module sram_compiled_array(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,din0,din1,din2,din3,din4,din5,din6,din7,din8,din9,din10,din11,din12,din13,din14,din15,din16,din17,din18,din19,din20,din21,din22,din23,din24,din25,din26,din27,din28,din29,din30,din31,dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7,dout8,dout9,dout10,dout11,dout12,dout13,dout14,dout15,dout16,dout17,dout18,dout19,dout20,dout21,dout22,dout23,dout24,dout25,dout26,dout27,dout28,dout29,dout30,dout31,clk,write_en,sense_en);
input addr0;
input addr1;
input addr2;
input addr3;
input addr4;
input addr5;
input addr6;
input addr7;
input din0;
input din1;
input din2;
input din3;
input din4;
input din5;
input din6;
input din7;
input din8;
input din9;
input din10;
input din11;
input din12;
input din13;
input din14;
input din15;
input din16;
input din17;
input din18;
input din19;
input din20;
input din21;
input din22;
input din23;
input din24;
input din25;
input din26;
input din27;
input din28;
input din29;
input din30;
input din31;
output dout0;
output dout1;
output dout2;
output dout3;
output dout4;
output dout5;
output dout6;
output dout7;
output dout8;
output dout9;
output dout10;
output dout11;
output dout12;
output dout13;
output dout14;
output dout15;
output dout16;
output dout17;
output dout18;
output dout19;
output dout20;
output dout21;
output dout22;
output dout23;
output dout24;
output dout25;
output dout26;
output dout27;
output dout28;
output dout29;
output dout30;
output dout31;
input clk;
input write_en;
input sense_en;
endmodule