// Verilog HDL and netlist files of
// "sram_compiled_20201119_153347_r64_c64_w8 sram_compiled_array schematic"
// Date Created : Apr 04 2021
// mrathore


// Netlisted models

// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell -
//colDecoder, View - schematic
// LAST TIME SAVED: Nov 19 15:34:19 2020
// NETLIST TIME: Apr  5 11:21:04 2021
`timescale 1ns / 1ps 

module colDecoder ( A0, A0_inv, A1, A1_inv, A2, A2_inv, CLK, YF0, YF1,
     YF2, YF3, YF4, YF5, YF6, YF7 );

output  YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7;

input  A0, A0_inv, A1, A1_inv, A2, A2_inv, CLK;


specify 
    specparam CDS_LIBNAME  =
     "sram_compiled_20201119_153347_r64_c64_w8";
    specparam CDS_CELLNAME = "colDecoder";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVC inst_clockedinv_b7_7 ( YF7, imd_YF7);
INVC inst_inv_b7_1_0 ( Y7, imd_Y7);
INVC inst_inv_b7_0_0 ( wire7_0_0, imd_wire7_0_0);
INVC inst_clockedinv_b6_6 ( YF6, imd_YF6);
INVC inst_inv_b6_1_0 ( Y6, imd_Y6);
INVC inst_inv_b6_0_0 ( wire6_0_0, imd_wire6_0_0);
INVC inst_clockedinv_b5_5 ( YF5, imd_YF5);
INVC inst_inv_b5_1_0 ( Y5, imd_Y5);
INVC inst_inv_b5_0_0 ( wire5_0_0, imd_wire5_0_0);
INVC inst_inv_b4_1_0 ( Y4, imd_Y4);
INVC inst_clockedinv_b4_4 ( YF4, imd_YF4);
INVC inst_inv_b4_0_0 ( wire4_0_0, imd_wire4_0_0);
INVC inst_clockedinv_b3_3 ( YF3, imd_YF3);
INVC inst_inv_b3_1_0 ( Y3, imd_Y3);
INVC inst_inv_b3_0_0 ( wire3_0_0, imd_wire3_0_0);
INVC inst_inv_b2_1_0 ( Y2, imd_Y2);
INVC inst_clockedinv_b2_2 ( YF2, imd_YF2);
INVC inst_inv_b2_0_0 ( wire2_0_0, imd_wire2_0_0);
INVC inst_inv_b1_1_0 ( Y1, imd_Y1);
INVC inst_clockedinv_b1_1 ( YF1, imd_YF1);
INVC inst_inv_b1_0_0 ( wire1_0_0, imd_wire1_0_0);
INVC inst_inv_b0_1_0 ( Y0, imd_Y0);
INVC inst_clockedinv_b0_0 ( YF0, imd_YF0);
INVC inst_inv_b0_0_0 ( wire0_0_0, imd_wire0_0_0);
NANDC2x1 inst_and_b7_1_0 ( imd_Y7, A2, wire7_0_0);
NANDC2x1 inst_and_b7_0_0 ( imd_wire7_0_0, A0, A1);
NANDC2x1 inst_clockedAND_b7_7 ( imd_YF7, CLK, Y7);
NANDC2x1 inst_and_b6_1_0 ( imd_Y6, A2, wire6_0_0);
NANDC2x1 inst_and_b6_0_0 ( imd_wire6_0_0, A0_inv, A1);
NANDC2x1 inst_clockedAND_b6_6 ( imd_YF6, CLK, Y6);
NANDC2x1 inst_and_b5_1_0 ( imd_Y5, A2, wire5_0_0);
NANDC2x1 inst_and_b5_0_0 ( imd_wire5_0_0, A0, A1_inv);
NANDC2x1 inst_clockedAND_b5_5 ( imd_YF5, CLK, Y5);
NANDC2x1 inst_clockedAND_b4_4 ( imd_YF4, CLK, Y4);
NANDC2x1 inst_and_b4_1_0 ( imd_Y4, A2, wire4_0_0);
NANDC2x1 inst_and_b4_0_0 ( imd_wire4_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b3_1_0 ( imd_Y3, A2_inv, wire3_0_0);
NANDC2x1 inst_and_b3_0_0 ( imd_wire3_0_0, A0, A1);
NANDC2x1 inst_clockedAND_b3_3 ( imd_YF3, CLK, Y3);
NANDC2x1 inst_and_b2_0_0 ( imd_wire2_0_0, A0_inv, A1);
NANDC2x1 inst_and_b2_1_0 ( imd_Y2, A2_inv, wire2_0_0);
NANDC2x1 inst_clockedAND_b2_2 ( imd_YF2, CLK, Y2);
NANDC2x1 inst_and_b1_0_0 ( imd_wire1_0_0, A0, A1_inv);
NANDC2x1 inst_and_b1_1_0 ( imd_Y1, A2_inv, wire1_0_0);
NANDC2x1 inst_clockedAND_b1_1 ( imd_YF1, CLK, Y1);
NANDC2x1 inst_and_b0_0_0 ( imd_wire0_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b0_1_0 ( imd_Y0, A2_inv, wire0_0_0);
NANDC2x1 inst_clockedAND_b0_0 ( imd_YF0, CLK, Y0);

endmodule
// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell - invCol,
//View - schematic
// LAST TIME SAVED: Nov 19 15:34:20 2020
// NETLIST TIME: Apr  5 11:21:04 2021
`timescale 1ns / 1ps 

module invCol ( A0, A1, A2, Abar0, Abar1, Abar2 );

output  Abar0, Abar1, Abar2;

input  A0, A1, A2;


specify 
    specparam CDS_LIBNAME  =
     "sram_compiled_20201119_153347_r64_c64_w8";
    specparam CDS_CELLNAME = "invCol";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVD wire2 ( Abar2, A2);
INVD wire1 ( Abar1, A1);
INVD wire0 ( Abar0, A0);

endmodule
// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell -
//columnMux, View - schematic
// LAST TIME SAVED: Nov 19 15:34:19 2020
// NETLIST TIME: Apr  5 11:21:04 2021
`timescale 1ns / 1ps 

module columnMux ( A0, Abar0, A1, Abar1, A2, Abar2, A3, Abar3, A4,
     Abar4, A5, Abar5, A6, Abar6, A7, Abar7, sel0, sel1, sel2, sel3,
     sel4, sel5, sel6, sel7, Y, Ybar );

output  Y, Ybar;

input  A0, A1, A2, A3, A4, A5, A6, A7, Abar0, Abar1, Abar2, Abar3,
     Abar4, Abar5, Abar6, Abar7, sel0, sel1, sel2, sel3, sel4, sel5,
     sel6, sel7;


specify 
    specparam CDS_LIBNAME  =
     "sram_compiled_20201119_153347_r64_c64_w8";
    specparam CDS_CELLNAME = "columnMux";
    specparam CDS_VIEWNAME = "schematic";
endspecify

muxTrans wire15 ( Abar7, Ybar, sel7);
muxTrans wire14 ( A7, Y, sel7);
muxTrans wire13 ( Abar6, Ybar, sel6);
muxTrans wire12 ( A6, Y, sel6);
muxTrans wire11 ( Abar5, Ybar, sel5);
muxTrans wire10 ( A5, Y, sel5);
muxTrans wire9 ( Abar4, Ybar, sel4);
muxTrans wire8 ( A4, Y, sel4);
muxTrans wire7 ( Abar3, Ybar, sel3);
muxTrans wire6 ( A3, Y, sel3);
muxTrans wire5 ( Abar2, Ybar, sel2);
muxTrans wire4 ( A2, Y, sel2);
muxTrans wire3 ( Abar1, Ybar, sel1);
muxTrans wire2 ( A1, Y, sel1);
muxTrans wire1 ( Abar0, Ybar, sel0);
muxTrans wire0 ( A0, Y, sel0);

endmodule
// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell - invRow,
//View - schematic
// LAST TIME SAVED: Nov 19 15:34:20 2020
// NETLIST TIME: Apr  5 11:21:04 2021
`timescale 1ns / 1ps 

module invRow ( A0, A1, A2, A3, A4, A5, Abar0, Abar1, Abar2, Abar3,
     Abar4, Abar5 );

output  Abar0, Abar1, Abar2, Abar3, Abar4, Abar5;

input  A0, A1, A2, A3, A4, A5;


specify 
    specparam CDS_LIBNAME  =
     "sram_compiled_20201119_153347_r64_c64_w8";
    specparam CDS_CELLNAME = "invRow";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVD wire5 ( Abar5, A5);
INVD wire4 ( Abar4, A4);
INVD wire3 ( Abar3, A3);
INVD wire2 ( Abar2, A2);
INVD wire1 ( Abar1, A1);
INVD wire0 ( Abar0, A0);

endmodule
// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell -
//rowDecoder, View - schematic
// LAST TIME SAVED: Nov 19 15:34:20 2020
// NETLIST TIME: Apr  5 11:21:04 2021
`timescale 1ns / 1ps 

module rowDecoder ( A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv, A4,
     A4_inv, A5, A5_inv, CLK, YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7,
     YF8, YF9, YF10, YF11, YF12, YF13, YF14, YF15, YF16, YF17, YF18,
     YF19, YF20, YF21, YF22, YF23, YF24, YF25, YF26, YF27, YF28, YF29,
     YF30, YF31, YF32, YF33, YF34, YF35, YF36, YF37, YF38, YF39, YF40,
     YF41, YF42, YF43, YF44, YF45, YF46, YF47, YF48, YF49, YF50, YF51,
     YF52, YF53, YF54, YF55, YF56, YF57, YF58, YF59, YF60, YF61, YF62,
     YF63 );

output  YF0, YF1, YF2, YF3, YF4, YF5, YF6, YF7, YF8, YF9, YF10, YF11,
     YF12, YF13, YF14, YF15, YF16, YF17, YF18, YF19, YF20, YF21, YF22,
     YF23, YF24, YF25, YF26, YF27, YF28, YF29, YF30, YF31, YF32, YF33,
     YF34, YF35, YF36, YF37, YF38, YF39, YF40, YF41, YF42, YF43, YF44,
     YF45, YF46, YF47, YF48, YF49, YF50, YF51, YF52, YF53, YF54, YF55,
     YF56, YF57, YF58, YF59, YF60, YF61, YF62, YF63;

input  A0, A0_inv, A1, A1_inv, A2, A2_inv, A3, A3_inv, A4, A4_inv, A5,
     A5_inv, CLK;


specify 
    specparam CDS_LIBNAME  =
     "sram_compiled_20201119_153347_r64_c64_w8";
    specparam CDS_CELLNAME = "rowDecoder";
    specparam CDS_VIEWNAME = "schematic";
endspecify

NANDC2x1 inst_clockedAND_b63_63 ( imd_YF63, CLK, Y63);
NANDC2x1 inst_and_b63_0_2 ( imd_wire63_0_2, A4, A5);
NANDC2x1 inst_and_b63_2_0 ( imd_Y63, wire63_0_2, wire63_1_0);
NANDC2x1 inst_and_b63_0_1 ( imd_wire63_0_1, A2, A3);
NANDC2x1 inst_and_b63_0_0 ( imd_wire63_0_0, A0, A1);
NANDC2x1 inst_and_b63_1_0 ( imd_wire63_1_0, wire63_0_0, wire63_0_1);
NANDC2x1 inst_clockedAND_b62_62 ( imd_YF62, CLK, Y62);
NANDC2x1 inst_and_b62_0_2 ( imd_wire62_0_2, A4, A5);
NANDC2x1 inst_and_b62_2_0 ( imd_Y62, wire62_0_2, wire62_1_0);
NANDC2x1 inst_and_b62_0_1 ( imd_wire62_0_1, A2, A3);
NANDC2x1 inst_and_b62_0_0 ( imd_wire62_0_0, A0_inv, A1);
NANDC2x1 inst_and_b62_1_0 ( imd_wire62_1_0, wire62_0_0, wire62_0_1);
NANDC2x1 inst_clockedAND_b61_61 ( imd_YF61, CLK, Y61);
NANDC2x1 inst_and_b61_0_2 ( imd_wire61_0_2, A4, A5);
NANDC2x1 inst_and_b61_2_0 ( imd_Y61, wire61_0_2, wire61_1_0);
NANDC2x1 inst_and_b61_0_1 ( imd_wire61_0_1, A2, A3);
NANDC2x1 inst_and_b61_0_0 ( imd_wire61_0_0, A0, A1_inv);
NANDC2x1 inst_and_b61_1_0 ( imd_wire61_1_0, wire61_0_0, wire61_0_1);
NANDC2x1 inst_clockedAND_b60_60 ( imd_YF60, CLK, Y60);
NANDC2x1 inst_and_b60_0_2 ( imd_wire60_0_2, A4, A5);
NANDC2x1 inst_and_b60_2_0 ( imd_Y60, wire60_0_2, wire60_1_0);
NANDC2x1 inst_and_b60_0_1 ( imd_wire60_0_1, A2, A3);
NANDC2x1 inst_and_b60_0_0 ( imd_wire60_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b60_1_0 ( imd_wire60_1_0, wire60_0_0, wire60_0_1);
NANDC2x1 inst_clockedAND_b59_59 ( imd_YF59, CLK, Y59);
NANDC2x1 inst_and_b59_0_2 ( imd_wire59_0_2, A4, A5);
NANDC2x1 inst_and_b59_2_0 ( imd_Y59, wire59_0_2, wire59_1_0);
NANDC2x1 inst_and_b59_0_1 ( imd_wire59_0_1, A2_inv, A3);
NANDC2x1 inst_and_b59_0_0 ( imd_wire59_0_0, A0, A1);
NANDC2x1 inst_and_b59_1_0 ( imd_wire59_1_0, wire59_0_0, wire59_0_1);
NANDC2x1 inst_clockedAND_b58_58 ( imd_YF58, CLK, Y58);
NANDC2x1 inst_and_b58_0_2 ( imd_wire58_0_2, A4, A5);
NANDC2x1 inst_and_b58_2_0 ( imd_Y58, wire58_0_2, wire58_1_0);
NANDC2x1 inst_and_b58_0_1 ( imd_wire58_0_1, A2_inv, A3);
NANDC2x1 inst_and_b58_0_0 ( imd_wire58_0_0, A0_inv, A1);
NANDC2x1 inst_and_b58_1_0 ( imd_wire58_1_0, wire58_0_0, wire58_0_1);
NANDC2x1 inst_clockedAND_b57_57 ( imd_YF57, CLK, Y57);
NANDC2x1 inst_and_b57_0_2 ( imd_wire57_0_2, A4, A5);
NANDC2x1 inst_and_b57_2_0 ( imd_Y57, wire57_0_2, wire57_1_0);
NANDC2x1 inst_and_b57_0_1 ( imd_wire57_0_1, A2_inv, A3);
NANDC2x1 inst_and_b57_0_0 ( imd_wire57_0_0, A0, A1_inv);
NANDC2x1 inst_and_b57_1_0 ( imd_wire57_1_0, wire57_0_0, wire57_0_1);
NANDC2x1 inst_clockedAND_b56_56 ( imd_YF56, CLK, Y56);
NANDC2x1 inst_and_b56_0_2 ( imd_wire56_0_2, A4, A5);
NANDC2x1 inst_and_b56_2_0 ( imd_Y56, wire56_0_2, wire56_1_0);
NANDC2x1 inst_and_b56_0_1 ( imd_wire56_0_1, A2_inv, A3);
NANDC2x1 inst_and_b56_0_0 ( imd_wire56_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b56_1_0 ( imd_wire56_1_0, wire56_0_0, wire56_0_1);
NANDC2x1 inst_clockedAND_b55_55 ( imd_YF55, CLK, Y55);
NANDC2x1 inst_and_b55_0_2 ( imd_wire55_0_2, A4, A5);
NANDC2x1 inst_and_b55_2_0 ( imd_Y55, wire55_0_2, wire55_1_0);
NANDC2x1 inst_and_b55_0_1 ( imd_wire55_0_1, A2, A3_inv);
NANDC2x1 inst_and_b54_0_1 ( imd_wire54_0_1, A2, A3_inv);
NANDC2x1 inst_and_b55_0_0 ( imd_wire55_0_0, A0, A1);
NANDC2x1 inst_and_b55_1_0 ( imd_wire55_1_0, wire55_0_0, wire55_0_1);
NANDC2x1 inst_clockedAND_b54_54 ( imd_YF54, CLK, Y54);
NANDC2x1 inst_and_b54_1_0 ( imd_wire54_1_0, wire54_0_0, wire54_0_1);
NANDC2x1 inst_and_b54_0_0 ( imd_wire54_0_0, A0_inv, A1);
NANDC2x1 inst_and_b54_0_2 ( imd_wire54_0_2, A4, A5);
NANDC2x1 inst_and_b54_2_0 ( imd_Y54, wire54_0_2, wire54_1_0);
NANDC2x1 inst_clockedAND_b53_53 ( imd_YF53, CLK, Y53);
NANDC2x1 inst_and_b53_0_2 ( imd_wire53_0_2, A4, A5);
NANDC2x1 inst_and_b53_2_0 ( imd_Y53, wire53_0_2, wire53_1_0);
NANDC2x1 inst_clockedAND_b52_52 ( imd_YF52, CLK, Y52);
NANDC2x1 inst_and_b52_0_2 ( imd_wire52_0_2, A4, A5);
NANDC2x1 inst_and_b52_2_0 ( imd_Y52, wire52_0_2, wire52_1_0);
NANDC2x1 inst_and_b52_0_1 ( imd_wire52_0_1, A2, A3_inv);
NANDC2x1 inst_and_b52_0_0 ( imd_wire52_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b52_1_0 ( imd_wire52_1_0, wire52_0_0, wire52_0_1);
NANDC2x1 inst_clockedAND_b51_51 ( imd_YF51, CLK, Y51);
NANDC2x1 inst_and_b51_0_2 ( imd_wire51_0_2, A4, A5);
NANDC2x1 inst_and_b51_2_0 ( imd_Y51, wire51_0_2, wire51_1_0);
NANDC2x1 inst_and_b51_0_1 ( imd_wire51_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b51_0_0 ( imd_wire51_0_0, A0, A1);
NANDC2x1 inst_and_b51_1_0 ( imd_wire51_1_0, wire51_0_0, wire51_0_1);
NANDC2x1 inst_clockedAND_b50_50 ( imd_YF50, CLK, Y50);
NANDC2x1 inst_and_b50_0_2 ( imd_wire50_0_2, A4, A5);
NANDC2x1 inst_and_b50_2_0 ( imd_Y50, wire50_0_2, wire50_1_0);
NANDC2x1 inst_and_b50_0_1 ( imd_wire50_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b50_0_0 ( imd_wire50_0_0, A0_inv, A1);
NANDC2x1 inst_and_b50_1_0 ( imd_wire50_1_0, wire50_0_0, wire50_0_1);
NANDC2x1 inst_clockedAND_b49_49 ( imd_YF49, CLK, Y49);
NANDC2x1 inst_and_b49_0_2 ( imd_wire49_0_2, A4, A5);
NANDC2x1 inst_and_b49_2_0 ( imd_Y49, wire49_0_2, wire49_1_0);
NANDC2x1 inst_and_b49_0_1 ( imd_wire49_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b49_0_0 ( imd_wire49_0_0, A0, A1_inv);
NANDC2x1 inst_and_b49_1_0 ( imd_wire49_1_0, wire49_0_0, wire49_0_1);
NANDC2x1 inst_clockedAND_b48_48 ( imd_YF48, CLK, Y48);
NANDC2x1 inst_and_b48_0_2 ( imd_wire48_0_2, A4, A5);
NANDC2x1 inst_and_b48_2_0 ( imd_Y48, wire48_0_2, wire48_1_0);
NANDC2x1 inst_and_b48_0_1 ( imd_wire48_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b48_0_0 ( imd_wire48_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b48_1_0 ( imd_wire48_1_0, wire48_0_0, wire48_0_1);
NANDC2x1 inst_clockedAND_b47_47 ( imd_YF47, CLK, Y47);
NANDC2x1 inst_and_b47_0_2 ( imd_wire47_0_2, A4_inv, A5);
NANDC2x1 inst_and_b47_2_0 ( imd_Y47, wire47_0_2, wire47_1_0);
NANDC2x1 inst_and_b47_0_1 ( imd_wire47_0_1, A2, A3);
NANDC2x1 inst_and_b47_0_0 ( imd_wire47_0_0, A0, A1);
NANDC2x1 inst_and_b47_1_0 ( imd_wire47_1_0, wire47_0_0, wire47_0_1);
NANDC2x1 inst_clockedAND_b46_46 ( imd_YF46, CLK, Y46);
NANDC2x1 inst_and_b46_0_2 ( imd_wire46_0_2, A4_inv, A5);
NANDC2x1 inst_and_b46_2_0 ( imd_Y46, wire46_0_2, wire46_1_0);
NANDC2x1 inst_and_b46_0_1 ( imd_wire46_0_1, A2, A3);
NANDC2x1 inst_and_b46_0_0 ( imd_wire46_0_0, A0_inv, A1);
NANDC2x1 inst_and_b46_1_0 ( imd_wire46_1_0, wire46_0_0, wire46_0_1);
NANDC2x1 inst_clockedAND_b45_45 ( imd_YF45, CLK, Y45);
NANDC2x1 inst_and_b45_0_2 ( imd_wire45_0_2, A4_inv, A5);
NANDC2x1 inst_and_b45_2_0 ( imd_Y45, wire45_0_2, wire45_1_0);
NANDC2x1 inst_and_b45_0_1 ( imd_wire45_0_1, A2, A3);
NANDC2x1 inst_and_b45_0_0 ( imd_wire45_0_0, A0, A1_inv);
NANDC2x1 inst_and_b45_1_0 ( imd_wire45_1_0, wire45_0_0, wire45_0_1);
NANDC2x1 inst_clockedAND_b44_44 ( imd_YF44, CLK, Y44);
NANDC2x1 inst_and_b44_0_2 ( imd_wire44_0_2, A4_inv, A5);
NANDC2x1 inst_and_b44_2_0 ( imd_Y44, wire44_0_2, wire44_1_0);
NANDC2x1 inst_and_b44_0_1 ( imd_wire44_0_1, A2, A3);
NANDC2x1 inst_and_b44_0_0 ( imd_wire44_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b44_1_0 ( imd_wire44_1_0, wire44_0_0, wire44_0_1);
NANDC2x1 inst_clockedAND_b43_43 ( imd_YF43, CLK, Y43);
NANDC2x1 inst_and_b43_0_2 ( imd_wire43_0_2, A4_inv, A5);
NANDC2x1 inst_and_b43_2_0 ( imd_Y43, wire43_0_2, wire43_1_0);
NANDC2x1 inst_and_b43_0_1 ( imd_wire43_0_1, A2_inv, A3);
NANDC2x1 inst_and_b43_0_0 ( imd_wire43_0_0, A0, A1);
NANDC2x1 inst_and_b43_1_0 ( imd_wire43_1_0, wire43_0_0, wire43_0_1);
NANDC2x1 inst_and_b53_1_0 ( imd_wire53_1_0, wire53_0_0, wire53_0_1);
NANDC2x1 inst_and_b53_0_0 ( imd_wire53_0_0, A0, A1_inv);
NANDC2x1 inst_and_b53_0_1 ( imd_wire53_0_1, A2, A3_inv);
NANDC2x1 inst_clockedAND_b42_42 ( imd_YF42, CLK, Y42);
NANDC2x1 inst_and_b42_2_0 ( imd_Y42, wire42_0_2, wire42_1_0);
NANDC2x1 inst_and_b42_0_2 ( imd_wire42_0_2, A4_inv, A5);
NANDC2x1 inst_and_b42_0_1 ( imd_wire42_0_1, A2_inv, A3);
NANDC2x1 inst_and_b42_0_0 ( imd_wire42_0_0, A0_inv, A1);
NANDC2x1 inst_and_b42_1_0 ( imd_wire42_1_0, wire42_0_0, wire42_0_1);
NANDC2x1 inst_clockedAND_b41_41 ( imd_YF41, CLK, Y41);
NANDC2x1 inst_and_b41_0_2 ( imd_wire41_0_2, A4_inv, A5);
NANDC2x1 inst_and_b41_2_0 ( imd_Y41, wire41_0_2, wire41_1_0);
NANDC2x1 inst_and_b41_0_1 ( imd_wire41_0_1, A2_inv, A3);
NANDC2x1 inst_and_b41_0_0 ( imd_wire41_0_0, A0, A1_inv);
NANDC2x1 inst_and_b41_1_0 ( imd_wire41_1_0, wire41_0_0, wire41_0_1);
NANDC2x1 inst_clockedAND_b40_40 ( imd_YF40, CLK, Y40);
NANDC2x1 inst_and_b40_0_2 ( imd_wire40_0_2, A4_inv, A5);
NANDC2x1 inst_and_b40_2_0 ( imd_Y40, wire40_0_2, wire40_1_0);
NANDC2x1 inst_and_b40_0_1 ( imd_wire40_0_1, A2_inv, A3);
NANDC2x1 inst_and_b40_0_0 ( imd_wire40_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b40_1_0 ( imd_wire40_1_0, wire40_0_0, wire40_0_1);
NANDC2x1 inst_clockedAND_b39_39 ( imd_YF39, CLK, Y39);
NANDC2x1 inst_and_b39_0_2 ( imd_wire39_0_2, A4_inv, A5);
NANDC2x1 inst_and_b39_2_0 ( imd_Y39, wire39_0_2, wire39_1_0);
NANDC2x1 inst_and_b39_0_1 ( imd_wire39_0_1, A2, A3_inv);
NANDC2x1 inst_and_b39_0_0 ( imd_wire39_0_0, A0, A1);
NANDC2x1 inst_and_b39_1_0 ( imd_wire39_1_0, wire39_0_0, wire39_0_1);
NANDC2x1 inst_clockedAND_b38_38 ( imd_YF38, CLK, Y38);
NANDC2x1 inst_and_b38_0_2 ( imd_wire38_0_2, A4_inv, A5);
NANDC2x1 inst_and_b38_2_0 ( imd_Y38, wire38_0_2, wire38_1_0);
NANDC2x1 inst_and_b38_0_1 ( imd_wire38_0_1, A2, A3_inv);
NANDC2x1 inst_and_b38_0_0 ( imd_wire38_0_0, A0_inv, A1);
NANDC2x1 inst_and_b38_1_0 ( imd_wire38_1_0, wire38_0_0, wire38_0_1);
NANDC2x1 inst_clockedAND_b37_37 ( imd_YF37, CLK, Y37);
NANDC2x1 inst_and_b37_0_2 ( imd_wire37_0_2, A4_inv, A5);
NANDC2x1 inst_and_b37_2_0 ( imd_Y37, wire37_0_2, wire37_1_0);
NANDC2x1 inst_and_b37_0_1 ( imd_wire37_0_1, A2, A3_inv);
NANDC2x1 inst_and_b37_0_0 ( imd_wire37_0_0, A0, A1_inv);
NANDC2x1 inst_and_b37_1_0 ( imd_wire37_1_0, wire37_0_0, wire37_0_1);
NANDC2x1 inst_clockedAND_b36_36 ( imd_YF36, CLK, Y36);
NANDC2x1 inst_and_b36_0_2 ( imd_wire36_0_2, A4_inv, A5);
NANDC2x1 inst_and_b36_2_0 ( imd_Y36, wire36_0_2, wire36_1_0);
NANDC2x1 inst_and_b36_0_1 ( imd_wire36_0_1, A2, A3_inv);
NANDC2x1 inst_and_b36_0_0 ( imd_wire36_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b36_1_0 ( imd_wire36_1_0, wire36_0_0, wire36_0_1);
NANDC2x1 inst_clockedAND_b35_35 ( imd_YF35, CLK, Y35);
NANDC2x1 inst_and_b35_0_2 ( imd_wire35_0_2, A4_inv, A5);
NANDC2x1 inst_and_b35_2_0 ( imd_Y35, wire35_0_2, wire35_1_0);
NANDC2x1 inst_and_b35_0_1 ( imd_wire35_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b35_0_0 ( imd_wire35_0_0, A0, A1);
NANDC2x1 inst_and_b35_1_0 ( imd_wire35_1_0, wire35_0_0, wire35_0_1);
NANDC2x1 inst_clockedAND_b34_34 ( imd_YF34, CLK, Y34);
NANDC2x1 inst_and_b34_0_2 ( imd_wire34_0_2, A4_inv, A5);
NANDC2x1 inst_and_b34_2_0 ( imd_Y34, wire34_0_2, wire34_1_0);
NANDC2x1 inst_and_b34_0_1 ( imd_wire34_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b34_0_0 ( imd_wire34_0_0, A0_inv, A1);
NANDC2x1 inst_and_b34_1_0 ( imd_wire34_1_0, wire34_0_0, wire34_0_1);
NANDC2x1 inst_clockedAND_b33_33 ( imd_YF33, CLK, Y33);
NANDC2x1 inst_and_b33_0_2 ( imd_wire33_0_2, A4_inv, A5);
NANDC2x1 inst_and_b33_2_0 ( imd_Y33, wire33_0_2, wire33_1_0);
NANDC2x1 inst_and_b33_0_1 ( imd_wire33_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b33_0_0 ( imd_wire33_0_0, A0, A1_inv);
NANDC2x1 inst_and_b33_1_0 ( imd_wire33_1_0, wire33_0_0, wire33_0_1);
NANDC2x1 inst_and_b32_0_2 ( imd_wire32_0_2, A4_inv, A5);
NANDC2x1 inst_clockedAND_b32_32 ( imd_YF32, CLK, Y32);
NANDC2x1 inst_and_b32_2_0 ( imd_Y32, wire32_0_2, wire32_1_0);
NANDC2x1 inst_and_b32_0_1 ( imd_wire32_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b32_0_0 ( imd_wire32_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b32_1_0 ( imd_wire32_1_0, wire32_0_0, wire32_0_1);
NANDC2x1 inst_clockedAND_b31_31 ( imd_YF31, CLK, Y31);
NANDC2x1 inst_and_b31_0_2 ( imd_wire31_0_2, A4, A5_inv);
NANDC2x1 inst_and_b31_2_0 ( imd_Y31, wire31_0_2, wire31_1_0);
NANDC2x1 inst_and_b31_0_1 ( imd_wire31_0_1, A2, A3);
NANDC2x1 inst_and_b31_0_0 ( imd_wire31_0_0, A0, A1);
NANDC2x1 inst_and_b31_1_0 ( imd_wire31_1_0, wire31_0_0, wire31_0_1);
NANDC2x1 inst_clockedAND_b30_30 ( imd_YF30, CLK, Y30);
NANDC2x1 inst_and_b30_0_2 ( imd_wire30_0_2, A4, A5_inv);
NANDC2x1 inst_and_b30_2_0 ( imd_Y30, wire30_0_2, wire30_1_0);
NANDC2x1 inst_and_b30_0_1 ( imd_wire30_0_1, A2, A3);
NANDC2x1 inst_and_b30_0_0 ( imd_wire30_0_0, A0_inv, A1);
NANDC2x1 inst_and_b30_1_0 ( imd_wire30_1_0, wire30_0_0, wire30_0_1);
NANDC2x1 inst_clockedAND_b29_29 ( imd_YF29, CLK, Y29);
NANDC2x1 inst_and_b29_0_2 ( imd_wire29_0_2, A4, A5_inv);
NANDC2x1 inst_and_b29_2_0 ( imd_Y29, wire29_0_2, wire29_1_0);
NANDC2x1 inst_and_b29_0_1 ( imd_wire29_0_1, A2, A3);
NANDC2x1 inst_and_b29_0_0 ( imd_wire29_0_0, A0, A1_inv);
NANDC2x1 inst_and_b29_1_0 ( imd_wire29_1_0, wire29_0_0, wire29_0_1);
NANDC2x1 inst_clockedAND_b28_28 ( imd_YF28, CLK, Y28);
NANDC2x1 inst_and_b28_0_2 ( imd_wire28_0_2, A4, A5_inv);
NANDC2x1 inst_and_b28_2_0 ( imd_Y28, wire28_0_2, wire28_1_0);
NANDC2x1 inst_and_b28_0_1 ( imd_wire28_0_1, A2, A3);
NANDC2x1 inst_and_b28_0_0 ( imd_wire28_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b28_1_0 ( imd_wire28_1_0, wire28_0_0, wire28_0_1);
NANDC2x1 inst_clockedAND_b27_27 ( imd_YF27, CLK, Y27);
NANDC2x1 inst_and_b27_0_2 ( imd_wire27_0_2, A4, A5_inv);
NANDC2x1 inst_and_b27_2_0 ( imd_Y27, wire27_0_2, wire27_1_0);
NANDC2x1 inst_and_b27_0_1 ( imd_wire27_0_1, A2_inv, A3);
NANDC2x1 inst_and_b27_0_0 ( imd_wire27_0_0, A0, A1);
NANDC2x1 inst_and_b27_1_0 ( imd_wire27_1_0, wire27_0_0, wire27_0_1);
NANDC2x1 inst_clockedAND_b26_26 ( imd_YF26, CLK, Y26);
NANDC2x1 inst_and_b26_0_2 ( imd_wire26_0_2, A4, A5_inv);
NANDC2x1 inst_and_b26_2_0 ( imd_Y26, wire26_0_2, wire26_1_0);
NANDC2x1 inst_and_b26_0_1 ( imd_wire26_0_1, A2_inv, A3);
NANDC2x1 inst_and_b26_0_0 ( imd_wire26_0_0, A0_inv, A1);
NANDC2x1 inst_and_b26_1_0 ( imd_wire26_1_0, wire26_0_0, wire26_0_1);
NANDC2x1 inst_clockedAND_b25_25 ( imd_YF25, CLK, Y25);
NANDC2x1 inst_and_b25_0_2 ( imd_wire25_0_2, A4, A5_inv);
NANDC2x1 inst_and_b25_2_0 ( imd_Y25, wire25_0_2, wire25_1_0);
NANDC2x1 inst_and_b25_0_1 ( imd_wire25_0_1, A2_inv, A3);
NANDC2x1 inst_and_b25_0_0 ( imd_wire25_0_0, A0, A1_inv);
NANDC2x1 inst_and_b25_1_0 ( imd_wire25_1_0, wire25_0_0, wire25_0_1);
NANDC2x1 inst_clockedAND_b24_24 ( imd_YF24, CLK, Y24);
NANDC2x1 inst_and_b24_0_2 ( imd_wire24_0_2, A4, A5_inv);
NANDC2x1 inst_and_b24_2_0 ( imd_Y24, wire24_0_2, wire24_1_0);
NANDC2x1 inst_and_b24_0_1 ( imd_wire24_0_1, A2_inv, A3);
NANDC2x1 inst_and_b24_0_0 ( imd_wire24_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b24_1_0 ( imd_wire24_1_0, wire24_0_0, wire24_0_1);
NANDC2x1 inst_clockedAND_b23_23 ( imd_YF23, CLK, Y23);
NANDC2x1 inst_and_b23_0_2 ( imd_wire23_0_2, A4, A5_inv);
NANDC2x1 inst_and_b23_2_0 ( imd_Y23, wire23_0_2, wire23_1_0);
NANDC2x1 inst_and_b23_0_1 ( imd_wire23_0_1, A2, A3_inv);
NANDC2x1 inst_and_b22_0_1 ( imd_wire22_0_1, A2, A3_inv);
NANDC2x1 inst_and_b23_0_0 ( imd_wire23_0_0, A0, A1);
NANDC2x1 inst_and_b23_1_0 ( imd_wire23_1_0, wire23_0_0, wire23_0_1);
NANDC2x1 inst_clockedAND_b22_22 ( imd_YF22, CLK, Y22);
NANDC2x1 inst_and_b22_1_0 ( imd_wire22_1_0, wire22_0_0, wire22_0_1);
NANDC2x1 inst_and_b22_0_0 ( imd_wire22_0_0, A0_inv, A1);
NANDC2x1 inst_and_b22_0_2 ( imd_wire22_0_2, A4, A5_inv);
NANDC2x1 inst_and_b22_2_0 ( imd_Y22, wire22_0_2, wire22_1_0);
NANDC2x1 inst_clockedAND_b21_21 ( imd_YF21, CLK, Y21);
NANDC2x1 inst_and_b21_0_2 ( imd_wire21_0_2, A4, A5_inv);
NANDC2x1 inst_and_b21_2_0 ( imd_Y21, wire21_0_2, wire21_1_0);
NANDC2x1 inst_clockedAND_b20_20 ( imd_YF20, CLK, Y20);
NANDC2x1 inst_and_b20_0_2 ( imd_wire20_0_2, A4, A5_inv);
NANDC2x1 inst_and_b20_2_0 ( imd_Y20, wire20_0_2, wire20_1_0);
NANDC2x1 inst_and_b20_0_1 ( imd_wire20_0_1, A2, A3_inv);
NANDC2x1 inst_and_b20_0_0 ( imd_wire20_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b20_1_0 ( imd_wire20_1_0, wire20_0_0, wire20_0_1);
NANDC2x1 inst_clockedAND_b19_19 ( imd_YF19, CLK, Y19);
NANDC2x1 inst_and_b19_0_2 ( imd_wire19_0_2, A4, A5_inv);
NANDC2x1 inst_and_b19_2_0 ( imd_Y19, wire19_0_2, wire19_1_0);
NANDC2x1 inst_and_b19_0_1 ( imd_wire19_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b19_0_0 ( imd_wire19_0_0, A0, A1);
NANDC2x1 inst_and_b19_1_0 ( imd_wire19_1_0, wire19_0_0, wire19_0_1);
NANDC2x1 inst_clockedAND_b18_18 ( imd_YF18, CLK, Y18);
NANDC2x1 inst_and_b18_0_2 ( imd_wire18_0_2, A4, A5_inv);
NANDC2x1 inst_and_b18_2_0 ( imd_Y18, wire18_0_2, wire18_1_0);
NANDC2x1 inst_and_b18_0_1 ( imd_wire18_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b18_0_0 ( imd_wire18_0_0, A0_inv, A1);
NANDC2x1 inst_and_b18_1_0 ( imd_wire18_1_0, wire18_0_0, wire18_0_1);
NANDC2x1 inst_clockedAND_b17_17 ( imd_YF17, CLK, Y17);
NANDC2x1 inst_and_b17_0_2 ( imd_wire17_0_2, A4, A5_inv);
NANDC2x1 inst_and_b17_2_0 ( imd_Y17, wire17_0_2, wire17_1_0);
NANDC2x1 inst_and_b17_0_1 ( imd_wire17_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b17_0_0 ( imd_wire17_0_0, A0, A1_inv);
NANDC2x1 inst_and_b17_1_0 ( imd_wire17_1_0, wire17_0_0, wire17_0_1);
NANDC2x1 inst_and_b16_0_2 ( imd_wire16_0_2, A4, A5_inv);
NANDC2x1 inst_clockedAND_b16_16 ( imd_YF16, CLK, Y16);
NANDC2x1 inst_and_b16_2_0 ( imd_Y16, wire16_0_2, wire16_1_0);
NANDC2x1 inst_and_b16_0_1 ( imd_wire16_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b16_0_0 ( imd_wire16_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b16_1_0 ( imd_wire16_1_0, wire16_0_0, wire16_0_1);
NANDC2x1 inst_clockedAND_b15_15 ( imd_YF15, CLK, Y15);
NANDC2x1 inst_and_b15_0_2 ( imd_wire15_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b15_2_0 ( imd_Y15, wire15_0_2, wire15_1_0);
NANDC2x1 inst_and_b15_0_1 ( imd_wire15_0_1, A2, A3);
NANDC2x1 inst_and_b15_0_0 ( imd_wire15_0_0, A0, A1);
NANDC2x1 inst_and_b15_1_0 ( imd_wire15_1_0, wire15_0_0, wire15_0_1);
NANDC2x1 inst_clockedAND_b14_14 ( imd_YF14, CLK, Y14);
NANDC2x1 inst_and_b14_0_2 ( imd_wire14_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b14_2_0 ( imd_Y14, wire14_0_2, wire14_1_0);
NANDC2x1 inst_and_b14_0_1 ( imd_wire14_0_1, A2, A3);
NANDC2x1 inst_and_b14_0_0 ( imd_wire14_0_0, A0_inv, A1);
NANDC2x1 inst_and_b14_1_0 ( imd_wire14_1_0, wire14_0_0, wire14_0_1);
NANDC2x1 inst_clockedAND_b13_13 ( imd_YF13, CLK, Y13);
NANDC2x1 inst_and_b13_0_2 ( imd_wire13_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b13_2_0 ( imd_Y13, wire13_0_2, wire13_1_0);
NANDC2x1 inst_and_b13_0_1 ( imd_wire13_0_1, A2, A3);
NANDC2x1 inst_and_b13_0_0 ( imd_wire13_0_0, A0, A1_inv);
NANDC2x1 inst_and_b13_1_0 ( imd_wire13_1_0, wire13_0_0, wire13_0_1);
NANDC2x1 inst_clockedAND_b12_12 ( imd_YF12, CLK, Y12);
NANDC2x1 inst_and_b12_0_2 ( imd_wire12_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b12_2_0 ( imd_Y12, wire12_0_2, wire12_1_0);
NANDC2x1 inst_and_b12_0_1 ( imd_wire12_0_1, A2, A3);
NANDC2x1 inst_and_b12_0_0 ( imd_wire12_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b12_1_0 ( imd_wire12_1_0, wire12_0_0, wire12_0_1);
NANDC2x1 inst_clockedAND_b11_11 ( imd_YF11, CLK, Y11);
NANDC2x1 inst_and_b11_0_2 ( imd_wire11_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b11_2_0 ( imd_Y11, wire11_0_2, wire11_1_0);
NANDC2x1 inst_and_b11_0_1 ( imd_wire11_0_1, A2_inv, A3);
NANDC2x1 inst_and_b11_0_0 ( imd_wire11_0_0, A0, A1);
NANDC2x1 inst_and_b11_1_0 ( imd_wire11_1_0, wire11_0_0, wire11_0_1);
NANDC2x1 inst_and_b21_1_0 ( imd_wire21_1_0, wire21_0_0, wire21_0_1);
NANDC2x1 inst_and_b21_0_0 ( imd_wire21_0_0, A0, A1_inv);
NANDC2x1 inst_and_b21_0_1 ( imd_wire21_0_1, A2, A3_inv);
NANDC2x1 inst_clockedAND_b10_10 ( imd_YF10, CLK, Y10);
NANDC2x1 inst_and_b10_2_0 ( imd_Y10, wire10_0_2, wire10_1_0);
NANDC2x1 inst_and_b10_0_2 ( imd_wire10_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b10_0_1 ( imd_wire10_0_1, A2_inv, A3);
NANDC2x1 inst_and_b10_0_0 ( imd_wire10_0_0, A0_inv, A1);
NANDC2x1 inst_and_b10_1_0 ( imd_wire10_1_0, wire10_0_0, wire10_0_1);
NANDC2x1 inst_clockedAND_b9_9 ( imd_YF9, CLK, Y9);
NANDC2x1 inst_and_b9_0_2 ( imd_wire9_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b9_2_0 ( imd_Y9, wire9_0_2, wire9_1_0);
NANDC2x1 inst_and_b9_0_1 ( imd_wire9_0_1, A2_inv, A3);
NANDC2x1 inst_and_b9_0_0 ( imd_wire9_0_0, A0, A1_inv);
NANDC2x1 inst_and_b9_1_0 ( imd_wire9_1_0, wire9_0_0, wire9_0_1);
NANDC2x1 inst_and_b8_0_1 ( imd_wire8_0_1, A2_inv, A3);
NANDC2x1 inst_and_b8_0_0 ( imd_wire8_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b8_1_0 ( imd_wire8_1_0, wire8_0_0, wire8_0_1);
NANDC2x1 inst_clockedAND_b8_8 ( imd_YF8, CLK, Y8);
NANDC2x1 inst_and_b8_0_2 ( imd_wire8_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b8_2_0 ( imd_Y8, wire8_0_2, wire8_1_0);
NANDC2x1 inst_clockedAND_b7_7 ( imd_YF7, CLK, Y7);
NANDC2x1 inst_and_b7_0_2 ( imd_wire7_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b7_2_0 ( imd_Y7, wire7_0_2, wire7_1_0);
NANDC2x1 inst_and_b7_0_1 ( imd_wire7_0_1, A2, A3_inv);
NANDC2x1 inst_and_b7_0_0 ( imd_wire7_0_0, A0, A1);
NANDC2x1 inst_and_b7_1_0 ( imd_wire7_1_0, wire7_0_0, wire7_0_1);
NANDC2x1 inst_clockedAND_b6_6 ( imd_YF6, CLK, Y6);
NANDC2x1 inst_and_b6_0_2 ( imd_wire6_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b6_2_0 ( imd_Y6, wire6_0_2, wire6_1_0);
NANDC2x1 inst_and_b6_0_1 ( imd_wire6_0_1, A2, A3_inv);
NANDC2x1 inst_and_b6_0_0 ( imd_wire6_0_0, A0_inv, A1);
NANDC2x1 inst_and_b6_1_0 ( imd_wire6_1_0, wire6_0_0, wire6_0_1);
NANDC2x1 inst_clockedAND_b5_5 ( imd_YF5, CLK, Y5);
NANDC2x1 inst_and_b5_0_2 ( imd_wire5_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b5_2_0 ( imd_Y5, wire5_0_2, wire5_1_0);
NANDC2x1 inst_and_b5_0_1 ( imd_wire5_0_1, A2, A3_inv);
NANDC2x1 inst_and_b5_0_0 ( imd_wire5_0_0, A0, A1_inv);
NANDC2x1 inst_and_b5_1_0 ( imd_wire5_1_0, wire5_0_0, wire5_0_1);
NANDC2x1 inst_and_b4_0_1 ( imd_wire4_0_1, A2, A3_inv);
NANDC2x1 inst_and_b4_0_0 ( imd_wire4_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b4_1_0 ( imd_wire4_1_0, wire4_0_0, wire4_0_1);
NANDC2x1 inst_clockedAND_b4_4 ( imd_YF4, CLK, Y4);
NANDC2x1 inst_and_b4_0_2 ( imd_wire4_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b4_2_0 ( imd_Y4, wire4_0_2, wire4_1_0);
NANDC2x1 inst_clockedAND_b3_3 ( imd_YF3, CLK, Y3);
NANDC2x1 inst_and_b3_0_2 ( imd_wire3_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b3_2_0 ( imd_Y3, wire3_0_2, wire3_1_0);
NANDC2x1 inst_and_b3_0_1 ( imd_wire3_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b3_0_0 ( imd_wire3_0_0, A0, A1);
NANDC2x1 inst_and_b3_1_0 ( imd_wire3_1_0, wire3_0_0, wire3_0_1);
NANDC2x1 inst_and_b2_0_0 ( imd_wire2_0_0, A0_inv, A1);
NANDC2x1 inst_and_b2_0_1 ( imd_wire2_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b2_1_0 ( imd_wire2_1_0, wire2_0_0, wire2_0_1);
NANDC2x1 inst_clockedAND_b2_2 ( imd_YF2, CLK, Y2);
NANDC2x1 inst_and_b2_0_2 ( imd_wire2_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b2_2_0 ( imd_Y2, wire2_0_2, wire2_1_0);
NANDC2x1 inst_and_b1_0_0 ( imd_wire1_0_0, A0, A1_inv);
NANDC2x1 inst_and_b1_0_1 ( imd_wire1_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b1_1_0 ( imd_wire1_1_0, wire1_0_0, wire1_0_1);
NANDC2x1 inst_and_b0_0_0 ( imd_wire0_0_0, A0_inv, A1_inv);
NANDC2x1 inst_and_b0_0_1 ( imd_wire0_0_1, A2_inv, A3_inv);
NANDC2x1 inst_and_b0_1_0 ( imd_wire0_1_0, wire0_0_0, wire0_0_1);
NANDC2x1 inst_clockedAND_b1_1 ( imd_YF1, CLK, Y1);
NANDC2x1 inst_and_b1_0_2 ( imd_wire1_0_2, A4_inv, A5_inv);
NANDC2x1 inst_and_b1_2_0 ( imd_Y1, wire1_0_2, wire1_1_0);
NANDC2x1 inst_and_b0_0_2 ( imd_wire0_0_2, A4_inv, A5_inv);
NANDC2x1 inst_clockedAND_b0_0 ( imd_YF0, CLK, Y0);
NANDC2x1 inst_and_b0_2_0 ( imd_Y0, wire0_0_2, wire0_1_0);
INVC inst_clockedinv_b63_63 ( YF63, imd_YF63);
INVC inst_inv_b63_2_0 ( Y63, imd_Y63);
INVC inst_inv_b63_1_0 ( wire63_1_0, imd_wire63_1_0);
INVC inst_inv_b63_0_2 ( wire63_0_2, imd_wire63_0_2);
INVC inst_inv_b63_0_1 ( wire63_0_1, imd_wire63_0_1);
INVC inst_inv_b63_0_0 ( wire63_0_0, imd_wire63_0_0);
INVC inst_clockedinv_b62_62 ( YF62, imd_YF62);
INVC inst_inv_b62_2_0 ( Y62, imd_Y62);
INVC inst_inv_b62_1_0 ( wire62_1_0, imd_wire62_1_0);
INVC inst_inv_b62_0_2 ( wire62_0_2, imd_wire62_0_2);
INVC inst_inv_b62_0_1 ( wire62_0_1, imd_wire62_0_1);
INVC inst_inv_b62_0_0 ( wire62_0_0, imd_wire62_0_0);
INVC inst_clockedinv_b61_61 ( YF61, imd_YF61);
INVC inst_inv_b61_2_0 ( Y61, imd_Y61);
INVC inst_inv_b61_1_0 ( wire61_1_0, imd_wire61_1_0);
INVC inst_inv_b61_0_2 ( wire61_0_2, imd_wire61_0_2);
INVC inst_inv_b61_0_1 ( wire61_0_1, imd_wire61_0_1);
INVC inst_inv_b61_0_0 ( wire61_0_0, imd_wire61_0_0);
INVC inst_clockedinv_b60_60 ( YF60, imd_YF60);
INVC inst_inv_b60_2_0 ( Y60, imd_Y60);
INVC inst_inv_b60_1_0 ( wire60_1_0, imd_wire60_1_0);
INVC inst_inv_b60_0_2 ( wire60_0_2, imd_wire60_0_2);
INVC inst_inv_b60_0_1 ( wire60_0_1, imd_wire60_0_1);
INVC inst_inv_b60_0_0 ( wire60_0_0, imd_wire60_0_0);
INVC inst_clockedinv_b59_59 ( YF59, imd_YF59);
INVC inst_inv_b59_2_0 ( Y59, imd_Y59);
INVC inst_inv_b59_1_0 ( wire59_1_0, imd_wire59_1_0);
INVC inst_inv_b59_0_2 ( wire59_0_2, imd_wire59_0_2);
INVC inst_inv_b59_0_1 ( wire59_0_1, imd_wire59_0_1);
INVC inst_inv_b59_0_0 ( wire59_0_0, imd_wire59_0_0);
INVC inst_clockedinv_b58_58 ( YF58, imd_YF58);
INVC inst_inv_b58_2_0 ( Y58, imd_Y58);
INVC inst_inv_b58_1_0 ( wire58_1_0, imd_wire58_1_0);
INVC inst_inv_b58_0_2 ( wire58_0_2, imd_wire58_0_2);
INVC inst_inv_b58_0_1 ( wire58_0_1, imd_wire58_0_1);
INVC inst_inv_b58_0_0 ( wire58_0_0, imd_wire58_0_0);
INVC inst_clockedinv_b57_57 ( YF57, imd_YF57);
INVC inst_inv_b57_2_0 ( Y57, imd_Y57);
INVC inst_inv_b57_1_0 ( wire57_1_0, imd_wire57_1_0);
INVC inst_inv_b57_0_2 ( wire57_0_2, imd_wire57_0_2);
INVC inst_inv_b57_0_1 ( wire57_0_1, imd_wire57_0_1);
INVC inst_inv_b57_0_0 ( wire57_0_0, imd_wire57_0_0);
INVC inst_clockedinv_b56_56 ( YF56, imd_YF56);
INVC inst_inv_b56_2_0 ( Y56, imd_Y56);
INVC inst_inv_b56_1_0 ( wire56_1_0, imd_wire56_1_0);
INVC inst_inv_b56_0_2 ( wire56_0_2, imd_wire56_0_2);
INVC inst_inv_b56_0_1 ( wire56_0_1, imd_wire56_0_1);
INVC inst_inv_b56_0_0 ( wire56_0_0, imd_wire56_0_0);
INVC inst_clockedinv_b55_55 ( YF55, imd_YF55);
INVC inst_inv_b55_2_0 ( Y55, imd_Y55);
INVC inst_inv_b55_1_0 ( wire55_1_0, imd_wire55_1_0);
INVC inst_inv_b55_0_2 ( wire55_0_2, imd_wire55_0_2);
INVC inst_inv_b55_0_1 ( wire55_0_1, imd_wire55_0_1);
INVC inst_inv_b55_0_0 ( wire55_0_0, imd_wire55_0_0);
INVC inst_clockedinv_b54_54 ( YF54, imd_YF54);
INVC inst_inv_b54_2_0 ( Y54, imd_Y54);
INVC inst_inv_b54_1_0 ( wire54_1_0, imd_wire54_1_0);
INVC inst_inv_b54_0_0 ( wire54_0_0, imd_wire54_0_0);
INVC inst_inv_b54_0_2 ( wire54_0_2, imd_wire54_0_2);
INVC inst_inv_b54_0_1 ( wire54_0_1, imd_wire54_0_1);
INVC inst_clockedinv_b53_53 ( YF53, imd_YF53);
INVC inst_inv_b53_2_0 ( Y53, imd_Y53);
INVC inst_inv_b53_1_0 ( wire53_1_0, imd_wire53_1_0);
INVC inst_inv_b53_0_2 ( wire53_0_2, imd_wire53_0_2);
INVC inst_clockedinv_b52_52 ( YF52, imd_YF52);
INVC inst_inv_b52_2_0 ( Y52, imd_Y52);
INVC inst_inv_b52_1_0 ( wire52_1_0, imd_wire52_1_0);
INVC inst_inv_b52_0_2 ( wire52_0_2, imd_wire52_0_2);
INVC inst_inv_b52_0_1 ( wire52_0_1, imd_wire52_0_1);
INVC inst_inv_b52_0_0 ( wire52_0_0, imd_wire52_0_0);
INVC inst_clockedinv_b51_51 ( YF51, imd_YF51);
INVC inst_inv_b51_2_0 ( Y51, imd_Y51);
INVC inst_inv_b51_1_0 ( wire51_1_0, imd_wire51_1_0);
INVC inst_inv_b51_0_2 ( wire51_0_2, imd_wire51_0_2);
INVC inst_inv_b51_0_1 ( wire51_0_1, imd_wire51_0_1);
INVC inst_inv_b51_0_0 ( wire51_0_0, imd_wire51_0_0);
INVC inst_clockedinv_b50_50 ( YF50, imd_YF50);
INVC inst_inv_b50_2_0 ( Y50, imd_Y50);
INVC inst_inv_b50_1_0 ( wire50_1_0, imd_wire50_1_0);
INVC inst_inv_b50_0_2 ( wire50_0_2, imd_wire50_0_2);
INVC inst_inv_b50_0_1 ( wire50_0_1, imd_wire50_0_1);
INVC inst_inv_b50_0_0 ( wire50_0_0, imd_wire50_0_0);
INVC inst_clockedinv_b49_49 ( YF49, imd_YF49);
INVC inst_inv_b49_2_0 ( Y49, imd_Y49);
INVC inst_inv_b49_1_0 ( wire49_1_0, imd_wire49_1_0);
INVC inst_inv_b49_0_2 ( wire49_0_2, imd_wire49_0_2);
INVC inst_inv_b49_0_1 ( wire49_0_1, imd_wire49_0_1);
INVC inst_inv_b49_0_0 ( wire49_0_0, imd_wire49_0_0);
INVC inst_clockedinv_b48_48 ( YF48, imd_YF48);
INVC inst_inv_b48_2_0 ( Y48, imd_Y48);
INVC inst_inv_b48_1_0 ( wire48_1_0, imd_wire48_1_0);
INVC inst_inv_b48_0_2 ( wire48_0_2, imd_wire48_0_2);
INVC inst_inv_b48_0_1 ( wire48_0_1, imd_wire48_0_1);
INVC inst_inv_b48_0_0 ( wire48_0_0, imd_wire48_0_0);
INVC inst_clockedinv_b47_47 ( YF47, imd_YF47);
INVC inst_inv_b47_2_0 ( Y47, imd_Y47);
INVC inst_inv_b47_1_0 ( wire47_1_0, imd_wire47_1_0);
INVC inst_inv_b47_0_2 ( wire47_0_2, imd_wire47_0_2);
INVC inst_inv_b47_0_1 ( wire47_0_1, imd_wire47_0_1);
INVC inst_inv_b47_0_0 ( wire47_0_0, imd_wire47_0_0);
INVC inst_clockedinv_b46_46 ( YF46, imd_YF46);
INVC inst_inv_b46_2_0 ( Y46, imd_Y46);
INVC inst_inv_b46_1_0 ( wire46_1_0, imd_wire46_1_0);
INVC inst_inv_b46_0_2 ( wire46_0_2, imd_wire46_0_2);
INVC inst_inv_b46_0_1 ( wire46_0_1, imd_wire46_0_1);
INVC inst_inv_b46_0_0 ( wire46_0_0, imd_wire46_0_0);
INVC inst_clockedinv_b45_45 ( YF45, imd_YF45);
INVC inst_inv_b45_2_0 ( Y45, imd_Y45);
INVC inst_inv_b45_1_0 ( wire45_1_0, imd_wire45_1_0);
INVC inst_inv_b45_0_2 ( wire45_0_2, imd_wire45_0_2);
INVC inst_inv_b45_0_1 ( wire45_0_1, imd_wire45_0_1);
INVC inst_inv_b45_0_0 ( wire45_0_0, imd_wire45_0_0);
INVC inst_clockedinv_b44_44 ( YF44, imd_YF44);
INVC inst_inv_b44_2_0 ( Y44, imd_Y44);
INVC inst_inv_b44_1_0 ( wire44_1_0, imd_wire44_1_0);
INVC inst_inv_b44_0_2 ( wire44_0_2, imd_wire44_0_2);
INVC inst_inv_b44_0_1 ( wire44_0_1, imd_wire44_0_1);
INVC inst_inv_b44_0_0 ( wire44_0_0, imd_wire44_0_0);
INVC inst_clockedinv_b43_43 ( YF43, imd_YF43);
INVC inst_inv_b43_2_0 ( Y43, imd_Y43);
INVC inst_inv_b43_1_0 ( wire43_1_0, imd_wire43_1_0);
INVC inst_inv_b43_0_2 ( wire43_0_2, imd_wire43_0_2);
INVC inst_inv_b43_0_1 ( wire43_0_1, imd_wire43_0_1);
INVC inst_inv_b43_0_0 ( wire43_0_0, imd_wire43_0_0);
INVC inst_inv_b53_0_1 ( wire53_0_1, imd_wire53_0_1);
INVC inst_inv_b53_0_0 ( wire53_0_0, imd_wire53_0_0);
INVC inst_clockedinv_b42_42 ( YF42, imd_YF42);
INVC inst_inv_b42_2_0 ( Y42, imd_Y42);
INVC inst_inv_b42_1_0 ( wire42_1_0, imd_wire42_1_0);
INVC inst_inv_b42_0_2 ( wire42_0_2, imd_wire42_0_2);
INVC inst_inv_b42_0_1 ( wire42_0_1, imd_wire42_0_1);
INVC inst_inv_b42_0_0 ( wire42_0_0, imd_wire42_0_0);
INVC inst_clockedinv_b41_41 ( YF41, imd_YF41);
INVC inst_inv_b41_2_0 ( Y41, imd_Y41);
INVC inst_inv_b41_1_0 ( wire41_1_0, imd_wire41_1_0);
INVC inst_inv_b41_0_2 ( wire41_0_2, imd_wire41_0_2);
INVC inst_inv_b41_0_1 ( wire41_0_1, imd_wire41_0_1);
INVC inst_inv_b41_0_0 ( wire41_0_0, imd_wire41_0_0);
INVC inst_clockedinv_b40_40 ( YF40, imd_YF40);
INVC inst_inv_b40_2_0 ( Y40, imd_Y40);
INVC inst_inv_b40_1_0 ( wire40_1_0, imd_wire40_1_0);
INVC inst_inv_b40_0_2 ( wire40_0_2, imd_wire40_0_2);
INVC inst_inv_b40_0_1 ( wire40_0_1, imd_wire40_0_1);
INVC inst_inv_b40_0_0 ( wire40_0_0, imd_wire40_0_0);
INVC inst_clockedinv_b39_39 ( YF39, imd_YF39);
INVC inst_inv_b39_2_0 ( Y39, imd_Y39);
INVC inst_inv_b39_1_0 ( wire39_1_0, imd_wire39_1_0);
INVC inst_inv_b39_0_2 ( wire39_0_2, imd_wire39_0_2);
INVC inst_inv_b39_0_1 ( wire39_0_1, imd_wire39_0_1);
INVC inst_inv_b39_0_0 ( wire39_0_0, imd_wire39_0_0);
INVC inst_clockedinv_b38_38 ( YF38, imd_YF38);
INVC inst_inv_b38_2_0 ( Y38, imd_Y38);
INVC inst_inv_b38_1_0 ( wire38_1_0, imd_wire38_1_0);
INVC inst_inv_b38_0_2 ( wire38_0_2, imd_wire38_0_2);
INVC inst_inv_b38_0_1 ( wire38_0_1, imd_wire38_0_1);
INVC inst_inv_b38_0_0 ( wire38_0_0, imd_wire38_0_0);
INVC inst_clockedinv_b37_37 ( YF37, imd_YF37);
INVC inst_inv_b37_2_0 ( Y37, imd_Y37);
INVC inst_inv_b37_1_0 ( wire37_1_0, imd_wire37_1_0);
INVC inst_inv_b37_0_2 ( wire37_0_2, imd_wire37_0_2);
INVC inst_inv_b37_0_1 ( wire37_0_1, imd_wire37_0_1);
INVC inst_inv_b37_0_0 ( wire37_0_0, imd_wire37_0_0);
INVC inst_clockedinv_b36_36 ( YF36, imd_YF36);
INVC inst_inv_b36_2_0 ( Y36, imd_Y36);
INVC inst_inv_b36_1_0 ( wire36_1_0, imd_wire36_1_0);
INVC inst_inv_b36_0_2 ( wire36_0_2, imd_wire36_0_2);
INVC inst_inv_b36_0_1 ( wire36_0_1, imd_wire36_0_1);
INVC inst_inv_b36_0_0 ( wire36_0_0, imd_wire36_0_0);
INVC inst_clockedinv_b35_35 ( YF35, imd_YF35);
INVC inst_inv_b35_2_0 ( Y35, imd_Y35);
INVC inst_inv_b35_1_0 ( wire35_1_0, imd_wire35_1_0);
INVC inst_inv_b35_0_2 ( wire35_0_2, imd_wire35_0_2);
INVC inst_inv_b35_0_1 ( wire35_0_1, imd_wire35_0_1);
INVC inst_inv_b35_0_0 ( wire35_0_0, imd_wire35_0_0);
INVC inst_clockedinv_b34_34 ( YF34, imd_YF34);
INVC inst_inv_b34_2_0 ( Y34, imd_Y34);
INVC inst_inv_b34_1_0 ( wire34_1_0, imd_wire34_1_0);
INVC inst_inv_b34_0_2 ( wire34_0_2, imd_wire34_0_2);
INVC inst_inv_b34_0_1 ( wire34_0_1, imd_wire34_0_1);
INVC inst_inv_b34_0_0 ( wire34_0_0, imd_wire34_0_0);
INVC inst_clockedinv_b33_33 ( YF33, imd_YF33);
INVC inst_inv_b33_2_0 ( Y33, imd_Y33);
INVC inst_inv_b33_1_0 ( wire33_1_0, imd_wire33_1_0);
INVC inst_inv_b33_0_2 ( wire33_0_2, imd_wire33_0_2);
INVC inst_inv_b33_0_1 ( wire33_0_1, imd_wire33_0_1);
INVC inst_inv_b33_0_0 ( wire33_0_0, imd_wire33_0_0);
INVC inst_inv_b32_0_2 ( wire32_0_2, imd_wire32_0_2);
INVC inst_inv_b32_2_0 ( Y32, imd_Y32);
INVC inst_clockedinv_b32_32 ( YF32, imd_YF32);
INVC inst_inv_b32_1_0 ( wire32_1_0, imd_wire32_1_0);
INVC inst_inv_b32_0_1 ( wire32_0_1, imd_wire32_0_1);
INVC inst_inv_b32_0_0 ( wire32_0_0, imd_wire32_0_0);
INVC inst_clockedinv_b31_31 ( YF31, imd_YF31);
INVC inst_inv_b31_2_0 ( Y31, imd_Y31);
INVC inst_inv_b31_1_0 ( wire31_1_0, imd_wire31_1_0);
INVC inst_inv_b31_0_2 ( wire31_0_2, imd_wire31_0_2);
INVC inst_inv_b31_0_1 ( wire31_0_1, imd_wire31_0_1);
INVC inst_inv_b31_0_0 ( wire31_0_0, imd_wire31_0_0);
INVC inst_clockedinv_b30_30 ( YF30, imd_YF30);
INVC inst_inv_b30_2_0 ( Y30, imd_Y30);
INVC inst_inv_b30_1_0 ( wire30_1_0, imd_wire30_1_0);
INVC inst_inv_b30_0_2 ( wire30_0_2, imd_wire30_0_2);
INVC inst_inv_b30_0_1 ( wire30_0_1, imd_wire30_0_1);
INVC inst_inv_b30_0_0 ( wire30_0_0, imd_wire30_0_0);
INVC inst_clockedinv_b29_29 ( YF29, imd_YF29);
INVC inst_inv_b29_2_0 ( Y29, imd_Y29);
INVC inst_inv_b29_1_0 ( wire29_1_0, imd_wire29_1_0);
INVC inst_inv_b29_0_2 ( wire29_0_2, imd_wire29_0_2);
INVC inst_inv_b29_0_1 ( wire29_0_1, imd_wire29_0_1);
INVC inst_inv_b29_0_0 ( wire29_0_0, imd_wire29_0_0);
INVC inst_clockedinv_b28_28 ( YF28, imd_YF28);
INVC inst_inv_b28_2_0 ( Y28, imd_Y28);
INVC inst_inv_b28_1_0 ( wire28_1_0, imd_wire28_1_0);
INVC inst_inv_b28_0_2 ( wire28_0_2, imd_wire28_0_2);
INVC inst_inv_b28_0_1 ( wire28_0_1, imd_wire28_0_1);
INVC inst_inv_b28_0_0 ( wire28_0_0, imd_wire28_0_0);
INVC inst_clockedinv_b27_27 ( YF27, imd_YF27);
INVC inst_inv_b27_2_0 ( Y27, imd_Y27);
INVC inst_inv_b27_1_0 ( wire27_1_0, imd_wire27_1_0);
INVC inst_inv_b27_0_2 ( wire27_0_2, imd_wire27_0_2);
INVC inst_inv_b27_0_1 ( wire27_0_1, imd_wire27_0_1);
INVC inst_inv_b27_0_0 ( wire27_0_0, imd_wire27_0_0);
INVC inst_clockedinv_b26_26 ( YF26, imd_YF26);
INVC inst_inv_b26_2_0 ( Y26, imd_Y26);
INVC inst_inv_b26_1_0 ( wire26_1_0, imd_wire26_1_0);
INVC inst_inv_b26_0_2 ( wire26_0_2, imd_wire26_0_2);
INVC inst_inv_b26_0_1 ( wire26_0_1, imd_wire26_0_1);
INVC inst_inv_b26_0_0 ( wire26_0_0, imd_wire26_0_0);
INVC inst_clockedinv_b25_25 ( YF25, imd_YF25);
INVC inst_inv_b25_2_0 ( Y25, imd_Y25);
INVC inst_inv_b25_1_0 ( wire25_1_0, imd_wire25_1_0);
INVC inst_inv_b25_0_2 ( wire25_0_2, imd_wire25_0_2);
INVC inst_inv_b25_0_1 ( wire25_0_1, imd_wire25_0_1);
INVC inst_inv_b25_0_0 ( wire25_0_0, imd_wire25_0_0);
INVC inst_clockedinv_b24_24 ( YF24, imd_YF24);
INVC inst_inv_b24_2_0 ( Y24, imd_Y24);
INVC inst_inv_b24_1_0 ( wire24_1_0, imd_wire24_1_0);
INVC inst_inv_b24_0_2 ( wire24_0_2, imd_wire24_0_2);
INVC inst_inv_b24_0_1 ( wire24_0_1, imd_wire24_0_1);
INVC inst_inv_b24_0_0 ( wire24_0_0, imd_wire24_0_0);
INVC inst_clockedinv_b23_23 ( YF23, imd_YF23);
INVC inst_inv_b23_2_0 ( Y23, imd_Y23);
INVC inst_inv_b23_1_0 ( wire23_1_0, imd_wire23_1_0);
INVC inst_inv_b23_0_2 ( wire23_0_2, imd_wire23_0_2);
INVC inst_inv_b23_0_1 ( wire23_0_1, imd_wire23_0_1);
INVC inst_inv_b23_0_0 ( wire23_0_0, imd_wire23_0_0);
INVC inst_clockedinv_b22_22 ( YF22, imd_YF22);
INVC inst_inv_b22_2_0 ( Y22, imd_Y22);
INVC inst_inv_b22_1_0 ( wire22_1_0, imd_wire22_1_0);
INVC inst_inv_b22_0_0 ( wire22_0_0, imd_wire22_0_0);
INVC inst_inv_b22_0_2 ( wire22_0_2, imd_wire22_0_2);
INVC inst_inv_b22_0_1 ( wire22_0_1, imd_wire22_0_1);
INVC inst_clockedinv_b21_21 ( YF21, imd_YF21);
INVC inst_inv_b21_2_0 ( Y21, imd_Y21);
INVC inst_inv_b21_1_0 ( wire21_1_0, imd_wire21_1_0);
INVC inst_inv_b21_0_2 ( wire21_0_2, imd_wire21_0_2);
INVC inst_clockedinv_b20_20 ( YF20, imd_YF20);
INVC inst_inv_b20_2_0 ( Y20, imd_Y20);
INVC inst_inv_b20_1_0 ( wire20_1_0, imd_wire20_1_0);
INVC inst_inv_b20_0_2 ( wire20_0_2, imd_wire20_0_2);
INVC inst_inv_b20_0_1 ( wire20_0_1, imd_wire20_0_1);
INVC inst_inv_b20_0_0 ( wire20_0_0, imd_wire20_0_0);
INVC inst_clockedinv_b19_19 ( YF19, imd_YF19);
INVC inst_inv_b19_2_0 ( Y19, imd_Y19);
INVC inst_inv_b19_1_0 ( wire19_1_0, imd_wire19_1_0);
INVC inst_inv_b19_0_2 ( wire19_0_2, imd_wire19_0_2);
INVC inst_inv_b19_0_1 ( wire19_0_1, imd_wire19_0_1);
INVC inst_inv_b19_0_0 ( wire19_0_0, imd_wire19_0_0);
INVC inst_clockedinv_b18_18 ( YF18, imd_YF18);
INVC inst_inv_b18_2_0 ( Y18, imd_Y18);
INVC inst_inv_b18_1_0 ( wire18_1_0, imd_wire18_1_0);
INVC inst_inv_b18_0_2 ( wire18_0_2, imd_wire18_0_2);
INVC inst_inv_b18_0_1 ( wire18_0_1, imd_wire18_0_1);
INVC inst_inv_b18_0_0 ( wire18_0_0, imd_wire18_0_0);
INVC inst_clockedinv_b17_17 ( YF17, imd_YF17);
INVC inst_inv_b17_2_0 ( Y17, imd_Y17);
INVC inst_inv_b17_1_0 ( wire17_1_0, imd_wire17_1_0);
INVC inst_inv_b17_0_2 ( wire17_0_2, imd_wire17_0_2);
INVC inst_inv_b17_0_1 ( wire17_0_1, imd_wire17_0_1);
INVC inst_inv_b17_0_0 ( wire17_0_0, imd_wire17_0_0);
INVC inst_inv_b16_0_2 ( wire16_0_2, imd_wire16_0_2);
INVC inst_inv_b16_2_0 ( Y16, imd_Y16);
INVC inst_clockedinv_b16_16 ( YF16, imd_YF16);
INVC inst_inv_b16_1_0 ( wire16_1_0, imd_wire16_1_0);
INVC inst_inv_b16_0_1 ( wire16_0_1, imd_wire16_0_1);
INVC inst_inv_b16_0_0 ( wire16_0_0, imd_wire16_0_0);
INVC inst_clockedinv_b15_15 ( YF15, imd_YF15);
INVC inst_inv_b15_2_0 ( Y15, imd_Y15);
INVC inst_inv_b15_1_0 ( wire15_1_0, imd_wire15_1_0);
INVC inst_inv_b15_0_2 ( wire15_0_2, imd_wire15_0_2);
INVC inst_inv_b15_0_1 ( wire15_0_1, imd_wire15_0_1);
INVC inst_inv_b15_0_0 ( wire15_0_0, imd_wire15_0_0);
INVC inst_clockedinv_b14_14 ( YF14, imd_YF14);
INVC inst_inv_b14_2_0 ( Y14, imd_Y14);
INVC inst_inv_b14_1_0 ( wire14_1_0, imd_wire14_1_0);
INVC inst_inv_b14_0_2 ( wire14_0_2, imd_wire14_0_2);
INVC inst_inv_b14_0_1 ( wire14_0_1, imd_wire14_0_1);
INVC inst_inv_b14_0_0 ( wire14_0_0, imd_wire14_0_0);
INVC inst_clockedinv_b13_13 ( YF13, imd_YF13);
INVC inst_inv_b13_2_0 ( Y13, imd_Y13);
INVC inst_inv_b13_1_0 ( wire13_1_0, imd_wire13_1_0);
INVC inst_inv_b13_0_2 ( wire13_0_2, imd_wire13_0_2);
INVC inst_inv_b13_0_1 ( wire13_0_1, imd_wire13_0_1);
INVC inst_inv_b13_0_0 ( wire13_0_0, imd_wire13_0_0);
INVC inst_clockedinv_b12_12 ( YF12, imd_YF12);
INVC inst_inv_b12_2_0 ( Y12, imd_Y12);
INVC inst_inv_b12_1_0 ( wire12_1_0, imd_wire12_1_0);
INVC inst_inv_b12_0_2 ( wire12_0_2, imd_wire12_0_2);
INVC inst_inv_b12_0_1 ( wire12_0_1, imd_wire12_0_1);
INVC inst_inv_b12_0_0 ( wire12_0_0, imd_wire12_0_0);
INVC inst_clockedinv_b11_11 ( YF11, imd_YF11);
INVC inst_inv_b11_2_0 ( Y11, imd_Y11);
INVC inst_inv_b11_1_0 ( wire11_1_0, imd_wire11_1_0);
INVC inst_inv_b11_0_2 ( wire11_0_2, imd_wire11_0_2);
INVC inst_inv_b11_0_1 ( wire11_0_1, imd_wire11_0_1);
INVC inst_inv_b11_0_0 ( wire11_0_0, imd_wire11_0_0);
INVC inst_inv_b21_0_1 ( wire21_0_1, imd_wire21_0_1);
INVC inst_inv_b21_0_0 ( wire21_0_0, imd_wire21_0_0);
INVC inst_clockedinv_b10_10 ( YF10, imd_YF10);
INVC inst_inv_b10_2_0 ( Y10, imd_Y10);
INVC inst_inv_b10_1_0 ( wire10_1_0, imd_wire10_1_0);
INVC inst_inv_b10_0_2 ( wire10_0_2, imd_wire10_0_2);
INVC inst_inv_b10_0_1 ( wire10_0_1, imd_wire10_0_1);
INVC inst_inv_b10_0_0 ( wire10_0_0, imd_wire10_0_0);
INVC inst_clockedinv_b9_9 ( YF9, imd_YF9);
INVC inst_inv_b9_2_0 ( Y9, imd_Y9);
INVC inst_inv_b9_1_0 ( wire9_1_0, imd_wire9_1_0);
INVC inst_inv_b9_0_2 ( wire9_0_2, imd_wire9_0_2);
INVC inst_inv_b9_0_1 ( wire9_0_1, imd_wire9_0_1);
INVC inst_inv_b9_0_0 ( wire9_0_0, imd_wire9_0_0);
INVC inst_inv_b8_0_1 ( wire8_0_1, imd_wire8_0_1);
INVC inst_inv_b8_1_0 ( wire8_1_0, imd_wire8_1_0);
INVC inst_inv_b8_0_0 ( wire8_0_0, imd_wire8_0_0);
INVC inst_inv_b8_2_0 ( Y8, imd_Y8);
INVC inst_clockedinv_b8_8 ( YF8, imd_YF8);
INVC inst_inv_b8_0_2 ( wire8_0_2, imd_wire8_0_2);
INVC inst_clockedinv_b7_7 ( YF7, imd_YF7);
INVC inst_inv_b7_2_0 ( Y7, imd_Y7);
INVC inst_inv_b7_1_0 ( wire7_1_0, imd_wire7_1_0);
INVC inst_inv_b7_0_2 ( wire7_0_2, imd_wire7_0_2);
INVC inst_inv_b7_0_1 ( wire7_0_1, imd_wire7_0_1);
INVC inst_inv_b7_0_0 ( wire7_0_0, imd_wire7_0_0);
INVC inst_clockedinv_b6_6 ( YF6, imd_YF6);
INVC inst_inv_b6_2_0 ( Y6, imd_Y6);
INVC inst_inv_b6_1_0 ( wire6_1_0, imd_wire6_1_0);
INVC inst_inv_b6_0_2 ( wire6_0_2, imd_wire6_0_2);
INVC inst_inv_b6_0_1 ( wire6_0_1, imd_wire6_0_1);
INVC inst_inv_b6_0_0 ( wire6_0_0, imd_wire6_0_0);
INVC inst_clockedinv_b5_5 ( YF5, imd_YF5);
INVC inst_inv_b5_2_0 ( Y5, imd_Y5);
INVC inst_inv_b5_1_0 ( wire5_1_0, imd_wire5_1_0);
INVC inst_inv_b5_0_2 ( wire5_0_2, imd_wire5_0_2);
INVC inst_inv_b5_0_1 ( wire5_0_1, imd_wire5_0_1);
INVC inst_inv_b5_0_0 ( wire5_0_0, imd_wire5_0_0);
INVC inst_inv_b4_0_1 ( wire4_0_1, imd_wire4_0_1);
INVC inst_inv_b4_1_0 ( wire4_1_0, imd_wire4_1_0);
INVC inst_inv_b4_0_0 ( wire4_0_0, imd_wire4_0_0);
INVC inst_inv_b4_2_0 ( Y4, imd_Y4);
INVC inst_clockedinv_b4_4 ( YF4, imd_YF4);
INVC inst_inv_b4_0_2 ( wire4_0_2, imd_wire4_0_2);
INVC inst_clockedinv_b3_3 ( YF3, imd_YF3);
INVC inst_inv_b3_2_0 ( Y3, imd_Y3);
INVC inst_inv_b3_1_0 ( wire3_1_0, imd_wire3_1_0);
INVC inst_inv_b3_0_2 ( wire3_0_2, imd_wire3_0_2);
INVC inst_inv_b3_0_1 ( wire3_0_1, imd_wire3_0_1);
INVC inst_inv_b3_0_0 ( wire3_0_0, imd_wire3_0_0);
INVC inst_inv_b2_0_0 ( wire2_0_0, imd_wire2_0_0);
INVC inst_inv_b2_1_0 ( wire2_1_0, imd_wire2_1_0);
INVC inst_inv_b2_0_1 ( wire2_0_1, imd_wire2_0_1);
INVC inst_inv_b2_2_0 ( Y2, imd_Y2);
INVC inst_clockedinv_b2_2 ( YF2, imd_YF2);
INVC inst_inv_b2_0_2 ( wire2_0_2, imd_wire2_0_2);
INVC inst_inv_b1_0_0 ( wire1_0_0, imd_wire1_0_0);
INVC inst_inv_b1_1_0 ( wire1_1_0, imd_wire1_1_0);
INVC inst_inv_b1_0_1 ( wire1_0_1, imd_wire1_0_1);
INVC inst_inv_b0_0_0 ( wire0_0_0, imd_wire0_0_0);
INVC inst_inv_b0_0_1 ( wire0_0_1, imd_wire0_0_1);
INVC inst_inv_b0_1_0 ( wire0_1_0, imd_wire0_1_0);
INVC inst_inv_b1_2_0 ( Y1, imd_Y1);
INVC inst_clockedinv_b1_1 ( YF1, imd_YF1);
INVC inst_inv_b1_0_2 ( wire1_0_2, imd_wire1_0_2);
INVC inst_inv_b0_0_2 ( wire0_0_2, imd_wire0_0_2);
INVC inst_inv_b0_2_0 ( Y0, imd_Y0);
INVC inst_clockedinv_b0_0 ( YF0, imd_YF0);

endmodule
// Library - sram_compiled_20201119_153347_r64_c64_w8, Cell -
//sram_compiled_array, View - schematic
// LAST TIME SAVED: Nov 19 15:34:19 2020
// NETLIST TIME: Apr  5 11:21:05 2021
`timescale 1ns / 1ps 

module sram_compiled_array ( addr0, addr1, addr2, addr3, addr4, addr5,
     addr6, addr7, addr8, din0, din1, din2, din3, din4, din5, din6,
     din7, dout0, dout1, dout2, dout3, dout4, dout5, dout6, dout7, clk,
     write_en, sense_en );

output  dout0, dout1, dout2, dout3, dout4, dout5, dout6, dout7;

input  addr0, addr1, addr2, addr3, addr4, addr5, addr6, addr7, addr8,
     clk, din0, din1, din2, din3, din4, din5, din6, din7, sense_en,
     write_en;


specify

    (sense_en  => dout0 ) = 0.6;   

    (sense_en  => dout1 ) = 0.7;   

    (sense_en  => dout2 ) = 0.7;   

    (sense_en  => dout3 ) = 0.6;  

    (sense_en  => dout4 ) = 0.6;   

    (sense_en  => dout5 ) = 0.7;   

    (sense_en  => dout6 ) = 0.7;   

    (sense_en  => dout7 ) = 0.6;  


endspecify

sram_cell_6t_3 inst_cell_63_63 ( BL63, BLN63, WL63);
sram_cell_6t_3 inst_cell_63_62 ( BL62, BLN62, WL63);
sram_cell_6t_3 inst_cell_63_61 ( BL61, BLN61, WL63);
sram_cell_6t_3 inst_cell_63_60 ( BL60, BLN60, WL63);
sram_cell_6t_3 inst_cell_63_59 ( BL59, BLN59, WL63);
sram_cell_6t_3 inst_cell_63_58 ( BL58, BLN58, WL63);
sram_cell_6t_3 inst_cell_63_57 ( BL57, BLN57, WL63);
sram_cell_6t_3 inst_cell_63_56 ( BL56, BLN56, WL63);
sram_cell_6t_3 inst_cell_63_55 ( BL55, BLN55, WL63);
sram_cell_6t_3 inst_cell_63_54 ( BL54, BLN54, WL63);
sram_cell_6t_3 inst_cell_63_53 ( BL53, BLN53, WL63);
sram_cell_6t_3 inst_cell_63_52 ( BL52, BLN52, WL63);
sram_cell_6t_3 inst_cell_63_51 ( BL51, BLN51, WL63);
sram_cell_6t_3 inst_cell_63_50 ( BL50, BLN50, WL63);
sram_cell_6t_3 inst_cell_63_49 ( BL49, BLN49, WL63);
sram_cell_6t_3 inst_cell_63_48 ( BL48, BLN48, WL63);
sram_cell_6t_3 inst_cell_63_47 ( BL47, BLN47, WL63);
sram_cell_6t_3 inst_cell_63_46 ( BL46, BLN46, WL63);
sram_cell_6t_3 inst_cell_63_45 ( BL45, BLN45, WL63);
sram_cell_6t_3 inst_cell_63_44 ( BL44, BLN44, WL63);
sram_cell_6t_3 inst_cell_63_43 ( BL43, BLN43, WL63);
sram_cell_6t_3 inst_cell_63_42 ( BL42, BLN42, WL63);
sram_cell_6t_3 inst_cell_63_41 ( BL41, BLN41, WL63);
sram_cell_6t_3 inst_cell_63_40 ( BL40, BLN40, WL63);
sram_cell_6t_3 inst_cell_63_39 ( BL39, BLN39, WL63);
sram_cell_6t_3 inst_cell_63_38 ( BL38, BLN38, WL63);
sram_cell_6t_3 inst_cell_63_37 ( BL37, BLN37, WL63);
sram_cell_6t_3 inst_cell_63_36 ( BL36, BLN36, WL63);
sram_cell_6t_3 inst_cell_63_35 ( BL35, BLN35, WL63);
sram_cell_6t_3 inst_cell_63_34 ( BL34, BLN34, WL63);
sram_cell_6t_3 inst_cell_62_55 ( BL55, BLN55, WL62);
sram_cell_6t_3 inst_cell_62_54 ( BL54, BLN54, WL62);
sram_cell_6t_3 inst_cell_62_53 ( BL53, BLN53, WL62);
sram_cell_6t_3 inst_cell_62_52 ( BL52, BLN52, WL62);
sram_cell_6t_3 inst_cell_62_51 ( BL51, BLN51, WL62);
sram_cell_6t_3 inst_cell_62_50 ( BL50, BLN50, WL62);
sram_cell_6t_3 inst_cell_62_49 ( BL49, BLN49, WL62);
sram_cell_6t_3 inst_cell_62_48 ( BL48, BLN48, WL62);
sram_cell_6t_3 inst_cell_63_33 ( BL33, BLN33, WL63);
sram_cell_6t_3 inst_cell_63_32 ( BL32, BLN32, WL63);
sram_cell_6t_3 inst_cell_63_31 ( BL31, BLN31, WL63);
sram_cell_6t_3 inst_cell_63_30 ( BL30, BLN30, WL63);
sram_cell_6t_3 inst_cell_63_29 ( BL29, BLN29, WL63);
sram_cell_6t_3 inst_cell_63_28 ( BL28, BLN28, WL63);
sram_cell_6t_3 inst_cell_63_27 ( BL27, BLN27, WL63);
sram_cell_6t_3 inst_cell_63_26 ( BL26, BLN26, WL63);
sram_cell_6t_3 inst_cell_63_25 ( BL25, BLN25, WL63);
sram_cell_6t_3 inst_cell_63_24 ( BL24, BLN24, WL63);
sram_cell_6t_3 inst_cell_63_23 ( BL23, BLN23, WL63);
sram_cell_6t_3 inst_cell_63_22 ( BL22, BLN22, WL63);
sram_cell_6t_3 inst_cell_63_21 ( BL21, BLN21, WL63);
sram_cell_6t_3 inst_cell_63_20 ( BL20, BLN20, WL63);
sram_cell_6t_3 inst_cell_63_19 ( BL19, BLN19, WL63);
sram_cell_6t_3 inst_cell_63_18 ( BL18, BLN18, WL63);
sram_cell_6t_3 inst_cell_63_17 ( BL17, BLN17, WL63);
sram_cell_6t_3 inst_cell_63_16 ( BL16, BLN16, WL63);
sram_cell_6t_3 inst_cell_63_15 ( BL15, BLN15, WL63);
sram_cell_6t_3 inst_cell_63_14 ( BL14, BLN14, WL63);
sram_cell_6t_3 inst_cell_63_13 ( BL13, BLN13, WL63);
sram_cell_6t_3 inst_cell_63_12 ( BL12, BLN12, WL63);
sram_cell_6t_3 inst_cell_63_11 ( BL11, BLN11, WL63);
sram_cell_6t_3 inst_cell_63_10 ( BL10, BLN10, WL63);
sram_cell_6t_3 inst_cell_63_9 ( BL9, BLN9, WL63);
sram_cell_6t_3 inst_cell_63_8 ( BL8, BLN8, WL63);
sram_cell_6t_3 inst_cell_63_7 ( BL7, BLN7, WL63);
sram_cell_6t_3 inst_cell_63_6 ( BL6, BLN6, WL63);
sram_cell_6t_3 inst_cell_63_5 ( BL5, BLN5, WL63);
sram_cell_6t_3 inst_cell_63_4 ( BL4, BLN4, WL63);
sram_cell_6t_3 inst_cell_63_3 ( BL3, BLN3, WL63);
sram_cell_6t_3 inst_cell_63_2 ( BL2, BLN2, WL63);
sram_cell_6t_3 inst_cell_63_1 ( BL1, BLN1, WL63);
sram_cell_6t_3 inst_cell_63_0 ( BL0, BLN0, WL63);
sram_cell_6t_3 inst_cell_62_63 ( BL63, BLN63, WL62);
sram_cell_6t_3 inst_cell_62_62 ( BL62, BLN62, WL62);
sram_cell_6t_3 inst_cell_62_61 ( BL61, BLN61, WL62);
sram_cell_6t_3 inst_cell_62_60 ( BL60, BLN60, WL62);
sram_cell_6t_3 inst_cell_62_59 ( BL59, BLN59, WL62);
sram_cell_6t_3 inst_cell_62_58 ( BL58, BLN58, WL62);
sram_cell_6t_3 inst_cell_62_57 ( BL57, BLN57, WL62);
sram_cell_6t_3 inst_cell_62_56 ( BL56, BLN56, WL62);
sram_cell_6t_3 inst_cell_62_47 ( BL47, BLN47, WL62);
sram_cell_6t_3 inst_cell_62_46 ( BL46, BLN46, WL62);
sram_cell_6t_3 inst_cell_62_45 ( BL45, BLN45, WL62);
sram_cell_6t_3 inst_cell_62_44 ( BL44, BLN44, WL62);
sram_cell_6t_3 inst_cell_62_43 ( BL43, BLN43, WL62);
sram_cell_6t_3 inst_cell_62_42 ( BL42, BLN42, WL62);
sram_cell_6t_3 inst_cell_62_41 ( BL41, BLN41, WL62);
sram_cell_6t_3 inst_cell_62_40 ( BL40, BLN40, WL62);
sram_cell_6t_3 inst_cell_62_39 ( BL39, BLN39, WL62);
sram_cell_6t_3 inst_cell_62_38 ( BL38, BLN38, WL62);
sram_cell_6t_3 inst_cell_62_37 ( BL37, BLN37, WL62);
sram_cell_6t_3 inst_cell_62_36 ( BL36, BLN36, WL62);
sram_cell_6t_3 inst_cell_62_35 ( BL35, BLN35, WL62);
sram_cell_6t_3 inst_cell_61_47 ( BL47, BLN47, WL61);
sram_cell_6t_3 inst_cell_61_46 ( BL46, BLN46, WL61);
sram_cell_6t_3 inst_cell_61_45 ( BL45, BLN45, WL61);
sram_cell_6t_3 inst_cell_61_44 ( BL44, BLN44, WL61);
sram_cell_6t_3 inst_cell_61_43 ( BL43, BLN43, WL61);
sram_cell_6t_3 inst_cell_61_42 ( BL42, BLN42, WL61);
sram_cell_6t_3 inst_cell_61_41 ( BL41, BLN41, WL61);
sram_cell_6t_3 inst_cell_61_40 ( BL40, BLN40, WL61);
sram_cell_6t_3 inst_cell_62_34 ( BL34, BLN34, WL62);
sram_cell_6t_3 inst_cell_62_33 ( BL33, BLN33, WL62);
sram_cell_6t_3 inst_cell_62_32 ( BL32, BLN32, WL62);
sram_cell_6t_3 inst_cell_62_31 ( BL31, BLN31, WL62);
sram_cell_6t_3 inst_cell_62_30 ( BL30, BLN30, WL62);
sram_cell_6t_3 inst_cell_62_29 ( BL29, BLN29, WL62);
sram_cell_6t_3 inst_cell_62_28 ( BL28, BLN28, WL62);
sram_cell_6t_3 inst_cell_62_27 ( BL27, BLN27, WL62);
sram_cell_6t_3 inst_cell_62_26 ( BL26, BLN26, WL62);
sram_cell_6t_3 inst_cell_62_25 ( BL25, BLN25, WL62);
sram_cell_6t_3 inst_cell_62_24 ( BL24, BLN24, WL62);
sram_cell_6t_3 inst_cell_62_23 ( BL23, BLN23, WL62);
sram_cell_6t_3 inst_cell_62_22 ( BL22, BLN22, WL62);
sram_cell_6t_3 inst_cell_62_21 ( BL21, BLN21, WL62);
sram_cell_6t_3 inst_cell_62_20 ( BL20, BLN20, WL62);
sram_cell_6t_3 inst_cell_62_19 ( BL19, BLN19, WL62);
sram_cell_6t_3 inst_cell_62_18 ( BL18, BLN18, WL62);
sram_cell_6t_3 inst_cell_62_17 ( BL17, BLN17, WL62);
sram_cell_6t_3 inst_cell_62_16 ( BL16, BLN16, WL62);
sram_cell_6t_3 inst_cell_62_15 ( BL15, BLN15, WL62);
sram_cell_6t_3 inst_cell_62_14 ( BL14, BLN14, WL62);
sram_cell_6t_3 inst_cell_62_13 ( BL13, BLN13, WL62);
sram_cell_6t_3 inst_cell_62_12 ( BL12, BLN12, WL62);
sram_cell_6t_3 inst_cell_62_11 ( BL11, BLN11, WL62);
sram_cell_6t_3 inst_cell_62_10 ( BL10, BLN10, WL62);
sram_cell_6t_3 inst_cell_62_9 ( BL9, BLN9, WL62);
sram_cell_6t_3 inst_cell_62_8 ( BL8, BLN8, WL62);
sram_cell_6t_3 inst_cell_62_7 ( BL7, BLN7, WL62);
sram_cell_6t_3 inst_cell_62_6 ( BL6, BLN6, WL62);
sram_cell_6t_3 inst_cell_62_5 ( BL5, BLN5, WL62);
sram_cell_6t_3 inst_cell_62_4 ( BL4, BLN4, WL62);
sram_cell_6t_3 inst_cell_62_3 ( BL3, BLN3, WL62);
sram_cell_6t_3 inst_cell_62_2 ( BL2, BLN2, WL62);
sram_cell_6t_3 inst_cell_62_1 ( BL1, BLN1, WL62);
sram_cell_6t_3 inst_cell_62_0 ( BL0, BLN0, WL62);
sram_cell_6t_3 inst_cell_61_63 ( BL63, BLN63, WL61);
sram_cell_6t_3 inst_cell_61_62 ( BL62, BLN62, WL61);
sram_cell_6t_3 inst_cell_61_61 ( BL61, BLN61, WL61);
sram_cell_6t_3 inst_cell_61_60 ( BL60, BLN60, WL61);
sram_cell_6t_3 inst_cell_61_59 ( BL59, BLN59, WL61);
sram_cell_6t_3 inst_cell_61_58 ( BL58, BLN58, WL61);
sram_cell_6t_3 inst_cell_61_57 ( BL57, BLN57, WL61);
sram_cell_6t_3 inst_cell_61_56 ( BL56, BLN56, WL61);
sram_cell_6t_3 inst_cell_61_55 ( BL55, BLN55, WL61);
sram_cell_6t_3 inst_cell_61_54 ( BL54, BLN54, WL61);
sram_cell_6t_3 inst_cell_61_53 ( BL53, BLN53, WL61);
sram_cell_6t_3 inst_cell_61_52 ( BL52, BLN52, WL61);
sram_cell_6t_3 inst_cell_61_51 ( BL51, BLN51, WL61);
sram_cell_6t_3 inst_cell_61_50 ( BL50, BLN50, WL61);
sram_cell_6t_3 inst_cell_61_49 ( BL49, BLN49, WL61);
sram_cell_6t_3 inst_cell_61_48 ( BL48, BLN48, WL61);
sram_cell_6t_3 inst_cell_61_39 ( BL39, BLN39, WL61);
sram_cell_6t_3 inst_cell_61_38 ( BL38, BLN38, WL61);
sram_cell_6t_3 inst_cell_61_37 ( BL37, BLN37, WL61);
sram_cell_6t_3 inst_cell_61_36 ( BL36, BLN36, WL61);
sram_cell_6t_3 inst_cell_61_35 ( BL35, BLN35, WL61);
sram_cell_6t_3 inst_cell_61_34 ( BL34, BLN34, WL61);
sram_cell_6t_3 inst_cell_61_33 ( BL33, BLN33, WL61);
sram_cell_6t_3 inst_cell_61_32 ( BL32, BLN32, WL61);
sram_cell_6t_3 inst_cell_61_31 ( BL31, BLN31, WL61);
sram_cell_6t_3 inst_cell_61_30 ( BL30, BLN30, WL61);
sram_cell_6t_3 inst_cell_61_29 ( BL29, BLN29, WL61);
sram_cell_6t_3 inst_cell_61_28 ( BL28, BLN28, WL61);
sram_cell_6t_3 inst_cell_61_27 ( BL27, BLN27, WL61);
sram_cell_6t_3 inst_cell_61_26 ( BL26, BLN26, WL61);
sram_cell_6t_3 inst_cell_61_25 ( BL25, BLN25, WL61);
sram_cell_6t_3 inst_cell_61_24 ( BL24, BLN24, WL61);
sram_cell_6t_3 inst_cell_61_23 ( BL23, BLN23, WL61);
sram_cell_6t_3 inst_cell_61_22 ( BL22, BLN22, WL61);
sram_cell_6t_3 inst_cell_61_21 ( BL21, BLN21, WL61);
sram_cell_6t_3 inst_cell_61_20 ( BL20, BLN20, WL61);
sram_cell_6t_3 inst_cell_61_19 ( BL19, BLN19, WL61);
sram_cell_6t_3 inst_cell_61_18 ( BL18, BLN18, WL61);
sram_cell_6t_3 inst_cell_61_17 ( BL17, BLN17, WL61);
sram_cell_6t_3 inst_cell_61_16 ( BL16, BLN16, WL61);
sram_cell_6t_3 inst_cell_61_15 ( BL15, BLN15, WL61);
sram_cell_6t_3 inst_cell_61_14 ( BL14, BLN14, WL61);
sram_cell_6t_3 inst_cell_61_13 ( BL13, BLN13, WL61);
sram_cell_6t_3 inst_cell_61_12 ( BL12, BLN12, WL61);
sram_cell_6t_3 inst_cell_61_11 ( BL11, BLN11, WL61);
sram_cell_6t_3 inst_cell_61_10 ( BL10, BLN10, WL61);
sram_cell_6t_3 inst_cell_61_9 ( BL9, BLN9, WL61);
sram_cell_6t_3 inst_cell_61_8 ( BL8, BLN8, WL61);
sram_cell_6t_3 inst_cell_61_7 ( BL7, BLN7, WL61);
sram_cell_6t_3 inst_cell_61_6 ( BL6, BLN6, WL61);
sram_cell_6t_3 inst_cell_61_5 ( BL5, BLN5, WL61);
sram_cell_6t_3 inst_cell_61_4 ( BL4, BLN4, WL61);
sram_cell_6t_3 inst_cell_61_3 ( BL3, BLN3, WL61);
sram_cell_6t_3 inst_cell_61_2 ( BL2, BLN2, WL61);
sram_cell_6t_3 inst_cell_61_1 ( BL1, BLN1, WL61);
sram_cell_6t_3 inst_cell_61_0 ( BL0, BLN0, WL61);
sram_cell_6t_3 inst_cell_60_63 ( BL63, BLN63, WL60);
sram_cell_6t_3 inst_cell_60_62 ( BL62, BLN62, WL60);
sram_cell_6t_3 inst_cell_60_61 ( BL61, BLN61, WL60);
sram_cell_6t_3 inst_cell_60_60 ( BL60, BLN60, WL60);
sram_cell_6t_3 inst_cell_60_59 ( BL59, BLN59, WL60);
sram_cell_6t_3 inst_cell_60_58 ( BL58, BLN58, WL60);
sram_cell_6t_3 inst_cell_60_57 ( BL57, BLN57, WL60);
sram_cell_6t_3 inst_cell_60_56 ( BL56, BLN56, WL60);
sram_cell_6t_3 inst_cell_60_55 ( BL55, BLN55, WL60);
sram_cell_6t_3 inst_cell_60_54 ( BL54, BLN54, WL60);
sram_cell_6t_3 inst_cell_60_53 ( BL53, BLN53, WL60);
sram_cell_6t_3 inst_cell_60_52 ( BL52, BLN52, WL60);
sram_cell_6t_3 inst_cell_60_51 ( BL51, BLN51, WL60);
sram_cell_6t_3 inst_cell_60_50 ( BL50, BLN50, WL60);
sram_cell_6t_3 inst_cell_60_49 ( BL49, BLN49, WL60);
sram_cell_6t_3 inst_cell_60_48 ( BL48, BLN48, WL60);
sram_cell_6t_3 inst_cell_60_47 ( BL47, BLN47, WL60);
sram_cell_6t_3 inst_cell_60_46 ( BL46, BLN46, WL60);
sram_cell_6t_3 inst_cell_60_45 ( BL45, BLN45, WL60);
sram_cell_6t_3 inst_cell_60_44 ( BL44, BLN44, WL60);
sram_cell_6t_3 inst_cell_60_43 ( BL43, BLN43, WL60);
sram_cell_6t_3 inst_cell_60_42 ( BL42, BLN42, WL60);
sram_cell_6t_3 inst_cell_60_41 ( BL41, BLN41, WL60);
sram_cell_6t_3 inst_cell_60_31 ( BL31, BLN31, WL60);
sram_cell_6t_3 inst_cell_60_30 ( BL30, BLN30, WL60);
sram_cell_6t_3 inst_cell_60_29 ( BL29, BLN29, WL60);
sram_cell_6t_3 inst_cell_60_28 ( BL28, BLN28, WL60);
sram_cell_6t_3 inst_cell_60_27 ( BL27, BLN27, WL60);
sram_cell_6t_3 inst_cell_60_26 ( BL26, BLN26, WL60);
sram_cell_6t_3 inst_cell_60_25 ( BL25, BLN25, WL60);
sram_cell_6t_3 inst_cell_60_24 ( BL24, BLN24, WL60);
sram_cell_6t_3 inst_cell_60_40 ( BL40, BLN40, WL60);
sram_cell_6t_3 inst_cell_60_39 ( BL39, BLN39, WL60);
sram_cell_6t_3 inst_cell_60_38 ( BL38, BLN38, WL60);
sram_cell_6t_3 inst_cell_60_37 ( BL37, BLN37, WL60);
sram_cell_6t_3 inst_cell_60_36 ( BL36, BLN36, WL60);
sram_cell_6t_3 inst_cell_60_35 ( BL35, BLN35, WL60);
sram_cell_6t_3 inst_cell_60_34 ( BL34, BLN34, WL60);
sram_cell_6t_3 inst_cell_60_33 ( BL33, BLN33, WL60);
sram_cell_6t_3 inst_cell_60_32 ( BL32, BLN32, WL60);
sram_cell_6t_3 inst_cell_60_23 ( BL23, BLN23, WL60);
sram_cell_6t_3 inst_cell_60_22 ( BL22, BLN22, WL60);
sram_cell_6t_3 inst_cell_60_21 ( BL21, BLN21, WL60);
sram_cell_6t_3 inst_cell_60_20 ( BL20, BLN20, WL60);
sram_cell_6t_3 inst_cell_60_19 ( BL19, BLN19, WL60);
sram_cell_6t_3 inst_cell_60_18 ( BL18, BLN18, WL60);
sram_cell_6t_3 inst_cell_60_17 ( BL17, BLN17, WL60);
sram_cell_6t_3 inst_cell_60_16 ( BL16, BLN16, WL60);
sram_cell_6t_3 inst_cell_60_15 ( BL15, BLN15, WL60);
sram_cell_6t_3 inst_cell_60_14 ( BL14, BLN14, WL60);
sram_cell_6t_3 inst_cell_60_13 ( BL13, BLN13, WL60);
sram_cell_6t_3 inst_cell_60_12 ( BL12, BLN12, WL60);
sram_cell_6t_3 inst_cell_60_11 ( BL11, BLN11, WL60);
sram_cell_6t_3 inst_cell_60_10 ( BL10, BLN10, WL60);
sram_cell_6t_3 inst_cell_60_9 ( BL9, BLN9, WL60);
sram_cell_6t_3 inst_cell_60_8 ( BL8, BLN8, WL60);
sram_cell_6t_3 inst_cell_60_7 ( BL7, BLN7, WL60);
sram_cell_6t_3 inst_cell_60_6 ( BL6, BLN6, WL60);
sram_cell_6t_3 inst_cell_60_5 ( BL5, BLN5, WL60);
sram_cell_6t_3 inst_cell_60_4 ( BL4, BLN4, WL60);
sram_cell_6t_3 inst_cell_60_3 ( BL3, BLN3, WL60);
sram_cell_6t_3 inst_cell_60_2 ( BL2, BLN2, WL60);
sram_cell_6t_3 inst_cell_60_1 ( BL1, BLN1, WL60);
sram_cell_6t_3 inst_cell_60_0 ( BL0, BLN0, WL60);
sram_cell_6t_3 inst_cell_59_63 ( BL63, BLN63, WL59);
sram_cell_6t_3 inst_cell_59_62 ( BL62, BLN62, WL59);
sram_cell_6t_3 inst_cell_59_61 ( BL61, BLN61, WL59);
sram_cell_6t_3 inst_cell_59_60 ( BL60, BLN60, WL59);
sram_cell_6t_3 inst_cell_59_59 ( BL59, BLN59, WL59);
sram_cell_6t_3 inst_cell_59_58 ( BL58, BLN58, WL59);
sram_cell_6t_3 inst_cell_59_57 ( BL57, BLN57, WL59);
sram_cell_6t_3 inst_cell_59_56 ( BL56, BLN56, WL59);
sram_cell_6t_3 inst_cell_59_55 ( BL55, BLN55, WL59);
sram_cell_6t_3 inst_cell_59_54 ( BL54, BLN54, WL59);
sram_cell_6t_3 inst_cell_59_53 ( BL53, BLN53, WL59);
sram_cell_6t_3 inst_cell_59_52 ( BL52, BLN52, WL59);
sram_cell_6t_3 inst_cell_59_51 ( BL51, BLN51, WL59);
sram_cell_6t_3 inst_cell_59_50 ( BL50, BLN50, WL59);
sram_cell_6t_3 inst_cell_59_49 ( BL49, BLN49, WL59);
sram_cell_6t_3 inst_cell_59_48 ( BL48, BLN48, WL59);
sram_cell_6t_3 inst_cell_59_47 ( BL47, BLN47, WL59);
sram_cell_6t_3 inst_cell_59_46 ( BL46, BLN46, WL59);
sram_cell_6t_3 inst_cell_59_45 ( BL45, BLN45, WL59);
sram_cell_6t_3 inst_cell_59_44 ( BL44, BLN44, WL59);
sram_cell_6t_3 inst_cell_59_43 ( BL43, BLN43, WL59);
sram_cell_6t_3 inst_cell_59_42 ( BL42, BLN42, WL59);
sram_cell_6t_3 inst_cell_59_23 ( BL23, BLN23, WL59);
sram_cell_6t_3 inst_cell_59_22 ( BL22, BLN22, WL59);
sram_cell_6t_3 inst_cell_59_21 ( BL21, BLN21, WL59);
sram_cell_6t_3 inst_cell_59_20 ( BL20, BLN20, WL59);
sram_cell_6t_3 inst_cell_59_19 ( BL19, BLN19, WL59);
sram_cell_6t_3 inst_cell_59_18 ( BL18, BLN18, WL59);
sram_cell_6t_3 inst_cell_59_17 ( BL17, BLN17, WL59);
sram_cell_6t_3 inst_cell_59_16 ( BL16, BLN16, WL59);
sram_cell_6t_3 inst_cell_59_41 ( BL41, BLN41, WL59);
sram_cell_6t_3 inst_cell_59_40 ( BL40, BLN40, WL59);
sram_cell_6t_3 inst_cell_59_39 ( BL39, BLN39, WL59);
sram_cell_6t_3 inst_cell_59_38 ( BL38, BLN38, WL59);
sram_cell_6t_3 inst_cell_59_37 ( BL37, BLN37, WL59);
sram_cell_6t_3 inst_cell_59_36 ( BL36, BLN36, WL59);
sram_cell_6t_3 inst_cell_59_35 ( BL35, BLN35, WL59);
sram_cell_6t_3 inst_cell_59_34 ( BL34, BLN34, WL59);
sram_cell_6t_3 inst_cell_59_33 ( BL33, BLN33, WL59);
sram_cell_6t_3 inst_cell_59_32 ( BL32, BLN32, WL59);
sram_cell_6t_3 inst_cell_59_31 ( BL31, BLN31, WL59);
sram_cell_6t_3 inst_cell_59_30 ( BL30, BLN30, WL59);
sram_cell_6t_3 inst_cell_59_29 ( BL29, BLN29, WL59);
sram_cell_6t_3 inst_cell_59_28 ( BL28, BLN28, WL59);
sram_cell_6t_3 inst_cell_59_27 ( BL27, BLN27, WL59);
sram_cell_6t_3 inst_cell_59_26 ( BL26, BLN26, WL59);
sram_cell_6t_3 inst_cell_59_25 ( BL25, BLN25, WL59);
sram_cell_6t_3 inst_cell_59_24 ( BL24, BLN24, WL59);
sram_cell_6t_3 inst_cell_59_15 ( BL15, BLN15, WL59);
sram_cell_6t_3 inst_cell_59_14 ( BL14, BLN14, WL59);
sram_cell_6t_3 inst_cell_59_13 ( BL13, BLN13, WL59);
sram_cell_6t_3 inst_cell_59_12 ( BL12, BLN12, WL59);
sram_cell_6t_3 inst_cell_59_11 ( BL11, BLN11, WL59);
sram_cell_6t_3 inst_cell_59_10 ( BL10, BLN10, WL59);
sram_cell_6t_3 inst_cell_59_9 ( BL9, BLN9, WL59);
sram_cell_6t_3 inst_cell_59_8 ( BL8, BLN8, WL59);
sram_cell_6t_3 inst_cell_59_7 ( BL7, BLN7, WL59);
sram_cell_6t_3 inst_cell_59_6 ( BL6, BLN6, WL59);
sram_cell_6t_3 inst_cell_59_5 ( BL5, BLN5, WL59);
sram_cell_6t_3 inst_cell_59_4 ( BL4, BLN4, WL59);
sram_cell_6t_3 inst_cell_59_3 ( BL3, BLN3, WL59);
sram_cell_6t_3 inst_cell_59_2 ( BL2, BLN2, WL59);
sram_cell_6t_3 inst_cell_59_1 ( BL1, BLN1, WL59);
sram_cell_6t_3 inst_cell_59_0 ( BL0, BLN0, WL59);
sram_cell_6t_3 inst_cell_58_63 ( BL63, BLN63, WL58);
sram_cell_6t_3 inst_cell_58_62 ( BL62, BLN62, WL58);
sram_cell_6t_3 inst_cell_58_61 ( BL61, BLN61, WL58);
sram_cell_6t_3 inst_cell_58_60 ( BL60, BLN60, WL58);
sram_cell_6t_3 inst_cell_58_59 ( BL59, BLN59, WL58);
sram_cell_6t_3 inst_cell_58_58 ( BL58, BLN58, WL58);
sram_cell_6t_3 inst_cell_58_57 ( BL57, BLN57, WL58);
sram_cell_6t_3 inst_cell_58_56 ( BL56, BLN56, WL58);
sram_cell_6t_3 inst_cell_58_55 ( BL55, BLN55, WL58);
sram_cell_6t_3 inst_cell_58_54 ( BL54, BLN54, WL58);
sram_cell_6t_3 inst_cell_58_53 ( BL53, BLN53, WL58);
sram_cell_6t_3 inst_cell_58_52 ( BL52, BLN52, WL58);
sram_cell_6t_3 inst_cell_58_51 ( BL51, BLN51, WL58);
sram_cell_6t_3 inst_cell_58_50 ( BL50, BLN50, WL58);
sram_cell_6t_3 inst_cell_58_49 ( BL49, BLN49, WL58);
sram_cell_6t_3 inst_cell_58_48 ( BL48, BLN48, WL58);
sram_cell_6t_3 inst_cell_58_47 ( BL47, BLN47, WL58);
sram_cell_6t_3 inst_cell_58_46 ( BL46, BLN46, WL58);
sram_cell_6t_3 inst_cell_58_45 ( BL45, BLN45, WL58);
sram_cell_6t_3 inst_cell_58_44 ( BL44, BLN44, WL58);
sram_cell_6t_3 inst_cell_58_43 ( BL43, BLN43, WL58);
sram_cell_6t_3 inst_cell_58_15 ( BL15, BLN15, WL58);
sram_cell_6t_3 inst_cell_58_14 ( BL14, BLN14, WL58);
sram_cell_6t_3 inst_cell_58_13 ( BL13, BLN13, WL58);
sram_cell_6t_3 inst_cell_58_12 ( BL12, BLN12, WL58);
sram_cell_6t_3 inst_cell_58_11 ( BL11, BLN11, WL58);
sram_cell_6t_3 inst_cell_58_10 ( BL10, BLN10, WL58);
sram_cell_6t_3 inst_cell_58_9 ( BL9, BLN9, WL58);
sram_cell_6t_3 inst_cell_58_8 ( BL8, BLN8, WL58);
sram_cell_6t_3 inst_cell_58_42 ( BL42, BLN42, WL58);
sram_cell_6t_3 inst_cell_58_41 ( BL41, BLN41, WL58);
sram_cell_6t_3 inst_cell_58_40 ( BL40, BLN40, WL58);
sram_cell_6t_3 inst_cell_58_39 ( BL39, BLN39, WL58);
sram_cell_6t_3 inst_cell_58_38 ( BL38, BLN38, WL58);
sram_cell_6t_3 inst_cell_58_37 ( BL37, BLN37, WL58);
sram_cell_6t_3 inst_cell_58_36 ( BL36, BLN36, WL58);
sram_cell_6t_3 inst_cell_58_35 ( BL35, BLN35, WL58);
sram_cell_6t_3 inst_cell_58_34 ( BL34, BLN34, WL58);
sram_cell_6t_3 inst_cell_58_33 ( BL33, BLN33, WL58);
sram_cell_6t_3 inst_cell_58_32 ( BL32, BLN32, WL58);
sram_cell_6t_3 inst_cell_58_31 ( BL31, BLN31, WL58);
sram_cell_6t_3 inst_cell_58_30 ( BL30, BLN30, WL58);
sram_cell_6t_3 inst_cell_58_29 ( BL29, BLN29, WL58);
sram_cell_6t_3 inst_cell_58_28 ( BL28, BLN28, WL58);
sram_cell_6t_3 inst_cell_58_27 ( BL27, BLN27, WL58);
sram_cell_6t_3 inst_cell_58_26 ( BL26, BLN26, WL58);
sram_cell_6t_3 inst_cell_58_25 ( BL25, BLN25, WL58);
sram_cell_6t_3 inst_cell_58_24 ( BL24, BLN24, WL58);
sram_cell_6t_3 inst_cell_58_23 ( BL23, BLN23, WL58);
sram_cell_6t_3 inst_cell_58_22 ( BL22, BLN22, WL58);
sram_cell_6t_3 inst_cell_58_21 ( BL21, BLN21, WL58);
sram_cell_6t_3 inst_cell_58_20 ( BL20, BLN20, WL58);
sram_cell_6t_3 inst_cell_58_19 ( BL19, BLN19, WL58);
sram_cell_6t_3 inst_cell_58_18 ( BL18, BLN18, WL58);
sram_cell_6t_3 inst_cell_58_17 ( BL17, BLN17, WL58);
sram_cell_6t_3 inst_cell_58_16 ( BL16, BLN16, WL58);
sram_cell_6t_3 inst_cell_58_7 ( BL7, BLN7, WL58);
sram_cell_6t_3 inst_cell_58_6 ( BL6, BLN6, WL58);
sram_cell_6t_3 inst_cell_58_5 ( BL5, BLN5, WL58);
sram_cell_6t_3 inst_cell_58_4 ( BL4, BLN4, WL58);
sram_cell_6t_3 inst_cell_58_3 ( BL3, BLN3, WL58);
sram_cell_6t_3 inst_cell_58_2 ( BL2, BLN2, WL58);
sram_cell_6t_3 inst_cell_58_1 ( BL1, BLN1, WL58);
sram_cell_6t_3 inst_cell_58_0 ( BL0, BLN0, WL58);
sram_cell_6t_3 inst_cell_57_63 ( BL63, BLN63, WL57);
sram_cell_6t_3 inst_cell_57_62 ( BL62, BLN62, WL57);
sram_cell_6t_3 inst_cell_57_61 ( BL61, BLN61, WL57);
sram_cell_6t_3 inst_cell_57_60 ( BL60, BLN60, WL57);
sram_cell_6t_3 inst_cell_57_59 ( BL59, BLN59, WL57);
sram_cell_6t_3 inst_cell_57_58 ( BL58, BLN58, WL57);
sram_cell_6t_3 inst_cell_57_57 ( BL57, BLN57, WL57);
sram_cell_6t_3 inst_cell_57_56 ( BL56, BLN56, WL57);
sram_cell_6t_3 inst_cell_57_55 ( BL55, BLN55, WL57);
sram_cell_6t_3 inst_cell_57_54 ( BL54, BLN54, WL57);
sram_cell_6t_3 inst_cell_57_53 ( BL53, BLN53, WL57);
sram_cell_6t_3 inst_cell_57_52 ( BL52, BLN52, WL57);
sram_cell_6t_3 inst_cell_57_51 ( BL51, BLN51, WL57);
sram_cell_6t_3 inst_cell_57_50 ( BL50, BLN50, WL57);
sram_cell_6t_3 inst_cell_57_49 ( BL49, BLN49, WL57);
sram_cell_6t_3 inst_cell_57_48 ( BL48, BLN48, WL57);
sram_cell_6t_3 inst_cell_57_47 ( BL47, BLN47, WL57);
sram_cell_6t_3 inst_cell_57_46 ( BL46, BLN46, WL57);
sram_cell_6t_3 inst_cell_57_45 ( BL45, BLN45, WL57);
sram_cell_6t_3 inst_cell_57_44 ( BL44, BLN44, WL57);
sram_cell_6t_3 inst_cell_57_7 ( BL7, BLN7, WL57);
sram_cell_6t_3 inst_cell_57_6 ( BL6, BLN6, WL57);
sram_cell_6t_3 inst_cell_57_5 ( BL5, BLN5, WL57);
sram_cell_6t_3 inst_cell_57_4 ( BL4, BLN4, WL57);
sram_cell_6t_3 inst_cell_57_3 ( BL3, BLN3, WL57);
sram_cell_6t_3 inst_cell_57_2 ( BL2, BLN2, WL57);
sram_cell_6t_3 inst_cell_57_1 ( BL1, BLN1, WL57);
sram_cell_6t_3 inst_cell_57_0 ( BL0, BLN0, WL57);
sram_cell_6t_3 inst_cell_57_43 ( BL43, BLN43, WL57);
sram_cell_6t_3 inst_cell_57_42 ( BL42, BLN42, WL57);
sram_cell_6t_3 inst_cell_57_41 ( BL41, BLN41, WL57);
sram_cell_6t_3 inst_cell_57_40 ( BL40, BLN40, WL57);
sram_cell_6t_3 inst_cell_57_39 ( BL39, BLN39, WL57);
sram_cell_6t_3 inst_cell_57_38 ( BL38, BLN38, WL57);
sram_cell_6t_3 inst_cell_57_37 ( BL37, BLN37, WL57);
sram_cell_6t_3 inst_cell_57_36 ( BL36, BLN36, WL57);
sram_cell_6t_3 inst_cell_57_35 ( BL35, BLN35, WL57);
sram_cell_6t_3 inst_cell_57_34 ( BL34, BLN34, WL57);
sram_cell_6t_3 inst_cell_57_33 ( BL33, BLN33, WL57);
sram_cell_6t_3 inst_cell_57_32 ( BL32, BLN32, WL57);
sram_cell_6t_3 inst_cell_57_31 ( BL31, BLN31, WL57);
sram_cell_6t_3 inst_cell_57_30 ( BL30, BLN30, WL57);
sram_cell_6t_3 inst_cell_57_29 ( BL29, BLN29, WL57);
sram_cell_6t_3 inst_cell_57_28 ( BL28, BLN28, WL57);
sram_cell_6t_3 inst_cell_57_27 ( BL27, BLN27, WL57);
sram_cell_6t_3 inst_cell_57_26 ( BL26, BLN26, WL57);
sram_cell_6t_3 inst_cell_57_25 ( BL25, BLN25, WL57);
sram_cell_6t_3 inst_cell_57_24 ( BL24, BLN24, WL57);
sram_cell_6t_3 inst_cell_57_23 ( BL23, BLN23, WL57);
sram_cell_6t_3 inst_cell_57_22 ( BL22, BLN22, WL57);
sram_cell_6t_3 inst_cell_57_21 ( BL21, BLN21, WL57);
sram_cell_6t_3 inst_cell_57_20 ( BL20, BLN20, WL57);
sram_cell_6t_3 inst_cell_57_19 ( BL19, BLN19, WL57);
sram_cell_6t_3 inst_cell_57_18 ( BL18, BLN18, WL57);
sram_cell_6t_3 inst_cell_57_17 ( BL17, BLN17, WL57);
sram_cell_6t_3 inst_cell_57_16 ( BL16, BLN16, WL57);
sram_cell_6t_3 inst_cell_57_15 ( BL15, BLN15, WL57);
sram_cell_6t_3 inst_cell_57_14 ( BL14, BLN14, WL57);
sram_cell_6t_3 inst_cell_57_13 ( BL13, BLN13, WL57);
sram_cell_6t_3 inst_cell_57_12 ( BL12, BLN12, WL57);
sram_cell_6t_3 inst_cell_57_11 ( BL11, BLN11, WL57);
sram_cell_6t_3 inst_cell_57_10 ( BL10, BLN10, WL57);
sram_cell_6t_3 inst_cell_57_9 ( BL9, BLN9, WL57);
sram_cell_6t_3 inst_cell_57_8 ( BL8, BLN8, WL57);
sram_cell_6t_3 inst_cell_56_63 ( BL63, BLN63, WL56);
sram_cell_6t_3 inst_cell_56_62 ( BL62, BLN62, WL56);
sram_cell_6t_3 inst_cell_56_61 ( BL61, BLN61, WL56);
sram_cell_6t_3 inst_cell_56_60 ( BL60, BLN60, WL56);
sram_cell_6t_3 inst_cell_56_59 ( BL59, BLN59, WL56);
sram_cell_6t_3 inst_cell_56_58 ( BL58, BLN58, WL56);
sram_cell_6t_3 inst_cell_56_57 ( BL57, BLN57, WL56);
sram_cell_6t_3 inst_cell_56_56 ( BL56, BLN56, WL56);
sram_cell_6t_3 inst_cell_56_55 ( BL55, BLN55, WL56);
sram_cell_6t_3 inst_cell_56_54 ( BL54, BLN54, WL56);
sram_cell_6t_3 inst_cell_56_53 ( BL53, BLN53, WL56);
sram_cell_6t_3 inst_cell_56_52 ( BL52, BLN52, WL56);
sram_cell_6t_3 inst_cell_56_51 ( BL51, BLN51, WL56);
sram_cell_6t_3 inst_cell_56_50 ( BL50, BLN50, WL56);
sram_cell_6t_3 inst_cell_56_49 ( BL49, BLN49, WL56);
sram_cell_6t_3 inst_cell_56_48 ( BL48, BLN48, WL56);
sram_cell_6t_3 inst_cell_56_47 ( BL47, BLN47, WL56);
sram_cell_6t_3 inst_cell_56_46 ( BL46, BLN46, WL56);
sram_cell_6t_3 inst_cell_56_45 ( BL45, BLN45, WL56);
sram_cell_6t_3 inst_cell_56_44 ( BL44, BLN44, WL56);
sram_cell_6t_3 inst_cell_56_43 ( BL43, BLN43, WL56);
sram_cell_6t_3 inst_cell_56_42 ( BL42, BLN42, WL56);
sram_cell_6t_3 inst_cell_56_41 ( BL41, BLN41, WL56);
sram_cell_6t_3 inst_cell_56_40 ( BL40, BLN40, WL56);
sram_cell_6t_3 inst_cell_56_39 ( BL39, BLN39, WL56);
sram_cell_6t_3 inst_cell_56_38 ( BL38, BLN38, WL56);
sram_cell_6t_3 inst_cell_56_37 ( BL37, BLN37, WL56);
sram_cell_6t_3 inst_cell_56_36 ( BL36, BLN36, WL56);
sram_cell_6t_3 inst_cell_56_35 ( BL35, BLN35, WL56);
sram_cell_6t_3 inst_cell_56_34 ( BL34, BLN34, WL56);
sram_cell_6t_3 inst_cell_56_33 ( BL33, BLN33, WL56);
sram_cell_6t_3 inst_cell_56_32 ( BL32, BLN32, WL56);
sram_cell_6t_3 inst_cell_56_31 ( BL31, BLN31, WL56);
sram_cell_6t_3 inst_cell_56_30 ( BL30, BLN30, WL56);
sram_cell_6t_3 inst_cell_56_29 ( BL29, BLN29, WL56);
sram_cell_6t_3 inst_cell_56_28 ( BL28, BLN28, WL56);
sram_cell_6t_3 inst_cell_56_27 ( BL27, BLN27, WL56);
sram_cell_6t_3 inst_cell_56_26 ( BL26, BLN26, WL56);
sram_cell_6t_3 inst_cell_56_25 ( BL25, BLN25, WL56);
sram_cell_6t_3 inst_cell_56_24 ( BL24, BLN24, WL56);
sram_cell_6t_3 inst_cell_56_23 ( BL23, BLN23, WL56);
sram_cell_6t_3 inst_cell_56_22 ( BL22, BLN22, WL56);
sram_cell_6t_3 inst_cell_56_21 ( BL21, BLN21, WL56);
sram_cell_6t_3 inst_cell_56_20 ( BL20, BLN20, WL56);
sram_cell_6t_3 inst_cell_56_19 ( BL19, BLN19, WL56);
sram_cell_6t_3 inst_cell_56_18 ( BL18, BLN18, WL56);
sram_cell_6t_3 inst_cell_56_17 ( BL17, BLN17, WL56);
sram_cell_6t_3 inst_cell_56_16 ( BL16, BLN16, WL56);
sram_cell_6t_3 inst_cell_56_15 ( BL15, BLN15, WL56);
sram_cell_6t_3 inst_cell_56_14 ( BL14, BLN14, WL56);
sram_cell_6t_3 inst_cell_56_13 ( BL13, BLN13, WL56);
sram_cell_6t_3 inst_cell_56_12 ( BL12, BLN12, WL56);
sram_cell_6t_3 inst_cell_56_11 ( BL11, BLN11, WL56);
sram_cell_6t_3 inst_cell_56_10 ( BL10, BLN10, WL56);
sram_cell_6t_3 inst_cell_56_9 ( BL9, BLN9, WL56);
sram_cell_6t_3 inst_cell_56_8 ( BL8, BLN8, WL56);
sram_cell_6t_3 inst_cell_56_7 ( BL7, BLN7, WL56);
sram_cell_6t_3 inst_cell_56_6 ( BL6, BLN6, WL56);
sram_cell_6t_3 inst_cell_56_5 ( BL5, BLN5, WL56);
sram_cell_6t_3 inst_cell_56_4 ( BL4, BLN4, WL56);
sram_cell_6t_3 inst_cell_56_3 ( BL3, BLN3, WL56);
sram_cell_6t_3 inst_cell_56_2 ( BL2, BLN2, WL56);
sram_cell_6t_3 inst_cell_56_1 ( BL1, BLN1, WL56);
sram_cell_6t_3 inst_cell_56_0 ( BL0, BLN0, WL56);
sram_cell_6t_3 inst_cell_55_63 ( BL63, BLN63, WL55);
sram_cell_6t_3 inst_cell_55_62 ( BL62, BLN62, WL55);
sram_cell_6t_3 inst_cell_55_61 ( BL61, BLN61, WL55);
sram_cell_6t_3 inst_cell_55_60 ( BL60, BLN60, WL55);
sram_cell_6t_3 inst_cell_55_59 ( BL59, BLN59, WL55);
sram_cell_6t_3 inst_cell_55_58 ( BL58, BLN58, WL55);
sram_cell_6t_3 inst_cell_55_57 ( BL57, BLN57, WL55);
sram_cell_6t_3 inst_cell_55_56 ( BL56, BLN56, WL55);
sram_cell_6t_3 inst_cell_55_55 ( BL55, BLN55, WL55);
sram_cell_6t_3 inst_cell_55_54 ( BL54, BLN54, WL55);
sram_cell_6t_3 inst_cell_55_53 ( BL53, BLN53, WL55);
sram_cell_6t_3 inst_cell_55_52 ( BL52, BLN52, WL55);
sram_cell_6t_3 inst_cell_55_51 ( BL51, BLN51, WL55);
sram_cell_6t_3 inst_cell_55_50 ( BL50, BLN50, WL55);
sram_cell_6t_3 inst_cell_55_49 ( BL49, BLN49, WL55);
sram_cell_6t_3 inst_cell_55_48 ( BL48, BLN48, WL55);
sram_cell_6t_3 inst_cell_55_47 ( BL47, BLN47, WL55);
sram_cell_6t_3 inst_cell_55_46 ( BL46, BLN46, WL55);
sram_cell_6t_3 inst_cell_55_45 ( BL45, BLN45, WL55);
sram_cell_6t_3 inst_cell_55_44 ( BL44, BLN44, WL55);
sram_cell_6t_3 inst_cell_55_43 ( BL43, BLN43, WL55);
sram_cell_6t_3 inst_cell_55_42 ( BL42, BLN42, WL55);
sram_cell_6t_3 inst_cell_55_41 ( BL41, BLN41, WL55);
sram_cell_6t_3 inst_cell_55_40 ( BL40, BLN40, WL55);
sram_cell_6t_3 inst_cell_55_39 ( BL39, BLN39, WL55);
sram_cell_6t_3 inst_cell_55_38 ( BL38, BLN38, WL55);
sram_cell_6t_3 inst_cell_55_37 ( BL37, BLN37, WL55);
sram_cell_6t_3 inst_cell_55_36 ( BL36, BLN36, WL55);
sram_cell_6t_3 inst_cell_55_35 ( BL35, BLN35, WL55);
sram_cell_6t_3 inst_cell_55_34 ( BL34, BLN34, WL55);
sram_cell_6t_3 inst_cell_55_33 ( BL33, BLN33, WL55);
sram_cell_6t_3 inst_cell_55_32 ( BL32, BLN32, WL55);
sram_cell_6t_3 inst_cell_55_31 ( BL31, BLN31, WL55);
sram_cell_6t_3 inst_cell_55_30 ( BL30, BLN30, WL55);
sram_cell_6t_3 inst_cell_55_29 ( BL29, BLN29, WL55);
sram_cell_6t_3 inst_cell_55_28 ( BL28, BLN28, WL55);
sram_cell_6t_3 inst_cell_55_27 ( BL27, BLN27, WL55);
sram_cell_6t_3 inst_cell_55_26 ( BL26, BLN26, WL55);
sram_cell_6t_3 inst_cell_55_25 ( BL25, BLN25, WL55);
sram_cell_6t_3 inst_cell_55_24 ( BL24, BLN24, WL55);
sram_cell_6t_3 inst_cell_55_23 ( BL23, BLN23, WL55);
sram_cell_6t_3 inst_cell_55_22 ( BL22, BLN22, WL55);
sram_cell_6t_3 inst_cell_55_21 ( BL21, BLN21, WL55);
sram_cell_6t_3 inst_cell_55_20 ( BL20, BLN20, WL55);
sram_cell_6t_3 inst_cell_55_19 ( BL19, BLN19, WL55);
sram_cell_6t_3 inst_cell_55_18 ( BL18, BLN18, WL55);
sram_cell_6t_3 inst_cell_55_17 ( BL17, BLN17, WL55);
sram_cell_6t_3 inst_cell_55_16 ( BL16, BLN16, WL55);
sram_cell_6t_3 inst_cell_55_15 ( BL15, BLN15, WL55);
sram_cell_6t_3 inst_cell_55_14 ( BL14, BLN14, WL55);
sram_cell_6t_3 inst_cell_55_13 ( BL13, BLN13, WL55);
sram_cell_6t_3 inst_cell_55_12 ( BL12, BLN12, WL55);
sram_cell_6t_3 inst_cell_55_11 ( BL11, BLN11, WL55);
sram_cell_6t_3 inst_cell_55_10 ( BL10, BLN10, WL55);
sram_cell_6t_3 inst_cell_55_9 ( BL9, BLN9, WL55);
sram_cell_6t_3 inst_cell_55_8 ( BL8, BLN8, WL55);
sram_cell_6t_3 inst_cell_55_7 ( BL7, BLN7, WL55);
sram_cell_6t_3 inst_cell_55_6 ( BL6, BLN6, WL55);
sram_cell_6t_3 inst_cell_55_5 ( BL5, BLN5, WL55);
sram_cell_6t_3 inst_cell_55_4 ( BL4, BLN4, WL55);
sram_cell_6t_3 inst_cell_55_3 ( BL3, BLN3, WL55);
sram_cell_6t_3 inst_cell_55_2 ( BL2, BLN2, WL55);
sram_cell_6t_3 inst_cell_55_1 ( BL1, BLN1, WL55);
sram_cell_6t_3 inst_cell_55_0 ( BL0, BLN0, WL55);
sram_cell_6t_3 inst_cell_54_63 ( BL63, BLN63, WL54);
sram_cell_6t_3 inst_cell_54_62 ( BL62, BLN62, WL54);
sram_cell_6t_3 inst_cell_54_61 ( BL61, BLN61, WL54);
sram_cell_6t_3 inst_cell_54_60 ( BL60, BLN60, WL54);
sram_cell_6t_3 inst_cell_54_59 ( BL59, BLN59, WL54);
sram_cell_6t_3 inst_cell_54_58 ( BL58, BLN58, WL54);
sram_cell_6t_3 inst_cell_54_57 ( BL57, BLN57, WL54);
sram_cell_6t_3 inst_cell_54_56 ( BL56, BLN56, WL54);
sram_cell_6t_3 inst_cell_54_55 ( BL55, BLN55, WL54);
sram_cell_6t_3 inst_cell_54_54 ( BL54, BLN54, WL54);
sram_cell_6t_3 inst_cell_54_53 ( BL53, BLN53, WL54);
sram_cell_6t_3 inst_cell_54_52 ( BL52, BLN52, WL54);
sram_cell_6t_3 inst_cell_54_51 ( BL51, BLN51, WL54);
sram_cell_6t_3 inst_cell_54_50 ( BL50, BLN50, WL54);
sram_cell_6t_3 inst_cell_54_49 ( BL49, BLN49, WL54);
sram_cell_6t_3 inst_cell_54_48 ( BL48, BLN48, WL54);
sram_cell_6t_3 inst_cell_54_47 ( BL47, BLN47, WL54);
sram_cell_6t_3 inst_cell_54_46 ( BL46, BLN46, WL54);
sram_cell_6t_3 inst_cell_54_45 ( BL45, BLN45, WL54);
sram_cell_6t_3 inst_cell_54_44 ( BL44, BLN44, WL54);
sram_cell_6t_3 inst_cell_54_43 ( BL43, BLN43, WL54);
sram_cell_6t_3 inst_cell_54_42 ( BL42, BLN42, WL54);
sram_cell_6t_3 inst_cell_54_41 ( BL41, BLN41, WL54);
sram_cell_6t_3 inst_cell_54_40 ( BL40, BLN40, WL54);
sram_cell_6t_3 inst_cell_54_39 ( BL39, BLN39, WL54);
sram_cell_6t_3 inst_cell_54_38 ( BL38, BLN38, WL54);
sram_cell_6t_3 inst_cell_54_37 ( BL37, BLN37, WL54);
sram_cell_6t_3 inst_cell_54_36 ( BL36, BLN36, WL54);
sram_cell_6t_3 inst_cell_54_35 ( BL35, BLN35, WL54);
sram_cell_6t_3 inst_cell_54_34 ( BL34, BLN34, WL54);
sram_cell_6t_3 inst_cell_54_33 ( BL33, BLN33, WL54);
sram_cell_6t_3 inst_cell_54_32 ( BL32, BLN32, WL54);
sram_cell_6t_3 inst_cell_54_31 ( BL31, BLN31, WL54);
sram_cell_6t_3 inst_cell_54_30 ( BL30, BLN30, WL54);
sram_cell_6t_3 inst_cell_54_29 ( BL29, BLN29, WL54);
sram_cell_6t_3 inst_cell_54_28 ( BL28, BLN28, WL54);
sram_cell_6t_3 inst_cell_54_27 ( BL27, BLN27, WL54);
sram_cell_6t_3 inst_cell_54_26 ( BL26, BLN26, WL54);
sram_cell_6t_3 inst_cell_54_25 ( BL25, BLN25, WL54);
sram_cell_6t_3 inst_cell_54_24 ( BL24, BLN24, WL54);
sram_cell_6t_3 inst_cell_54_23 ( BL23, BLN23, WL54);
sram_cell_6t_3 inst_cell_54_22 ( BL22, BLN22, WL54);
sram_cell_6t_3 inst_cell_54_21 ( BL21, BLN21, WL54);
sram_cell_6t_3 inst_cell_54_20 ( BL20, BLN20, WL54);
sram_cell_6t_3 inst_cell_54_19 ( BL19, BLN19, WL54);
sram_cell_6t_3 inst_cell_54_18 ( BL18, BLN18, WL54);
sram_cell_6t_3 inst_cell_54_17 ( BL17, BLN17, WL54);
sram_cell_6t_3 inst_cell_54_16 ( BL16, BLN16, WL54);
sram_cell_6t_3 inst_cell_54_15 ( BL15, BLN15, WL54);
sram_cell_6t_3 inst_cell_54_14 ( BL14, BLN14, WL54);
sram_cell_6t_3 inst_cell_54_13 ( BL13, BLN13, WL54);
sram_cell_6t_3 inst_cell_54_12 ( BL12, BLN12, WL54);
sram_cell_6t_3 inst_cell_54_11 ( BL11, BLN11, WL54);
sram_cell_6t_3 inst_cell_54_10 ( BL10, BLN10, WL54);
sram_cell_6t_3 inst_cell_54_9 ( BL9, BLN9, WL54);
sram_cell_6t_3 inst_cell_54_8 ( BL8, BLN8, WL54);
sram_cell_6t_3 inst_cell_54_7 ( BL7, BLN7, WL54);
sram_cell_6t_3 inst_cell_54_6 ( BL6, BLN6, WL54);
sram_cell_6t_3 inst_cell_54_5 ( BL5, BLN5, WL54);
sram_cell_6t_3 inst_cell_54_4 ( BL4, BLN4, WL54);
sram_cell_6t_3 inst_cell_54_3 ( BL3, BLN3, WL54);
sram_cell_6t_3 inst_cell_54_2 ( BL2, BLN2, WL54);
sram_cell_6t_3 inst_cell_54_1 ( BL1, BLN1, WL54);
sram_cell_6t_3 inst_cell_54_0 ( BL0, BLN0, WL54);
sram_cell_6t_3 inst_cell_53_63 ( BL63, BLN63, WL53);
sram_cell_6t_3 inst_cell_53_62 ( BL62, BLN62, WL53);
sram_cell_6t_3 inst_cell_53_61 ( BL61, BLN61, WL53);
sram_cell_6t_3 inst_cell_53_60 ( BL60, BLN60, WL53);
sram_cell_6t_3 inst_cell_53_59 ( BL59, BLN59, WL53);
sram_cell_6t_3 inst_cell_53_58 ( BL58, BLN58, WL53);
sram_cell_6t_3 inst_cell_53_57 ( BL57, BLN57, WL53);
sram_cell_6t_3 inst_cell_53_56 ( BL56, BLN56, WL53);
sram_cell_6t_3 inst_cell_53_55 ( BL55, BLN55, WL53);
sram_cell_6t_3 inst_cell_53_54 ( BL54, BLN54, WL53);
sram_cell_6t_3 inst_cell_53_53 ( BL53, BLN53, WL53);
sram_cell_6t_3 inst_cell_53_52 ( BL52, BLN52, WL53);
sram_cell_6t_3 inst_cell_53_51 ( BL51, BLN51, WL53);
sram_cell_6t_3 inst_cell_53_50 ( BL50, BLN50, WL53);
sram_cell_6t_3 inst_cell_53_49 ( BL49, BLN49, WL53);
sram_cell_6t_3 inst_cell_53_48 ( BL48, BLN48, WL53);
sram_cell_6t_3 inst_cell_53_47 ( BL47, BLN47, WL53);
sram_cell_6t_3 inst_cell_53_46 ( BL46, BLN46, WL53);
sram_cell_6t_3 inst_cell_53_45 ( BL45, BLN45, WL53);
sram_cell_6t_3 inst_cell_53_44 ( BL44, BLN44, WL53);
sram_cell_6t_3 inst_cell_53_43 ( BL43, BLN43, WL53);
sram_cell_6t_3 inst_cell_53_42 ( BL42, BLN42, WL53);
sram_cell_6t_3 inst_cell_53_41 ( BL41, BLN41, WL53);
sram_cell_6t_3 inst_cell_53_40 ( BL40, BLN40, WL53);
sram_cell_6t_3 inst_cell_53_39 ( BL39, BLN39, WL53);
sram_cell_6t_3 inst_cell_53_38 ( BL38, BLN38, WL53);
sram_cell_6t_3 inst_cell_53_37 ( BL37, BLN37, WL53);
sram_cell_6t_3 inst_cell_53_36 ( BL36, BLN36, WL53);
sram_cell_6t_3 inst_cell_53_35 ( BL35, BLN35, WL53);
sram_cell_6t_3 inst_cell_53_34 ( BL34, BLN34, WL53);
sram_cell_6t_3 inst_cell_53_33 ( BL33, BLN33, WL53);
sram_cell_6t_3 inst_cell_53_32 ( BL32, BLN32, WL53);
sram_cell_6t_3 inst_cell_53_31 ( BL31, BLN31, WL53);
sram_cell_6t_3 inst_cell_53_30 ( BL30, BLN30, WL53);
sram_cell_6t_3 inst_cell_53_29 ( BL29, BLN29, WL53);
sram_cell_6t_3 inst_cell_53_28 ( BL28, BLN28, WL53);
sram_cell_6t_3 inst_cell_53_27 ( BL27, BLN27, WL53);
sram_cell_6t_3 inst_cell_53_26 ( BL26, BLN26, WL53);
sram_cell_6t_3 inst_cell_53_25 ( BL25, BLN25, WL53);
sram_cell_6t_3 inst_cell_53_24 ( BL24, BLN24, WL53);
sram_cell_6t_3 inst_cell_53_23 ( BL23, BLN23, WL53);
sram_cell_6t_3 inst_cell_53_22 ( BL22, BLN22, WL53);
sram_cell_6t_3 inst_cell_53_21 ( BL21, BLN21, WL53);
sram_cell_6t_3 inst_cell_53_20 ( BL20, BLN20, WL53);
sram_cell_6t_3 inst_cell_53_19 ( BL19, BLN19, WL53);
sram_cell_6t_3 inst_cell_53_18 ( BL18, BLN18, WL53);
sram_cell_6t_3 inst_cell_53_17 ( BL17, BLN17, WL53);
sram_cell_6t_3 inst_cell_53_16 ( BL16, BLN16, WL53);
sram_cell_6t_3 inst_cell_53_15 ( BL15, BLN15, WL53);
sram_cell_6t_3 inst_cell_53_14 ( BL14, BLN14, WL53);
sram_cell_6t_3 inst_cell_53_13 ( BL13, BLN13, WL53);
sram_cell_6t_3 inst_cell_53_12 ( BL12, BLN12, WL53);
sram_cell_6t_3 inst_cell_53_11 ( BL11, BLN11, WL53);
sram_cell_6t_3 inst_cell_53_10 ( BL10, BLN10, WL53);
sram_cell_6t_3 inst_cell_53_9 ( BL9, BLN9, WL53);
sram_cell_6t_3 inst_cell_53_8 ( BL8, BLN8, WL53);
sram_cell_6t_3 inst_cell_53_7 ( BL7, BLN7, WL53);
sram_cell_6t_3 inst_cell_53_6 ( BL6, BLN6, WL53);
sram_cell_6t_3 inst_cell_53_5 ( BL5, BLN5, WL53);
sram_cell_6t_3 inst_cell_53_4 ( BL4, BLN4, WL53);
sram_cell_6t_3 inst_cell_53_3 ( BL3, BLN3, WL53);
sram_cell_6t_3 inst_cell_53_2 ( BL2, BLN2, WL53);
sram_cell_6t_3 inst_cell_53_1 ( BL1, BLN1, WL53);
sram_cell_6t_3 inst_cell_53_0 ( BL0, BLN0, WL53);
sram_cell_6t_3 inst_cell_52_63 ( BL63, BLN63, WL52);
sram_cell_6t_3 inst_cell_52_62 ( BL62, BLN62, WL52);
sram_cell_6t_3 inst_cell_52_61 ( BL61, BLN61, WL52);
sram_cell_6t_3 inst_cell_52_60 ( BL60, BLN60, WL52);
sram_cell_6t_3 inst_cell_52_59 ( BL59, BLN59, WL52);
sram_cell_6t_3 inst_cell_52_58 ( BL58, BLN58, WL52);
sram_cell_6t_3 inst_cell_52_57 ( BL57, BLN57, WL52);
sram_cell_6t_3 inst_cell_52_56 ( BL56, BLN56, WL52);
sram_cell_6t_3 inst_cell_52_55 ( BL55, BLN55, WL52);
sram_cell_6t_3 inst_cell_52_54 ( BL54, BLN54, WL52);
sram_cell_6t_3 inst_cell_52_53 ( BL53, BLN53, WL52);
sram_cell_6t_3 inst_cell_52_52 ( BL52, BLN52, WL52);
sram_cell_6t_3 inst_cell_52_51 ( BL51, BLN51, WL52);
sram_cell_6t_3 inst_cell_52_50 ( BL50, BLN50, WL52);
sram_cell_6t_3 inst_cell_52_49 ( BL49, BLN49, WL52);
sram_cell_6t_3 inst_cell_52_48 ( BL48, BLN48, WL52);
sram_cell_6t_3 inst_cell_52_47 ( BL47, BLN47, WL52);
sram_cell_6t_3 inst_cell_52_46 ( BL46, BLN46, WL52);
sram_cell_6t_3 inst_cell_52_45 ( BL45, BLN45, WL52);
sram_cell_6t_3 inst_cell_52_44 ( BL44, BLN44, WL52);
sram_cell_6t_3 inst_cell_52_43 ( BL43, BLN43, WL52);
sram_cell_6t_3 inst_cell_52_42 ( BL42, BLN42, WL52);
sram_cell_6t_3 inst_cell_52_41 ( BL41, BLN41, WL52);
sram_cell_6t_3 inst_cell_52_40 ( BL40, BLN40, WL52);
sram_cell_6t_3 inst_cell_52_39 ( BL39, BLN39, WL52);
sram_cell_6t_3 inst_cell_52_38 ( BL38, BLN38, WL52);
sram_cell_6t_3 inst_cell_52_37 ( BL37, BLN37, WL52);
sram_cell_6t_3 inst_cell_52_36 ( BL36, BLN36, WL52);
sram_cell_6t_3 inst_cell_52_35 ( BL35, BLN35, WL52);
sram_cell_6t_3 inst_cell_52_34 ( BL34, BLN34, WL52);
sram_cell_6t_3 inst_cell_52_33 ( BL33, BLN33, WL52);
sram_cell_6t_3 inst_cell_52_32 ( BL32, BLN32, WL52);
sram_cell_6t_3 inst_cell_52_31 ( BL31, BLN31, WL52);
sram_cell_6t_3 inst_cell_52_30 ( BL30, BLN30, WL52);
sram_cell_6t_3 inst_cell_52_29 ( BL29, BLN29, WL52);
sram_cell_6t_3 inst_cell_52_28 ( BL28, BLN28, WL52);
sram_cell_6t_3 inst_cell_52_27 ( BL27, BLN27, WL52);
sram_cell_6t_3 inst_cell_52_26 ( BL26, BLN26, WL52);
sram_cell_6t_3 inst_cell_52_25 ( BL25, BLN25, WL52);
sram_cell_6t_3 inst_cell_52_24 ( BL24, BLN24, WL52);
sram_cell_6t_3 inst_cell_52_23 ( BL23, BLN23, WL52);
sram_cell_6t_3 inst_cell_52_22 ( BL22, BLN22, WL52);
sram_cell_6t_3 inst_cell_52_21 ( BL21, BLN21, WL52);
sram_cell_6t_3 inst_cell_52_20 ( BL20, BLN20, WL52);
sram_cell_6t_3 inst_cell_52_19 ( BL19, BLN19, WL52);
sram_cell_6t_3 inst_cell_52_18 ( BL18, BLN18, WL52);
sram_cell_6t_3 inst_cell_52_17 ( BL17, BLN17, WL52);
sram_cell_6t_3 inst_cell_52_16 ( BL16, BLN16, WL52);
sram_cell_6t_3 inst_cell_52_15 ( BL15, BLN15, WL52);
sram_cell_6t_3 inst_cell_52_14 ( BL14, BLN14, WL52);
sram_cell_6t_3 inst_cell_52_13 ( BL13, BLN13, WL52);
sram_cell_6t_3 inst_cell_52_12 ( BL12, BLN12, WL52);
sram_cell_6t_3 inst_cell_52_11 ( BL11, BLN11, WL52);
sram_cell_6t_3 inst_cell_52_10 ( BL10, BLN10, WL52);
sram_cell_6t_3 inst_cell_52_9 ( BL9, BLN9, WL52);
sram_cell_6t_3 inst_cell_52_8 ( BL8, BLN8, WL52);
sram_cell_6t_3 inst_cell_52_7 ( BL7, BLN7, WL52);
sram_cell_6t_3 inst_cell_52_6 ( BL6, BLN6, WL52);
sram_cell_6t_3 inst_cell_52_5 ( BL5, BLN5, WL52);
sram_cell_6t_3 inst_cell_52_4 ( BL4, BLN4, WL52);
sram_cell_6t_3 inst_cell_52_3 ( BL3, BLN3, WL52);
sram_cell_6t_3 inst_cell_52_2 ( BL2, BLN2, WL52);
sram_cell_6t_3 inst_cell_52_1 ( BL1, BLN1, WL52);
sram_cell_6t_3 inst_cell_52_0 ( BL0, BLN0, WL52);
sram_cell_6t_3 inst_cell_51_63 ( BL63, BLN63, WL51);
sram_cell_6t_3 inst_cell_51_62 ( BL62, BLN62, WL51);
sram_cell_6t_3 inst_cell_51_61 ( BL61, BLN61, WL51);
sram_cell_6t_3 inst_cell_51_60 ( BL60, BLN60, WL51);
sram_cell_6t_3 inst_cell_51_59 ( BL59, BLN59, WL51);
sram_cell_6t_3 inst_cell_51_58 ( BL58, BLN58, WL51);
sram_cell_6t_3 inst_cell_51_57 ( BL57, BLN57, WL51);
sram_cell_6t_3 inst_cell_51_56 ( BL56, BLN56, WL51);
sram_cell_6t_3 inst_cell_51_55 ( BL55, BLN55, WL51);
sram_cell_6t_3 inst_cell_51_54 ( BL54, BLN54, WL51);
sram_cell_6t_3 inst_cell_51_53 ( BL53, BLN53, WL51);
sram_cell_6t_3 inst_cell_51_52 ( BL52, BLN52, WL51);
sram_cell_6t_3 inst_cell_51_51 ( BL51, BLN51, WL51);
sram_cell_6t_3 inst_cell_51_50 ( BL50, BLN50, WL51);
sram_cell_6t_3 inst_cell_51_49 ( BL49, BLN49, WL51);
sram_cell_6t_3 inst_cell_51_48 ( BL48, BLN48, WL51);
sram_cell_6t_3 inst_cell_51_47 ( BL47, BLN47, WL51);
sram_cell_6t_3 inst_cell_51_46 ( BL46, BLN46, WL51);
sram_cell_6t_3 inst_cell_51_45 ( BL45, BLN45, WL51);
sram_cell_6t_3 inst_cell_51_44 ( BL44, BLN44, WL51);
sram_cell_6t_3 inst_cell_51_43 ( BL43, BLN43, WL51);
sram_cell_6t_3 inst_cell_51_42 ( BL42, BLN42, WL51);
sram_cell_6t_3 inst_cell_51_41 ( BL41, BLN41, WL51);
sram_cell_6t_3 inst_cell_51_40 ( BL40, BLN40, WL51);
sram_cell_6t_3 inst_cell_51_39 ( BL39, BLN39, WL51);
sram_cell_6t_3 inst_cell_51_38 ( BL38, BLN38, WL51);
sram_cell_6t_3 inst_cell_51_37 ( BL37, BLN37, WL51);
sram_cell_6t_3 inst_cell_51_36 ( BL36, BLN36, WL51);
sram_cell_6t_3 inst_cell_51_35 ( BL35, BLN35, WL51);
sram_cell_6t_3 inst_cell_51_34 ( BL34, BLN34, WL51);
sram_cell_6t_3 inst_cell_51_33 ( BL33, BLN33, WL51);
sram_cell_6t_3 inst_cell_51_32 ( BL32, BLN32, WL51);
sram_cell_6t_3 inst_cell_51_31 ( BL31, BLN31, WL51);
sram_cell_6t_3 inst_cell_51_30 ( BL30, BLN30, WL51);
sram_cell_6t_3 inst_cell_51_29 ( BL29, BLN29, WL51);
sram_cell_6t_3 inst_cell_51_28 ( BL28, BLN28, WL51);
sram_cell_6t_3 inst_cell_51_27 ( BL27, BLN27, WL51);
sram_cell_6t_3 inst_cell_51_26 ( BL26, BLN26, WL51);
sram_cell_6t_3 inst_cell_51_25 ( BL25, BLN25, WL51);
sram_cell_6t_3 inst_cell_51_24 ( BL24, BLN24, WL51);
sram_cell_6t_3 inst_cell_51_23 ( BL23, BLN23, WL51);
sram_cell_6t_3 inst_cell_51_22 ( BL22, BLN22, WL51);
sram_cell_6t_3 inst_cell_51_21 ( BL21, BLN21, WL51);
sram_cell_6t_3 inst_cell_51_20 ( BL20, BLN20, WL51);
sram_cell_6t_3 inst_cell_51_19 ( BL19, BLN19, WL51);
sram_cell_6t_3 inst_cell_51_18 ( BL18, BLN18, WL51);
sram_cell_6t_3 inst_cell_51_17 ( BL17, BLN17, WL51);
sram_cell_6t_3 inst_cell_51_16 ( BL16, BLN16, WL51);
sram_cell_6t_3 inst_cell_51_15 ( BL15, BLN15, WL51);
sram_cell_6t_3 inst_cell_51_14 ( BL14, BLN14, WL51);
sram_cell_6t_3 inst_cell_51_13 ( BL13, BLN13, WL51);
sram_cell_6t_3 inst_cell_51_12 ( BL12, BLN12, WL51);
sram_cell_6t_3 inst_cell_51_11 ( BL11, BLN11, WL51);
sram_cell_6t_3 inst_cell_51_10 ( BL10, BLN10, WL51);
sram_cell_6t_3 inst_cell_51_9 ( BL9, BLN9, WL51);
sram_cell_6t_3 inst_cell_51_8 ( BL8, BLN8, WL51);
sram_cell_6t_3 inst_cell_51_7 ( BL7, BLN7, WL51);
sram_cell_6t_3 inst_cell_51_6 ( BL6, BLN6, WL51);
sram_cell_6t_3 inst_cell_51_5 ( BL5, BLN5, WL51);
sram_cell_6t_3 inst_cell_51_4 ( BL4, BLN4, WL51);
sram_cell_6t_3 inst_cell_51_3 ( BL3, BLN3, WL51);
sram_cell_6t_3 inst_cell_51_2 ( BL2, BLN2, WL51);
sram_cell_6t_3 inst_cell_51_1 ( BL1, BLN1, WL51);
sram_cell_6t_3 inst_cell_51_0 ( BL0, BLN0, WL51);
sram_cell_6t_3 inst_cell_50_63 ( BL63, BLN63, WL50);
sram_cell_6t_3 inst_cell_50_62 ( BL62, BLN62, WL50);
sram_cell_6t_3 inst_cell_50_61 ( BL61, BLN61, WL50);
sram_cell_6t_3 inst_cell_50_60 ( BL60, BLN60, WL50);
sram_cell_6t_3 inst_cell_50_59 ( BL59, BLN59, WL50);
sram_cell_6t_3 inst_cell_50_58 ( BL58, BLN58, WL50);
sram_cell_6t_3 inst_cell_50_57 ( BL57, BLN57, WL50);
sram_cell_6t_3 inst_cell_50_56 ( BL56, BLN56, WL50);
sram_cell_6t_3 inst_cell_50_55 ( BL55, BLN55, WL50);
sram_cell_6t_3 inst_cell_50_54 ( BL54, BLN54, WL50);
sram_cell_6t_3 inst_cell_50_53 ( BL53, BLN53, WL50);
sram_cell_6t_3 inst_cell_50_52 ( BL52, BLN52, WL50);
sram_cell_6t_3 inst_cell_50_51 ( BL51, BLN51, WL50);
sram_cell_6t_3 inst_cell_50_50 ( BL50, BLN50, WL50);
sram_cell_6t_3 inst_cell_50_49 ( BL49, BLN49, WL50);
sram_cell_6t_3 inst_cell_50_48 ( BL48, BLN48, WL50);
sram_cell_6t_3 inst_cell_50_47 ( BL47, BLN47, WL50);
sram_cell_6t_3 inst_cell_50_46 ( BL46, BLN46, WL50);
sram_cell_6t_3 inst_cell_50_45 ( BL45, BLN45, WL50);
sram_cell_6t_3 inst_cell_50_44 ( BL44, BLN44, WL50);
sram_cell_6t_3 inst_cell_50_43 ( BL43, BLN43, WL50);
sram_cell_6t_3 inst_cell_50_42 ( BL42, BLN42, WL50);
sram_cell_6t_3 inst_cell_50_41 ( BL41, BLN41, WL50);
sram_cell_6t_3 inst_cell_50_40 ( BL40, BLN40, WL50);
sram_cell_6t_3 inst_cell_50_39 ( BL39, BLN39, WL50);
sram_cell_6t_3 inst_cell_50_38 ( BL38, BLN38, WL50);
sram_cell_6t_3 inst_cell_50_37 ( BL37, BLN37, WL50);
sram_cell_6t_3 inst_cell_50_36 ( BL36, BLN36, WL50);
sram_cell_6t_3 inst_cell_50_35 ( BL35, BLN35, WL50);
sram_cell_6t_3 inst_cell_50_34 ( BL34, BLN34, WL50);
sram_cell_6t_3 inst_cell_50_33 ( BL33, BLN33, WL50);
sram_cell_6t_3 inst_cell_50_32 ( BL32, BLN32, WL50);
sram_cell_6t_3 inst_cell_50_31 ( BL31, BLN31, WL50);
sram_cell_6t_3 inst_cell_50_30 ( BL30, BLN30, WL50);
sram_cell_6t_3 inst_cell_50_29 ( BL29, BLN29, WL50);
sram_cell_6t_3 inst_cell_50_28 ( BL28, BLN28, WL50);
sram_cell_6t_3 inst_cell_50_27 ( BL27, BLN27, WL50);
sram_cell_6t_3 inst_cell_50_26 ( BL26, BLN26, WL50);
sram_cell_6t_3 inst_cell_50_25 ( BL25, BLN25, WL50);
sram_cell_6t_3 inst_cell_50_24 ( BL24, BLN24, WL50);
sram_cell_6t_3 inst_cell_50_23 ( BL23, BLN23, WL50);
sram_cell_6t_3 inst_cell_50_22 ( BL22, BLN22, WL50);
sram_cell_6t_3 inst_cell_50_21 ( BL21, BLN21, WL50);
sram_cell_6t_3 inst_cell_50_20 ( BL20, BLN20, WL50);
sram_cell_6t_3 inst_cell_50_19 ( BL19, BLN19, WL50);
sram_cell_6t_3 inst_cell_50_18 ( BL18, BLN18, WL50);
sram_cell_6t_3 inst_cell_50_17 ( BL17, BLN17, WL50);
sram_cell_6t_3 inst_cell_50_16 ( BL16, BLN16, WL50);
sram_cell_6t_3 inst_cell_50_15 ( BL15, BLN15, WL50);
sram_cell_6t_3 inst_cell_50_14 ( BL14, BLN14, WL50);
sram_cell_6t_3 inst_cell_50_13 ( BL13, BLN13, WL50);
sram_cell_6t_3 inst_cell_50_12 ( BL12, BLN12, WL50);
sram_cell_6t_3 inst_cell_50_11 ( BL11, BLN11, WL50);
sram_cell_6t_3 inst_cell_50_10 ( BL10, BLN10, WL50);
sram_cell_6t_3 inst_cell_50_9 ( BL9, BLN9, WL50);
sram_cell_6t_3 inst_cell_50_8 ( BL8, BLN8, WL50);
sram_cell_6t_3 inst_cell_50_7 ( BL7, BLN7, WL50);
sram_cell_6t_3 inst_cell_50_6 ( BL6, BLN6, WL50);
sram_cell_6t_3 inst_cell_50_5 ( BL5, BLN5, WL50);
sram_cell_6t_3 inst_cell_50_4 ( BL4, BLN4, WL50);
sram_cell_6t_3 inst_cell_50_3 ( BL3, BLN3, WL50);
sram_cell_6t_3 inst_cell_50_2 ( BL2, BLN2, WL50);
sram_cell_6t_3 inst_cell_50_1 ( BL1, BLN1, WL50);
sram_cell_6t_3 inst_cell_50_0 ( BL0, BLN0, WL50);
sram_cell_6t_3 inst_cell_49_63 ( BL63, BLN63, WL49);
sram_cell_6t_3 inst_cell_49_62 ( BL62, BLN62, WL49);
sram_cell_6t_3 inst_cell_49_61 ( BL61, BLN61, WL49);
sram_cell_6t_3 inst_cell_49_60 ( BL60, BLN60, WL49);
sram_cell_6t_3 inst_cell_49_59 ( BL59, BLN59, WL49);
sram_cell_6t_3 inst_cell_49_58 ( BL58, BLN58, WL49);
sram_cell_6t_3 inst_cell_49_57 ( BL57, BLN57, WL49);
sram_cell_6t_3 inst_cell_49_56 ( BL56, BLN56, WL49);
sram_cell_6t_3 inst_cell_49_55 ( BL55, BLN55, WL49);
sram_cell_6t_3 inst_cell_49_54 ( BL54, BLN54, WL49);
sram_cell_6t_3 inst_cell_49_53 ( BL53, BLN53, WL49);
sram_cell_6t_3 inst_cell_49_52 ( BL52, BLN52, WL49);
sram_cell_6t_3 inst_cell_49_51 ( BL51, BLN51, WL49);
sram_cell_6t_3 inst_cell_49_50 ( BL50, BLN50, WL49);
sram_cell_6t_3 inst_cell_49_23 ( BL23, BLN23, WL49);
sram_cell_6t_3 inst_cell_48_23 ( BL23, BLN23, WL48);
sram_cell_6t_3 inst_cell_49_22 ( BL22, BLN22, WL49);
sram_cell_6t_3 inst_cell_48_22 ( BL22, BLN22, WL48);
sram_cell_6t_3 inst_cell_49_21 ( BL21, BLN21, WL49);
sram_cell_6t_3 inst_cell_48_21 ( BL21, BLN21, WL48);
sram_cell_6t_3 inst_cell_49_20 ( BL20, BLN20, WL49);
sram_cell_6t_3 inst_cell_48_20 ( BL20, BLN20, WL48);
sram_cell_6t_3 inst_cell_49_19 ( BL19, BLN19, WL49);
sram_cell_6t_3 inst_cell_48_19 ( BL19, BLN19, WL48);
sram_cell_6t_3 inst_cell_49_18 ( BL18, BLN18, WL49);
sram_cell_6t_3 inst_cell_48_18 ( BL18, BLN18, WL48);
sram_cell_6t_3 inst_cell_49_17 ( BL17, BLN17, WL49);
sram_cell_6t_3 inst_cell_48_17 ( BL17, BLN17, WL48);
sram_cell_6t_3 inst_cell_49_16 ( BL16, BLN16, WL49);
sram_cell_6t_3 inst_cell_48_16 ( BL16, BLN16, WL48);
sram_cell_6t_3 inst_cell_49_15 ( BL15, BLN15, WL49);
sram_cell_6t_3 inst_cell_48_15 ( BL15, BLN15, WL48);
sram_cell_6t_3 inst_cell_49_14 ( BL14, BLN14, WL49);
sram_cell_6t_3 inst_cell_48_14 ( BL14, BLN14, WL48);
sram_cell_6t_3 inst_cell_49_13 ( BL13, BLN13, WL49);
sram_cell_6t_3 inst_cell_48_13 ( BL13, BLN13, WL48);
sram_cell_6t_3 inst_cell_49_12 ( BL12, BLN12, WL49);
sram_cell_6t_3 inst_cell_48_12 ( BL12, BLN12, WL48);
sram_cell_6t_3 inst_cell_49_11 ( BL11, BLN11, WL49);
sram_cell_6t_3 inst_cell_48_11 ( BL11, BLN11, WL48);
sram_cell_6t_3 inst_cell_49_10 ( BL10, BLN10, WL49);
sram_cell_6t_3 inst_cell_48_10 ( BL10, BLN10, WL48);
sram_cell_6t_3 inst_cell_49_9 ( BL9, BLN9, WL49);
sram_cell_6t_3 inst_cell_48_9 ( BL9, BLN9, WL48);
sram_cell_6t_3 inst_cell_49_8 ( BL8, BLN8, WL49);
sram_cell_6t_3 inst_cell_48_8 ( BL8, BLN8, WL48);
sram_cell_6t_3 inst_cell_49_7 ( BL7, BLN7, WL49);
sram_cell_6t_3 inst_cell_48_7 ( BL7, BLN7, WL48);
sram_cell_6t_3 inst_cell_49_6 ( BL6, BLN6, WL49);
sram_cell_6t_3 inst_cell_48_6 ( BL6, BLN6, WL48);
sram_cell_6t_3 inst_cell_49_5 ( BL5, BLN5, WL49);
sram_cell_6t_3 inst_cell_48_5 ( BL5, BLN5, WL48);
sram_cell_6t_3 inst_cell_49_4 ( BL4, BLN4, WL49);
sram_cell_6t_3 inst_cell_48_4 ( BL4, BLN4, WL48);
sram_cell_6t_3 inst_cell_49_3 ( BL3, BLN3, WL49);
sram_cell_6t_3 inst_cell_48_3 ( BL3, BLN3, WL48);
sram_cell_6t_3 inst_cell_49_2 ( BL2, BLN2, WL49);
sram_cell_6t_3 inst_cell_48_2 ( BL2, BLN2, WL48);
sram_cell_6t_3 inst_cell_49_1 ( BL1, BLN1, WL49);
sram_cell_6t_3 inst_cell_48_1 ( BL1, BLN1, WL48);
sram_cell_6t_3 inst_cell_49_0 ( BL0, BLN0, WL49);
sram_cell_6t_3 inst_cell_48_0 ( BL0, BLN0, WL48);
sram_cell_6t_3 inst_cell_48_63 ( BL63, BLN63, WL48);
sram_cell_6t_3 inst_cell_47_63 ( BL63, BLN63, WL47);
sram_cell_6t_3 inst_cell_48_62 ( BL62, BLN62, WL48);
sram_cell_6t_3 inst_cell_47_62 ( BL62, BLN62, WL47);
sram_cell_6t_3 inst_cell_48_61 ( BL61, BLN61, WL48);
sram_cell_6t_3 inst_cell_47_61 ( BL61, BLN61, WL47);
sram_cell_6t_3 inst_cell_48_60 ( BL60, BLN60, WL48);
sram_cell_6t_3 inst_cell_47_60 ( BL60, BLN60, WL47);
sram_cell_6t_3 inst_cell_48_59 ( BL59, BLN59, WL48);
sram_cell_6t_3 inst_cell_47_59 ( BL59, BLN59, WL47);
sram_cell_6t_3 inst_cell_48_58 ( BL58, BLN58, WL48);
sram_cell_6t_3 inst_cell_47_58 ( BL58, BLN58, WL47);
sram_cell_6t_3 inst_cell_48_57 ( BL57, BLN57, WL48);
sram_cell_6t_3 inst_cell_47_57 ( BL57, BLN57, WL47);
sram_cell_6t_3 inst_cell_48_56 ( BL56, BLN56, WL48);
sram_cell_6t_3 inst_cell_47_56 ( BL56, BLN56, WL47);
sram_cell_6t_3 inst_cell_48_55 ( BL55, BLN55, WL48);
sram_cell_6t_3 inst_cell_47_55 ( BL55, BLN55, WL47);
sram_cell_6t_3 inst_cell_48_54 ( BL54, BLN54, WL48);
sram_cell_6t_3 inst_cell_47_54 ( BL54, BLN54, WL47);
sram_cell_6t_3 inst_cell_48_53 ( BL53, BLN53, WL48);
sram_cell_6t_3 inst_cell_47_53 ( BL53, BLN53, WL47);
sram_cell_6t_3 inst_cell_48_52 ( BL52, BLN52, WL48);
sram_cell_6t_3 inst_cell_47_52 ( BL52, BLN52, WL47);
sram_cell_6t_3 inst_cell_48_51 ( BL51, BLN51, WL48);
sram_cell_6t_3 inst_cell_47_51 ( BL51, BLN51, WL47);
sram_cell_6t_3 inst_cell_48_50 ( BL50, BLN50, WL48);
sram_cell_6t_3 inst_cell_47_50 ( BL50, BLN50, WL47);
sram_cell_6t_3 inst_cell_49_49 ( BL49, BLN49, WL49);
sram_cell_6t_3 inst_cell_49_48 ( BL48, BLN48, WL49);
sram_cell_6t_3 inst_cell_49_47 ( BL47, BLN47, WL49);
sram_cell_6t_3 inst_cell_49_46 ( BL46, BLN46, WL49);
sram_cell_6t_3 inst_cell_49_45 ( BL45, BLN45, WL49);
sram_cell_6t_3 inst_cell_49_44 ( BL44, BLN44, WL49);
sram_cell_6t_3 inst_cell_49_43 ( BL43, BLN43, WL49);
sram_cell_6t_3 inst_cell_49_42 ( BL42, BLN42, WL49);
sram_cell_6t_3 inst_cell_49_41 ( BL41, BLN41, WL49);
sram_cell_6t_3 inst_cell_49_40 ( BL40, BLN40, WL49);
sram_cell_6t_3 inst_cell_49_39 ( BL39, BLN39, WL49);
sram_cell_6t_3 inst_cell_49_38 ( BL38, BLN38, WL49);
sram_cell_6t_3 inst_cell_49_37 ( BL37, BLN37, WL49);
sram_cell_6t_3 inst_cell_49_36 ( BL36, BLN36, WL49);
sram_cell_6t_3 inst_cell_49_35 ( BL35, BLN35, WL49);
sram_cell_6t_3 inst_cell_49_34 ( BL34, BLN34, WL49);
sram_cell_6t_3 inst_cell_49_33 ( BL33, BLN33, WL49);
sram_cell_6t_3 inst_cell_49_32 ( BL32, BLN32, WL49);
sram_cell_6t_3 inst_cell_49_31 ( BL31, BLN31, WL49);
sram_cell_6t_3 inst_cell_49_30 ( BL30, BLN30, WL49);
sram_cell_6t_3 inst_cell_49_29 ( BL29, BLN29, WL49);
sram_cell_6t_3 inst_cell_49_28 ( BL28, BLN28, WL49);
sram_cell_6t_3 inst_cell_49_27 ( BL27, BLN27, WL49);
sram_cell_6t_3 inst_cell_49_26 ( BL26, BLN26, WL49);
sram_cell_6t_3 inst_cell_49_25 ( BL25, BLN25, WL49);
sram_cell_6t_3 inst_cell_49_24 ( BL24, BLN24, WL49);
sram_cell_6t_3 inst_cell_48_49 ( BL49, BLN49, WL48);
sram_cell_6t_3 inst_cell_48_48 ( BL48, BLN48, WL48);
sram_cell_6t_3 inst_cell_48_47 ( BL47, BLN47, WL48);
sram_cell_6t_3 inst_cell_48_46 ( BL46, BLN46, WL48);
sram_cell_6t_3 inst_cell_48_45 ( BL45, BLN45, WL48);
sram_cell_6t_3 inst_cell_48_44 ( BL44, BLN44, WL48);
sram_cell_6t_3 inst_cell_48_43 ( BL43, BLN43, WL48);
sram_cell_6t_3 inst_cell_48_42 ( BL42, BLN42, WL48);
sram_cell_6t_3 inst_cell_48_41 ( BL41, BLN41, WL48);
sram_cell_6t_3 inst_cell_48_40 ( BL40, BLN40, WL48);
sram_cell_6t_3 inst_cell_48_39 ( BL39, BLN39, WL48);
sram_cell_6t_3 inst_cell_48_38 ( BL38, BLN38, WL48);
sram_cell_6t_3 inst_cell_48_37 ( BL37, BLN37, WL48);
sram_cell_6t_3 inst_cell_48_36 ( BL36, BLN36, WL48);
sram_cell_6t_3 inst_cell_48_35 ( BL35, BLN35, WL48);
sram_cell_6t_3 inst_cell_48_34 ( BL34, BLN34, WL48);
sram_cell_6t_3 inst_cell_48_33 ( BL33, BLN33, WL48);
sram_cell_6t_3 inst_cell_48_32 ( BL32, BLN32, WL48);
sram_cell_6t_3 inst_cell_48_31 ( BL31, BLN31, WL48);
sram_cell_6t_3 inst_cell_48_30 ( BL30, BLN30, WL48);
sram_cell_6t_3 inst_cell_48_29 ( BL29, BLN29, WL48);
sram_cell_6t_3 inst_cell_48_28 ( BL28, BLN28, WL48);
sram_cell_6t_3 inst_cell_48_27 ( BL27, BLN27, WL48);
sram_cell_6t_3 inst_cell_48_26 ( BL26, BLN26, WL48);
sram_cell_6t_3 inst_cell_48_25 ( BL25, BLN25, WL48);
sram_cell_6t_3 inst_cell_48_24 ( BL24, BLN24, WL48);
sram_cell_6t_3 inst_cell_47_49 ( BL49, BLN49, WL47);
sram_cell_6t_3 inst_cell_47_48 ( BL48, BLN48, WL47);
sram_cell_6t_3 inst_cell_47_47 ( BL47, BLN47, WL47);
sram_cell_6t_3 inst_cell_47_46 ( BL46, BLN46, WL47);
sram_cell_6t_3 inst_cell_47_45 ( BL45, BLN45, WL47);
sram_cell_6t_3 inst_cell_47_44 ( BL44, BLN44, WL47);
sram_cell_6t_3 inst_cell_47_43 ( BL43, BLN43, WL47);
sram_cell_6t_3 inst_cell_47_42 ( BL42, BLN42, WL47);
sram_cell_6t_3 inst_cell_47_41 ( BL41, BLN41, WL47);
sram_cell_6t_3 inst_cell_47_40 ( BL40, BLN40, WL47);
sram_cell_6t_3 inst_cell_47_39 ( BL39, BLN39, WL47);
sram_cell_6t_3 inst_cell_47_38 ( BL38, BLN38, WL47);
sram_cell_6t_3 inst_cell_47_37 ( BL37, BLN37, WL47);
sram_cell_6t_3 inst_cell_47_36 ( BL36, BLN36, WL47);
sram_cell_6t_3 inst_cell_47_35 ( BL35, BLN35, WL47);
sram_cell_6t_3 inst_cell_47_34 ( BL34, BLN34, WL47);
sram_cell_6t_3 inst_cell_47_33 ( BL33, BLN33, WL47);
sram_cell_6t_3 inst_cell_47_32 ( BL32, BLN32, WL47);
sram_cell_6t_3 inst_cell_47_31 ( BL31, BLN31, WL47);
sram_cell_6t_3 inst_cell_47_30 ( BL30, BLN30, WL47);
sram_cell_6t_3 inst_cell_47_29 ( BL29, BLN29, WL47);
sram_cell_6t_3 inst_cell_47_28 ( BL28, BLN28, WL47);
sram_cell_6t_3 inst_cell_47_27 ( BL27, BLN27, WL47);
sram_cell_6t_3 inst_cell_47_26 ( BL26, BLN26, WL47);
sram_cell_6t_3 inst_cell_47_25 ( BL25, BLN25, WL47);
sram_cell_6t_3 inst_cell_47_24 ( BL24, BLN24, WL47);
sram_cell_6t_3 inst_cell_46_63 ( BL63, BLN63, WL46);
sram_cell_6t_3 inst_cell_45_63 ( BL63, BLN63, WL45);
sram_cell_6t_3 inst_cell_46_62 ( BL62, BLN62, WL46);
sram_cell_6t_3 inst_cell_45_62 ( BL62, BLN62, WL45);
sram_cell_6t_3 inst_cell_46_61 ( BL61, BLN61, WL46);
sram_cell_6t_3 inst_cell_45_61 ( BL61, BLN61, WL45);
sram_cell_6t_3 inst_cell_46_60 ( BL60, BLN60, WL46);
sram_cell_6t_3 inst_cell_45_60 ( BL60, BLN60, WL45);
sram_cell_6t_3 inst_cell_46_59 ( BL59, BLN59, WL46);
sram_cell_6t_3 inst_cell_45_59 ( BL59, BLN59, WL45);
sram_cell_6t_3 inst_cell_46_58 ( BL58, BLN58, WL46);
sram_cell_6t_3 inst_cell_45_58 ( BL58, BLN58, WL45);
sram_cell_6t_3 inst_cell_46_57 ( BL57, BLN57, WL46);
sram_cell_6t_3 inst_cell_45_57 ( BL57, BLN57, WL45);
sram_cell_6t_3 inst_cell_46_56 ( BL56, BLN56, WL46);
sram_cell_6t_3 inst_cell_45_56 ( BL56, BLN56, WL45);
sram_cell_6t_3 inst_cell_46_55 ( BL55, BLN55, WL46);
sram_cell_6t_3 inst_cell_45_55 ( BL55, BLN55, WL45);
sram_cell_6t_3 inst_cell_46_54 ( BL54, BLN54, WL46);
sram_cell_6t_3 inst_cell_45_54 ( BL54, BLN54, WL45);
sram_cell_6t_3 inst_cell_46_53 ( BL53, BLN53, WL46);
sram_cell_6t_3 inst_cell_45_53 ( BL53, BLN53, WL45);
sram_cell_6t_3 inst_cell_46_52 ( BL52, BLN52, WL46);
sram_cell_6t_3 inst_cell_45_52 ( BL52, BLN52, WL45);
sram_cell_6t_3 inst_cell_46_51 ( BL51, BLN51, WL46);
sram_cell_6t_3 inst_cell_45_51 ( BL51, BLN51, WL45);
sram_cell_6t_3 inst_cell_46_50 ( BL50, BLN50, WL46);
sram_cell_6t_3 inst_cell_45_50 ( BL50, BLN50, WL45);
sram_cell_6t_3 inst_cell_46_49 ( BL49, BLN49, WL46);
sram_cell_6t_3 inst_cell_45_49 ( BL49, BLN49, WL45);
sram_cell_6t_3 inst_cell_46_48 ( BL48, BLN48, WL46);
sram_cell_6t_3 inst_cell_45_48 ( BL48, BLN48, WL45);
sram_cell_6t_3 inst_cell_46_47 ( BL47, BLN47, WL46);
sram_cell_6t_3 inst_cell_45_47 ( BL47, BLN47, WL45);
sram_cell_6t_3 inst_cell_46_46 ( BL46, BLN46, WL46);
sram_cell_6t_3 inst_cell_45_46 ( BL46, BLN46, WL45);
sram_cell_6t_3 inst_cell_46_45 ( BL45, BLN45, WL46);
sram_cell_6t_3 inst_cell_45_45 ( BL45, BLN45, WL45);
sram_cell_6t_3 inst_cell_46_44 ( BL44, BLN44, WL46);
sram_cell_6t_3 inst_cell_45_44 ( BL44, BLN44, WL45);
sram_cell_6t_3 inst_cell_46_43 ( BL43, BLN43, WL46);
sram_cell_6t_3 inst_cell_45_43 ( BL43, BLN43, WL45);
sram_cell_6t_3 inst_cell_46_42 ( BL42, BLN42, WL46);
sram_cell_6t_3 inst_cell_45_42 ( BL42, BLN42, WL45);
sram_cell_6t_3 inst_cell_46_41 ( BL41, BLN41, WL46);
sram_cell_6t_3 inst_cell_45_41 ( BL41, BLN41, WL45);
sram_cell_6t_3 inst_cell_46_40 ( BL40, BLN40, WL46);
sram_cell_6t_3 inst_cell_45_40 ( BL40, BLN40, WL45);
sram_cell_6t_3 inst_cell_46_39 ( BL39, BLN39, WL46);
sram_cell_6t_3 inst_cell_45_39 ( BL39, BLN39, WL45);
sram_cell_6t_3 inst_cell_46_38 ( BL38, BLN38, WL46);
sram_cell_6t_3 inst_cell_45_38 ( BL38, BLN38, WL45);
sram_cell_6t_3 inst_cell_46_37 ( BL37, BLN37, WL46);
sram_cell_6t_3 inst_cell_45_37 ( BL37, BLN37, WL45);
sram_cell_6t_3 inst_cell_46_36 ( BL36, BLN36, WL46);
sram_cell_6t_3 inst_cell_45_36 ( BL36, BLN36, WL45);
sram_cell_6t_3 inst_cell_46_35 ( BL35, BLN35, WL46);
sram_cell_6t_3 inst_cell_45_35 ( BL35, BLN35, WL45);
sram_cell_6t_3 inst_cell_46_34 ( BL34, BLN34, WL46);
sram_cell_6t_3 inst_cell_45_34 ( BL34, BLN34, WL45);
sram_cell_6t_3 inst_cell_46_33 ( BL33, BLN33, WL46);
sram_cell_6t_3 inst_cell_45_33 ( BL33, BLN33, WL45);
sram_cell_6t_3 inst_cell_46_32 ( BL32, BLN32, WL46);
sram_cell_6t_3 inst_cell_45_32 ( BL32, BLN32, WL45);
sram_cell_6t_3 inst_cell_46_31 ( BL31, BLN31, WL46);
sram_cell_6t_3 inst_cell_45_31 ( BL31, BLN31, WL45);
sram_cell_6t_3 inst_cell_46_30 ( BL30, BLN30, WL46);
sram_cell_6t_3 inst_cell_45_30 ( BL30, BLN30, WL45);
sram_cell_6t_3 inst_cell_46_29 ( BL29, BLN29, WL46);
sram_cell_6t_3 inst_cell_45_29 ( BL29, BLN29, WL45);
sram_cell_6t_3 inst_cell_46_28 ( BL28, BLN28, WL46);
sram_cell_6t_3 inst_cell_45_28 ( BL28, BLN28, WL45);
sram_cell_6t_3 inst_cell_46_27 ( BL27, BLN27, WL46);
sram_cell_6t_3 inst_cell_45_27 ( BL27, BLN27, WL45);
sram_cell_6t_3 inst_cell_46_26 ( BL26, BLN26, WL46);
sram_cell_6t_3 inst_cell_45_26 ( BL26, BLN26, WL45);
sram_cell_6t_3 inst_cell_46_25 ( BL25, BLN25, WL46);
sram_cell_6t_3 inst_cell_45_25 ( BL25, BLN25, WL45);
sram_cell_6t_3 inst_cell_46_24 ( BL24, BLN24, WL46);
sram_cell_6t_3 inst_cell_45_24 ( BL24, BLN24, WL45);
sram_cell_6t_3 inst_cell_47_23 ( BL23, BLN23, WL47);
sram_cell_6t_3 inst_cell_47_22 ( BL22, BLN22, WL47);
sram_cell_6t_3 inst_cell_47_21 ( BL21, BLN21, WL47);
sram_cell_6t_3 inst_cell_47_20 ( BL20, BLN20, WL47);
sram_cell_6t_3 inst_cell_47_19 ( BL19, BLN19, WL47);
sram_cell_6t_3 inst_cell_47_18 ( BL18, BLN18, WL47);
sram_cell_6t_3 inst_cell_47_17 ( BL17, BLN17, WL47);
sram_cell_6t_3 inst_cell_47_16 ( BL16, BLN16, WL47);
sram_cell_6t_3 inst_cell_47_15 ( BL15, BLN15, WL47);
sram_cell_6t_3 inst_cell_47_14 ( BL14, BLN14, WL47);
sram_cell_6t_3 inst_cell_47_13 ( BL13, BLN13, WL47);
sram_cell_6t_3 inst_cell_47_12 ( BL12, BLN12, WL47);
sram_cell_6t_3 inst_cell_47_11 ( BL11, BLN11, WL47);
sram_cell_6t_3 inst_cell_47_10 ( BL10, BLN10, WL47);
sram_cell_6t_3 inst_cell_47_9 ( BL9, BLN9, WL47);
sram_cell_6t_3 inst_cell_47_8 ( BL8, BLN8, WL47);
sram_cell_6t_3 inst_cell_47_7 ( BL7, BLN7, WL47);
sram_cell_6t_3 inst_cell_47_6 ( BL6, BLN6, WL47);
sram_cell_6t_3 inst_cell_47_5 ( BL5, BLN5, WL47);
sram_cell_6t_3 inst_cell_47_4 ( BL4, BLN4, WL47);
sram_cell_6t_3 inst_cell_47_3 ( BL3, BLN3, WL47);
sram_cell_6t_3 inst_cell_47_2 ( BL2, BLN2, WL47);
sram_cell_6t_3 inst_cell_47_1 ( BL1, BLN1, WL47);
sram_cell_6t_3 inst_cell_47_0 ( BL0, BLN0, WL47);
sram_cell_6t_3 inst_cell_46_23 ( BL23, BLN23, WL46);
sram_cell_6t_3 inst_cell_46_22 ( BL22, BLN22, WL46);
sram_cell_6t_3 inst_cell_46_21 ( BL21, BLN21, WL46);
sram_cell_6t_3 inst_cell_46_20 ( BL20, BLN20, WL46);
sram_cell_6t_3 inst_cell_46_19 ( BL19, BLN19, WL46);
sram_cell_6t_3 inst_cell_46_18 ( BL18, BLN18, WL46);
sram_cell_6t_3 inst_cell_46_17 ( BL17, BLN17, WL46);
sram_cell_6t_3 inst_cell_46_16 ( BL16, BLN16, WL46);
sram_cell_6t_3 inst_cell_46_15 ( BL15, BLN15, WL46);
sram_cell_6t_3 inst_cell_46_14 ( BL14, BLN14, WL46);
sram_cell_6t_3 inst_cell_46_13 ( BL13, BLN13, WL46);
sram_cell_6t_3 inst_cell_46_12 ( BL12, BLN12, WL46);
sram_cell_6t_3 inst_cell_46_11 ( BL11, BLN11, WL46);
sram_cell_6t_3 inst_cell_46_10 ( BL10, BLN10, WL46);
sram_cell_6t_3 inst_cell_46_9 ( BL9, BLN9, WL46);
sram_cell_6t_3 inst_cell_46_8 ( BL8, BLN8, WL46);
sram_cell_6t_3 inst_cell_46_7 ( BL7, BLN7, WL46);
sram_cell_6t_3 inst_cell_46_6 ( BL6, BLN6, WL46);
sram_cell_6t_3 inst_cell_46_5 ( BL5, BLN5, WL46);
sram_cell_6t_3 inst_cell_46_4 ( BL4, BLN4, WL46);
sram_cell_6t_3 inst_cell_46_3 ( BL3, BLN3, WL46);
sram_cell_6t_3 inst_cell_46_2 ( BL2, BLN2, WL46);
sram_cell_6t_3 inst_cell_46_1 ( BL1, BLN1, WL46);
sram_cell_6t_3 inst_cell_46_0 ( BL0, BLN0, WL46);
sram_cell_6t_3 inst_cell_45_23 ( BL23, BLN23, WL45);
sram_cell_6t_3 inst_cell_45_22 ( BL22, BLN22, WL45);
sram_cell_6t_3 inst_cell_45_21 ( BL21, BLN21, WL45);
sram_cell_6t_3 inst_cell_45_20 ( BL20, BLN20, WL45);
sram_cell_6t_3 inst_cell_45_19 ( BL19, BLN19, WL45);
sram_cell_6t_3 inst_cell_45_18 ( BL18, BLN18, WL45);
sram_cell_6t_3 inst_cell_45_17 ( BL17, BLN17, WL45);
sram_cell_6t_3 inst_cell_45_16 ( BL16, BLN16, WL45);
sram_cell_6t_3 inst_cell_45_15 ( BL15, BLN15, WL45);
sram_cell_6t_3 inst_cell_45_14 ( BL14, BLN14, WL45);
sram_cell_6t_3 inst_cell_45_13 ( BL13, BLN13, WL45);
sram_cell_6t_3 inst_cell_45_12 ( BL12, BLN12, WL45);
sram_cell_6t_3 inst_cell_45_11 ( BL11, BLN11, WL45);
sram_cell_6t_3 inst_cell_45_10 ( BL10, BLN10, WL45);
sram_cell_6t_3 inst_cell_45_9 ( BL9, BLN9, WL45);
sram_cell_6t_3 inst_cell_45_8 ( BL8, BLN8, WL45);
sram_cell_6t_3 inst_cell_45_7 ( BL7, BLN7, WL45);
sram_cell_6t_3 inst_cell_45_6 ( BL6, BLN6, WL45);
sram_cell_6t_3 inst_cell_45_5 ( BL5, BLN5, WL45);
sram_cell_6t_3 inst_cell_45_4 ( BL4, BLN4, WL45);
sram_cell_6t_3 inst_cell_45_3 ( BL3, BLN3, WL45);
sram_cell_6t_3 inst_cell_45_2 ( BL2, BLN2, WL45);
sram_cell_6t_3 inst_cell_45_1 ( BL1, BLN1, WL45);
sram_cell_6t_3 inst_cell_45_0 ( BL0, BLN0, WL45);
sram_cell_6t_3 inst_cell_44_39 ( BL39, BLN39, WL44);
sram_cell_6t_3 inst_cell_43_39 ( BL39, BLN39, WL43);
sram_cell_6t_3 inst_cell_44_38 ( BL38, BLN38, WL44);
sram_cell_6t_3 inst_cell_43_38 ( BL38, BLN38, WL43);
sram_cell_6t_3 inst_cell_44_37 ( BL37, BLN37, WL44);
sram_cell_6t_3 inst_cell_43_37 ( BL37, BLN37, WL43);
sram_cell_6t_3 inst_cell_44_36 ( BL36, BLN36, WL44);
sram_cell_6t_3 inst_cell_43_36 ( BL36, BLN36, WL43);
sram_cell_6t_3 inst_cell_44_35 ( BL35, BLN35, WL44);
sram_cell_6t_3 inst_cell_43_35 ( BL35, BLN35, WL43);
sram_cell_6t_3 inst_cell_44_34 ( BL34, BLN34, WL44);
sram_cell_6t_3 inst_cell_43_34 ( BL34, BLN34, WL43);
sram_cell_6t_3 inst_cell_44_33 ( BL33, BLN33, WL44);
sram_cell_6t_3 inst_cell_43_33 ( BL33, BLN33, WL43);
sram_cell_6t_3 inst_cell_44_32 ( BL32, BLN32, WL44);
sram_cell_6t_3 inst_cell_43_32 ( BL32, BLN32, WL43);
sram_cell_6t_3 inst_cell_44_31 ( BL31, BLN31, WL44);
sram_cell_6t_3 inst_cell_43_31 ( BL31, BLN31, WL43);
sram_cell_6t_3 inst_cell_44_30 ( BL30, BLN30, WL44);
sram_cell_6t_3 inst_cell_43_30 ( BL30, BLN30, WL43);
sram_cell_6t_3 inst_cell_44_29 ( BL29, BLN29, WL44);
sram_cell_6t_3 inst_cell_43_29 ( BL29, BLN29, WL43);
sram_cell_6t_3 inst_cell_44_28 ( BL28, BLN28, WL44);
sram_cell_6t_3 inst_cell_43_28 ( BL28, BLN28, WL43);
sram_cell_6t_3 inst_cell_44_27 ( BL27, BLN27, WL44);
sram_cell_6t_3 inst_cell_43_27 ( BL27, BLN27, WL43);
sram_cell_6t_3 inst_cell_44_26 ( BL26, BLN26, WL44);
sram_cell_6t_3 inst_cell_43_26 ( BL26, BLN26, WL43);
sram_cell_6t_3 inst_cell_44_25 ( BL25, BLN25, WL44);
sram_cell_6t_3 inst_cell_43_25 ( BL25, BLN25, WL43);
sram_cell_6t_3 inst_cell_44_24 ( BL24, BLN24, WL44);
sram_cell_6t_3 inst_cell_43_24 ( BL24, BLN24, WL43);
sram_cell_6t_3 inst_cell_44_23 ( BL23, BLN23, WL44);
sram_cell_6t_3 inst_cell_43_23 ( BL23, BLN23, WL43);
sram_cell_6t_3 inst_cell_44_22 ( BL22, BLN22, WL44);
sram_cell_6t_3 inst_cell_43_22 ( BL22, BLN22, WL43);
sram_cell_6t_3 inst_cell_44_21 ( BL21, BLN21, WL44);
sram_cell_6t_3 inst_cell_43_21 ( BL21, BLN21, WL43);
sram_cell_6t_3 inst_cell_44_20 ( BL20, BLN20, WL44);
sram_cell_6t_3 inst_cell_43_20 ( BL20, BLN20, WL43);
sram_cell_6t_3 inst_cell_44_19 ( BL19, BLN19, WL44);
sram_cell_6t_3 inst_cell_43_19 ( BL19, BLN19, WL43);
sram_cell_6t_3 inst_cell_44_18 ( BL18, BLN18, WL44);
sram_cell_6t_3 inst_cell_43_18 ( BL18, BLN18, WL43);
sram_cell_6t_3 inst_cell_44_17 ( BL17, BLN17, WL44);
sram_cell_6t_3 inst_cell_43_17 ( BL17, BLN17, WL43);
sram_cell_6t_3 inst_cell_44_16 ( BL16, BLN16, WL44);
sram_cell_6t_3 inst_cell_43_16 ( BL16, BLN16, WL43);
sram_cell_6t_3 inst_cell_44_15 ( BL15, BLN15, WL44);
sram_cell_6t_3 inst_cell_43_15 ( BL15, BLN15, WL43);
sram_cell_6t_3 inst_cell_44_14 ( BL14, BLN14, WL44);
sram_cell_6t_3 inst_cell_43_14 ( BL14, BLN14, WL43);
sram_cell_6t_3 inst_cell_44_13 ( BL13, BLN13, WL44);
sram_cell_6t_3 inst_cell_43_13 ( BL13, BLN13, WL43);
sram_cell_6t_3 inst_cell_44_12 ( BL12, BLN12, WL44);
sram_cell_6t_3 inst_cell_43_12 ( BL12, BLN12, WL43);
sram_cell_6t_3 inst_cell_44_11 ( BL11, BLN11, WL44);
sram_cell_6t_3 inst_cell_43_11 ( BL11, BLN11, WL43);
sram_cell_6t_3 inst_cell_44_10 ( BL10, BLN10, WL44);
sram_cell_6t_3 inst_cell_43_10 ( BL10, BLN10, WL43);
sram_cell_6t_3 inst_cell_44_9 ( BL9, BLN9, WL44);
sram_cell_6t_3 inst_cell_43_9 ( BL9, BLN9, WL43);
sram_cell_6t_3 inst_cell_44_8 ( BL8, BLN8, WL44);
sram_cell_6t_3 inst_cell_43_8 ( BL8, BLN8, WL43);
sram_cell_6t_3 inst_cell_44_7 ( BL7, BLN7, WL44);
sram_cell_6t_3 inst_cell_43_7 ( BL7, BLN7, WL43);
sram_cell_6t_3 inst_cell_44_6 ( BL6, BLN6, WL44);
sram_cell_6t_3 inst_cell_43_6 ( BL6, BLN6, WL43);
sram_cell_6t_3 inst_cell_44_5 ( BL5, BLN5, WL44);
sram_cell_6t_3 inst_cell_43_5 ( BL5, BLN5, WL43);
sram_cell_6t_3 inst_cell_44_4 ( BL4, BLN4, WL44);
sram_cell_6t_3 inst_cell_43_4 ( BL4, BLN4, WL43);
sram_cell_6t_3 inst_cell_44_3 ( BL3, BLN3, WL44);
sram_cell_6t_3 inst_cell_43_3 ( BL3, BLN3, WL43);
sram_cell_6t_3 inst_cell_44_2 ( BL2, BLN2, WL44);
sram_cell_6t_3 inst_cell_43_2 ( BL2, BLN2, WL43);
sram_cell_6t_3 inst_cell_44_1 ( BL1, BLN1, WL44);
sram_cell_6t_3 inst_cell_43_1 ( BL1, BLN1, WL43);
sram_cell_6t_3 inst_cell_44_0 ( BL0, BLN0, WL44);
sram_cell_6t_3 inst_cell_43_0 ( BL0, BLN0, WL43);
sram_cell_6t_3 inst_cell_44_63 ( BL63, BLN63, WL44);
sram_cell_6t_3 inst_cell_44_62 ( BL62, BLN62, WL44);
sram_cell_6t_3 inst_cell_44_61 ( BL61, BLN61, WL44);
sram_cell_6t_3 inst_cell_44_60 ( BL60, BLN60, WL44);
sram_cell_6t_3 inst_cell_44_59 ( BL59, BLN59, WL44);
sram_cell_6t_3 inst_cell_44_58 ( BL58, BLN58, WL44);
sram_cell_6t_3 inst_cell_44_57 ( BL57, BLN57, WL44);
sram_cell_6t_3 inst_cell_44_56 ( BL56, BLN56, WL44);
sram_cell_6t_3 inst_cell_44_55 ( BL55, BLN55, WL44);
sram_cell_6t_3 inst_cell_44_54 ( BL54, BLN54, WL44);
sram_cell_6t_3 inst_cell_44_53 ( BL53, BLN53, WL44);
sram_cell_6t_3 inst_cell_44_52 ( BL52, BLN52, WL44);
sram_cell_6t_3 inst_cell_44_51 ( BL51, BLN51, WL44);
sram_cell_6t_3 inst_cell_44_50 ( BL50, BLN50, WL44);
sram_cell_6t_3 inst_cell_44_49 ( BL49, BLN49, WL44);
sram_cell_6t_3 inst_cell_44_48 ( BL48, BLN48, WL44);
sram_cell_6t_3 inst_cell_44_47 ( BL47, BLN47, WL44);
sram_cell_6t_3 inst_cell_44_46 ( BL46, BLN46, WL44);
sram_cell_6t_3 inst_cell_44_45 ( BL45, BLN45, WL44);
sram_cell_6t_3 inst_cell_44_44 ( BL44, BLN44, WL44);
sram_cell_6t_3 inst_cell_44_43 ( BL43, BLN43, WL44);
sram_cell_6t_3 inst_cell_44_42 ( BL42, BLN42, WL44);
sram_cell_6t_3 inst_cell_44_41 ( BL41, BLN41, WL44);
sram_cell_6t_3 inst_cell_44_40 ( BL40, BLN40, WL44);
sram_cell_6t_3 inst_cell_43_63 ( BL63, BLN63, WL43);
sram_cell_6t_3 inst_cell_43_62 ( BL62, BLN62, WL43);
sram_cell_6t_3 inst_cell_43_61 ( BL61, BLN61, WL43);
sram_cell_6t_3 inst_cell_43_60 ( BL60, BLN60, WL43);
sram_cell_6t_3 inst_cell_43_59 ( BL59, BLN59, WL43);
sram_cell_6t_3 inst_cell_43_58 ( BL58, BLN58, WL43);
sram_cell_6t_3 inst_cell_43_57 ( BL57, BLN57, WL43);
sram_cell_6t_3 inst_cell_43_56 ( BL56, BLN56, WL43);
sram_cell_6t_3 inst_cell_43_55 ( BL55, BLN55, WL43);
sram_cell_6t_3 inst_cell_43_54 ( BL54, BLN54, WL43);
sram_cell_6t_3 inst_cell_43_53 ( BL53, BLN53, WL43);
sram_cell_6t_3 inst_cell_43_52 ( BL52, BLN52, WL43);
sram_cell_6t_3 inst_cell_43_51 ( BL51, BLN51, WL43);
sram_cell_6t_3 inst_cell_43_50 ( BL50, BLN50, WL43);
sram_cell_6t_3 inst_cell_43_49 ( BL49, BLN49, WL43);
sram_cell_6t_3 inst_cell_43_48 ( BL48, BLN48, WL43);
sram_cell_6t_3 inst_cell_43_47 ( BL47, BLN47, WL43);
sram_cell_6t_3 inst_cell_43_46 ( BL46, BLN46, WL43);
sram_cell_6t_3 inst_cell_43_45 ( BL45, BLN45, WL43);
sram_cell_6t_3 inst_cell_43_44 ( BL44, BLN44, WL43);
sram_cell_6t_3 inst_cell_43_43 ( BL43, BLN43, WL43);
sram_cell_6t_3 inst_cell_43_42 ( BL42, BLN42, WL43);
sram_cell_6t_3 inst_cell_43_41 ( BL41, BLN41, WL43);
sram_cell_6t_3 inst_cell_43_40 ( BL40, BLN40, WL43);
sram_cell_6t_3 inst_cell_42_63 ( BL63, BLN63, WL42);
sram_cell_6t_3 inst_cell_42_62 ( BL62, BLN62, WL42);
sram_cell_6t_3 inst_cell_42_61 ( BL61, BLN61, WL42);
sram_cell_6t_3 inst_cell_42_60 ( BL60, BLN60, WL42);
sram_cell_6t_3 inst_cell_42_59 ( BL59, BLN59, WL42);
sram_cell_6t_3 inst_cell_42_58 ( BL58, BLN58, WL42);
sram_cell_6t_3 inst_cell_42_57 ( BL57, BLN57, WL42);
sram_cell_6t_3 inst_cell_42_56 ( BL56, BLN56, WL42);
sram_cell_6t_3 inst_cell_42_55 ( BL55, BLN55, WL42);
sram_cell_6t_3 inst_cell_42_54 ( BL54, BLN54, WL42);
sram_cell_6t_3 inst_cell_42_53 ( BL53, BLN53, WL42);
sram_cell_6t_3 inst_cell_42_52 ( BL52, BLN52, WL42);
sram_cell_6t_3 inst_cell_42_51 ( BL51, BLN51, WL42);
sram_cell_6t_3 inst_cell_42_50 ( BL50, BLN50, WL42);
sram_cell_6t_3 inst_cell_42_49 ( BL49, BLN49, WL42);
sram_cell_6t_3 inst_cell_42_48 ( BL48, BLN48, WL42);
sram_cell_6t_3 inst_cell_42_47 ( BL47, BLN47, WL42);
sram_cell_6t_3 inst_cell_42_46 ( BL46, BLN46, WL42);
sram_cell_6t_3 inst_cell_42_45 ( BL45, BLN45, WL42);
sram_cell_6t_3 inst_cell_42_44 ( BL44, BLN44, WL42);
sram_cell_6t_3 inst_cell_42_43 ( BL43, BLN43, WL42);
sram_cell_6t_3 inst_cell_42_42 ( BL42, BLN42, WL42);
sram_cell_6t_3 inst_cell_42_41 ( BL41, BLN41, WL42);
sram_cell_6t_3 inst_cell_42_40 ( BL40, BLN40, WL42);
sram_cell_6t_3 inst_cell_42_15 ( BL15, BLN15, WL42);
sram_cell_6t_3 inst_cell_41_15 ( BL15, BLN15, WL41);
sram_cell_6t_3 inst_cell_42_14 ( BL14, BLN14, WL42);
sram_cell_6t_3 inst_cell_41_14 ( BL14, BLN14, WL41);
sram_cell_6t_3 inst_cell_42_13 ( BL13, BLN13, WL42);
sram_cell_6t_3 inst_cell_41_13 ( BL13, BLN13, WL41);
sram_cell_6t_3 inst_cell_42_12 ( BL12, BLN12, WL42);
sram_cell_6t_3 inst_cell_41_12 ( BL12, BLN12, WL41);
sram_cell_6t_3 inst_cell_42_11 ( BL11, BLN11, WL42);
sram_cell_6t_3 inst_cell_41_11 ( BL11, BLN11, WL41);
sram_cell_6t_3 inst_cell_42_10 ( BL10, BLN10, WL42);
sram_cell_6t_3 inst_cell_41_10 ( BL10, BLN10, WL41);
sram_cell_6t_3 inst_cell_42_9 ( BL9, BLN9, WL42);
sram_cell_6t_3 inst_cell_41_9 ( BL9, BLN9, WL41);
sram_cell_6t_3 inst_cell_42_8 ( BL8, BLN8, WL42);
sram_cell_6t_3 inst_cell_41_8 ( BL8, BLN8, WL41);
sram_cell_6t_3 inst_cell_42_7 ( BL7, BLN7, WL42);
sram_cell_6t_3 inst_cell_41_7 ( BL7, BLN7, WL41);
sram_cell_6t_3 inst_cell_42_6 ( BL6, BLN6, WL42);
sram_cell_6t_3 inst_cell_41_6 ( BL6, BLN6, WL41);
sram_cell_6t_3 inst_cell_42_5 ( BL5, BLN5, WL42);
sram_cell_6t_3 inst_cell_41_5 ( BL5, BLN5, WL41);
sram_cell_6t_3 inst_cell_42_4 ( BL4, BLN4, WL42);
sram_cell_6t_3 inst_cell_41_4 ( BL4, BLN4, WL41);
sram_cell_6t_3 inst_cell_42_3 ( BL3, BLN3, WL42);
sram_cell_6t_3 inst_cell_41_3 ( BL3, BLN3, WL41);
sram_cell_6t_3 inst_cell_42_2 ( BL2, BLN2, WL42);
sram_cell_6t_3 inst_cell_41_2 ( BL2, BLN2, WL41);
sram_cell_6t_3 inst_cell_42_1 ( BL1, BLN1, WL42);
sram_cell_6t_3 inst_cell_41_1 ( BL1, BLN1, WL41);
sram_cell_6t_3 inst_cell_42_0 ( BL0, BLN0, WL42);
sram_cell_6t_3 inst_cell_41_0 ( BL0, BLN0, WL41);
sram_cell_6t_3 inst_cell_41_63 ( BL63, BLN63, WL41);
sram_cell_6t_3 inst_cell_40_63 ( BL63, BLN63, WL40);
sram_cell_6t_3 inst_cell_41_62 ( BL62, BLN62, WL41);
sram_cell_6t_3 inst_cell_40_62 ( BL62, BLN62, WL40);
sram_cell_6t_3 inst_cell_41_61 ( BL61, BLN61, WL41);
sram_cell_6t_3 inst_cell_40_61 ( BL61, BLN61, WL40);
sram_cell_6t_3 inst_cell_41_60 ( BL60, BLN60, WL41);
sram_cell_6t_3 inst_cell_40_60 ( BL60, BLN60, WL40);
sram_cell_6t_3 inst_cell_41_59 ( BL59, BLN59, WL41);
sram_cell_6t_3 inst_cell_40_59 ( BL59, BLN59, WL40);
sram_cell_6t_3 inst_cell_41_58 ( BL58, BLN58, WL41);
sram_cell_6t_3 inst_cell_40_58 ( BL58, BLN58, WL40);
sram_cell_6t_3 inst_cell_41_57 ( BL57, BLN57, WL41);
sram_cell_6t_3 inst_cell_40_57 ( BL57, BLN57, WL40);
sram_cell_6t_3 inst_cell_41_56 ( BL56, BLN56, WL41);
sram_cell_6t_3 inst_cell_40_56 ( BL56, BLN56, WL40);
sram_cell_6t_3 inst_cell_41_55 ( BL55, BLN55, WL41);
sram_cell_6t_3 inst_cell_40_55 ( BL55, BLN55, WL40);
sram_cell_6t_3 inst_cell_41_54 ( BL54, BLN54, WL41);
sram_cell_6t_3 inst_cell_40_54 ( BL54, BLN54, WL40);
sram_cell_6t_3 inst_cell_41_53 ( BL53, BLN53, WL41);
sram_cell_6t_3 inst_cell_40_53 ( BL53, BLN53, WL40);
sram_cell_6t_3 inst_cell_41_52 ( BL52, BLN52, WL41);
sram_cell_6t_3 inst_cell_40_52 ( BL52, BLN52, WL40);
sram_cell_6t_3 inst_cell_41_51 ( BL51, BLN51, WL41);
sram_cell_6t_3 inst_cell_40_51 ( BL51, BLN51, WL40);
sram_cell_6t_3 inst_cell_41_50 ( BL50, BLN50, WL41);
sram_cell_6t_3 inst_cell_40_50 ( BL50, BLN50, WL40);
sram_cell_6t_3 inst_cell_41_49 ( BL49, BLN49, WL41);
sram_cell_6t_3 inst_cell_40_49 ( BL49, BLN49, WL40);
sram_cell_6t_3 inst_cell_41_48 ( BL48, BLN48, WL41);
sram_cell_6t_3 inst_cell_40_48 ( BL48, BLN48, WL40);
sram_cell_6t_3 inst_cell_41_47 ( BL47, BLN47, WL41);
sram_cell_6t_3 inst_cell_40_47 ( BL47, BLN47, WL40);
sram_cell_6t_3 inst_cell_41_46 ( BL46, BLN46, WL41);
sram_cell_6t_3 inst_cell_40_46 ( BL46, BLN46, WL40);
sram_cell_6t_3 inst_cell_41_45 ( BL45, BLN45, WL41);
sram_cell_6t_3 inst_cell_40_45 ( BL45, BLN45, WL40);
sram_cell_6t_3 inst_cell_41_44 ( BL44, BLN44, WL41);
sram_cell_6t_3 inst_cell_40_44 ( BL44, BLN44, WL40);
sram_cell_6t_3 inst_cell_41_43 ( BL43, BLN43, WL41);
sram_cell_6t_3 inst_cell_40_43 ( BL43, BLN43, WL40);
sram_cell_6t_3 inst_cell_41_42 ( BL42, BLN42, WL41);
sram_cell_6t_3 inst_cell_40_42 ( BL42, BLN42, WL40);
sram_cell_6t_3 inst_cell_41_41 ( BL41, BLN41, WL41);
sram_cell_6t_3 inst_cell_40_41 ( BL41, BLN41, WL40);
sram_cell_6t_3 inst_cell_41_40 ( BL40, BLN40, WL41);
sram_cell_6t_3 inst_cell_40_40 ( BL40, BLN40, WL40);
sram_cell_6t_3 inst_cell_42_39 ( BL39, BLN39, WL42);
sram_cell_6t_3 inst_cell_42_38 ( BL38, BLN38, WL42);
sram_cell_6t_3 inst_cell_42_37 ( BL37, BLN37, WL42);
sram_cell_6t_3 inst_cell_42_36 ( BL36, BLN36, WL42);
sram_cell_6t_3 inst_cell_42_35 ( BL35, BLN35, WL42);
sram_cell_6t_3 inst_cell_42_34 ( BL34, BLN34, WL42);
sram_cell_6t_3 inst_cell_42_33 ( BL33, BLN33, WL42);
sram_cell_6t_3 inst_cell_42_32 ( BL32, BLN32, WL42);
sram_cell_6t_3 inst_cell_42_31 ( BL31, BLN31, WL42);
sram_cell_6t_3 inst_cell_42_30 ( BL30, BLN30, WL42);
sram_cell_6t_3 inst_cell_42_29 ( BL29, BLN29, WL42);
sram_cell_6t_3 inst_cell_42_28 ( BL28, BLN28, WL42);
sram_cell_6t_3 inst_cell_42_27 ( BL27, BLN27, WL42);
sram_cell_6t_3 inst_cell_42_26 ( BL26, BLN26, WL42);
sram_cell_6t_3 inst_cell_42_25 ( BL25, BLN25, WL42);
sram_cell_6t_3 inst_cell_42_24 ( BL24, BLN24, WL42);
sram_cell_6t_3 inst_cell_42_23 ( BL23, BLN23, WL42);
sram_cell_6t_3 inst_cell_42_22 ( BL22, BLN22, WL42);
sram_cell_6t_3 inst_cell_42_21 ( BL21, BLN21, WL42);
sram_cell_6t_3 inst_cell_42_20 ( BL20, BLN20, WL42);
sram_cell_6t_3 inst_cell_42_19 ( BL19, BLN19, WL42);
sram_cell_6t_3 inst_cell_42_18 ( BL18, BLN18, WL42);
sram_cell_6t_3 inst_cell_42_17 ( BL17, BLN17, WL42);
sram_cell_6t_3 inst_cell_42_16 ( BL16, BLN16, WL42);
sram_cell_6t_3 inst_cell_41_39 ( BL39, BLN39, WL41);
sram_cell_6t_3 inst_cell_41_38 ( BL38, BLN38, WL41);
sram_cell_6t_3 inst_cell_41_37 ( BL37, BLN37, WL41);
sram_cell_6t_3 inst_cell_41_36 ( BL36, BLN36, WL41);
sram_cell_6t_3 inst_cell_41_35 ( BL35, BLN35, WL41);
sram_cell_6t_3 inst_cell_41_34 ( BL34, BLN34, WL41);
sram_cell_6t_3 inst_cell_41_33 ( BL33, BLN33, WL41);
sram_cell_6t_3 inst_cell_41_32 ( BL32, BLN32, WL41);
sram_cell_6t_3 inst_cell_41_31 ( BL31, BLN31, WL41);
sram_cell_6t_3 inst_cell_41_30 ( BL30, BLN30, WL41);
sram_cell_6t_3 inst_cell_41_29 ( BL29, BLN29, WL41);
sram_cell_6t_3 inst_cell_41_28 ( BL28, BLN28, WL41);
sram_cell_6t_3 inst_cell_41_27 ( BL27, BLN27, WL41);
sram_cell_6t_3 inst_cell_41_26 ( BL26, BLN26, WL41);
sram_cell_6t_3 inst_cell_41_25 ( BL25, BLN25, WL41);
sram_cell_6t_3 inst_cell_41_24 ( BL24, BLN24, WL41);
sram_cell_6t_3 inst_cell_41_23 ( BL23, BLN23, WL41);
sram_cell_6t_3 inst_cell_41_22 ( BL22, BLN22, WL41);
sram_cell_6t_3 inst_cell_41_21 ( BL21, BLN21, WL41);
sram_cell_6t_3 inst_cell_41_20 ( BL20, BLN20, WL41);
sram_cell_6t_3 inst_cell_41_19 ( BL19, BLN19, WL41);
sram_cell_6t_3 inst_cell_41_18 ( BL18, BLN18, WL41);
sram_cell_6t_3 inst_cell_41_17 ( BL17, BLN17, WL41);
sram_cell_6t_3 inst_cell_41_16 ( BL16, BLN16, WL41);
sram_cell_6t_3 inst_cell_40_39 ( BL39, BLN39, WL40);
sram_cell_6t_3 inst_cell_40_38 ( BL38, BLN38, WL40);
sram_cell_6t_3 inst_cell_40_37 ( BL37, BLN37, WL40);
sram_cell_6t_3 inst_cell_40_36 ( BL36, BLN36, WL40);
sram_cell_6t_3 inst_cell_40_35 ( BL35, BLN35, WL40);
sram_cell_6t_3 inst_cell_40_34 ( BL34, BLN34, WL40);
sram_cell_6t_3 inst_cell_40_33 ( BL33, BLN33, WL40);
sram_cell_6t_3 inst_cell_40_32 ( BL32, BLN32, WL40);
sram_cell_6t_3 inst_cell_40_31 ( BL31, BLN31, WL40);
sram_cell_6t_3 inst_cell_40_30 ( BL30, BLN30, WL40);
sram_cell_6t_3 inst_cell_40_29 ( BL29, BLN29, WL40);
sram_cell_6t_3 inst_cell_40_28 ( BL28, BLN28, WL40);
sram_cell_6t_3 inst_cell_40_27 ( BL27, BLN27, WL40);
sram_cell_6t_3 inst_cell_40_26 ( BL26, BLN26, WL40);
sram_cell_6t_3 inst_cell_40_25 ( BL25, BLN25, WL40);
sram_cell_6t_3 inst_cell_40_24 ( BL24, BLN24, WL40);
sram_cell_6t_3 inst_cell_40_23 ( BL23, BLN23, WL40);
sram_cell_6t_3 inst_cell_40_22 ( BL22, BLN22, WL40);
sram_cell_6t_3 inst_cell_40_21 ( BL21, BLN21, WL40);
sram_cell_6t_3 inst_cell_40_20 ( BL20, BLN20, WL40);
sram_cell_6t_3 inst_cell_40_19 ( BL19, BLN19, WL40);
sram_cell_6t_3 inst_cell_40_18 ( BL18, BLN18, WL40);
sram_cell_6t_3 inst_cell_40_17 ( BL17, BLN17, WL40);
sram_cell_6t_3 inst_cell_40_16 ( BL16, BLN16, WL40);
sram_cell_6t_3 inst_cell_39_62 ( BL62, BLN62, WL39);
sram_cell_6t_3 inst_cell_38_62 ( BL62, BLN62, WL38);
sram_cell_6t_3 inst_cell_39_61 ( BL61, BLN61, WL39);
sram_cell_6t_3 inst_cell_38_61 ( BL61, BLN61, WL38);
sram_cell_6t_3 inst_cell_39_60 ( BL60, BLN60, WL39);
sram_cell_6t_3 inst_cell_38_60 ( BL60, BLN60, WL38);
sram_cell_6t_3 inst_cell_39_59 ( BL59, BLN59, WL39);
sram_cell_6t_3 inst_cell_38_59 ( BL59, BLN59, WL38);
sram_cell_6t_3 inst_cell_39_58 ( BL58, BLN58, WL39);
sram_cell_6t_3 inst_cell_38_58 ( BL58, BLN58, WL38);
sram_cell_6t_3 inst_cell_39_57 ( BL57, BLN57, WL39);
sram_cell_6t_3 inst_cell_38_57 ( BL57, BLN57, WL38);
sram_cell_6t_3 inst_cell_39_56 ( BL56, BLN56, WL39);
sram_cell_6t_3 inst_cell_38_56 ( BL56, BLN56, WL38);
sram_cell_6t_3 inst_cell_39_55 ( BL55, BLN55, WL39);
sram_cell_6t_3 inst_cell_38_55 ( BL55, BLN55, WL38);
sram_cell_6t_3 inst_cell_39_54 ( BL54, BLN54, WL39);
sram_cell_6t_3 inst_cell_38_54 ( BL54, BLN54, WL38);
sram_cell_6t_3 inst_cell_39_53 ( BL53, BLN53, WL39);
sram_cell_6t_3 inst_cell_38_53 ( BL53, BLN53, WL38);
sram_cell_6t_3 inst_cell_39_52 ( BL52, BLN52, WL39);
sram_cell_6t_3 inst_cell_38_52 ( BL52, BLN52, WL38);
sram_cell_6t_3 inst_cell_39_51 ( BL51, BLN51, WL39);
sram_cell_6t_3 inst_cell_38_51 ( BL51, BLN51, WL38);
sram_cell_6t_3 inst_cell_39_50 ( BL50, BLN50, WL39);
sram_cell_6t_3 inst_cell_38_50 ( BL50, BLN50, WL38);
sram_cell_6t_3 inst_cell_39_49 ( BL49, BLN49, WL39);
sram_cell_6t_3 inst_cell_38_49 ( BL49, BLN49, WL38);
sram_cell_6t_3 inst_cell_39_48 ( BL48, BLN48, WL39);
sram_cell_6t_3 inst_cell_38_48 ( BL48, BLN48, WL38);
sram_cell_6t_3 inst_cell_39_47 ( BL47, BLN47, WL39);
sram_cell_6t_3 inst_cell_38_47 ( BL47, BLN47, WL38);
sram_cell_6t_3 inst_cell_39_46 ( BL46, BLN46, WL39);
sram_cell_6t_3 inst_cell_38_46 ( BL46, BLN46, WL38);
sram_cell_6t_3 inst_cell_39_45 ( BL45, BLN45, WL39);
sram_cell_6t_3 inst_cell_38_45 ( BL45, BLN45, WL38);
sram_cell_6t_3 inst_cell_39_44 ( BL44, BLN44, WL39);
sram_cell_6t_3 inst_cell_38_44 ( BL44, BLN44, WL38);
sram_cell_6t_3 inst_cell_39_43 ( BL43, BLN43, WL39);
sram_cell_6t_3 inst_cell_38_43 ( BL43, BLN43, WL38);
sram_cell_6t_3 inst_cell_39_42 ( BL42, BLN42, WL39);
sram_cell_6t_3 inst_cell_38_42 ( BL42, BLN42, WL38);
sram_cell_6t_3 inst_cell_39_41 ( BL41, BLN41, WL39);
sram_cell_6t_3 inst_cell_38_41 ( BL41, BLN41, WL38);
sram_cell_6t_3 inst_cell_39_40 ( BL40, BLN40, WL39);
sram_cell_6t_3 inst_cell_38_40 ( BL40, BLN40, WL38);
sram_cell_6t_3 inst_cell_39_39 ( BL39, BLN39, WL39);
sram_cell_6t_3 inst_cell_38_39 ( BL39, BLN39, WL38);
sram_cell_6t_3 inst_cell_39_38 ( BL38, BLN38, WL39);
sram_cell_6t_3 inst_cell_38_38 ( BL38, BLN38, WL38);
sram_cell_6t_3 inst_cell_39_37 ( BL37, BLN37, WL39);
sram_cell_6t_3 inst_cell_38_37 ( BL37, BLN37, WL38);
sram_cell_6t_3 inst_cell_39_36 ( BL36, BLN36, WL39);
sram_cell_6t_3 inst_cell_38_36 ( BL36, BLN36, WL38);
sram_cell_6t_3 inst_cell_39_35 ( BL35, BLN35, WL39);
sram_cell_6t_3 inst_cell_38_35 ( BL35, BLN35, WL38);
sram_cell_6t_3 inst_cell_39_34 ( BL34, BLN34, WL39);
sram_cell_6t_3 inst_cell_38_34 ( BL34, BLN34, WL38);
sram_cell_6t_3 inst_cell_39_33 ( BL33, BLN33, WL39);
sram_cell_6t_3 inst_cell_38_33 ( BL33, BLN33, WL38);
sram_cell_6t_3 inst_cell_39_32 ( BL32, BLN32, WL39);
sram_cell_6t_3 inst_cell_38_32 ( BL32, BLN32, WL38);
sram_cell_6t_3 inst_cell_39_31 ( BL31, BLN31, WL39);
sram_cell_6t_3 inst_cell_38_31 ( BL31, BLN31, WL38);
sram_cell_6t_3 inst_cell_39_30 ( BL30, BLN30, WL39);
sram_cell_6t_3 inst_cell_38_30 ( BL30, BLN30, WL38);
sram_cell_6t_3 inst_cell_39_29 ( BL29, BLN29, WL39);
sram_cell_6t_3 inst_cell_38_29 ( BL29, BLN29, WL38);
sram_cell_6t_3 inst_cell_39_28 ( BL28, BLN28, WL39);
sram_cell_6t_3 inst_cell_38_28 ( BL28, BLN28, WL38);
sram_cell_6t_3 inst_cell_39_27 ( BL27, BLN27, WL39);
sram_cell_6t_3 inst_cell_38_27 ( BL27, BLN27, WL38);
sram_cell_6t_3 inst_cell_39_26 ( BL26, BLN26, WL39);
sram_cell_6t_3 inst_cell_38_26 ( BL26, BLN26, WL38);
sram_cell_6t_3 inst_cell_39_25 ( BL25, BLN25, WL39);
sram_cell_6t_3 inst_cell_38_25 ( BL25, BLN25, WL38);
sram_cell_6t_3 inst_cell_39_24 ( BL24, BLN24, WL39);
sram_cell_6t_3 inst_cell_38_24 ( BL24, BLN24, WL38);
sram_cell_6t_3 inst_cell_39_23 ( BL23, BLN23, WL39);
sram_cell_6t_3 inst_cell_38_23 ( BL23, BLN23, WL38);
sram_cell_6t_3 inst_cell_39_22 ( BL22, BLN22, WL39);
sram_cell_6t_3 inst_cell_38_22 ( BL22, BLN22, WL38);
sram_cell_6t_3 inst_cell_39_21 ( BL21, BLN21, WL39);
sram_cell_6t_3 inst_cell_38_21 ( BL21, BLN21, WL38);
sram_cell_6t_3 inst_cell_39_20 ( BL20, BLN20, WL39);
sram_cell_6t_3 inst_cell_38_20 ( BL20, BLN20, WL38);
sram_cell_6t_3 inst_cell_39_19 ( BL19, BLN19, WL39);
sram_cell_6t_3 inst_cell_38_19 ( BL19, BLN19, WL38);
sram_cell_6t_3 inst_cell_39_18 ( BL18, BLN18, WL39);
sram_cell_6t_3 inst_cell_38_18 ( BL18, BLN18, WL38);
sram_cell_6t_3 inst_cell_39_17 ( BL17, BLN17, WL39);
sram_cell_6t_3 inst_cell_38_17 ( BL17, BLN17, WL38);
sram_cell_6t_3 inst_cell_39_16 ( BL16, BLN16, WL39);
sram_cell_6t_3 inst_cell_38_16 ( BL16, BLN16, WL38);
sram_cell_6t_3 inst_cell_40_15 ( BL15, BLN15, WL40);
sram_cell_6t_3 inst_cell_40_14 ( BL14, BLN14, WL40);
sram_cell_6t_3 inst_cell_40_13 ( BL13, BLN13, WL40);
sram_cell_6t_3 inst_cell_40_12 ( BL12, BLN12, WL40);
sram_cell_6t_3 inst_cell_40_11 ( BL11, BLN11, WL40);
sram_cell_6t_3 inst_cell_40_10 ( BL10, BLN10, WL40);
sram_cell_6t_3 inst_cell_40_9 ( BL9, BLN9, WL40);
sram_cell_6t_3 inst_cell_40_8 ( BL8, BLN8, WL40);
sram_cell_6t_3 inst_cell_40_7 ( BL7, BLN7, WL40);
sram_cell_6t_3 inst_cell_40_6 ( BL6, BLN6, WL40);
sram_cell_6t_3 inst_cell_40_5 ( BL5, BLN5, WL40);
sram_cell_6t_3 inst_cell_40_4 ( BL4, BLN4, WL40);
sram_cell_6t_3 inst_cell_40_3 ( BL3, BLN3, WL40);
sram_cell_6t_3 inst_cell_40_2 ( BL2, BLN2, WL40);
sram_cell_6t_3 inst_cell_40_1 ( BL1, BLN1, WL40);
sram_cell_6t_3 inst_cell_40_0 ( BL0, BLN0, WL40);
sram_cell_6t_3 inst_cell_39_63 ( BL63, BLN63, WL39);
sram_cell_6t_3 inst_cell_39_15 ( BL15, BLN15, WL39);
sram_cell_6t_3 inst_cell_39_14 ( BL14, BLN14, WL39);
sram_cell_6t_3 inst_cell_39_13 ( BL13, BLN13, WL39);
sram_cell_6t_3 inst_cell_39_12 ( BL12, BLN12, WL39);
sram_cell_6t_3 inst_cell_39_11 ( BL11, BLN11, WL39);
sram_cell_6t_3 inst_cell_39_10 ( BL10, BLN10, WL39);
sram_cell_6t_3 inst_cell_39_9 ( BL9, BLN9, WL39);
sram_cell_6t_3 inst_cell_39_8 ( BL8, BLN8, WL39);
sram_cell_6t_3 inst_cell_39_7 ( BL7, BLN7, WL39);
sram_cell_6t_3 inst_cell_39_6 ( BL6, BLN6, WL39);
sram_cell_6t_3 inst_cell_39_5 ( BL5, BLN5, WL39);
sram_cell_6t_3 inst_cell_39_4 ( BL4, BLN4, WL39);
sram_cell_6t_3 inst_cell_39_3 ( BL3, BLN3, WL39);
sram_cell_6t_3 inst_cell_39_2 ( BL2, BLN2, WL39);
sram_cell_6t_3 inst_cell_39_1 ( BL1, BLN1, WL39);
sram_cell_6t_3 inst_cell_39_0 ( BL0, BLN0, WL39);
sram_cell_6t_3 inst_cell_38_63 ( BL63, BLN63, WL38);
sram_cell_6t_3 inst_cell_38_15 ( BL15, BLN15, WL38);
sram_cell_6t_3 inst_cell_38_14 ( BL14, BLN14, WL38);
sram_cell_6t_3 inst_cell_38_13 ( BL13, BLN13, WL38);
sram_cell_6t_3 inst_cell_38_12 ( BL12, BLN12, WL38);
sram_cell_6t_3 inst_cell_38_11 ( BL11, BLN11, WL38);
sram_cell_6t_3 inst_cell_38_10 ( BL10, BLN10, WL38);
sram_cell_6t_3 inst_cell_38_9 ( BL9, BLN9, WL38);
sram_cell_6t_3 inst_cell_38_8 ( BL8, BLN8, WL38);
sram_cell_6t_3 inst_cell_38_7 ( BL7, BLN7, WL38);
sram_cell_6t_3 inst_cell_38_6 ( BL6, BLN6, WL38);
sram_cell_6t_3 inst_cell_38_5 ( BL5, BLN5, WL38);
sram_cell_6t_3 inst_cell_38_4 ( BL4, BLN4, WL38);
sram_cell_6t_3 inst_cell_38_3 ( BL3, BLN3, WL38);
sram_cell_6t_3 inst_cell_38_2 ( BL2, BLN2, WL38);
sram_cell_6t_3 inst_cell_38_1 ( BL1, BLN1, WL38);
sram_cell_6t_3 inst_cell_38_0 ( BL0, BLN0, WL38);
sram_cell_6t_3 inst_cell_37_63 ( BL63, BLN63, WL37);
sram_cell_6t_3 inst_cell_37_31 ( BL31, BLN31, WL37);
sram_cell_6t_3 inst_cell_36_31 ( BL31, BLN31, WL36);
sram_cell_6t_3 inst_cell_37_30 ( BL30, BLN30, WL37);
sram_cell_6t_3 inst_cell_36_30 ( BL30, BLN30, WL36);
sram_cell_6t_3 inst_cell_37_29 ( BL29, BLN29, WL37);
sram_cell_6t_3 inst_cell_36_29 ( BL29, BLN29, WL36);
sram_cell_6t_3 inst_cell_37_28 ( BL28, BLN28, WL37);
sram_cell_6t_3 inst_cell_36_28 ( BL28, BLN28, WL36);
sram_cell_6t_3 inst_cell_37_27 ( BL27, BLN27, WL37);
sram_cell_6t_3 inst_cell_36_27 ( BL27, BLN27, WL36);
sram_cell_6t_3 inst_cell_37_26 ( BL26, BLN26, WL37);
sram_cell_6t_3 inst_cell_36_26 ( BL26, BLN26, WL36);
sram_cell_6t_3 inst_cell_37_25 ( BL25, BLN25, WL37);
sram_cell_6t_3 inst_cell_36_25 ( BL25, BLN25, WL36);
sram_cell_6t_3 inst_cell_37_24 ( BL24, BLN24, WL37);
sram_cell_6t_3 inst_cell_36_24 ( BL24, BLN24, WL36);
sram_cell_6t_3 inst_cell_37_23 ( BL23, BLN23, WL37);
sram_cell_6t_3 inst_cell_36_23 ( BL23, BLN23, WL36);
sram_cell_6t_3 inst_cell_37_22 ( BL22, BLN22, WL37);
sram_cell_6t_3 inst_cell_36_22 ( BL22, BLN22, WL36);
sram_cell_6t_3 inst_cell_37_21 ( BL21, BLN21, WL37);
sram_cell_6t_3 inst_cell_36_21 ( BL21, BLN21, WL36);
sram_cell_6t_3 inst_cell_37_20 ( BL20, BLN20, WL37);
sram_cell_6t_3 inst_cell_36_20 ( BL20, BLN20, WL36);
sram_cell_6t_3 inst_cell_37_19 ( BL19, BLN19, WL37);
sram_cell_6t_3 inst_cell_36_19 ( BL19, BLN19, WL36);
sram_cell_6t_3 inst_cell_37_18 ( BL18, BLN18, WL37);
sram_cell_6t_3 inst_cell_36_18 ( BL18, BLN18, WL36);
sram_cell_6t_3 inst_cell_37_17 ( BL17, BLN17, WL37);
sram_cell_6t_3 inst_cell_36_17 ( BL17, BLN17, WL36);
sram_cell_6t_3 inst_cell_37_16 ( BL16, BLN16, WL37);
sram_cell_6t_3 inst_cell_36_16 ( BL16, BLN16, WL36);
sram_cell_6t_3 inst_cell_37_15 ( BL15, BLN15, WL37);
sram_cell_6t_3 inst_cell_36_15 ( BL15, BLN15, WL36);
sram_cell_6t_3 inst_cell_37_14 ( BL14, BLN14, WL37);
sram_cell_6t_3 inst_cell_36_14 ( BL14, BLN14, WL36);
sram_cell_6t_3 inst_cell_37_13 ( BL13, BLN13, WL37);
sram_cell_6t_3 inst_cell_36_13 ( BL13, BLN13, WL36);
sram_cell_6t_3 inst_cell_37_12 ( BL12, BLN12, WL37);
sram_cell_6t_3 inst_cell_36_12 ( BL12, BLN12, WL36);
sram_cell_6t_3 inst_cell_37_11 ( BL11, BLN11, WL37);
sram_cell_6t_3 inst_cell_36_11 ( BL11, BLN11, WL36);
sram_cell_6t_3 inst_cell_37_10 ( BL10, BLN10, WL37);
sram_cell_6t_3 inst_cell_36_10 ( BL10, BLN10, WL36);
sram_cell_6t_3 inst_cell_37_9 ( BL9, BLN9, WL37);
sram_cell_6t_3 inst_cell_36_9 ( BL9, BLN9, WL36);
sram_cell_6t_3 inst_cell_37_8 ( BL8, BLN8, WL37);
sram_cell_6t_3 inst_cell_36_8 ( BL8, BLN8, WL36);
sram_cell_6t_3 inst_cell_37_7 ( BL7, BLN7, WL37);
sram_cell_6t_3 inst_cell_36_7 ( BL7, BLN7, WL36);
sram_cell_6t_3 inst_cell_37_6 ( BL6, BLN6, WL37);
sram_cell_6t_3 inst_cell_36_6 ( BL6, BLN6, WL36);
sram_cell_6t_3 inst_cell_37_5 ( BL5, BLN5, WL37);
sram_cell_6t_3 inst_cell_36_5 ( BL5, BLN5, WL36);
sram_cell_6t_3 inst_cell_37_4 ( BL4, BLN4, WL37);
sram_cell_6t_3 inst_cell_36_4 ( BL4, BLN4, WL36);
sram_cell_6t_3 inst_cell_37_3 ( BL3, BLN3, WL37);
sram_cell_6t_3 inst_cell_36_3 ( BL3, BLN3, WL36);
sram_cell_6t_3 inst_cell_37_2 ( BL2, BLN2, WL37);
sram_cell_6t_3 inst_cell_36_2 ( BL2, BLN2, WL36);
sram_cell_6t_3 inst_cell_37_1 ( BL1, BLN1, WL37);
sram_cell_6t_3 inst_cell_36_1 ( BL1, BLN1, WL36);
sram_cell_6t_3 inst_cell_37_0 ( BL0, BLN0, WL37);
sram_cell_6t_3 inst_cell_36_0 ( BL0, BLN0, WL36);
sram_cell_6t_3 inst_cell_36_63 ( BL63, BLN63, WL36);
sram_cell_6t_3 inst_cell_35_63 ( BL63, BLN63, WL35);
sram_cell_6t_3 inst_cell_37_62 ( BL62, BLN62, WL37);
sram_cell_6t_3 inst_cell_37_61 ( BL61, BLN61, WL37);
sram_cell_6t_3 inst_cell_37_60 ( BL60, BLN60, WL37);
sram_cell_6t_3 inst_cell_37_59 ( BL59, BLN59, WL37);
sram_cell_6t_3 inst_cell_37_58 ( BL58, BLN58, WL37);
sram_cell_6t_3 inst_cell_37_57 ( BL57, BLN57, WL37);
sram_cell_6t_3 inst_cell_37_56 ( BL56, BLN56, WL37);
sram_cell_6t_3 inst_cell_37_55 ( BL55, BLN55, WL37);
sram_cell_6t_3 inst_cell_37_54 ( BL54, BLN54, WL37);
sram_cell_6t_3 inst_cell_37_53 ( BL53, BLN53, WL37);
sram_cell_6t_3 inst_cell_37_52 ( BL52, BLN52, WL37);
sram_cell_6t_3 inst_cell_37_51 ( BL51, BLN51, WL37);
sram_cell_6t_3 inst_cell_37_50 ( BL50, BLN50, WL37);
sram_cell_6t_3 inst_cell_37_49 ( BL49, BLN49, WL37);
sram_cell_6t_3 inst_cell_37_48 ( BL48, BLN48, WL37);
sram_cell_6t_3 inst_cell_37_47 ( BL47, BLN47, WL37);
sram_cell_6t_3 inst_cell_37_46 ( BL46, BLN46, WL37);
sram_cell_6t_3 inst_cell_37_45 ( BL45, BLN45, WL37);
sram_cell_6t_3 inst_cell_37_44 ( BL44, BLN44, WL37);
sram_cell_6t_3 inst_cell_37_43 ( BL43, BLN43, WL37);
sram_cell_6t_3 inst_cell_37_42 ( BL42, BLN42, WL37);
sram_cell_6t_3 inst_cell_37_41 ( BL41, BLN41, WL37);
sram_cell_6t_3 inst_cell_37_40 ( BL40, BLN40, WL37);
sram_cell_6t_3 inst_cell_37_39 ( BL39, BLN39, WL37);
sram_cell_6t_3 inst_cell_37_38 ( BL38, BLN38, WL37);
sram_cell_6t_3 inst_cell_37_37 ( BL37, BLN37, WL37);
sram_cell_6t_3 inst_cell_37_36 ( BL36, BLN36, WL37);
sram_cell_6t_3 inst_cell_37_35 ( BL35, BLN35, WL37);
sram_cell_6t_3 inst_cell_37_34 ( BL34, BLN34, WL37);
sram_cell_6t_3 inst_cell_37_33 ( BL33, BLN33, WL37);
sram_cell_6t_3 inst_cell_37_32 ( BL32, BLN32, WL37);
sram_cell_6t_3 inst_cell_36_62 ( BL62, BLN62, WL36);
sram_cell_6t_3 inst_cell_36_61 ( BL61, BLN61, WL36);
sram_cell_6t_3 inst_cell_36_60 ( BL60, BLN60, WL36);
sram_cell_6t_3 inst_cell_36_59 ( BL59, BLN59, WL36);
sram_cell_6t_3 inst_cell_36_58 ( BL58, BLN58, WL36);
sram_cell_6t_3 inst_cell_36_57 ( BL57, BLN57, WL36);
sram_cell_6t_3 inst_cell_36_56 ( BL56, BLN56, WL36);
sram_cell_6t_3 inst_cell_36_55 ( BL55, BLN55, WL36);
sram_cell_6t_3 inst_cell_36_54 ( BL54, BLN54, WL36);
sram_cell_6t_3 inst_cell_36_53 ( BL53, BLN53, WL36);
sram_cell_6t_3 inst_cell_36_52 ( BL52, BLN52, WL36);
sram_cell_6t_3 inst_cell_36_51 ( BL51, BLN51, WL36);
sram_cell_6t_3 inst_cell_36_50 ( BL50, BLN50, WL36);
sram_cell_6t_3 inst_cell_36_49 ( BL49, BLN49, WL36);
sram_cell_6t_3 inst_cell_36_48 ( BL48, BLN48, WL36);
sram_cell_6t_3 inst_cell_36_47 ( BL47, BLN47, WL36);
sram_cell_6t_3 inst_cell_36_46 ( BL46, BLN46, WL36);
sram_cell_6t_3 inst_cell_36_45 ( BL45, BLN45, WL36);
sram_cell_6t_3 inst_cell_36_44 ( BL44, BLN44, WL36);
sram_cell_6t_3 inst_cell_36_43 ( BL43, BLN43, WL36);
sram_cell_6t_3 inst_cell_36_42 ( BL42, BLN42, WL36);
sram_cell_6t_3 inst_cell_36_41 ( BL41, BLN41, WL36);
sram_cell_6t_3 inst_cell_36_40 ( BL40, BLN40, WL36);
sram_cell_6t_3 inst_cell_36_39 ( BL39, BLN39, WL36);
sram_cell_6t_3 inst_cell_36_38 ( BL38, BLN38, WL36);
sram_cell_6t_3 inst_cell_36_37 ( BL37, BLN37, WL36);
sram_cell_6t_3 inst_cell_36_36 ( BL36, BLN36, WL36);
sram_cell_6t_3 inst_cell_36_35 ( BL35, BLN35, WL36);
sram_cell_6t_3 inst_cell_36_34 ( BL34, BLN34, WL36);
sram_cell_6t_3 inst_cell_36_33 ( BL33, BLN33, WL36);
sram_cell_6t_3 inst_cell_36_32 ( BL32, BLN32, WL36);
sram_cell_6t_3 inst_cell_35_62 ( BL62, BLN62, WL35);
sram_cell_6t_3 inst_cell_35_61 ( BL61, BLN61, WL35);
sram_cell_6t_3 inst_cell_35_60 ( BL60, BLN60, WL35);
sram_cell_6t_3 inst_cell_35_59 ( BL59, BLN59, WL35);
sram_cell_6t_3 inst_cell_35_58 ( BL58, BLN58, WL35);
sram_cell_6t_3 inst_cell_35_57 ( BL57, BLN57, WL35);
sram_cell_6t_3 inst_cell_35_56 ( BL56, BLN56, WL35);
sram_cell_6t_3 inst_cell_35_55 ( BL55, BLN55, WL35);
sram_cell_6t_3 inst_cell_35_54 ( BL54, BLN54, WL35);
sram_cell_6t_3 inst_cell_35_53 ( BL53, BLN53, WL35);
sram_cell_6t_3 inst_cell_35_52 ( BL52, BLN52, WL35);
sram_cell_6t_3 inst_cell_35_51 ( BL51, BLN51, WL35);
sram_cell_6t_3 inst_cell_35_50 ( BL50, BLN50, WL35);
sram_cell_6t_3 inst_cell_35_49 ( BL49, BLN49, WL35);
sram_cell_6t_3 inst_cell_35_48 ( BL48, BLN48, WL35);
sram_cell_6t_3 inst_cell_35_47 ( BL47, BLN47, WL35);
sram_cell_6t_3 inst_cell_35_46 ( BL46, BLN46, WL35);
sram_cell_6t_3 inst_cell_35_45 ( BL45, BLN45, WL35);
sram_cell_6t_3 inst_cell_35_44 ( BL44, BLN44, WL35);
sram_cell_6t_3 inst_cell_35_43 ( BL43, BLN43, WL35);
sram_cell_6t_3 inst_cell_35_42 ( BL42, BLN42, WL35);
sram_cell_6t_3 inst_cell_35_41 ( BL41, BLN41, WL35);
sram_cell_6t_3 inst_cell_35_40 ( BL40, BLN40, WL35);
sram_cell_6t_3 inst_cell_35_39 ( BL39, BLN39, WL35);
sram_cell_6t_3 inst_cell_35_38 ( BL38, BLN38, WL35);
sram_cell_6t_3 inst_cell_35_37 ( BL37, BLN37, WL35);
sram_cell_6t_3 inst_cell_35_36 ( BL36, BLN36, WL35);
sram_cell_6t_3 inst_cell_35_35 ( BL35, BLN35, WL35);
sram_cell_6t_3 inst_cell_35_34 ( BL34, BLN34, WL35);
sram_cell_6t_3 inst_cell_35_33 ( BL33, BLN33, WL35);
sram_cell_6t_3 inst_cell_35_32 ( BL32, BLN32, WL35);
sram_cell_6t_3 inst_cell_35_7 ( BL7, BLN7, WL35);
sram_cell_6t_3 inst_cell_34_7 ( BL7, BLN7, WL34);
sram_cell_6t_3 inst_cell_35_6 ( BL6, BLN6, WL35);
sram_cell_6t_3 inst_cell_34_6 ( BL6, BLN6, WL34);
sram_cell_6t_3 inst_cell_35_5 ( BL5, BLN5, WL35);
sram_cell_6t_3 inst_cell_34_5 ( BL5, BLN5, WL34);
sram_cell_6t_3 inst_cell_35_4 ( BL4, BLN4, WL35);
sram_cell_6t_3 inst_cell_34_4 ( BL4, BLN4, WL34);
sram_cell_6t_3 inst_cell_35_3 ( BL3, BLN3, WL35);
sram_cell_6t_3 inst_cell_34_3 ( BL3, BLN3, WL34);
sram_cell_6t_3 inst_cell_35_2 ( BL2, BLN2, WL35);
sram_cell_6t_3 inst_cell_34_2 ( BL2, BLN2, WL34);
sram_cell_6t_3 inst_cell_35_1 ( BL1, BLN1, WL35);
sram_cell_6t_3 inst_cell_34_1 ( BL1, BLN1, WL34);
sram_cell_6t_3 inst_cell_35_0 ( BL0, BLN0, WL35);
sram_cell_6t_3 inst_cell_34_0 ( BL0, BLN0, WL34);
sram_cell_6t_3 inst_cell_34_63 ( BL63, BLN63, WL34);
sram_cell_6t_3 inst_cell_33_63 ( BL63, BLN63, WL33);
sram_cell_6t_3 inst_cell_34_62 ( BL62, BLN62, WL34);
sram_cell_6t_3 inst_cell_33_62 ( BL62, BLN62, WL33);
sram_cell_6t_3 inst_cell_34_61 ( BL61, BLN61, WL34);
sram_cell_6t_3 inst_cell_33_61 ( BL61, BLN61, WL33);
sram_cell_6t_3 inst_cell_34_60 ( BL60, BLN60, WL34);
sram_cell_6t_3 inst_cell_33_60 ( BL60, BLN60, WL33);
sram_cell_6t_3 inst_cell_34_59 ( BL59, BLN59, WL34);
sram_cell_6t_3 inst_cell_33_59 ( BL59, BLN59, WL33);
sram_cell_6t_3 inst_cell_34_58 ( BL58, BLN58, WL34);
sram_cell_6t_3 inst_cell_33_58 ( BL58, BLN58, WL33);
sram_cell_6t_3 inst_cell_34_57 ( BL57, BLN57, WL34);
sram_cell_6t_3 inst_cell_33_57 ( BL57, BLN57, WL33);
sram_cell_6t_3 inst_cell_34_56 ( BL56, BLN56, WL34);
sram_cell_6t_3 inst_cell_33_56 ( BL56, BLN56, WL33);
sram_cell_6t_3 inst_cell_34_55 ( BL55, BLN55, WL34);
sram_cell_6t_3 inst_cell_33_55 ( BL55, BLN55, WL33);
sram_cell_6t_3 inst_cell_34_54 ( BL54, BLN54, WL34);
sram_cell_6t_3 inst_cell_33_54 ( BL54, BLN54, WL33);
sram_cell_6t_3 inst_cell_34_53 ( BL53, BLN53, WL34);
sram_cell_6t_3 inst_cell_33_53 ( BL53, BLN53, WL33);
sram_cell_6t_3 inst_cell_34_52 ( BL52, BLN52, WL34);
sram_cell_6t_3 inst_cell_33_52 ( BL52, BLN52, WL33);
sram_cell_6t_3 inst_cell_34_51 ( BL51, BLN51, WL34);
sram_cell_6t_3 inst_cell_33_51 ( BL51, BLN51, WL33);
sram_cell_6t_3 inst_cell_34_50 ( BL50, BLN50, WL34);
sram_cell_6t_3 inst_cell_33_50 ( BL50, BLN50, WL33);
sram_cell_6t_3 inst_cell_34_49 ( BL49, BLN49, WL34);
sram_cell_6t_3 inst_cell_33_49 ( BL49, BLN49, WL33);
sram_cell_6t_3 inst_cell_34_48 ( BL48, BLN48, WL34);
sram_cell_6t_3 inst_cell_33_48 ( BL48, BLN48, WL33);
sram_cell_6t_3 inst_cell_34_47 ( BL47, BLN47, WL34);
sram_cell_6t_3 inst_cell_33_47 ( BL47, BLN47, WL33);
sram_cell_6t_3 inst_cell_34_46 ( BL46, BLN46, WL34);
sram_cell_6t_3 inst_cell_33_46 ( BL46, BLN46, WL33);
sram_cell_6t_3 inst_cell_34_45 ( BL45, BLN45, WL34);
sram_cell_6t_3 inst_cell_33_45 ( BL45, BLN45, WL33);
sram_cell_6t_3 inst_cell_34_44 ( BL44, BLN44, WL34);
sram_cell_6t_3 inst_cell_33_44 ( BL44, BLN44, WL33);
sram_cell_6t_3 inst_cell_34_43 ( BL43, BLN43, WL34);
sram_cell_6t_3 inst_cell_33_43 ( BL43, BLN43, WL33);
sram_cell_6t_3 inst_cell_34_42 ( BL42, BLN42, WL34);
sram_cell_6t_3 inst_cell_33_42 ( BL42, BLN42, WL33);
sram_cell_6t_3 inst_cell_34_41 ( BL41, BLN41, WL34);
sram_cell_6t_3 inst_cell_33_41 ( BL41, BLN41, WL33);
sram_cell_6t_3 inst_cell_34_40 ( BL40, BLN40, WL34);
sram_cell_6t_3 inst_cell_33_40 ( BL40, BLN40, WL33);
sram_cell_6t_3 inst_cell_34_39 ( BL39, BLN39, WL34);
sram_cell_6t_3 inst_cell_33_39 ( BL39, BLN39, WL33);
sram_cell_6t_3 inst_cell_34_38 ( BL38, BLN38, WL34);
sram_cell_6t_3 inst_cell_33_38 ( BL38, BLN38, WL33);
sram_cell_6t_3 inst_cell_34_37 ( BL37, BLN37, WL34);
sram_cell_6t_3 inst_cell_33_37 ( BL37, BLN37, WL33);
sram_cell_6t_3 inst_cell_34_36 ( BL36, BLN36, WL34);
sram_cell_6t_3 inst_cell_33_36 ( BL36, BLN36, WL33);
sram_cell_6t_3 inst_cell_34_35 ( BL35, BLN35, WL34);
sram_cell_6t_3 inst_cell_33_35 ( BL35, BLN35, WL33);
sram_cell_6t_3 inst_cell_34_34 ( BL34, BLN34, WL34);
sram_cell_6t_3 inst_cell_33_34 ( BL34, BLN34, WL33);
sram_cell_6t_3 inst_cell_34_33 ( BL33, BLN33, WL34);
sram_cell_6t_3 inst_cell_33_33 ( BL33, BLN33, WL33);
sram_cell_6t_3 inst_cell_34_32 ( BL32, BLN32, WL34);
sram_cell_6t_3 inst_cell_33_32 ( BL32, BLN32, WL33);
sram_cell_6t_3 inst_cell_35_31 ( BL31, BLN31, WL35);
sram_cell_6t_3 inst_cell_35_30 ( BL30, BLN30, WL35);
sram_cell_6t_3 inst_cell_35_29 ( BL29, BLN29, WL35);
sram_cell_6t_3 inst_cell_35_28 ( BL28, BLN28, WL35);
sram_cell_6t_3 inst_cell_35_27 ( BL27, BLN27, WL35);
sram_cell_6t_3 inst_cell_35_26 ( BL26, BLN26, WL35);
sram_cell_6t_3 inst_cell_35_25 ( BL25, BLN25, WL35);
sram_cell_6t_3 inst_cell_35_24 ( BL24, BLN24, WL35);
sram_cell_6t_3 inst_cell_35_23 ( BL23, BLN23, WL35);
sram_cell_6t_3 inst_cell_35_22 ( BL22, BLN22, WL35);
sram_cell_6t_3 inst_cell_35_21 ( BL21, BLN21, WL35);
sram_cell_6t_3 inst_cell_35_20 ( BL20, BLN20, WL35);
sram_cell_6t_3 inst_cell_35_19 ( BL19, BLN19, WL35);
sram_cell_6t_3 inst_cell_35_18 ( BL18, BLN18, WL35);
sram_cell_6t_3 inst_cell_35_17 ( BL17, BLN17, WL35);
sram_cell_6t_3 inst_cell_35_16 ( BL16, BLN16, WL35);
sram_cell_6t_3 inst_cell_35_15 ( BL15, BLN15, WL35);
sram_cell_6t_3 inst_cell_35_14 ( BL14, BLN14, WL35);
sram_cell_6t_3 inst_cell_35_13 ( BL13, BLN13, WL35);
sram_cell_6t_3 inst_cell_35_12 ( BL12, BLN12, WL35);
sram_cell_6t_3 inst_cell_35_11 ( BL11, BLN11, WL35);
sram_cell_6t_3 inst_cell_35_10 ( BL10, BLN10, WL35);
sram_cell_6t_3 inst_cell_35_9 ( BL9, BLN9, WL35);
sram_cell_6t_3 inst_cell_35_8 ( BL8, BLN8, WL35);
sram_cell_6t_3 inst_cell_34_31 ( BL31, BLN31, WL34);
sram_cell_6t_3 inst_cell_34_30 ( BL30, BLN30, WL34);
sram_cell_6t_3 inst_cell_34_29 ( BL29, BLN29, WL34);
sram_cell_6t_3 inst_cell_34_28 ( BL28, BLN28, WL34);
sram_cell_6t_3 inst_cell_34_27 ( BL27, BLN27, WL34);
sram_cell_6t_3 inst_cell_34_26 ( BL26, BLN26, WL34);
sram_cell_6t_3 inst_cell_34_25 ( BL25, BLN25, WL34);
sram_cell_6t_3 inst_cell_34_24 ( BL24, BLN24, WL34);
sram_cell_6t_3 inst_cell_34_23 ( BL23, BLN23, WL34);
sram_cell_6t_3 inst_cell_34_22 ( BL22, BLN22, WL34);
sram_cell_6t_3 inst_cell_34_21 ( BL21, BLN21, WL34);
sram_cell_6t_3 inst_cell_34_20 ( BL20, BLN20, WL34);
sram_cell_6t_3 inst_cell_34_19 ( BL19, BLN19, WL34);
sram_cell_6t_3 inst_cell_34_18 ( BL18, BLN18, WL34);
sram_cell_6t_3 inst_cell_34_17 ( BL17, BLN17, WL34);
sram_cell_6t_3 inst_cell_34_16 ( BL16, BLN16, WL34);
sram_cell_6t_3 inst_cell_34_15 ( BL15, BLN15, WL34);
sram_cell_6t_3 inst_cell_34_14 ( BL14, BLN14, WL34);
sram_cell_6t_3 inst_cell_34_13 ( BL13, BLN13, WL34);
sram_cell_6t_3 inst_cell_34_12 ( BL12, BLN12, WL34);
sram_cell_6t_3 inst_cell_34_11 ( BL11, BLN11, WL34);
sram_cell_6t_3 inst_cell_34_10 ( BL10, BLN10, WL34);
sram_cell_6t_3 inst_cell_34_9 ( BL9, BLN9, WL34);
sram_cell_6t_3 inst_cell_34_8 ( BL8, BLN8, WL34);
sram_cell_6t_3 inst_cell_33_31 ( BL31, BLN31, WL33);
sram_cell_6t_3 inst_cell_33_30 ( BL30, BLN30, WL33);
sram_cell_6t_3 inst_cell_33_29 ( BL29, BLN29, WL33);
sram_cell_6t_3 inst_cell_33_28 ( BL28, BLN28, WL33);
sram_cell_6t_3 inst_cell_33_27 ( BL27, BLN27, WL33);
sram_cell_6t_3 inst_cell_33_26 ( BL26, BLN26, WL33);
sram_cell_6t_3 inst_cell_33_25 ( BL25, BLN25, WL33);
sram_cell_6t_3 inst_cell_33_24 ( BL24, BLN24, WL33);
sram_cell_6t_3 inst_cell_33_23 ( BL23, BLN23, WL33);
sram_cell_6t_3 inst_cell_33_22 ( BL22, BLN22, WL33);
sram_cell_6t_3 inst_cell_33_21 ( BL21, BLN21, WL33);
sram_cell_6t_3 inst_cell_33_20 ( BL20, BLN20, WL33);
sram_cell_6t_3 inst_cell_33_19 ( BL19, BLN19, WL33);
sram_cell_6t_3 inst_cell_33_18 ( BL18, BLN18, WL33);
sram_cell_6t_3 inst_cell_33_17 ( BL17, BLN17, WL33);
sram_cell_6t_3 inst_cell_33_16 ( BL16, BLN16, WL33);
sram_cell_6t_3 inst_cell_33_15 ( BL15, BLN15, WL33);
sram_cell_6t_3 inst_cell_33_14 ( BL14, BLN14, WL33);
sram_cell_6t_3 inst_cell_33_13 ( BL13, BLN13, WL33);
sram_cell_6t_3 inst_cell_33_12 ( BL12, BLN12, WL33);
sram_cell_6t_3 inst_cell_33_11 ( BL11, BLN11, WL33);
sram_cell_6t_3 inst_cell_33_10 ( BL10, BLN10, WL33);
sram_cell_6t_3 inst_cell_33_9 ( BL9, BLN9, WL33);
sram_cell_6t_3 inst_cell_33_8 ( BL8, BLN8, WL33);
sram_cell_6t_3 inst_cell_32_62 ( BL62, BLN62, WL32);
sram_cell_6t_3 inst_cell_31_62 ( BL62, BLN62, WL31);
sram_cell_6t_3 inst_cell_32_61 ( BL61, BLN61, WL32);
sram_cell_6t_3 inst_cell_31_61 ( BL61, BLN61, WL31);
sram_cell_6t_3 inst_cell_32_60 ( BL60, BLN60, WL32);
sram_cell_6t_3 inst_cell_31_60 ( BL60, BLN60, WL31);
sram_cell_6t_3 inst_cell_32_59 ( BL59, BLN59, WL32);
sram_cell_6t_3 inst_cell_31_59 ( BL59, BLN59, WL31);
sram_cell_6t_3 inst_cell_32_58 ( BL58, BLN58, WL32);
sram_cell_6t_3 inst_cell_31_58 ( BL58, BLN58, WL31);
sram_cell_6t_3 inst_cell_32_57 ( BL57, BLN57, WL32);
sram_cell_6t_3 inst_cell_31_57 ( BL57, BLN57, WL31);
sram_cell_6t_3 inst_cell_32_56 ( BL56, BLN56, WL32);
sram_cell_6t_3 inst_cell_31_56 ( BL56, BLN56, WL31);
sram_cell_6t_3 inst_cell_32_55 ( BL55, BLN55, WL32);
sram_cell_6t_3 inst_cell_31_55 ( BL55, BLN55, WL31);
sram_cell_6t_3 inst_cell_32_54 ( BL54, BLN54, WL32);
sram_cell_6t_3 inst_cell_31_54 ( BL54, BLN54, WL31);
sram_cell_6t_3 inst_cell_32_53 ( BL53, BLN53, WL32);
sram_cell_6t_3 inst_cell_31_53 ( BL53, BLN53, WL31);
sram_cell_6t_3 inst_cell_32_52 ( BL52, BLN52, WL32);
sram_cell_6t_3 inst_cell_31_52 ( BL52, BLN52, WL31);
sram_cell_6t_3 inst_cell_32_51 ( BL51, BLN51, WL32);
sram_cell_6t_3 inst_cell_31_51 ( BL51, BLN51, WL31);
sram_cell_6t_3 inst_cell_32_50 ( BL50, BLN50, WL32);
sram_cell_6t_3 inst_cell_31_50 ( BL50, BLN50, WL31);
sram_cell_6t_3 inst_cell_32_49 ( BL49, BLN49, WL32);
sram_cell_6t_3 inst_cell_31_49 ( BL49, BLN49, WL31);
sram_cell_6t_3 inst_cell_32_48 ( BL48, BLN48, WL32);
sram_cell_6t_3 inst_cell_31_48 ( BL48, BLN48, WL31);
sram_cell_6t_3 inst_cell_32_47 ( BL47, BLN47, WL32);
sram_cell_6t_3 inst_cell_31_47 ( BL47, BLN47, WL31);
sram_cell_6t_3 inst_cell_32_46 ( BL46, BLN46, WL32);
sram_cell_6t_3 inst_cell_31_46 ( BL46, BLN46, WL31);
sram_cell_6t_3 inst_cell_32_45 ( BL45, BLN45, WL32);
sram_cell_6t_3 inst_cell_31_45 ( BL45, BLN45, WL31);
sram_cell_6t_3 inst_cell_32_44 ( BL44, BLN44, WL32);
sram_cell_6t_3 inst_cell_31_44 ( BL44, BLN44, WL31);
sram_cell_6t_3 inst_cell_32_43 ( BL43, BLN43, WL32);
sram_cell_6t_3 inst_cell_31_43 ( BL43, BLN43, WL31);
sram_cell_6t_3 inst_cell_32_42 ( BL42, BLN42, WL32);
sram_cell_6t_3 inst_cell_31_42 ( BL42, BLN42, WL31);
sram_cell_6t_3 inst_cell_32_41 ( BL41, BLN41, WL32);
sram_cell_6t_3 inst_cell_31_41 ( BL41, BLN41, WL31);
sram_cell_6t_3 inst_cell_32_40 ( BL40, BLN40, WL32);
sram_cell_6t_3 inst_cell_31_40 ( BL40, BLN40, WL31);
sram_cell_6t_3 inst_cell_32_39 ( BL39, BLN39, WL32);
sram_cell_6t_3 inst_cell_31_39 ( BL39, BLN39, WL31);
sram_cell_6t_3 inst_cell_32_38 ( BL38, BLN38, WL32);
sram_cell_6t_3 inst_cell_31_38 ( BL38, BLN38, WL31);
sram_cell_6t_3 inst_cell_32_37 ( BL37, BLN37, WL32);
sram_cell_6t_3 inst_cell_31_37 ( BL37, BLN37, WL31);
sram_cell_6t_3 inst_cell_32_36 ( BL36, BLN36, WL32);
sram_cell_6t_3 inst_cell_31_36 ( BL36, BLN36, WL31);
sram_cell_6t_3 inst_cell_32_35 ( BL35, BLN35, WL32);
sram_cell_6t_3 inst_cell_31_35 ( BL35, BLN35, WL31);
sram_cell_6t_3 inst_cell_32_34 ( BL34, BLN34, WL32);
sram_cell_6t_3 inst_cell_31_34 ( BL34, BLN34, WL31);
sram_cell_6t_3 inst_cell_32_33 ( BL33, BLN33, WL32);
sram_cell_6t_3 inst_cell_31_33 ( BL33, BLN33, WL31);
sram_cell_6t_3 inst_cell_32_32 ( BL32, BLN32, WL32);
sram_cell_6t_3 inst_cell_31_32 ( BL32, BLN32, WL31);
sram_cell_6t_3 inst_cell_32_31 ( BL31, BLN31, WL32);
sram_cell_6t_3 inst_cell_31_31 ( BL31, BLN31, WL31);
sram_cell_6t_3 inst_cell_32_30 ( BL30, BLN30, WL32);
sram_cell_6t_3 inst_cell_31_30 ( BL30, BLN30, WL31);
sram_cell_6t_3 inst_cell_32_29 ( BL29, BLN29, WL32);
sram_cell_6t_3 inst_cell_31_29 ( BL29, BLN29, WL31);
sram_cell_6t_3 inst_cell_32_28 ( BL28, BLN28, WL32);
sram_cell_6t_3 inst_cell_31_28 ( BL28, BLN28, WL31);
sram_cell_6t_3 inst_cell_32_27 ( BL27, BLN27, WL32);
sram_cell_6t_3 inst_cell_31_27 ( BL27, BLN27, WL31);
sram_cell_6t_3 inst_cell_32_26 ( BL26, BLN26, WL32);
sram_cell_6t_3 inst_cell_31_26 ( BL26, BLN26, WL31);
sram_cell_6t_3 inst_cell_32_25 ( BL25, BLN25, WL32);
sram_cell_6t_3 inst_cell_31_25 ( BL25, BLN25, WL31);
sram_cell_6t_3 inst_cell_32_24 ( BL24, BLN24, WL32);
sram_cell_6t_3 inst_cell_31_24 ( BL24, BLN24, WL31);
sram_cell_6t_3 inst_cell_32_23 ( BL23, BLN23, WL32);
sram_cell_6t_3 inst_cell_31_23 ( BL23, BLN23, WL31);
sram_cell_6t_3 inst_cell_32_22 ( BL22, BLN22, WL32);
sram_cell_6t_3 inst_cell_31_22 ( BL22, BLN22, WL31);
sram_cell_6t_3 inst_cell_32_21 ( BL21, BLN21, WL32);
sram_cell_6t_3 inst_cell_31_21 ( BL21, BLN21, WL31);
sram_cell_6t_3 inst_cell_32_20 ( BL20, BLN20, WL32);
sram_cell_6t_3 inst_cell_31_20 ( BL20, BLN20, WL31);
sram_cell_6t_3 inst_cell_32_19 ( BL19, BLN19, WL32);
sram_cell_6t_3 inst_cell_31_19 ( BL19, BLN19, WL31);
sram_cell_6t_3 inst_cell_32_18 ( BL18, BLN18, WL32);
sram_cell_6t_3 inst_cell_31_18 ( BL18, BLN18, WL31);
sram_cell_6t_3 inst_cell_32_17 ( BL17, BLN17, WL32);
sram_cell_6t_3 inst_cell_31_17 ( BL17, BLN17, WL31);
sram_cell_6t_3 inst_cell_32_16 ( BL16, BLN16, WL32);
sram_cell_6t_3 inst_cell_31_16 ( BL16, BLN16, WL31);
sram_cell_6t_3 inst_cell_32_15 ( BL15, BLN15, WL32);
sram_cell_6t_3 inst_cell_31_15 ( BL15, BLN15, WL31);
sram_cell_6t_3 inst_cell_32_14 ( BL14, BLN14, WL32);
sram_cell_6t_3 inst_cell_31_14 ( BL14, BLN14, WL31);
sram_cell_6t_3 inst_cell_32_13 ( BL13, BLN13, WL32);
sram_cell_6t_3 inst_cell_31_13 ( BL13, BLN13, WL31);
sram_cell_6t_3 inst_cell_32_12 ( BL12, BLN12, WL32);
sram_cell_6t_3 inst_cell_31_12 ( BL12, BLN12, WL31);
sram_cell_6t_3 inst_cell_32_11 ( BL11, BLN11, WL32);
sram_cell_6t_3 inst_cell_31_11 ( BL11, BLN11, WL31);
sram_cell_6t_3 inst_cell_32_10 ( BL10, BLN10, WL32);
sram_cell_6t_3 inst_cell_31_10 ( BL10, BLN10, WL31);
sram_cell_6t_3 inst_cell_32_9 ( BL9, BLN9, WL32);
sram_cell_6t_3 inst_cell_31_9 ( BL9, BLN9, WL31);
sram_cell_6t_3 inst_cell_32_8 ( BL8, BLN8, WL32);
sram_cell_6t_3 inst_cell_31_8 ( BL8, BLN8, WL31);
sram_cell_6t_3 inst_cell_33_7 ( BL7, BLN7, WL33);
sram_cell_6t_3 inst_cell_33_6 ( BL6, BLN6, WL33);
sram_cell_6t_3 inst_cell_33_5 ( BL5, BLN5, WL33);
sram_cell_6t_3 inst_cell_33_4 ( BL4, BLN4, WL33);
sram_cell_6t_3 inst_cell_33_3 ( BL3, BLN3, WL33);
sram_cell_6t_3 inst_cell_33_2 ( BL2, BLN2, WL33);
sram_cell_6t_3 inst_cell_33_1 ( BL1, BLN1, WL33);
sram_cell_6t_3 inst_cell_33_0 ( BL0, BLN0, WL33);
sram_cell_6t_3 inst_cell_32_63 ( BL63, BLN63, WL32);
sram_cell_6t_3 inst_cell_32_7 ( BL7, BLN7, WL32);
sram_cell_6t_3 inst_cell_32_6 ( BL6, BLN6, WL32);
sram_cell_6t_3 inst_cell_32_5 ( BL5, BLN5, WL32);
sram_cell_6t_3 inst_cell_32_4 ( BL4, BLN4, WL32);
sram_cell_6t_3 inst_cell_32_3 ( BL3, BLN3, WL32);
sram_cell_6t_3 inst_cell_32_2 ( BL2, BLN2, WL32);
sram_cell_6t_3 inst_cell_32_1 ( BL1, BLN1, WL32);
sram_cell_6t_3 inst_cell_32_0 ( BL0, BLN0, WL32);
sram_cell_6t_3 inst_cell_31_63 ( BL63, BLN63, WL31);
sram_cell_6t_3 inst_cell_31_7 ( BL7, BLN7, WL31);
sram_cell_6t_3 inst_cell_31_6 ( BL6, BLN6, WL31);
sram_cell_6t_3 inst_cell_31_5 ( BL5, BLN5, WL31);
sram_cell_6t_3 inst_cell_31_4 ( BL4, BLN4, WL31);
sram_cell_6t_3 inst_cell_31_3 ( BL3, BLN3, WL31);
sram_cell_6t_3 inst_cell_31_2 ( BL2, BLN2, WL31);
sram_cell_6t_3 inst_cell_31_1 ( BL1, BLN1, WL31);
sram_cell_6t_3 inst_cell_31_0 ( BL0, BLN0, WL31);
sram_cell_6t_3 inst_cell_30_63 ( BL63, BLN63, WL30);
sram_cell_6t_3 inst_cell_30_31 ( BL31, BLN31, WL30);
sram_cell_6t_3 inst_cell_29_31 ( BL31, BLN31, WL29);
sram_cell_6t_3 inst_cell_30_30 ( BL30, BLN30, WL30);
sram_cell_6t_3 inst_cell_29_30 ( BL30, BLN30, WL29);
sram_cell_6t_3 inst_cell_30_29 ( BL29, BLN29, WL30);
sram_cell_6t_3 inst_cell_29_29 ( BL29, BLN29, WL29);
sram_cell_6t_3 inst_cell_30_28 ( BL28, BLN28, WL30);
sram_cell_6t_3 inst_cell_29_28 ( BL28, BLN28, WL29);
sram_cell_6t_3 inst_cell_30_27 ( BL27, BLN27, WL30);
sram_cell_6t_3 inst_cell_29_27 ( BL27, BLN27, WL29);
sram_cell_6t_3 inst_cell_30_26 ( BL26, BLN26, WL30);
sram_cell_6t_3 inst_cell_29_26 ( BL26, BLN26, WL29);
sram_cell_6t_3 inst_cell_30_25 ( BL25, BLN25, WL30);
sram_cell_6t_3 inst_cell_29_25 ( BL25, BLN25, WL29);
sram_cell_6t_3 inst_cell_30_24 ( BL24, BLN24, WL30);
sram_cell_6t_3 inst_cell_29_24 ( BL24, BLN24, WL29);
sram_cell_6t_3 inst_cell_30_23 ( BL23, BLN23, WL30);
sram_cell_6t_3 inst_cell_29_23 ( BL23, BLN23, WL29);
sram_cell_6t_3 inst_cell_30_22 ( BL22, BLN22, WL30);
sram_cell_6t_3 inst_cell_29_22 ( BL22, BLN22, WL29);
sram_cell_6t_3 inst_cell_30_21 ( BL21, BLN21, WL30);
sram_cell_6t_3 inst_cell_29_21 ( BL21, BLN21, WL29);
sram_cell_6t_3 inst_cell_30_20 ( BL20, BLN20, WL30);
sram_cell_6t_3 inst_cell_29_20 ( BL20, BLN20, WL29);
sram_cell_6t_3 inst_cell_30_19 ( BL19, BLN19, WL30);
sram_cell_6t_3 inst_cell_29_19 ( BL19, BLN19, WL29);
sram_cell_6t_3 inst_cell_30_18 ( BL18, BLN18, WL30);
sram_cell_6t_3 inst_cell_29_18 ( BL18, BLN18, WL29);
sram_cell_6t_3 inst_cell_30_17 ( BL17, BLN17, WL30);
sram_cell_6t_3 inst_cell_29_17 ( BL17, BLN17, WL29);
sram_cell_6t_3 inst_cell_30_16 ( BL16, BLN16, WL30);
sram_cell_6t_3 inst_cell_29_16 ( BL16, BLN16, WL29);
sram_cell_6t_3 inst_cell_30_15 ( BL15, BLN15, WL30);
sram_cell_6t_3 inst_cell_29_15 ( BL15, BLN15, WL29);
sram_cell_6t_3 inst_cell_30_14 ( BL14, BLN14, WL30);
sram_cell_6t_3 inst_cell_29_14 ( BL14, BLN14, WL29);
sram_cell_6t_3 inst_cell_30_13 ( BL13, BLN13, WL30);
sram_cell_6t_3 inst_cell_29_13 ( BL13, BLN13, WL29);
sram_cell_6t_3 inst_cell_30_12 ( BL12, BLN12, WL30);
sram_cell_6t_3 inst_cell_29_12 ( BL12, BLN12, WL29);
sram_cell_6t_3 inst_cell_30_11 ( BL11, BLN11, WL30);
sram_cell_6t_3 inst_cell_29_11 ( BL11, BLN11, WL29);
sram_cell_6t_3 inst_cell_30_10 ( BL10, BLN10, WL30);
sram_cell_6t_3 inst_cell_29_10 ( BL10, BLN10, WL29);
sram_cell_6t_3 inst_cell_30_9 ( BL9, BLN9, WL30);
sram_cell_6t_3 inst_cell_29_9 ( BL9, BLN9, WL29);
sram_cell_6t_3 inst_cell_30_8 ( BL8, BLN8, WL30);
sram_cell_6t_3 inst_cell_29_8 ( BL8, BLN8, WL29);
sram_cell_6t_3 inst_cell_30_7 ( BL7, BLN7, WL30);
sram_cell_6t_3 inst_cell_29_7 ( BL7, BLN7, WL29);
sram_cell_6t_3 inst_cell_30_6 ( BL6, BLN6, WL30);
sram_cell_6t_3 inst_cell_29_6 ( BL6, BLN6, WL29);
sram_cell_6t_3 inst_cell_30_5 ( BL5, BLN5, WL30);
sram_cell_6t_3 inst_cell_29_5 ( BL5, BLN5, WL29);
sram_cell_6t_3 inst_cell_30_4 ( BL4, BLN4, WL30);
sram_cell_6t_3 inst_cell_29_4 ( BL4, BLN4, WL29);
sram_cell_6t_3 inst_cell_30_3 ( BL3, BLN3, WL30);
sram_cell_6t_3 inst_cell_29_3 ( BL3, BLN3, WL29);
sram_cell_6t_3 inst_cell_30_2 ( BL2, BLN2, WL30);
sram_cell_6t_3 inst_cell_29_2 ( BL2, BLN2, WL29);
sram_cell_6t_3 inst_cell_30_1 ( BL1, BLN1, WL30);
sram_cell_6t_3 inst_cell_29_1 ( BL1, BLN1, WL29);
sram_cell_6t_3 inst_cell_30_0 ( BL0, BLN0, WL30);
sram_cell_6t_3 inst_cell_29_0 ( BL0, BLN0, WL29);
sram_cell_6t_3 inst_cell_29_63 ( BL63, BLN63, WL29);
sram_cell_6t_3 inst_cell_28_63 ( BL63, BLN63, WL28);
sram_cell_6t_3 inst_cell_30_62 ( BL62, BLN62, WL30);
sram_cell_6t_3 inst_cell_30_61 ( BL61, BLN61, WL30);
sram_cell_6t_3 inst_cell_30_60 ( BL60, BLN60, WL30);
sram_cell_6t_3 inst_cell_30_59 ( BL59, BLN59, WL30);
sram_cell_6t_3 inst_cell_30_58 ( BL58, BLN58, WL30);
sram_cell_6t_3 inst_cell_30_57 ( BL57, BLN57, WL30);
sram_cell_6t_3 inst_cell_30_56 ( BL56, BLN56, WL30);
sram_cell_6t_3 inst_cell_30_55 ( BL55, BLN55, WL30);
sram_cell_6t_3 inst_cell_30_54 ( BL54, BLN54, WL30);
sram_cell_6t_3 inst_cell_30_53 ( BL53, BLN53, WL30);
sram_cell_6t_3 inst_cell_30_52 ( BL52, BLN52, WL30);
sram_cell_6t_3 inst_cell_30_51 ( BL51, BLN51, WL30);
sram_cell_6t_3 inst_cell_30_50 ( BL50, BLN50, WL30);
sram_cell_6t_3 inst_cell_30_49 ( BL49, BLN49, WL30);
sram_cell_6t_3 inst_cell_30_48 ( BL48, BLN48, WL30);
sram_cell_6t_3 inst_cell_30_47 ( BL47, BLN47, WL30);
sram_cell_6t_3 inst_cell_30_46 ( BL46, BLN46, WL30);
sram_cell_6t_3 inst_cell_30_45 ( BL45, BLN45, WL30);
sram_cell_6t_3 inst_cell_30_44 ( BL44, BLN44, WL30);
sram_cell_6t_3 inst_cell_30_43 ( BL43, BLN43, WL30);
sram_cell_6t_3 inst_cell_30_42 ( BL42, BLN42, WL30);
sram_cell_6t_3 inst_cell_30_41 ( BL41, BLN41, WL30);
sram_cell_6t_3 inst_cell_30_40 ( BL40, BLN40, WL30);
sram_cell_6t_3 inst_cell_30_39 ( BL39, BLN39, WL30);
sram_cell_6t_3 inst_cell_30_38 ( BL38, BLN38, WL30);
sram_cell_6t_3 inst_cell_30_37 ( BL37, BLN37, WL30);
sram_cell_6t_3 inst_cell_30_36 ( BL36, BLN36, WL30);
sram_cell_6t_3 inst_cell_30_35 ( BL35, BLN35, WL30);
sram_cell_6t_3 inst_cell_30_34 ( BL34, BLN34, WL30);
sram_cell_6t_3 inst_cell_30_33 ( BL33, BLN33, WL30);
sram_cell_6t_3 inst_cell_30_32 ( BL32, BLN32, WL30);
sram_cell_6t_3 inst_cell_29_62 ( BL62, BLN62, WL29);
sram_cell_6t_3 inst_cell_29_61 ( BL61, BLN61, WL29);
sram_cell_6t_3 inst_cell_29_60 ( BL60, BLN60, WL29);
sram_cell_6t_3 inst_cell_29_59 ( BL59, BLN59, WL29);
sram_cell_6t_3 inst_cell_29_58 ( BL58, BLN58, WL29);
sram_cell_6t_3 inst_cell_29_57 ( BL57, BLN57, WL29);
sram_cell_6t_3 inst_cell_29_56 ( BL56, BLN56, WL29);
sram_cell_6t_3 inst_cell_29_55 ( BL55, BLN55, WL29);
sram_cell_6t_3 inst_cell_29_54 ( BL54, BLN54, WL29);
sram_cell_6t_3 inst_cell_29_53 ( BL53, BLN53, WL29);
sram_cell_6t_3 inst_cell_29_52 ( BL52, BLN52, WL29);
sram_cell_6t_3 inst_cell_29_51 ( BL51, BLN51, WL29);
sram_cell_6t_3 inst_cell_29_50 ( BL50, BLN50, WL29);
sram_cell_6t_3 inst_cell_29_49 ( BL49, BLN49, WL29);
sram_cell_6t_3 inst_cell_29_48 ( BL48, BLN48, WL29);
sram_cell_6t_3 inst_cell_29_47 ( BL47, BLN47, WL29);
sram_cell_6t_3 inst_cell_29_46 ( BL46, BLN46, WL29);
sram_cell_6t_3 inst_cell_29_45 ( BL45, BLN45, WL29);
sram_cell_6t_3 inst_cell_29_44 ( BL44, BLN44, WL29);
sram_cell_6t_3 inst_cell_29_43 ( BL43, BLN43, WL29);
sram_cell_6t_3 inst_cell_29_42 ( BL42, BLN42, WL29);
sram_cell_6t_3 inst_cell_29_41 ( BL41, BLN41, WL29);
sram_cell_6t_3 inst_cell_29_40 ( BL40, BLN40, WL29);
sram_cell_6t_3 inst_cell_29_39 ( BL39, BLN39, WL29);
sram_cell_6t_3 inst_cell_29_38 ( BL38, BLN38, WL29);
sram_cell_6t_3 inst_cell_29_37 ( BL37, BLN37, WL29);
sram_cell_6t_3 inst_cell_29_36 ( BL36, BLN36, WL29);
sram_cell_6t_3 inst_cell_29_35 ( BL35, BLN35, WL29);
sram_cell_6t_3 inst_cell_29_34 ( BL34, BLN34, WL29);
sram_cell_6t_3 inst_cell_29_33 ( BL33, BLN33, WL29);
sram_cell_6t_3 inst_cell_29_32 ( BL32, BLN32, WL29);
sram_cell_6t_3 inst_cell_28_62 ( BL62, BLN62, WL28);
sram_cell_6t_3 inst_cell_28_61 ( BL61, BLN61, WL28);
sram_cell_6t_3 inst_cell_28_60 ( BL60, BLN60, WL28);
sram_cell_6t_3 inst_cell_28_59 ( BL59, BLN59, WL28);
sram_cell_6t_3 inst_cell_28_58 ( BL58, BLN58, WL28);
sram_cell_6t_3 inst_cell_28_57 ( BL57, BLN57, WL28);
sram_cell_6t_3 inst_cell_28_56 ( BL56, BLN56, WL28);
sram_cell_6t_3 inst_cell_28_55 ( BL55, BLN55, WL28);
sram_cell_6t_3 inst_cell_28_54 ( BL54, BLN54, WL28);
sram_cell_6t_3 inst_cell_28_53 ( BL53, BLN53, WL28);
sram_cell_6t_3 inst_cell_28_52 ( BL52, BLN52, WL28);
sram_cell_6t_3 inst_cell_28_51 ( BL51, BLN51, WL28);
sram_cell_6t_3 inst_cell_28_50 ( BL50, BLN50, WL28);
sram_cell_6t_3 inst_cell_28_49 ( BL49, BLN49, WL28);
sram_cell_6t_3 inst_cell_28_48 ( BL48, BLN48, WL28);
sram_cell_6t_3 inst_cell_28_47 ( BL47, BLN47, WL28);
sram_cell_6t_3 inst_cell_28_46 ( BL46, BLN46, WL28);
sram_cell_6t_3 inst_cell_28_45 ( BL45, BLN45, WL28);
sram_cell_6t_3 inst_cell_28_44 ( BL44, BLN44, WL28);
sram_cell_6t_3 inst_cell_28_43 ( BL43, BLN43, WL28);
sram_cell_6t_3 inst_cell_28_42 ( BL42, BLN42, WL28);
sram_cell_6t_3 inst_cell_28_41 ( BL41, BLN41, WL28);
sram_cell_6t_3 inst_cell_28_40 ( BL40, BLN40, WL28);
sram_cell_6t_3 inst_cell_28_39 ( BL39, BLN39, WL28);
sram_cell_6t_3 inst_cell_28_38 ( BL38, BLN38, WL28);
sram_cell_6t_3 inst_cell_28_37 ( BL37, BLN37, WL28);
sram_cell_6t_3 inst_cell_28_36 ( BL36, BLN36, WL28);
sram_cell_6t_3 inst_cell_28_35 ( BL35, BLN35, WL28);
sram_cell_6t_3 inst_cell_28_34 ( BL34, BLN34, WL28);
sram_cell_6t_3 inst_cell_28_33 ( BL33, BLN33, WL28);
sram_cell_6t_3 inst_cell_28_32 ( BL32, BLN32, WL28);
sram_cell_6t_3 inst_cell_28_7 ( BL7, BLN7, WL28);
sram_cell_6t_3 inst_cell_27_7 ( BL7, BLN7, WL27);
sram_cell_6t_3 inst_cell_28_6 ( BL6, BLN6, WL28);
sram_cell_6t_3 inst_cell_27_6 ( BL6, BLN6, WL27);
sram_cell_6t_3 inst_cell_28_5 ( BL5, BLN5, WL28);
sram_cell_6t_3 inst_cell_27_5 ( BL5, BLN5, WL27);
sram_cell_6t_3 inst_cell_28_4 ( BL4, BLN4, WL28);
sram_cell_6t_3 inst_cell_27_4 ( BL4, BLN4, WL27);
sram_cell_6t_3 inst_cell_28_3 ( BL3, BLN3, WL28);
sram_cell_6t_3 inst_cell_27_3 ( BL3, BLN3, WL27);
sram_cell_6t_3 inst_cell_28_2 ( BL2, BLN2, WL28);
sram_cell_6t_3 inst_cell_27_2 ( BL2, BLN2, WL27);
sram_cell_6t_3 inst_cell_28_1 ( BL1, BLN1, WL28);
sram_cell_6t_3 inst_cell_27_1 ( BL1, BLN1, WL27);
sram_cell_6t_3 inst_cell_28_0 ( BL0, BLN0, WL28);
sram_cell_6t_3 inst_cell_27_0 ( BL0, BLN0, WL27);
sram_cell_6t_3 inst_cell_27_63 ( BL63, BLN63, WL27);
sram_cell_6t_3 inst_cell_26_63 ( BL63, BLN63, WL26);
sram_cell_6t_3 inst_cell_27_62 ( BL62, BLN62, WL27);
sram_cell_6t_3 inst_cell_26_62 ( BL62, BLN62, WL26);
sram_cell_6t_3 inst_cell_27_61 ( BL61, BLN61, WL27);
sram_cell_6t_3 inst_cell_26_61 ( BL61, BLN61, WL26);
sram_cell_6t_3 inst_cell_27_60 ( BL60, BLN60, WL27);
sram_cell_6t_3 inst_cell_26_60 ( BL60, BLN60, WL26);
sram_cell_6t_3 inst_cell_27_59 ( BL59, BLN59, WL27);
sram_cell_6t_3 inst_cell_26_59 ( BL59, BLN59, WL26);
sram_cell_6t_3 inst_cell_27_58 ( BL58, BLN58, WL27);
sram_cell_6t_3 inst_cell_26_58 ( BL58, BLN58, WL26);
sram_cell_6t_3 inst_cell_27_57 ( BL57, BLN57, WL27);
sram_cell_6t_3 inst_cell_26_57 ( BL57, BLN57, WL26);
sram_cell_6t_3 inst_cell_27_56 ( BL56, BLN56, WL27);
sram_cell_6t_3 inst_cell_26_56 ( BL56, BLN56, WL26);
sram_cell_6t_3 inst_cell_27_55 ( BL55, BLN55, WL27);
sram_cell_6t_3 inst_cell_26_55 ( BL55, BLN55, WL26);
sram_cell_6t_3 inst_cell_27_54 ( BL54, BLN54, WL27);
sram_cell_6t_3 inst_cell_26_54 ( BL54, BLN54, WL26);
sram_cell_6t_3 inst_cell_27_53 ( BL53, BLN53, WL27);
sram_cell_6t_3 inst_cell_26_53 ( BL53, BLN53, WL26);
sram_cell_6t_3 inst_cell_27_52 ( BL52, BLN52, WL27);
sram_cell_6t_3 inst_cell_26_52 ( BL52, BLN52, WL26);
sram_cell_6t_3 inst_cell_27_51 ( BL51, BLN51, WL27);
sram_cell_6t_3 inst_cell_26_51 ( BL51, BLN51, WL26);
sram_cell_6t_3 inst_cell_27_50 ( BL50, BLN50, WL27);
sram_cell_6t_3 inst_cell_26_50 ( BL50, BLN50, WL26);
sram_cell_6t_3 inst_cell_27_49 ( BL49, BLN49, WL27);
sram_cell_6t_3 inst_cell_26_49 ( BL49, BLN49, WL26);
sram_cell_6t_3 inst_cell_27_48 ( BL48, BLN48, WL27);
sram_cell_6t_3 inst_cell_26_48 ( BL48, BLN48, WL26);
sram_cell_6t_3 inst_cell_27_47 ( BL47, BLN47, WL27);
sram_cell_6t_3 inst_cell_26_47 ( BL47, BLN47, WL26);
sram_cell_6t_3 inst_cell_27_46 ( BL46, BLN46, WL27);
sram_cell_6t_3 inst_cell_26_46 ( BL46, BLN46, WL26);
sram_cell_6t_3 inst_cell_27_45 ( BL45, BLN45, WL27);
sram_cell_6t_3 inst_cell_26_45 ( BL45, BLN45, WL26);
sram_cell_6t_3 inst_cell_27_44 ( BL44, BLN44, WL27);
sram_cell_6t_3 inst_cell_26_44 ( BL44, BLN44, WL26);
sram_cell_6t_3 inst_cell_27_43 ( BL43, BLN43, WL27);
sram_cell_6t_3 inst_cell_26_43 ( BL43, BLN43, WL26);
sram_cell_6t_3 inst_cell_27_42 ( BL42, BLN42, WL27);
sram_cell_6t_3 inst_cell_26_42 ( BL42, BLN42, WL26);
sram_cell_6t_3 inst_cell_27_41 ( BL41, BLN41, WL27);
sram_cell_6t_3 inst_cell_26_41 ( BL41, BLN41, WL26);
sram_cell_6t_3 inst_cell_27_40 ( BL40, BLN40, WL27);
sram_cell_6t_3 inst_cell_26_40 ( BL40, BLN40, WL26);
sram_cell_6t_3 inst_cell_27_39 ( BL39, BLN39, WL27);
sram_cell_6t_3 inst_cell_26_39 ( BL39, BLN39, WL26);
sram_cell_6t_3 inst_cell_27_38 ( BL38, BLN38, WL27);
sram_cell_6t_3 inst_cell_26_38 ( BL38, BLN38, WL26);
sram_cell_6t_3 inst_cell_27_37 ( BL37, BLN37, WL27);
sram_cell_6t_3 inst_cell_26_37 ( BL37, BLN37, WL26);
sram_cell_6t_3 inst_cell_27_36 ( BL36, BLN36, WL27);
sram_cell_6t_3 inst_cell_26_36 ( BL36, BLN36, WL26);
sram_cell_6t_3 inst_cell_27_35 ( BL35, BLN35, WL27);
sram_cell_6t_3 inst_cell_26_35 ( BL35, BLN35, WL26);
sram_cell_6t_3 inst_cell_27_34 ( BL34, BLN34, WL27);
sram_cell_6t_3 inst_cell_26_34 ( BL34, BLN34, WL26);
sram_cell_6t_3 inst_cell_27_33 ( BL33, BLN33, WL27);
sram_cell_6t_3 inst_cell_26_33 ( BL33, BLN33, WL26);
sram_cell_6t_3 inst_cell_27_32 ( BL32, BLN32, WL27);
sram_cell_6t_3 inst_cell_26_32 ( BL32, BLN32, WL26);
sram_cell_6t_3 inst_cell_28_31 ( BL31, BLN31, WL28);
sram_cell_6t_3 inst_cell_28_30 ( BL30, BLN30, WL28);
sram_cell_6t_3 inst_cell_28_29 ( BL29, BLN29, WL28);
sram_cell_6t_3 inst_cell_28_28 ( BL28, BLN28, WL28);
sram_cell_6t_3 inst_cell_28_27 ( BL27, BLN27, WL28);
sram_cell_6t_3 inst_cell_28_26 ( BL26, BLN26, WL28);
sram_cell_6t_3 inst_cell_28_25 ( BL25, BLN25, WL28);
sram_cell_6t_3 inst_cell_28_24 ( BL24, BLN24, WL28);
sram_cell_6t_3 inst_cell_28_23 ( BL23, BLN23, WL28);
sram_cell_6t_3 inst_cell_28_22 ( BL22, BLN22, WL28);
sram_cell_6t_3 inst_cell_28_21 ( BL21, BLN21, WL28);
sram_cell_6t_3 inst_cell_28_20 ( BL20, BLN20, WL28);
sram_cell_6t_3 inst_cell_28_19 ( BL19, BLN19, WL28);
sram_cell_6t_3 inst_cell_28_18 ( BL18, BLN18, WL28);
sram_cell_6t_3 inst_cell_28_17 ( BL17, BLN17, WL28);
sram_cell_6t_3 inst_cell_28_16 ( BL16, BLN16, WL28);
sram_cell_6t_3 inst_cell_28_15 ( BL15, BLN15, WL28);
sram_cell_6t_3 inst_cell_28_14 ( BL14, BLN14, WL28);
sram_cell_6t_3 inst_cell_28_13 ( BL13, BLN13, WL28);
sram_cell_6t_3 inst_cell_28_12 ( BL12, BLN12, WL28);
sram_cell_6t_3 inst_cell_28_11 ( BL11, BLN11, WL28);
sram_cell_6t_3 inst_cell_28_10 ( BL10, BLN10, WL28);
sram_cell_6t_3 inst_cell_28_9 ( BL9, BLN9, WL28);
sram_cell_6t_3 inst_cell_28_8 ( BL8, BLN8, WL28);
sram_cell_6t_3 inst_cell_27_31 ( BL31, BLN31, WL27);
sram_cell_6t_3 inst_cell_27_30 ( BL30, BLN30, WL27);
sram_cell_6t_3 inst_cell_27_29 ( BL29, BLN29, WL27);
sram_cell_6t_3 inst_cell_27_28 ( BL28, BLN28, WL27);
sram_cell_6t_3 inst_cell_27_27 ( BL27, BLN27, WL27);
sram_cell_6t_3 inst_cell_27_26 ( BL26, BLN26, WL27);
sram_cell_6t_3 inst_cell_27_25 ( BL25, BLN25, WL27);
sram_cell_6t_3 inst_cell_27_24 ( BL24, BLN24, WL27);
sram_cell_6t_3 inst_cell_27_23 ( BL23, BLN23, WL27);
sram_cell_6t_3 inst_cell_27_22 ( BL22, BLN22, WL27);
sram_cell_6t_3 inst_cell_27_21 ( BL21, BLN21, WL27);
sram_cell_6t_3 inst_cell_27_20 ( BL20, BLN20, WL27);
sram_cell_6t_3 inst_cell_27_19 ( BL19, BLN19, WL27);
sram_cell_6t_3 inst_cell_27_18 ( BL18, BLN18, WL27);
sram_cell_6t_3 inst_cell_27_17 ( BL17, BLN17, WL27);
sram_cell_6t_3 inst_cell_27_16 ( BL16, BLN16, WL27);
sram_cell_6t_3 inst_cell_27_15 ( BL15, BLN15, WL27);
sram_cell_6t_3 inst_cell_27_14 ( BL14, BLN14, WL27);
sram_cell_6t_3 inst_cell_27_13 ( BL13, BLN13, WL27);
sram_cell_6t_3 inst_cell_27_12 ( BL12, BLN12, WL27);
sram_cell_6t_3 inst_cell_27_11 ( BL11, BLN11, WL27);
sram_cell_6t_3 inst_cell_27_10 ( BL10, BLN10, WL27);
sram_cell_6t_3 inst_cell_27_9 ( BL9, BLN9, WL27);
sram_cell_6t_3 inst_cell_27_8 ( BL8, BLN8, WL27);
sram_cell_6t_3 inst_cell_26_31 ( BL31, BLN31, WL26);
sram_cell_6t_3 inst_cell_26_30 ( BL30, BLN30, WL26);
sram_cell_6t_3 inst_cell_26_29 ( BL29, BLN29, WL26);
sram_cell_6t_3 inst_cell_26_28 ( BL28, BLN28, WL26);
sram_cell_6t_3 inst_cell_26_27 ( BL27, BLN27, WL26);
sram_cell_6t_3 inst_cell_26_26 ( BL26, BLN26, WL26);
sram_cell_6t_3 inst_cell_26_25 ( BL25, BLN25, WL26);
sram_cell_6t_3 inst_cell_26_24 ( BL24, BLN24, WL26);
sram_cell_6t_3 inst_cell_26_23 ( BL23, BLN23, WL26);
sram_cell_6t_3 inst_cell_26_22 ( BL22, BLN22, WL26);
sram_cell_6t_3 inst_cell_26_21 ( BL21, BLN21, WL26);
sram_cell_6t_3 inst_cell_26_20 ( BL20, BLN20, WL26);
sram_cell_6t_3 inst_cell_26_19 ( BL19, BLN19, WL26);
sram_cell_6t_3 inst_cell_26_18 ( BL18, BLN18, WL26);
sram_cell_6t_3 inst_cell_26_17 ( BL17, BLN17, WL26);
sram_cell_6t_3 inst_cell_26_16 ( BL16, BLN16, WL26);
sram_cell_6t_3 inst_cell_26_15 ( BL15, BLN15, WL26);
sram_cell_6t_3 inst_cell_26_14 ( BL14, BLN14, WL26);
sram_cell_6t_3 inst_cell_26_13 ( BL13, BLN13, WL26);
sram_cell_6t_3 inst_cell_26_12 ( BL12, BLN12, WL26);
sram_cell_6t_3 inst_cell_26_11 ( BL11, BLN11, WL26);
sram_cell_6t_3 inst_cell_26_10 ( BL10, BLN10, WL26);
sram_cell_6t_3 inst_cell_26_9 ( BL9, BLN9, WL26);
sram_cell_6t_3 inst_cell_26_8 ( BL8, BLN8, WL26);
sram_cell_6t_3 inst_cell_25_62 ( BL62, BLN62, WL25);
sram_cell_6t_3 inst_cell_24_62 ( BL62, BLN62, WL24);
sram_cell_6t_3 inst_cell_25_61 ( BL61, BLN61, WL25);
sram_cell_6t_3 inst_cell_24_61 ( BL61, BLN61, WL24);
sram_cell_6t_3 inst_cell_25_60 ( BL60, BLN60, WL25);
sram_cell_6t_3 inst_cell_24_60 ( BL60, BLN60, WL24);
sram_cell_6t_3 inst_cell_25_59 ( BL59, BLN59, WL25);
sram_cell_6t_3 inst_cell_24_59 ( BL59, BLN59, WL24);
sram_cell_6t_3 inst_cell_25_58 ( BL58, BLN58, WL25);
sram_cell_6t_3 inst_cell_24_58 ( BL58, BLN58, WL24);
sram_cell_6t_3 inst_cell_25_57 ( BL57, BLN57, WL25);
sram_cell_6t_3 inst_cell_24_57 ( BL57, BLN57, WL24);
sram_cell_6t_3 inst_cell_25_56 ( BL56, BLN56, WL25);
sram_cell_6t_3 inst_cell_24_56 ( BL56, BLN56, WL24);
sram_cell_6t_3 inst_cell_25_55 ( BL55, BLN55, WL25);
sram_cell_6t_3 inst_cell_24_55 ( BL55, BLN55, WL24);
sram_cell_6t_3 inst_cell_25_54 ( BL54, BLN54, WL25);
sram_cell_6t_3 inst_cell_24_54 ( BL54, BLN54, WL24);
sram_cell_6t_3 inst_cell_25_53 ( BL53, BLN53, WL25);
sram_cell_6t_3 inst_cell_24_53 ( BL53, BLN53, WL24);
sram_cell_6t_3 inst_cell_25_52 ( BL52, BLN52, WL25);
sram_cell_6t_3 inst_cell_24_52 ( BL52, BLN52, WL24);
sram_cell_6t_3 inst_cell_25_51 ( BL51, BLN51, WL25);
sram_cell_6t_3 inst_cell_24_51 ( BL51, BLN51, WL24);
sram_cell_6t_3 inst_cell_25_50 ( BL50, BLN50, WL25);
sram_cell_6t_3 inst_cell_24_50 ( BL50, BLN50, WL24);
sram_cell_6t_3 inst_cell_25_49 ( BL49, BLN49, WL25);
sram_cell_6t_3 inst_cell_24_49 ( BL49, BLN49, WL24);
sram_cell_6t_3 inst_cell_25_48 ( BL48, BLN48, WL25);
sram_cell_6t_3 inst_cell_24_48 ( BL48, BLN48, WL24);
sram_cell_6t_3 inst_cell_25_47 ( BL47, BLN47, WL25);
sram_cell_6t_3 inst_cell_24_47 ( BL47, BLN47, WL24);
sram_cell_6t_3 inst_cell_25_46 ( BL46, BLN46, WL25);
sram_cell_6t_3 inst_cell_24_46 ( BL46, BLN46, WL24);
sram_cell_6t_3 inst_cell_25_45 ( BL45, BLN45, WL25);
sram_cell_6t_3 inst_cell_24_45 ( BL45, BLN45, WL24);
sram_cell_6t_3 inst_cell_25_44 ( BL44, BLN44, WL25);
sram_cell_6t_3 inst_cell_24_44 ( BL44, BLN44, WL24);
sram_cell_6t_3 inst_cell_25_43 ( BL43, BLN43, WL25);
sram_cell_6t_3 inst_cell_24_43 ( BL43, BLN43, WL24);
sram_cell_6t_3 inst_cell_25_42 ( BL42, BLN42, WL25);
sram_cell_6t_3 inst_cell_24_42 ( BL42, BLN42, WL24);
sram_cell_6t_3 inst_cell_25_41 ( BL41, BLN41, WL25);
sram_cell_6t_3 inst_cell_24_41 ( BL41, BLN41, WL24);
sram_cell_6t_3 inst_cell_25_40 ( BL40, BLN40, WL25);
sram_cell_6t_3 inst_cell_24_40 ( BL40, BLN40, WL24);
sram_cell_6t_3 inst_cell_25_39 ( BL39, BLN39, WL25);
sram_cell_6t_3 inst_cell_24_39 ( BL39, BLN39, WL24);
sram_cell_6t_3 inst_cell_25_38 ( BL38, BLN38, WL25);
sram_cell_6t_3 inst_cell_24_38 ( BL38, BLN38, WL24);
sram_cell_6t_3 inst_cell_25_37 ( BL37, BLN37, WL25);
sram_cell_6t_3 inst_cell_24_37 ( BL37, BLN37, WL24);
sram_cell_6t_3 inst_cell_25_36 ( BL36, BLN36, WL25);
sram_cell_6t_3 inst_cell_24_36 ( BL36, BLN36, WL24);
sram_cell_6t_3 inst_cell_25_35 ( BL35, BLN35, WL25);
sram_cell_6t_3 inst_cell_24_35 ( BL35, BLN35, WL24);
sram_cell_6t_3 inst_cell_25_34 ( BL34, BLN34, WL25);
sram_cell_6t_3 inst_cell_24_34 ( BL34, BLN34, WL24);
sram_cell_6t_3 inst_cell_25_33 ( BL33, BLN33, WL25);
sram_cell_6t_3 inst_cell_24_33 ( BL33, BLN33, WL24);
sram_cell_6t_3 inst_cell_25_32 ( BL32, BLN32, WL25);
sram_cell_6t_3 inst_cell_24_32 ( BL32, BLN32, WL24);
sram_cell_6t_3 inst_cell_25_31 ( BL31, BLN31, WL25);
sram_cell_6t_3 inst_cell_24_31 ( BL31, BLN31, WL24);
sram_cell_6t_3 inst_cell_25_30 ( BL30, BLN30, WL25);
sram_cell_6t_3 inst_cell_24_30 ( BL30, BLN30, WL24);
sram_cell_6t_3 inst_cell_25_29 ( BL29, BLN29, WL25);
sram_cell_6t_3 inst_cell_24_29 ( BL29, BLN29, WL24);
sram_cell_6t_3 inst_cell_25_28 ( BL28, BLN28, WL25);
sram_cell_6t_3 inst_cell_24_28 ( BL28, BLN28, WL24);
sram_cell_6t_3 inst_cell_25_27 ( BL27, BLN27, WL25);
sram_cell_6t_3 inst_cell_24_27 ( BL27, BLN27, WL24);
sram_cell_6t_3 inst_cell_25_26 ( BL26, BLN26, WL25);
sram_cell_6t_3 inst_cell_24_26 ( BL26, BLN26, WL24);
sram_cell_6t_3 inst_cell_25_25 ( BL25, BLN25, WL25);
sram_cell_6t_3 inst_cell_24_25 ( BL25, BLN25, WL24);
sram_cell_6t_3 inst_cell_25_24 ( BL24, BLN24, WL25);
sram_cell_6t_3 inst_cell_24_24 ( BL24, BLN24, WL24);
sram_cell_6t_3 inst_cell_25_23 ( BL23, BLN23, WL25);
sram_cell_6t_3 inst_cell_24_23 ( BL23, BLN23, WL24);
sram_cell_6t_3 inst_cell_25_22 ( BL22, BLN22, WL25);
sram_cell_6t_3 inst_cell_24_22 ( BL22, BLN22, WL24);
sram_cell_6t_3 inst_cell_25_21 ( BL21, BLN21, WL25);
sram_cell_6t_3 inst_cell_24_21 ( BL21, BLN21, WL24);
sram_cell_6t_3 inst_cell_25_20 ( BL20, BLN20, WL25);
sram_cell_6t_3 inst_cell_24_20 ( BL20, BLN20, WL24);
sram_cell_6t_3 inst_cell_25_19 ( BL19, BLN19, WL25);
sram_cell_6t_3 inst_cell_24_19 ( BL19, BLN19, WL24);
sram_cell_6t_3 inst_cell_25_18 ( BL18, BLN18, WL25);
sram_cell_6t_3 inst_cell_24_18 ( BL18, BLN18, WL24);
sram_cell_6t_3 inst_cell_25_17 ( BL17, BLN17, WL25);
sram_cell_6t_3 inst_cell_24_17 ( BL17, BLN17, WL24);
sram_cell_6t_3 inst_cell_25_16 ( BL16, BLN16, WL25);
sram_cell_6t_3 inst_cell_24_16 ( BL16, BLN16, WL24);
sram_cell_6t_3 inst_cell_25_15 ( BL15, BLN15, WL25);
sram_cell_6t_3 inst_cell_24_15 ( BL15, BLN15, WL24);
sram_cell_6t_3 inst_cell_25_14 ( BL14, BLN14, WL25);
sram_cell_6t_3 inst_cell_24_14 ( BL14, BLN14, WL24);
sram_cell_6t_3 inst_cell_25_13 ( BL13, BLN13, WL25);
sram_cell_6t_3 inst_cell_24_13 ( BL13, BLN13, WL24);
sram_cell_6t_3 inst_cell_25_12 ( BL12, BLN12, WL25);
sram_cell_6t_3 inst_cell_24_12 ( BL12, BLN12, WL24);
sram_cell_6t_3 inst_cell_25_11 ( BL11, BLN11, WL25);
sram_cell_6t_3 inst_cell_24_11 ( BL11, BLN11, WL24);
sram_cell_6t_3 inst_cell_25_10 ( BL10, BLN10, WL25);
sram_cell_6t_3 inst_cell_24_10 ( BL10, BLN10, WL24);
sram_cell_6t_3 inst_cell_25_9 ( BL9, BLN9, WL25);
sram_cell_6t_3 inst_cell_24_9 ( BL9, BLN9, WL24);
sram_cell_6t_3 inst_cell_25_8 ( BL8, BLN8, WL25);
sram_cell_6t_3 inst_cell_24_8 ( BL8, BLN8, WL24);
sram_cell_6t_3 inst_cell_26_7 ( BL7, BLN7, WL26);
sram_cell_6t_3 inst_cell_26_6 ( BL6, BLN6, WL26);
sram_cell_6t_3 inst_cell_26_5 ( BL5, BLN5, WL26);
sram_cell_6t_3 inst_cell_26_4 ( BL4, BLN4, WL26);
sram_cell_6t_3 inst_cell_26_3 ( BL3, BLN3, WL26);
sram_cell_6t_3 inst_cell_26_2 ( BL2, BLN2, WL26);
sram_cell_6t_3 inst_cell_26_1 ( BL1, BLN1, WL26);
sram_cell_6t_3 inst_cell_26_0 ( BL0, BLN0, WL26);
sram_cell_6t_3 inst_cell_25_63 ( BL63, BLN63, WL25);
sram_cell_6t_3 inst_cell_25_7 ( BL7, BLN7, WL25);
sram_cell_6t_3 inst_cell_25_6 ( BL6, BLN6, WL25);
sram_cell_6t_3 inst_cell_25_5 ( BL5, BLN5, WL25);
sram_cell_6t_3 inst_cell_25_4 ( BL4, BLN4, WL25);
sram_cell_6t_3 inst_cell_25_3 ( BL3, BLN3, WL25);
sram_cell_6t_3 inst_cell_25_2 ( BL2, BLN2, WL25);
sram_cell_6t_3 inst_cell_25_1 ( BL1, BLN1, WL25);
sram_cell_6t_3 inst_cell_25_0 ( BL0, BLN0, WL25);
sram_cell_6t_3 inst_cell_24_63 ( BL63, BLN63, WL24);
sram_cell_6t_3 inst_cell_24_7 ( BL7, BLN7, WL24);
sram_cell_6t_3 inst_cell_24_6 ( BL6, BLN6, WL24);
sram_cell_6t_3 inst_cell_24_5 ( BL5, BLN5, WL24);
sram_cell_6t_3 inst_cell_24_4 ( BL4, BLN4, WL24);
sram_cell_6t_3 inst_cell_24_3 ( BL3, BLN3, WL24);
sram_cell_6t_3 inst_cell_24_2 ( BL2, BLN2, WL24);
sram_cell_6t_3 inst_cell_24_1 ( BL1, BLN1, WL24);
sram_cell_6t_3 inst_cell_24_0 ( BL0, BLN0, WL24);
sram_cell_6t_3 inst_cell_23_63 ( BL63, BLN63, WL23);
sram_cell_6t_3 inst_cell_23_31 ( BL31, BLN31, WL23);
sram_cell_6t_3 inst_cell_22_31 ( BL31, BLN31, WL22);
sram_cell_6t_3 inst_cell_23_30 ( BL30, BLN30, WL23);
sram_cell_6t_3 inst_cell_22_30 ( BL30, BLN30, WL22);
sram_cell_6t_3 inst_cell_23_29 ( BL29, BLN29, WL23);
sram_cell_6t_3 inst_cell_22_29 ( BL29, BLN29, WL22);
sram_cell_6t_3 inst_cell_23_28 ( BL28, BLN28, WL23);
sram_cell_6t_3 inst_cell_22_28 ( BL28, BLN28, WL22);
sram_cell_6t_3 inst_cell_23_27 ( BL27, BLN27, WL23);
sram_cell_6t_3 inst_cell_22_27 ( BL27, BLN27, WL22);
sram_cell_6t_3 inst_cell_23_26 ( BL26, BLN26, WL23);
sram_cell_6t_3 inst_cell_22_26 ( BL26, BLN26, WL22);
sram_cell_6t_3 inst_cell_23_25 ( BL25, BLN25, WL23);
sram_cell_6t_3 inst_cell_22_25 ( BL25, BLN25, WL22);
sram_cell_6t_3 inst_cell_23_24 ( BL24, BLN24, WL23);
sram_cell_6t_3 inst_cell_22_24 ( BL24, BLN24, WL22);
sram_cell_6t_3 inst_cell_23_23 ( BL23, BLN23, WL23);
sram_cell_6t_3 inst_cell_22_23 ( BL23, BLN23, WL22);
sram_cell_6t_3 inst_cell_23_22 ( BL22, BLN22, WL23);
sram_cell_6t_3 inst_cell_22_22 ( BL22, BLN22, WL22);
sram_cell_6t_3 inst_cell_23_21 ( BL21, BLN21, WL23);
sram_cell_6t_3 inst_cell_22_21 ( BL21, BLN21, WL22);
sram_cell_6t_3 inst_cell_23_20 ( BL20, BLN20, WL23);
sram_cell_6t_3 inst_cell_22_20 ( BL20, BLN20, WL22);
sram_cell_6t_3 inst_cell_23_19 ( BL19, BLN19, WL23);
sram_cell_6t_3 inst_cell_22_19 ( BL19, BLN19, WL22);
sram_cell_6t_3 inst_cell_23_18 ( BL18, BLN18, WL23);
sram_cell_6t_3 inst_cell_22_18 ( BL18, BLN18, WL22);
sram_cell_6t_3 inst_cell_23_17 ( BL17, BLN17, WL23);
sram_cell_6t_3 inst_cell_22_17 ( BL17, BLN17, WL22);
sram_cell_6t_3 inst_cell_23_16 ( BL16, BLN16, WL23);
sram_cell_6t_3 inst_cell_22_16 ( BL16, BLN16, WL22);
sram_cell_6t_3 inst_cell_23_15 ( BL15, BLN15, WL23);
sram_cell_6t_3 inst_cell_22_15 ( BL15, BLN15, WL22);
sram_cell_6t_3 inst_cell_23_14 ( BL14, BLN14, WL23);
sram_cell_6t_3 inst_cell_22_14 ( BL14, BLN14, WL22);
sram_cell_6t_3 inst_cell_23_13 ( BL13, BLN13, WL23);
sram_cell_6t_3 inst_cell_22_13 ( BL13, BLN13, WL22);
sram_cell_6t_3 inst_cell_23_12 ( BL12, BLN12, WL23);
sram_cell_6t_3 inst_cell_22_12 ( BL12, BLN12, WL22);
sram_cell_6t_3 inst_cell_23_11 ( BL11, BLN11, WL23);
sram_cell_6t_3 inst_cell_22_11 ( BL11, BLN11, WL22);
sram_cell_6t_3 inst_cell_23_10 ( BL10, BLN10, WL23);
sram_cell_6t_3 inst_cell_22_10 ( BL10, BLN10, WL22);
sram_cell_6t_3 inst_cell_23_9 ( BL9, BLN9, WL23);
sram_cell_6t_3 inst_cell_22_9 ( BL9, BLN9, WL22);
sram_cell_6t_3 inst_cell_23_8 ( BL8, BLN8, WL23);
sram_cell_6t_3 inst_cell_22_8 ( BL8, BLN8, WL22);
sram_cell_6t_3 inst_cell_23_7 ( BL7, BLN7, WL23);
sram_cell_6t_3 inst_cell_22_7 ( BL7, BLN7, WL22);
sram_cell_6t_3 inst_cell_23_6 ( BL6, BLN6, WL23);
sram_cell_6t_3 inst_cell_22_6 ( BL6, BLN6, WL22);
sram_cell_6t_3 inst_cell_23_5 ( BL5, BLN5, WL23);
sram_cell_6t_3 inst_cell_22_5 ( BL5, BLN5, WL22);
sram_cell_6t_3 inst_cell_23_4 ( BL4, BLN4, WL23);
sram_cell_6t_3 inst_cell_22_4 ( BL4, BLN4, WL22);
sram_cell_6t_3 inst_cell_23_3 ( BL3, BLN3, WL23);
sram_cell_6t_3 inst_cell_22_3 ( BL3, BLN3, WL22);
sram_cell_6t_3 inst_cell_23_2 ( BL2, BLN2, WL23);
sram_cell_6t_3 inst_cell_22_2 ( BL2, BLN2, WL22);
sram_cell_6t_3 inst_cell_23_1 ( BL1, BLN1, WL23);
sram_cell_6t_3 inst_cell_22_1 ( BL1, BLN1, WL22);
sram_cell_6t_3 inst_cell_23_0 ( BL0, BLN0, WL23);
sram_cell_6t_3 inst_cell_22_0 ( BL0, BLN0, WL22);
sram_cell_6t_3 inst_cell_22_63 ( BL63, BLN63, WL22);
sram_cell_6t_3 inst_cell_21_63 ( BL63, BLN63, WL21);
sram_cell_6t_3 inst_cell_23_62 ( BL62, BLN62, WL23);
sram_cell_6t_3 inst_cell_23_61 ( BL61, BLN61, WL23);
sram_cell_6t_3 inst_cell_23_60 ( BL60, BLN60, WL23);
sram_cell_6t_3 inst_cell_23_59 ( BL59, BLN59, WL23);
sram_cell_6t_3 inst_cell_23_58 ( BL58, BLN58, WL23);
sram_cell_6t_3 inst_cell_23_57 ( BL57, BLN57, WL23);
sram_cell_6t_3 inst_cell_23_56 ( BL56, BLN56, WL23);
sram_cell_6t_3 inst_cell_23_55 ( BL55, BLN55, WL23);
sram_cell_6t_3 inst_cell_23_54 ( BL54, BLN54, WL23);
sram_cell_6t_3 inst_cell_23_53 ( BL53, BLN53, WL23);
sram_cell_6t_3 inst_cell_23_52 ( BL52, BLN52, WL23);
sram_cell_6t_3 inst_cell_23_51 ( BL51, BLN51, WL23);
sram_cell_6t_3 inst_cell_23_50 ( BL50, BLN50, WL23);
sram_cell_6t_3 inst_cell_23_49 ( BL49, BLN49, WL23);
sram_cell_6t_3 inst_cell_23_48 ( BL48, BLN48, WL23);
sram_cell_6t_3 inst_cell_23_47 ( BL47, BLN47, WL23);
sram_cell_6t_3 inst_cell_23_46 ( BL46, BLN46, WL23);
sram_cell_6t_3 inst_cell_23_45 ( BL45, BLN45, WL23);
sram_cell_6t_3 inst_cell_23_44 ( BL44, BLN44, WL23);
sram_cell_6t_3 inst_cell_23_43 ( BL43, BLN43, WL23);
sram_cell_6t_3 inst_cell_23_42 ( BL42, BLN42, WL23);
sram_cell_6t_3 inst_cell_23_41 ( BL41, BLN41, WL23);
sram_cell_6t_3 inst_cell_23_40 ( BL40, BLN40, WL23);
sram_cell_6t_3 inst_cell_23_39 ( BL39, BLN39, WL23);
sram_cell_6t_3 inst_cell_23_38 ( BL38, BLN38, WL23);
sram_cell_6t_3 inst_cell_23_37 ( BL37, BLN37, WL23);
sram_cell_6t_3 inst_cell_23_36 ( BL36, BLN36, WL23);
sram_cell_6t_3 inst_cell_23_35 ( BL35, BLN35, WL23);
sram_cell_6t_3 inst_cell_23_34 ( BL34, BLN34, WL23);
sram_cell_6t_3 inst_cell_23_33 ( BL33, BLN33, WL23);
sram_cell_6t_3 inst_cell_23_32 ( BL32, BLN32, WL23);
sram_cell_6t_3 inst_cell_22_62 ( BL62, BLN62, WL22);
sram_cell_6t_3 inst_cell_22_61 ( BL61, BLN61, WL22);
sram_cell_6t_3 inst_cell_22_60 ( BL60, BLN60, WL22);
sram_cell_6t_3 inst_cell_22_59 ( BL59, BLN59, WL22);
sram_cell_6t_3 inst_cell_22_58 ( BL58, BLN58, WL22);
sram_cell_6t_3 inst_cell_22_57 ( BL57, BLN57, WL22);
sram_cell_6t_3 inst_cell_22_56 ( BL56, BLN56, WL22);
sram_cell_6t_3 inst_cell_22_55 ( BL55, BLN55, WL22);
sram_cell_6t_3 inst_cell_22_54 ( BL54, BLN54, WL22);
sram_cell_6t_3 inst_cell_22_53 ( BL53, BLN53, WL22);
sram_cell_6t_3 inst_cell_22_52 ( BL52, BLN52, WL22);
sram_cell_6t_3 inst_cell_22_51 ( BL51, BLN51, WL22);
sram_cell_6t_3 inst_cell_22_50 ( BL50, BLN50, WL22);
sram_cell_6t_3 inst_cell_22_49 ( BL49, BLN49, WL22);
sram_cell_6t_3 inst_cell_22_48 ( BL48, BLN48, WL22);
sram_cell_6t_3 inst_cell_22_47 ( BL47, BLN47, WL22);
sram_cell_6t_3 inst_cell_22_46 ( BL46, BLN46, WL22);
sram_cell_6t_3 inst_cell_22_45 ( BL45, BLN45, WL22);
sram_cell_6t_3 inst_cell_22_44 ( BL44, BLN44, WL22);
sram_cell_6t_3 inst_cell_22_43 ( BL43, BLN43, WL22);
sram_cell_6t_3 inst_cell_22_42 ( BL42, BLN42, WL22);
sram_cell_6t_3 inst_cell_22_41 ( BL41, BLN41, WL22);
sram_cell_6t_3 inst_cell_22_40 ( BL40, BLN40, WL22);
sram_cell_6t_3 inst_cell_22_39 ( BL39, BLN39, WL22);
sram_cell_6t_3 inst_cell_22_38 ( BL38, BLN38, WL22);
sram_cell_6t_3 inst_cell_22_37 ( BL37, BLN37, WL22);
sram_cell_6t_3 inst_cell_22_36 ( BL36, BLN36, WL22);
sram_cell_6t_3 inst_cell_22_35 ( BL35, BLN35, WL22);
sram_cell_6t_3 inst_cell_22_34 ( BL34, BLN34, WL22);
sram_cell_6t_3 inst_cell_22_33 ( BL33, BLN33, WL22);
sram_cell_6t_3 inst_cell_22_32 ( BL32, BLN32, WL22);
sram_cell_6t_3 inst_cell_21_62 ( BL62, BLN62, WL21);
sram_cell_6t_3 inst_cell_21_61 ( BL61, BLN61, WL21);
sram_cell_6t_3 inst_cell_21_60 ( BL60, BLN60, WL21);
sram_cell_6t_3 inst_cell_21_59 ( BL59, BLN59, WL21);
sram_cell_6t_3 inst_cell_21_58 ( BL58, BLN58, WL21);
sram_cell_6t_3 inst_cell_21_57 ( BL57, BLN57, WL21);
sram_cell_6t_3 inst_cell_21_56 ( BL56, BLN56, WL21);
sram_cell_6t_3 inst_cell_21_55 ( BL55, BLN55, WL21);
sram_cell_6t_3 inst_cell_21_54 ( BL54, BLN54, WL21);
sram_cell_6t_3 inst_cell_21_53 ( BL53, BLN53, WL21);
sram_cell_6t_3 inst_cell_21_52 ( BL52, BLN52, WL21);
sram_cell_6t_3 inst_cell_21_51 ( BL51, BLN51, WL21);
sram_cell_6t_3 inst_cell_21_50 ( BL50, BLN50, WL21);
sram_cell_6t_3 inst_cell_21_49 ( BL49, BLN49, WL21);
sram_cell_6t_3 inst_cell_21_48 ( BL48, BLN48, WL21);
sram_cell_6t_3 inst_cell_21_47 ( BL47, BLN47, WL21);
sram_cell_6t_3 inst_cell_21_46 ( BL46, BLN46, WL21);
sram_cell_6t_3 inst_cell_21_45 ( BL45, BLN45, WL21);
sram_cell_6t_3 inst_cell_21_44 ( BL44, BLN44, WL21);
sram_cell_6t_3 inst_cell_21_43 ( BL43, BLN43, WL21);
sram_cell_6t_3 inst_cell_21_42 ( BL42, BLN42, WL21);
sram_cell_6t_3 inst_cell_21_41 ( BL41, BLN41, WL21);
sram_cell_6t_3 inst_cell_21_40 ( BL40, BLN40, WL21);
sram_cell_6t_3 inst_cell_21_39 ( BL39, BLN39, WL21);
sram_cell_6t_3 inst_cell_21_38 ( BL38, BLN38, WL21);
sram_cell_6t_3 inst_cell_21_37 ( BL37, BLN37, WL21);
sram_cell_6t_3 inst_cell_21_36 ( BL36, BLN36, WL21);
sram_cell_6t_3 inst_cell_21_35 ( BL35, BLN35, WL21);
sram_cell_6t_3 inst_cell_21_34 ( BL34, BLN34, WL21);
sram_cell_6t_3 inst_cell_21_33 ( BL33, BLN33, WL21);
sram_cell_6t_3 inst_cell_21_32 ( BL32, BLN32, WL21);
sram_cell_6t_3 inst_cell_21_7 ( BL7, BLN7, WL21);
sram_cell_6t_3 inst_cell_20_7 ( BL7, BLN7, WL20);
sram_cell_6t_3 inst_cell_21_6 ( BL6, BLN6, WL21);
sram_cell_6t_3 inst_cell_20_6 ( BL6, BLN6, WL20);
sram_cell_6t_3 inst_cell_21_5 ( BL5, BLN5, WL21);
sram_cell_6t_3 inst_cell_20_5 ( BL5, BLN5, WL20);
sram_cell_6t_3 inst_cell_21_4 ( BL4, BLN4, WL21);
sram_cell_6t_3 inst_cell_20_4 ( BL4, BLN4, WL20);
sram_cell_6t_3 inst_cell_21_3 ( BL3, BLN3, WL21);
sram_cell_6t_3 inst_cell_20_3 ( BL3, BLN3, WL20);
sram_cell_6t_3 inst_cell_21_2 ( BL2, BLN2, WL21);
sram_cell_6t_3 inst_cell_20_2 ( BL2, BLN2, WL20);
sram_cell_6t_3 inst_cell_21_1 ( BL1, BLN1, WL21);
sram_cell_6t_3 inst_cell_20_1 ( BL1, BLN1, WL20);
sram_cell_6t_3 inst_cell_21_0 ( BL0, BLN0, WL21);
sram_cell_6t_3 inst_cell_20_0 ( BL0, BLN0, WL20);
sram_cell_6t_3 inst_cell_20_63 ( BL63, BLN63, WL20);
sram_cell_6t_3 inst_cell_19_63 ( BL63, BLN63, WL19);
sram_cell_6t_3 inst_cell_20_62 ( BL62, BLN62, WL20);
sram_cell_6t_3 inst_cell_19_62 ( BL62, BLN62, WL19);
sram_cell_6t_3 inst_cell_20_61 ( BL61, BLN61, WL20);
sram_cell_6t_3 inst_cell_19_61 ( BL61, BLN61, WL19);
sram_cell_6t_3 inst_cell_20_60 ( BL60, BLN60, WL20);
sram_cell_6t_3 inst_cell_19_60 ( BL60, BLN60, WL19);
sram_cell_6t_3 inst_cell_20_59 ( BL59, BLN59, WL20);
sram_cell_6t_3 inst_cell_19_59 ( BL59, BLN59, WL19);
sram_cell_6t_3 inst_cell_20_58 ( BL58, BLN58, WL20);
sram_cell_6t_3 inst_cell_19_58 ( BL58, BLN58, WL19);
sram_cell_6t_3 inst_cell_20_57 ( BL57, BLN57, WL20);
sram_cell_6t_3 inst_cell_19_57 ( BL57, BLN57, WL19);
sram_cell_6t_3 inst_cell_20_56 ( BL56, BLN56, WL20);
sram_cell_6t_3 inst_cell_19_56 ( BL56, BLN56, WL19);
sram_cell_6t_3 inst_cell_20_55 ( BL55, BLN55, WL20);
sram_cell_6t_3 inst_cell_19_55 ( BL55, BLN55, WL19);
sram_cell_6t_3 inst_cell_20_54 ( BL54, BLN54, WL20);
sram_cell_6t_3 inst_cell_19_54 ( BL54, BLN54, WL19);
sram_cell_6t_3 inst_cell_20_53 ( BL53, BLN53, WL20);
sram_cell_6t_3 inst_cell_19_53 ( BL53, BLN53, WL19);
sram_cell_6t_3 inst_cell_20_52 ( BL52, BLN52, WL20);
sram_cell_6t_3 inst_cell_19_52 ( BL52, BLN52, WL19);
sram_cell_6t_3 inst_cell_20_51 ( BL51, BLN51, WL20);
sram_cell_6t_3 inst_cell_19_51 ( BL51, BLN51, WL19);
sram_cell_6t_3 inst_cell_20_50 ( BL50, BLN50, WL20);
sram_cell_6t_3 inst_cell_19_50 ( BL50, BLN50, WL19);
sram_cell_6t_3 inst_cell_20_49 ( BL49, BLN49, WL20);
sram_cell_6t_3 inst_cell_19_49 ( BL49, BLN49, WL19);
sram_cell_6t_3 inst_cell_20_48 ( BL48, BLN48, WL20);
sram_cell_6t_3 inst_cell_19_48 ( BL48, BLN48, WL19);
sram_cell_6t_3 inst_cell_20_47 ( BL47, BLN47, WL20);
sram_cell_6t_3 inst_cell_19_47 ( BL47, BLN47, WL19);
sram_cell_6t_3 inst_cell_20_46 ( BL46, BLN46, WL20);
sram_cell_6t_3 inst_cell_19_46 ( BL46, BLN46, WL19);
sram_cell_6t_3 inst_cell_20_45 ( BL45, BLN45, WL20);
sram_cell_6t_3 inst_cell_19_45 ( BL45, BLN45, WL19);
sram_cell_6t_3 inst_cell_20_44 ( BL44, BLN44, WL20);
sram_cell_6t_3 inst_cell_19_44 ( BL44, BLN44, WL19);
sram_cell_6t_3 inst_cell_20_43 ( BL43, BLN43, WL20);
sram_cell_6t_3 inst_cell_19_43 ( BL43, BLN43, WL19);
sram_cell_6t_3 inst_cell_20_42 ( BL42, BLN42, WL20);
sram_cell_6t_3 inst_cell_19_42 ( BL42, BLN42, WL19);
sram_cell_6t_3 inst_cell_20_41 ( BL41, BLN41, WL20);
sram_cell_6t_3 inst_cell_19_41 ( BL41, BLN41, WL19);
sram_cell_6t_3 inst_cell_20_40 ( BL40, BLN40, WL20);
sram_cell_6t_3 inst_cell_19_40 ( BL40, BLN40, WL19);
sram_cell_6t_3 inst_cell_20_39 ( BL39, BLN39, WL20);
sram_cell_6t_3 inst_cell_19_39 ( BL39, BLN39, WL19);
sram_cell_6t_3 inst_cell_20_38 ( BL38, BLN38, WL20);
sram_cell_6t_3 inst_cell_19_38 ( BL38, BLN38, WL19);
sram_cell_6t_3 inst_cell_20_37 ( BL37, BLN37, WL20);
sram_cell_6t_3 inst_cell_19_37 ( BL37, BLN37, WL19);
sram_cell_6t_3 inst_cell_20_36 ( BL36, BLN36, WL20);
sram_cell_6t_3 inst_cell_19_36 ( BL36, BLN36, WL19);
sram_cell_6t_3 inst_cell_20_35 ( BL35, BLN35, WL20);
sram_cell_6t_3 inst_cell_19_35 ( BL35, BLN35, WL19);
sram_cell_6t_3 inst_cell_20_34 ( BL34, BLN34, WL20);
sram_cell_6t_3 inst_cell_19_34 ( BL34, BLN34, WL19);
sram_cell_6t_3 inst_cell_20_33 ( BL33, BLN33, WL20);
sram_cell_6t_3 inst_cell_19_33 ( BL33, BLN33, WL19);
sram_cell_6t_3 inst_cell_20_32 ( BL32, BLN32, WL20);
sram_cell_6t_3 inst_cell_19_32 ( BL32, BLN32, WL19);
sram_cell_6t_3 inst_cell_21_31 ( BL31, BLN31, WL21);
sram_cell_6t_3 inst_cell_21_30 ( BL30, BLN30, WL21);
sram_cell_6t_3 inst_cell_21_29 ( BL29, BLN29, WL21);
sram_cell_6t_3 inst_cell_21_28 ( BL28, BLN28, WL21);
sram_cell_6t_3 inst_cell_21_27 ( BL27, BLN27, WL21);
sram_cell_6t_3 inst_cell_21_26 ( BL26, BLN26, WL21);
sram_cell_6t_3 inst_cell_21_25 ( BL25, BLN25, WL21);
sram_cell_6t_3 inst_cell_21_24 ( BL24, BLN24, WL21);
sram_cell_6t_3 inst_cell_21_23 ( BL23, BLN23, WL21);
sram_cell_6t_3 inst_cell_21_22 ( BL22, BLN22, WL21);
sram_cell_6t_3 inst_cell_21_21 ( BL21, BLN21, WL21);
sram_cell_6t_3 inst_cell_21_20 ( BL20, BLN20, WL21);
sram_cell_6t_3 inst_cell_21_19 ( BL19, BLN19, WL21);
sram_cell_6t_3 inst_cell_21_18 ( BL18, BLN18, WL21);
sram_cell_6t_3 inst_cell_21_17 ( BL17, BLN17, WL21);
sram_cell_6t_3 inst_cell_21_16 ( BL16, BLN16, WL21);
sram_cell_6t_3 inst_cell_21_15 ( BL15, BLN15, WL21);
sram_cell_6t_3 inst_cell_21_14 ( BL14, BLN14, WL21);
sram_cell_6t_3 inst_cell_21_13 ( BL13, BLN13, WL21);
sram_cell_6t_3 inst_cell_21_12 ( BL12, BLN12, WL21);
sram_cell_6t_3 inst_cell_21_11 ( BL11, BLN11, WL21);
sram_cell_6t_3 inst_cell_21_10 ( BL10, BLN10, WL21);
sram_cell_6t_3 inst_cell_21_9 ( BL9, BLN9, WL21);
sram_cell_6t_3 inst_cell_21_8 ( BL8, BLN8, WL21);
sram_cell_6t_3 inst_cell_20_31 ( BL31, BLN31, WL20);
sram_cell_6t_3 inst_cell_20_30 ( BL30, BLN30, WL20);
sram_cell_6t_3 inst_cell_20_29 ( BL29, BLN29, WL20);
sram_cell_6t_3 inst_cell_20_28 ( BL28, BLN28, WL20);
sram_cell_6t_3 inst_cell_20_27 ( BL27, BLN27, WL20);
sram_cell_6t_3 inst_cell_20_26 ( BL26, BLN26, WL20);
sram_cell_6t_3 inst_cell_20_25 ( BL25, BLN25, WL20);
sram_cell_6t_3 inst_cell_20_24 ( BL24, BLN24, WL20);
sram_cell_6t_3 inst_cell_20_23 ( BL23, BLN23, WL20);
sram_cell_6t_3 inst_cell_20_22 ( BL22, BLN22, WL20);
sram_cell_6t_3 inst_cell_20_21 ( BL21, BLN21, WL20);
sram_cell_6t_3 inst_cell_20_20 ( BL20, BLN20, WL20);
sram_cell_6t_3 inst_cell_20_19 ( BL19, BLN19, WL20);
sram_cell_6t_3 inst_cell_20_18 ( BL18, BLN18, WL20);
sram_cell_6t_3 inst_cell_20_17 ( BL17, BLN17, WL20);
sram_cell_6t_3 inst_cell_20_16 ( BL16, BLN16, WL20);
sram_cell_6t_3 inst_cell_20_15 ( BL15, BLN15, WL20);
sram_cell_6t_3 inst_cell_20_14 ( BL14, BLN14, WL20);
sram_cell_6t_3 inst_cell_20_13 ( BL13, BLN13, WL20);
sram_cell_6t_3 inst_cell_20_12 ( BL12, BLN12, WL20);
sram_cell_6t_3 inst_cell_20_11 ( BL11, BLN11, WL20);
sram_cell_6t_3 inst_cell_20_10 ( BL10, BLN10, WL20);
sram_cell_6t_3 inst_cell_20_9 ( BL9, BLN9, WL20);
sram_cell_6t_3 inst_cell_20_8 ( BL8, BLN8, WL20);
sram_cell_6t_3 inst_cell_19_31 ( BL31, BLN31, WL19);
sram_cell_6t_3 inst_cell_19_30 ( BL30, BLN30, WL19);
sram_cell_6t_3 inst_cell_19_29 ( BL29, BLN29, WL19);
sram_cell_6t_3 inst_cell_19_28 ( BL28, BLN28, WL19);
sram_cell_6t_3 inst_cell_19_27 ( BL27, BLN27, WL19);
sram_cell_6t_3 inst_cell_19_26 ( BL26, BLN26, WL19);
sram_cell_6t_3 inst_cell_19_25 ( BL25, BLN25, WL19);
sram_cell_6t_3 inst_cell_19_24 ( BL24, BLN24, WL19);
sram_cell_6t_3 inst_cell_19_23 ( BL23, BLN23, WL19);
sram_cell_6t_3 inst_cell_19_22 ( BL22, BLN22, WL19);
sram_cell_6t_3 inst_cell_19_21 ( BL21, BLN21, WL19);
sram_cell_6t_3 inst_cell_19_20 ( BL20, BLN20, WL19);
sram_cell_6t_3 inst_cell_19_19 ( BL19, BLN19, WL19);
sram_cell_6t_3 inst_cell_19_18 ( BL18, BLN18, WL19);
sram_cell_6t_3 inst_cell_19_17 ( BL17, BLN17, WL19);
sram_cell_6t_3 inst_cell_19_16 ( BL16, BLN16, WL19);
sram_cell_6t_3 inst_cell_19_15 ( BL15, BLN15, WL19);
sram_cell_6t_3 inst_cell_19_14 ( BL14, BLN14, WL19);
sram_cell_6t_3 inst_cell_19_13 ( BL13, BLN13, WL19);
sram_cell_6t_3 inst_cell_19_12 ( BL12, BLN12, WL19);
sram_cell_6t_3 inst_cell_19_11 ( BL11, BLN11, WL19);
sram_cell_6t_3 inst_cell_19_10 ( BL10, BLN10, WL19);
sram_cell_6t_3 inst_cell_19_9 ( BL9, BLN9, WL19);
sram_cell_6t_3 inst_cell_19_8 ( BL8, BLN8, WL19);
sram_cell_6t_3 inst_cell_18_62 ( BL62, BLN62, WL18);
sram_cell_6t_3 inst_cell_17_62 ( BL62, BLN62, WL17);
sram_cell_6t_3 inst_cell_18_61 ( BL61, BLN61, WL18);
sram_cell_6t_3 inst_cell_17_61 ( BL61, BLN61, WL17);
sram_cell_6t_3 inst_cell_18_60 ( BL60, BLN60, WL18);
sram_cell_6t_3 inst_cell_17_60 ( BL60, BLN60, WL17);
sram_cell_6t_3 inst_cell_18_59 ( BL59, BLN59, WL18);
sram_cell_6t_3 inst_cell_17_59 ( BL59, BLN59, WL17);
sram_cell_6t_3 inst_cell_18_58 ( BL58, BLN58, WL18);
sram_cell_6t_3 inst_cell_17_58 ( BL58, BLN58, WL17);
sram_cell_6t_3 inst_cell_18_57 ( BL57, BLN57, WL18);
sram_cell_6t_3 inst_cell_17_57 ( BL57, BLN57, WL17);
sram_cell_6t_3 inst_cell_18_56 ( BL56, BLN56, WL18);
sram_cell_6t_3 inst_cell_17_56 ( BL56, BLN56, WL17);
sram_cell_6t_3 inst_cell_18_55 ( BL55, BLN55, WL18);
sram_cell_6t_3 inst_cell_17_55 ( BL55, BLN55, WL17);
sram_cell_6t_3 inst_cell_18_54 ( BL54, BLN54, WL18);
sram_cell_6t_3 inst_cell_17_54 ( BL54, BLN54, WL17);
sram_cell_6t_3 inst_cell_18_53 ( BL53, BLN53, WL18);
sram_cell_6t_3 inst_cell_17_53 ( BL53, BLN53, WL17);
sram_cell_6t_3 inst_cell_18_52 ( BL52, BLN52, WL18);
sram_cell_6t_3 inst_cell_17_52 ( BL52, BLN52, WL17);
sram_cell_6t_3 inst_cell_18_51 ( BL51, BLN51, WL18);
sram_cell_6t_3 inst_cell_17_51 ( BL51, BLN51, WL17);
sram_cell_6t_3 inst_cell_18_50 ( BL50, BLN50, WL18);
sram_cell_6t_3 inst_cell_17_50 ( BL50, BLN50, WL17);
sram_cell_6t_3 inst_cell_18_49 ( BL49, BLN49, WL18);
sram_cell_6t_3 inst_cell_17_49 ( BL49, BLN49, WL17);
sram_cell_6t_3 inst_cell_18_48 ( BL48, BLN48, WL18);
sram_cell_6t_3 inst_cell_17_48 ( BL48, BLN48, WL17);
sram_cell_6t_3 inst_cell_18_47 ( BL47, BLN47, WL18);
sram_cell_6t_3 inst_cell_17_47 ( BL47, BLN47, WL17);
sram_cell_6t_3 inst_cell_18_46 ( BL46, BLN46, WL18);
sram_cell_6t_3 inst_cell_17_46 ( BL46, BLN46, WL17);
sram_cell_6t_3 inst_cell_18_45 ( BL45, BLN45, WL18);
sram_cell_6t_3 inst_cell_17_45 ( BL45, BLN45, WL17);
sram_cell_6t_3 inst_cell_18_44 ( BL44, BLN44, WL18);
sram_cell_6t_3 inst_cell_17_44 ( BL44, BLN44, WL17);
sram_cell_6t_3 inst_cell_18_43 ( BL43, BLN43, WL18);
sram_cell_6t_3 inst_cell_17_43 ( BL43, BLN43, WL17);
sram_cell_6t_3 inst_cell_18_42 ( BL42, BLN42, WL18);
sram_cell_6t_3 inst_cell_17_42 ( BL42, BLN42, WL17);
sram_cell_6t_3 inst_cell_18_41 ( BL41, BLN41, WL18);
sram_cell_6t_3 inst_cell_17_41 ( BL41, BLN41, WL17);
sram_cell_6t_3 inst_cell_18_40 ( BL40, BLN40, WL18);
sram_cell_6t_3 inst_cell_17_40 ( BL40, BLN40, WL17);
sram_cell_6t_3 inst_cell_18_39 ( BL39, BLN39, WL18);
sram_cell_6t_3 inst_cell_17_39 ( BL39, BLN39, WL17);
sram_cell_6t_3 inst_cell_18_38 ( BL38, BLN38, WL18);
sram_cell_6t_3 inst_cell_17_38 ( BL38, BLN38, WL17);
sram_cell_6t_3 inst_cell_18_37 ( BL37, BLN37, WL18);
sram_cell_6t_3 inst_cell_17_37 ( BL37, BLN37, WL17);
sram_cell_6t_3 inst_cell_18_36 ( BL36, BLN36, WL18);
sram_cell_6t_3 inst_cell_17_36 ( BL36, BLN36, WL17);
sram_cell_6t_3 inst_cell_18_35 ( BL35, BLN35, WL18);
sram_cell_6t_3 inst_cell_17_35 ( BL35, BLN35, WL17);
sram_cell_6t_3 inst_cell_18_34 ( BL34, BLN34, WL18);
sram_cell_6t_3 inst_cell_17_34 ( BL34, BLN34, WL17);
sram_cell_6t_3 inst_cell_18_33 ( BL33, BLN33, WL18);
sram_cell_6t_3 inst_cell_17_33 ( BL33, BLN33, WL17);
sram_cell_6t_3 inst_cell_18_32 ( BL32, BLN32, WL18);
sram_cell_6t_3 inst_cell_17_32 ( BL32, BLN32, WL17);
sram_cell_6t_3 inst_cell_18_31 ( BL31, BLN31, WL18);
sram_cell_6t_3 inst_cell_17_31 ( BL31, BLN31, WL17);
sram_cell_6t_3 inst_cell_18_30 ( BL30, BLN30, WL18);
sram_cell_6t_3 inst_cell_17_30 ( BL30, BLN30, WL17);
sram_cell_6t_3 inst_cell_18_29 ( BL29, BLN29, WL18);
sram_cell_6t_3 inst_cell_17_29 ( BL29, BLN29, WL17);
sram_cell_6t_3 inst_cell_18_28 ( BL28, BLN28, WL18);
sram_cell_6t_3 inst_cell_17_28 ( BL28, BLN28, WL17);
sram_cell_6t_3 inst_cell_18_27 ( BL27, BLN27, WL18);
sram_cell_6t_3 inst_cell_17_27 ( BL27, BLN27, WL17);
sram_cell_6t_3 inst_cell_18_26 ( BL26, BLN26, WL18);
sram_cell_6t_3 inst_cell_17_26 ( BL26, BLN26, WL17);
sram_cell_6t_3 inst_cell_18_25 ( BL25, BLN25, WL18);
sram_cell_6t_3 inst_cell_17_25 ( BL25, BLN25, WL17);
sram_cell_6t_3 inst_cell_18_24 ( BL24, BLN24, WL18);
sram_cell_6t_3 inst_cell_17_24 ( BL24, BLN24, WL17);
sram_cell_6t_3 inst_cell_18_23 ( BL23, BLN23, WL18);
sram_cell_6t_3 inst_cell_17_23 ( BL23, BLN23, WL17);
sram_cell_6t_3 inst_cell_18_22 ( BL22, BLN22, WL18);
sram_cell_6t_3 inst_cell_17_22 ( BL22, BLN22, WL17);
sram_cell_6t_3 inst_cell_18_21 ( BL21, BLN21, WL18);
sram_cell_6t_3 inst_cell_17_21 ( BL21, BLN21, WL17);
sram_cell_6t_3 inst_cell_18_20 ( BL20, BLN20, WL18);
sram_cell_6t_3 inst_cell_17_20 ( BL20, BLN20, WL17);
sram_cell_6t_3 inst_cell_18_19 ( BL19, BLN19, WL18);
sram_cell_6t_3 inst_cell_17_19 ( BL19, BLN19, WL17);
sram_cell_6t_3 inst_cell_18_18 ( BL18, BLN18, WL18);
sram_cell_6t_3 inst_cell_17_18 ( BL18, BLN18, WL17);
sram_cell_6t_3 inst_cell_18_17 ( BL17, BLN17, WL18);
sram_cell_6t_3 inst_cell_17_17 ( BL17, BLN17, WL17);
sram_cell_6t_3 inst_cell_18_16 ( BL16, BLN16, WL18);
sram_cell_6t_3 inst_cell_17_16 ( BL16, BLN16, WL17);
sram_cell_6t_3 inst_cell_18_15 ( BL15, BLN15, WL18);
sram_cell_6t_3 inst_cell_17_15 ( BL15, BLN15, WL17);
sram_cell_6t_3 inst_cell_18_14 ( BL14, BLN14, WL18);
sram_cell_6t_3 inst_cell_17_14 ( BL14, BLN14, WL17);
sram_cell_6t_3 inst_cell_18_13 ( BL13, BLN13, WL18);
sram_cell_6t_3 inst_cell_17_13 ( BL13, BLN13, WL17);
sram_cell_6t_3 inst_cell_18_12 ( BL12, BLN12, WL18);
sram_cell_6t_3 inst_cell_17_12 ( BL12, BLN12, WL17);
sram_cell_6t_3 inst_cell_18_11 ( BL11, BLN11, WL18);
sram_cell_6t_3 inst_cell_17_11 ( BL11, BLN11, WL17);
sram_cell_6t_3 inst_cell_18_10 ( BL10, BLN10, WL18);
sram_cell_6t_3 inst_cell_17_10 ( BL10, BLN10, WL17);
sram_cell_6t_3 inst_cell_18_9 ( BL9, BLN9, WL18);
sram_cell_6t_3 inst_cell_17_9 ( BL9, BLN9, WL17);
sram_cell_6t_3 inst_cell_18_8 ( BL8, BLN8, WL18);
sram_cell_6t_3 inst_cell_17_8 ( BL8, BLN8, WL17);
sram_cell_6t_3 inst_cell_19_7 ( BL7, BLN7, WL19);
sram_cell_6t_3 inst_cell_19_6 ( BL6, BLN6, WL19);
sram_cell_6t_3 inst_cell_19_5 ( BL5, BLN5, WL19);
sram_cell_6t_3 inst_cell_19_4 ( BL4, BLN4, WL19);
sram_cell_6t_3 inst_cell_19_3 ( BL3, BLN3, WL19);
sram_cell_6t_3 inst_cell_19_2 ( BL2, BLN2, WL19);
sram_cell_6t_3 inst_cell_19_1 ( BL1, BLN1, WL19);
sram_cell_6t_3 inst_cell_19_0 ( BL0, BLN0, WL19);
sram_cell_6t_3 inst_cell_18_63 ( BL63, BLN63, WL18);
sram_cell_6t_3 inst_cell_18_7 ( BL7, BLN7, WL18);
sram_cell_6t_3 inst_cell_18_6 ( BL6, BLN6, WL18);
sram_cell_6t_3 inst_cell_18_5 ( BL5, BLN5, WL18);
sram_cell_6t_3 inst_cell_18_4 ( BL4, BLN4, WL18);
sram_cell_6t_3 inst_cell_18_3 ( BL3, BLN3, WL18);
sram_cell_6t_3 inst_cell_18_2 ( BL2, BLN2, WL18);
sram_cell_6t_3 inst_cell_18_1 ( BL1, BLN1, WL18);
sram_cell_6t_3 inst_cell_18_0 ( BL0, BLN0, WL18);
sram_cell_6t_3 inst_cell_17_63 ( BL63, BLN63, WL17);
sram_cell_6t_3 inst_cell_17_7 ( BL7, BLN7, WL17);
sram_cell_6t_3 inst_cell_17_6 ( BL6, BLN6, WL17);
sram_cell_6t_3 inst_cell_17_5 ( BL5, BLN5, WL17);
sram_cell_6t_3 inst_cell_17_4 ( BL4, BLN4, WL17);
sram_cell_6t_3 inst_cell_17_3 ( BL3, BLN3, WL17);
sram_cell_6t_3 inst_cell_17_2 ( BL2, BLN2, WL17);
sram_cell_6t_3 inst_cell_17_1 ( BL1, BLN1, WL17);
sram_cell_6t_3 inst_cell_17_0 ( BL0, BLN0, WL17);
sram_cell_6t_3 inst_cell_16_63 ( BL63, BLN63, WL16);
sram_cell_6t_3 inst_cell_16_31 ( BL31, BLN31, WL16);
sram_cell_6t_3 inst_cell_15_31 ( BL31, BLN31, WL15);
sram_cell_6t_3 inst_cell_16_30 ( BL30, BLN30, WL16);
sram_cell_6t_3 inst_cell_15_30 ( BL30, BLN30, WL15);
sram_cell_6t_3 inst_cell_16_29 ( BL29, BLN29, WL16);
sram_cell_6t_3 inst_cell_15_29 ( BL29, BLN29, WL15);
sram_cell_6t_3 inst_cell_16_28 ( BL28, BLN28, WL16);
sram_cell_6t_3 inst_cell_15_28 ( BL28, BLN28, WL15);
sram_cell_6t_3 inst_cell_16_27 ( BL27, BLN27, WL16);
sram_cell_6t_3 inst_cell_15_27 ( BL27, BLN27, WL15);
sram_cell_6t_3 inst_cell_16_26 ( BL26, BLN26, WL16);
sram_cell_6t_3 inst_cell_15_26 ( BL26, BLN26, WL15);
sram_cell_6t_3 inst_cell_16_25 ( BL25, BLN25, WL16);
sram_cell_6t_3 inst_cell_15_25 ( BL25, BLN25, WL15);
sram_cell_6t_3 inst_cell_16_24 ( BL24, BLN24, WL16);
sram_cell_6t_3 inst_cell_15_24 ( BL24, BLN24, WL15);
sram_cell_6t_3 inst_cell_16_23 ( BL23, BLN23, WL16);
sram_cell_6t_3 inst_cell_15_23 ( BL23, BLN23, WL15);
sram_cell_6t_3 inst_cell_16_22 ( BL22, BLN22, WL16);
sram_cell_6t_3 inst_cell_15_22 ( BL22, BLN22, WL15);
sram_cell_6t_3 inst_cell_16_21 ( BL21, BLN21, WL16);
sram_cell_6t_3 inst_cell_15_21 ( BL21, BLN21, WL15);
sram_cell_6t_3 inst_cell_16_20 ( BL20, BLN20, WL16);
sram_cell_6t_3 inst_cell_15_20 ( BL20, BLN20, WL15);
sram_cell_6t_3 inst_cell_16_19 ( BL19, BLN19, WL16);
sram_cell_6t_3 inst_cell_15_19 ( BL19, BLN19, WL15);
sram_cell_6t_3 inst_cell_16_18 ( BL18, BLN18, WL16);
sram_cell_6t_3 inst_cell_15_18 ( BL18, BLN18, WL15);
sram_cell_6t_3 inst_cell_16_17 ( BL17, BLN17, WL16);
sram_cell_6t_3 inst_cell_15_17 ( BL17, BLN17, WL15);
sram_cell_6t_3 inst_cell_16_16 ( BL16, BLN16, WL16);
sram_cell_6t_3 inst_cell_15_16 ( BL16, BLN16, WL15);
sram_cell_6t_3 inst_cell_16_15 ( BL15, BLN15, WL16);
sram_cell_6t_3 inst_cell_15_15 ( BL15, BLN15, WL15);
sram_cell_6t_3 inst_cell_16_14 ( BL14, BLN14, WL16);
sram_cell_6t_3 inst_cell_15_14 ( BL14, BLN14, WL15);
sram_cell_6t_3 inst_cell_16_13 ( BL13, BLN13, WL16);
sram_cell_6t_3 inst_cell_15_13 ( BL13, BLN13, WL15);
sram_cell_6t_3 inst_cell_16_12 ( BL12, BLN12, WL16);
sram_cell_6t_3 inst_cell_15_12 ( BL12, BLN12, WL15);
sram_cell_6t_3 inst_cell_16_11 ( BL11, BLN11, WL16);
sram_cell_6t_3 inst_cell_15_11 ( BL11, BLN11, WL15);
sram_cell_6t_3 inst_cell_16_10 ( BL10, BLN10, WL16);
sram_cell_6t_3 inst_cell_15_10 ( BL10, BLN10, WL15);
sram_cell_6t_3 inst_cell_16_9 ( BL9, BLN9, WL16);
sram_cell_6t_3 inst_cell_15_9 ( BL9, BLN9, WL15);
sram_cell_6t_3 inst_cell_16_8 ( BL8, BLN8, WL16);
sram_cell_6t_3 inst_cell_15_8 ( BL8, BLN8, WL15);
sram_cell_6t_3 inst_cell_16_7 ( BL7, BLN7, WL16);
sram_cell_6t_3 inst_cell_15_7 ( BL7, BLN7, WL15);
sram_cell_6t_3 inst_cell_16_6 ( BL6, BLN6, WL16);
sram_cell_6t_3 inst_cell_15_6 ( BL6, BLN6, WL15);
sram_cell_6t_3 inst_cell_16_5 ( BL5, BLN5, WL16);
sram_cell_6t_3 inst_cell_15_5 ( BL5, BLN5, WL15);
sram_cell_6t_3 inst_cell_16_4 ( BL4, BLN4, WL16);
sram_cell_6t_3 inst_cell_15_4 ( BL4, BLN4, WL15);
sram_cell_6t_3 inst_cell_16_3 ( BL3, BLN3, WL16);
sram_cell_6t_3 inst_cell_15_3 ( BL3, BLN3, WL15);
sram_cell_6t_3 inst_cell_16_2 ( BL2, BLN2, WL16);
sram_cell_6t_3 inst_cell_15_2 ( BL2, BLN2, WL15);
sram_cell_6t_3 inst_cell_16_1 ( BL1, BLN1, WL16);
sram_cell_6t_3 inst_cell_15_1 ( BL1, BLN1, WL15);
sram_cell_6t_3 inst_cell_16_0 ( BL0, BLN0, WL16);
sram_cell_6t_3 inst_cell_15_0 ( BL0, BLN0, WL15);
sram_cell_6t_3 inst_cell_15_63 ( BL63, BLN63, WL15);
sram_cell_6t_3 inst_cell_14_63 ( BL63, BLN63, WL14);
sram_cell_6t_3 inst_cell_16_62 ( BL62, BLN62, WL16);
sram_cell_6t_3 inst_cell_16_61 ( BL61, BLN61, WL16);
sram_cell_6t_3 inst_cell_16_60 ( BL60, BLN60, WL16);
sram_cell_6t_3 inst_cell_16_59 ( BL59, BLN59, WL16);
sram_cell_6t_3 inst_cell_16_58 ( BL58, BLN58, WL16);
sram_cell_6t_3 inst_cell_16_57 ( BL57, BLN57, WL16);
sram_cell_6t_3 inst_cell_16_56 ( BL56, BLN56, WL16);
sram_cell_6t_3 inst_cell_16_55 ( BL55, BLN55, WL16);
sram_cell_6t_3 inst_cell_16_54 ( BL54, BLN54, WL16);
sram_cell_6t_3 inst_cell_16_53 ( BL53, BLN53, WL16);
sram_cell_6t_3 inst_cell_16_52 ( BL52, BLN52, WL16);
sram_cell_6t_3 inst_cell_16_51 ( BL51, BLN51, WL16);
sram_cell_6t_3 inst_cell_16_50 ( BL50, BLN50, WL16);
sram_cell_6t_3 inst_cell_16_49 ( BL49, BLN49, WL16);
sram_cell_6t_3 inst_cell_16_48 ( BL48, BLN48, WL16);
sram_cell_6t_3 inst_cell_16_47 ( BL47, BLN47, WL16);
sram_cell_6t_3 inst_cell_16_46 ( BL46, BLN46, WL16);
sram_cell_6t_3 inst_cell_16_45 ( BL45, BLN45, WL16);
sram_cell_6t_3 inst_cell_16_44 ( BL44, BLN44, WL16);
sram_cell_6t_3 inst_cell_16_43 ( BL43, BLN43, WL16);
sram_cell_6t_3 inst_cell_16_42 ( BL42, BLN42, WL16);
sram_cell_6t_3 inst_cell_16_41 ( BL41, BLN41, WL16);
sram_cell_6t_3 inst_cell_16_40 ( BL40, BLN40, WL16);
sram_cell_6t_3 inst_cell_16_39 ( BL39, BLN39, WL16);
sram_cell_6t_3 inst_cell_16_38 ( BL38, BLN38, WL16);
sram_cell_6t_3 inst_cell_16_37 ( BL37, BLN37, WL16);
sram_cell_6t_3 inst_cell_16_36 ( BL36, BLN36, WL16);
sram_cell_6t_3 inst_cell_16_35 ( BL35, BLN35, WL16);
sram_cell_6t_3 inst_cell_16_34 ( BL34, BLN34, WL16);
sram_cell_6t_3 inst_cell_16_33 ( BL33, BLN33, WL16);
sram_cell_6t_3 inst_cell_16_32 ( BL32, BLN32, WL16);
sram_cell_6t_3 inst_cell_15_62 ( BL62, BLN62, WL15);
sram_cell_6t_3 inst_cell_15_61 ( BL61, BLN61, WL15);
sram_cell_6t_3 inst_cell_15_60 ( BL60, BLN60, WL15);
sram_cell_6t_3 inst_cell_15_59 ( BL59, BLN59, WL15);
sram_cell_6t_3 inst_cell_15_58 ( BL58, BLN58, WL15);
sram_cell_6t_3 inst_cell_15_57 ( BL57, BLN57, WL15);
sram_cell_6t_3 inst_cell_15_56 ( BL56, BLN56, WL15);
sram_cell_6t_3 inst_cell_15_55 ( BL55, BLN55, WL15);
sram_cell_6t_3 inst_cell_15_54 ( BL54, BLN54, WL15);
sram_cell_6t_3 inst_cell_15_53 ( BL53, BLN53, WL15);
sram_cell_6t_3 inst_cell_15_52 ( BL52, BLN52, WL15);
sram_cell_6t_3 inst_cell_15_51 ( BL51, BLN51, WL15);
sram_cell_6t_3 inst_cell_15_50 ( BL50, BLN50, WL15);
sram_cell_6t_3 inst_cell_15_49 ( BL49, BLN49, WL15);
sram_cell_6t_3 inst_cell_15_48 ( BL48, BLN48, WL15);
sram_cell_6t_3 inst_cell_15_47 ( BL47, BLN47, WL15);
sram_cell_6t_3 inst_cell_15_46 ( BL46, BLN46, WL15);
sram_cell_6t_3 inst_cell_15_45 ( BL45, BLN45, WL15);
sram_cell_6t_3 inst_cell_15_44 ( BL44, BLN44, WL15);
sram_cell_6t_3 inst_cell_15_43 ( BL43, BLN43, WL15);
sram_cell_6t_3 inst_cell_15_42 ( BL42, BLN42, WL15);
sram_cell_6t_3 inst_cell_15_41 ( BL41, BLN41, WL15);
sram_cell_6t_3 inst_cell_15_40 ( BL40, BLN40, WL15);
sram_cell_6t_3 inst_cell_15_39 ( BL39, BLN39, WL15);
sram_cell_6t_3 inst_cell_15_38 ( BL38, BLN38, WL15);
sram_cell_6t_3 inst_cell_15_37 ( BL37, BLN37, WL15);
sram_cell_6t_3 inst_cell_15_36 ( BL36, BLN36, WL15);
sram_cell_6t_3 inst_cell_15_35 ( BL35, BLN35, WL15);
sram_cell_6t_3 inst_cell_15_34 ( BL34, BLN34, WL15);
sram_cell_6t_3 inst_cell_15_33 ( BL33, BLN33, WL15);
sram_cell_6t_3 inst_cell_15_32 ( BL32, BLN32, WL15);
sram_cell_6t_3 inst_cell_14_62 ( BL62, BLN62, WL14);
sram_cell_6t_3 inst_cell_14_61 ( BL61, BLN61, WL14);
sram_cell_6t_3 inst_cell_14_60 ( BL60, BLN60, WL14);
sram_cell_6t_3 inst_cell_14_59 ( BL59, BLN59, WL14);
sram_cell_6t_3 inst_cell_14_58 ( BL58, BLN58, WL14);
sram_cell_6t_3 inst_cell_14_57 ( BL57, BLN57, WL14);
sram_cell_6t_3 inst_cell_14_56 ( BL56, BLN56, WL14);
sram_cell_6t_3 inst_cell_14_55 ( BL55, BLN55, WL14);
sram_cell_6t_3 inst_cell_14_54 ( BL54, BLN54, WL14);
sram_cell_6t_3 inst_cell_14_53 ( BL53, BLN53, WL14);
sram_cell_6t_3 inst_cell_14_52 ( BL52, BLN52, WL14);
sram_cell_6t_3 inst_cell_14_51 ( BL51, BLN51, WL14);
sram_cell_6t_3 inst_cell_14_50 ( BL50, BLN50, WL14);
sram_cell_6t_3 inst_cell_14_49 ( BL49, BLN49, WL14);
sram_cell_6t_3 inst_cell_14_48 ( BL48, BLN48, WL14);
sram_cell_6t_3 inst_cell_14_47 ( BL47, BLN47, WL14);
sram_cell_6t_3 inst_cell_14_46 ( BL46, BLN46, WL14);
sram_cell_6t_3 inst_cell_14_45 ( BL45, BLN45, WL14);
sram_cell_6t_3 inst_cell_14_44 ( BL44, BLN44, WL14);
sram_cell_6t_3 inst_cell_14_43 ( BL43, BLN43, WL14);
sram_cell_6t_3 inst_cell_14_42 ( BL42, BLN42, WL14);
sram_cell_6t_3 inst_cell_14_41 ( BL41, BLN41, WL14);
sram_cell_6t_3 inst_cell_14_40 ( BL40, BLN40, WL14);
sram_cell_6t_3 inst_cell_14_39 ( BL39, BLN39, WL14);
sram_cell_6t_3 inst_cell_14_38 ( BL38, BLN38, WL14);
sram_cell_6t_3 inst_cell_14_37 ( BL37, BLN37, WL14);
sram_cell_6t_3 inst_cell_14_36 ( BL36, BLN36, WL14);
sram_cell_6t_3 inst_cell_14_35 ( BL35, BLN35, WL14);
sram_cell_6t_3 inst_cell_14_34 ( BL34, BLN34, WL14);
sram_cell_6t_3 inst_cell_14_33 ( BL33, BLN33, WL14);
sram_cell_6t_3 inst_cell_14_32 ( BL32, BLN32, WL14);
sram_cell_6t_3 inst_cell_14_31 ( BL31, BLN31, WL14);
sram_cell_6t_3 inst_cell_14_30 ( BL30, BLN30, WL14);
sram_cell_6t_3 inst_cell_14_29 ( BL29, BLN29, WL14);
sram_cell_6t_3 inst_cell_14_28 ( BL28, BLN28, WL14);
sram_cell_6t_3 inst_cell_14_27 ( BL27, BLN27, WL14);
sram_cell_6t_3 inst_cell_14_26 ( BL26, BLN26, WL14);
sram_cell_6t_3 inst_cell_14_25 ( BL25, BLN25, WL14);
sram_cell_6t_3 inst_cell_14_24 ( BL24, BLN24, WL14);
sram_cell_6t_3 inst_cell_14_23 ( BL23, BLN23, WL14);
sram_cell_6t_3 inst_cell_14_22 ( BL22, BLN22, WL14);
sram_cell_6t_3 inst_cell_14_21 ( BL21, BLN21, WL14);
sram_cell_6t_3 inst_cell_14_20 ( BL20, BLN20, WL14);
sram_cell_6t_3 inst_cell_14_19 ( BL19, BLN19, WL14);
sram_cell_6t_3 inst_cell_14_18 ( BL18, BLN18, WL14);
sram_cell_6t_3 inst_cell_14_17 ( BL17, BLN17, WL14);
sram_cell_6t_3 inst_cell_14_16 ( BL16, BLN16, WL14);
sram_cell_6t_3 inst_cell_14_15 ( BL15, BLN15, WL14);
sram_cell_6t_3 inst_cell_14_14 ( BL14, BLN14, WL14);
sram_cell_6t_3 inst_cell_14_13 ( BL13, BLN13, WL14);
sram_cell_6t_3 inst_cell_14_12 ( BL12, BLN12, WL14);
sram_cell_6t_3 inst_cell_14_11 ( BL11, BLN11, WL14);
sram_cell_6t_3 inst_cell_14_10 ( BL10, BLN10, WL14);
sram_cell_6t_3 inst_cell_14_9 ( BL9, BLN9, WL14);
sram_cell_6t_3 inst_cell_14_8 ( BL8, BLN8, WL14);
sram_cell_6t_3 inst_cell_14_7 ( BL7, BLN7, WL14);
sram_cell_6t_3 inst_cell_14_6 ( BL6, BLN6, WL14);
sram_cell_6t_3 inst_cell_14_5 ( BL5, BLN5, WL14);
sram_cell_6t_3 inst_cell_14_4 ( BL4, BLN4, WL14);
sram_cell_6t_3 inst_cell_14_3 ( BL3, BLN3, WL14);
sram_cell_6t_3 inst_cell_14_2 ( BL2, BLN2, WL14);
sram_cell_6t_3 inst_cell_14_1 ( BL1, BLN1, WL14);
sram_cell_6t_3 inst_cell_14_0 ( BL0, BLN0, WL14);
sram_cell_6t_3 inst_cell_13_31 ( BL31, BLN31, WL13);
sram_cell_6t_3 inst_cell_13_30 ( BL30, BLN30, WL13);
sram_cell_6t_3 inst_cell_13_29 ( BL29, BLN29, WL13);
sram_cell_6t_3 inst_cell_13_28 ( BL28, BLN28, WL13);
sram_cell_6t_3 inst_cell_13_27 ( BL27, BLN27, WL13);
sram_cell_6t_3 inst_cell_13_26 ( BL26, BLN26, WL13);
sram_cell_6t_3 inst_cell_13_25 ( BL25, BLN25, WL13);
sram_cell_6t_3 inst_cell_13_24 ( BL24, BLN24, WL13);
sram_cell_6t_3 inst_cell_13_23 ( BL23, BLN23, WL13);
sram_cell_6t_3 inst_cell_13_22 ( BL22, BLN22, WL13);
sram_cell_6t_3 inst_cell_13_21 ( BL21, BLN21, WL13);
sram_cell_6t_3 inst_cell_13_20 ( BL20, BLN20, WL13);
sram_cell_6t_3 inst_cell_13_19 ( BL19, BLN19, WL13);
sram_cell_6t_3 inst_cell_13_18 ( BL18, BLN18, WL13);
sram_cell_6t_3 inst_cell_13_17 ( BL17, BLN17, WL13);
sram_cell_6t_3 inst_cell_13_16 ( BL16, BLN16, WL13);
sram_cell_6t_3 inst_cell_13_15 ( BL15, BLN15, WL13);
sram_cell_6t_3 inst_cell_13_14 ( BL14, BLN14, WL13);
sram_cell_6t_3 inst_cell_13_13 ( BL13, BLN13, WL13);
sram_cell_6t_3 inst_cell_13_12 ( BL12, BLN12, WL13);
sram_cell_6t_3 inst_cell_13_11 ( BL11, BLN11, WL13);
sram_cell_6t_3 inst_cell_13_10 ( BL10, BLN10, WL13);
sram_cell_6t_3 inst_cell_13_9 ( BL9, BLN9, WL13);
sram_cell_6t_3 inst_cell_13_8 ( BL8, BLN8, WL13);
sram_cell_6t_3 inst_cell_13_7 ( BL7, BLN7, WL13);
sram_cell_6t_3 inst_cell_13_6 ( BL6, BLN6, WL13);
sram_cell_6t_3 inst_cell_13_5 ( BL5, BLN5, WL13);
sram_cell_6t_3 inst_cell_13_4 ( BL4, BLN4, WL13);
sram_cell_6t_3 inst_cell_13_3 ( BL3, BLN3, WL13);
sram_cell_6t_3 inst_cell_13_2 ( BL2, BLN2, WL13);
sram_cell_6t_3 inst_cell_13_1 ( BL1, BLN1, WL13);
sram_cell_6t_3 inst_cell_13_0 ( BL0, BLN0, WL13);
sram_cell_6t_3 inst_cell_12_31 ( BL31, BLN31, WL12);
sram_cell_6t_3 inst_cell_12_30 ( BL30, BLN30, WL12);
sram_cell_6t_3 inst_cell_12_29 ( BL29, BLN29, WL12);
sram_cell_6t_3 inst_cell_12_28 ( BL28, BLN28, WL12);
sram_cell_6t_3 inst_cell_12_27 ( BL27, BLN27, WL12);
sram_cell_6t_3 inst_cell_12_26 ( BL26, BLN26, WL12);
sram_cell_6t_3 inst_cell_12_25 ( BL25, BLN25, WL12);
sram_cell_6t_3 inst_cell_12_24 ( BL24, BLN24, WL12);
sram_cell_6t_3 inst_cell_12_23 ( BL23, BLN23, WL12);
sram_cell_6t_3 inst_cell_12_22 ( BL22, BLN22, WL12);
sram_cell_6t_3 inst_cell_12_21 ( BL21, BLN21, WL12);
sram_cell_6t_3 inst_cell_12_20 ( BL20, BLN20, WL12);
sram_cell_6t_3 inst_cell_12_19 ( BL19, BLN19, WL12);
sram_cell_6t_3 inst_cell_12_18 ( BL18, BLN18, WL12);
sram_cell_6t_3 inst_cell_12_17 ( BL17, BLN17, WL12);
sram_cell_6t_3 inst_cell_12_16 ( BL16, BLN16, WL12);
sram_cell_6t_3 inst_cell_12_15 ( BL15, BLN15, WL12);
sram_cell_6t_3 inst_cell_12_14 ( BL14, BLN14, WL12);
sram_cell_6t_3 inst_cell_12_13 ( BL13, BLN13, WL12);
sram_cell_6t_3 inst_cell_12_12 ( BL12, BLN12, WL12);
sram_cell_6t_3 inst_cell_12_11 ( BL11, BLN11, WL12);
sram_cell_6t_3 inst_cell_12_10 ( BL10, BLN10, WL12);
sram_cell_6t_3 inst_cell_12_9 ( BL9, BLN9, WL12);
sram_cell_6t_3 inst_cell_12_8 ( BL8, BLN8, WL12);
sram_cell_6t_3 inst_cell_12_7 ( BL7, BLN7, WL12);
sram_cell_6t_3 inst_cell_12_6 ( BL6, BLN6, WL12);
sram_cell_6t_3 inst_cell_12_5 ( BL5, BLN5, WL12);
sram_cell_6t_3 inst_cell_12_4 ( BL4, BLN4, WL12);
sram_cell_6t_3 inst_cell_12_3 ( BL3, BLN3, WL12);
sram_cell_6t_3 inst_cell_12_2 ( BL2, BLN2, WL12);
sram_cell_6t_3 inst_cell_12_1 ( BL1, BLN1, WL12);
sram_cell_6t_3 inst_cell_12_0 ( BL0, BLN0, WL12);
sram_cell_6t_3 inst_cell_11_31 ( BL31, BLN31, WL11);
sram_cell_6t_3 inst_cell_11_30 ( BL30, BLN30, WL11);
sram_cell_6t_3 inst_cell_11_29 ( BL29, BLN29, WL11);
sram_cell_6t_3 inst_cell_11_28 ( BL28, BLN28, WL11);
sram_cell_6t_3 inst_cell_11_27 ( BL27, BLN27, WL11);
sram_cell_6t_3 inst_cell_11_26 ( BL26, BLN26, WL11);
sram_cell_6t_3 inst_cell_11_25 ( BL25, BLN25, WL11);
sram_cell_6t_3 inst_cell_11_24 ( BL24, BLN24, WL11);
sram_cell_6t_3 inst_cell_11_23 ( BL23, BLN23, WL11);
sram_cell_6t_3 inst_cell_11_22 ( BL22, BLN22, WL11);
sram_cell_6t_3 inst_cell_11_21 ( BL21, BLN21, WL11);
sram_cell_6t_3 inst_cell_11_20 ( BL20, BLN20, WL11);
sram_cell_6t_3 inst_cell_11_19 ( BL19, BLN19, WL11);
sram_cell_6t_3 inst_cell_11_18 ( BL18, BLN18, WL11);
sram_cell_6t_3 inst_cell_11_17 ( BL17, BLN17, WL11);
sram_cell_6t_3 inst_cell_11_16 ( BL16, BLN16, WL11);
sram_cell_6t_3 inst_cell_11_15 ( BL15, BLN15, WL11);
sram_cell_6t_3 inst_cell_11_14 ( BL14, BLN14, WL11);
sram_cell_6t_3 inst_cell_11_13 ( BL13, BLN13, WL11);
sram_cell_6t_3 inst_cell_11_12 ( BL12, BLN12, WL11);
sram_cell_6t_3 inst_cell_11_11 ( BL11, BLN11, WL11);
sram_cell_6t_3 inst_cell_11_10 ( BL10, BLN10, WL11);
sram_cell_6t_3 inst_cell_11_9 ( BL9, BLN9, WL11);
sram_cell_6t_3 inst_cell_11_8 ( BL8, BLN8, WL11);
sram_cell_6t_3 inst_cell_11_7 ( BL7, BLN7, WL11);
sram_cell_6t_3 inst_cell_11_6 ( BL6, BLN6, WL11);
sram_cell_6t_3 inst_cell_11_5 ( BL5, BLN5, WL11);
sram_cell_6t_3 inst_cell_11_4 ( BL4, BLN4, WL11);
sram_cell_6t_3 inst_cell_11_3 ( BL3, BLN3, WL11);
sram_cell_6t_3 inst_cell_11_2 ( BL2, BLN2, WL11);
sram_cell_6t_3 inst_cell_11_1 ( BL1, BLN1, WL11);
sram_cell_6t_3 inst_cell_11_0 ( BL0, BLN0, WL11);
sram_cell_6t_3 inst_cell_10_31 ( BL31, BLN31, WL10);
sram_cell_6t_3 inst_cell_10_30 ( BL30, BLN30, WL10);
sram_cell_6t_3 inst_cell_10_29 ( BL29, BLN29, WL10);
sram_cell_6t_3 inst_cell_10_28 ( BL28, BLN28, WL10);
sram_cell_6t_3 inst_cell_10_27 ( BL27, BLN27, WL10);
sram_cell_6t_3 inst_cell_10_26 ( BL26, BLN26, WL10);
sram_cell_6t_3 inst_cell_10_25 ( BL25, BLN25, WL10);
sram_cell_6t_3 inst_cell_10_24 ( BL24, BLN24, WL10);
sram_cell_6t_3 inst_cell_10_23 ( BL23, BLN23, WL10);
sram_cell_6t_3 inst_cell_10_22 ( BL22, BLN22, WL10);
sram_cell_6t_3 inst_cell_10_21 ( BL21, BLN21, WL10);
sram_cell_6t_3 inst_cell_10_20 ( BL20, BLN20, WL10);
sram_cell_6t_3 inst_cell_10_19 ( BL19, BLN19, WL10);
sram_cell_6t_3 inst_cell_10_18 ( BL18, BLN18, WL10);
sram_cell_6t_3 inst_cell_10_17 ( BL17, BLN17, WL10);
sram_cell_6t_3 inst_cell_10_16 ( BL16, BLN16, WL10);
sram_cell_6t_3 inst_cell_10_15 ( BL15, BLN15, WL10);
sram_cell_6t_3 inst_cell_10_14 ( BL14, BLN14, WL10);
sram_cell_6t_3 inst_cell_10_13 ( BL13, BLN13, WL10);
sram_cell_6t_3 inst_cell_10_12 ( BL12, BLN12, WL10);
sram_cell_6t_3 inst_cell_10_11 ( BL11, BLN11, WL10);
sram_cell_6t_3 inst_cell_10_10 ( BL10, BLN10, WL10);
sram_cell_6t_3 inst_cell_10_9 ( BL9, BLN9, WL10);
sram_cell_6t_3 inst_cell_10_8 ( BL8, BLN8, WL10);
sram_cell_6t_3 inst_cell_10_7 ( BL7, BLN7, WL10);
sram_cell_6t_3 inst_cell_10_6 ( BL6, BLN6, WL10);
sram_cell_6t_3 inst_cell_10_5 ( BL5, BLN5, WL10);
sram_cell_6t_3 inst_cell_10_4 ( BL4, BLN4, WL10);
sram_cell_6t_3 inst_cell_10_3 ( BL3, BLN3, WL10);
sram_cell_6t_3 inst_cell_10_2 ( BL2, BLN2, WL10);
sram_cell_6t_3 inst_cell_10_1 ( BL1, BLN1, WL10);
sram_cell_6t_3 inst_cell_10_0 ( BL0, BLN0, WL10);
sram_cell_6t_3 inst_cell_9_31 ( BL31, BLN31, WL9);
sram_cell_6t_3 inst_cell_9_30 ( BL30, BLN30, WL9);
sram_cell_6t_3 inst_cell_9_29 ( BL29, BLN29, WL9);
sram_cell_6t_3 inst_cell_9_28 ( BL28, BLN28, WL9);
sram_cell_6t_3 inst_cell_9_27 ( BL27, BLN27, WL9);
sram_cell_6t_3 inst_cell_9_26 ( BL26, BLN26, WL9);
sram_cell_6t_3 inst_cell_9_25 ( BL25, BLN25, WL9);
sram_cell_6t_3 inst_cell_9_24 ( BL24, BLN24, WL9);
sram_cell_6t_3 inst_cell_9_23 ( BL23, BLN23, WL9);
sram_cell_6t_3 inst_cell_9_22 ( BL22, BLN22, WL9);
sram_cell_6t_3 inst_cell_9_21 ( BL21, BLN21, WL9);
sram_cell_6t_3 inst_cell_9_20 ( BL20, BLN20, WL9);
sram_cell_6t_3 inst_cell_9_19 ( BL19, BLN19, WL9);
sram_cell_6t_3 inst_cell_9_18 ( BL18, BLN18, WL9);
sram_cell_6t_3 inst_cell_9_17 ( BL17, BLN17, WL9);
sram_cell_6t_3 inst_cell_9_16 ( BL16, BLN16, WL9);
sram_cell_6t_3 inst_cell_9_15 ( BL15, BLN15, WL9);
sram_cell_6t_3 inst_cell_9_14 ( BL14, BLN14, WL9);
sram_cell_6t_3 inst_cell_9_13 ( BL13, BLN13, WL9);
sram_cell_6t_3 inst_cell_9_12 ( BL12, BLN12, WL9);
sram_cell_6t_3 inst_cell_9_11 ( BL11, BLN11, WL9);
sram_cell_6t_3 inst_cell_9_10 ( BL10, BLN10, WL9);
sram_cell_6t_3 inst_cell_9_9 ( BL9, BLN9, WL9);
sram_cell_6t_3 inst_cell_9_8 ( BL8, BLN8, WL9);
sram_cell_6t_3 inst_cell_9_7 ( BL7, BLN7, WL9);
sram_cell_6t_3 inst_cell_9_6 ( BL6, BLN6, WL9);
sram_cell_6t_3 inst_cell_9_5 ( BL5, BLN5, WL9);
sram_cell_6t_3 inst_cell_9_4 ( BL4, BLN4, WL9);
sram_cell_6t_3 inst_cell_9_3 ( BL3, BLN3, WL9);
sram_cell_6t_3 inst_cell_9_2 ( BL2, BLN2, WL9);
sram_cell_6t_3 inst_cell_9_1 ( BL1, BLN1, WL9);
sram_cell_6t_3 inst_cell_9_0 ( BL0, BLN0, WL9);
sram_cell_6t_3 inst_cell_8_31 ( BL31, BLN31, WL8);
sram_cell_6t_3 inst_cell_8_30 ( BL30, BLN30, WL8);
sram_cell_6t_3 inst_cell_8_29 ( BL29, BLN29, WL8);
sram_cell_6t_3 inst_cell_8_28 ( BL28, BLN28, WL8);
sram_cell_6t_3 inst_cell_8_27 ( BL27, BLN27, WL8);
sram_cell_6t_3 inst_cell_8_26 ( BL26, BLN26, WL8);
sram_cell_6t_3 inst_cell_8_25 ( BL25, BLN25, WL8);
sram_cell_6t_3 inst_cell_8_24 ( BL24, BLN24, WL8);
sram_cell_6t_3 inst_cell_8_23 ( BL23, BLN23, WL8);
sram_cell_6t_3 inst_cell_8_22 ( BL22, BLN22, WL8);
sram_cell_6t_3 inst_cell_8_21 ( BL21, BLN21, WL8);
sram_cell_6t_3 inst_cell_8_20 ( BL20, BLN20, WL8);
sram_cell_6t_3 inst_cell_8_19 ( BL19, BLN19, WL8);
sram_cell_6t_3 inst_cell_8_18 ( BL18, BLN18, WL8);
sram_cell_6t_3 inst_cell_8_17 ( BL17, BLN17, WL8);
sram_cell_6t_3 inst_cell_8_16 ( BL16, BLN16, WL8);
sram_cell_6t_3 inst_cell_8_15 ( BL15, BLN15, WL8);
sram_cell_6t_3 inst_cell_8_14 ( BL14, BLN14, WL8);
sram_cell_6t_3 inst_cell_8_13 ( BL13, BLN13, WL8);
sram_cell_6t_3 inst_cell_8_12 ( BL12, BLN12, WL8);
sram_cell_6t_3 inst_cell_8_11 ( BL11, BLN11, WL8);
sram_cell_6t_3 inst_cell_8_10 ( BL10, BLN10, WL8);
sram_cell_6t_3 inst_cell_8_9 ( BL9, BLN9, WL8);
sram_cell_6t_3 inst_cell_8_8 ( BL8, BLN8, WL8);
sram_cell_6t_3 inst_cell_8_7 ( BL7, BLN7, WL8);
sram_cell_6t_3 inst_cell_8_6 ( BL6, BLN6, WL8);
sram_cell_6t_3 inst_cell_8_5 ( BL5, BLN5, WL8);
sram_cell_6t_3 inst_cell_8_4 ( BL4, BLN4, WL8);
sram_cell_6t_3 inst_cell_8_3 ( BL3, BLN3, WL8);
sram_cell_6t_3 inst_cell_8_2 ( BL2, BLN2, WL8);
sram_cell_6t_3 inst_cell_8_1 ( BL1, BLN1, WL8);
sram_cell_6t_3 inst_cell_8_0 ( BL0, BLN0, WL8);
sram_cell_6t_3 inst_cell_7_31 ( BL31, BLN31, WL7);
sram_cell_6t_3 inst_cell_7_30 ( BL30, BLN30, WL7);
sram_cell_6t_3 inst_cell_7_29 ( BL29, BLN29, WL7);
sram_cell_6t_3 inst_cell_7_28 ( BL28, BLN28, WL7);
sram_cell_6t_3 inst_cell_7_27 ( BL27, BLN27, WL7);
sram_cell_6t_3 inst_cell_7_26 ( BL26, BLN26, WL7);
sram_cell_6t_3 inst_cell_7_25 ( BL25, BLN25, WL7);
sram_cell_6t_3 inst_cell_7_24 ( BL24, BLN24, WL7);
sram_cell_6t_3 inst_cell_7_23 ( BL23, BLN23, WL7);
sram_cell_6t_3 inst_cell_7_22 ( BL22, BLN22, WL7);
sram_cell_6t_3 inst_cell_7_21 ( BL21, BLN21, WL7);
sram_cell_6t_3 inst_cell_7_20 ( BL20, BLN20, WL7);
sram_cell_6t_3 inst_cell_7_19 ( BL19, BLN19, WL7);
sram_cell_6t_3 inst_cell_7_18 ( BL18, BLN18, WL7);
sram_cell_6t_3 inst_cell_7_17 ( BL17, BLN17, WL7);
sram_cell_6t_3 inst_cell_7_16 ( BL16, BLN16, WL7);
sram_cell_6t_3 inst_cell_7_15 ( BL15, BLN15, WL7);
sram_cell_6t_3 inst_cell_7_14 ( BL14, BLN14, WL7);
sram_cell_6t_3 inst_cell_7_13 ( BL13, BLN13, WL7);
sram_cell_6t_3 inst_cell_7_12 ( BL12, BLN12, WL7);
sram_cell_6t_3 inst_cell_7_11 ( BL11, BLN11, WL7);
sram_cell_6t_3 inst_cell_7_10 ( BL10, BLN10, WL7);
sram_cell_6t_3 inst_cell_7_9 ( BL9, BLN9, WL7);
sram_cell_6t_3 inst_cell_7_8 ( BL8, BLN8, WL7);
sram_cell_6t_3 inst_cell_7_7 ( BL7, BLN7, WL7);
sram_cell_6t_3 inst_cell_7_6 ( BL6, BLN6, WL7);
sram_cell_6t_3 inst_cell_7_5 ( BL5, BLN5, WL7);
sram_cell_6t_3 inst_cell_7_4 ( BL4, BLN4, WL7);
sram_cell_6t_3 inst_cell_7_3 ( BL3, BLN3, WL7);
sram_cell_6t_3 inst_cell_7_2 ( BL2, BLN2, WL7);
sram_cell_6t_3 inst_cell_7_1 ( BL1, BLN1, WL7);
sram_cell_6t_3 inst_cell_7_0 ( BL0, BLN0, WL7);
sram_cell_6t_3 inst_cell_6_31 ( BL31, BLN31, WL6);
sram_cell_6t_3 inst_cell_6_30 ( BL30, BLN30, WL6);
sram_cell_6t_3 inst_cell_6_29 ( BL29, BLN29, WL6);
sram_cell_6t_3 inst_cell_6_28 ( BL28, BLN28, WL6);
sram_cell_6t_3 inst_cell_6_27 ( BL27, BLN27, WL6);
sram_cell_6t_3 inst_cell_6_26 ( BL26, BLN26, WL6);
sram_cell_6t_3 inst_cell_6_25 ( BL25, BLN25, WL6);
sram_cell_6t_3 inst_cell_6_24 ( BL24, BLN24, WL6);
sram_cell_6t_3 inst_cell_6_23 ( BL23, BLN23, WL6);
sram_cell_6t_3 inst_cell_6_22 ( BL22, BLN22, WL6);
sram_cell_6t_3 inst_cell_6_21 ( BL21, BLN21, WL6);
sram_cell_6t_3 inst_cell_6_20 ( BL20, BLN20, WL6);
sram_cell_6t_3 inst_cell_6_19 ( BL19, BLN19, WL6);
sram_cell_6t_3 inst_cell_6_18 ( BL18, BLN18, WL6);
sram_cell_6t_3 inst_cell_6_17 ( BL17, BLN17, WL6);
sram_cell_6t_3 inst_cell_6_16 ( BL16, BLN16, WL6);
sram_cell_6t_3 inst_cell_6_15 ( BL15, BLN15, WL6);
sram_cell_6t_3 inst_cell_6_14 ( BL14, BLN14, WL6);
sram_cell_6t_3 inst_cell_6_13 ( BL13, BLN13, WL6);
sram_cell_6t_3 inst_cell_6_12 ( BL12, BLN12, WL6);
sram_cell_6t_3 inst_cell_6_11 ( BL11, BLN11, WL6);
sram_cell_6t_3 inst_cell_6_10 ( BL10, BLN10, WL6);
sram_cell_6t_3 inst_cell_6_9 ( BL9, BLN9, WL6);
sram_cell_6t_3 inst_cell_6_8 ( BL8, BLN8, WL6);
sram_cell_6t_3 inst_cell_6_7 ( BL7, BLN7, WL6);
sram_cell_6t_3 inst_cell_6_6 ( BL6, BLN6, WL6);
sram_cell_6t_3 inst_cell_6_5 ( BL5, BLN5, WL6);
sram_cell_6t_3 inst_cell_6_4 ( BL4, BLN4, WL6);
sram_cell_6t_3 inst_cell_6_3 ( BL3, BLN3, WL6);
sram_cell_6t_3 inst_cell_6_2 ( BL2, BLN2, WL6);
sram_cell_6t_3 inst_cell_6_1 ( BL1, BLN1, WL6);
sram_cell_6t_3 inst_cell_6_0 ( BL0, BLN0, WL6);
sram_cell_6t_3 inst_cell_5_31 ( BL31, BLN31, WL5);
sram_cell_6t_3 inst_cell_5_30 ( BL30, BLN30, WL5);
sram_cell_6t_3 inst_cell_5_29 ( BL29, BLN29, WL5);
sram_cell_6t_3 inst_cell_5_28 ( BL28, BLN28, WL5);
sram_cell_6t_3 inst_cell_5_27 ( BL27, BLN27, WL5);
sram_cell_6t_3 inst_cell_5_26 ( BL26, BLN26, WL5);
sram_cell_6t_3 inst_cell_5_25 ( BL25, BLN25, WL5);
sram_cell_6t_3 inst_cell_5_24 ( BL24, BLN24, WL5);
sram_cell_6t_3 inst_cell_5_23 ( BL23, BLN23, WL5);
sram_cell_6t_3 inst_cell_5_22 ( BL22, BLN22, WL5);
sram_cell_6t_3 inst_cell_5_21 ( BL21, BLN21, WL5);
sram_cell_6t_3 inst_cell_5_20 ( BL20, BLN20, WL5);
sram_cell_6t_3 inst_cell_5_19 ( BL19, BLN19, WL5);
sram_cell_6t_3 inst_cell_5_18 ( BL18, BLN18, WL5);
sram_cell_6t_3 inst_cell_5_17 ( BL17, BLN17, WL5);
sram_cell_6t_3 inst_cell_5_16 ( BL16, BLN16, WL5);
sram_cell_6t_3 inst_cell_5_15 ( BL15, BLN15, WL5);
sram_cell_6t_3 inst_cell_5_14 ( BL14, BLN14, WL5);
sram_cell_6t_3 inst_cell_5_13 ( BL13, BLN13, WL5);
sram_cell_6t_3 inst_cell_5_12 ( BL12, BLN12, WL5);
sram_cell_6t_3 inst_cell_5_11 ( BL11, BLN11, WL5);
sram_cell_6t_3 inst_cell_5_10 ( BL10, BLN10, WL5);
sram_cell_6t_3 inst_cell_5_9 ( BL9, BLN9, WL5);
sram_cell_6t_3 inst_cell_5_8 ( BL8, BLN8, WL5);
sram_cell_6t_3 inst_cell_5_7 ( BL7, BLN7, WL5);
sram_cell_6t_3 inst_cell_5_6 ( BL6, BLN6, WL5);
sram_cell_6t_3 inst_cell_5_5 ( BL5, BLN5, WL5);
sram_cell_6t_3 inst_cell_5_4 ( BL4, BLN4, WL5);
sram_cell_6t_3 inst_cell_5_3 ( BL3, BLN3, WL5);
sram_cell_6t_3 inst_cell_5_2 ( BL2, BLN2, WL5);
sram_cell_6t_3 inst_cell_5_1 ( BL1, BLN1, WL5);
sram_cell_6t_3 inst_cell_5_0 ( BL0, BLN0, WL5);
sram_cell_6t_3 inst_cell_4_31 ( BL31, BLN31, WL4);
sram_cell_6t_3 inst_cell_4_30 ( BL30, BLN30, WL4);
sram_cell_6t_3 inst_cell_4_29 ( BL29, BLN29, WL4);
sram_cell_6t_3 inst_cell_4_28 ( BL28, BLN28, WL4);
sram_cell_6t_3 inst_cell_4_27 ( BL27, BLN27, WL4);
sram_cell_6t_3 inst_cell_4_26 ( BL26, BLN26, WL4);
sram_cell_6t_3 inst_cell_4_25 ( BL25, BLN25, WL4);
sram_cell_6t_3 inst_cell_4_24 ( BL24, BLN24, WL4);
sram_cell_6t_3 inst_cell_4_23 ( BL23, BLN23, WL4);
sram_cell_6t_3 inst_cell_4_22 ( BL22, BLN22, WL4);
sram_cell_6t_3 inst_cell_4_21 ( BL21, BLN21, WL4);
sram_cell_6t_3 inst_cell_4_20 ( BL20, BLN20, WL4);
sram_cell_6t_3 inst_cell_4_19 ( BL19, BLN19, WL4);
sram_cell_6t_3 inst_cell_4_18 ( BL18, BLN18, WL4);
sram_cell_6t_3 inst_cell_4_17 ( BL17, BLN17, WL4);
sram_cell_6t_3 inst_cell_4_16 ( BL16, BLN16, WL4);
sram_cell_6t_3 inst_cell_4_15 ( BL15, BLN15, WL4);
sram_cell_6t_3 inst_cell_4_14 ( BL14, BLN14, WL4);
sram_cell_6t_3 inst_cell_4_13 ( BL13, BLN13, WL4);
sram_cell_6t_3 inst_cell_4_12 ( BL12, BLN12, WL4);
sram_cell_6t_3 inst_cell_4_11 ( BL11, BLN11, WL4);
sram_cell_6t_3 inst_cell_4_10 ( BL10, BLN10, WL4);
sram_cell_6t_3 inst_cell_4_9 ( BL9, BLN9, WL4);
sram_cell_6t_3 inst_cell_4_8 ( BL8, BLN8, WL4);
sram_cell_6t_3 inst_cell_4_7 ( BL7, BLN7, WL4);
sram_cell_6t_3 inst_cell_4_6 ( BL6, BLN6, WL4);
sram_cell_6t_3 inst_cell_4_5 ( BL5, BLN5, WL4);
sram_cell_6t_3 inst_cell_4_4 ( BL4, BLN4, WL4);
sram_cell_6t_3 inst_cell_4_3 ( BL3, BLN3, WL4);
sram_cell_6t_3 inst_cell_4_2 ( BL2, BLN2, WL4);
sram_cell_6t_3 inst_cell_4_1 ( BL1, BLN1, WL4);
sram_cell_6t_3 inst_cell_4_0 ( BL0, BLN0, WL4);
sram_cell_6t_3 inst_cell_3_31 ( BL31, BLN31, WL3);
sram_cell_6t_3 inst_cell_3_30 ( BL30, BLN30, WL3);
sram_cell_6t_3 inst_cell_3_29 ( BL29, BLN29, WL3);
sram_cell_6t_3 inst_cell_3_28 ( BL28, BLN28, WL3);
sram_cell_6t_3 inst_cell_3_27 ( BL27, BLN27, WL3);
sram_cell_6t_3 inst_cell_3_26 ( BL26, BLN26, WL3);
sram_cell_6t_3 inst_cell_3_25 ( BL25, BLN25, WL3);
sram_cell_6t_3 inst_cell_3_24 ( BL24, BLN24, WL3);
sram_cell_6t_3 inst_cell_3_23 ( BL23, BLN23, WL3);
sram_cell_6t_3 inst_cell_3_22 ( BL22, BLN22, WL3);
sram_cell_6t_3 inst_cell_3_21 ( BL21, BLN21, WL3);
sram_cell_6t_3 inst_cell_3_20 ( BL20, BLN20, WL3);
sram_cell_6t_3 inst_cell_3_19 ( BL19, BLN19, WL3);
sram_cell_6t_3 inst_cell_3_18 ( BL18, BLN18, WL3);
sram_cell_6t_3 inst_cell_3_17 ( BL17, BLN17, WL3);
sram_cell_6t_3 inst_cell_3_16 ( BL16, BLN16, WL3);
sram_cell_6t_3 inst_cell_3_15 ( BL15, BLN15, WL3);
sram_cell_6t_3 inst_cell_3_14 ( BL14, BLN14, WL3);
sram_cell_6t_3 inst_cell_3_13 ( BL13, BLN13, WL3);
sram_cell_6t_3 inst_cell_3_12 ( BL12, BLN12, WL3);
sram_cell_6t_3 inst_cell_3_11 ( BL11, BLN11, WL3);
sram_cell_6t_3 inst_cell_3_10 ( BL10, BLN10, WL3);
sram_cell_6t_3 inst_cell_3_9 ( BL9, BLN9, WL3);
sram_cell_6t_3 inst_cell_3_8 ( BL8, BLN8, WL3);
sram_cell_6t_3 inst_cell_3_7 ( BL7, BLN7, WL3);
sram_cell_6t_3 inst_cell_3_6 ( BL6, BLN6, WL3);
sram_cell_6t_3 inst_cell_3_5 ( BL5, BLN5, WL3);
sram_cell_6t_3 inst_cell_3_4 ( BL4, BLN4, WL3);
sram_cell_6t_3 inst_cell_3_3 ( BL3, BLN3, WL3);
sram_cell_6t_3 inst_cell_3_2 ( BL2, BLN2, WL3);
sram_cell_6t_3 inst_cell_3_1 ( BL1, BLN1, WL3);
sram_cell_6t_3 inst_cell_3_0 ( BL0, BLN0, WL3);
sram_cell_6t_3 inst_cell_2_31 ( BL31, BLN31, WL2);
sram_cell_6t_3 inst_cell_2_30 ( BL30, BLN30, WL2);
sram_cell_6t_3 inst_cell_2_29 ( BL29, BLN29, WL2);
sram_cell_6t_3 inst_cell_2_28 ( BL28, BLN28, WL2);
sram_cell_6t_3 inst_cell_2_27 ( BL27, BLN27, WL2);
sram_cell_6t_3 inst_cell_2_26 ( BL26, BLN26, WL2);
sram_cell_6t_3 inst_cell_2_25 ( BL25, BLN25, WL2);
sram_cell_6t_3 inst_cell_2_24 ( BL24, BLN24, WL2);
sram_cell_6t_3 inst_cell_2_23 ( BL23, BLN23, WL2);
sram_cell_6t_3 inst_cell_2_22 ( BL22, BLN22, WL2);
sram_cell_6t_3 inst_cell_2_21 ( BL21, BLN21, WL2);
sram_cell_6t_3 inst_cell_2_20 ( BL20, BLN20, WL2);
sram_cell_6t_3 inst_cell_2_19 ( BL19, BLN19, WL2);
sram_cell_6t_3 inst_cell_2_18 ( BL18, BLN18, WL2);
sram_cell_6t_3 inst_cell_2_17 ( BL17, BLN17, WL2);
sram_cell_6t_3 inst_cell_2_16 ( BL16, BLN16, WL2);
sram_cell_6t_3 inst_cell_2_15 ( BL15, BLN15, WL2);
sram_cell_6t_3 inst_cell_2_14 ( BL14, BLN14, WL2);
sram_cell_6t_3 inst_cell_2_13 ( BL13, BLN13, WL2);
sram_cell_6t_3 inst_cell_2_12 ( BL12, BLN12, WL2);
sram_cell_6t_3 inst_cell_2_11 ( BL11, BLN11, WL2);
sram_cell_6t_3 inst_cell_2_10 ( BL10, BLN10, WL2);
sram_cell_6t_3 inst_cell_2_9 ( BL9, BLN9, WL2);
sram_cell_6t_3 inst_cell_2_8 ( BL8, BLN8, WL2);
sram_cell_6t_3 inst_cell_2_7 ( BL7, BLN7, WL2);
sram_cell_6t_3 inst_cell_2_6 ( BL6, BLN6, WL2);
sram_cell_6t_3 inst_cell_2_5 ( BL5, BLN5, WL2);
sram_cell_6t_3 inst_cell_2_4 ( BL4, BLN4, WL2);
sram_cell_6t_3 inst_cell_2_3 ( BL3, BLN3, WL2);
sram_cell_6t_3 inst_cell_2_2 ( BL2, BLN2, WL2);
sram_cell_6t_3 inst_cell_2_1 ( BL1, BLN1, WL2);
sram_cell_6t_3 inst_cell_2_0 ( BL0, BLN0, WL2);
sram_cell_6t_3 inst_cell_1_31 ( BL31, BLN31, WL1);
sram_cell_6t_3 inst_cell_0_31 ( BL31, BLN31, WL0);
sram_cell_6t_3 inst_cell_1_30 ( BL30, BLN30, WL1);
sram_cell_6t_3 inst_cell_0_30 ( BL30, BLN30, WL0);
sram_cell_6t_3 inst_cell_1_29 ( BL29, BLN29, WL1);
sram_cell_6t_3 inst_cell_0_29 ( BL29, BLN29, WL0);
sram_cell_6t_3 inst_cell_1_28 ( BL28, BLN28, WL1);
sram_cell_6t_3 inst_cell_0_28 ( BL28, BLN28, WL0);
sram_cell_6t_3 inst_cell_1_27 ( BL27, BLN27, WL1);
sram_cell_6t_3 inst_cell_0_27 ( BL27, BLN27, WL0);
sram_cell_6t_3 inst_cell_1_26 ( BL26, BLN26, WL1);
sram_cell_6t_3 inst_cell_0_26 ( BL26, BLN26, WL0);
sram_cell_6t_3 inst_cell_1_25 ( BL25, BLN25, WL1);
sram_cell_6t_3 inst_cell_0_25 ( BL25, BLN25, WL0);
sram_cell_6t_3 inst_cell_1_24 ( BL24, BLN24, WL1);
sram_cell_6t_3 inst_cell_0_24 ( BL24, BLN24, WL0);
sram_cell_6t_3 inst_cell_1_23 ( BL23, BLN23, WL1);
sram_cell_6t_3 inst_cell_0_23 ( BL23, BLN23, WL0);
sram_cell_6t_3 inst_cell_1_22 ( BL22, BLN22, WL1);
sram_cell_6t_3 inst_cell_0_22 ( BL22, BLN22, WL0);
sram_cell_6t_3 inst_cell_1_21 ( BL21, BLN21, WL1);
sram_cell_6t_3 inst_cell_0_21 ( BL21, BLN21, WL0);
sram_cell_6t_3 inst_cell_1_20 ( BL20, BLN20, WL1);
sram_cell_6t_3 inst_cell_0_20 ( BL20, BLN20, WL0);
sram_cell_6t_3 inst_cell_1_19 ( BL19, BLN19, WL1);
sram_cell_6t_3 inst_cell_0_19 ( BL19, BLN19, WL0);
sram_cell_6t_3 inst_cell_1_18 ( BL18, BLN18, WL1);
sram_cell_6t_3 inst_cell_0_18 ( BL18, BLN18, WL0);
sram_cell_6t_3 inst_cell_1_17 ( BL17, BLN17, WL1);
sram_cell_6t_3 inst_cell_0_17 ( BL17, BLN17, WL0);
sram_cell_6t_3 inst_cell_1_16 ( BL16, BLN16, WL1);
sram_cell_6t_3 inst_cell_0_16 ( BL16, BLN16, WL0);
sram_cell_6t_3 inst_cell_1_15 ( BL15, BLN15, WL1);
sram_cell_6t_3 inst_cell_0_15 ( BL15, BLN15, WL0);
sram_cell_6t_3 inst_cell_1_14 ( BL14, BLN14, WL1);
sram_cell_6t_3 inst_cell_0_14 ( BL14, BLN14, WL0);
sram_cell_6t_3 inst_cell_1_13 ( BL13, BLN13, WL1);
sram_cell_6t_3 inst_cell_0_13 ( BL13, BLN13, WL0);
sram_cell_6t_3 inst_cell_1_12 ( BL12, BLN12, WL1);
sram_cell_6t_3 inst_cell_0_12 ( BL12, BLN12, WL0);
sram_cell_6t_3 inst_cell_1_11 ( BL11, BLN11, WL1);
sram_cell_6t_3 inst_cell_0_11 ( BL11, BLN11, WL0);
sram_cell_6t_3 inst_cell_1_10 ( BL10, BLN10, WL1);
sram_cell_6t_3 inst_cell_0_10 ( BL10, BLN10, WL0);
sram_cell_6t_3 inst_cell_1_9 ( BL9, BLN9, WL1);
sram_cell_6t_3 inst_cell_0_9 ( BL9, BLN9, WL0);
sram_cell_6t_3 inst_cell_1_8 ( BL8, BLN8, WL1);
sram_cell_6t_3 inst_cell_0_8 ( BL8, BLN8, WL0);
sram_cell_6t_3 inst_cell_1_7 ( BL7, BLN7, WL1);
sram_cell_6t_3 inst_cell_0_7 ( BL7, BLN7, WL0);
sram_cell_6t_3 inst_cell_1_6 ( BL6, BLN6, WL1);
sram_cell_6t_3 inst_cell_0_6 ( BL6, BLN6, WL0);
sram_cell_6t_3 inst_cell_1_5 ( BL5, BLN5, WL1);
sram_cell_6t_3 inst_cell_0_5 ( BL5, BLN5, WL0);
sram_cell_6t_3 inst_cell_1_4 ( BL4, BLN4, WL1);
sram_cell_6t_3 inst_cell_0_4 ( BL4, BLN4, WL0);
sram_cell_6t_3 inst_cell_1_3 ( BL3, BLN3, WL1);
sram_cell_6t_3 inst_cell_0_3 ( BL3, BLN3, WL0);
sram_cell_6t_3 inst_cell_1_2 ( BL2, BLN2, WL1);
sram_cell_6t_3 inst_cell_0_2 ( BL2, BLN2, WL0);
sram_cell_6t_3 inst_cell_1_1 ( BL1, BLN1, WL1);
sram_cell_6t_3 inst_cell_0_1 ( BL1, BLN1, WL0);
sram_cell_6t_3 inst_cell_1_0 ( BL0, BLN0, WL1);
sram_cell_6t_3 inst_cell_0_0 ( BL0, BLN0, WL0);
sram_cell_6t_3 inst_cell_13_63 ( BL63, BLN63, WL13);
sram_cell_6t_3 inst_cell_12_63 ( BL63, BLN63, WL12);
sram_cell_6t_3 inst_cell_11_63 ( BL63, BLN63, WL11);
sram_cell_6t_3 inst_cell_10_63 ( BL63, BLN63, WL10);
sram_cell_6t_3 inst_cell_9_63 ( BL63, BLN63, WL9);
sram_cell_6t_3 inst_cell_8_63 ( BL63, BLN63, WL8);
sram_cell_6t_3 inst_cell_7_63 ( BL63, BLN63, WL7);
sram_cell_6t_3 inst_cell_6_63 ( BL63, BLN63, WL6);
sram_cell_6t_3 inst_cell_5_63 ( BL63, BLN63, WL5);
sram_cell_6t_3 inst_cell_4_63 ( BL63, BLN63, WL4);
sram_cell_6t_3 inst_cell_3_63 ( BL63, BLN63, WL3);
sram_cell_6t_3 inst_cell_2_63 ( BL63, BLN63, WL2);
sram_cell_6t_3 inst_cell_1_63 ( BL63, BLN63, WL1);
sram_cell_6t_3 inst_cell_0_63 ( BL63, BLN63, WL0);
sram_cell_6t_3 inst_cell_13_62 ( BL62, BLN62, WL13);
sram_cell_6t_3 inst_cell_12_62 ( BL62, BLN62, WL12);
sram_cell_6t_3 inst_cell_11_62 ( BL62, BLN62, WL11);
sram_cell_6t_3 inst_cell_10_62 ( BL62, BLN62, WL10);
sram_cell_6t_3 inst_cell_9_62 ( BL62, BLN62, WL9);
sram_cell_6t_3 inst_cell_8_62 ( BL62, BLN62, WL8);
sram_cell_6t_3 inst_cell_7_62 ( BL62, BLN62, WL7);
sram_cell_6t_3 inst_cell_6_62 ( BL62, BLN62, WL6);
sram_cell_6t_3 inst_cell_5_62 ( BL62, BLN62, WL5);
sram_cell_6t_3 inst_cell_4_62 ( BL62, BLN62, WL4);
sram_cell_6t_3 inst_cell_3_62 ( BL62, BLN62, WL3);
sram_cell_6t_3 inst_cell_2_62 ( BL62, BLN62, WL2);
sram_cell_6t_3 inst_cell_1_62 ( BL62, BLN62, WL1);
sram_cell_6t_3 inst_cell_0_62 ( BL62, BLN62, WL0);
sram_cell_6t_3 inst_cell_13_61 ( BL61, BLN61, WL13);
sram_cell_6t_3 inst_cell_12_61 ( BL61, BLN61, WL12);
sram_cell_6t_3 inst_cell_11_61 ( BL61, BLN61, WL11);
sram_cell_6t_3 inst_cell_10_61 ( BL61, BLN61, WL10);
sram_cell_6t_3 inst_cell_9_61 ( BL61, BLN61, WL9);
sram_cell_6t_3 inst_cell_8_61 ( BL61, BLN61, WL8);
sram_cell_6t_3 inst_cell_7_61 ( BL61, BLN61, WL7);
sram_cell_6t_3 inst_cell_6_61 ( BL61, BLN61, WL6);
sram_cell_6t_3 inst_cell_5_61 ( BL61, BLN61, WL5);
sram_cell_6t_3 inst_cell_4_61 ( BL61, BLN61, WL4);
sram_cell_6t_3 inst_cell_3_61 ( BL61, BLN61, WL3);
sram_cell_6t_3 inst_cell_2_61 ( BL61, BLN61, WL2);
sram_cell_6t_3 inst_cell_1_61 ( BL61, BLN61, WL1);
sram_cell_6t_3 inst_cell_0_61 ( BL61, BLN61, WL0);
sram_cell_6t_3 inst_cell_13_60 ( BL60, BLN60, WL13);
sram_cell_6t_3 inst_cell_12_60 ( BL60, BLN60, WL12);
sram_cell_6t_3 inst_cell_11_60 ( BL60, BLN60, WL11);
sram_cell_6t_3 inst_cell_10_60 ( BL60, BLN60, WL10);
sram_cell_6t_3 inst_cell_9_60 ( BL60, BLN60, WL9);
sram_cell_6t_3 inst_cell_8_60 ( BL60, BLN60, WL8);
sram_cell_6t_3 inst_cell_7_60 ( BL60, BLN60, WL7);
sram_cell_6t_3 inst_cell_6_60 ( BL60, BLN60, WL6);
sram_cell_6t_3 inst_cell_5_60 ( BL60, BLN60, WL5);
sram_cell_6t_3 inst_cell_4_60 ( BL60, BLN60, WL4);
sram_cell_6t_3 inst_cell_3_60 ( BL60, BLN60, WL3);
sram_cell_6t_3 inst_cell_2_60 ( BL60, BLN60, WL2);
sram_cell_6t_3 inst_cell_1_60 ( BL60, BLN60, WL1);
sram_cell_6t_3 inst_cell_0_60 ( BL60, BLN60, WL0);
sram_cell_6t_3 inst_cell_13_59 ( BL59, BLN59, WL13);
sram_cell_6t_3 inst_cell_12_59 ( BL59, BLN59, WL12);
sram_cell_6t_3 inst_cell_11_59 ( BL59, BLN59, WL11);
sram_cell_6t_3 inst_cell_10_59 ( BL59, BLN59, WL10);
sram_cell_6t_3 inst_cell_9_59 ( BL59, BLN59, WL9);
sram_cell_6t_3 inst_cell_8_59 ( BL59, BLN59, WL8);
sram_cell_6t_3 inst_cell_7_59 ( BL59, BLN59, WL7);
sram_cell_6t_3 inst_cell_6_59 ( BL59, BLN59, WL6);
sram_cell_6t_3 inst_cell_5_59 ( BL59, BLN59, WL5);
sram_cell_6t_3 inst_cell_4_59 ( BL59, BLN59, WL4);
sram_cell_6t_3 inst_cell_3_59 ( BL59, BLN59, WL3);
sram_cell_6t_3 inst_cell_2_59 ( BL59, BLN59, WL2);
sram_cell_6t_3 inst_cell_1_59 ( BL59, BLN59, WL1);
sram_cell_6t_3 inst_cell_0_59 ( BL59, BLN59, WL0);
sram_cell_6t_3 inst_cell_13_58 ( BL58, BLN58, WL13);
sram_cell_6t_3 inst_cell_12_58 ( BL58, BLN58, WL12);
sram_cell_6t_3 inst_cell_11_58 ( BL58, BLN58, WL11);
sram_cell_6t_3 inst_cell_10_58 ( BL58, BLN58, WL10);
sram_cell_6t_3 inst_cell_9_58 ( BL58, BLN58, WL9);
sram_cell_6t_3 inst_cell_8_58 ( BL58, BLN58, WL8);
sram_cell_6t_3 inst_cell_7_58 ( BL58, BLN58, WL7);
sram_cell_6t_3 inst_cell_6_58 ( BL58, BLN58, WL6);
sram_cell_6t_3 inst_cell_5_58 ( BL58, BLN58, WL5);
sram_cell_6t_3 inst_cell_4_58 ( BL58, BLN58, WL4);
sram_cell_6t_3 inst_cell_3_58 ( BL58, BLN58, WL3);
sram_cell_6t_3 inst_cell_2_58 ( BL58, BLN58, WL2);
sram_cell_6t_3 inst_cell_1_58 ( BL58, BLN58, WL1);
sram_cell_6t_3 inst_cell_0_58 ( BL58, BLN58, WL0);
sram_cell_6t_3 inst_cell_13_57 ( BL57, BLN57, WL13);
sram_cell_6t_3 inst_cell_12_57 ( BL57, BLN57, WL12);
sram_cell_6t_3 inst_cell_11_57 ( BL57, BLN57, WL11);
sram_cell_6t_3 inst_cell_10_57 ( BL57, BLN57, WL10);
sram_cell_6t_3 inst_cell_9_57 ( BL57, BLN57, WL9);
sram_cell_6t_3 inst_cell_8_57 ( BL57, BLN57, WL8);
sram_cell_6t_3 inst_cell_7_57 ( BL57, BLN57, WL7);
sram_cell_6t_3 inst_cell_6_57 ( BL57, BLN57, WL6);
sram_cell_6t_3 inst_cell_5_57 ( BL57, BLN57, WL5);
sram_cell_6t_3 inst_cell_4_57 ( BL57, BLN57, WL4);
sram_cell_6t_3 inst_cell_3_57 ( BL57, BLN57, WL3);
sram_cell_6t_3 inst_cell_2_57 ( BL57, BLN57, WL2);
sram_cell_6t_3 inst_cell_1_57 ( BL57, BLN57, WL1);
sram_cell_6t_3 inst_cell_0_57 ( BL57, BLN57, WL0);
sram_cell_6t_3 inst_cell_13_56 ( BL56, BLN56, WL13);
sram_cell_6t_3 inst_cell_12_56 ( BL56, BLN56, WL12);
sram_cell_6t_3 inst_cell_11_56 ( BL56, BLN56, WL11);
sram_cell_6t_3 inst_cell_10_56 ( BL56, BLN56, WL10);
sram_cell_6t_3 inst_cell_9_56 ( BL56, BLN56, WL9);
sram_cell_6t_3 inst_cell_8_56 ( BL56, BLN56, WL8);
sram_cell_6t_3 inst_cell_7_56 ( BL56, BLN56, WL7);
sram_cell_6t_3 inst_cell_6_56 ( BL56, BLN56, WL6);
sram_cell_6t_3 inst_cell_5_56 ( BL56, BLN56, WL5);
sram_cell_6t_3 inst_cell_4_56 ( BL56, BLN56, WL4);
sram_cell_6t_3 inst_cell_3_56 ( BL56, BLN56, WL3);
sram_cell_6t_3 inst_cell_2_56 ( BL56, BLN56, WL2);
sram_cell_6t_3 inst_cell_1_56 ( BL56, BLN56, WL1);
sram_cell_6t_3 inst_cell_0_56 ( BL56, BLN56, WL0);
sram_cell_6t_3 inst_cell_13_55 ( BL55, BLN55, WL13);
sram_cell_6t_3 inst_cell_12_55 ( BL55, BLN55, WL12);
sram_cell_6t_3 inst_cell_11_55 ( BL55, BLN55, WL11);
sram_cell_6t_3 inst_cell_10_55 ( BL55, BLN55, WL10);
sram_cell_6t_3 inst_cell_9_55 ( BL55, BLN55, WL9);
sram_cell_6t_3 inst_cell_8_55 ( BL55, BLN55, WL8);
sram_cell_6t_3 inst_cell_7_55 ( BL55, BLN55, WL7);
sram_cell_6t_3 inst_cell_6_55 ( BL55, BLN55, WL6);
sram_cell_6t_3 inst_cell_5_55 ( BL55, BLN55, WL5);
sram_cell_6t_3 inst_cell_4_55 ( BL55, BLN55, WL4);
sram_cell_6t_3 inst_cell_3_55 ( BL55, BLN55, WL3);
sram_cell_6t_3 inst_cell_2_55 ( BL55, BLN55, WL2);
sram_cell_6t_3 inst_cell_1_55 ( BL55, BLN55, WL1);
sram_cell_6t_3 inst_cell_0_55 ( BL55, BLN55, WL0);
sram_cell_6t_3 inst_cell_13_54 ( BL54, BLN54, WL13);
sram_cell_6t_3 inst_cell_12_54 ( BL54, BLN54, WL12);
sram_cell_6t_3 inst_cell_11_54 ( BL54, BLN54, WL11);
sram_cell_6t_3 inst_cell_10_54 ( BL54, BLN54, WL10);
sram_cell_6t_3 inst_cell_9_54 ( BL54, BLN54, WL9);
sram_cell_6t_3 inst_cell_8_54 ( BL54, BLN54, WL8);
sram_cell_6t_3 inst_cell_7_54 ( BL54, BLN54, WL7);
sram_cell_6t_3 inst_cell_6_54 ( BL54, BLN54, WL6);
sram_cell_6t_3 inst_cell_5_54 ( BL54, BLN54, WL5);
sram_cell_6t_3 inst_cell_4_54 ( BL54, BLN54, WL4);
sram_cell_6t_3 inst_cell_3_54 ( BL54, BLN54, WL3);
sram_cell_6t_3 inst_cell_2_54 ( BL54, BLN54, WL2);
sram_cell_6t_3 inst_cell_1_54 ( BL54, BLN54, WL1);
sram_cell_6t_3 inst_cell_0_54 ( BL54, BLN54, WL0);
sram_cell_6t_3 inst_cell_13_53 ( BL53, BLN53, WL13);
sram_cell_6t_3 inst_cell_12_53 ( BL53, BLN53, WL12);
sram_cell_6t_3 inst_cell_11_53 ( BL53, BLN53, WL11);
sram_cell_6t_3 inst_cell_10_53 ( BL53, BLN53, WL10);
sram_cell_6t_3 inst_cell_9_53 ( BL53, BLN53, WL9);
sram_cell_6t_3 inst_cell_8_53 ( BL53, BLN53, WL8);
sram_cell_6t_3 inst_cell_7_53 ( BL53, BLN53, WL7);
sram_cell_6t_3 inst_cell_6_53 ( BL53, BLN53, WL6);
sram_cell_6t_3 inst_cell_5_53 ( BL53, BLN53, WL5);
sram_cell_6t_3 inst_cell_4_53 ( BL53, BLN53, WL4);
sram_cell_6t_3 inst_cell_3_53 ( BL53, BLN53, WL3);
sram_cell_6t_3 inst_cell_2_53 ( BL53, BLN53, WL2);
sram_cell_6t_3 inst_cell_1_53 ( BL53, BLN53, WL1);
sram_cell_6t_3 inst_cell_0_53 ( BL53, BLN53, WL0);
sram_cell_6t_3 inst_cell_13_52 ( BL52, BLN52, WL13);
sram_cell_6t_3 inst_cell_12_52 ( BL52, BLN52, WL12);
sram_cell_6t_3 inst_cell_11_52 ( BL52, BLN52, WL11);
sram_cell_6t_3 inst_cell_10_52 ( BL52, BLN52, WL10);
sram_cell_6t_3 inst_cell_9_52 ( BL52, BLN52, WL9);
sram_cell_6t_3 inst_cell_8_52 ( BL52, BLN52, WL8);
sram_cell_6t_3 inst_cell_7_52 ( BL52, BLN52, WL7);
sram_cell_6t_3 inst_cell_6_52 ( BL52, BLN52, WL6);
sram_cell_6t_3 inst_cell_5_52 ( BL52, BLN52, WL5);
sram_cell_6t_3 inst_cell_4_52 ( BL52, BLN52, WL4);
sram_cell_6t_3 inst_cell_3_52 ( BL52, BLN52, WL3);
sram_cell_6t_3 inst_cell_2_52 ( BL52, BLN52, WL2);
sram_cell_6t_3 inst_cell_1_52 ( BL52, BLN52, WL1);
sram_cell_6t_3 inst_cell_0_52 ( BL52, BLN52, WL0);
sram_cell_6t_3 inst_cell_13_51 ( BL51, BLN51, WL13);
sram_cell_6t_3 inst_cell_12_51 ( BL51, BLN51, WL12);
sram_cell_6t_3 inst_cell_11_51 ( BL51, BLN51, WL11);
sram_cell_6t_3 inst_cell_10_51 ( BL51, BLN51, WL10);
sram_cell_6t_3 inst_cell_9_51 ( BL51, BLN51, WL9);
sram_cell_6t_3 inst_cell_8_51 ( BL51, BLN51, WL8);
sram_cell_6t_3 inst_cell_7_51 ( BL51, BLN51, WL7);
sram_cell_6t_3 inst_cell_6_51 ( BL51, BLN51, WL6);
sram_cell_6t_3 inst_cell_5_51 ( BL51, BLN51, WL5);
sram_cell_6t_3 inst_cell_4_51 ( BL51, BLN51, WL4);
sram_cell_6t_3 inst_cell_3_51 ( BL51, BLN51, WL3);
sram_cell_6t_3 inst_cell_2_51 ( BL51, BLN51, WL2);
sram_cell_6t_3 inst_cell_1_51 ( BL51, BLN51, WL1);
sram_cell_6t_3 inst_cell_0_51 ( BL51, BLN51, WL0);
sram_cell_6t_3 inst_cell_13_50 ( BL50, BLN50, WL13);
sram_cell_6t_3 inst_cell_12_50 ( BL50, BLN50, WL12);
sram_cell_6t_3 inst_cell_11_50 ( BL50, BLN50, WL11);
sram_cell_6t_3 inst_cell_10_50 ( BL50, BLN50, WL10);
sram_cell_6t_3 inst_cell_9_50 ( BL50, BLN50, WL9);
sram_cell_6t_3 inst_cell_8_50 ( BL50, BLN50, WL8);
sram_cell_6t_3 inst_cell_7_50 ( BL50, BLN50, WL7);
sram_cell_6t_3 inst_cell_6_50 ( BL50, BLN50, WL6);
sram_cell_6t_3 inst_cell_5_50 ( BL50, BLN50, WL5);
sram_cell_6t_3 inst_cell_4_50 ( BL50, BLN50, WL4);
sram_cell_6t_3 inst_cell_3_50 ( BL50, BLN50, WL3);
sram_cell_6t_3 inst_cell_2_50 ( BL50, BLN50, WL2);
sram_cell_6t_3 inst_cell_1_50 ( BL50, BLN50, WL1);
sram_cell_6t_3 inst_cell_0_50 ( BL50, BLN50, WL0);
sram_cell_6t_3 inst_cell_13_49 ( BL49, BLN49, WL13);
sram_cell_6t_3 inst_cell_12_49 ( BL49, BLN49, WL12);
sram_cell_6t_3 inst_cell_11_49 ( BL49, BLN49, WL11);
sram_cell_6t_3 inst_cell_10_49 ( BL49, BLN49, WL10);
sram_cell_6t_3 inst_cell_9_49 ( BL49, BLN49, WL9);
sram_cell_6t_3 inst_cell_8_49 ( BL49, BLN49, WL8);
sram_cell_6t_3 inst_cell_7_49 ( BL49, BLN49, WL7);
sram_cell_6t_3 inst_cell_6_49 ( BL49, BLN49, WL6);
sram_cell_6t_3 inst_cell_5_49 ( BL49, BLN49, WL5);
sram_cell_6t_3 inst_cell_4_49 ( BL49, BLN49, WL4);
sram_cell_6t_3 inst_cell_3_49 ( BL49, BLN49, WL3);
sram_cell_6t_3 inst_cell_2_49 ( BL49, BLN49, WL2);
sram_cell_6t_3 inst_cell_1_49 ( BL49, BLN49, WL1);
sram_cell_6t_3 inst_cell_0_49 ( BL49, BLN49, WL0);
sram_cell_6t_3 inst_cell_13_48 ( BL48, BLN48, WL13);
sram_cell_6t_3 inst_cell_12_48 ( BL48, BLN48, WL12);
sram_cell_6t_3 inst_cell_11_48 ( BL48, BLN48, WL11);
sram_cell_6t_3 inst_cell_10_48 ( BL48, BLN48, WL10);
sram_cell_6t_3 inst_cell_9_48 ( BL48, BLN48, WL9);
sram_cell_6t_3 inst_cell_8_48 ( BL48, BLN48, WL8);
sram_cell_6t_3 inst_cell_7_48 ( BL48, BLN48, WL7);
sram_cell_6t_3 inst_cell_6_48 ( BL48, BLN48, WL6);
sram_cell_6t_3 inst_cell_5_48 ( BL48, BLN48, WL5);
sram_cell_6t_3 inst_cell_4_48 ( BL48, BLN48, WL4);
sram_cell_6t_3 inst_cell_3_48 ( BL48, BLN48, WL3);
sram_cell_6t_3 inst_cell_2_48 ( BL48, BLN48, WL2);
sram_cell_6t_3 inst_cell_1_48 ( BL48, BLN48, WL1);
sram_cell_6t_3 inst_cell_0_48 ( BL48, BLN48, WL0);
sram_cell_6t_3 inst_cell_13_47 ( BL47, BLN47, WL13);
sram_cell_6t_3 inst_cell_12_47 ( BL47, BLN47, WL12);
sram_cell_6t_3 inst_cell_11_47 ( BL47, BLN47, WL11);
sram_cell_6t_3 inst_cell_10_47 ( BL47, BLN47, WL10);
sram_cell_6t_3 inst_cell_9_47 ( BL47, BLN47, WL9);
sram_cell_6t_3 inst_cell_8_47 ( BL47, BLN47, WL8);
sram_cell_6t_3 inst_cell_7_47 ( BL47, BLN47, WL7);
sram_cell_6t_3 inst_cell_6_47 ( BL47, BLN47, WL6);
sram_cell_6t_3 inst_cell_5_47 ( BL47, BLN47, WL5);
sram_cell_6t_3 inst_cell_4_47 ( BL47, BLN47, WL4);
sram_cell_6t_3 inst_cell_3_47 ( BL47, BLN47, WL3);
sram_cell_6t_3 inst_cell_2_47 ( BL47, BLN47, WL2);
sram_cell_6t_3 inst_cell_1_47 ( BL47, BLN47, WL1);
sram_cell_6t_3 inst_cell_0_47 ( BL47, BLN47, WL0);
sram_cell_6t_3 inst_cell_13_46 ( BL46, BLN46, WL13);
sram_cell_6t_3 inst_cell_12_46 ( BL46, BLN46, WL12);
sram_cell_6t_3 inst_cell_11_46 ( BL46, BLN46, WL11);
sram_cell_6t_3 inst_cell_10_46 ( BL46, BLN46, WL10);
sram_cell_6t_3 inst_cell_9_46 ( BL46, BLN46, WL9);
sram_cell_6t_3 inst_cell_8_46 ( BL46, BLN46, WL8);
sram_cell_6t_3 inst_cell_7_46 ( BL46, BLN46, WL7);
sram_cell_6t_3 inst_cell_6_46 ( BL46, BLN46, WL6);
sram_cell_6t_3 inst_cell_5_46 ( BL46, BLN46, WL5);
sram_cell_6t_3 inst_cell_4_46 ( BL46, BLN46, WL4);
sram_cell_6t_3 inst_cell_3_46 ( BL46, BLN46, WL3);
sram_cell_6t_3 inst_cell_2_46 ( BL46, BLN46, WL2);
sram_cell_6t_3 inst_cell_1_46 ( BL46, BLN46, WL1);
sram_cell_6t_3 inst_cell_0_46 ( BL46, BLN46, WL0);
sram_cell_6t_3 inst_cell_13_45 ( BL45, BLN45, WL13);
sram_cell_6t_3 inst_cell_12_45 ( BL45, BLN45, WL12);
sram_cell_6t_3 inst_cell_11_45 ( BL45, BLN45, WL11);
sram_cell_6t_3 inst_cell_10_45 ( BL45, BLN45, WL10);
sram_cell_6t_3 inst_cell_9_45 ( BL45, BLN45, WL9);
sram_cell_6t_3 inst_cell_8_45 ( BL45, BLN45, WL8);
sram_cell_6t_3 inst_cell_7_45 ( BL45, BLN45, WL7);
sram_cell_6t_3 inst_cell_6_45 ( BL45, BLN45, WL6);
sram_cell_6t_3 inst_cell_5_45 ( BL45, BLN45, WL5);
sram_cell_6t_3 inst_cell_4_45 ( BL45, BLN45, WL4);
sram_cell_6t_3 inst_cell_3_45 ( BL45, BLN45, WL3);
sram_cell_6t_3 inst_cell_2_45 ( BL45, BLN45, WL2);
sram_cell_6t_3 inst_cell_1_45 ( BL45, BLN45, WL1);
sram_cell_6t_3 inst_cell_0_45 ( BL45, BLN45, WL0);
sram_cell_6t_3 inst_cell_13_44 ( BL44, BLN44, WL13);
sram_cell_6t_3 inst_cell_12_44 ( BL44, BLN44, WL12);
sram_cell_6t_3 inst_cell_11_44 ( BL44, BLN44, WL11);
sram_cell_6t_3 inst_cell_10_44 ( BL44, BLN44, WL10);
sram_cell_6t_3 inst_cell_9_44 ( BL44, BLN44, WL9);
sram_cell_6t_3 inst_cell_8_44 ( BL44, BLN44, WL8);
sram_cell_6t_3 inst_cell_7_44 ( BL44, BLN44, WL7);
sram_cell_6t_3 inst_cell_6_44 ( BL44, BLN44, WL6);
sram_cell_6t_3 inst_cell_5_44 ( BL44, BLN44, WL5);
sram_cell_6t_3 inst_cell_4_44 ( BL44, BLN44, WL4);
sram_cell_6t_3 inst_cell_3_44 ( BL44, BLN44, WL3);
sram_cell_6t_3 inst_cell_2_44 ( BL44, BLN44, WL2);
sram_cell_6t_3 inst_cell_1_44 ( BL44, BLN44, WL1);
sram_cell_6t_3 inst_cell_0_44 ( BL44, BLN44, WL0);
sram_cell_6t_3 inst_cell_13_43 ( BL43, BLN43, WL13);
sram_cell_6t_3 inst_cell_12_43 ( BL43, BLN43, WL12);
sram_cell_6t_3 inst_cell_11_43 ( BL43, BLN43, WL11);
sram_cell_6t_3 inst_cell_10_43 ( BL43, BLN43, WL10);
sram_cell_6t_3 inst_cell_9_43 ( BL43, BLN43, WL9);
sram_cell_6t_3 inst_cell_8_43 ( BL43, BLN43, WL8);
sram_cell_6t_3 inst_cell_7_43 ( BL43, BLN43, WL7);
sram_cell_6t_3 inst_cell_6_43 ( BL43, BLN43, WL6);
sram_cell_6t_3 inst_cell_5_43 ( BL43, BLN43, WL5);
sram_cell_6t_3 inst_cell_4_43 ( BL43, BLN43, WL4);
sram_cell_6t_3 inst_cell_3_43 ( BL43, BLN43, WL3);
sram_cell_6t_3 inst_cell_2_43 ( BL43, BLN43, WL2);
sram_cell_6t_3 inst_cell_1_43 ( BL43, BLN43, WL1);
sram_cell_6t_3 inst_cell_0_43 ( BL43, BLN43, WL0);
sram_cell_6t_3 inst_cell_13_42 ( BL42, BLN42, WL13);
sram_cell_6t_3 inst_cell_12_42 ( BL42, BLN42, WL12);
sram_cell_6t_3 inst_cell_11_42 ( BL42, BLN42, WL11);
sram_cell_6t_3 inst_cell_10_42 ( BL42, BLN42, WL10);
sram_cell_6t_3 inst_cell_9_42 ( BL42, BLN42, WL9);
sram_cell_6t_3 inst_cell_8_42 ( BL42, BLN42, WL8);
sram_cell_6t_3 inst_cell_7_42 ( BL42, BLN42, WL7);
sram_cell_6t_3 inst_cell_6_42 ( BL42, BLN42, WL6);
sram_cell_6t_3 inst_cell_5_42 ( BL42, BLN42, WL5);
sram_cell_6t_3 inst_cell_4_42 ( BL42, BLN42, WL4);
sram_cell_6t_3 inst_cell_3_42 ( BL42, BLN42, WL3);
sram_cell_6t_3 inst_cell_2_42 ( BL42, BLN42, WL2);
sram_cell_6t_3 inst_cell_1_42 ( BL42, BLN42, WL1);
sram_cell_6t_3 inst_cell_0_42 ( BL42, BLN42, WL0);
sram_cell_6t_3 inst_cell_13_41 ( BL41, BLN41, WL13);
sram_cell_6t_3 inst_cell_12_41 ( BL41, BLN41, WL12);
sram_cell_6t_3 inst_cell_11_41 ( BL41, BLN41, WL11);
sram_cell_6t_3 inst_cell_10_41 ( BL41, BLN41, WL10);
sram_cell_6t_3 inst_cell_9_41 ( BL41, BLN41, WL9);
sram_cell_6t_3 inst_cell_8_41 ( BL41, BLN41, WL8);
sram_cell_6t_3 inst_cell_7_41 ( BL41, BLN41, WL7);
sram_cell_6t_3 inst_cell_6_41 ( BL41, BLN41, WL6);
sram_cell_6t_3 inst_cell_5_41 ( BL41, BLN41, WL5);
sram_cell_6t_3 inst_cell_4_41 ( BL41, BLN41, WL4);
sram_cell_6t_3 inst_cell_3_41 ( BL41, BLN41, WL3);
sram_cell_6t_3 inst_cell_2_41 ( BL41, BLN41, WL2);
sram_cell_6t_3 inst_cell_1_41 ( BL41, BLN41, WL1);
sram_cell_6t_3 inst_cell_0_41 ( BL41, BLN41, WL0);
sram_cell_6t_3 inst_cell_13_40 ( BL40, BLN40, WL13);
sram_cell_6t_3 inst_cell_12_40 ( BL40, BLN40, WL12);
sram_cell_6t_3 inst_cell_11_40 ( BL40, BLN40, WL11);
sram_cell_6t_3 inst_cell_10_40 ( BL40, BLN40, WL10);
sram_cell_6t_3 inst_cell_9_40 ( BL40, BLN40, WL9);
sram_cell_6t_3 inst_cell_8_40 ( BL40, BLN40, WL8);
sram_cell_6t_3 inst_cell_7_40 ( BL40, BLN40, WL7);
sram_cell_6t_3 inst_cell_6_40 ( BL40, BLN40, WL6);
sram_cell_6t_3 inst_cell_5_40 ( BL40, BLN40, WL5);
sram_cell_6t_3 inst_cell_4_40 ( BL40, BLN40, WL4);
sram_cell_6t_3 inst_cell_3_40 ( BL40, BLN40, WL3);
sram_cell_6t_3 inst_cell_2_40 ( BL40, BLN40, WL2);
sram_cell_6t_3 inst_cell_1_40 ( BL40, BLN40, WL1);
sram_cell_6t_3 inst_cell_0_40 ( BL40, BLN40, WL0);
sram_cell_6t_3 inst_cell_13_39 ( BL39, BLN39, WL13);
sram_cell_6t_3 inst_cell_12_39 ( BL39, BLN39, WL12);
sram_cell_6t_3 inst_cell_11_39 ( BL39, BLN39, WL11);
sram_cell_6t_3 inst_cell_10_39 ( BL39, BLN39, WL10);
sram_cell_6t_3 inst_cell_9_39 ( BL39, BLN39, WL9);
sram_cell_6t_3 inst_cell_8_39 ( BL39, BLN39, WL8);
sram_cell_6t_3 inst_cell_7_39 ( BL39, BLN39, WL7);
sram_cell_6t_3 inst_cell_6_39 ( BL39, BLN39, WL6);
sram_cell_6t_3 inst_cell_5_39 ( BL39, BLN39, WL5);
sram_cell_6t_3 inst_cell_4_39 ( BL39, BLN39, WL4);
sram_cell_6t_3 inst_cell_3_39 ( BL39, BLN39, WL3);
sram_cell_6t_3 inst_cell_2_39 ( BL39, BLN39, WL2);
sram_cell_6t_3 inst_cell_1_39 ( BL39, BLN39, WL1);
sram_cell_6t_3 inst_cell_0_39 ( BL39, BLN39, WL0);
sram_cell_6t_3 inst_cell_13_38 ( BL38, BLN38, WL13);
sram_cell_6t_3 inst_cell_12_38 ( BL38, BLN38, WL12);
sram_cell_6t_3 inst_cell_11_38 ( BL38, BLN38, WL11);
sram_cell_6t_3 inst_cell_10_38 ( BL38, BLN38, WL10);
sram_cell_6t_3 inst_cell_9_38 ( BL38, BLN38, WL9);
sram_cell_6t_3 inst_cell_8_38 ( BL38, BLN38, WL8);
sram_cell_6t_3 inst_cell_7_38 ( BL38, BLN38, WL7);
sram_cell_6t_3 inst_cell_6_38 ( BL38, BLN38, WL6);
sram_cell_6t_3 inst_cell_5_38 ( BL38, BLN38, WL5);
sram_cell_6t_3 inst_cell_4_38 ( BL38, BLN38, WL4);
sram_cell_6t_3 inst_cell_3_38 ( BL38, BLN38, WL3);
sram_cell_6t_3 inst_cell_2_38 ( BL38, BLN38, WL2);
sram_cell_6t_3 inst_cell_1_38 ( BL38, BLN38, WL1);
sram_cell_6t_3 inst_cell_0_38 ( BL38, BLN38, WL0);
sram_cell_6t_3 inst_cell_13_37 ( BL37, BLN37, WL13);
sram_cell_6t_3 inst_cell_12_37 ( BL37, BLN37, WL12);
sram_cell_6t_3 inst_cell_11_37 ( BL37, BLN37, WL11);
sram_cell_6t_3 inst_cell_10_37 ( BL37, BLN37, WL10);
sram_cell_6t_3 inst_cell_9_37 ( BL37, BLN37, WL9);
sram_cell_6t_3 inst_cell_8_37 ( BL37, BLN37, WL8);
sram_cell_6t_3 inst_cell_7_37 ( BL37, BLN37, WL7);
sram_cell_6t_3 inst_cell_6_37 ( BL37, BLN37, WL6);
sram_cell_6t_3 inst_cell_5_37 ( BL37, BLN37, WL5);
sram_cell_6t_3 inst_cell_4_37 ( BL37, BLN37, WL4);
sram_cell_6t_3 inst_cell_3_37 ( BL37, BLN37, WL3);
sram_cell_6t_3 inst_cell_2_37 ( BL37, BLN37, WL2);
sram_cell_6t_3 inst_cell_1_37 ( BL37, BLN37, WL1);
sram_cell_6t_3 inst_cell_0_37 ( BL37, BLN37, WL0);
sram_cell_6t_3 inst_cell_13_36 ( BL36, BLN36, WL13);
sram_cell_6t_3 inst_cell_12_36 ( BL36, BLN36, WL12);
sram_cell_6t_3 inst_cell_11_36 ( BL36, BLN36, WL11);
sram_cell_6t_3 inst_cell_10_36 ( BL36, BLN36, WL10);
sram_cell_6t_3 inst_cell_9_36 ( BL36, BLN36, WL9);
sram_cell_6t_3 inst_cell_8_36 ( BL36, BLN36, WL8);
sram_cell_6t_3 inst_cell_7_36 ( BL36, BLN36, WL7);
sram_cell_6t_3 inst_cell_6_36 ( BL36, BLN36, WL6);
sram_cell_6t_3 inst_cell_5_36 ( BL36, BLN36, WL5);
sram_cell_6t_3 inst_cell_4_36 ( BL36, BLN36, WL4);
sram_cell_6t_3 inst_cell_3_36 ( BL36, BLN36, WL3);
sram_cell_6t_3 inst_cell_2_36 ( BL36, BLN36, WL2);
sram_cell_6t_3 inst_cell_1_36 ( BL36, BLN36, WL1);
sram_cell_6t_3 inst_cell_0_36 ( BL36, BLN36, WL0);
sram_cell_6t_3 inst_cell_13_35 ( BL35, BLN35, WL13);
sram_cell_6t_3 inst_cell_12_35 ( BL35, BLN35, WL12);
sram_cell_6t_3 inst_cell_11_35 ( BL35, BLN35, WL11);
sram_cell_6t_3 inst_cell_10_35 ( BL35, BLN35, WL10);
sram_cell_6t_3 inst_cell_9_35 ( BL35, BLN35, WL9);
sram_cell_6t_3 inst_cell_8_35 ( BL35, BLN35, WL8);
sram_cell_6t_3 inst_cell_7_35 ( BL35, BLN35, WL7);
sram_cell_6t_3 inst_cell_6_35 ( BL35, BLN35, WL6);
sram_cell_6t_3 inst_cell_5_35 ( BL35, BLN35, WL5);
sram_cell_6t_3 inst_cell_4_35 ( BL35, BLN35, WL4);
sram_cell_6t_3 inst_cell_3_35 ( BL35, BLN35, WL3);
sram_cell_6t_3 inst_cell_2_35 ( BL35, BLN35, WL2);
sram_cell_6t_3 inst_cell_1_35 ( BL35, BLN35, WL1);
sram_cell_6t_3 inst_cell_0_35 ( BL35, BLN35, WL0);
sram_cell_6t_3 inst_cell_13_34 ( BL34, BLN34, WL13);
sram_cell_6t_3 inst_cell_12_34 ( BL34, BLN34, WL12);
sram_cell_6t_3 inst_cell_11_34 ( BL34, BLN34, WL11);
sram_cell_6t_3 inst_cell_10_34 ( BL34, BLN34, WL10);
sram_cell_6t_3 inst_cell_9_34 ( BL34, BLN34, WL9);
sram_cell_6t_3 inst_cell_8_34 ( BL34, BLN34, WL8);
sram_cell_6t_3 inst_cell_7_34 ( BL34, BLN34, WL7);
sram_cell_6t_3 inst_cell_6_34 ( BL34, BLN34, WL6);
sram_cell_6t_3 inst_cell_5_34 ( BL34, BLN34, WL5);
sram_cell_6t_3 inst_cell_4_34 ( BL34, BLN34, WL4);
sram_cell_6t_3 inst_cell_3_34 ( BL34, BLN34, WL3);
sram_cell_6t_3 inst_cell_2_34 ( BL34, BLN34, WL2);
sram_cell_6t_3 inst_cell_1_34 ( BL34, BLN34, WL1);
sram_cell_6t_3 inst_cell_0_34 ( BL34, BLN34, WL0);
sram_cell_6t_3 inst_cell_13_33 ( BL33, BLN33, WL13);
sram_cell_6t_3 inst_cell_13_32 ( BL32, BLN32, WL13);
sram_cell_6t_3 inst_cell_12_33 ( BL33, BLN33, WL12);
sram_cell_6t_3 inst_cell_12_32 ( BL32, BLN32, WL12);
sram_cell_6t_3 inst_cell_11_33 ( BL33, BLN33, WL11);
sram_cell_6t_3 inst_cell_11_32 ( BL32, BLN32, WL11);
sram_cell_6t_3 inst_cell_10_33 ( BL33, BLN33, WL10);
sram_cell_6t_3 inst_cell_10_32 ( BL32, BLN32, WL10);
sram_cell_6t_3 inst_cell_9_33 ( BL33, BLN33, WL9);
sram_cell_6t_3 inst_cell_9_32 ( BL32, BLN32, WL9);
sram_cell_6t_3 inst_cell_8_33 ( BL33, BLN33, WL8);
sram_cell_6t_3 inst_cell_8_32 ( BL32, BLN32, WL8);
sram_cell_6t_3 inst_cell_7_33 ( BL33, BLN33, WL7);
sram_cell_6t_3 inst_cell_7_32 ( BL32, BLN32, WL7);
sram_cell_6t_3 inst_cell_6_33 ( BL33, BLN33, WL6);
sram_cell_6t_3 inst_cell_6_32 ( BL32, BLN32, WL6);
sram_cell_6t_3 inst_cell_5_33 ( BL33, BLN33, WL5);
sram_cell_6t_3 inst_cell_5_32 ( BL32, BLN32, WL5);
sram_cell_6t_3 inst_cell_4_33 ( BL33, BLN33, WL4);
sram_cell_6t_3 inst_cell_4_32 ( BL32, BLN32, WL4);
sram_cell_6t_3 inst_cell_3_33 ( BL33, BLN33, WL3);
sram_cell_6t_3 inst_cell_3_32 ( BL32, BLN32, WL3);
sram_cell_6t_3 inst_cell_2_33 ( BL33, BLN33, WL2);
sram_cell_6t_3 inst_cell_2_32 ( BL32, BLN32, WL2);
sram_cell_6t_3 inst_cell_1_33 ( BL33, BLN33, WL1);
sram_cell_6t_3 inst_cell_0_33 ( BL33, BLN33, WL0);
sram_cell_6t_3 inst_cell_1_32 ( BL32, BLN32, WL1);
sram_cell_6t_3 inst_cell_0_32 ( BL32, BLN32, WL0);
inverter_compiler inst_invComp ( clk_bar, clk);
sense_amp_clocked_compiler inst_senAmp7 ( dout7, net7274, DL7, DLN7,
     sense_en);
sense_amp_clocked_compiler inst_senAmp6 ( dout6, net7275, DL6, DLN6,
     sense_en);
sense_amp_clocked_compiler inst_senAmp5 ( dout5, net7276, DL5, DLN5,
     sense_en);
sense_amp_clocked_compiler inst_senAmp4 ( dout4, net7277, DL4, DLN4,
     sense_en);
sense_amp_clocked_compiler inst_senAmp3 ( dout3, net7278, DL3, DLN3,
     sense_en);
sense_amp_clocked_compiler inst_senAmp2 ( dout2, net7279, DL2, DLN2,
     sense_en);
sense_amp_clocked_compiler inst_senAmp0 ( dout0, net7280, DL0, DLN0,
     sense_en);
sense_amp_clocked_compiler inst_senAmp1 ( dout1, net7281, DL1, DLN1,
     sense_en);
write_driver_compiler inst_writeDriver7 ( DL7, DLN7, clk_bar, din7,
     write_en);
write_driver_compiler inst_writeDriver6 ( DL6, DLN6, clk_bar, din6,
     write_en);
write_driver_compiler inst_writeDriver5 ( DL5, DLN5, clk_bar, din5,
     write_en);
write_driver_compiler inst_writeDriver4 ( DL4, DLN4, clk_bar, din4,
     write_en);
write_driver_compiler inst_writeDriver3 ( DL3, DLN3, clk_bar, din3,
     write_en);
write_driver_compiler inst_writeDriver2 ( DL2, DLN2, clk_bar, din2,
     write_en);
write_driver_compiler inst_writeDriver0 ( DL0, DLN0, clk_bar, din0,
     write_en);
write_driver_compiler inst_writeDriver1 ( DL1, DLN1, clk_bar, din1,
     write_en);
colDecoder inst_colDec ( .YF7(SL7), .YF6(SL6), .YF5(SL5), .YF4(SL4),
     .YF3(SL3), .YF2(SL2), .YF1(SL1), .YF0(SL0), .CLK(clk_bar),
     .A2_inv(inv_addr8), .A2(addr8), .A1_inv(inv_addr7), .A1(addr7),
     .A0_inv(inv_addr6), .A0(addr6));
invCol inst_invCol ( .Abar2(inv_addr8), .Abar1(inv_addr7),
     .Abar0(inv_addr6), .A2(addr8), .A1(addr7), .A0(addr6));
precharge_compiler inst_precharge63 ( BL63, BLN63, clk_bar);
precharge_compiler inst_precharge62 ( BL62, BLN62, clk_bar);
precharge_compiler inst_precharge61 ( BL61, BLN61, clk_bar);
precharge_compiler inst_precharge60 ( BL60, BLN60, clk_bar);
precharge_compiler inst_precharge59 ( BL59, BLN59, clk_bar);
precharge_compiler inst_precharge58 ( BL58, BLN58, clk_bar);
precharge_compiler inst_precharge57 ( BL57, BLN57, clk_bar);
precharge_compiler inst_precharge56 ( BL56, BLN56, clk_bar);
precharge_compiler inst_precharge55 ( BL55, BLN55, clk_bar);
precharge_compiler inst_precharge54 ( BL54, BLN54, clk_bar);
precharge_compiler inst_precharge53 ( BL53, BLN53, clk_bar);
precharge_compiler inst_precharge52 ( BL52, BLN52, clk_bar);
precharge_compiler inst_precharge51 ( BL51, BLN51, clk_bar);
precharge_compiler inst_precharge50 ( BL50, BLN50, clk_bar);
precharge_compiler inst_precharge49 ( BL49, BLN49, clk_bar);
precharge_compiler inst_precharge48 ( BL48, BLN48, clk_bar);
precharge_compiler inst_precharge47 ( BL47, BLN47, clk_bar);
precharge_compiler inst_precharge46 ( BL46, BLN46, clk_bar);
precharge_compiler inst_precharge45 ( BL45, BLN45, clk_bar);
precharge_compiler inst_precharge44 ( BL44, BLN44, clk_bar);
precharge_compiler inst_precharge43 ( BL43, BLN43, clk_bar);
precharge_compiler inst_precharge42 ( BL42, BLN42, clk_bar);
precharge_compiler inst_precharge41 ( BL41, BLN41, clk_bar);
precharge_compiler inst_precharge40 ( BL40, BLN40, clk_bar);
precharge_compiler inst_precharge39 ( BL39, BLN39, clk_bar);
precharge_compiler inst_precharge38 ( BL38, BLN38, clk_bar);
precharge_compiler inst_precharge37 ( BL37, BLN37, clk_bar);
precharge_compiler inst_precharge36 ( BL36, BLN36, clk_bar);
precharge_compiler inst_precharge35 ( BL35, BLN35, clk_bar);
precharge_compiler inst_precharge34 ( BL34, BLN34, clk_bar);
precharge_compiler inst_precharge33 ( BL33, BLN33, clk_bar);
precharge_compiler inst_precharge32 ( BL32, BLN32, clk_bar);
precharge_compiler inst_precharge31 ( BL31, BLN31, clk_bar);
precharge_compiler inst_precharge30 ( BL30, BLN30, clk_bar);
precharge_compiler inst_precharge29 ( BL29, BLN29, clk_bar);
precharge_compiler inst_precharge28 ( BL28, BLN28, clk_bar);
precharge_compiler inst_precharge27 ( BL27, BLN27, clk_bar);
precharge_compiler inst_precharge26 ( BL26, BLN26, clk_bar);
precharge_compiler inst_precharge25 ( BL25, BLN25, clk_bar);
precharge_compiler inst_precharge24 ( BL24, BLN24, clk_bar);
precharge_compiler inst_precharge23 ( BL23, BLN23, clk_bar);
precharge_compiler inst_precharge22 ( BL22, BLN22, clk_bar);
precharge_compiler inst_precharge21 ( BL21, BLN21, clk_bar);
precharge_compiler inst_precharge20 ( BL20, BLN20, clk_bar);
precharge_compiler inst_precharge19 ( BL19, BLN19, clk_bar);
precharge_compiler inst_precharge18 ( BL18, BLN18, clk_bar);
precharge_compiler inst_precharge17 ( BL17, BLN17, clk_bar);
precharge_compiler inst_precharge16 ( BL16, BLN16, clk_bar);
precharge_compiler inst_precharge15 ( BL15, BLN15, clk_bar);
precharge_compiler inst_precharge14 ( BL14, BLN14, clk_bar);
precharge_compiler inst_precharge13 ( BL13, BLN13, clk_bar);
precharge_compiler inst_precharge12 ( BL12, BLN12, clk_bar);
precharge_compiler inst_precharge11 ( BL11, BLN11, clk_bar);
precharge_compiler inst_precharge10 ( BL10, BLN10, clk_bar);
precharge_compiler inst_precharge9 ( BL9, BLN9, clk_bar);
precharge_compiler inst_precharge8 ( BL8, BLN8, clk_bar);
precharge_compiler inst_precharge7 ( BL7, BLN7, clk_bar);
precharge_compiler inst_precharge6 ( BL6, BLN6, clk_bar);
precharge_compiler inst_precharge5 ( BL5, BLN5, clk_bar);
precharge_compiler inst_precharge4 ( BL4, BLN4, clk_bar);
precharge_compiler inst_precharge3 ( BL3, BLN3, clk_bar);
precharge_compiler inst_precharge2 ( BL2, BLN2, clk_bar);
precharge_compiler inst_precharge1 ( BL1, BLN1, clk_bar);
precharge_compiler inst_precharge0 ( BL0, BLN0, clk_bar);
columnMux inst_colMux7 ( .Ybar(DLN7), .Y(DL7), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN63), .A7(BL63), .Abar6(BLN62), .A6(BL62),
     .Abar5(BLN61), .A5(BL61), .Abar4(BLN60), .A4(BL60), .Abar3(BLN59),
     .A3(BL59), .Abar2(BLN58), .A2(BL58), .Abar1(BLN57), .A1(BL57),
     .Abar0(BLN56), .A0(BL56));
columnMux inst_colMux6 ( .Ybar(DLN6), .Y(DL6), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN55), .A7(BL55), .Abar6(BLN54), .A6(BL54),
     .Abar5(BLN53), .A5(BL53), .Abar4(BLN52), .A4(BL52), .Abar3(BLN51),
     .A3(BL51), .Abar2(BLN50), .A2(BL50), .Abar1(BLN49), .A1(BL49),
     .Abar0(BLN48), .A0(BL48));
columnMux inst_colMux5 ( .Ybar(DLN5), .Y(DL5), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN47), .A7(BL47), .Abar6(BLN46), .A6(BL46),
     .Abar5(BLN45), .A5(BL45), .Abar4(BLN44), .A4(BL44), .Abar3(BLN43),
     .A3(BL43), .Abar2(BLN42), .A2(BL42), .Abar1(BLN41), .A1(BL41),
     .Abar0(BLN40), .A0(BL40));
columnMux inst_colMux4 ( .Ybar(DLN4), .Y(DL4), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN39), .A7(BL39), .Abar6(BLN38), .A6(BL38),
     .Abar5(BLN37), .A5(BL37), .Abar4(BLN36), .A4(BL36), .Abar3(BLN35),
     .A3(BL35), .Abar2(BLN34), .A2(BL34), .Abar1(BLN33), .A1(BL33),
     .Abar0(BLN32), .A0(BL32));
columnMux inst_colMux3 ( .Ybar(DLN3), .Y(DL3), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN31), .A7(BL31), .Abar6(BLN30), .A6(BL30),
     .Abar5(BLN29), .A5(BL29), .Abar4(BLN28), .A4(BL28), .Abar3(BLN27),
     .A3(BL27), .Abar2(BLN26), .A2(BL26), .Abar1(BLN25), .A1(BL25),
     .Abar0(BLN24), .A0(BL24));
columnMux inst_colMux2 ( .Ybar(DLN2), .Y(DL2), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN23), .A7(BL23), .Abar6(BLN22), .A6(BL22),
     .Abar5(BLN21), .A5(BL21), .Abar4(BLN20), .A4(BL20), .Abar3(BLN19),
     .A3(BL19), .Abar2(BLN18), .A2(BL18), .Abar1(BLN17), .A1(BL17),
     .Abar0(BLN16), .A0(BL16));
columnMux inst_colMux1 ( .Ybar(DLN1), .Y(DL1), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN15), .A7(BL15), .Abar6(BLN14), .A6(BL14),
     .Abar5(BLN13), .A5(BL13), .Abar4(BLN12), .A4(BL12), .Abar3(BLN11),
     .A3(BL11), .Abar2(BLN10), .A2(BL10), .Abar1(BLN9), .A1(BL9),
     .Abar0(BLN8), .A0(BL8));
columnMux inst_colMux0 ( .Ybar(DLN0), .Y(DL0), .sel7(SL7), .sel6(SL6),
     .sel5(SL5), .sel4(SL4), .sel3(SL3), .sel2(SL2), .sel1(SL1),
     .sel0(SL0), .Abar7(BLN7), .A7(BL7), .Abar6(BLN6), .A6(BL6),
     .Abar5(BLN5), .A5(BL5), .Abar4(BLN4), .A4(BL4), .Abar3(BLN3),
     .A3(BL3), .Abar2(BLN2), .A2(BL2), .Abar1(BLN1), .A1(BL1),
     .Abar0(BLN0), .A0(BL0));
invRow inst_invRow ( .Abar5(inv_addr5), .Abar4(inv_addr4),
     .Abar3(inv_addr3), .Abar2(inv_addr2), .Abar1(inv_addr1),
     .Abar0(inv_addr0), .A5(addr5), .A4(addr4), .A3(addr3), .A2(addr2),
     .A1(addr1), .A0(addr0));
rowDecoder inst_rowDec ( .YF63(WL63), .YF62(WL62), .YF61(WL61),
     .YF60(WL60), .YF59(WL59), .YF58(WL58), .YF57(WL57), .YF56(WL56),
     .YF55(WL55), .YF54(WL54), .YF53(WL53), .YF52(WL52), .YF51(WL51),
     .YF50(WL50), .YF49(WL49), .YF48(WL48), .YF47(WL47), .YF46(WL46),
     .YF45(WL45), .YF44(WL44), .YF43(WL43), .YF42(WL42), .YF41(WL41),
     .YF40(WL40), .YF39(WL39), .YF38(WL38), .YF37(WL37), .YF36(WL36),
     .YF35(WL35), .YF34(WL34), .YF33(WL33), .YF32(WL32), .YF31(WL31),
     .YF30(WL30), .YF29(WL29), .YF28(WL28), .YF27(WL27), .YF26(WL26),
     .YF25(WL25), .YF24(WL24), .YF23(WL23), .YF22(WL22), .YF21(WL21),
     .YF20(WL20), .YF19(WL19), .YF18(WL18), .YF17(WL17), .YF16(WL16),
     .YF15(WL15), .YF14(WL14), .YF13(WL13), .YF12(WL12), .YF11(WL11),
     .YF10(WL10), .YF9(WL9), .YF8(WL8), .YF7(WL7), .YF6(WL6),
     .YF5(WL5), .YF4(WL4), .YF3(WL3), .YF2(WL2), .YF1(WL1), .YF0(WL0),
     .CLK(clk_bar), .A5_inv(inv_addr5), .A5(addr5), .A4_inv(inv_addr4),
     .A4(addr4), .A3_inv(inv_addr3), .A3(addr3), .A2_inv(inv_addr2),
     .A2(addr2), .A1_inv(inv_addr1), .A1(addr1), .A0_inv(inv_addr0),
     .A0(addr0));

endmodule


// End HDL models
