`timescale 1ns / 1ps 

module invRow(A0,A1,A2,A3,A4,A5,A6,Abar0,Abar1,Abar2,Abar3,Abar4,Abar5,Abar6);
input A0;
input A1;
input A2;
input A3;
input A4;
input A5;
input A6;
output Abar0;
output Abar1;
output Abar2;
output Abar3;
output Abar4;
output Abar5;
output Abar6;
INVD wire0 (.A(A0),.Y(Abar0));
INVD wire1 (.A(A1),.Y(Abar1));
INVD wire2 (.A(A2),.Y(Abar2));
INVD wire3 (.A(A3),.Y(Abar3));
INVD wire4 (.A(A4),.Y(Abar4));
INVD wire5 (.A(A5),.Y(Abar5));
INVD wire6 (.A(A6),.Y(Abar6));
endmodule
module invCol(A0,A1,Abar0,Abar1);
input A0;
input A1;
output Abar0;
output Abar1;
INVD wire0 (.A(A0),.Y(Abar0));
INVD wire1 (.A(A1),.Y(Abar1));
endmodule
module rowDecoder(A0,A0_inv,A1,A1_inv,A2,A2_inv,A3,A3_inv,A4,A4_inv,A5,A5_inv,A6,A6_inv,CLK,YF0,YF1,YF2,YF3,YF4,YF5,YF6,YF7,YF8,YF9,YF10,YF11,YF12,YF13,YF14,YF15,YF16,YF17,YF18,YF19,YF20,YF21,YF22,YF23,YF24,YF25,YF26,YF27,YF28,YF29,YF30,YF31,YF32,YF33,YF34,YF35,YF36,YF37,YF38,YF39,YF40,YF41,YF42,YF43,YF44,YF45,YF46,YF47,YF48,YF49,YF50,YF51,YF52,YF53,YF54,YF55,YF56,YF57,YF58,YF59,YF60,YF61,YF62,YF63,YF64,YF65,YF66,YF67,YF68,YF69,YF70,YF71,YF72,YF73,YF74,YF75,YF76,YF77,YF78,YF79,YF80,YF81,YF82,YF83,YF84,YF85,YF86,YF87,YF88,YF89,YF90,YF91,YF92,YF93,YF94,YF95,YF96,YF97,YF98,YF99,YF100,YF101,YF102,YF103,YF104,YF105,YF106,YF107,YF108,YF109,YF110,YF111,YF112,YF113,YF114,YF115,YF116,YF117,YF118,YF119,YF120,YF121,YF122,YF123,YF124,YF125,YF126,YF127);
input A0;
input A0_inv;
input A1;
input A1_inv;
input A2;
input A2_inv;
input A3;
input A3_inv;
input A4;
input A4_inv;
input A5;
input A5_inv;
input A6;
input A6_inv;
input CLK;
output YF0;
output YF1;
output YF2;
output YF3;
output YF4;
output YF5;
output YF6;
output YF7;
output YF8;
output YF9;
output YF10;
output YF11;
output YF12;
output YF13;
output YF14;
output YF15;
output YF16;
output YF17;
output YF18;
output YF19;
output YF20;
output YF21;
output YF22;
output YF23;
output YF24;
output YF25;
output YF26;
output YF27;
output YF28;
output YF29;
output YF30;
output YF31;
output YF32;
output YF33;
output YF34;
output YF35;
output YF36;
output YF37;
output YF38;
output YF39;
output YF40;
output YF41;
output YF42;
output YF43;
output YF44;
output YF45;
output YF46;
output YF47;
output YF48;
output YF49;
output YF50;
output YF51;
output YF52;
output YF53;
output YF54;
output YF55;
output YF56;
output YF57;
output YF58;
output YF59;
output YF60;
output YF61;
output YF62;
output YF63;
output YF64;
output YF65;
output YF66;
output YF67;
output YF68;
output YF69;
output YF70;
output YF71;
output YF72;
output YF73;
output YF74;
output YF75;
output YF76;
output YF77;
output YF78;
output YF79;
output YF80;
output YF81;
output YF82;
output YF83;
output YF84;
output YF85;
output YF86;
output YF87;
output YF88;
output YF89;
output YF90;
output YF91;
output YF92;
output YF93;
output YF94;
output YF95;
output YF96;
output YF97;
output YF98;
output YF99;
output YF100;
output YF101;
output YF102;
output YF103;
output YF104;
output YF105;
output YF106;
output YF107;
output YF108;
output YF109;
output YF110;
output YF111;
output YF112;
output YF113;
output YF114;
output YF115;
output YF116;
output YF117;
output YF118;
output YF119;
output YF120;
output YF121;
output YF122;
output YF123;
output YF124;
output YF125;
output YF126;
output YF127;
NANDC2x1 inst_and_b0_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire0_0_0));
INVC inst_inv_b0_0_0 (.A(imd_wire0_0_0),.Y(wire0_0_0));
NANDC2x1 inst_and_b0_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire0_0_1));
INVC inst_inv_b0_0_1 (.A(imd_wire0_0_1),.Y(wire0_0_1));
NANDC2x1 inst_and_b0_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire0_0_2));
INVC inst_inv_b0_0_2 (.A(imd_wire0_0_2),.Y(wire0_0_2));
NANDC2x1 inst_and_b0_1_0 (.A(wire0_0_0),.B(wire0_0_1),.Y(imd_wire0_1_0));
INVC inst_inv_b0_1_0 (.A(imd_wire0_1_0),.Y(wire0_1_0));
NANDC2x1 inst_and_b0_1_1 (.A(A6_inv),.B(wire0_0_2),.Y(imd_wire0_1_1));
INVC inst_inv_b0_1_1 (.A(imd_wire0_1_1),.Y(wire0_1_1));
NANDC2x1 inst_and_b0_2_0 (.A(wire0_1_0),.B(wire0_1_1),.Y(imd_Y0));
INVC inst_inv_b0_2_0 (.A(imd_Y0),.Y(Y0));
NANDC2x1 inst_clockedAND_b0_0 (.A(CLK),.B(Y0),.Y(imd_YF0));
INVC inst_clockedinv_b0_0 (.A(imd_YF0),.Y(YF0));


NANDC2x1 inst_and_b1_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire1_0_0));
INVC inst_inv_b1_0_0 (.A(imd_wire1_0_0),.Y(wire1_0_0));
NANDC2x1 inst_and_b1_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire1_0_1));
INVC inst_inv_b1_0_1 (.A(imd_wire1_0_1),.Y(wire1_0_1));
NANDC2x1 inst_and_b1_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire1_0_2));
INVC inst_inv_b1_0_2 (.A(imd_wire1_0_2),.Y(wire1_0_2));
NANDC2x1 inst_and_b1_1_0 (.A(wire1_0_0),.B(wire1_0_1),.Y(imd_wire1_1_0));
INVC inst_inv_b1_1_0 (.A(imd_wire1_1_0),.Y(wire1_1_0));
NANDC2x1 inst_and_b1_1_1 (.A(A6_inv),.B(wire1_0_2),.Y(imd_wire1_1_1));
INVC inst_inv_b1_1_1 (.A(imd_wire1_1_1),.Y(wire1_1_1));
NANDC2x1 inst_and_b1_2_0 (.A(wire1_1_0),.B(wire1_1_1),.Y(imd_Y1));
INVC inst_inv_b1_2_0 (.A(imd_Y1),.Y(Y1));
NANDC2x1 inst_clockedAND_b1_1 (.A(CLK),.B(Y1),.Y(imd_YF1));
INVC inst_clockedinv_b1_1 (.A(imd_YF1),.Y(YF1));


NANDC2x1 inst_and_b2_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire2_0_0));
INVC inst_inv_b2_0_0 (.A(imd_wire2_0_0),.Y(wire2_0_0));
NANDC2x1 inst_and_b2_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire2_0_1));
INVC inst_inv_b2_0_1 (.A(imd_wire2_0_1),.Y(wire2_0_1));
NANDC2x1 inst_and_b2_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire2_0_2));
INVC inst_inv_b2_0_2 (.A(imd_wire2_0_2),.Y(wire2_0_2));
NANDC2x1 inst_and_b2_1_0 (.A(wire2_0_0),.B(wire2_0_1),.Y(imd_wire2_1_0));
INVC inst_inv_b2_1_0 (.A(imd_wire2_1_0),.Y(wire2_1_0));
NANDC2x1 inst_and_b2_1_1 (.A(A6_inv),.B(wire2_0_2),.Y(imd_wire2_1_1));
INVC inst_inv_b2_1_1 (.A(imd_wire2_1_1),.Y(wire2_1_1));
NANDC2x1 inst_and_b2_2_0 (.A(wire2_1_0),.B(wire2_1_1),.Y(imd_Y2));
INVC inst_inv_b2_2_0 (.A(imd_Y2),.Y(Y2));
NANDC2x1 inst_clockedAND_b2_2 (.A(CLK),.B(Y2),.Y(imd_YF2));
INVC inst_clockedinv_b2_2 (.A(imd_YF2),.Y(YF2));


NANDC2x1 inst_and_b3_0_0 (.A(A0),.B(A1),.Y(imd_wire3_0_0));
INVC inst_inv_b3_0_0 (.A(imd_wire3_0_0),.Y(wire3_0_0));
NANDC2x1 inst_and_b3_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire3_0_1));
INVC inst_inv_b3_0_1 (.A(imd_wire3_0_1),.Y(wire3_0_1));
NANDC2x1 inst_and_b3_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire3_0_2));
INVC inst_inv_b3_0_2 (.A(imd_wire3_0_2),.Y(wire3_0_2));
NANDC2x1 inst_and_b3_1_0 (.A(wire3_0_0),.B(wire3_0_1),.Y(imd_wire3_1_0));
INVC inst_inv_b3_1_0 (.A(imd_wire3_1_0),.Y(wire3_1_0));
NANDC2x1 inst_and_b3_1_1 (.A(A6_inv),.B(wire3_0_2),.Y(imd_wire3_1_1));
INVC inst_inv_b3_1_1 (.A(imd_wire3_1_1),.Y(wire3_1_1));
NANDC2x1 inst_and_b3_2_0 (.A(wire3_1_0),.B(wire3_1_1),.Y(imd_Y3));
INVC inst_inv_b3_2_0 (.A(imd_Y3),.Y(Y3));
NANDC2x1 inst_clockedAND_b3_3 (.A(CLK),.B(Y3),.Y(imd_YF3));
INVC inst_clockedinv_b3_3 (.A(imd_YF3),.Y(YF3));


NANDC2x1 inst_and_b4_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire4_0_0));
INVC inst_inv_b4_0_0 (.A(imd_wire4_0_0),.Y(wire4_0_0));
NANDC2x1 inst_and_b4_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire4_0_1));
INVC inst_inv_b4_0_1 (.A(imd_wire4_0_1),.Y(wire4_0_1));
NANDC2x1 inst_and_b4_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire4_0_2));
INVC inst_inv_b4_0_2 (.A(imd_wire4_0_2),.Y(wire4_0_2));
NANDC2x1 inst_and_b4_1_0 (.A(wire4_0_0),.B(wire4_0_1),.Y(imd_wire4_1_0));
INVC inst_inv_b4_1_0 (.A(imd_wire4_1_0),.Y(wire4_1_0));
NANDC2x1 inst_and_b4_1_1 (.A(A6_inv),.B(wire4_0_2),.Y(imd_wire4_1_1));
INVC inst_inv_b4_1_1 (.A(imd_wire4_1_1),.Y(wire4_1_1));
NANDC2x1 inst_and_b4_2_0 (.A(wire4_1_0),.B(wire4_1_1),.Y(imd_Y4));
INVC inst_inv_b4_2_0 (.A(imd_Y4),.Y(Y4));
NANDC2x1 inst_clockedAND_b4_4 (.A(CLK),.B(Y4),.Y(imd_YF4));
INVC inst_clockedinv_b4_4 (.A(imd_YF4),.Y(YF4));


NANDC2x1 inst_and_b5_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire5_0_0));
INVC inst_inv_b5_0_0 (.A(imd_wire5_0_0),.Y(wire5_0_0));
NANDC2x1 inst_and_b5_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire5_0_1));
INVC inst_inv_b5_0_1 (.A(imd_wire5_0_1),.Y(wire5_0_1));
NANDC2x1 inst_and_b5_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire5_0_2));
INVC inst_inv_b5_0_2 (.A(imd_wire5_0_2),.Y(wire5_0_2));
NANDC2x1 inst_and_b5_1_0 (.A(wire5_0_0),.B(wire5_0_1),.Y(imd_wire5_1_0));
INVC inst_inv_b5_1_0 (.A(imd_wire5_1_0),.Y(wire5_1_0));
NANDC2x1 inst_and_b5_1_1 (.A(A6_inv),.B(wire5_0_2),.Y(imd_wire5_1_1));
INVC inst_inv_b5_1_1 (.A(imd_wire5_1_1),.Y(wire5_1_1));
NANDC2x1 inst_and_b5_2_0 (.A(wire5_1_0),.B(wire5_1_1),.Y(imd_Y5));
INVC inst_inv_b5_2_0 (.A(imd_Y5),.Y(Y5));
NANDC2x1 inst_clockedAND_b5_5 (.A(CLK),.B(Y5),.Y(imd_YF5));
INVC inst_clockedinv_b5_5 (.A(imd_YF5),.Y(YF5));


NANDC2x1 inst_and_b6_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire6_0_0));
INVC inst_inv_b6_0_0 (.A(imd_wire6_0_0),.Y(wire6_0_0));
NANDC2x1 inst_and_b6_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire6_0_1));
INVC inst_inv_b6_0_1 (.A(imd_wire6_0_1),.Y(wire6_0_1));
NANDC2x1 inst_and_b6_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire6_0_2));
INVC inst_inv_b6_0_2 (.A(imd_wire6_0_2),.Y(wire6_0_2));
NANDC2x1 inst_and_b6_1_0 (.A(wire6_0_0),.B(wire6_0_1),.Y(imd_wire6_1_0));
INVC inst_inv_b6_1_0 (.A(imd_wire6_1_0),.Y(wire6_1_0));
NANDC2x1 inst_and_b6_1_1 (.A(A6_inv),.B(wire6_0_2),.Y(imd_wire6_1_1));
INVC inst_inv_b6_1_1 (.A(imd_wire6_1_1),.Y(wire6_1_1));
NANDC2x1 inst_and_b6_2_0 (.A(wire6_1_0),.B(wire6_1_1),.Y(imd_Y6));
INVC inst_inv_b6_2_0 (.A(imd_Y6),.Y(Y6));
NANDC2x1 inst_clockedAND_b6_6 (.A(CLK),.B(Y6),.Y(imd_YF6));
INVC inst_clockedinv_b6_6 (.A(imd_YF6),.Y(YF6));


NANDC2x1 inst_and_b7_0_0 (.A(A0),.B(A1),.Y(imd_wire7_0_0));
INVC inst_inv_b7_0_0 (.A(imd_wire7_0_0),.Y(wire7_0_0));
NANDC2x1 inst_and_b7_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire7_0_1));
INVC inst_inv_b7_0_1 (.A(imd_wire7_0_1),.Y(wire7_0_1));
NANDC2x1 inst_and_b7_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire7_0_2));
INVC inst_inv_b7_0_2 (.A(imd_wire7_0_2),.Y(wire7_0_2));
NANDC2x1 inst_and_b7_1_0 (.A(wire7_0_0),.B(wire7_0_1),.Y(imd_wire7_1_0));
INVC inst_inv_b7_1_0 (.A(imd_wire7_1_0),.Y(wire7_1_0));
NANDC2x1 inst_and_b7_1_1 (.A(A6_inv),.B(wire7_0_2),.Y(imd_wire7_1_1));
INVC inst_inv_b7_1_1 (.A(imd_wire7_1_1),.Y(wire7_1_1));
NANDC2x1 inst_and_b7_2_0 (.A(wire7_1_0),.B(wire7_1_1),.Y(imd_Y7));
INVC inst_inv_b7_2_0 (.A(imd_Y7),.Y(Y7));
NANDC2x1 inst_clockedAND_b7_7 (.A(CLK),.B(Y7),.Y(imd_YF7));
INVC inst_clockedinv_b7_7 (.A(imd_YF7),.Y(YF7));


NANDC2x1 inst_and_b8_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire8_0_0));
INVC inst_inv_b8_0_0 (.A(imd_wire8_0_0),.Y(wire8_0_0));
NANDC2x1 inst_and_b8_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire8_0_1));
INVC inst_inv_b8_0_1 (.A(imd_wire8_0_1),.Y(wire8_0_1));
NANDC2x1 inst_and_b8_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire8_0_2));
INVC inst_inv_b8_0_2 (.A(imd_wire8_0_2),.Y(wire8_0_2));
NANDC2x1 inst_and_b8_1_0 (.A(wire8_0_0),.B(wire8_0_1),.Y(imd_wire8_1_0));
INVC inst_inv_b8_1_0 (.A(imd_wire8_1_0),.Y(wire8_1_0));
NANDC2x1 inst_and_b8_1_1 (.A(A6_inv),.B(wire8_0_2),.Y(imd_wire8_1_1));
INVC inst_inv_b8_1_1 (.A(imd_wire8_1_1),.Y(wire8_1_1));
NANDC2x1 inst_and_b8_2_0 (.A(wire8_1_0),.B(wire8_1_1),.Y(imd_Y8));
INVC inst_inv_b8_2_0 (.A(imd_Y8),.Y(Y8));
NANDC2x1 inst_clockedAND_b8_8 (.A(CLK),.B(Y8),.Y(imd_YF8));
INVC inst_clockedinv_b8_8 (.A(imd_YF8),.Y(YF8));


NANDC2x1 inst_and_b9_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire9_0_0));
INVC inst_inv_b9_0_0 (.A(imd_wire9_0_0),.Y(wire9_0_0));
NANDC2x1 inst_and_b9_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire9_0_1));
INVC inst_inv_b9_0_1 (.A(imd_wire9_0_1),.Y(wire9_0_1));
NANDC2x1 inst_and_b9_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire9_0_2));
INVC inst_inv_b9_0_2 (.A(imd_wire9_0_2),.Y(wire9_0_2));
NANDC2x1 inst_and_b9_1_0 (.A(wire9_0_0),.B(wire9_0_1),.Y(imd_wire9_1_0));
INVC inst_inv_b9_1_0 (.A(imd_wire9_1_0),.Y(wire9_1_0));
NANDC2x1 inst_and_b9_1_1 (.A(A6_inv),.B(wire9_0_2),.Y(imd_wire9_1_1));
INVC inst_inv_b9_1_1 (.A(imd_wire9_1_1),.Y(wire9_1_1));
NANDC2x1 inst_and_b9_2_0 (.A(wire9_1_0),.B(wire9_1_1),.Y(imd_Y9));
INVC inst_inv_b9_2_0 (.A(imd_Y9),.Y(Y9));
NANDC2x1 inst_clockedAND_b9_9 (.A(CLK),.B(Y9),.Y(imd_YF9));
INVC inst_clockedinv_b9_9 (.A(imd_YF9),.Y(YF9));


NANDC2x1 inst_and_b10_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire10_0_0));
INVC inst_inv_b10_0_0 (.A(imd_wire10_0_0),.Y(wire10_0_0));
NANDC2x1 inst_and_b10_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire10_0_1));
INVC inst_inv_b10_0_1 (.A(imd_wire10_0_1),.Y(wire10_0_1));
NANDC2x1 inst_and_b10_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire10_0_2));
INVC inst_inv_b10_0_2 (.A(imd_wire10_0_2),.Y(wire10_0_2));
NANDC2x1 inst_and_b10_1_0 (.A(wire10_0_0),.B(wire10_0_1),.Y(imd_wire10_1_0));
INVC inst_inv_b10_1_0 (.A(imd_wire10_1_0),.Y(wire10_1_0));
NANDC2x1 inst_and_b10_1_1 (.A(A6_inv),.B(wire10_0_2),.Y(imd_wire10_1_1));
INVC inst_inv_b10_1_1 (.A(imd_wire10_1_1),.Y(wire10_1_1));
NANDC2x1 inst_and_b10_2_0 (.A(wire10_1_0),.B(wire10_1_1),.Y(imd_Y10));
INVC inst_inv_b10_2_0 (.A(imd_Y10),.Y(Y10));
NANDC2x1 inst_clockedAND_b10_10 (.A(CLK),.B(Y10),.Y(imd_YF10));
INVC inst_clockedinv_b10_10 (.A(imd_YF10),.Y(YF10));


NANDC2x1 inst_and_b11_0_0 (.A(A0),.B(A1),.Y(imd_wire11_0_0));
INVC inst_inv_b11_0_0 (.A(imd_wire11_0_0),.Y(wire11_0_0));
NANDC2x1 inst_and_b11_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire11_0_1));
INVC inst_inv_b11_0_1 (.A(imd_wire11_0_1),.Y(wire11_0_1));
NANDC2x1 inst_and_b11_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire11_0_2));
INVC inst_inv_b11_0_2 (.A(imd_wire11_0_2),.Y(wire11_0_2));
NANDC2x1 inst_and_b11_1_0 (.A(wire11_0_0),.B(wire11_0_1),.Y(imd_wire11_1_0));
INVC inst_inv_b11_1_0 (.A(imd_wire11_1_0),.Y(wire11_1_0));
NANDC2x1 inst_and_b11_1_1 (.A(A6_inv),.B(wire11_0_2),.Y(imd_wire11_1_1));
INVC inst_inv_b11_1_1 (.A(imd_wire11_1_1),.Y(wire11_1_1));
NANDC2x1 inst_and_b11_2_0 (.A(wire11_1_0),.B(wire11_1_1),.Y(imd_Y11));
INVC inst_inv_b11_2_0 (.A(imd_Y11),.Y(Y11));
NANDC2x1 inst_clockedAND_b11_11 (.A(CLK),.B(Y11),.Y(imd_YF11));
INVC inst_clockedinv_b11_11 (.A(imd_YF11),.Y(YF11));


NANDC2x1 inst_and_b12_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire12_0_0));
INVC inst_inv_b12_0_0 (.A(imd_wire12_0_0),.Y(wire12_0_0));
NANDC2x1 inst_and_b12_0_1 (.A(A2),.B(A3),.Y(imd_wire12_0_1));
INVC inst_inv_b12_0_1 (.A(imd_wire12_0_1),.Y(wire12_0_1));
NANDC2x1 inst_and_b12_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire12_0_2));
INVC inst_inv_b12_0_2 (.A(imd_wire12_0_2),.Y(wire12_0_2));
NANDC2x1 inst_and_b12_1_0 (.A(wire12_0_0),.B(wire12_0_1),.Y(imd_wire12_1_0));
INVC inst_inv_b12_1_0 (.A(imd_wire12_1_0),.Y(wire12_1_0));
NANDC2x1 inst_and_b12_1_1 (.A(A6_inv),.B(wire12_0_2),.Y(imd_wire12_1_1));
INVC inst_inv_b12_1_1 (.A(imd_wire12_1_1),.Y(wire12_1_1));
NANDC2x1 inst_and_b12_2_0 (.A(wire12_1_0),.B(wire12_1_1),.Y(imd_Y12));
INVC inst_inv_b12_2_0 (.A(imd_Y12),.Y(Y12));
NANDC2x1 inst_clockedAND_b12_12 (.A(CLK),.B(Y12),.Y(imd_YF12));
INVC inst_clockedinv_b12_12 (.A(imd_YF12),.Y(YF12));


NANDC2x1 inst_and_b13_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire13_0_0));
INVC inst_inv_b13_0_0 (.A(imd_wire13_0_0),.Y(wire13_0_0));
NANDC2x1 inst_and_b13_0_1 (.A(A2),.B(A3),.Y(imd_wire13_0_1));
INVC inst_inv_b13_0_1 (.A(imd_wire13_0_1),.Y(wire13_0_1));
NANDC2x1 inst_and_b13_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire13_0_2));
INVC inst_inv_b13_0_2 (.A(imd_wire13_0_2),.Y(wire13_0_2));
NANDC2x1 inst_and_b13_1_0 (.A(wire13_0_0),.B(wire13_0_1),.Y(imd_wire13_1_0));
INVC inst_inv_b13_1_0 (.A(imd_wire13_1_0),.Y(wire13_1_0));
NANDC2x1 inst_and_b13_1_1 (.A(A6_inv),.B(wire13_0_2),.Y(imd_wire13_1_1));
INVC inst_inv_b13_1_1 (.A(imd_wire13_1_1),.Y(wire13_1_1));
NANDC2x1 inst_and_b13_2_0 (.A(wire13_1_0),.B(wire13_1_1),.Y(imd_Y13));
INVC inst_inv_b13_2_0 (.A(imd_Y13),.Y(Y13));
NANDC2x1 inst_clockedAND_b13_13 (.A(CLK),.B(Y13),.Y(imd_YF13));
INVC inst_clockedinv_b13_13 (.A(imd_YF13),.Y(YF13));


NANDC2x1 inst_and_b14_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire14_0_0));
INVC inst_inv_b14_0_0 (.A(imd_wire14_0_0),.Y(wire14_0_0));
NANDC2x1 inst_and_b14_0_1 (.A(A2),.B(A3),.Y(imd_wire14_0_1));
INVC inst_inv_b14_0_1 (.A(imd_wire14_0_1),.Y(wire14_0_1));
NANDC2x1 inst_and_b14_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire14_0_2));
INVC inst_inv_b14_0_2 (.A(imd_wire14_0_2),.Y(wire14_0_2));
NANDC2x1 inst_and_b14_1_0 (.A(wire14_0_0),.B(wire14_0_1),.Y(imd_wire14_1_0));
INVC inst_inv_b14_1_0 (.A(imd_wire14_1_0),.Y(wire14_1_0));
NANDC2x1 inst_and_b14_1_1 (.A(A6_inv),.B(wire14_0_2),.Y(imd_wire14_1_1));
INVC inst_inv_b14_1_1 (.A(imd_wire14_1_1),.Y(wire14_1_1));
NANDC2x1 inst_and_b14_2_0 (.A(wire14_1_0),.B(wire14_1_1),.Y(imd_Y14));
INVC inst_inv_b14_2_0 (.A(imd_Y14),.Y(Y14));
NANDC2x1 inst_clockedAND_b14_14 (.A(CLK),.B(Y14),.Y(imd_YF14));
INVC inst_clockedinv_b14_14 (.A(imd_YF14),.Y(YF14));


NANDC2x1 inst_and_b15_0_0 (.A(A0),.B(A1),.Y(imd_wire15_0_0));
INVC inst_inv_b15_0_0 (.A(imd_wire15_0_0),.Y(wire15_0_0));
NANDC2x1 inst_and_b15_0_1 (.A(A2),.B(A3),.Y(imd_wire15_0_1));
INVC inst_inv_b15_0_1 (.A(imd_wire15_0_1),.Y(wire15_0_1));
NANDC2x1 inst_and_b15_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire15_0_2));
INVC inst_inv_b15_0_2 (.A(imd_wire15_0_2),.Y(wire15_0_2));
NANDC2x1 inst_and_b15_1_0 (.A(wire15_0_0),.B(wire15_0_1),.Y(imd_wire15_1_0));
INVC inst_inv_b15_1_0 (.A(imd_wire15_1_0),.Y(wire15_1_0));
NANDC2x1 inst_and_b15_1_1 (.A(A6_inv),.B(wire15_0_2),.Y(imd_wire15_1_1));
INVC inst_inv_b15_1_1 (.A(imd_wire15_1_1),.Y(wire15_1_1));
NANDC2x1 inst_and_b15_2_0 (.A(wire15_1_0),.B(wire15_1_1),.Y(imd_Y15));
INVC inst_inv_b15_2_0 (.A(imd_Y15),.Y(Y15));
NANDC2x1 inst_clockedAND_b15_15 (.A(CLK),.B(Y15),.Y(imd_YF15));
INVC inst_clockedinv_b15_15 (.A(imd_YF15),.Y(YF15));


NANDC2x1 inst_and_b16_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire16_0_0));
INVC inst_inv_b16_0_0 (.A(imd_wire16_0_0),.Y(wire16_0_0));
NANDC2x1 inst_and_b16_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire16_0_1));
INVC inst_inv_b16_0_1 (.A(imd_wire16_0_1),.Y(wire16_0_1));
NANDC2x1 inst_and_b16_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire16_0_2));
INVC inst_inv_b16_0_2 (.A(imd_wire16_0_2),.Y(wire16_0_2));
NANDC2x1 inst_and_b16_1_0 (.A(wire16_0_0),.B(wire16_0_1),.Y(imd_wire16_1_0));
INVC inst_inv_b16_1_0 (.A(imd_wire16_1_0),.Y(wire16_1_0));
NANDC2x1 inst_and_b16_1_1 (.A(A6_inv),.B(wire16_0_2),.Y(imd_wire16_1_1));
INVC inst_inv_b16_1_1 (.A(imd_wire16_1_1),.Y(wire16_1_1));
NANDC2x1 inst_and_b16_2_0 (.A(wire16_1_0),.B(wire16_1_1),.Y(imd_Y16));
INVC inst_inv_b16_2_0 (.A(imd_Y16),.Y(Y16));
NANDC2x1 inst_clockedAND_b16_16 (.A(CLK),.B(Y16),.Y(imd_YF16));
INVC inst_clockedinv_b16_16 (.A(imd_YF16),.Y(YF16));


NANDC2x1 inst_and_b17_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire17_0_0));
INVC inst_inv_b17_0_0 (.A(imd_wire17_0_0),.Y(wire17_0_0));
NANDC2x1 inst_and_b17_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire17_0_1));
INVC inst_inv_b17_0_1 (.A(imd_wire17_0_1),.Y(wire17_0_1));
NANDC2x1 inst_and_b17_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire17_0_2));
INVC inst_inv_b17_0_2 (.A(imd_wire17_0_2),.Y(wire17_0_2));
NANDC2x1 inst_and_b17_1_0 (.A(wire17_0_0),.B(wire17_0_1),.Y(imd_wire17_1_0));
INVC inst_inv_b17_1_0 (.A(imd_wire17_1_0),.Y(wire17_1_0));
NANDC2x1 inst_and_b17_1_1 (.A(A6_inv),.B(wire17_0_2),.Y(imd_wire17_1_1));
INVC inst_inv_b17_1_1 (.A(imd_wire17_1_1),.Y(wire17_1_1));
NANDC2x1 inst_and_b17_2_0 (.A(wire17_1_0),.B(wire17_1_1),.Y(imd_Y17));
INVC inst_inv_b17_2_0 (.A(imd_Y17),.Y(Y17));
NANDC2x1 inst_clockedAND_b17_17 (.A(CLK),.B(Y17),.Y(imd_YF17));
INVC inst_clockedinv_b17_17 (.A(imd_YF17),.Y(YF17));


NANDC2x1 inst_and_b18_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire18_0_0));
INVC inst_inv_b18_0_0 (.A(imd_wire18_0_0),.Y(wire18_0_0));
NANDC2x1 inst_and_b18_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire18_0_1));
INVC inst_inv_b18_0_1 (.A(imd_wire18_0_1),.Y(wire18_0_1));
NANDC2x1 inst_and_b18_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire18_0_2));
INVC inst_inv_b18_0_2 (.A(imd_wire18_0_2),.Y(wire18_0_2));
NANDC2x1 inst_and_b18_1_0 (.A(wire18_0_0),.B(wire18_0_1),.Y(imd_wire18_1_0));
INVC inst_inv_b18_1_0 (.A(imd_wire18_1_0),.Y(wire18_1_0));
NANDC2x1 inst_and_b18_1_1 (.A(A6_inv),.B(wire18_0_2),.Y(imd_wire18_1_1));
INVC inst_inv_b18_1_1 (.A(imd_wire18_1_1),.Y(wire18_1_1));
NANDC2x1 inst_and_b18_2_0 (.A(wire18_1_0),.B(wire18_1_1),.Y(imd_Y18));
INVC inst_inv_b18_2_0 (.A(imd_Y18),.Y(Y18));
NANDC2x1 inst_clockedAND_b18_18 (.A(CLK),.B(Y18),.Y(imd_YF18));
INVC inst_clockedinv_b18_18 (.A(imd_YF18),.Y(YF18));


NANDC2x1 inst_and_b19_0_0 (.A(A0),.B(A1),.Y(imd_wire19_0_0));
INVC inst_inv_b19_0_0 (.A(imd_wire19_0_0),.Y(wire19_0_0));
NANDC2x1 inst_and_b19_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire19_0_1));
INVC inst_inv_b19_0_1 (.A(imd_wire19_0_1),.Y(wire19_0_1));
NANDC2x1 inst_and_b19_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire19_0_2));
INVC inst_inv_b19_0_2 (.A(imd_wire19_0_2),.Y(wire19_0_2));
NANDC2x1 inst_and_b19_1_0 (.A(wire19_0_0),.B(wire19_0_1),.Y(imd_wire19_1_0));
INVC inst_inv_b19_1_0 (.A(imd_wire19_1_0),.Y(wire19_1_0));
NANDC2x1 inst_and_b19_1_1 (.A(A6_inv),.B(wire19_0_2),.Y(imd_wire19_1_1));
INVC inst_inv_b19_1_1 (.A(imd_wire19_1_1),.Y(wire19_1_1));
NANDC2x1 inst_and_b19_2_0 (.A(wire19_1_0),.B(wire19_1_1),.Y(imd_Y19));
INVC inst_inv_b19_2_0 (.A(imd_Y19),.Y(Y19));
NANDC2x1 inst_clockedAND_b19_19 (.A(CLK),.B(Y19),.Y(imd_YF19));
INVC inst_clockedinv_b19_19 (.A(imd_YF19),.Y(YF19));


NANDC2x1 inst_and_b20_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire20_0_0));
INVC inst_inv_b20_0_0 (.A(imd_wire20_0_0),.Y(wire20_0_0));
NANDC2x1 inst_and_b20_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire20_0_1));
INVC inst_inv_b20_0_1 (.A(imd_wire20_0_1),.Y(wire20_0_1));
NANDC2x1 inst_and_b20_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire20_0_2));
INVC inst_inv_b20_0_2 (.A(imd_wire20_0_2),.Y(wire20_0_2));
NANDC2x1 inst_and_b20_1_0 (.A(wire20_0_0),.B(wire20_0_1),.Y(imd_wire20_1_0));
INVC inst_inv_b20_1_0 (.A(imd_wire20_1_0),.Y(wire20_1_0));
NANDC2x1 inst_and_b20_1_1 (.A(A6_inv),.B(wire20_0_2),.Y(imd_wire20_1_1));
INVC inst_inv_b20_1_1 (.A(imd_wire20_1_1),.Y(wire20_1_1));
NANDC2x1 inst_and_b20_2_0 (.A(wire20_1_0),.B(wire20_1_1),.Y(imd_Y20));
INVC inst_inv_b20_2_0 (.A(imd_Y20),.Y(Y20));
NANDC2x1 inst_clockedAND_b20_20 (.A(CLK),.B(Y20),.Y(imd_YF20));
INVC inst_clockedinv_b20_20 (.A(imd_YF20),.Y(YF20));


NANDC2x1 inst_and_b21_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire21_0_0));
INVC inst_inv_b21_0_0 (.A(imd_wire21_0_0),.Y(wire21_0_0));
NANDC2x1 inst_and_b21_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire21_0_1));
INVC inst_inv_b21_0_1 (.A(imd_wire21_0_1),.Y(wire21_0_1));
NANDC2x1 inst_and_b21_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire21_0_2));
INVC inst_inv_b21_0_2 (.A(imd_wire21_0_2),.Y(wire21_0_2));
NANDC2x1 inst_and_b21_1_0 (.A(wire21_0_0),.B(wire21_0_1),.Y(imd_wire21_1_0));
INVC inst_inv_b21_1_0 (.A(imd_wire21_1_0),.Y(wire21_1_0));
NANDC2x1 inst_and_b21_1_1 (.A(A6_inv),.B(wire21_0_2),.Y(imd_wire21_1_1));
INVC inst_inv_b21_1_1 (.A(imd_wire21_1_1),.Y(wire21_1_1));
NANDC2x1 inst_and_b21_2_0 (.A(wire21_1_0),.B(wire21_1_1),.Y(imd_Y21));
INVC inst_inv_b21_2_0 (.A(imd_Y21),.Y(Y21));
NANDC2x1 inst_clockedAND_b21_21 (.A(CLK),.B(Y21),.Y(imd_YF21));
INVC inst_clockedinv_b21_21 (.A(imd_YF21),.Y(YF21));


NANDC2x1 inst_and_b22_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire22_0_0));
INVC inst_inv_b22_0_0 (.A(imd_wire22_0_0),.Y(wire22_0_0));
NANDC2x1 inst_and_b22_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire22_0_1));
INVC inst_inv_b22_0_1 (.A(imd_wire22_0_1),.Y(wire22_0_1));
NANDC2x1 inst_and_b22_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire22_0_2));
INVC inst_inv_b22_0_2 (.A(imd_wire22_0_2),.Y(wire22_0_2));
NANDC2x1 inst_and_b22_1_0 (.A(wire22_0_0),.B(wire22_0_1),.Y(imd_wire22_1_0));
INVC inst_inv_b22_1_0 (.A(imd_wire22_1_0),.Y(wire22_1_0));
NANDC2x1 inst_and_b22_1_1 (.A(A6_inv),.B(wire22_0_2),.Y(imd_wire22_1_1));
INVC inst_inv_b22_1_1 (.A(imd_wire22_1_1),.Y(wire22_1_1));
NANDC2x1 inst_and_b22_2_0 (.A(wire22_1_0),.B(wire22_1_1),.Y(imd_Y22));
INVC inst_inv_b22_2_0 (.A(imd_Y22),.Y(Y22));
NANDC2x1 inst_clockedAND_b22_22 (.A(CLK),.B(Y22),.Y(imd_YF22));
INVC inst_clockedinv_b22_22 (.A(imd_YF22),.Y(YF22));


NANDC2x1 inst_and_b23_0_0 (.A(A0),.B(A1),.Y(imd_wire23_0_0));
INVC inst_inv_b23_0_0 (.A(imd_wire23_0_0),.Y(wire23_0_0));
NANDC2x1 inst_and_b23_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire23_0_1));
INVC inst_inv_b23_0_1 (.A(imd_wire23_0_1),.Y(wire23_0_1));
NANDC2x1 inst_and_b23_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire23_0_2));
INVC inst_inv_b23_0_2 (.A(imd_wire23_0_2),.Y(wire23_0_2));
NANDC2x1 inst_and_b23_1_0 (.A(wire23_0_0),.B(wire23_0_1),.Y(imd_wire23_1_0));
INVC inst_inv_b23_1_0 (.A(imd_wire23_1_0),.Y(wire23_1_0));
NANDC2x1 inst_and_b23_1_1 (.A(A6_inv),.B(wire23_0_2),.Y(imd_wire23_1_1));
INVC inst_inv_b23_1_1 (.A(imd_wire23_1_1),.Y(wire23_1_1));
NANDC2x1 inst_and_b23_2_0 (.A(wire23_1_0),.B(wire23_1_1),.Y(imd_Y23));
INVC inst_inv_b23_2_0 (.A(imd_Y23),.Y(Y23));
NANDC2x1 inst_clockedAND_b23_23 (.A(CLK),.B(Y23),.Y(imd_YF23));
INVC inst_clockedinv_b23_23 (.A(imd_YF23),.Y(YF23));


NANDC2x1 inst_and_b24_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire24_0_0));
INVC inst_inv_b24_0_0 (.A(imd_wire24_0_0),.Y(wire24_0_0));
NANDC2x1 inst_and_b24_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire24_0_1));
INVC inst_inv_b24_0_1 (.A(imd_wire24_0_1),.Y(wire24_0_1));
NANDC2x1 inst_and_b24_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire24_0_2));
INVC inst_inv_b24_0_2 (.A(imd_wire24_0_2),.Y(wire24_0_2));
NANDC2x1 inst_and_b24_1_0 (.A(wire24_0_0),.B(wire24_0_1),.Y(imd_wire24_1_0));
INVC inst_inv_b24_1_0 (.A(imd_wire24_1_0),.Y(wire24_1_0));
NANDC2x1 inst_and_b24_1_1 (.A(A6_inv),.B(wire24_0_2),.Y(imd_wire24_1_1));
INVC inst_inv_b24_1_1 (.A(imd_wire24_1_1),.Y(wire24_1_1));
NANDC2x1 inst_and_b24_2_0 (.A(wire24_1_0),.B(wire24_1_1),.Y(imd_Y24));
INVC inst_inv_b24_2_0 (.A(imd_Y24),.Y(Y24));
NANDC2x1 inst_clockedAND_b24_24 (.A(CLK),.B(Y24),.Y(imd_YF24));
INVC inst_clockedinv_b24_24 (.A(imd_YF24),.Y(YF24));


NANDC2x1 inst_and_b25_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire25_0_0));
INVC inst_inv_b25_0_0 (.A(imd_wire25_0_0),.Y(wire25_0_0));
NANDC2x1 inst_and_b25_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire25_0_1));
INVC inst_inv_b25_0_1 (.A(imd_wire25_0_1),.Y(wire25_0_1));
NANDC2x1 inst_and_b25_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire25_0_2));
INVC inst_inv_b25_0_2 (.A(imd_wire25_0_2),.Y(wire25_0_2));
NANDC2x1 inst_and_b25_1_0 (.A(wire25_0_0),.B(wire25_0_1),.Y(imd_wire25_1_0));
INVC inst_inv_b25_1_0 (.A(imd_wire25_1_0),.Y(wire25_1_0));
NANDC2x1 inst_and_b25_1_1 (.A(A6_inv),.B(wire25_0_2),.Y(imd_wire25_1_1));
INVC inst_inv_b25_1_1 (.A(imd_wire25_1_1),.Y(wire25_1_1));
NANDC2x1 inst_and_b25_2_0 (.A(wire25_1_0),.B(wire25_1_1),.Y(imd_Y25));
INVC inst_inv_b25_2_0 (.A(imd_Y25),.Y(Y25));
NANDC2x1 inst_clockedAND_b25_25 (.A(CLK),.B(Y25),.Y(imd_YF25));
INVC inst_clockedinv_b25_25 (.A(imd_YF25),.Y(YF25));


NANDC2x1 inst_and_b26_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire26_0_0));
INVC inst_inv_b26_0_0 (.A(imd_wire26_0_0),.Y(wire26_0_0));
NANDC2x1 inst_and_b26_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire26_0_1));
INVC inst_inv_b26_0_1 (.A(imd_wire26_0_1),.Y(wire26_0_1));
NANDC2x1 inst_and_b26_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire26_0_2));
INVC inst_inv_b26_0_2 (.A(imd_wire26_0_2),.Y(wire26_0_2));
NANDC2x1 inst_and_b26_1_0 (.A(wire26_0_0),.B(wire26_0_1),.Y(imd_wire26_1_0));
INVC inst_inv_b26_1_0 (.A(imd_wire26_1_0),.Y(wire26_1_0));
NANDC2x1 inst_and_b26_1_1 (.A(A6_inv),.B(wire26_0_2),.Y(imd_wire26_1_1));
INVC inst_inv_b26_1_1 (.A(imd_wire26_1_1),.Y(wire26_1_1));
NANDC2x1 inst_and_b26_2_0 (.A(wire26_1_0),.B(wire26_1_1),.Y(imd_Y26));
INVC inst_inv_b26_2_0 (.A(imd_Y26),.Y(Y26));
NANDC2x1 inst_clockedAND_b26_26 (.A(CLK),.B(Y26),.Y(imd_YF26));
INVC inst_clockedinv_b26_26 (.A(imd_YF26),.Y(YF26));


NANDC2x1 inst_and_b27_0_0 (.A(A0),.B(A1),.Y(imd_wire27_0_0));
INVC inst_inv_b27_0_0 (.A(imd_wire27_0_0),.Y(wire27_0_0));
NANDC2x1 inst_and_b27_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire27_0_1));
INVC inst_inv_b27_0_1 (.A(imd_wire27_0_1),.Y(wire27_0_1));
NANDC2x1 inst_and_b27_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire27_0_2));
INVC inst_inv_b27_0_2 (.A(imd_wire27_0_2),.Y(wire27_0_2));
NANDC2x1 inst_and_b27_1_0 (.A(wire27_0_0),.B(wire27_0_1),.Y(imd_wire27_1_0));
INVC inst_inv_b27_1_0 (.A(imd_wire27_1_0),.Y(wire27_1_0));
NANDC2x1 inst_and_b27_1_1 (.A(A6_inv),.B(wire27_0_2),.Y(imd_wire27_1_1));
INVC inst_inv_b27_1_1 (.A(imd_wire27_1_1),.Y(wire27_1_1));
NANDC2x1 inst_and_b27_2_0 (.A(wire27_1_0),.B(wire27_1_1),.Y(imd_Y27));
INVC inst_inv_b27_2_0 (.A(imd_Y27),.Y(Y27));
NANDC2x1 inst_clockedAND_b27_27 (.A(CLK),.B(Y27),.Y(imd_YF27));
INVC inst_clockedinv_b27_27 (.A(imd_YF27),.Y(YF27));


NANDC2x1 inst_and_b28_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire28_0_0));
INVC inst_inv_b28_0_0 (.A(imd_wire28_0_0),.Y(wire28_0_0));
NANDC2x1 inst_and_b28_0_1 (.A(A2),.B(A3),.Y(imd_wire28_0_1));
INVC inst_inv_b28_0_1 (.A(imd_wire28_0_1),.Y(wire28_0_1));
NANDC2x1 inst_and_b28_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire28_0_2));
INVC inst_inv_b28_0_2 (.A(imd_wire28_0_2),.Y(wire28_0_2));
NANDC2x1 inst_and_b28_1_0 (.A(wire28_0_0),.B(wire28_0_1),.Y(imd_wire28_1_0));
INVC inst_inv_b28_1_0 (.A(imd_wire28_1_0),.Y(wire28_1_0));
NANDC2x1 inst_and_b28_1_1 (.A(A6_inv),.B(wire28_0_2),.Y(imd_wire28_1_1));
INVC inst_inv_b28_1_1 (.A(imd_wire28_1_1),.Y(wire28_1_1));
NANDC2x1 inst_and_b28_2_0 (.A(wire28_1_0),.B(wire28_1_1),.Y(imd_Y28));
INVC inst_inv_b28_2_0 (.A(imd_Y28),.Y(Y28));
NANDC2x1 inst_clockedAND_b28_28 (.A(CLK),.B(Y28),.Y(imd_YF28));
INVC inst_clockedinv_b28_28 (.A(imd_YF28),.Y(YF28));


NANDC2x1 inst_and_b29_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire29_0_0));
INVC inst_inv_b29_0_0 (.A(imd_wire29_0_0),.Y(wire29_0_0));
NANDC2x1 inst_and_b29_0_1 (.A(A2),.B(A3),.Y(imd_wire29_0_1));
INVC inst_inv_b29_0_1 (.A(imd_wire29_0_1),.Y(wire29_0_1));
NANDC2x1 inst_and_b29_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire29_0_2));
INVC inst_inv_b29_0_2 (.A(imd_wire29_0_2),.Y(wire29_0_2));
NANDC2x1 inst_and_b29_1_0 (.A(wire29_0_0),.B(wire29_0_1),.Y(imd_wire29_1_0));
INVC inst_inv_b29_1_0 (.A(imd_wire29_1_0),.Y(wire29_1_0));
NANDC2x1 inst_and_b29_1_1 (.A(A6_inv),.B(wire29_0_2),.Y(imd_wire29_1_1));
INVC inst_inv_b29_1_1 (.A(imd_wire29_1_1),.Y(wire29_1_1));
NANDC2x1 inst_and_b29_2_0 (.A(wire29_1_0),.B(wire29_1_1),.Y(imd_Y29));
INVC inst_inv_b29_2_0 (.A(imd_Y29),.Y(Y29));
NANDC2x1 inst_clockedAND_b29_29 (.A(CLK),.B(Y29),.Y(imd_YF29));
INVC inst_clockedinv_b29_29 (.A(imd_YF29),.Y(YF29));


NANDC2x1 inst_and_b30_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire30_0_0));
INVC inst_inv_b30_0_0 (.A(imd_wire30_0_0),.Y(wire30_0_0));
NANDC2x1 inst_and_b30_0_1 (.A(A2),.B(A3),.Y(imd_wire30_0_1));
INVC inst_inv_b30_0_1 (.A(imd_wire30_0_1),.Y(wire30_0_1));
NANDC2x1 inst_and_b30_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire30_0_2));
INVC inst_inv_b30_0_2 (.A(imd_wire30_0_2),.Y(wire30_0_2));
NANDC2x1 inst_and_b30_1_0 (.A(wire30_0_0),.B(wire30_0_1),.Y(imd_wire30_1_0));
INVC inst_inv_b30_1_0 (.A(imd_wire30_1_0),.Y(wire30_1_0));
NANDC2x1 inst_and_b30_1_1 (.A(A6_inv),.B(wire30_0_2),.Y(imd_wire30_1_1));
INVC inst_inv_b30_1_1 (.A(imd_wire30_1_1),.Y(wire30_1_1));
NANDC2x1 inst_and_b30_2_0 (.A(wire30_1_0),.B(wire30_1_1),.Y(imd_Y30));
INVC inst_inv_b30_2_0 (.A(imd_Y30),.Y(Y30));
NANDC2x1 inst_clockedAND_b30_30 (.A(CLK),.B(Y30),.Y(imd_YF30));
INVC inst_clockedinv_b30_30 (.A(imd_YF30),.Y(YF30));


NANDC2x1 inst_and_b31_0_0 (.A(A0),.B(A1),.Y(imd_wire31_0_0));
INVC inst_inv_b31_0_0 (.A(imd_wire31_0_0),.Y(wire31_0_0));
NANDC2x1 inst_and_b31_0_1 (.A(A2),.B(A3),.Y(imd_wire31_0_1));
INVC inst_inv_b31_0_1 (.A(imd_wire31_0_1),.Y(wire31_0_1));
NANDC2x1 inst_and_b31_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire31_0_2));
INVC inst_inv_b31_0_2 (.A(imd_wire31_0_2),.Y(wire31_0_2));
NANDC2x1 inst_and_b31_1_0 (.A(wire31_0_0),.B(wire31_0_1),.Y(imd_wire31_1_0));
INVC inst_inv_b31_1_0 (.A(imd_wire31_1_0),.Y(wire31_1_0));
NANDC2x1 inst_and_b31_1_1 (.A(A6_inv),.B(wire31_0_2),.Y(imd_wire31_1_1));
INVC inst_inv_b31_1_1 (.A(imd_wire31_1_1),.Y(wire31_1_1));
NANDC2x1 inst_and_b31_2_0 (.A(wire31_1_0),.B(wire31_1_1),.Y(imd_Y31));
INVC inst_inv_b31_2_0 (.A(imd_Y31),.Y(Y31));
NANDC2x1 inst_clockedAND_b31_31 (.A(CLK),.B(Y31),.Y(imd_YF31));
INVC inst_clockedinv_b31_31 (.A(imd_YF31),.Y(YF31));


NANDC2x1 inst_and_b32_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire32_0_0));
INVC inst_inv_b32_0_0 (.A(imd_wire32_0_0),.Y(wire32_0_0));
NANDC2x1 inst_and_b32_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire32_0_1));
INVC inst_inv_b32_0_1 (.A(imd_wire32_0_1),.Y(wire32_0_1));
NANDC2x1 inst_and_b32_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire32_0_2));
INVC inst_inv_b32_0_2 (.A(imd_wire32_0_2),.Y(wire32_0_2));
NANDC2x1 inst_and_b32_1_0 (.A(wire32_0_0),.B(wire32_0_1),.Y(imd_wire32_1_0));
INVC inst_inv_b32_1_0 (.A(imd_wire32_1_0),.Y(wire32_1_0));
NANDC2x1 inst_and_b32_1_1 (.A(A6_inv),.B(wire32_0_2),.Y(imd_wire32_1_1));
INVC inst_inv_b32_1_1 (.A(imd_wire32_1_1),.Y(wire32_1_1));
NANDC2x1 inst_and_b32_2_0 (.A(wire32_1_0),.B(wire32_1_1),.Y(imd_Y32));
INVC inst_inv_b32_2_0 (.A(imd_Y32),.Y(Y32));
NANDC2x1 inst_clockedAND_b32_32 (.A(CLK),.B(Y32),.Y(imd_YF32));
INVC inst_clockedinv_b32_32 (.A(imd_YF32),.Y(YF32));


NANDC2x1 inst_and_b33_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire33_0_0));
INVC inst_inv_b33_0_0 (.A(imd_wire33_0_0),.Y(wire33_0_0));
NANDC2x1 inst_and_b33_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire33_0_1));
INVC inst_inv_b33_0_1 (.A(imd_wire33_0_1),.Y(wire33_0_1));
NANDC2x1 inst_and_b33_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire33_0_2));
INVC inst_inv_b33_0_2 (.A(imd_wire33_0_2),.Y(wire33_0_2));
NANDC2x1 inst_and_b33_1_0 (.A(wire33_0_0),.B(wire33_0_1),.Y(imd_wire33_1_0));
INVC inst_inv_b33_1_0 (.A(imd_wire33_1_0),.Y(wire33_1_0));
NANDC2x1 inst_and_b33_1_1 (.A(A6_inv),.B(wire33_0_2),.Y(imd_wire33_1_1));
INVC inst_inv_b33_1_1 (.A(imd_wire33_1_1),.Y(wire33_1_1));
NANDC2x1 inst_and_b33_2_0 (.A(wire33_1_0),.B(wire33_1_1),.Y(imd_Y33));
INVC inst_inv_b33_2_0 (.A(imd_Y33),.Y(Y33));
NANDC2x1 inst_clockedAND_b33_33 (.A(CLK),.B(Y33),.Y(imd_YF33));
INVC inst_clockedinv_b33_33 (.A(imd_YF33),.Y(YF33));


NANDC2x1 inst_and_b34_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire34_0_0));
INVC inst_inv_b34_0_0 (.A(imd_wire34_0_0),.Y(wire34_0_0));
NANDC2x1 inst_and_b34_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire34_0_1));
INVC inst_inv_b34_0_1 (.A(imd_wire34_0_1),.Y(wire34_0_1));
NANDC2x1 inst_and_b34_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire34_0_2));
INVC inst_inv_b34_0_2 (.A(imd_wire34_0_2),.Y(wire34_0_2));
NANDC2x1 inst_and_b34_1_0 (.A(wire34_0_0),.B(wire34_0_1),.Y(imd_wire34_1_0));
INVC inst_inv_b34_1_0 (.A(imd_wire34_1_0),.Y(wire34_1_0));
NANDC2x1 inst_and_b34_1_1 (.A(A6_inv),.B(wire34_0_2),.Y(imd_wire34_1_1));
INVC inst_inv_b34_1_1 (.A(imd_wire34_1_1),.Y(wire34_1_1));
NANDC2x1 inst_and_b34_2_0 (.A(wire34_1_0),.B(wire34_1_1),.Y(imd_Y34));
INVC inst_inv_b34_2_0 (.A(imd_Y34),.Y(Y34));
NANDC2x1 inst_clockedAND_b34_34 (.A(CLK),.B(Y34),.Y(imd_YF34));
INVC inst_clockedinv_b34_34 (.A(imd_YF34),.Y(YF34));


NANDC2x1 inst_and_b35_0_0 (.A(A0),.B(A1),.Y(imd_wire35_0_0));
INVC inst_inv_b35_0_0 (.A(imd_wire35_0_0),.Y(wire35_0_0));
NANDC2x1 inst_and_b35_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire35_0_1));
INVC inst_inv_b35_0_1 (.A(imd_wire35_0_1),.Y(wire35_0_1));
NANDC2x1 inst_and_b35_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire35_0_2));
INVC inst_inv_b35_0_2 (.A(imd_wire35_0_2),.Y(wire35_0_2));
NANDC2x1 inst_and_b35_1_0 (.A(wire35_0_0),.B(wire35_0_1),.Y(imd_wire35_1_0));
INVC inst_inv_b35_1_0 (.A(imd_wire35_1_0),.Y(wire35_1_0));
NANDC2x1 inst_and_b35_1_1 (.A(A6_inv),.B(wire35_0_2),.Y(imd_wire35_1_1));
INVC inst_inv_b35_1_1 (.A(imd_wire35_1_1),.Y(wire35_1_1));
NANDC2x1 inst_and_b35_2_0 (.A(wire35_1_0),.B(wire35_1_1),.Y(imd_Y35));
INVC inst_inv_b35_2_0 (.A(imd_Y35),.Y(Y35));
NANDC2x1 inst_clockedAND_b35_35 (.A(CLK),.B(Y35),.Y(imd_YF35));
INVC inst_clockedinv_b35_35 (.A(imd_YF35),.Y(YF35));


NANDC2x1 inst_and_b36_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire36_0_0));
INVC inst_inv_b36_0_0 (.A(imd_wire36_0_0),.Y(wire36_0_0));
NANDC2x1 inst_and_b36_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire36_0_1));
INVC inst_inv_b36_0_1 (.A(imd_wire36_0_1),.Y(wire36_0_1));
NANDC2x1 inst_and_b36_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire36_0_2));
INVC inst_inv_b36_0_2 (.A(imd_wire36_0_2),.Y(wire36_0_2));
NANDC2x1 inst_and_b36_1_0 (.A(wire36_0_0),.B(wire36_0_1),.Y(imd_wire36_1_0));
INVC inst_inv_b36_1_0 (.A(imd_wire36_1_0),.Y(wire36_1_0));
NANDC2x1 inst_and_b36_1_1 (.A(A6_inv),.B(wire36_0_2),.Y(imd_wire36_1_1));
INVC inst_inv_b36_1_1 (.A(imd_wire36_1_1),.Y(wire36_1_1));
NANDC2x1 inst_and_b36_2_0 (.A(wire36_1_0),.B(wire36_1_1),.Y(imd_Y36));
INVC inst_inv_b36_2_0 (.A(imd_Y36),.Y(Y36));
NANDC2x1 inst_clockedAND_b36_36 (.A(CLK),.B(Y36),.Y(imd_YF36));
INVC inst_clockedinv_b36_36 (.A(imd_YF36),.Y(YF36));


NANDC2x1 inst_and_b37_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire37_0_0));
INVC inst_inv_b37_0_0 (.A(imd_wire37_0_0),.Y(wire37_0_0));
NANDC2x1 inst_and_b37_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire37_0_1));
INVC inst_inv_b37_0_1 (.A(imd_wire37_0_1),.Y(wire37_0_1));
NANDC2x1 inst_and_b37_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire37_0_2));
INVC inst_inv_b37_0_2 (.A(imd_wire37_0_2),.Y(wire37_0_2));
NANDC2x1 inst_and_b37_1_0 (.A(wire37_0_0),.B(wire37_0_1),.Y(imd_wire37_1_0));
INVC inst_inv_b37_1_0 (.A(imd_wire37_1_0),.Y(wire37_1_0));
NANDC2x1 inst_and_b37_1_1 (.A(A6_inv),.B(wire37_0_2),.Y(imd_wire37_1_1));
INVC inst_inv_b37_1_1 (.A(imd_wire37_1_1),.Y(wire37_1_1));
NANDC2x1 inst_and_b37_2_0 (.A(wire37_1_0),.B(wire37_1_1),.Y(imd_Y37));
INVC inst_inv_b37_2_0 (.A(imd_Y37),.Y(Y37));
NANDC2x1 inst_clockedAND_b37_37 (.A(CLK),.B(Y37),.Y(imd_YF37));
INVC inst_clockedinv_b37_37 (.A(imd_YF37),.Y(YF37));


NANDC2x1 inst_and_b38_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire38_0_0));
INVC inst_inv_b38_0_0 (.A(imd_wire38_0_0),.Y(wire38_0_0));
NANDC2x1 inst_and_b38_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire38_0_1));
INVC inst_inv_b38_0_1 (.A(imd_wire38_0_1),.Y(wire38_0_1));
NANDC2x1 inst_and_b38_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire38_0_2));
INVC inst_inv_b38_0_2 (.A(imd_wire38_0_2),.Y(wire38_0_2));
NANDC2x1 inst_and_b38_1_0 (.A(wire38_0_0),.B(wire38_0_1),.Y(imd_wire38_1_0));
INVC inst_inv_b38_1_0 (.A(imd_wire38_1_0),.Y(wire38_1_0));
NANDC2x1 inst_and_b38_1_1 (.A(A6_inv),.B(wire38_0_2),.Y(imd_wire38_1_1));
INVC inst_inv_b38_1_1 (.A(imd_wire38_1_1),.Y(wire38_1_1));
NANDC2x1 inst_and_b38_2_0 (.A(wire38_1_0),.B(wire38_1_1),.Y(imd_Y38));
INVC inst_inv_b38_2_0 (.A(imd_Y38),.Y(Y38));
NANDC2x1 inst_clockedAND_b38_38 (.A(CLK),.B(Y38),.Y(imd_YF38));
INVC inst_clockedinv_b38_38 (.A(imd_YF38),.Y(YF38));


NANDC2x1 inst_and_b39_0_0 (.A(A0),.B(A1),.Y(imd_wire39_0_0));
INVC inst_inv_b39_0_0 (.A(imd_wire39_0_0),.Y(wire39_0_0));
NANDC2x1 inst_and_b39_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire39_0_1));
INVC inst_inv_b39_0_1 (.A(imd_wire39_0_1),.Y(wire39_0_1));
NANDC2x1 inst_and_b39_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire39_0_2));
INVC inst_inv_b39_0_2 (.A(imd_wire39_0_2),.Y(wire39_0_2));
NANDC2x1 inst_and_b39_1_0 (.A(wire39_0_0),.B(wire39_0_1),.Y(imd_wire39_1_0));
INVC inst_inv_b39_1_0 (.A(imd_wire39_1_0),.Y(wire39_1_0));
NANDC2x1 inst_and_b39_1_1 (.A(A6_inv),.B(wire39_0_2),.Y(imd_wire39_1_1));
INVC inst_inv_b39_1_1 (.A(imd_wire39_1_1),.Y(wire39_1_1));
NANDC2x1 inst_and_b39_2_0 (.A(wire39_1_0),.B(wire39_1_1),.Y(imd_Y39));
INVC inst_inv_b39_2_0 (.A(imd_Y39),.Y(Y39));
NANDC2x1 inst_clockedAND_b39_39 (.A(CLK),.B(Y39),.Y(imd_YF39));
INVC inst_clockedinv_b39_39 (.A(imd_YF39),.Y(YF39));


NANDC2x1 inst_and_b40_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire40_0_0));
INVC inst_inv_b40_0_0 (.A(imd_wire40_0_0),.Y(wire40_0_0));
NANDC2x1 inst_and_b40_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire40_0_1));
INVC inst_inv_b40_0_1 (.A(imd_wire40_0_1),.Y(wire40_0_1));
NANDC2x1 inst_and_b40_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire40_0_2));
INVC inst_inv_b40_0_2 (.A(imd_wire40_0_2),.Y(wire40_0_2));
NANDC2x1 inst_and_b40_1_0 (.A(wire40_0_0),.B(wire40_0_1),.Y(imd_wire40_1_0));
INVC inst_inv_b40_1_0 (.A(imd_wire40_1_0),.Y(wire40_1_0));
NANDC2x1 inst_and_b40_1_1 (.A(A6_inv),.B(wire40_0_2),.Y(imd_wire40_1_1));
INVC inst_inv_b40_1_1 (.A(imd_wire40_1_1),.Y(wire40_1_1));
NANDC2x1 inst_and_b40_2_0 (.A(wire40_1_0),.B(wire40_1_1),.Y(imd_Y40));
INVC inst_inv_b40_2_0 (.A(imd_Y40),.Y(Y40));
NANDC2x1 inst_clockedAND_b40_40 (.A(CLK),.B(Y40),.Y(imd_YF40));
INVC inst_clockedinv_b40_40 (.A(imd_YF40),.Y(YF40));


NANDC2x1 inst_and_b41_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire41_0_0));
INVC inst_inv_b41_0_0 (.A(imd_wire41_0_0),.Y(wire41_0_0));
NANDC2x1 inst_and_b41_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire41_0_1));
INVC inst_inv_b41_0_1 (.A(imd_wire41_0_1),.Y(wire41_0_1));
NANDC2x1 inst_and_b41_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire41_0_2));
INVC inst_inv_b41_0_2 (.A(imd_wire41_0_2),.Y(wire41_0_2));
NANDC2x1 inst_and_b41_1_0 (.A(wire41_0_0),.B(wire41_0_1),.Y(imd_wire41_1_0));
INVC inst_inv_b41_1_0 (.A(imd_wire41_1_0),.Y(wire41_1_0));
NANDC2x1 inst_and_b41_1_1 (.A(A6_inv),.B(wire41_0_2),.Y(imd_wire41_1_1));
INVC inst_inv_b41_1_1 (.A(imd_wire41_1_1),.Y(wire41_1_1));
NANDC2x1 inst_and_b41_2_0 (.A(wire41_1_0),.B(wire41_1_1),.Y(imd_Y41));
INVC inst_inv_b41_2_0 (.A(imd_Y41),.Y(Y41));
NANDC2x1 inst_clockedAND_b41_41 (.A(CLK),.B(Y41),.Y(imd_YF41));
INVC inst_clockedinv_b41_41 (.A(imd_YF41),.Y(YF41));


NANDC2x1 inst_and_b42_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire42_0_0));
INVC inst_inv_b42_0_0 (.A(imd_wire42_0_0),.Y(wire42_0_0));
NANDC2x1 inst_and_b42_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire42_0_1));
INVC inst_inv_b42_0_1 (.A(imd_wire42_0_1),.Y(wire42_0_1));
NANDC2x1 inst_and_b42_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire42_0_2));
INVC inst_inv_b42_0_2 (.A(imd_wire42_0_2),.Y(wire42_0_2));
NANDC2x1 inst_and_b42_1_0 (.A(wire42_0_0),.B(wire42_0_1),.Y(imd_wire42_1_0));
INVC inst_inv_b42_1_0 (.A(imd_wire42_1_0),.Y(wire42_1_0));
NANDC2x1 inst_and_b42_1_1 (.A(A6_inv),.B(wire42_0_2),.Y(imd_wire42_1_1));
INVC inst_inv_b42_1_1 (.A(imd_wire42_1_1),.Y(wire42_1_1));
NANDC2x1 inst_and_b42_2_0 (.A(wire42_1_0),.B(wire42_1_1),.Y(imd_Y42));
INVC inst_inv_b42_2_0 (.A(imd_Y42),.Y(Y42));
NANDC2x1 inst_clockedAND_b42_42 (.A(CLK),.B(Y42),.Y(imd_YF42));
INVC inst_clockedinv_b42_42 (.A(imd_YF42),.Y(YF42));


NANDC2x1 inst_and_b43_0_0 (.A(A0),.B(A1),.Y(imd_wire43_0_0));
INVC inst_inv_b43_0_0 (.A(imd_wire43_0_0),.Y(wire43_0_0));
NANDC2x1 inst_and_b43_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire43_0_1));
INVC inst_inv_b43_0_1 (.A(imd_wire43_0_1),.Y(wire43_0_1));
NANDC2x1 inst_and_b43_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire43_0_2));
INVC inst_inv_b43_0_2 (.A(imd_wire43_0_2),.Y(wire43_0_2));
NANDC2x1 inst_and_b43_1_0 (.A(wire43_0_0),.B(wire43_0_1),.Y(imd_wire43_1_0));
INVC inst_inv_b43_1_0 (.A(imd_wire43_1_0),.Y(wire43_1_0));
NANDC2x1 inst_and_b43_1_1 (.A(A6_inv),.B(wire43_0_2),.Y(imd_wire43_1_1));
INVC inst_inv_b43_1_1 (.A(imd_wire43_1_1),.Y(wire43_1_1));
NANDC2x1 inst_and_b43_2_0 (.A(wire43_1_0),.B(wire43_1_1),.Y(imd_Y43));
INVC inst_inv_b43_2_0 (.A(imd_Y43),.Y(Y43));
NANDC2x1 inst_clockedAND_b43_43 (.A(CLK),.B(Y43),.Y(imd_YF43));
INVC inst_clockedinv_b43_43 (.A(imd_YF43),.Y(YF43));


NANDC2x1 inst_and_b44_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire44_0_0));
INVC inst_inv_b44_0_0 (.A(imd_wire44_0_0),.Y(wire44_0_0));
NANDC2x1 inst_and_b44_0_1 (.A(A2),.B(A3),.Y(imd_wire44_0_1));
INVC inst_inv_b44_0_1 (.A(imd_wire44_0_1),.Y(wire44_0_1));
NANDC2x1 inst_and_b44_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire44_0_2));
INVC inst_inv_b44_0_2 (.A(imd_wire44_0_2),.Y(wire44_0_2));
NANDC2x1 inst_and_b44_1_0 (.A(wire44_0_0),.B(wire44_0_1),.Y(imd_wire44_1_0));
INVC inst_inv_b44_1_0 (.A(imd_wire44_1_0),.Y(wire44_1_0));
NANDC2x1 inst_and_b44_1_1 (.A(A6_inv),.B(wire44_0_2),.Y(imd_wire44_1_1));
INVC inst_inv_b44_1_1 (.A(imd_wire44_1_1),.Y(wire44_1_1));
NANDC2x1 inst_and_b44_2_0 (.A(wire44_1_0),.B(wire44_1_1),.Y(imd_Y44));
INVC inst_inv_b44_2_0 (.A(imd_Y44),.Y(Y44));
NANDC2x1 inst_clockedAND_b44_44 (.A(CLK),.B(Y44),.Y(imd_YF44));
INVC inst_clockedinv_b44_44 (.A(imd_YF44),.Y(YF44));


NANDC2x1 inst_and_b45_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire45_0_0));
INVC inst_inv_b45_0_0 (.A(imd_wire45_0_0),.Y(wire45_0_0));
NANDC2x1 inst_and_b45_0_1 (.A(A2),.B(A3),.Y(imd_wire45_0_1));
INVC inst_inv_b45_0_1 (.A(imd_wire45_0_1),.Y(wire45_0_1));
NANDC2x1 inst_and_b45_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire45_0_2));
INVC inst_inv_b45_0_2 (.A(imd_wire45_0_2),.Y(wire45_0_2));
NANDC2x1 inst_and_b45_1_0 (.A(wire45_0_0),.B(wire45_0_1),.Y(imd_wire45_1_0));
INVC inst_inv_b45_1_0 (.A(imd_wire45_1_0),.Y(wire45_1_0));
NANDC2x1 inst_and_b45_1_1 (.A(A6_inv),.B(wire45_0_2),.Y(imd_wire45_1_1));
INVC inst_inv_b45_1_1 (.A(imd_wire45_1_1),.Y(wire45_1_1));
NANDC2x1 inst_and_b45_2_0 (.A(wire45_1_0),.B(wire45_1_1),.Y(imd_Y45));
INVC inst_inv_b45_2_0 (.A(imd_Y45),.Y(Y45));
NANDC2x1 inst_clockedAND_b45_45 (.A(CLK),.B(Y45),.Y(imd_YF45));
INVC inst_clockedinv_b45_45 (.A(imd_YF45),.Y(YF45));


NANDC2x1 inst_and_b46_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire46_0_0));
INVC inst_inv_b46_0_0 (.A(imd_wire46_0_0),.Y(wire46_0_0));
NANDC2x1 inst_and_b46_0_1 (.A(A2),.B(A3),.Y(imd_wire46_0_1));
INVC inst_inv_b46_0_1 (.A(imd_wire46_0_1),.Y(wire46_0_1));
NANDC2x1 inst_and_b46_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire46_0_2));
INVC inst_inv_b46_0_2 (.A(imd_wire46_0_2),.Y(wire46_0_2));
NANDC2x1 inst_and_b46_1_0 (.A(wire46_0_0),.B(wire46_0_1),.Y(imd_wire46_1_0));
INVC inst_inv_b46_1_0 (.A(imd_wire46_1_0),.Y(wire46_1_0));
NANDC2x1 inst_and_b46_1_1 (.A(A6_inv),.B(wire46_0_2),.Y(imd_wire46_1_1));
INVC inst_inv_b46_1_1 (.A(imd_wire46_1_1),.Y(wire46_1_1));
NANDC2x1 inst_and_b46_2_0 (.A(wire46_1_0),.B(wire46_1_1),.Y(imd_Y46));
INVC inst_inv_b46_2_0 (.A(imd_Y46),.Y(Y46));
NANDC2x1 inst_clockedAND_b46_46 (.A(CLK),.B(Y46),.Y(imd_YF46));
INVC inst_clockedinv_b46_46 (.A(imd_YF46),.Y(YF46));


NANDC2x1 inst_and_b47_0_0 (.A(A0),.B(A1),.Y(imd_wire47_0_0));
INVC inst_inv_b47_0_0 (.A(imd_wire47_0_0),.Y(wire47_0_0));
NANDC2x1 inst_and_b47_0_1 (.A(A2),.B(A3),.Y(imd_wire47_0_1));
INVC inst_inv_b47_0_1 (.A(imd_wire47_0_1),.Y(wire47_0_1));
NANDC2x1 inst_and_b47_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire47_0_2));
INVC inst_inv_b47_0_2 (.A(imd_wire47_0_2),.Y(wire47_0_2));
NANDC2x1 inst_and_b47_1_0 (.A(wire47_0_0),.B(wire47_0_1),.Y(imd_wire47_1_0));
INVC inst_inv_b47_1_0 (.A(imd_wire47_1_0),.Y(wire47_1_0));
NANDC2x1 inst_and_b47_1_1 (.A(A6_inv),.B(wire47_0_2),.Y(imd_wire47_1_1));
INVC inst_inv_b47_1_1 (.A(imd_wire47_1_1),.Y(wire47_1_1));
NANDC2x1 inst_and_b47_2_0 (.A(wire47_1_0),.B(wire47_1_1),.Y(imd_Y47));
INVC inst_inv_b47_2_0 (.A(imd_Y47),.Y(Y47));
NANDC2x1 inst_clockedAND_b47_47 (.A(CLK),.B(Y47),.Y(imd_YF47));
INVC inst_clockedinv_b47_47 (.A(imd_YF47),.Y(YF47));


NANDC2x1 inst_and_b48_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire48_0_0));
INVC inst_inv_b48_0_0 (.A(imd_wire48_0_0),.Y(wire48_0_0));
NANDC2x1 inst_and_b48_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire48_0_1));
INVC inst_inv_b48_0_1 (.A(imd_wire48_0_1),.Y(wire48_0_1));
NANDC2x1 inst_and_b48_0_2 (.A(A4),.B(A5),.Y(imd_wire48_0_2));
INVC inst_inv_b48_0_2 (.A(imd_wire48_0_2),.Y(wire48_0_2));
NANDC2x1 inst_and_b48_1_0 (.A(wire48_0_0),.B(wire48_0_1),.Y(imd_wire48_1_0));
INVC inst_inv_b48_1_0 (.A(imd_wire48_1_0),.Y(wire48_1_0));
NANDC2x1 inst_and_b48_1_1 (.A(A6_inv),.B(wire48_0_2),.Y(imd_wire48_1_1));
INVC inst_inv_b48_1_1 (.A(imd_wire48_1_1),.Y(wire48_1_1));
NANDC2x1 inst_and_b48_2_0 (.A(wire48_1_0),.B(wire48_1_1),.Y(imd_Y48));
INVC inst_inv_b48_2_0 (.A(imd_Y48),.Y(Y48));
NANDC2x1 inst_clockedAND_b48_48 (.A(CLK),.B(Y48),.Y(imd_YF48));
INVC inst_clockedinv_b48_48 (.A(imd_YF48),.Y(YF48));


NANDC2x1 inst_and_b49_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire49_0_0));
INVC inst_inv_b49_0_0 (.A(imd_wire49_0_0),.Y(wire49_0_0));
NANDC2x1 inst_and_b49_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire49_0_1));
INVC inst_inv_b49_0_1 (.A(imd_wire49_0_1),.Y(wire49_0_1));
NANDC2x1 inst_and_b49_0_2 (.A(A4),.B(A5),.Y(imd_wire49_0_2));
INVC inst_inv_b49_0_2 (.A(imd_wire49_0_2),.Y(wire49_0_2));
NANDC2x1 inst_and_b49_1_0 (.A(wire49_0_0),.B(wire49_0_1),.Y(imd_wire49_1_0));
INVC inst_inv_b49_1_0 (.A(imd_wire49_1_0),.Y(wire49_1_0));
NANDC2x1 inst_and_b49_1_1 (.A(A6_inv),.B(wire49_0_2),.Y(imd_wire49_1_1));
INVC inst_inv_b49_1_1 (.A(imd_wire49_1_1),.Y(wire49_1_1));
NANDC2x1 inst_and_b49_2_0 (.A(wire49_1_0),.B(wire49_1_1),.Y(imd_Y49));
INVC inst_inv_b49_2_0 (.A(imd_Y49),.Y(Y49));
NANDC2x1 inst_clockedAND_b49_49 (.A(CLK),.B(Y49),.Y(imd_YF49));
INVC inst_clockedinv_b49_49 (.A(imd_YF49),.Y(YF49));


NANDC2x1 inst_and_b50_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire50_0_0));
INVC inst_inv_b50_0_0 (.A(imd_wire50_0_0),.Y(wire50_0_0));
NANDC2x1 inst_and_b50_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire50_0_1));
INVC inst_inv_b50_0_1 (.A(imd_wire50_0_1),.Y(wire50_0_1));
NANDC2x1 inst_and_b50_0_2 (.A(A4),.B(A5),.Y(imd_wire50_0_2));
INVC inst_inv_b50_0_2 (.A(imd_wire50_0_2),.Y(wire50_0_2));
NANDC2x1 inst_and_b50_1_0 (.A(wire50_0_0),.B(wire50_0_1),.Y(imd_wire50_1_0));
INVC inst_inv_b50_1_0 (.A(imd_wire50_1_0),.Y(wire50_1_0));
NANDC2x1 inst_and_b50_1_1 (.A(A6_inv),.B(wire50_0_2),.Y(imd_wire50_1_1));
INVC inst_inv_b50_1_1 (.A(imd_wire50_1_1),.Y(wire50_1_1));
NANDC2x1 inst_and_b50_2_0 (.A(wire50_1_0),.B(wire50_1_1),.Y(imd_Y50));
INVC inst_inv_b50_2_0 (.A(imd_Y50),.Y(Y50));
NANDC2x1 inst_clockedAND_b50_50 (.A(CLK),.B(Y50),.Y(imd_YF50));
INVC inst_clockedinv_b50_50 (.A(imd_YF50),.Y(YF50));


NANDC2x1 inst_and_b51_0_0 (.A(A0),.B(A1),.Y(imd_wire51_0_0));
INVC inst_inv_b51_0_0 (.A(imd_wire51_0_0),.Y(wire51_0_0));
NANDC2x1 inst_and_b51_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire51_0_1));
INVC inst_inv_b51_0_1 (.A(imd_wire51_0_1),.Y(wire51_0_1));
NANDC2x1 inst_and_b51_0_2 (.A(A4),.B(A5),.Y(imd_wire51_0_2));
INVC inst_inv_b51_0_2 (.A(imd_wire51_0_2),.Y(wire51_0_2));
NANDC2x1 inst_and_b51_1_0 (.A(wire51_0_0),.B(wire51_0_1),.Y(imd_wire51_1_0));
INVC inst_inv_b51_1_0 (.A(imd_wire51_1_0),.Y(wire51_1_0));
NANDC2x1 inst_and_b51_1_1 (.A(A6_inv),.B(wire51_0_2),.Y(imd_wire51_1_1));
INVC inst_inv_b51_1_1 (.A(imd_wire51_1_1),.Y(wire51_1_1));
NANDC2x1 inst_and_b51_2_0 (.A(wire51_1_0),.B(wire51_1_1),.Y(imd_Y51));
INVC inst_inv_b51_2_0 (.A(imd_Y51),.Y(Y51));
NANDC2x1 inst_clockedAND_b51_51 (.A(CLK),.B(Y51),.Y(imd_YF51));
INVC inst_clockedinv_b51_51 (.A(imd_YF51),.Y(YF51));


NANDC2x1 inst_and_b52_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire52_0_0));
INVC inst_inv_b52_0_0 (.A(imd_wire52_0_0),.Y(wire52_0_0));
NANDC2x1 inst_and_b52_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire52_0_1));
INVC inst_inv_b52_0_1 (.A(imd_wire52_0_1),.Y(wire52_0_1));
NANDC2x1 inst_and_b52_0_2 (.A(A4),.B(A5),.Y(imd_wire52_0_2));
INVC inst_inv_b52_0_2 (.A(imd_wire52_0_2),.Y(wire52_0_2));
NANDC2x1 inst_and_b52_1_0 (.A(wire52_0_0),.B(wire52_0_1),.Y(imd_wire52_1_0));
INVC inst_inv_b52_1_0 (.A(imd_wire52_1_0),.Y(wire52_1_0));
NANDC2x1 inst_and_b52_1_1 (.A(A6_inv),.B(wire52_0_2),.Y(imd_wire52_1_1));
INVC inst_inv_b52_1_1 (.A(imd_wire52_1_1),.Y(wire52_1_1));
NANDC2x1 inst_and_b52_2_0 (.A(wire52_1_0),.B(wire52_1_1),.Y(imd_Y52));
INVC inst_inv_b52_2_0 (.A(imd_Y52),.Y(Y52));
NANDC2x1 inst_clockedAND_b52_52 (.A(CLK),.B(Y52),.Y(imd_YF52));
INVC inst_clockedinv_b52_52 (.A(imd_YF52),.Y(YF52));


NANDC2x1 inst_and_b53_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire53_0_0));
INVC inst_inv_b53_0_0 (.A(imd_wire53_0_0),.Y(wire53_0_0));
NANDC2x1 inst_and_b53_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire53_0_1));
INVC inst_inv_b53_0_1 (.A(imd_wire53_0_1),.Y(wire53_0_1));
NANDC2x1 inst_and_b53_0_2 (.A(A4),.B(A5),.Y(imd_wire53_0_2));
INVC inst_inv_b53_0_2 (.A(imd_wire53_0_2),.Y(wire53_0_2));
NANDC2x1 inst_and_b53_1_0 (.A(wire53_0_0),.B(wire53_0_1),.Y(imd_wire53_1_0));
INVC inst_inv_b53_1_0 (.A(imd_wire53_1_0),.Y(wire53_1_0));
NANDC2x1 inst_and_b53_1_1 (.A(A6_inv),.B(wire53_0_2),.Y(imd_wire53_1_1));
INVC inst_inv_b53_1_1 (.A(imd_wire53_1_1),.Y(wire53_1_1));
NANDC2x1 inst_and_b53_2_0 (.A(wire53_1_0),.B(wire53_1_1),.Y(imd_Y53));
INVC inst_inv_b53_2_0 (.A(imd_Y53),.Y(Y53));
NANDC2x1 inst_clockedAND_b53_53 (.A(CLK),.B(Y53),.Y(imd_YF53));
INVC inst_clockedinv_b53_53 (.A(imd_YF53),.Y(YF53));


NANDC2x1 inst_and_b54_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire54_0_0));
INVC inst_inv_b54_0_0 (.A(imd_wire54_0_0),.Y(wire54_0_0));
NANDC2x1 inst_and_b54_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire54_0_1));
INVC inst_inv_b54_0_1 (.A(imd_wire54_0_1),.Y(wire54_0_1));
NANDC2x1 inst_and_b54_0_2 (.A(A4),.B(A5),.Y(imd_wire54_0_2));
INVC inst_inv_b54_0_2 (.A(imd_wire54_0_2),.Y(wire54_0_2));
NANDC2x1 inst_and_b54_1_0 (.A(wire54_0_0),.B(wire54_0_1),.Y(imd_wire54_1_0));
INVC inst_inv_b54_1_0 (.A(imd_wire54_1_0),.Y(wire54_1_0));
NANDC2x1 inst_and_b54_1_1 (.A(A6_inv),.B(wire54_0_2),.Y(imd_wire54_1_1));
INVC inst_inv_b54_1_1 (.A(imd_wire54_1_1),.Y(wire54_1_1));
NANDC2x1 inst_and_b54_2_0 (.A(wire54_1_0),.B(wire54_1_1),.Y(imd_Y54));
INVC inst_inv_b54_2_0 (.A(imd_Y54),.Y(Y54));
NANDC2x1 inst_clockedAND_b54_54 (.A(CLK),.B(Y54),.Y(imd_YF54));
INVC inst_clockedinv_b54_54 (.A(imd_YF54),.Y(YF54));


NANDC2x1 inst_and_b55_0_0 (.A(A0),.B(A1),.Y(imd_wire55_0_0));
INVC inst_inv_b55_0_0 (.A(imd_wire55_0_0),.Y(wire55_0_0));
NANDC2x1 inst_and_b55_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire55_0_1));
INVC inst_inv_b55_0_1 (.A(imd_wire55_0_1),.Y(wire55_0_1));
NANDC2x1 inst_and_b55_0_2 (.A(A4),.B(A5),.Y(imd_wire55_0_2));
INVC inst_inv_b55_0_2 (.A(imd_wire55_0_2),.Y(wire55_0_2));
NANDC2x1 inst_and_b55_1_0 (.A(wire55_0_0),.B(wire55_0_1),.Y(imd_wire55_1_0));
INVC inst_inv_b55_1_0 (.A(imd_wire55_1_0),.Y(wire55_1_0));
NANDC2x1 inst_and_b55_1_1 (.A(A6_inv),.B(wire55_0_2),.Y(imd_wire55_1_1));
INVC inst_inv_b55_1_1 (.A(imd_wire55_1_1),.Y(wire55_1_1));
NANDC2x1 inst_and_b55_2_0 (.A(wire55_1_0),.B(wire55_1_1),.Y(imd_Y55));
INVC inst_inv_b55_2_0 (.A(imd_Y55),.Y(Y55));
NANDC2x1 inst_clockedAND_b55_55 (.A(CLK),.B(Y55),.Y(imd_YF55));
INVC inst_clockedinv_b55_55 (.A(imd_YF55),.Y(YF55));


NANDC2x1 inst_and_b56_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire56_0_0));
INVC inst_inv_b56_0_0 (.A(imd_wire56_0_0),.Y(wire56_0_0));
NANDC2x1 inst_and_b56_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire56_0_1));
INVC inst_inv_b56_0_1 (.A(imd_wire56_0_1),.Y(wire56_0_1));
NANDC2x1 inst_and_b56_0_2 (.A(A4),.B(A5),.Y(imd_wire56_0_2));
INVC inst_inv_b56_0_2 (.A(imd_wire56_0_2),.Y(wire56_0_2));
NANDC2x1 inst_and_b56_1_0 (.A(wire56_0_0),.B(wire56_0_1),.Y(imd_wire56_1_0));
INVC inst_inv_b56_1_0 (.A(imd_wire56_1_0),.Y(wire56_1_0));
NANDC2x1 inst_and_b56_1_1 (.A(A6_inv),.B(wire56_0_2),.Y(imd_wire56_1_1));
INVC inst_inv_b56_1_1 (.A(imd_wire56_1_1),.Y(wire56_1_1));
NANDC2x1 inst_and_b56_2_0 (.A(wire56_1_0),.B(wire56_1_1),.Y(imd_Y56));
INVC inst_inv_b56_2_0 (.A(imd_Y56),.Y(Y56));
NANDC2x1 inst_clockedAND_b56_56 (.A(CLK),.B(Y56),.Y(imd_YF56));
INVC inst_clockedinv_b56_56 (.A(imd_YF56),.Y(YF56));


NANDC2x1 inst_and_b57_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire57_0_0));
INVC inst_inv_b57_0_0 (.A(imd_wire57_0_0),.Y(wire57_0_0));
NANDC2x1 inst_and_b57_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire57_0_1));
INVC inst_inv_b57_0_1 (.A(imd_wire57_0_1),.Y(wire57_0_1));
NANDC2x1 inst_and_b57_0_2 (.A(A4),.B(A5),.Y(imd_wire57_0_2));
INVC inst_inv_b57_0_2 (.A(imd_wire57_0_2),.Y(wire57_0_2));
NANDC2x1 inst_and_b57_1_0 (.A(wire57_0_0),.B(wire57_0_1),.Y(imd_wire57_1_0));
INVC inst_inv_b57_1_0 (.A(imd_wire57_1_0),.Y(wire57_1_0));
NANDC2x1 inst_and_b57_1_1 (.A(A6_inv),.B(wire57_0_2),.Y(imd_wire57_1_1));
INVC inst_inv_b57_1_1 (.A(imd_wire57_1_1),.Y(wire57_1_1));
NANDC2x1 inst_and_b57_2_0 (.A(wire57_1_0),.B(wire57_1_1),.Y(imd_Y57));
INVC inst_inv_b57_2_0 (.A(imd_Y57),.Y(Y57));
NANDC2x1 inst_clockedAND_b57_57 (.A(CLK),.B(Y57),.Y(imd_YF57));
INVC inst_clockedinv_b57_57 (.A(imd_YF57),.Y(YF57));


NANDC2x1 inst_and_b58_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire58_0_0));
INVC inst_inv_b58_0_0 (.A(imd_wire58_0_0),.Y(wire58_0_0));
NANDC2x1 inst_and_b58_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire58_0_1));
INVC inst_inv_b58_0_1 (.A(imd_wire58_0_1),.Y(wire58_0_1));
NANDC2x1 inst_and_b58_0_2 (.A(A4),.B(A5),.Y(imd_wire58_0_2));
INVC inst_inv_b58_0_2 (.A(imd_wire58_0_2),.Y(wire58_0_2));
NANDC2x1 inst_and_b58_1_0 (.A(wire58_0_0),.B(wire58_0_1),.Y(imd_wire58_1_0));
INVC inst_inv_b58_1_0 (.A(imd_wire58_1_0),.Y(wire58_1_0));
NANDC2x1 inst_and_b58_1_1 (.A(A6_inv),.B(wire58_0_2),.Y(imd_wire58_1_1));
INVC inst_inv_b58_1_1 (.A(imd_wire58_1_1),.Y(wire58_1_1));
NANDC2x1 inst_and_b58_2_0 (.A(wire58_1_0),.B(wire58_1_1),.Y(imd_Y58));
INVC inst_inv_b58_2_0 (.A(imd_Y58),.Y(Y58));
NANDC2x1 inst_clockedAND_b58_58 (.A(CLK),.B(Y58),.Y(imd_YF58));
INVC inst_clockedinv_b58_58 (.A(imd_YF58),.Y(YF58));


NANDC2x1 inst_and_b59_0_0 (.A(A0),.B(A1),.Y(imd_wire59_0_0));
INVC inst_inv_b59_0_0 (.A(imd_wire59_0_0),.Y(wire59_0_0));
NANDC2x1 inst_and_b59_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire59_0_1));
INVC inst_inv_b59_0_1 (.A(imd_wire59_0_1),.Y(wire59_0_1));
NANDC2x1 inst_and_b59_0_2 (.A(A4),.B(A5),.Y(imd_wire59_0_2));
INVC inst_inv_b59_0_2 (.A(imd_wire59_0_2),.Y(wire59_0_2));
NANDC2x1 inst_and_b59_1_0 (.A(wire59_0_0),.B(wire59_0_1),.Y(imd_wire59_1_0));
INVC inst_inv_b59_1_0 (.A(imd_wire59_1_0),.Y(wire59_1_0));
NANDC2x1 inst_and_b59_1_1 (.A(A6_inv),.B(wire59_0_2),.Y(imd_wire59_1_1));
INVC inst_inv_b59_1_1 (.A(imd_wire59_1_1),.Y(wire59_1_1));
NANDC2x1 inst_and_b59_2_0 (.A(wire59_1_0),.B(wire59_1_1),.Y(imd_Y59));
INVC inst_inv_b59_2_0 (.A(imd_Y59),.Y(Y59));
NANDC2x1 inst_clockedAND_b59_59 (.A(CLK),.B(Y59),.Y(imd_YF59));
INVC inst_clockedinv_b59_59 (.A(imd_YF59),.Y(YF59));


NANDC2x1 inst_and_b60_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire60_0_0));
INVC inst_inv_b60_0_0 (.A(imd_wire60_0_0),.Y(wire60_0_0));
NANDC2x1 inst_and_b60_0_1 (.A(A2),.B(A3),.Y(imd_wire60_0_1));
INVC inst_inv_b60_0_1 (.A(imd_wire60_0_1),.Y(wire60_0_1));
NANDC2x1 inst_and_b60_0_2 (.A(A4),.B(A5),.Y(imd_wire60_0_2));
INVC inst_inv_b60_0_2 (.A(imd_wire60_0_2),.Y(wire60_0_2));
NANDC2x1 inst_and_b60_1_0 (.A(wire60_0_0),.B(wire60_0_1),.Y(imd_wire60_1_0));
INVC inst_inv_b60_1_0 (.A(imd_wire60_1_0),.Y(wire60_1_0));
NANDC2x1 inst_and_b60_1_1 (.A(A6_inv),.B(wire60_0_2),.Y(imd_wire60_1_1));
INVC inst_inv_b60_1_1 (.A(imd_wire60_1_1),.Y(wire60_1_1));
NANDC2x1 inst_and_b60_2_0 (.A(wire60_1_0),.B(wire60_1_1),.Y(imd_Y60));
INVC inst_inv_b60_2_0 (.A(imd_Y60),.Y(Y60));
NANDC2x1 inst_clockedAND_b60_60 (.A(CLK),.B(Y60),.Y(imd_YF60));
INVC inst_clockedinv_b60_60 (.A(imd_YF60),.Y(YF60));


NANDC2x1 inst_and_b61_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire61_0_0));
INVC inst_inv_b61_0_0 (.A(imd_wire61_0_0),.Y(wire61_0_0));
NANDC2x1 inst_and_b61_0_1 (.A(A2),.B(A3),.Y(imd_wire61_0_1));
INVC inst_inv_b61_0_1 (.A(imd_wire61_0_1),.Y(wire61_0_1));
NANDC2x1 inst_and_b61_0_2 (.A(A4),.B(A5),.Y(imd_wire61_0_2));
INVC inst_inv_b61_0_2 (.A(imd_wire61_0_2),.Y(wire61_0_2));
NANDC2x1 inst_and_b61_1_0 (.A(wire61_0_0),.B(wire61_0_1),.Y(imd_wire61_1_0));
INVC inst_inv_b61_1_0 (.A(imd_wire61_1_0),.Y(wire61_1_0));
NANDC2x1 inst_and_b61_1_1 (.A(A6_inv),.B(wire61_0_2),.Y(imd_wire61_1_1));
INVC inst_inv_b61_1_1 (.A(imd_wire61_1_1),.Y(wire61_1_1));
NANDC2x1 inst_and_b61_2_0 (.A(wire61_1_0),.B(wire61_1_1),.Y(imd_Y61));
INVC inst_inv_b61_2_0 (.A(imd_Y61),.Y(Y61));
NANDC2x1 inst_clockedAND_b61_61 (.A(CLK),.B(Y61),.Y(imd_YF61));
INVC inst_clockedinv_b61_61 (.A(imd_YF61),.Y(YF61));


NANDC2x1 inst_and_b62_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire62_0_0));
INVC inst_inv_b62_0_0 (.A(imd_wire62_0_0),.Y(wire62_0_0));
NANDC2x1 inst_and_b62_0_1 (.A(A2),.B(A3),.Y(imd_wire62_0_1));
INVC inst_inv_b62_0_1 (.A(imd_wire62_0_1),.Y(wire62_0_1));
NANDC2x1 inst_and_b62_0_2 (.A(A4),.B(A5),.Y(imd_wire62_0_2));
INVC inst_inv_b62_0_2 (.A(imd_wire62_0_2),.Y(wire62_0_2));
NANDC2x1 inst_and_b62_1_0 (.A(wire62_0_0),.B(wire62_0_1),.Y(imd_wire62_1_0));
INVC inst_inv_b62_1_0 (.A(imd_wire62_1_0),.Y(wire62_1_0));
NANDC2x1 inst_and_b62_1_1 (.A(A6_inv),.B(wire62_0_2),.Y(imd_wire62_1_1));
INVC inst_inv_b62_1_1 (.A(imd_wire62_1_1),.Y(wire62_1_1));
NANDC2x1 inst_and_b62_2_0 (.A(wire62_1_0),.B(wire62_1_1),.Y(imd_Y62));
INVC inst_inv_b62_2_0 (.A(imd_Y62),.Y(Y62));
NANDC2x1 inst_clockedAND_b62_62 (.A(CLK),.B(Y62),.Y(imd_YF62));
INVC inst_clockedinv_b62_62 (.A(imd_YF62),.Y(YF62));


NANDC2x1 inst_and_b63_0_0 (.A(A0),.B(A1),.Y(imd_wire63_0_0));
INVC inst_inv_b63_0_0 (.A(imd_wire63_0_0),.Y(wire63_0_0));
NANDC2x1 inst_and_b63_0_1 (.A(A2),.B(A3),.Y(imd_wire63_0_1));
INVC inst_inv_b63_0_1 (.A(imd_wire63_0_1),.Y(wire63_0_1));
NANDC2x1 inst_and_b63_0_2 (.A(A4),.B(A5),.Y(imd_wire63_0_2));
INVC inst_inv_b63_0_2 (.A(imd_wire63_0_2),.Y(wire63_0_2));
NANDC2x1 inst_and_b63_1_0 (.A(wire63_0_0),.B(wire63_0_1),.Y(imd_wire63_1_0));
INVC inst_inv_b63_1_0 (.A(imd_wire63_1_0),.Y(wire63_1_0));
NANDC2x1 inst_and_b63_1_1 (.A(A6_inv),.B(wire63_0_2),.Y(imd_wire63_1_1));
INVC inst_inv_b63_1_1 (.A(imd_wire63_1_1),.Y(wire63_1_1));
NANDC2x1 inst_and_b63_2_0 (.A(wire63_1_0),.B(wire63_1_1),.Y(imd_Y63));
INVC inst_inv_b63_2_0 (.A(imd_Y63),.Y(Y63));
NANDC2x1 inst_clockedAND_b63_63 (.A(CLK),.B(Y63),.Y(imd_YF63));
INVC inst_clockedinv_b63_63 (.A(imd_YF63),.Y(YF63));


NANDC2x1 inst_and_b64_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire64_0_0));
INVC inst_inv_b64_0_0 (.A(imd_wire64_0_0),.Y(wire64_0_0));
NANDC2x1 inst_and_b64_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire64_0_1));
INVC inst_inv_b64_0_1 (.A(imd_wire64_0_1),.Y(wire64_0_1));
NANDC2x1 inst_and_b64_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire64_0_2));
INVC inst_inv_b64_0_2 (.A(imd_wire64_0_2),.Y(wire64_0_2));
NANDC2x1 inst_and_b64_1_0 (.A(wire64_0_0),.B(wire64_0_1),.Y(imd_wire64_1_0));
INVC inst_inv_b64_1_0 (.A(imd_wire64_1_0),.Y(wire64_1_0));
NANDC2x1 inst_and_b64_1_1 (.A(A6),.B(wire64_0_2),.Y(imd_wire64_1_1));
INVC inst_inv_b64_1_1 (.A(imd_wire64_1_1),.Y(wire64_1_1));
NANDC2x1 inst_and_b64_2_0 (.A(wire64_1_0),.B(wire64_1_1),.Y(imd_Y64));
INVC inst_inv_b64_2_0 (.A(imd_Y64),.Y(Y64));
NANDC2x1 inst_clockedAND_b64_64 (.A(CLK),.B(Y64),.Y(imd_YF64));
INVC inst_clockedinv_b64_64 (.A(imd_YF64),.Y(YF64));


NANDC2x1 inst_and_b65_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire65_0_0));
INVC inst_inv_b65_0_0 (.A(imd_wire65_0_0),.Y(wire65_0_0));
NANDC2x1 inst_and_b65_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire65_0_1));
INVC inst_inv_b65_0_1 (.A(imd_wire65_0_1),.Y(wire65_0_1));
NANDC2x1 inst_and_b65_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire65_0_2));
INVC inst_inv_b65_0_2 (.A(imd_wire65_0_2),.Y(wire65_0_2));
NANDC2x1 inst_and_b65_1_0 (.A(wire65_0_0),.B(wire65_0_1),.Y(imd_wire65_1_0));
INVC inst_inv_b65_1_0 (.A(imd_wire65_1_0),.Y(wire65_1_0));
NANDC2x1 inst_and_b65_1_1 (.A(A6),.B(wire65_0_2),.Y(imd_wire65_1_1));
INVC inst_inv_b65_1_1 (.A(imd_wire65_1_1),.Y(wire65_1_1));
NANDC2x1 inst_and_b65_2_0 (.A(wire65_1_0),.B(wire65_1_1),.Y(imd_Y65));
INVC inst_inv_b65_2_0 (.A(imd_Y65),.Y(Y65));
NANDC2x1 inst_clockedAND_b65_65 (.A(CLK),.B(Y65),.Y(imd_YF65));
INVC inst_clockedinv_b65_65 (.A(imd_YF65),.Y(YF65));


NANDC2x1 inst_and_b66_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire66_0_0));
INVC inst_inv_b66_0_0 (.A(imd_wire66_0_0),.Y(wire66_0_0));
NANDC2x1 inst_and_b66_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire66_0_1));
INVC inst_inv_b66_0_1 (.A(imd_wire66_0_1),.Y(wire66_0_1));
NANDC2x1 inst_and_b66_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire66_0_2));
INVC inst_inv_b66_0_2 (.A(imd_wire66_0_2),.Y(wire66_0_2));
NANDC2x1 inst_and_b66_1_0 (.A(wire66_0_0),.B(wire66_0_1),.Y(imd_wire66_1_0));
INVC inst_inv_b66_1_0 (.A(imd_wire66_1_0),.Y(wire66_1_0));
NANDC2x1 inst_and_b66_1_1 (.A(A6),.B(wire66_0_2),.Y(imd_wire66_1_1));
INVC inst_inv_b66_1_1 (.A(imd_wire66_1_1),.Y(wire66_1_1));
NANDC2x1 inst_and_b66_2_0 (.A(wire66_1_0),.B(wire66_1_1),.Y(imd_Y66));
INVC inst_inv_b66_2_0 (.A(imd_Y66),.Y(Y66));
NANDC2x1 inst_clockedAND_b66_66 (.A(CLK),.B(Y66),.Y(imd_YF66));
INVC inst_clockedinv_b66_66 (.A(imd_YF66),.Y(YF66));


NANDC2x1 inst_and_b67_0_0 (.A(A0),.B(A1),.Y(imd_wire67_0_0));
INVC inst_inv_b67_0_0 (.A(imd_wire67_0_0),.Y(wire67_0_0));
NANDC2x1 inst_and_b67_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire67_0_1));
INVC inst_inv_b67_0_1 (.A(imd_wire67_0_1),.Y(wire67_0_1));
NANDC2x1 inst_and_b67_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire67_0_2));
INVC inst_inv_b67_0_2 (.A(imd_wire67_0_2),.Y(wire67_0_2));
NANDC2x1 inst_and_b67_1_0 (.A(wire67_0_0),.B(wire67_0_1),.Y(imd_wire67_1_0));
INVC inst_inv_b67_1_0 (.A(imd_wire67_1_0),.Y(wire67_1_0));
NANDC2x1 inst_and_b67_1_1 (.A(A6),.B(wire67_0_2),.Y(imd_wire67_1_1));
INVC inst_inv_b67_1_1 (.A(imd_wire67_1_1),.Y(wire67_1_1));
NANDC2x1 inst_and_b67_2_0 (.A(wire67_1_0),.B(wire67_1_1),.Y(imd_Y67));
INVC inst_inv_b67_2_0 (.A(imd_Y67),.Y(Y67));
NANDC2x1 inst_clockedAND_b67_67 (.A(CLK),.B(Y67),.Y(imd_YF67));
INVC inst_clockedinv_b67_67 (.A(imd_YF67),.Y(YF67));


NANDC2x1 inst_and_b68_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire68_0_0));
INVC inst_inv_b68_0_0 (.A(imd_wire68_0_0),.Y(wire68_0_0));
NANDC2x1 inst_and_b68_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire68_0_1));
INVC inst_inv_b68_0_1 (.A(imd_wire68_0_1),.Y(wire68_0_1));
NANDC2x1 inst_and_b68_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire68_0_2));
INVC inst_inv_b68_0_2 (.A(imd_wire68_0_2),.Y(wire68_0_2));
NANDC2x1 inst_and_b68_1_0 (.A(wire68_0_0),.B(wire68_0_1),.Y(imd_wire68_1_0));
INVC inst_inv_b68_1_0 (.A(imd_wire68_1_0),.Y(wire68_1_0));
NANDC2x1 inst_and_b68_1_1 (.A(A6),.B(wire68_0_2),.Y(imd_wire68_1_1));
INVC inst_inv_b68_1_1 (.A(imd_wire68_1_1),.Y(wire68_1_1));
NANDC2x1 inst_and_b68_2_0 (.A(wire68_1_0),.B(wire68_1_1),.Y(imd_Y68));
INVC inst_inv_b68_2_0 (.A(imd_Y68),.Y(Y68));
NANDC2x1 inst_clockedAND_b68_68 (.A(CLK),.B(Y68),.Y(imd_YF68));
INVC inst_clockedinv_b68_68 (.A(imd_YF68),.Y(YF68));


NANDC2x1 inst_and_b69_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire69_0_0));
INVC inst_inv_b69_0_0 (.A(imd_wire69_0_0),.Y(wire69_0_0));
NANDC2x1 inst_and_b69_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire69_0_1));
INVC inst_inv_b69_0_1 (.A(imd_wire69_0_1),.Y(wire69_0_1));
NANDC2x1 inst_and_b69_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire69_0_2));
INVC inst_inv_b69_0_2 (.A(imd_wire69_0_2),.Y(wire69_0_2));
NANDC2x1 inst_and_b69_1_0 (.A(wire69_0_0),.B(wire69_0_1),.Y(imd_wire69_1_0));
INVC inst_inv_b69_1_0 (.A(imd_wire69_1_0),.Y(wire69_1_0));
NANDC2x1 inst_and_b69_1_1 (.A(A6),.B(wire69_0_2),.Y(imd_wire69_1_1));
INVC inst_inv_b69_1_1 (.A(imd_wire69_1_1),.Y(wire69_1_1));
NANDC2x1 inst_and_b69_2_0 (.A(wire69_1_0),.B(wire69_1_1),.Y(imd_Y69));
INVC inst_inv_b69_2_0 (.A(imd_Y69),.Y(Y69));
NANDC2x1 inst_clockedAND_b69_69 (.A(CLK),.B(Y69),.Y(imd_YF69));
INVC inst_clockedinv_b69_69 (.A(imd_YF69),.Y(YF69));


NANDC2x1 inst_and_b70_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire70_0_0));
INVC inst_inv_b70_0_0 (.A(imd_wire70_0_0),.Y(wire70_0_0));
NANDC2x1 inst_and_b70_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire70_0_1));
INVC inst_inv_b70_0_1 (.A(imd_wire70_0_1),.Y(wire70_0_1));
NANDC2x1 inst_and_b70_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire70_0_2));
INVC inst_inv_b70_0_2 (.A(imd_wire70_0_2),.Y(wire70_0_2));
NANDC2x1 inst_and_b70_1_0 (.A(wire70_0_0),.B(wire70_0_1),.Y(imd_wire70_1_0));
INVC inst_inv_b70_1_0 (.A(imd_wire70_1_0),.Y(wire70_1_0));
NANDC2x1 inst_and_b70_1_1 (.A(A6),.B(wire70_0_2),.Y(imd_wire70_1_1));
INVC inst_inv_b70_1_1 (.A(imd_wire70_1_1),.Y(wire70_1_1));
NANDC2x1 inst_and_b70_2_0 (.A(wire70_1_0),.B(wire70_1_1),.Y(imd_Y70));
INVC inst_inv_b70_2_0 (.A(imd_Y70),.Y(Y70));
NANDC2x1 inst_clockedAND_b70_70 (.A(CLK),.B(Y70),.Y(imd_YF70));
INVC inst_clockedinv_b70_70 (.A(imd_YF70),.Y(YF70));


NANDC2x1 inst_and_b71_0_0 (.A(A0),.B(A1),.Y(imd_wire71_0_0));
INVC inst_inv_b71_0_0 (.A(imd_wire71_0_0),.Y(wire71_0_0));
NANDC2x1 inst_and_b71_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire71_0_1));
INVC inst_inv_b71_0_1 (.A(imd_wire71_0_1),.Y(wire71_0_1));
NANDC2x1 inst_and_b71_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire71_0_2));
INVC inst_inv_b71_0_2 (.A(imd_wire71_0_2),.Y(wire71_0_2));
NANDC2x1 inst_and_b71_1_0 (.A(wire71_0_0),.B(wire71_0_1),.Y(imd_wire71_1_0));
INVC inst_inv_b71_1_0 (.A(imd_wire71_1_0),.Y(wire71_1_0));
NANDC2x1 inst_and_b71_1_1 (.A(A6),.B(wire71_0_2),.Y(imd_wire71_1_1));
INVC inst_inv_b71_1_1 (.A(imd_wire71_1_1),.Y(wire71_1_1));
NANDC2x1 inst_and_b71_2_0 (.A(wire71_1_0),.B(wire71_1_1),.Y(imd_Y71));
INVC inst_inv_b71_2_0 (.A(imd_Y71),.Y(Y71));
NANDC2x1 inst_clockedAND_b71_71 (.A(CLK),.B(Y71),.Y(imd_YF71));
INVC inst_clockedinv_b71_71 (.A(imd_YF71),.Y(YF71));


NANDC2x1 inst_and_b72_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire72_0_0));
INVC inst_inv_b72_0_0 (.A(imd_wire72_0_0),.Y(wire72_0_0));
NANDC2x1 inst_and_b72_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire72_0_1));
INVC inst_inv_b72_0_1 (.A(imd_wire72_0_1),.Y(wire72_0_1));
NANDC2x1 inst_and_b72_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire72_0_2));
INVC inst_inv_b72_0_2 (.A(imd_wire72_0_2),.Y(wire72_0_2));
NANDC2x1 inst_and_b72_1_0 (.A(wire72_0_0),.B(wire72_0_1),.Y(imd_wire72_1_0));
INVC inst_inv_b72_1_0 (.A(imd_wire72_1_0),.Y(wire72_1_0));
NANDC2x1 inst_and_b72_1_1 (.A(A6),.B(wire72_0_2),.Y(imd_wire72_1_1));
INVC inst_inv_b72_1_1 (.A(imd_wire72_1_1),.Y(wire72_1_1));
NANDC2x1 inst_and_b72_2_0 (.A(wire72_1_0),.B(wire72_1_1),.Y(imd_Y72));
INVC inst_inv_b72_2_0 (.A(imd_Y72),.Y(Y72));
NANDC2x1 inst_clockedAND_b72_72 (.A(CLK),.B(Y72),.Y(imd_YF72));
INVC inst_clockedinv_b72_72 (.A(imd_YF72),.Y(YF72));


NANDC2x1 inst_and_b73_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire73_0_0));
INVC inst_inv_b73_0_0 (.A(imd_wire73_0_0),.Y(wire73_0_0));
NANDC2x1 inst_and_b73_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire73_0_1));
INVC inst_inv_b73_0_1 (.A(imd_wire73_0_1),.Y(wire73_0_1));
NANDC2x1 inst_and_b73_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire73_0_2));
INVC inst_inv_b73_0_2 (.A(imd_wire73_0_2),.Y(wire73_0_2));
NANDC2x1 inst_and_b73_1_0 (.A(wire73_0_0),.B(wire73_0_1),.Y(imd_wire73_1_0));
INVC inst_inv_b73_1_0 (.A(imd_wire73_1_0),.Y(wire73_1_0));
NANDC2x1 inst_and_b73_1_1 (.A(A6),.B(wire73_0_2),.Y(imd_wire73_1_1));
INVC inst_inv_b73_1_1 (.A(imd_wire73_1_1),.Y(wire73_1_1));
NANDC2x1 inst_and_b73_2_0 (.A(wire73_1_0),.B(wire73_1_1),.Y(imd_Y73));
INVC inst_inv_b73_2_0 (.A(imd_Y73),.Y(Y73));
NANDC2x1 inst_clockedAND_b73_73 (.A(CLK),.B(Y73),.Y(imd_YF73));
INVC inst_clockedinv_b73_73 (.A(imd_YF73),.Y(YF73));


NANDC2x1 inst_and_b74_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire74_0_0));
INVC inst_inv_b74_0_0 (.A(imd_wire74_0_0),.Y(wire74_0_0));
NANDC2x1 inst_and_b74_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire74_0_1));
INVC inst_inv_b74_0_1 (.A(imd_wire74_0_1),.Y(wire74_0_1));
NANDC2x1 inst_and_b74_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire74_0_2));
INVC inst_inv_b74_0_2 (.A(imd_wire74_0_2),.Y(wire74_0_2));
NANDC2x1 inst_and_b74_1_0 (.A(wire74_0_0),.B(wire74_0_1),.Y(imd_wire74_1_0));
INVC inst_inv_b74_1_0 (.A(imd_wire74_1_0),.Y(wire74_1_0));
NANDC2x1 inst_and_b74_1_1 (.A(A6),.B(wire74_0_2),.Y(imd_wire74_1_1));
INVC inst_inv_b74_1_1 (.A(imd_wire74_1_1),.Y(wire74_1_1));
NANDC2x1 inst_and_b74_2_0 (.A(wire74_1_0),.B(wire74_1_1),.Y(imd_Y74));
INVC inst_inv_b74_2_0 (.A(imd_Y74),.Y(Y74));
NANDC2x1 inst_clockedAND_b74_74 (.A(CLK),.B(Y74),.Y(imd_YF74));
INVC inst_clockedinv_b74_74 (.A(imd_YF74),.Y(YF74));


NANDC2x1 inst_and_b75_0_0 (.A(A0),.B(A1),.Y(imd_wire75_0_0));
INVC inst_inv_b75_0_0 (.A(imd_wire75_0_0),.Y(wire75_0_0));
NANDC2x1 inst_and_b75_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire75_0_1));
INVC inst_inv_b75_0_1 (.A(imd_wire75_0_1),.Y(wire75_0_1));
NANDC2x1 inst_and_b75_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire75_0_2));
INVC inst_inv_b75_0_2 (.A(imd_wire75_0_2),.Y(wire75_0_2));
NANDC2x1 inst_and_b75_1_0 (.A(wire75_0_0),.B(wire75_0_1),.Y(imd_wire75_1_0));
INVC inst_inv_b75_1_0 (.A(imd_wire75_1_0),.Y(wire75_1_0));
NANDC2x1 inst_and_b75_1_1 (.A(A6),.B(wire75_0_2),.Y(imd_wire75_1_1));
INVC inst_inv_b75_1_1 (.A(imd_wire75_1_1),.Y(wire75_1_1));
NANDC2x1 inst_and_b75_2_0 (.A(wire75_1_0),.B(wire75_1_1),.Y(imd_Y75));
INVC inst_inv_b75_2_0 (.A(imd_Y75),.Y(Y75));
NANDC2x1 inst_clockedAND_b75_75 (.A(CLK),.B(Y75),.Y(imd_YF75));
INVC inst_clockedinv_b75_75 (.A(imd_YF75),.Y(YF75));


NANDC2x1 inst_and_b76_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire76_0_0));
INVC inst_inv_b76_0_0 (.A(imd_wire76_0_0),.Y(wire76_0_0));
NANDC2x1 inst_and_b76_0_1 (.A(A2),.B(A3),.Y(imd_wire76_0_1));
INVC inst_inv_b76_0_1 (.A(imd_wire76_0_1),.Y(wire76_0_1));
NANDC2x1 inst_and_b76_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire76_0_2));
INVC inst_inv_b76_0_2 (.A(imd_wire76_0_2),.Y(wire76_0_2));
NANDC2x1 inst_and_b76_1_0 (.A(wire76_0_0),.B(wire76_0_1),.Y(imd_wire76_1_0));
INVC inst_inv_b76_1_0 (.A(imd_wire76_1_0),.Y(wire76_1_0));
NANDC2x1 inst_and_b76_1_1 (.A(A6),.B(wire76_0_2),.Y(imd_wire76_1_1));
INVC inst_inv_b76_1_1 (.A(imd_wire76_1_1),.Y(wire76_1_1));
NANDC2x1 inst_and_b76_2_0 (.A(wire76_1_0),.B(wire76_1_1),.Y(imd_Y76));
INVC inst_inv_b76_2_0 (.A(imd_Y76),.Y(Y76));
NANDC2x1 inst_clockedAND_b76_76 (.A(CLK),.B(Y76),.Y(imd_YF76));
INVC inst_clockedinv_b76_76 (.A(imd_YF76),.Y(YF76));


NANDC2x1 inst_and_b77_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire77_0_0));
INVC inst_inv_b77_0_0 (.A(imd_wire77_0_0),.Y(wire77_0_0));
NANDC2x1 inst_and_b77_0_1 (.A(A2),.B(A3),.Y(imd_wire77_0_1));
INVC inst_inv_b77_0_1 (.A(imd_wire77_0_1),.Y(wire77_0_1));
NANDC2x1 inst_and_b77_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire77_0_2));
INVC inst_inv_b77_0_2 (.A(imd_wire77_0_2),.Y(wire77_0_2));
NANDC2x1 inst_and_b77_1_0 (.A(wire77_0_0),.B(wire77_0_1),.Y(imd_wire77_1_0));
INVC inst_inv_b77_1_0 (.A(imd_wire77_1_0),.Y(wire77_1_0));
NANDC2x1 inst_and_b77_1_1 (.A(A6),.B(wire77_0_2),.Y(imd_wire77_1_1));
INVC inst_inv_b77_1_1 (.A(imd_wire77_1_1),.Y(wire77_1_1));
NANDC2x1 inst_and_b77_2_0 (.A(wire77_1_0),.B(wire77_1_1),.Y(imd_Y77));
INVC inst_inv_b77_2_0 (.A(imd_Y77),.Y(Y77));
NANDC2x1 inst_clockedAND_b77_77 (.A(CLK),.B(Y77),.Y(imd_YF77));
INVC inst_clockedinv_b77_77 (.A(imd_YF77),.Y(YF77));


NANDC2x1 inst_and_b78_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire78_0_0));
INVC inst_inv_b78_0_0 (.A(imd_wire78_0_0),.Y(wire78_0_0));
NANDC2x1 inst_and_b78_0_1 (.A(A2),.B(A3),.Y(imd_wire78_0_1));
INVC inst_inv_b78_0_1 (.A(imd_wire78_0_1),.Y(wire78_0_1));
NANDC2x1 inst_and_b78_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire78_0_2));
INVC inst_inv_b78_0_2 (.A(imd_wire78_0_2),.Y(wire78_0_2));
NANDC2x1 inst_and_b78_1_0 (.A(wire78_0_0),.B(wire78_0_1),.Y(imd_wire78_1_0));
INVC inst_inv_b78_1_0 (.A(imd_wire78_1_0),.Y(wire78_1_0));
NANDC2x1 inst_and_b78_1_1 (.A(A6),.B(wire78_0_2),.Y(imd_wire78_1_1));
INVC inst_inv_b78_1_1 (.A(imd_wire78_1_1),.Y(wire78_1_1));
NANDC2x1 inst_and_b78_2_0 (.A(wire78_1_0),.B(wire78_1_1),.Y(imd_Y78));
INVC inst_inv_b78_2_0 (.A(imd_Y78),.Y(Y78));
NANDC2x1 inst_clockedAND_b78_78 (.A(CLK),.B(Y78),.Y(imd_YF78));
INVC inst_clockedinv_b78_78 (.A(imd_YF78),.Y(YF78));


NANDC2x1 inst_and_b79_0_0 (.A(A0),.B(A1),.Y(imd_wire79_0_0));
INVC inst_inv_b79_0_0 (.A(imd_wire79_0_0),.Y(wire79_0_0));
NANDC2x1 inst_and_b79_0_1 (.A(A2),.B(A3),.Y(imd_wire79_0_1));
INVC inst_inv_b79_0_1 (.A(imd_wire79_0_1),.Y(wire79_0_1));
NANDC2x1 inst_and_b79_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire79_0_2));
INVC inst_inv_b79_0_2 (.A(imd_wire79_0_2),.Y(wire79_0_2));
NANDC2x1 inst_and_b79_1_0 (.A(wire79_0_0),.B(wire79_0_1),.Y(imd_wire79_1_0));
INVC inst_inv_b79_1_0 (.A(imd_wire79_1_0),.Y(wire79_1_0));
NANDC2x1 inst_and_b79_1_1 (.A(A6),.B(wire79_0_2),.Y(imd_wire79_1_1));
INVC inst_inv_b79_1_1 (.A(imd_wire79_1_1),.Y(wire79_1_1));
NANDC2x1 inst_and_b79_2_0 (.A(wire79_1_0),.B(wire79_1_1),.Y(imd_Y79));
INVC inst_inv_b79_2_0 (.A(imd_Y79),.Y(Y79));
NANDC2x1 inst_clockedAND_b79_79 (.A(CLK),.B(Y79),.Y(imd_YF79));
INVC inst_clockedinv_b79_79 (.A(imd_YF79),.Y(YF79));


NANDC2x1 inst_and_b80_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire80_0_0));
INVC inst_inv_b80_0_0 (.A(imd_wire80_0_0),.Y(wire80_0_0));
NANDC2x1 inst_and_b80_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire80_0_1));
INVC inst_inv_b80_0_1 (.A(imd_wire80_0_1),.Y(wire80_0_1));
NANDC2x1 inst_and_b80_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire80_0_2));
INVC inst_inv_b80_0_2 (.A(imd_wire80_0_2),.Y(wire80_0_2));
NANDC2x1 inst_and_b80_1_0 (.A(wire80_0_0),.B(wire80_0_1),.Y(imd_wire80_1_0));
INVC inst_inv_b80_1_0 (.A(imd_wire80_1_0),.Y(wire80_1_0));
NANDC2x1 inst_and_b80_1_1 (.A(A6),.B(wire80_0_2),.Y(imd_wire80_1_1));
INVC inst_inv_b80_1_1 (.A(imd_wire80_1_1),.Y(wire80_1_1));
NANDC2x1 inst_and_b80_2_0 (.A(wire80_1_0),.B(wire80_1_1),.Y(imd_Y80));
INVC inst_inv_b80_2_0 (.A(imd_Y80),.Y(Y80));
NANDC2x1 inst_clockedAND_b80_80 (.A(CLK),.B(Y80),.Y(imd_YF80));
INVC inst_clockedinv_b80_80 (.A(imd_YF80),.Y(YF80));


NANDC2x1 inst_and_b81_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire81_0_0));
INVC inst_inv_b81_0_0 (.A(imd_wire81_0_0),.Y(wire81_0_0));
NANDC2x1 inst_and_b81_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire81_0_1));
INVC inst_inv_b81_0_1 (.A(imd_wire81_0_1),.Y(wire81_0_1));
NANDC2x1 inst_and_b81_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire81_0_2));
INVC inst_inv_b81_0_2 (.A(imd_wire81_0_2),.Y(wire81_0_2));
NANDC2x1 inst_and_b81_1_0 (.A(wire81_0_0),.B(wire81_0_1),.Y(imd_wire81_1_0));
INVC inst_inv_b81_1_0 (.A(imd_wire81_1_0),.Y(wire81_1_0));
NANDC2x1 inst_and_b81_1_1 (.A(A6),.B(wire81_0_2),.Y(imd_wire81_1_1));
INVC inst_inv_b81_1_1 (.A(imd_wire81_1_1),.Y(wire81_1_1));
NANDC2x1 inst_and_b81_2_0 (.A(wire81_1_0),.B(wire81_1_1),.Y(imd_Y81));
INVC inst_inv_b81_2_0 (.A(imd_Y81),.Y(Y81));
NANDC2x1 inst_clockedAND_b81_81 (.A(CLK),.B(Y81),.Y(imd_YF81));
INVC inst_clockedinv_b81_81 (.A(imd_YF81),.Y(YF81));


NANDC2x1 inst_and_b82_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire82_0_0));
INVC inst_inv_b82_0_0 (.A(imd_wire82_0_0),.Y(wire82_0_0));
NANDC2x1 inst_and_b82_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire82_0_1));
INVC inst_inv_b82_0_1 (.A(imd_wire82_0_1),.Y(wire82_0_1));
NANDC2x1 inst_and_b82_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire82_0_2));
INVC inst_inv_b82_0_2 (.A(imd_wire82_0_2),.Y(wire82_0_2));
NANDC2x1 inst_and_b82_1_0 (.A(wire82_0_0),.B(wire82_0_1),.Y(imd_wire82_1_0));
INVC inst_inv_b82_1_0 (.A(imd_wire82_1_0),.Y(wire82_1_0));
NANDC2x1 inst_and_b82_1_1 (.A(A6),.B(wire82_0_2),.Y(imd_wire82_1_1));
INVC inst_inv_b82_1_1 (.A(imd_wire82_1_1),.Y(wire82_1_1));
NANDC2x1 inst_and_b82_2_0 (.A(wire82_1_0),.B(wire82_1_1),.Y(imd_Y82));
INVC inst_inv_b82_2_0 (.A(imd_Y82),.Y(Y82));
NANDC2x1 inst_clockedAND_b82_82 (.A(CLK),.B(Y82),.Y(imd_YF82));
INVC inst_clockedinv_b82_82 (.A(imd_YF82),.Y(YF82));


NANDC2x1 inst_and_b83_0_0 (.A(A0),.B(A1),.Y(imd_wire83_0_0));
INVC inst_inv_b83_0_0 (.A(imd_wire83_0_0),.Y(wire83_0_0));
NANDC2x1 inst_and_b83_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire83_0_1));
INVC inst_inv_b83_0_1 (.A(imd_wire83_0_1),.Y(wire83_0_1));
NANDC2x1 inst_and_b83_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire83_0_2));
INVC inst_inv_b83_0_2 (.A(imd_wire83_0_2),.Y(wire83_0_2));
NANDC2x1 inst_and_b83_1_0 (.A(wire83_0_0),.B(wire83_0_1),.Y(imd_wire83_1_0));
INVC inst_inv_b83_1_0 (.A(imd_wire83_1_0),.Y(wire83_1_0));
NANDC2x1 inst_and_b83_1_1 (.A(A6),.B(wire83_0_2),.Y(imd_wire83_1_1));
INVC inst_inv_b83_1_1 (.A(imd_wire83_1_1),.Y(wire83_1_1));
NANDC2x1 inst_and_b83_2_0 (.A(wire83_1_0),.B(wire83_1_1),.Y(imd_Y83));
INVC inst_inv_b83_2_0 (.A(imd_Y83),.Y(Y83));
NANDC2x1 inst_clockedAND_b83_83 (.A(CLK),.B(Y83),.Y(imd_YF83));
INVC inst_clockedinv_b83_83 (.A(imd_YF83),.Y(YF83));


NANDC2x1 inst_and_b84_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire84_0_0));
INVC inst_inv_b84_0_0 (.A(imd_wire84_0_0),.Y(wire84_0_0));
NANDC2x1 inst_and_b84_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire84_0_1));
INVC inst_inv_b84_0_1 (.A(imd_wire84_0_1),.Y(wire84_0_1));
NANDC2x1 inst_and_b84_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire84_0_2));
INVC inst_inv_b84_0_2 (.A(imd_wire84_0_2),.Y(wire84_0_2));
NANDC2x1 inst_and_b84_1_0 (.A(wire84_0_0),.B(wire84_0_1),.Y(imd_wire84_1_0));
INVC inst_inv_b84_1_0 (.A(imd_wire84_1_0),.Y(wire84_1_0));
NANDC2x1 inst_and_b84_1_1 (.A(A6),.B(wire84_0_2),.Y(imd_wire84_1_1));
INVC inst_inv_b84_1_1 (.A(imd_wire84_1_1),.Y(wire84_1_1));
NANDC2x1 inst_and_b84_2_0 (.A(wire84_1_0),.B(wire84_1_1),.Y(imd_Y84));
INVC inst_inv_b84_2_0 (.A(imd_Y84),.Y(Y84));
NANDC2x1 inst_clockedAND_b84_84 (.A(CLK),.B(Y84),.Y(imd_YF84));
INVC inst_clockedinv_b84_84 (.A(imd_YF84),.Y(YF84));


NANDC2x1 inst_and_b85_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire85_0_0));
INVC inst_inv_b85_0_0 (.A(imd_wire85_0_0),.Y(wire85_0_0));
NANDC2x1 inst_and_b85_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire85_0_1));
INVC inst_inv_b85_0_1 (.A(imd_wire85_0_1),.Y(wire85_0_1));
NANDC2x1 inst_and_b85_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire85_0_2));
INVC inst_inv_b85_0_2 (.A(imd_wire85_0_2),.Y(wire85_0_2));
NANDC2x1 inst_and_b85_1_0 (.A(wire85_0_0),.B(wire85_0_1),.Y(imd_wire85_1_0));
INVC inst_inv_b85_1_0 (.A(imd_wire85_1_0),.Y(wire85_1_0));
NANDC2x1 inst_and_b85_1_1 (.A(A6),.B(wire85_0_2),.Y(imd_wire85_1_1));
INVC inst_inv_b85_1_1 (.A(imd_wire85_1_1),.Y(wire85_1_1));
NANDC2x1 inst_and_b85_2_0 (.A(wire85_1_0),.B(wire85_1_1),.Y(imd_Y85));
INVC inst_inv_b85_2_0 (.A(imd_Y85),.Y(Y85));
NANDC2x1 inst_clockedAND_b85_85 (.A(CLK),.B(Y85),.Y(imd_YF85));
INVC inst_clockedinv_b85_85 (.A(imd_YF85),.Y(YF85));


NANDC2x1 inst_and_b86_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire86_0_0));
INVC inst_inv_b86_0_0 (.A(imd_wire86_0_0),.Y(wire86_0_0));
NANDC2x1 inst_and_b86_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire86_0_1));
INVC inst_inv_b86_0_1 (.A(imd_wire86_0_1),.Y(wire86_0_1));
NANDC2x1 inst_and_b86_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire86_0_2));
INVC inst_inv_b86_0_2 (.A(imd_wire86_0_2),.Y(wire86_0_2));
NANDC2x1 inst_and_b86_1_0 (.A(wire86_0_0),.B(wire86_0_1),.Y(imd_wire86_1_0));
INVC inst_inv_b86_1_0 (.A(imd_wire86_1_0),.Y(wire86_1_0));
NANDC2x1 inst_and_b86_1_1 (.A(A6),.B(wire86_0_2),.Y(imd_wire86_1_1));
INVC inst_inv_b86_1_1 (.A(imd_wire86_1_1),.Y(wire86_1_1));
NANDC2x1 inst_and_b86_2_0 (.A(wire86_1_0),.B(wire86_1_1),.Y(imd_Y86));
INVC inst_inv_b86_2_0 (.A(imd_Y86),.Y(Y86));
NANDC2x1 inst_clockedAND_b86_86 (.A(CLK),.B(Y86),.Y(imd_YF86));
INVC inst_clockedinv_b86_86 (.A(imd_YF86),.Y(YF86));


NANDC2x1 inst_and_b87_0_0 (.A(A0),.B(A1),.Y(imd_wire87_0_0));
INVC inst_inv_b87_0_0 (.A(imd_wire87_0_0),.Y(wire87_0_0));
NANDC2x1 inst_and_b87_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire87_0_1));
INVC inst_inv_b87_0_1 (.A(imd_wire87_0_1),.Y(wire87_0_1));
NANDC2x1 inst_and_b87_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire87_0_2));
INVC inst_inv_b87_0_2 (.A(imd_wire87_0_2),.Y(wire87_0_2));
NANDC2x1 inst_and_b87_1_0 (.A(wire87_0_0),.B(wire87_0_1),.Y(imd_wire87_1_0));
INVC inst_inv_b87_1_0 (.A(imd_wire87_1_0),.Y(wire87_1_0));
NANDC2x1 inst_and_b87_1_1 (.A(A6),.B(wire87_0_2),.Y(imd_wire87_1_1));
INVC inst_inv_b87_1_1 (.A(imd_wire87_1_1),.Y(wire87_1_1));
NANDC2x1 inst_and_b87_2_0 (.A(wire87_1_0),.B(wire87_1_1),.Y(imd_Y87));
INVC inst_inv_b87_2_0 (.A(imd_Y87),.Y(Y87));
NANDC2x1 inst_clockedAND_b87_87 (.A(CLK),.B(Y87),.Y(imd_YF87));
INVC inst_clockedinv_b87_87 (.A(imd_YF87),.Y(YF87));


NANDC2x1 inst_and_b88_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire88_0_0));
INVC inst_inv_b88_0_0 (.A(imd_wire88_0_0),.Y(wire88_0_0));
NANDC2x1 inst_and_b88_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire88_0_1));
INVC inst_inv_b88_0_1 (.A(imd_wire88_0_1),.Y(wire88_0_1));
NANDC2x1 inst_and_b88_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire88_0_2));
INVC inst_inv_b88_0_2 (.A(imd_wire88_0_2),.Y(wire88_0_2));
NANDC2x1 inst_and_b88_1_0 (.A(wire88_0_0),.B(wire88_0_1),.Y(imd_wire88_1_0));
INVC inst_inv_b88_1_0 (.A(imd_wire88_1_0),.Y(wire88_1_0));
NANDC2x1 inst_and_b88_1_1 (.A(A6),.B(wire88_0_2),.Y(imd_wire88_1_1));
INVC inst_inv_b88_1_1 (.A(imd_wire88_1_1),.Y(wire88_1_1));
NANDC2x1 inst_and_b88_2_0 (.A(wire88_1_0),.B(wire88_1_1),.Y(imd_Y88));
INVC inst_inv_b88_2_0 (.A(imd_Y88),.Y(Y88));
NANDC2x1 inst_clockedAND_b88_88 (.A(CLK),.B(Y88),.Y(imd_YF88));
INVC inst_clockedinv_b88_88 (.A(imd_YF88),.Y(YF88));


NANDC2x1 inst_and_b89_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire89_0_0));
INVC inst_inv_b89_0_0 (.A(imd_wire89_0_0),.Y(wire89_0_0));
NANDC2x1 inst_and_b89_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire89_0_1));
INVC inst_inv_b89_0_1 (.A(imd_wire89_0_1),.Y(wire89_0_1));
NANDC2x1 inst_and_b89_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire89_0_2));
INVC inst_inv_b89_0_2 (.A(imd_wire89_0_2),.Y(wire89_0_2));
NANDC2x1 inst_and_b89_1_0 (.A(wire89_0_0),.B(wire89_0_1),.Y(imd_wire89_1_0));
INVC inst_inv_b89_1_0 (.A(imd_wire89_1_0),.Y(wire89_1_0));
NANDC2x1 inst_and_b89_1_1 (.A(A6),.B(wire89_0_2),.Y(imd_wire89_1_1));
INVC inst_inv_b89_1_1 (.A(imd_wire89_1_1),.Y(wire89_1_1));
NANDC2x1 inst_and_b89_2_0 (.A(wire89_1_0),.B(wire89_1_1),.Y(imd_Y89));
INVC inst_inv_b89_2_0 (.A(imd_Y89),.Y(Y89));
NANDC2x1 inst_clockedAND_b89_89 (.A(CLK),.B(Y89),.Y(imd_YF89));
INVC inst_clockedinv_b89_89 (.A(imd_YF89),.Y(YF89));


NANDC2x1 inst_and_b90_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire90_0_0));
INVC inst_inv_b90_0_0 (.A(imd_wire90_0_0),.Y(wire90_0_0));
NANDC2x1 inst_and_b90_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire90_0_1));
INVC inst_inv_b90_0_1 (.A(imd_wire90_0_1),.Y(wire90_0_1));
NANDC2x1 inst_and_b90_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire90_0_2));
INVC inst_inv_b90_0_2 (.A(imd_wire90_0_2),.Y(wire90_0_2));
NANDC2x1 inst_and_b90_1_0 (.A(wire90_0_0),.B(wire90_0_1),.Y(imd_wire90_1_0));
INVC inst_inv_b90_1_0 (.A(imd_wire90_1_0),.Y(wire90_1_0));
NANDC2x1 inst_and_b90_1_1 (.A(A6),.B(wire90_0_2),.Y(imd_wire90_1_1));
INVC inst_inv_b90_1_1 (.A(imd_wire90_1_1),.Y(wire90_1_1));
NANDC2x1 inst_and_b90_2_0 (.A(wire90_1_0),.B(wire90_1_1),.Y(imd_Y90));
INVC inst_inv_b90_2_0 (.A(imd_Y90),.Y(Y90));
NANDC2x1 inst_clockedAND_b90_90 (.A(CLK),.B(Y90),.Y(imd_YF90));
INVC inst_clockedinv_b90_90 (.A(imd_YF90),.Y(YF90));


NANDC2x1 inst_and_b91_0_0 (.A(A0),.B(A1),.Y(imd_wire91_0_0));
INVC inst_inv_b91_0_0 (.A(imd_wire91_0_0),.Y(wire91_0_0));
NANDC2x1 inst_and_b91_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire91_0_1));
INVC inst_inv_b91_0_1 (.A(imd_wire91_0_1),.Y(wire91_0_1));
NANDC2x1 inst_and_b91_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire91_0_2));
INVC inst_inv_b91_0_2 (.A(imd_wire91_0_2),.Y(wire91_0_2));
NANDC2x1 inst_and_b91_1_0 (.A(wire91_0_0),.B(wire91_0_1),.Y(imd_wire91_1_0));
INVC inst_inv_b91_1_0 (.A(imd_wire91_1_0),.Y(wire91_1_0));
NANDC2x1 inst_and_b91_1_1 (.A(A6),.B(wire91_0_2),.Y(imd_wire91_1_1));
INVC inst_inv_b91_1_1 (.A(imd_wire91_1_1),.Y(wire91_1_1));
NANDC2x1 inst_and_b91_2_0 (.A(wire91_1_0),.B(wire91_1_1),.Y(imd_Y91));
INVC inst_inv_b91_2_0 (.A(imd_Y91),.Y(Y91));
NANDC2x1 inst_clockedAND_b91_91 (.A(CLK),.B(Y91),.Y(imd_YF91));
INVC inst_clockedinv_b91_91 (.A(imd_YF91),.Y(YF91));


NANDC2x1 inst_and_b92_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire92_0_0));
INVC inst_inv_b92_0_0 (.A(imd_wire92_0_0),.Y(wire92_0_0));
NANDC2x1 inst_and_b92_0_1 (.A(A2),.B(A3),.Y(imd_wire92_0_1));
INVC inst_inv_b92_0_1 (.A(imd_wire92_0_1),.Y(wire92_0_1));
NANDC2x1 inst_and_b92_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire92_0_2));
INVC inst_inv_b92_0_2 (.A(imd_wire92_0_2),.Y(wire92_0_2));
NANDC2x1 inst_and_b92_1_0 (.A(wire92_0_0),.B(wire92_0_1),.Y(imd_wire92_1_0));
INVC inst_inv_b92_1_0 (.A(imd_wire92_1_0),.Y(wire92_1_0));
NANDC2x1 inst_and_b92_1_1 (.A(A6),.B(wire92_0_2),.Y(imd_wire92_1_1));
INVC inst_inv_b92_1_1 (.A(imd_wire92_1_1),.Y(wire92_1_1));
NANDC2x1 inst_and_b92_2_0 (.A(wire92_1_0),.B(wire92_1_1),.Y(imd_Y92));
INVC inst_inv_b92_2_0 (.A(imd_Y92),.Y(Y92));
NANDC2x1 inst_clockedAND_b92_92 (.A(CLK),.B(Y92),.Y(imd_YF92));
INVC inst_clockedinv_b92_92 (.A(imd_YF92),.Y(YF92));


NANDC2x1 inst_and_b93_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire93_0_0));
INVC inst_inv_b93_0_0 (.A(imd_wire93_0_0),.Y(wire93_0_0));
NANDC2x1 inst_and_b93_0_1 (.A(A2),.B(A3),.Y(imd_wire93_0_1));
INVC inst_inv_b93_0_1 (.A(imd_wire93_0_1),.Y(wire93_0_1));
NANDC2x1 inst_and_b93_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire93_0_2));
INVC inst_inv_b93_0_2 (.A(imd_wire93_0_2),.Y(wire93_0_2));
NANDC2x1 inst_and_b93_1_0 (.A(wire93_0_0),.B(wire93_0_1),.Y(imd_wire93_1_0));
INVC inst_inv_b93_1_0 (.A(imd_wire93_1_0),.Y(wire93_1_0));
NANDC2x1 inst_and_b93_1_1 (.A(A6),.B(wire93_0_2),.Y(imd_wire93_1_1));
INVC inst_inv_b93_1_1 (.A(imd_wire93_1_1),.Y(wire93_1_1));
NANDC2x1 inst_and_b93_2_0 (.A(wire93_1_0),.B(wire93_1_1),.Y(imd_Y93));
INVC inst_inv_b93_2_0 (.A(imd_Y93),.Y(Y93));
NANDC2x1 inst_clockedAND_b93_93 (.A(CLK),.B(Y93),.Y(imd_YF93));
INVC inst_clockedinv_b93_93 (.A(imd_YF93),.Y(YF93));


NANDC2x1 inst_and_b94_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire94_0_0));
INVC inst_inv_b94_0_0 (.A(imd_wire94_0_0),.Y(wire94_0_0));
NANDC2x1 inst_and_b94_0_1 (.A(A2),.B(A3),.Y(imd_wire94_0_1));
INVC inst_inv_b94_0_1 (.A(imd_wire94_0_1),.Y(wire94_0_1));
NANDC2x1 inst_and_b94_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire94_0_2));
INVC inst_inv_b94_0_2 (.A(imd_wire94_0_2),.Y(wire94_0_2));
NANDC2x1 inst_and_b94_1_0 (.A(wire94_0_0),.B(wire94_0_1),.Y(imd_wire94_1_0));
INVC inst_inv_b94_1_0 (.A(imd_wire94_1_0),.Y(wire94_1_0));
NANDC2x1 inst_and_b94_1_1 (.A(A6),.B(wire94_0_2),.Y(imd_wire94_1_1));
INVC inst_inv_b94_1_1 (.A(imd_wire94_1_1),.Y(wire94_1_1));
NANDC2x1 inst_and_b94_2_0 (.A(wire94_1_0),.B(wire94_1_1),.Y(imd_Y94));
INVC inst_inv_b94_2_0 (.A(imd_Y94),.Y(Y94));
NANDC2x1 inst_clockedAND_b94_94 (.A(CLK),.B(Y94),.Y(imd_YF94));
INVC inst_clockedinv_b94_94 (.A(imd_YF94),.Y(YF94));


NANDC2x1 inst_and_b95_0_0 (.A(A0),.B(A1),.Y(imd_wire95_0_0));
INVC inst_inv_b95_0_0 (.A(imd_wire95_0_0),.Y(wire95_0_0));
NANDC2x1 inst_and_b95_0_1 (.A(A2),.B(A3),.Y(imd_wire95_0_1));
INVC inst_inv_b95_0_1 (.A(imd_wire95_0_1),.Y(wire95_0_1));
NANDC2x1 inst_and_b95_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire95_0_2));
INVC inst_inv_b95_0_2 (.A(imd_wire95_0_2),.Y(wire95_0_2));
NANDC2x1 inst_and_b95_1_0 (.A(wire95_0_0),.B(wire95_0_1),.Y(imd_wire95_1_0));
INVC inst_inv_b95_1_0 (.A(imd_wire95_1_0),.Y(wire95_1_0));
NANDC2x1 inst_and_b95_1_1 (.A(A6),.B(wire95_0_2),.Y(imd_wire95_1_1));
INVC inst_inv_b95_1_1 (.A(imd_wire95_1_1),.Y(wire95_1_1));
NANDC2x1 inst_and_b95_2_0 (.A(wire95_1_0),.B(wire95_1_1),.Y(imd_Y95));
INVC inst_inv_b95_2_0 (.A(imd_Y95),.Y(Y95));
NANDC2x1 inst_clockedAND_b95_95 (.A(CLK),.B(Y95),.Y(imd_YF95));
INVC inst_clockedinv_b95_95 (.A(imd_YF95),.Y(YF95));


NANDC2x1 inst_and_b96_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire96_0_0));
INVC inst_inv_b96_0_0 (.A(imd_wire96_0_0),.Y(wire96_0_0));
NANDC2x1 inst_and_b96_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire96_0_1));
INVC inst_inv_b96_0_1 (.A(imd_wire96_0_1),.Y(wire96_0_1));
NANDC2x1 inst_and_b96_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire96_0_2));
INVC inst_inv_b96_0_2 (.A(imd_wire96_0_2),.Y(wire96_0_2));
NANDC2x1 inst_and_b96_1_0 (.A(wire96_0_0),.B(wire96_0_1),.Y(imd_wire96_1_0));
INVC inst_inv_b96_1_0 (.A(imd_wire96_1_0),.Y(wire96_1_0));
NANDC2x1 inst_and_b96_1_1 (.A(A6),.B(wire96_0_2),.Y(imd_wire96_1_1));
INVC inst_inv_b96_1_1 (.A(imd_wire96_1_1),.Y(wire96_1_1));
NANDC2x1 inst_and_b96_2_0 (.A(wire96_1_0),.B(wire96_1_1),.Y(imd_Y96));
INVC inst_inv_b96_2_0 (.A(imd_Y96),.Y(Y96));
NANDC2x1 inst_clockedAND_b96_96 (.A(CLK),.B(Y96),.Y(imd_YF96));
INVC inst_clockedinv_b96_96 (.A(imd_YF96),.Y(YF96));


NANDC2x1 inst_and_b97_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire97_0_0));
INVC inst_inv_b97_0_0 (.A(imd_wire97_0_0),.Y(wire97_0_0));
NANDC2x1 inst_and_b97_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire97_0_1));
INVC inst_inv_b97_0_1 (.A(imd_wire97_0_1),.Y(wire97_0_1));
NANDC2x1 inst_and_b97_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire97_0_2));
INVC inst_inv_b97_0_2 (.A(imd_wire97_0_2),.Y(wire97_0_2));
NANDC2x1 inst_and_b97_1_0 (.A(wire97_0_0),.B(wire97_0_1),.Y(imd_wire97_1_0));
INVC inst_inv_b97_1_0 (.A(imd_wire97_1_0),.Y(wire97_1_0));
NANDC2x1 inst_and_b97_1_1 (.A(A6),.B(wire97_0_2),.Y(imd_wire97_1_1));
INVC inst_inv_b97_1_1 (.A(imd_wire97_1_1),.Y(wire97_1_1));
NANDC2x1 inst_and_b97_2_0 (.A(wire97_1_0),.B(wire97_1_1),.Y(imd_Y97));
INVC inst_inv_b97_2_0 (.A(imd_Y97),.Y(Y97));
NANDC2x1 inst_clockedAND_b97_97 (.A(CLK),.B(Y97),.Y(imd_YF97));
INVC inst_clockedinv_b97_97 (.A(imd_YF97),.Y(YF97));


NANDC2x1 inst_and_b98_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire98_0_0));
INVC inst_inv_b98_0_0 (.A(imd_wire98_0_0),.Y(wire98_0_0));
NANDC2x1 inst_and_b98_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire98_0_1));
INVC inst_inv_b98_0_1 (.A(imd_wire98_0_1),.Y(wire98_0_1));
NANDC2x1 inst_and_b98_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire98_0_2));
INVC inst_inv_b98_0_2 (.A(imd_wire98_0_2),.Y(wire98_0_2));
NANDC2x1 inst_and_b98_1_0 (.A(wire98_0_0),.B(wire98_0_1),.Y(imd_wire98_1_0));
INVC inst_inv_b98_1_0 (.A(imd_wire98_1_0),.Y(wire98_1_0));
NANDC2x1 inst_and_b98_1_1 (.A(A6),.B(wire98_0_2),.Y(imd_wire98_1_1));
INVC inst_inv_b98_1_1 (.A(imd_wire98_1_1),.Y(wire98_1_1));
NANDC2x1 inst_and_b98_2_0 (.A(wire98_1_0),.B(wire98_1_1),.Y(imd_Y98));
INVC inst_inv_b98_2_0 (.A(imd_Y98),.Y(Y98));
NANDC2x1 inst_clockedAND_b98_98 (.A(CLK),.B(Y98),.Y(imd_YF98));
INVC inst_clockedinv_b98_98 (.A(imd_YF98),.Y(YF98));


NANDC2x1 inst_and_b99_0_0 (.A(A0),.B(A1),.Y(imd_wire99_0_0));
INVC inst_inv_b99_0_0 (.A(imd_wire99_0_0),.Y(wire99_0_0));
NANDC2x1 inst_and_b99_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire99_0_1));
INVC inst_inv_b99_0_1 (.A(imd_wire99_0_1),.Y(wire99_0_1));
NANDC2x1 inst_and_b99_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire99_0_2));
INVC inst_inv_b99_0_2 (.A(imd_wire99_0_2),.Y(wire99_0_2));
NANDC2x1 inst_and_b99_1_0 (.A(wire99_0_0),.B(wire99_0_1),.Y(imd_wire99_1_0));
INVC inst_inv_b99_1_0 (.A(imd_wire99_1_0),.Y(wire99_1_0));
NANDC2x1 inst_and_b99_1_1 (.A(A6),.B(wire99_0_2),.Y(imd_wire99_1_1));
INVC inst_inv_b99_1_1 (.A(imd_wire99_1_1),.Y(wire99_1_1));
NANDC2x1 inst_and_b99_2_0 (.A(wire99_1_0),.B(wire99_1_1),.Y(imd_Y99));
INVC inst_inv_b99_2_0 (.A(imd_Y99),.Y(Y99));
NANDC2x1 inst_clockedAND_b99_99 (.A(CLK),.B(Y99),.Y(imd_YF99));
INVC inst_clockedinv_b99_99 (.A(imd_YF99),.Y(YF99));


NANDC2x1 inst_and_b100_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire100_0_0));
INVC inst_inv_b100_0_0 (.A(imd_wire100_0_0),.Y(wire100_0_0));
NANDC2x1 inst_and_b100_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire100_0_1));
INVC inst_inv_b100_0_1 (.A(imd_wire100_0_1),.Y(wire100_0_1));
NANDC2x1 inst_and_b100_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire100_0_2));
INVC inst_inv_b100_0_2 (.A(imd_wire100_0_2),.Y(wire100_0_2));
NANDC2x1 inst_and_b100_1_0 (.A(wire100_0_0),.B(wire100_0_1),.Y(imd_wire100_1_0));
INVC inst_inv_b100_1_0 (.A(imd_wire100_1_0),.Y(wire100_1_0));
NANDC2x1 inst_and_b100_1_1 (.A(A6),.B(wire100_0_2),.Y(imd_wire100_1_1));
INVC inst_inv_b100_1_1 (.A(imd_wire100_1_1),.Y(wire100_1_1));
NANDC2x1 inst_and_b100_2_0 (.A(wire100_1_0),.B(wire100_1_1),.Y(imd_Y100));
INVC inst_inv_b100_2_0 (.A(imd_Y100),.Y(Y100));
NANDC2x1 inst_clockedAND_b100_100 (.A(CLK),.B(Y100),.Y(imd_YF100));
INVC inst_clockedinv_b100_100 (.A(imd_YF100),.Y(YF100));


NANDC2x1 inst_and_b101_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire101_0_0));
INVC inst_inv_b101_0_0 (.A(imd_wire101_0_0),.Y(wire101_0_0));
NANDC2x1 inst_and_b101_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire101_0_1));
INVC inst_inv_b101_0_1 (.A(imd_wire101_0_1),.Y(wire101_0_1));
NANDC2x1 inst_and_b101_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire101_0_2));
INVC inst_inv_b101_0_2 (.A(imd_wire101_0_2),.Y(wire101_0_2));
NANDC2x1 inst_and_b101_1_0 (.A(wire101_0_0),.B(wire101_0_1),.Y(imd_wire101_1_0));
INVC inst_inv_b101_1_0 (.A(imd_wire101_1_0),.Y(wire101_1_0));
NANDC2x1 inst_and_b101_1_1 (.A(A6),.B(wire101_0_2),.Y(imd_wire101_1_1));
INVC inst_inv_b101_1_1 (.A(imd_wire101_1_1),.Y(wire101_1_1));
NANDC2x1 inst_and_b101_2_0 (.A(wire101_1_0),.B(wire101_1_1),.Y(imd_Y101));
INVC inst_inv_b101_2_0 (.A(imd_Y101),.Y(Y101));
NANDC2x1 inst_clockedAND_b101_101 (.A(CLK),.B(Y101),.Y(imd_YF101));
INVC inst_clockedinv_b101_101 (.A(imd_YF101),.Y(YF101));


NANDC2x1 inst_and_b102_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire102_0_0));
INVC inst_inv_b102_0_0 (.A(imd_wire102_0_0),.Y(wire102_0_0));
NANDC2x1 inst_and_b102_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire102_0_1));
INVC inst_inv_b102_0_1 (.A(imd_wire102_0_1),.Y(wire102_0_1));
NANDC2x1 inst_and_b102_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire102_0_2));
INVC inst_inv_b102_0_2 (.A(imd_wire102_0_2),.Y(wire102_0_2));
NANDC2x1 inst_and_b102_1_0 (.A(wire102_0_0),.B(wire102_0_1),.Y(imd_wire102_1_0));
INVC inst_inv_b102_1_0 (.A(imd_wire102_1_0),.Y(wire102_1_0));
NANDC2x1 inst_and_b102_1_1 (.A(A6),.B(wire102_0_2),.Y(imd_wire102_1_1));
INVC inst_inv_b102_1_1 (.A(imd_wire102_1_1),.Y(wire102_1_1));
NANDC2x1 inst_and_b102_2_0 (.A(wire102_1_0),.B(wire102_1_1),.Y(imd_Y102));
INVC inst_inv_b102_2_0 (.A(imd_Y102),.Y(Y102));
NANDC2x1 inst_clockedAND_b102_102 (.A(CLK),.B(Y102),.Y(imd_YF102));
INVC inst_clockedinv_b102_102 (.A(imd_YF102),.Y(YF102));


NANDC2x1 inst_and_b103_0_0 (.A(A0),.B(A1),.Y(imd_wire103_0_0));
INVC inst_inv_b103_0_0 (.A(imd_wire103_0_0),.Y(wire103_0_0));
NANDC2x1 inst_and_b103_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire103_0_1));
INVC inst_inv_b103_0_1 (.A(imd_wire103_0_1),.Y(wire103_0_1));
NANDC2x1 inst_and_b103_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire103_0_2));
INVC inst_inv_b103_0_2 (.A(imd_wire103_0_2),.Y(wire103_0_2));
NANDC2x1 inst_and_b103_1_0 (.A(wire103_0_0),.B(wire103_0_1),.Y(imd_wire103_1_0));
INVC inst_inv_b103_1_0 (.A(imd_wire103_1_0),.Y(wire103_1_0));
NANDC2x1 inst_and_b103_1_1 (.A(A6),.B(wire103_0_2),.Y(imd_wire103_1_1));
INVC inst_inv_b103_1_1 (.A(imd_wire103_1_1),.Y(wire103_1_1));
NANDC2x1 inst_and_b103_2_0 (.A(wire103_1_0),.B(wire103_1_1),.Y(imd_Y103));
INVC inst_inv_b103_2_0 (.A(imd_Y103),.Y(Y103));
NANDC2x1 inst_clockedAND_b103_103 (.A(CLK),.B(Y103),.Y(imd_YF103));
INVC inst_clockedinv_b103_103 (.A(imd_YF103),.Y(YF103));


NANDC2x1 inst_and_b104_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire104_0_0));
INVC inst_inv_b104_0_0 (.A(imd_wire104_0_0),.Y(wire104_0_0));
NANDC2x1 inst_and_b104_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire104_0_1));
INVC inst_inv_b104_0_1 (.A(imd_wire104_0_1),.Y(wire104_0_1));
NANDC2x1 inst_and_b104_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire104_0_2));
INVC inst_inv_b104_0_2 (.A(imd_wire104_0_2),.Y(wire104_0_2));
NANDC2x1 inst_and_b104_1_0 (.A(wire104_0_0),.B(wire104_0_1),.Y(imd_wire104_1_0));
INVC inst_inv_b104_1_0 (.A(imd_wire104_1_0),.Y(wire104_1_0));
NANDC2x1 inst_and_b104_1_1 (.A(A6),.B(wire104_0_2),.Y(imd_wire104_1_1));
INVC inst_inv_b104_1_1 (.A(imd_wire104_1_1),.Y(wire104_1_1));
NANDC2x1 inst_and_b104_2_0 (.A(wire104_1_0),.B(wire104_1_1),.Y(imd_Y104));
INVC inst_inv_b104_2_0 (.A(imd_Y104),.Y(Y104));
NANDC2x1 inst_clockedAND_b104_104 (.A(CLK),.B(Y104),.Y(imd_YF104));
INVC inst_clockedinv_b104_104 (.A(imd_YF104),.Y(YF104));


NANDC2x1 inst_and_b105_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire105_0_0));
INVC inst_inv_b105_0_0 (.A(imd_wire105_0_0),.Y(wire105_0_0));
NANDC2x1 inst_and_b105_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire105_0_1));
INVC inst_inv_b105_0_1 (.A(imd_wire105_0_1),.Y(wire105_0_1));
NANDC2x1 inst_and_b105_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire105_0_2));
INVC inst_inv_b105_0_2 (.A(imd_wire105_0_2),.Y(wire105_0_2));
NANDC2x1 inst_and_b105_1_0 (.A(wire105_0_0),.B(wire105_0_1),.Y(imd_wire105_1_0));
INVC inst_inv_b105_1_0 (.A(imd_wire105_1_0),.Y(wire105_1_0));
NANDC2x1 inst_and_b105_1_1 (.A(A6),.B(wire105_0_2),.Y(imd_wire105_1_1));
INVC inst_inv_b105_1_1 (.A(imd_wire105_1_1),.Y(wire105_1_1));
NANDC2x1 inst_and_b105_2_0 (.A(wire105_1_0),.B(wire105_1_1),.Y(imd_Y105));
INVC inst_inv_b105_2_0 (.A(imd_Y105),.Y(Y105));
NANDC2x1 inst_clockedAND_b105_105 (.A(CLK),.B(Y105),.Y(imd_YF105));
INVC inst_clockedinv_b105_105 (.A(imd_YF105),.Y(YF105));


NANDC2x1 inst_and_b106_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire106_0_0));
INVC inst_inv_b106_0_0 (.A(imd_wire106_0_0),.Y(wire106_0_0));
NANDC2x1 inst_and_b106_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire106_0_1));
INVC inst_inv_b106_0_1 (.A(imd_wire106_0_1),.Y(wire106_0_1));
NANDC2x1 inst_and_b106_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire106_0_2));
INVC inst_inv_b106_0_2 (.A(imd_wire106_0_2),.Y(wire106_0_2));
NANDC2x1 inst_and_b106_1_0 (.A(wire106_0_0),.B(wire106_0_1),.Y(imd_wire106_1_0));
INVC inst_inv_b106_1_0 (.A(imd_wire106_1_0),.Y(wire106_1_0));
NANDC2x1 inst_and_b106_1_1 (.A(A6),.B(wire106_0_2),.Y(imd_wire106_1_1));
INVC inst_inv_b106_1_1 (.A(imd_wire106_1_1),.Y(wire106_1_1));
NANDC2x1 inst_and_b106_2_0 (.A(wire106_1_0),.B(wire106_1_1),.Y(imd_Y106));
INVC inst_inv_b106_2_0 (.A(imd_Y106),.Y(Y106));
NANDC2x1 inst_clockedAND_b106_106 (.A(CLK),.B(Y106),.Y(imd_YF106));
INVC inst_clockedinv_b106_106 (.A(imd_YF106),.Y(YF106));


NANDC2x1 inst_and_b107_0_0 (.A(A0),.B(A1),.Y(imd_wire107_0_0));
INVC inst_inv_b107_0_0 (.A(imd_wire107_0_0),.Y(wire107_0_0));
NANDC2x1 inst_and_b107_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire107_0_1));
INVC inst_inv_b107_0_1 (.A(imd_wire107_0_1),.Y(wire107_0_1));
NANDC2x1 inst_and_b107_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire107_0_2));
INVC inst_inv_b107_0_2 (.A(imd_wire107_0_2),.Y(wire107_0_2));
NANDC2x1 inst_and_b107_1_0 (.A(wire107_0_0),.B(wire107_0_1),.Y(imd_wire107_1_0));
INVC inst_inv_b107_1_0 (.A(imd_wire107_1_0),.Y(wire107_1_0));
NANDC2x1 inst_and_b107_1_1 (.A(A6),.B(wire107_0_2),.Y(imd_wire107_1_1));
INVC inst_inv_b107_1_1 (.A(imd_wire107_1_1),.Y(wire107_1_1));
NANDC2x1 inst_and_b107_2_0 (.A(wire107_1_0),.B(wire107_1_1),.Y(imd_Y107));
INVC inst_inv_b107_2_0 (.A(imd_Y107),.Y(Y107));
NANDC2x1 inst_clockedAND_b107_107 (.A(CLK),.B(Y107),.Y(imd_YF107));
INVC inst_clockedinv_b107_107 (.A(imd_YF107),.Y(YF107));


NANDC2x1 inst_and_b108_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire108_0_0));
INVC inst_inv_b108_0_0 (.A(imd_wire108_0_0),.Y(wire108_0_0));
NANDC2x1 inst_and_b108_0_1 (.A(A2),.B(A3),.Y(imd_wire108_0_1));
INVC inst_inv_b108_0_1 (.A(imd_wire108_0_1),.Y(wire108_0_1));
NANDC2x1 inst_and_b108_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire108_0_2));
INVC inst_inv_b108_0_2 (.A(imd_wire108_0_2),.Y(wire108_0_2));
NANDC2x1 inst_and_b108_1_0 (.A(wire108_0_0),.B(wire108_0_1),.Y(imd_wire108_1_0));
INVC inst_inv_b108_1_0 (.A(imd_wire108_1_0),.Y(wire108_1_0));
NANDC2x1 inst_and_b108_1_1 (.A(A6),.B(wire108_0_2),.Y(imd_wire108_1_1));
INVC inst_inv_b108_1_1 (.A(imd_wire108_1_1),.Y(wire108_1_1));
NANDC2x1 inst_and_b108_2_0 (.A(wire108_1_0),.B(wire108_1_1),.Y(imd_Y108));
INVC inst_inv_b108_2_0 (.A(imd_Y108),.Y(Y108));
NANDC2x1 inst_clockedAND_b108_108 (.A(CLK),.B(Y108),.Y(imd_YF108));
INVC inst_clockedinv_b108_108 (.A(imd_YF108),.Y(YF108));


NANDC2x1 inst_and_b109_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire109_0_0));
INVC inst_inv_b109_0_0 (.A(imd_wire109_0_0),.Y(wire109_0_0));
NANDC2x1 inst_and_b109_0_1 (.A(A2),.B(A3),.Y(imd_wire109_0_1));
INVC inst_inv_b109_0_1 (.A(imd_wire109_0_1),.Y(wire109_0_1));
NANDC2x1 inst_and_b109_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire109_0_2));
INVC inst_inv_b109_0_2 (.A(imd_wire109_0_2),.Y(wire109_0_2));
NANDC2x1 inst_and_b109_1_0 (.A(wire109_0_0),.B(wire109_0_1),.Y(imd_wire109_1_0));
INVC inst_inv_b109_1_0 (.A(imd_wire109_1_0),.Y(wire109_1_0));
NANDC2x1 inst_and_b109_1_1 (.A(A6),.B(wire109_0_2),.Y(imd_wire109_1_1));
INVC inst_inv_b109_1_1 (.A(imd_wire109_1_1),.Y(wire109_1_1));
NANDC2x1 inst_and_b109_2_0 (.A(wire109_1_0),.B(wire109_1_1),.Y(imd_Y109));
INVC inst_inv_b109_2_0 (.A(imd_Y109),.Y(Y109));
NANDC2x1 inst_clockedAND_b109_109 (.A(CLK),.B(Y109),.Y(imd_YF109));
INVC inst_clockedinv_b109_109 (.A(imd_YF109),.Y(YF109));


NANDC2x1 inst_and_b110_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire110_0_0));
INVC inst_inv_b110_0_0 (.A(imd_wire110_0_0),.Y(wire110_0_0));
NANDC2x1 inst_and_b110_0_1 (.A(A2),.B(A3),.Y(imd_wire110_0_1));
INVC inst_inv_b110_0_1 (.A(imd_wire110_0_1),.Y(wire110_0_1));
NANDC2x1 inst_and_b110_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire110_0_2));
INVC inst_inv_b110_0_2 (.A(imd_wire110_0_2),.Y(wire110_0_2));
NANDC2x1 inst_and_b110_1_0 (.A(wire110_0_0),.B(wire110_0_1),.Y(imd_wire110_1_0));
INVC inst_inv_b110_1_0 (.A(imd_wire110_1_0),.Y(wire110_1_0));
NANDC2x1 inst_and_b110_1_1 (.A(A6),.B(wire110_0_2),.Y(imd_wire110_1_1));
INVC inst_inv_b110_1_1 (.A(imd_wire110_1_1),.Y(wire110_1_1));
NANDC2x1 inst_and_b110_2_0 (.A(wire110_1_0),.B(wire110_1_1),.Y(imd_Y110));
INVC inst_inv_b110_2_0 (.A(imd_Y110),.Y(Y110));
NANDC2x1 inst_clockedAND_b110_110 (.A(CLK),.B(Y110),.Y(imd_YF110));
INVC inst_clockedinv_b110_110 (.A(imd_YF110),.Y(YF110));


NANDC2x1 inst_and_b111_0_0 (.A(A0),.B(A1),.Y(imd_wire111_0_0));
INVC inst_inv_b111_0_0 (.A(imd_wire111_0_0),.Y(wire111_0_0));
NANDC2x1 inst_and_b111_0_1 (.A(A2),.B(A3),.Y(imd_wire111_0_1));
INVC inst_inv_b111_0_1 (.A(imd_wire111_0_1),.Y(wire111_0_1));
NANDC2x1 inst_and_b111_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire111_0_2));
INVC inst_inv_b111_0_2 (.A(imd_wire111_0_2),.Y(wire111_0_2));
NANDC2x1 inst_and_b111_1_0 (.A(wire111_0_0),.B(wire111_0_1),.Y(imd_wire111_1_0));
INVC inst_inv_b111_1_0 (.A(imd_wire111_1_0),.Y(wire111_1_0));
NANDC2x1 inst_and_b111_1_1 (.A(A6),.B(wire111_0_2),.Y(imd_wire111_1_1));
INVC inst_inv_b111_1_1 (.A(imd_wire111_1_1),.Y(wire111_1_1));
NANDC2x1 inst_and_b111_2_0 (.A(wire111_1_0),.B(wire111_1_1),.Y(imd_Y111));
INVC inst_inv_b111_2_0 (.A(imd_Y111),.Y(Y111));
NANDC2x1 inst_clockedAND_b111_111 (.A(CLK),.B(Y111),.Y(imd_YF111));
INVC inst_clockedinv_b111_111 (.A(imd_YF111),.Y(YF111));


NANDC2x1 inst_and_b112_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire112_0_0));
INVC inst_inv_b112_0_0 (.A(imd_wire112_0_0),.Y(wire112_0_0));
NANDC2x1 inst_and_b112_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire112_0_1));
INVC inst_inv_b112_0_1 (.A(imd_wire112_0_1),.Y(wire112_0_1));
NANDC2x1 inst_and_b112_0_2 (.A(A4),.B(A5),.Y(imd_wire112_0_2));
INVC inst_inv_b112_0_2 (.A(imd_wire112_0_2),.Y(wire112_0_2));
NANDC2x1 inst_and_b112_1_0 (.A(wire112_0_0),.B(wire112_0_1),.Y(imd_wire112_1_0));
INVC inst_inv_b112_1_0 (.A(imd_wire112_1_0),.Y(wire112_1_0));
NANDC2x1 inst_and_b112_1_1 (.A(A6),.B(wire112_0_2),.Y(imd_wire112_1_1));
INVC inst_inv_b112_1_1 (.A(imd_wire112_1_1),.Y(wire112_1_1));
NANDC2x1 inst_and_b112_2_0 (.A(wire112_1_0),.B(wire112_1_1),.Y(imd_Y112));
INVC inst_inv_b112_2_0 (.A(imd_Y112),.Y(Y112));
NANDC2x1 inst_clockedAND_b112_112 (.A(CLK),.B(Y112),.Y(imd_YF112));
INVC inst_clockedinv_b112_112 (.A(imd_YF112),.Y(YF112));


NANDC2x1 inst_and_b113_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire113_0_0));
INVC inst_inv_b113_0_0 (.A(imd_wire113_0_0),.Y(wire113_0_0));
NANDC2x1 inst_and_b113_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire113_0_1));
INVC inst_inv_b113_0_1 (.A(imd_wire113_0_1),.Y(wire113_0_1));
NANDC2x1 inst_and_b113_0_2 (.A(A4),.B(A5),.Y(imd_wire113_0_2));
INVC inst_inv_b113_0_2 (.A(imd_wire113_0_2),.Y(wire113_0_2));
NANDC2x1 inst_and_b113_1_0 (.A(wire113_0_0),.B(wire113_0_1),.Y(imd_wire113_1_0));
INVC inst_inv_b113_1_0 (.A(imd_wire113_1_0),.Y(wire113_1_0));
NANDC2x1 inst_and_b113_1_1 (.A(A6),.B(wire113_0_2),.Y(imd_wire113_1_1));
INVC inst_inv_b113_1_1 (.A(imd_wire113_1_1),.Y(wire113_1_1));
NANDC2x1 inst_and_b113_2_0 (.A(wire113_1_0),.B(wire113_1_1),.Y(imd_Y113));
INVC inst_inv_b113_2_0 (.A(imd_Y113),.Y(Y113));
NANDC2x1 inst_clockedAND_b113_113 (.A(CLK),.B(Y113),.Y(imd_YF113));
INVC inst_clockedinv_b113_113 (.A(imd_YF113),.Y(YF113));


NANDC2x1 inst_and_b114_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire114_0_0));
INVC inst_inv_b114_0_0 (.A(imd_wire114_0_0),.Y(wire114_0_0));
NANDC2x1 inst_and_b114_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire114_0_1));
INVC inst_inv_b114_0_1 (.A(imd_wire114_0_1),.Y(wire114_0_1));
NANDC2x1 inst_and_b114_0_2 (.A(A4),.B(A5),.Y(imd_wire114_0_2));
INVC inst_inv_b114_0_2 (.A(imd_wire114_0_2),.Y(wire114_0_2));
NANDC2x1 inst_and_b114_1_0 (.A(wire114_0_0),.B(wire114_0_1),.Y(imd_wire114_1_0));
INVC inst_inv_b114_1_0 (.A(imd_wire114_1_0),.Y(wire114_1_0));
NANDC2x1 inst_and_b114_1_1 (.A(A6),.B(wire114_0_2),.Y(imd_wire114_1_1));
INVC inst_inv_b114_1_1 (.A(imd_wire114_1_1),.Y(wire114_1_1));
NANDC2x1 inst_and_b114_2_0 (.A(wire114_1_0),.B(wire114_1_1),.Y(imd_Y114));
INVC inst_inv_b114_2_0 (.A(imd_Y114),.Y(Y114));
NANDC2x1 inst_clockedAND_b114_114 (.A(CLK),.B(Y114),.Y(imd_YF114));
INVC inst_clockedinv_b114_114 (.A(imd_YF114),.Y(YF114));


NANDC2x1 inst_and_b115_0_0 (.A(A0),.B(A1),.Y(imd_wire115_0_0));
INVC inst_inv_b115_0_0 (.A(imd_wire115_0_0),.Y(wire115_0_0));
NANDC2x1 inst_and_b115_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire115_0_1));
INVC inst_inv_b115_0_1 (.A(imd_wire115_0_1),.Y(wire115_0_1));
NANDC2x1 inst_and_b115_0_2 (.A(A4),.B(A5),.Y(imd_wire115_0_2));
INVC inst_inv_b115_0_2 (.A(imd_wire115_0_2),.Y(wire115_0_2));
NANDC2x1 inst_and_b115_1_0 (.A(wire115_0_0),.B(wire115_0_1),.Y(imd_wire115_1_0));
INVC inst_inv_b115_1_0 (.A(imd_wire115_1_0),.Y(wire115_1_0));
NANDC2x1 inst_and_b115_1_1 (.A(A6),.B(wire115_0_2),.Y(imd_wire115_1_1));
INVC inst_inv_b115_1_1 (.A(imd_wire115_1_1),.Y(wire115_1_1));
NANDC2x1 inst_and_b115_2_0 (.A(wire115_1_0),.B(wire115_1_1),.Y(imd_Y115));
INVC inst_inv_b115_2_0 (.A(imd_Y115),.Y(Y115));
NANDC2x1 inst_clockedAND_b115_115 (.A(CLK),.B(Y115),.Y(imd_YF115));
INVC inst_clockedinv_b115_115 (.A(imd_YF115),.Y(YF115));


NANDC2x1 inst_and_b116_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire116_0_0));
INVC inst_inv_b116_0_0 (.A(imd_wire116_0_0),.Y(wire116_0_0));
NANDC2x1 inst_and_b116_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire116_0_1));
INVC inst_inv_b116_0_1 (.A(imd_wire116_0_1),.Y(wire116_0_1));
NANDC2x1 inst_and_b116_0_2 (.A(A4),.B(A5),.Y(imd_wire116_0_2));
INVC inst_inv_b116_0_2 (.A(imd_wire116_0_2),.Y(wire116_0_2));
NANDC2x1 inst_and_b116_1_0 (.A(wire116_0_0),.B(wire116_0_1),.Y(imd_wire116_1_0));
INVC inst_inv_b116_1_0 (.A(imd_wire116_1_0),.Y(wire116_1_0));
NANDC2x1 inst_and_b116_1_1 (.A(A6),.B(wire116_0_2),.Y(imd_wire116_1_1));
INVC inst_inv_b116_1_1 (.A(imd_wire116_1_1),.Y(wire116_1_1));
NANDC2x1 inst_and_b116_2_0 (.A(wire116_1_0),.B(wire116_1_1),.Y(imd_Y116));
INVC inst_inv_b116_2_0 (.A(imd_Y116),.Y(Y116));
NANDC2x1 inst_clockedAND_b116_116 (.A(CLK),.B(Y116),.Y(imd_YF116));
INVC inst_clockedinv_b116_116 (.A(imd_YF116),.Y(YF116));


NANDC2x1 inst_and_b117_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire117_0_0));
INVC inst_inv_b117_0_0 (.A(imd_wire117_0_0),.Y(wire117_0_0));
NANDC2x1 inst_and_b117_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire117_0_1));
INVC inst_inv_b117_0_1 (.A(imd_wire117_0_1),.Y(wire117_0_1));
NANDC2x1 inst_and_b117_0_2 (.A(A4),.B(A5),.Y(imd_wire117_0_2));
INVC inst_inv_b117_0_2 (.A(imd_wire117_0_2),.Y(wire117_0_2));
NANDC2x1 inst_and_b117_1_0 (.A(wire117_0_0),.B(wire117_0_1),.Y(imd_wire117_1_0));
INVC inst_inv_b117_1_0 (.A(imd_wire117_1_0),.Y(wire117_1_0));
NANDC2x1 inst_and_b117_1_1 (.A(A6),.B(wire117_0_2),.Y(imd_wire117_1_1));
INVC inst_inv_b117_1_1 (.A(imd_wire117_1_1),.Y(wire117_1_1));
NANDC2x1 inst_and_b117_2_0 (.A(wire117_1_0),.B(wire117_1_1),.Y(imd_Y117));
INVC inst_inv_b117_2_0 (.A(imd_Y117),.Y(Y117));
NANDC2x1 inst_clockedAND_b117_117 (.A(CLK),.B(Y117),.Y(imd_YF117));
INVC inst_clockedinv_b117_117 (.A(imd_YF117),.Y(YF117));


NANDC2x1 inst_and_b118_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire118_0_0));
INVC inst_inv_b118_0_0 (.A(imd_wire118_0_0),.Y(wire118_0_0));
NANDC2x1 inst_and_b118_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire118_0_1));
INVC inst_inv_b118_0_1 (.A(imd_wire118_0_1),.Y(wire118_0_1));
NANDC2x1 inst_and_b118_0_2 (.A(A4),.B(A5),.Y(imd_wire118_0_2));
INVC inst_inv_b118_0_2 (.A(imd_wire118_0_2),.Y(wire118_0_2));
NANDC2x1 inst_and_b118_1_0 (.A(wire118_0_0),.B(wire118_0_1),.Y(imd_wire118_1_0));
INVC inst_inv_b118_1_0 (.A(imd_wire118_1_0),.Y(wire118_1_0));
NANDC2x1 inst_and_b118_1_1 (.A(A6),.B(wire118_0_2),.Y(imd_wire118_1_1));
INVC inst_inv_b118_1_1 (.A(imd_wire118_1_1),.Y(wire118_1_1));
NANDC2x1 inst_and_b118_2_0 (.A(wire118_1_0),.B(wire118_1_1),.Y(imd_Y118));
INVC inst_inv_b118_2_0 (.A(imd_Y118),.Y(Y118));
NANDC2x1 inst_clockedAND_b118_118 (.A(CLK),.B(Y118),.Y(imd_YF118));
INVC inst_clockedinv_b118_118 (.A(imd_YF118),.Y(YF118));


NANDC2x1 inst_and_b119_0_0 (.A(A0),.B(A1),.Y(imd_wire119_0_0));
INVC inst_inv_b119_0_0 (.A(imd_wire119_0_0),.Y(wire119_0_0));
NANDC2x1 inst_and_b119_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire119_0_1));
INVC inst_inv_b119_0_1 (.A(imd_wire119_0_1),.Y(wire119_0_1));
NANDC2x1 inst_and_b119_0_2 (.A(A4),.B(A5),.Y(imd_wire119_0_2));
INVC inst_inv_b119_0_2 (.A(imd_wire119_0_2),.Y(wire119_0_2));
NANDC2x1 inst_and_b119_1_0 (.A(wire119_0_0),.B(wire119_0_1),.Y(imd_wire119_1_0));
INVC inst_inv_b119_1_0 (.A(imd_wire119_1_0),.Y(wire119_1_0));
NANDC2x1 inst_and_b119_1_1 (.A(A6),.B(wire119_0_2),.Y(imd_wire119_1_1));
INVC inst_inv_b119_1_1 (.A(imd_wire119_1_1),.Y(wire119_1_1));
NANDC2x1 inst_and_b119_2_0 (.A(wire119_1_0),.B(wire119_1_1),.Y(imd_Y119));
INVC inst_inv_b119_2_0 (.A(imd_Y119),.Y(Y119));
NANDC2x1 inst_clockedAND_b119_119 (.A(CLK),.B(Y119),.Y(imd_YF119));
INVC inst_clockedinv_b119_119 (.A(imd_YF119),.Y(YF119));


NANDC2x1 inst_and_b120_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire120_0_0));
INVC inst_inv_b120_0_0 (.A(imd_wire120_0_0),.Y(wire120_0_0));
NANDC2x1 inst_and_b120_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire120_0_1));
INVC inst_inv_b120_0_1 (.A(imd_wire120_0_1),.Y(wire120_0_1));
NANDC2x1 inst_and_b120_0_2 (.A(A4),.B(A5),.Y(imd_wire120_0_2));
INVC inst_inv_b120_0_2 (.A(imd_wire120_0_2),.Y(wire120_0_2));
NANDC2x1 inst_and_b120_1_0 (.A(wire120_0_0),.B(wire120_0_1),.Y(imd_wire120_1_0));
INVC inst_inv_b120_1_0 (.A(imd_wire120_1_0),.Y(wire120_1_0));
NANDC2x1 inst_and_b120_1_1 (.A(A6),.B(wire120_0_2),.Y(imd_wire120_1_1));
INVC inst_inv_b120_1_1 (.A(imd_wire120_1_1),.Y(wire120_1_1));
NANDC2x1 inst_and_b120_2_0 (.A(wire120_1_0),.B(wire120_1_1),.Y(imd_Y120));
INVC inst_inv_b120_2_0 (.A(imd_Y120),.Y(Y120));
NANDC2x1 inst_clockedAND_b120_120 (.A(CLK),.B(Y120),.Y(imd_YF120));
INVC inst_clockedinv_b120_120 (.A(imd_YF120),.Y(YF120));


NANDC2x1 inst_and_b121_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire121_0_0));
INVC inst_inv_b121_0_0 (.A(imd_wire121_0_0),.Y(wire121_0_0));
NANDC2x1 inst_and_b121_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire121_0_1));
INVC inst_inv_b121_0_1 (.A(imd_wire121_0_1),.Y(wire121_0_1));
NANDC2x1 inst_and_b121_0_2 (.A(A4),.B(A5),.Y(imd_wire121_0_2));
INVC inst_inv_b121_0_2 (.A(imd_wire121_0_2),.Y(wire121_0_2));
NANDC2x1 inst_and_b121_1_0 (.A(wire121_0_0),.B(wire121_0_1),.Y(imd_wire121_1_0));
INVC inst_inv_b121_1_0 (.A(imd_wire121_1_0),.Y(wire121_1_0));
NANDC2x1 inst_and_b121_1_1 (.A(A6),.B(wire121_0_2),.Y(imd_wire121_1_1));
INVC inst_inv_b121_1_1 (.A(imd_wire121_1_1),.Y(wire121_1_1));
NANDC2x1 inst_and_b121_2_0 (.A(wire121_1_0),.B(wire121_1_1),.Y(imd_Y121));
INVC inst_inv_b121_2_0 (.A(imd_Y121),.Y(Y121));
NANDC2x1 inst_clockedAND_b121_121 (.A(CLK),.B(Y121),.Y(imd_YF121));
INVC inst_clockedinv_b121_121 (.A(imd_YF121),.Y(YF121));


NANDC2x1 inst_and_b122_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire122_0_0));
INVC inst_inv_b122_0_0 (.A(imd_wire122_0_0),.Y(wire122_0_0));
NANDC2x1 inst_and_b122_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire122_0_1));
INVC inst_inv_b122_0_1 (.A(imd_wire122_0_1),.Y(wire122_0_1));
NANDC2x1 inst_and_b122_0_2 (.A(A4),.B(A5),.Y(imd_wire122_0_2));
INVC inst_inv_b122_0_2 (.A(imd_wire122_0_2),.Y(wire122_0_2));
NANDC2x1 inst_and_b122_1_0 (.A(wire122_0_0),.B(wire122_0_1),.Y(imd_wire122_1_0));
INVC inst_inv_b122_1_0 (.A(imd_wire122_1_0),.Y(wire122_1_0));
NANDC2x1 inst_and_b122_1_1 (.A(A6),.B(wire122_0_2),.Y(imd_wire122_1_1));
INVC inst_inv_b122_1_1 (.A(imd_wire122_1_1),.Y(wire122_1_1));
NANDC2x1 inst_and_b122_2_0 (.A(wire122_1_0),.B(wire122_1_1),.Y(imd_Y122));
INVC inst_inv_b122_2_0 (.A(imd_Y122),.Y(Y122));
NANDC2x1 inst_clockedAND_b122_122 (.A(CLK),.B(Y122),.Y(imd_YF122));
INVC inst_clockedinv_b122_122 (.A(imd_YF122),.Y(YF122));


NANDC2x1 inst_and_b123_0_0 (.A(A0),.B(A1),.Y(imd_wire123_0_0));
INVC inst_inv_b123_0_0 (.A(imd_wire123_0_0),.Y(wire123_0_0));
NANDC2x1 inst_and_b123_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire123_0_1));
INVC inst_inv_b123_0_1 (.A(imd_wire123_0_1),.Y(wire123_0_1));
NANDC2x1 inst_and_b123_0_2 (.A(A4),.B(A5),.Y(imd_wire123_0_2));
INVC inst_inv_b123_0_2 (.A(imd_wire123_0_2),.Y(wire123_0_2));
NANDC2x1 inst_and_b123_1_0 (.A(wire123_0_0),.B(wire123_0_1),.Y(imd_wire123_1_0));
INVC inst_inv_b123_1_0 (.A(imd_wire123_1_0),.Y(wire123_1_0));
NANDC2x1 inst_and_b123_1_1 (.A(A6),.B(wire123_0_2),.Y(imd_wire123_1_1));
INVC inst_inv_b123_1_1 (.A(imd_wire123_1_1),.Y(wire123_1_1));
NANDC2x1 inst_and_b123_2_0 (.A(wire123_1_0),.B(wire123_1_1),.Y(imd_Y123));
INVC inst_inv_b123_2_0 (.A(imd_Y123),.Y(Y123));
NANDC2x1 inst_clockedAND_b123_123 (.A(CLK),.B(Y123),.Y(imd_YF123));
INVC inst_clockedinv_b123_123 (.A(imd_YF123),.Y(YF123));


NANDC2x1 inst_and_b124_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire124_0_0));
INVC inst_inv_b124_0_0 (.A(imd_wire124_0_0),.Y(wire124_0_0));
NANDC2x1 inst_and_b124_0_1 (.A(A2),.B(A3),.Y(imd_wire124_0_1));
INVC inst_inv_b124_0_1 (.A(imd_wire124_0_1),.Y(wire124_0_1));
NANDC2x1 inst_and_b124_0_2 (.A(A4),.B(A5),.Y(imd_wire124_0_2));
INVC inst_inv_b124_0_2 (.A(imd_wire124_0_2),.Y(wire124_0_2));
NANDC2x1 inst_and_b124_1_0 (.A(wire124_0_0),.B(wire124_0_1),.Y(imd_wire124_1_0));
INVC inst_inv_b124_1_0 (.A(imd_wire124_1_0),.Y(wire124_1_0));
NANDC2x1 inst_and_b124_1_1 (.A(A6),.B(wire124_0_2),.Y(imd_wire124_1_1));
INVC inst_inv_b124_1_1 (.A(imd_wire124_1_1),.Y(wire124_1_1));
NANDC2x1 inst_and_b124_2_0 (.A(wire124_1_0),.B(wire124_1_1),.Y(imd_Y124));
INVC inst_inv_b124_2_0 (.A(imd_Y124),.Y(Y124));
NANDC2x1 inst_clockedAND_b124_124 (.A(CLK),.B(Y124),.Y(imd_YF124));
INVC inst_clockedinv_b124_124 (.A(imd_YF124),.Y(YF124));


NANDC2x1 inst_and_b125_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire125_0_0));
INVC inst_inv_b125_0_0 (.A(imd_wire125_0_0),.Y(wire125_0_0));
NANDC2x1 inst_and_b125_0_1 (.A(A2),.B(A3),.Y(imd_wire125_0_1));
INVC inst_inv_b125_0_1 (.A(imd_wire125_0_1),.Y(wire125_0_1));
NANDC2x1 inst_and_b125_0_2 (.A(A4),.B(A5),.Y(imd_wire125_0_2));
INVC inst_inv_b125_0_2 (.A(imd_wire125_0_2),.Y(wire125_0_2));
NANDC2x1 inst_and_b125_1_0 (.A(wire125_0_0),.B(wire125_0_1),.Y(imd_wire125_1_0));
INVC inst_inv_b125_1_0 (.A(imd_wire125_1_0),.Y(wire125_1_0));
NANDC2x1 inst_and_b125_1_1 (.A(A6),.B(wire125_0_2),.Y(imd_wire125_1_1));
INVC inst_inv_b125_1_1 (.A(imd_wire125_1_1),.Y(wire125_1_1));
NANDC2x1 inst_and_b125_2_0 (.A(wire125_1_0),.B(wire125_1_1),.Y(imd_Y125));
INVC inst_inv_b125_2_0 (.A(imd_Y125),.Y(Y125));
NANDC2x1 inst_clockedAND_b125_125 (.A(CLK),.B(Y125),.Y(imd_YF125));
INVC inst_clockedinv_b125_125 (.A(imd_YF125),.Y(YF125));


NANDC2x1 inst_and_b126_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire126_0_0));
INVC inst_inv_b126_0_0 (.A(imd_wire126_0_0),.Y(wire126_0_0));
NANDC2x1 inst_and_b126_0_1 (.A(A2),.B(A3),.Y(imd_wire126_0_1));
INVC inst_inv_b126_0_1 (.A(imd_wire126_0_1),.Y(wire126_0_1));
NANDC2x1 inst_and_b126_0_2 (.A(A4),.B(A5),.Y(imd_wire126_0_2));
INVC inst_inv_b126_0_2 (.A(imd_wire126_0_2),.Y(wire126_0_2));
NANDC2x1 inst_and_b126_1_0 (.A(wire126_0_0),.B(wire126_0_1),.Y(imd_wire126_1_0));
INVC inst_inv_b126_1_0 (.A(imd_wire126_1_0),.Y(wire126_1_0));
NANDC2x1 inst_and_b126_1_1 (.A(A6),.B(wire126_0_2),.Y(imd_wire126_1_1));
INVC inst_inv_b126_1_1 (.A(imd_wire126_1_1),.Y(wire126_1_1));
NANDC2x1 inst_and_b126_2_0 (.A(wire126_1_0),.B(wire126_1_1),.Y(imd_Y126));
INVC inst_inv_b126_2_0 (.A(imd_Y126),.Y(Y126));
NANDC2x1 inst_clockedAND_b126_126 (.A(CLK),.B(Y126),.Y(imd_YF126));
INVC inst_clockedinv_b126_126 (.A(imd_YF126),.Y(YF126));


NANDC2x1 inst_and_b127_0_0 (.A(A0),.B(A1),.Y(imd_wire127_0_0));
INVC inst_inv_b127_0_0 (.A(imd_wire127_0_0),.Y(wire127_0_0));
NANDC2x1 inst_and_b127_0_1 (.A(A2),.B(A3),.Y(imd_wire127_0_1));
INVC inst_inv_b127_0_1 (.A(imd_wire127_0_1),.Y(wire127_0_1));
NANDC2x1 inst_and_b127_0_2 (.A(A4),.B(A5),.Y(imd_wire127_0_2));
INVC inst_inv_b127_0_2 (.A(imd_wire127_0_2),.Y(wire127_0_2));
NANDC2x1 inst_and_b127_1_0 (.A(wire127_0_0),.B(wire127_0_1),.Y(imd_wire127_1_0));
INVC inst_inv_b127_1_0 (.A(imd_wire127_1_0),.Y(wire127_1_0));
NANDC2x1 inst_and_b127_1_1 (.A(A6),.B(wire127_0_2),.Y(imd_wire127_1_1));
INVC inst_inv_b127_1_1 (.A(imd_wire127_1_1),.Y(wire127_1_1));
NANDC2x1 inst_and_b127_2_0 (.A(wire127_1_0),.B(wire127_1_1),.Y(imd_Y127));
INVC inst_inv_b127_2_0 (.A(imd_Y127),.Y(Y127));
NANDC2x1 inst_clockedAND_b127_127 (.A(CLK),.B(Y127),.Y(imd_YF127));
INVC inst_clockedinv_b127_127 (.A(imd_YF127),.Y(YF127));


endmodule
module colDecoder(A0,A0_inv,A1,A1_inv,CLK,YF0,YF1,YF2,YF3);
input A0;
input A0_inv;
input A1;
input A1_inv;
input CLK;
output YF0;
output YF1;
output YF2;
output YF3;
NANDC2x1 inst_and_b0_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_Y0));
INVC inst_inv_b0_0_0 (.A(imd_Y0),.Y(Y0));
NANDC2x1 inst_clockedAND_b0_0 (.A(CLK),.B(Y0),.Y(imd_YF0));
INVC inst_clockedinv_b0_0 (.A(imd_YF0),.Y(YF0));


NANDC2x1 inst_and_b1_0_0 (.A(A0),.B(A1_inv),.Y(imd_Y1));
INVC inst_inv_b1_0_0 (.A(imd_Y1),.Y(Y1));
NANDC2x1 inst_clockedAND_b1_1 (.A(CLK),.B(Y1),.Y(imd_YF1));
INVC inst_clockedinv_b1_1 (.A(imd_YF1),.Y(YF1));


NANDC2x1 inst_and_b2_0_0 (.A(A0_inv),.B(A1),.Y(imd_Y2));
INVC inst_inv_b2_0_0 (.A(imd_Y2),.Y(Y2));
NANDC2x1 inst_clockedAND_b2_2 (.A(CLK),.B(Y2),.Y(imd_YF2));
INVC inst_clockedinv_b2_2 (.A(imd_YF2),.Y(YF2));


NANDC2x1 inst_and_b3_0_0 (.A(A0),.B(A1),.Y(imd_Y3));
INVC inst_inv_b3_0_0 (.A(imd_Y3),.Y(Y3));
NANDC2x1 inst_clockedAND_b3_3 (.A(CLK),.B(Y3),.Y(imd_YF3));
INVC inst_clockedinv_b3_3 (.A(imd_YF3),.Y(YF3));


endmodule
module columnMux(A0,Abar0,A1,Abar1,A2,Abar2,A3,Abar3,sel0,sel1,sel2,sel3,Y,Ybar);
input A0;
input Abar0;
input A1;
input Abar1;
input A2;
input Abar2;
input A3;
input Abar3;
input sel0;
input sel1;
input sel2;
input sel3;
output Y;
output Ybar;
muxTrans wire0 (.A(A0),.S(sel0),.Y(Y));
muxTrans wire1 (.A(Abar0),.S(sel0),.Y(Ybar));
muxTrans wire2 (.A(A1),.S(sel1),.Y(Y));
muxTrans wire3 (.A(Abar1),.S(sel1),.Y(Ybar));
muxTrans wire4 (.A(A2),.S(sel2),.Y(Y));
muxTrans wire5 (.A(Abar2),.S(sel2),.Y(Ybar));
muxTrans wire6 (.A(A3),.S(sel3),.Y(Y));
muxTrans wire7 (.A(Abar3),.S(sel3),.Y(Ybar));
endmodule
module sram_2kb_128x128x32(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,addr8,din0,din1,din2,din3,din4,din5,din6,din7,din8,din9,din10,din11,din12,din13,din14,din15,din16,din17,din18,din19,din20,din21,din22,din23,din24,din25,din26,din27,din28,din29,din30,din31,dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7,dout8,dout9,dout10,dout11,dout12,dout13,dout14,dout15,dout16,dout17,dout18,dout19,dout20,dout21,dout22,dout23,dout24,dout25,dout26,dout27,dout28,dout29,dout30,dout31,clk,write_en,sense_en);
input addr0;
input addr1;
input addr2;
input addr3;
input addr4;
input addr5;
input addr6;
input addr7;
input addr8;
input din0;
input din1;
input din2;
input din3;
input din4;
input din5;
input din6;
input din7;
input din8;
input din9;
input din10;
input din11;
input din12;
input din13;
input din14;
input din15;
input din16;
input din17;
input din18;
input din19;
input din20;
input din21;
input din22;
input din23;
input din24;
input din25;
input din26;
input din27;
input din28;
input din29;
input din30;
input din31;
output dout0;
output dout1;
output dout2;
output dout3;
output dout4;
output dout5;
output dout6;
output dout7;
output dout8;
output dout9;
output dout10;
output dout11;
output dout12;
output dout13;
output dout14;
output dout15;
output dout16;
output dout17;
output dout18;
output dout19;
output dout20;
output dout21;
output dout22;
output dout23;
output dout24;
output dout25;
output dout26;
output dout27;
output dout28;
output dout29;
output dout30;
output dout31;
input clk;
input write_en;
input sense_en;


specify

    (sense_en  => dout0  ) = 0.6;   
    (sense_en  => dout1  ) = 1.6;   
    (sense_en  => dout2  ) = 12.6;   
    (sense_en  => dout3  ) = 10.6;   
    (sense_en  => dout4  ) = 8.1;   
    (sense_en  => dout5  ) = 11.6;   
    (sense_en  => dout6  ) = 1.6;   
    (sense_en  => dout7  ) = 5.6;   
    (sense_en  => dout8  ) = 7.6;   
    (sense_en  => dout9  ) = 9.6;   
    (sense_en  => dout10 ) = 4.6;   
    (sense_en  => dout11 ) = 1.6; 
    (sense_en  => dout12 ) = 1.6;   
    (sense_en  => dout13 ) = 5;   
    (sense_en  => dout14 ) = 3;   
    (sense_en  => dout15 ) = 2;   
    (sense_en  => dout16 ) = 0.9;   
    (sense_en  => dout17 ) = 5; 
    (sense_en  => dout18 ) = 6;   
    (sense_en  => dout19 ) = 4;   
    (sense_en  => dout20 ) = 2;   
    (sense_en  => dout21 ) = 8;   
    (sense_en  => dout22 ) = 3;   
    (sense_en  => dout23 ) = 8;   
    (sense_en  => dout24 ) = 1;   
    (sense_en  => dout25 ) = 7;   
    (sense_en  => dout26 ) = 9.6;   
    (sense_en  => dout27 ) = 4.6;   
    (sense_en  => dout28 ) = 1.6;   
    (sense_en  => dout29 ) = 8.6; 
    (sense_en  => dout30 ) = 0;   
    (sense_en  => dout31 ) = 3.6;   

endspecify


inverter_compiler inst_invComp (.A0(clk),.A0_bar(clk_bar));
invRow inst_invRow(addr0,addr1,addr2,addr3,addr4,addr5,addr6,inv_addr0,inv_addr1,inv_addr2,inv_addr3,inv_addr4,inv_addr5,inv_addr6);
invCol inst_invCol(addr7,addr8,inv_addr7,inv_addr8);
rowDecoder inst_rowDec (addr0,inv_addr0,addr1,inv_addr1,addr2,inv_addr2,addr3,inv_addr3,addr4,inv_addr4,addr5,inv_addr5,addr6,inv_addr6,clk_bar,WL0,WL1,WL2,WL3,WL4,WL5,WL6,WL7,WL8,WL9,WL10,WL11,WL12,WL13,WL14,WL15,WL16,WL17,WL18,WL19,WL20,WL21,WL22,WL23,WL24,WL25,WL26,WL27,WL28,WL29,WL30,WL31,WL32,WL33,WL34,WL35,WL36,WL37,WL38,WL39,WL40,WL41,WL42,WL43,WL44,WL45,WL46,WL47,WL48,WL49,WL50,WL51,WL52,WL53,WL54,WL55,WL56,WL57,WL58,WL59,WL60,WL61,WL62,WL63,WL64,WL65,WL66,WL67,WL68,WL69,WL70,WL71,WL72,WL73,WL74,WL75,WL76,WL77,WL78,WL79,WL80,WL81,WL82,WL83,WL84,WL85,WL86,WL87,WL88,WL89,WL90,WL91,WL92,WL93,WL94,WL95,WL96,WL97,WL98,WL99,WL100,WL101,WL102,WL103,WL104,WL105,WL106,WL107,WL108,WL109,WL110,WL111,WL112,WL113,WL114,WL115,WL116,WL117,WL118,WL119,WL120,WL121,WL122,WL123,WL124,WL125,WL126,WL127);
colDecoder inst_colDec (addr7,inv_addr7,addr8,inv_addr8,clk_bar,SL0,SL1,SL2,SL3);
sram_cell_6t_5 inst_cell_0_0 (.BL(BL0),.BLN(BLN0),.WL(WL0));
sram_cell_6t_5 inst_cell_0_1 (.BL(BL1),.BLN(BLN1),.WL(WL0));
sram_cell_6t_5 inst_cell_0_2 (.BL(BL2),.BLN(BLN2),.WL(WL0));
sram_cell_6t_5 inst_cell_0_3 (.BL(BL3),.BLN(BLN3),.WL(WL0));
sram_cell_6t_5 inst_cell_0_4 (.BL(BL4),.BLN(BLN4),.WL(WL0));
sram_cell_6t_5 inst_cell_0_5 (.BL(BL5),.BLN(BLN5),.WL(WL0));
sram_cell_6t_5 inst_cell_0_6 (.BL(BL6),.BLN(BLN6),.WL(WL0));
sram_cell_6t_5 inst_cell_0_7 (.BL(BL7),.BLN(BLN7),.WL(WL0));
sram_cell_6t_5 inst_cell_0_8 (.BL(BL8),.BLN(BLN8),.WL(WL0));
sram_cell_6t_5 inst_cell_0_9 (.BL(BL9),.BLN(BLN9),.WL(WL0));
sram_cell_6t_5 inst_cell_0_10 (.BL(BL10),.BLN(BLN10),.WL(WL0));
sram_cell_6t_5 inst_cell_0_11 (.BL(BL11),.BLN(BLN11),.WL(WL0));
sram_cell_6t_5 inst_cell_0_12 (.BL(BL12),.BLN(BLN12),.WL(WL0));
sram_cell_6t_5 inst_cell_0_13 (.BL(BL13),.BLN(BLN13),.WL(WL0));
sram_cell_6t_5 inst_cell_0_14 (.BL(BL14),.BLN(BLN14),.WL(WL0));
sram_cell_6t_5 inst_cell_0_15 (.BL(BL15),.BLN(BLN15),.WL(WL0));
sram_cell_6t_5 inst_cell_0_16 (.BL(BL16),.BLN(BLN16),.WL(WL0));
sram_cell_6t_5 inst_cell_0_17 (.BL(BL17),.BLN(BLN17),.WL(WL0));
sram_cell_6t_5 inst_cell_0_18 (.BL(BL18),.BLN(BLN18),.WL(WL0));
sram_cell_6t_5 inst_cell_0_19 (.BL(BL19),.BLN(BLN19),.WL(WL0));
sram_cell_6t_5 inst_cell_0_20 (.BL(BL20),.BLN(BLN20),.WL(WL0));
sram_cell_6t_5 inst_cell_0_21 (.BL(BL21),.BLN(BLN21),.WL(WL0));
sram_cell_6t_5 inst_cell_0_22 (.BL(BL22),.BLN(BLN22),.WL(WL0));
sram_cell_6t_5 inst_cell_0_23 (.BL(BL23),.BLN(BLN23),.WL(WL0));
sram_cell_6t_5 inst_cell_0_24 (.BL(BL24),.BLN(BLN24),.WL(WL0));
sram_cell_6t_5 inst_cell_0_25 (.BL(BL25),.BLN(BLN25),.WL(WL0));
sram_cell_6t_5 inst_cell_0_26 (.BL(BL26),.BLN(BLN26),.WL(WL0));
sram_cell_6t_5 inst_cell_0_27 (.BL(BL27),.BLN(BLN27),.WL(WL0));
sram_cell_6t_5 inst_cell_0_28 (.BL(BL28),.BLN(BLN28),.WL(WL0));
sram_cell_6t_5 inst_cell_0_29 (.BL(BL29),.BLN(BLN29),.WL(WL0));
sram_cell_6t_5 inst_cell_0_30 (.BL(BL30),.BLN(BLN30),.WL(WL0));
sram_cell_6t_5 inst_cell_0_31 (.BL(BL31),.BLN(BLN31),.WL(WL0));
sram_cell_6t_5 inst_cell_0_32 (.BL(BL32),.BLN(BLN32),.WL(WL0));
sram_cell_6t_5 inst_cell_0_33 (.BL(BL33),.BLN(BLN33),.WL(WL0));
sram_cell_6t_5 inst_cell_0_34 (.BL(BL34),.BLN(BLN34),.WL(WL0));
sram_cell_6t_5 inst_cell_0_35 (.BL(BL35),.BLN(BLN35),.WL(WL0));
sram_cell_6t_5 inst_cell_0_36 (.BL(BL36),.BLN(BLN36),.WL(WL0));
sram_cell_6t_5 inst_cell_0_37 (.BL(BL37),.BLN(BLN37),.WL(WL0));
sram_cell_6t_5 inst_cell_0_38 (.BL(BL38),.BLN(BLN38),.WL(WL0));
sram_cell_6t_5 inst_cell_0_39 (.BL(BL39),.BLN(BLN39),.WL(WL0));
sram_cell_6t_5 inst_cell_0_40 (.BL(BL40),.BLN(BLN40),.WL(WL0));
sram_cell_6t_5 inst_cell_0_41 (.BL(BL41),.BLN(BLN41),.WL(WL0));
sram_cell_6t_5 inst_cell_0_42 (.BL(BL42),.BLN(BLN42),.WL(WL0));
sram_cell_6t_5 inst_cell_0_43 (.BL(BL43),.BLN(BLN43),.WL(WL0));
sram_cell_6t_5 inst_cell_0_44 (.BL(BL44),.BLN(BLN44),.WL(WL0));
sram_cell_6t_5 inst_cell_0_45 (.BL(BL45),.BLN(BLN45),.WL(WL0));
sram_cell_6t_5 inst_cell_0_46 (.BL(BL46),.BLN(BLN46),.WL(WL0));
sram_cell_6t_5 inst_cell_0_47 (.BL(BL47),.BLN(BLN47),.WL(WL0));
sram_cell_6t_5 inst_cell_0_48 (.BL(BL48),.BLN(BLN48),.WL(WL0));
sram_cell_6t_5 inst_cell_0_49 (.BL(BL49),.BLN(BLN49),.WL(WL0));
sram_cell_6t_5 inst_cell_0_50 (.BL(BL50),.BLN(BLN50),.WL(WL0));
sram_cell_6t_5 inst_cell_0_51 (.BL(BL51),.BLN(BLN51),.WL(WL0));
sram_cell_6t_5 inst_cell_0_52 (.BL(BL52),.BLN(BLN52),.WL(WL0));
sram_cell_6t_5 inst_cell_0_53 (.BL(BL53),.BLN(BLN53),.WL(WL0));
sram_cell_6t_5 inst_cell_0_54 (.BL(BL54),.BLN(BLN54),.WL(WL0));
sram_cell_6t_5 inst_cell_0_55 (.BL(BL55),.BLN(BLN55),.WL(WL0));
sram_cell_6t_5 inst_cell_0_56 (.BL(BL56),.BLN(BLN56),.WL(WL0));
sram_cell_6t_5 inst_cell_0_57 (.BL(BL57),.BLN(BLN57),.WL(WL0));
sram_cell_6t_5 inst_cell_0_58 (.BL(BL58),.BLN(BLN58),.WL(WL0));
sram_cell_6t_5 inst_cell_0_59 (.BL(BL59),.BLN(BLN59),.WL(WL0));
sram_cell_6t_5 inst_cell_0_60 (.BL(BL60),.BLN(BLN60),.WL(WL0));
sram_cell_6t_5 inst_cell_0_61 (.BL(BL61),.BLN(BLN61),.WL(WL0));
sram_cell_6t_5 inst_cell_0_62 (.BL(BL62),.BLN(BLN62),.WL(WL0));
sram_cell_6t_5 inst_cell_0_63 (.BL(BL63),.BLN(BLN63),.WL(WL0));
sram_cell_6t_5 inst_cell_0_64 (.BL(BL64),.BLN(BLN64),.WL(WL0));
sram_cell_6t_5 inst_cell_0_65 (.BL(BL65),.BLN(BLN65),.WL(WL0));
sram_cell_6t_5 inst_cell_0_66 (.BL(BL66),.BLN(BLN66),.WL(WL0));
sram_cell_6t_5 inst_cell_0_67 (.BL(BL67),.BLN(BLN67),.WL(WL0));
sram_cell_6t_5 inst_cell_0_68 (.BL(BL68),.BLN(BLN68),.WL(WL0));
sram_cell_6t_5 inst_cell_0_69 (.BL(BL69),.BLN(BLN69),.WL(WL0));
sram_cell_6t_5 inst_cell_0_70 (.BL(BL70),.BLN(BLN70),.WL(WL0));
sram_cell_6t_5 inst_cell_0_71 (.BL(BL71),.BLN(BLN71),.WL(WL0));
sram_cell_6t_5 inst_cell_0_72 (.BL(BL72),.BLN(BLN72),.WL(WL0));
sram_cell_6t_5 inst_cell_0_73 (.BL(BL73),.BLN(BLN73),.WL(WL0));
sram_cell_6t_5 inst_cell_0_74 (.BL(BL74),.BLN(BLN74),.WL(WL0));
sram_cell_6t_5 inst_cell_0_75 (.BL(BL75),.BLN(BLN75),.WL(WL0));
sram_cell_6t_5 inst_cell_0_76 (.BL(BL76),.BLN(BLN76),.WL(WL0));
sram_cell_6t_5 inst_cell_0_77 (.BL(BL77),.BLN(BLN77),.WL(WL0));
sram_cell_6t_5 inst_cell_0_78 (.BL(BL78),.BLN(BLN78),.WL(WL0));
sram_cell_6t_5 inst_cell_0_79 (.BL(BL79),.BLN(BLN79),.WL(WL0));
sram_cell_6t_5 inst_cell_0_80 (.BL(BL80),.BLN(BLN80),.WL(WL0));
sram_cell_6t_5 inst_cell_0_81 (.BL(BL81),.BLN(BLN81),.WL(WL0));
sram_cell_6t_5 inst_cell_0_82 (.BL(BL82),.BLN(BLN82),.WL(WL0));
sram_cell_6t_5 inst_cell_0_83 (.BL(BL83),.BLN(BLN83),.WL(WL0));
sram_cell_6t_5 inst_cell_0_84 (.BL(BL84),.BLN(BLN84),.WL(WL0));
sram_cell_6t_5 inst_cell_0_85 (.BL(BL85),.BLN(BLN85),.WL(WL0));
sram_cell_6t_5 inst_cell_0_86 (.BL(BL86),.BLN(BLN86),.WL(WL0));
sram_cell_6t_5 inst_cell_0_87 (.BL(BL87),.BLN(BLN87),.WL(WL0));
sram_cell_6t_5 inst_cell_0_88 (.BL(BL88),.BLN(BLN88),.WL(WL0));
sram_cell_6t_5 inst_cell_0_89 (.BL(BL89),.BLN(BLN89),.WL(WL0));
sram_cell_6t_5 inst_cell_0_90 (.BL(BL90),.BLN(BLN90),.WL(WL0));
sram_cell_6t_5 inst_cell_0_91 (.BL(BL91),.BLN(BLN91),.WL(WL0));
sram_cell_6t_5 inst_cell_0_92 (.BL(BL92),.BLN(BLN92),.WL(WL0));
sram_cell_6t_5 inst_cell_0_93 (.BL(BL93),.BLN(BLN93),.WL(WL0));
sram_cell_6t_5 inst_cell_0_94 (.BL(BL94),.BLN(BLN94),.WL(WL0));
sram_cell_6t_5 inst_cell_0_95 (.BL(BL95),.BLN(BLN95),.WL(WL0));
sram_cell_6t_5 inst_cell_0_96 (.BL(BL96),.BLN(BLN96),.WL(WL0));
sram_cell_6t_5 inst_cell_0_97 (.BL(BL97),.BLN(BLN97),.WL(WL0));
sram_cell_6t_5 inst_cell_0_98 (.BL(BL98),.BLN(BLN98),.WL(WL0));
sram_cell_6t_5 inst_cell_0_99 (.BL(BL99),.BLN(BLN99),.WL(WL0));
sram_cell_6t_5 inst_cell_0_100 (.BL(BL100),.BLN(BLN100),.WL(WL0));
sram_cell_6t_5 inst_cell_0_101 (.BL(BL101),.BLN(BLN101),.WL(WL0));
sram_cell_6t_5 inst_cell_0_102 (.BL(BL102),.BLN(BLN102),.WL(WL0));
sram_cell_6t_5 inst_cell_0_103 (.BL(BL103),.BLN(BLN103),.WL(WL0));
sram_cell_6t_5 inst_cell_0_104 (.BL(BL104),.BLN(BLN104),.WL(WL0));
sram_cell_6t_5 inst_cell_0_105 (.BL(BL105),.BLN(BLN105),.WL(WL0));
sram_cell_6t_5 inst_cell_0_106 (.BL(BL106),.BLN(BLN106),.WL(WL0));
sram_cell_6t_5 inst_cell_0_107 (.BL(BL107),.BLN(BLN107),.WL(WL0));
sram_cell_6t_5 inst_cell_0_108 (.BL(BL108),.BLN(BLN108),.WL(WL0));
sram_cell_6t_5 inst_cell_0_109 (.BL(BL109),.BLN(BLN109),.WL(WL0));
sram_cell_6t_5 inst_cell_0_110 (.BL(BL110),.BLN(BLN110),.WL(WL0));
sram_cell_6t_5 inst_cell_0_111 (.BL(BL111),.BLN(BLN111),.WL(WL0));
sram_cell_6t_5 inst_cell_0_112 (.BL(BL112),.BLN(BLN112),.WL(WL0));
sram_cell_6t_5 inst_cell_0_113 (.BL(BL113),.BLN(BLN113),.WL(WL0));
sram_cell_6t_5 inst_cell_0_114 (.BL(BL114),.BLN(BLN114),.WL(WL0));
sram_cell_6t_5 inst_cell_0_115 (.BL(BL115),.BLN(BLN115),.WL(WL0));
sram_cell_6t_5 inst_cell_0_116 (.BL(BL116),.BLN(BLN116),.WL(WL0));
sram_cell_6t_5 inst_cell_0_117 (.BL(BL117),.BLN(BLN117),.WL(WL0));
sram_cell_6t_5 inst_cell_0_118 (.BL(BL118),.BLN(BLN118),.WL(WL0));
sram_cell_6t_5 inst_cell_0_119 (.BL(BL119),.BLN(BLN119),.WL(WL0));
sram_cell_6t_5 inst_cell_0_120 (.BL(BL120),.BLN(BLN120),.WL(WL0));
sram_cell_6t_5 inst_cell_0_121 (.BL(BL121),.BLN(BLN121),.WL(WL0));
sram_cell_6t_5 inst_cell_0_122 (.BL(BL122),.BLN(BLN122),.WL(WL0));
sram_cell_6t_5 inst_cell_0_123 (.BL(BL123),.BLN(BLN123),.WL(WL0));
sram_cell_6t_5 inst_cell_0_124 (.BL(BL124),.BLN(BLN124),.WL(WL0));
sram_cell_6t_5 inst_cell_0_125 (.BL(BL125),.BLN(BLN125),.WL(WL0));
sram_cell_6t_5 inst_cell_0_126 (.BL(BL126),.BLN(BLN126),.WL(WL0));
sram_cell_6t_5 inst_cell_0_127 (.BL(BL127),.BLN(BLN127),.WL(WL0));
sram_cell_6t_5 inst_cell_1_0 (.BL(BL0),.BLN(BLN0),.WL(WL1));
sram_cell_6t_5 inst_cell_1_1 (.BL(BL1),.BLN(BLN1),.WL(WL1));
sram_cell_6t_5 inst_cell_1_2 (.BL(BL2),.BLN(BLN2),.WL(WL1));
sram_cell_6t_5 inst_cell_1_3 (.BL(BL3),.BLN(BLN3),.WL(WL1));
sram_cell_6t_5 inst_cell_1_4 (.BL(BL4),.BLN(BLN4),.WL(WL1));
sram_cell_6t_5 inst_cell_1_5 (.BL(BL5),.BLN(BLN5),.WL(WL1));
sram_cell_6t_5 inst_cell_1_6 (.BL(BL6),.BLN(BLN6),.WL(WL1));
sram_cell_6t_5 inst_cell_1_7 (.BL(BL7),.BLN(BLN7),.WL(WL1));
sram_cell_6t_5 inst_cell_1_8 (.BL(BL8),.BLN(BLN8),.WL(WL1));
sram_cell_6t_5 inst_cell_1_9 (.BL(BL9),.BLN(BLN9),.WL(WL1));
sram_cell_6t_5 inst_cell_1_10 (.BL(BL10),.BLN(BLN10),.WL(WL1));
sram_cell_6t_5 inst_cell_1_11 (.BL(BL11),.BLN(BLN11),.WL(WL1));
sram_cell_6t_5 inst_cell_1_12 (.BL(BL12),.BLN(BLN12),.WL(WL1));
sram_cell_6t_5 inst_cell_1_13 (.BL(BL13),.BLN(BLN13),.WL(WL1));
sram_cell_6t_5 inst_cell_1_14 (.BL(BL14),.BLN(BLN14),.WL(WL1));
sram_cell_6t_5 inst_cell_1_15 (.BL(BL15),.BLN(BLN15),.WL(WL1));
sram_cell_6t_5 inst_cell_1_16 (.BL(BL16),.BLN(BLN16),.WL(WL1));
sram_cell_6t_5 inst_cell_1_17 (.BL(BL17),.BLN(BLN17),.WL(WL1));
sram_cell_6t_5 inst_cell_1_18 (.BL(BL18),.BLN(BLN18),.WL(WL1));
sram_cell_6t_5 inst_cell_1_19 (.BL(BL19),.BLN(BLN19),.WL(WL1));
sram_cell_6t_5 inst_cell_1_20 (.BL(BL20),.BLN(BLN20),.WL(WL1));
sram_cell_6t_5 inst_cell_1_21 (.BL(BL21),.BLN(BLN21),.WL(WL1));
sram_cell_6t_5 inst_cell_1_22 (.BL(BL22),.BLN(BLN22),.WL(WL1));
sram_cell_6t_5 inst_cell_1_23 (.BL(BL23),.BLN(BLN23),.WL(WL1));
sram_cell_6t_5 inst_cell_1_24 (.BL(BL24),.BLN(BLN24),.WL(WL1));
sram_cell_6t_5 inst_cell_1_25 (.BL(BL25),.BLN(BLN25),.WL(WL1));
sram_cell_6t_5 inst_cell_1_26 (.BL(BL26),.BLN(BLN26),.WL(WL1));
sram_cell_6t_5 inst_cell_1_27 (.BL(BL27),.BLN(BLN27),.WL(WL1));
sram_cell_6t_5 inst_cell_1_28 (.BL(BL28),.BLN(BLN28),.WL(WL1));
sram_cell_6t_5 inst_cell_1_29 (.BL(BL29),.BLN(BLN29),.WL(WL1));
sram_cell_6t_5 inst_cell_1_30 (.BL(BL30),.BLN(BLN30),.WL(WL1));
sram_cell_6t_5 inst_cell_1_31 (.BL(BL31),.BLN(BLN31),.WL(WL1));
sram_cell_6t_5 inst_cell_1_32 (.BL(BL32),.BLN(BLN32),.WL(WL1));
sram_cell_6t_5 inst_cell_1_33 (.BL(BL33),.BLN(BLN33),.WL(WL1));
sram_cell_6t_5 inst_cell_1_34 (.BL(BL34),.BLN(BLN34),.WL(WL1));
sram_cell_6t_5 inst_cell_1_35 (.BL(BL35),.BLN(BLN35),.WL(WL1));
sram_cell_6t_5 inst_cell_1_36 (.BL(BL36),.BLN(BLN36),.WL(WL1));
sram_cell_6t_5 inst_cell_1_37 (.BL(BL37),.BLN(BLN37),.WL(WL1));
sram_cell_6t_5 inst_cell_1_38 (.BL(BL38),.BLN(BLN38),.WL(WL1));
sram_cell_6t_5 inst_cell_1_39 (.BL(BL39),.BLN(BLN39),.WL(WL1));
sram_cell_6t_5 inst_cell_1_40 (.BL(BL40),.BLN(BLN40),.WL(WL1));
sram_cell_6t_5 inst_cell_1_41 (.BL(BL41),.BLN(BLN41),.WL(WL1));
sram_cell_6t_5 inst_cell_1_42 (.BL(BL42),.BLN(BLN42),.WL(WL1));
sram_cell_6t_5 inst_cell_1_43 (.BL(BL43),.BLN(BLN43),.WL(WL1));
sram_cell_6t_5 inst_cell_1_44 (.BL(BL44),.BLN(BLN44),.WL(WL1));
sram_cell_6t_5 inst_cell_1_45 (.BL(BL45),.BLN(BLN45),.WL(WL1));
sram_cell_6t_5 inst_cell_1_46 (.BL(BL46),.BLN(BLN46),.WL(WL1));
sram_cell_6t_5 inst_cell_1_47 (.BL(BL47),.BLN(BLN47),.WL(WL1));
sram_cell_6t_5 inst_cell_1_48 (.BL(BL48),.BLN(BLN48),.WL(WL1));
sram_cell_6t_5 inst_cell_1_49 (.BL(BL49),.BLN(BLN49),.WL(WL1));
sram_cell_6t_5 inst_cell_1_50 (.BL(BL50),.BLN(BLN50),.WL(WL1));
sram_cell_6t_5 inst_cell_1_51 (.BL(BL51),.BLN(BLN51),.WL(WL1));
sram_cell_6t_5 inst_cell_1_52 (.BL(BL52),.BLN(BLN52),.WL(WL1));
sram_cell_6t_5 inst_cell_1_53 (.BL(BL53),.BLN(BLN53),.WL(WL1));
sram_cell_6t_5 inst_cell_1_54 (.BL(BL54),.BLN(BLN54),.WL(WL1));
sram_cell_6t_5 inst_cell_1_55 (.BL(BL55),.BLN(BLN55),.WL(WL1));
sram_cell_6t_5 inst_cell_1_56 (.BL(BL56),.BLN(BLN56),.WL(WL1));
sram_cell_6t_5 inst_cell_1_57 (.BL(BL57),.BLN(BLN57),.WL(WL1));
sram_cell_6t_5 inst_cell_1_58 (.BL(BL58),.BLN(BLN58),.WL(WL1));
sram_cell_6t_5 inst_cell_1_59 (.BL(BL59),.BLN(BLN59),.WL(WL1));
sram_cell_6t_5 inst_cell_1_60 (.BL(BL60),.BLN(BLN60),.WL(WL1));
sram_cell_6t_5 inst_cell_1_61 (.BL(BL61),.BLN(BLN61),.WL(WL1));
sram_cell_6t_5 inst_cell_1_62 (.BL(BL62),.BLN(BLN62),.WL(WL1));
sram_cell_6t_5 inst_cell_1_63 (.BL(BL63),.BLN(BLN63),.WL(WL1));
sram_cell_6t_5 inst_cell_1_64 (.BL(BL64),.BLN(BLN64),.WL(WL1));
sram_cell_6t_5 inst_cell_1_65 (.BL(BL65),.BLN(BLN65),.WL(WL1));
sram_cell_6t_5 inst_cell_1_66 (.BL(BL66),.BLN(BLN66),.WL(WL1));
sram_cell_6t_5 inst_cell_1_67 (.BL(BL67),.BLN(BLN67),.WL(WL1));
sram_cell_6t_5 inst_cell_1_68 (.BL(BL68),.BLN(BLN68),.WL(WL1));
sram_cell_6t_5 inst_cell_1_69 (.BL(BL69),.BLN(BLN69),.WL(WL1));
sram_cell_6t_5 inst_cell_1_70 (.BL(BL70),.BLN(BLN70),.WL(WL1));
sram_cell_6t_5 inst_cell_1_71 (.BL(BL71),.BLN(BLN71),.WL(WL1));
sram_cell_6t_5 inst_cell_1_72 (.BL(BL72),.BLN(BLN72),.WL(WL1));
sram_cell_6t_5 inst_cell_1_73 (.BL(BL73),.BLN(BLN73),.WL(WL1));
sram_cell_6t_5 inst_cell_1_74 (.BL(BL74),.BLN(BLN74),.WL(WL1));
sram_cell_6t_5 inst_cell_1_75 (.BL(BL75),.BLN(BLN75),.WL(WL1));
sram_cell_6t_5 inst_cell_1_76 (.BL(BL76),.BLN(BLN76),.WL(WL1));
sram_cell_6t_5 inst_cell_1_77 (.BL(BL77),.BLN(BLN77),.WL(WL1));
sram_cell_6t_5 inst_cell_1_78 (.BL(BL78),.BLN(BLN78),.WL(WL1));
sram_cell_6t_5 inst_cell_1_79 (.BL(BL79),.BLN(BLN79),.WL(WL1));
sram_cell_6t_5 inst_cell_1_80 (.BL(BL80),.BLN(BLN80),.WL(WL1));
sram_cell_6t_5 inst_cell_1_81 (.BL(BL81),.BLN(BLN81),.WL(WL1));
sram_cell_6t_5 inst_cell_1_82 (.BL(BL82),.BLN(BLN82),.WL(WL1));
sram_cell_6t_5 inst_cell_1_83 (.BL(BL83),.BLN(BLN83),.WL(WL1));
sram_cell_6t_5 inst_cell_1_84 (.BL(BL84),.BLN(BLN84),.WL(WL1));
sram_cell_6t_5 inst_cell_1_85 (.BL(BL85),.BLN(BLN85),.WL(WL1));
sram_cell_6t_5 inst_cell_1_86 (.BL(BL86),.BLN(BLN86),.WL(WL1));
sram_cell_6t_5 inst_cell_1_87 (.BL(BL87),.BLN(BLN87),.WL(WL1));
sram_cell_6t_5 inst_cell_1_88 (.BL(BL88),.BLN(BLN88),.WL(WL1));
sram_cell_6t_5 inst_cell_1_89 (.BL(BL89),.BLN(BLN89),.WL(WL1));
sram_cell_6t_5 inst_cell_1_90 (.BL(BL90),.BLN(BLN90),.WL(WL1));
sram_cell_6t_5 inst_cell_1_91 (.BL(BL91),.BLN(BLN91),.WL(WL1));
sram_cell_6t_5 inst_cell_1_92 (.BL(BL92),.BLN(BLN92),.WL(WL1));
sram_cell_6t_5 inst_cell_1_93 (.BL(BL93),.BLN(BLN93),.WL(WL1));
sram_cell_6t_5 inst_cell_1_94 (.BL(BL94),.BLN(BLN94),.WL(WL1));
sram_cell_6t_5 inst_cell_1_95 (.BL(BL95),.BLN(BLN95),.WL(WL1));
sram_cell_6t_5 inst_cell_1_96 (.BL(BL96),.BLN(BLN96),.WL(WL1));
sram_cell_6t_5 inst_cell_1_97 (.BL(BL97),.BLN(BLN97),.WL(WL1));
sram_cell_6t_5 inst_cell_1_98 (.BL(BL98),.BLN(BLN98),.WL(WL1));
sram_cell_6t_5 inst_cell_1_99 (.BL(BL99),.BLN(BLN99),.WL(WL1));
sram_cell_6t_5 inst_cell_1_100 (.BL(BL100),.BLN(BLN100),.WL(WL1));
sram_cell_6t_5 inst_cell_1_101 (.BL(BL101),.BLN(BLN101),.WL(WL1));
sram_cell_6t_5 inst_cell_1_102 (.BL(BL102),.BLN(BLN102),.WL(WL1));
sram_cell_6t_5 inst_cell_1_103 (.BL(BL103),.BLN(BLN103),.WL(WL1));
sram_cell_6t_5 inst_cell_1_104 (.BL(BL104),.BLN(BLN104),.WL(WL1));
sram_cell_6t_5 inst_cell_1_105 (.BL(BL105),.BLN(BLN105),.WL(WL1));
sram_cell_6t_5 inst_cell_1_106 (.BL(BL106),.BLN(BLN106),.WL(WL1));
sram_cell_6t_5 inst_cell_1_107 (.BL(BL107),.BLN(BLN107),.WL(WL1));
sram_cell_6t_5 inst_cell_1_108 (.BL(BL108),.BLN(BLN108),.WL(WL1));
sram_cell_6t_5 inst_cell_1_109 (.BL(BL109),.BLN(BLN109),.WL(WL1));
sram_cell_6t_5 inst_cell_1_110 (.BL(BL110),.BLN(BLN110),.WL(WL1));
sram_cell_6t_5 inst_cell_1_111 (.BL(BL111),.BLN(BLN111),.WL(WL1));
sram_cell_6t_5 inst_cell_1_112 (.BL(BL112),.BLN(BLN112),.WL(WL1));
sram_cell_6t_5 inst_cell_1_113 (.BL(BL113),.BLN(BLN113),.WL(WL1));
sram_cell_6t_5 inst_cell_1_114 (.BL(BL114),.BLN(BLN114),.WL(WL1));
sram_cell_6t_5 inst_cell_1_115 (.BL(BL115),.BLN(BLN115),.WL(WL1));
sram_cell_6t_5 inst_cell_1_116 (.BL(BL116),.BLN(BLN116),.WL(WL1));
sram_cell_6t_5 inst_cell_1_117 (.BL(BL117),.BLN(BLN117),.WL(WL1));
sram_cell_6t_5 inst_cell_1_118 (.BL(BL118),.BLN(BLN118),.WL(WL1));
sram_cell_6t_5 inst_cell_1_119 (.BL(BL119),.BLN(BLN119),.WL(WL1));
sram_cell_6t_5 inst_cell_1_120 (.BL(BL120),.BLN(BLN120),.WL(WL1));
sram_cell_6t_5 inst_cell_1_121 (.BL(BL121),.BLN(BLN121),.WL(WL1));
sram_cell_6t_5 inst_cell_1_122 (.BL(BL122),.BLN(BLN122),.WL(WL1));
sram_cell_6t_5 inst_cell_1_123 (.BL(BL123),.BLN(BLN123),.WL(WL1));
sram_cell_6t_5 inst_cell_1_124 (.BL(BL124),.BLN(BLN124),.WL(WL1));
sram_cell_6t_5 inst_cell_1_125 (.BL(BL125),.BLN(BLN125),.WL(WL1));
sram_cell_6t_5 inst_cell_1_126 (.BL(BL126),.BLN(BLN126),.WL(WL1));
sram_cell_6t_5 inst_cell_1_127 (.BL(BL127),.BLN(BLN127),.WL(WL1));
sram_cell_6t_5 inst_cell_2_0 (.BL(BL0),.BLN(BLN0),.WL(WL2));
sram_cell_6t_5 inst_cell_2_1 (.BL(BL1),.BLN(BLN1),.WL(WL2));
sram_cell_6t_5 inst_cell_2_2 (.BL(BL2),.BLN(BLN2),.WL(WL2));
sram_cell_6t_5 inst_cell_2_3 (.BL(BL3),.BLN(BLN3),.WL(WL2));
sram_cell_6t_5 inst_cell_2_4 (.BL(BL4),.BLN(BLN4),.WL(WL2));
sram_cell_6t_5 inst_cell_2_5 (.BL(BL5),.BLN(BLN5),.WL(WL2));
sram_cell_6t_5 inst_cell_2_6 (.BL(BL6),.BLN(BLN6),.WL(WL2));
sram_cell_6t_5 inst_cell_2_7 (.BL(BL7),.BLN(BLN7),.WL(WL2));
sram_cell_6t_5 inst_cell_2_8 (.BL(BL8),.BLN(BLN8),.WL(WL2));
sram_cell_6t_5 inst_cell_2_9 (.BL(BL9),.BLN(BLN9),.WL(WL2));
sram_cell_6t_5 inst_cell_2_10 (.BL(BL10),.BLN(BLN10),.WL(WL2));
sram_cell_6t_5 inst_cell_2_11 (.BL(BL11),.BLN(BLN11),.WL(WL2));
sram_cell_6t_5 inst_cell_2_12 (.BL(BL12),.BLN(BLN12),.WL(WL2));
sram_cell_6t_5 inst_cell_2_13 (.BL(BL13),.BLN(BLN13),.WL(WL2));
sram_cell_6t_5 inst_cell_2_14 (.BL(BL14),.BLN(BLN14),.WL(WL2));
sram_cell_6t_5 inst_cell_2_15 (.BL(BL15),.BLN(BLN15),.WL(WL2));
sram_cell_6t_5 inst_cell_2_16 (.BL(BL16),.BLN(BLN16),.WL(WL2));
sram_cell_6t_5 inst_cell_2_17 (.BL(BL17),.BLN(BLN17),.WL(WL2));
sram_cell_6t_5 inst_cell_2_18 (.BL(BL18),.BLN(BLN18),.WL(WL2));
sram_cell_6t_5 inst_cell_2_19 (.BL(BL19),.BLN(BLN19),.WL(WL2));
sram_cell_6t_5 inst_cell_2_20 (.BL(BL20),.BLN(BLN20),.WL(WL2));
sram_cell_6t_5 inst_cell_2_21 (.BL(BL21),.BLN(BLN21),.WL(WL2));
sram_cell_6t_5 inst_cell_2_22 (.BL(BL22),.BLN(BLN22),.WL(WL2));
sram_cell_6t_5 inst_cell_2_23 (.BL(BL23),.BLN(BLN23),.WL(WL2));
sram_cell_6t_5 inst_cell_2_24 (.BL(BL24),.BLN(BLN24),.WL(WL2));
sram_cell_6t_5 inst_cell_2_25 (.BL(BL25),.BLN(BLN25),.WL(WL2));
sram_cell_6t_5 inst_cell_2_26 (.BL(BL26),.BLN(BLN26),.WL(WL2));
sram_cell_6t_5 inst_cell_2_27 (.BL(BL27),.BLN(BLN27),.WL(WL2));
sram_cell_6t_5 inst_cell_2_28 (.BL(BL28),.BLN(BLN28),.WL(WL2));
sram_cell_6t_5 inst_cell_2_29 (.BL(BL29),.BLN(BLN29),.WL(WL2));
sram_cell_6t_5 inst_cell_2_30 (.BL(BL30),.BLN(BLN30),.WL(WL2));
sram_cell_6t_5 inst_cell_2_31 (.BL(BL31),.BLN(BLN31),.WL(WL2));
sram_cell_6t_5 inst_cell_2_32 (.BL(BL32),.BLN(BLN32),.WL(WL2));
sram_cell_6t_5 inst_cell_2_33 (.BL(BL33),.BLN(BLN33),.WL(WL2));
sram_cell_6t_5 inst_cell_2_34 (.BL(BL34),.BLN(BLN34),.WL(WL2));
sram_cell_6t_5 inst_cell_2_35 (.BL(BL35),.BLN(BLN35),.WL(WL2));
sram_cell_6t_5 inst_cell_2_36 (.BL(BL36),.BLN(BLN36),.WL(WL2));
sram_cell_6t_5 inst_cell_2_37 (.BL(BL37),.BLN(BLN37),.WL(WL2));
sram_cell_6t_5 inst_cell_2_38 (.BL(BL38),.BLN(BLN38),.WL(WL2));
sram_cell_6t_5 inst_cell_2_39 (.BL(BL39),.BLN(BLN39),.WL(WL2));
sram_cell_6t_5 inst_cell_2_40 (.BL(BL40),.BLN(BLN40),.WL(WL2));
sram_cell_6t_5 inst_cell_2_41 (.BL(BL41),.BLN(BLN41),.WL(WL2));
sram_cell_6t_5 inst_cell_2_42 (.BL(BL42),.BLN(BLN42),.WL(WL2));
sram_cell_6t_5 inst_cell_2_43 (.BL(BL43),.BLN(BLN43),.WL(WL2));
sram_cell_6t_5 inst_cell_2_44 (.BL(BL44),.BLN(BLN44),.WL(WL2));
sram_cell_6t_5 inst_cell_2_45 (.BL(BL45),.BLN(BLN45),.WL(WL2));
sram_cell_6t_5 inst_cell_2_46 (.BL(BL46),.BLN(BLN46),.WL(WL2));
sram_cell_6t_5 inst_cell_2_47 (.BL(BL47),.BLN(BLN47),.WL(WL2));
sram_cell_6t_5 inst_cell_2_48 (.BL(BL48),.BLN(BLN48),.WL(WL2));
sram_cell_6t_5 inst_cell_2_49 (.BL(BL49),.BLN(BLN49),.WL(WL2));
sram_cell_6t_5 inst_cell_2_50 (.BL(BL50),.BLN(BLN50),.WL(WL2));
sram_cell_6t_5 inst_cell_2_51 (.BL(BL51),.BLN(BLN51),.WL(WL2));
sram_cell_6t_5 inst_cell_2_52 (.BL(BL52),.BLN(BLN52),.WL(WL2));
sram_cell_6t_5 inst_cell_2_53 (.BL(BL53),.BLN(BLN53),.WL(WL2));
sram_cell_6t_5 inst_cell_2_54 (.BL(BL54),.BLN(BLN54),.WL(WL2));
sram_cell_6t_5 inst_cell_2_55 (.BL(BL55),.BLN(BLN55),.WL(WL2));
sram_cell_6t_5 inst_cell_2_56 (.BL(BL56),.BLN(BLN56),.WL(WL2));
sram_cell_6t_5 inst_cell_2_57 (.BL(BL57),.BLN(BLN57),.WL(WL2));
sram_cell_6t_5 inst_cell_2_58 (.BL(BL58),.BLN(BLN58),.WL(WL2));
sram_cell_6t_5 inst_cell_2_59 (.BL(BL59),.BLN(BLN59),.WL(WL2));
sram_cell_6t_5 inst_cell_2_60 (.BL(BL60),.BLN(BLN60),.WL(WL2));
sram_cell_6t_5 inst_cell_2_61 (.BL(BL61),.BLN(BLN61),.WL(WL2));
sram_cell_6t_5 inst_cell_2_62 (.BL(BL62),.BLN(BLN62),.WL(WL2));
sram_cell_6t_5 inst_cell_2_63 (.BL(BL63),.BLN(BLN63),.WL(WL2));
sram_cell_6t_5 inst_cell_2_64 (.BL(BL64),.BLN(BLN64),.WL(WL2));
sram_cell_6t_5 inst_cell_2_65 (.BL(BL65),.BLN(BLN65),.WL(WL2));
sram_cell_6t_5 inst_cell_2_66 (.BL(BL66),.BLN(BLN66),.WL(WL2));
sram_cell_6t_5 inst_cell_2_67 (.BL(BL67),.BLN(BLN67),.WL(WL2));
sram_cell_6t_5 inst_cell_2_68 (.BL(BL68),.BLN(BLN68),.WL(WL2));
sram_cell_6t_5 inst_cell_2_69 (.BL(BL69),.BLN(BLN69),.WL(WL2));
sram_cell_6t_5 inst_cell_2_70 (.BL(BL70),.BLN(BLN70),.WL(WL2));
sram_cell_6t_5 inst_cell_2_71 (.BL(BL71),.BLN(BLN71),.WL(WL2));
sram_cell_6t_5 inst_cell_2_72 (.BL(BL72),.BLN(BLN72),.WL(WL2));
sram_cell_6t_5 inst_cell_2_73 (.BL(BL73),.BLN(BLN73),.WL(WL2));
sram_cell_6t_5 inst_cell_2_74 (.BL(BL74),.BLN(BLN74),.WL(WL2));
sram_cell_6t_5 inst_cell_2_75 (.BL(BL75),.BLN(BLN75),.WL(WL2));
sram_cell_6t_5 inst_cell_2_76 (.BL(BL76),.BLN(BLN76),.WL(WL2));
sram_cell_6t_5 inst_cell_2_77 (.BL(BL77),.BLN(BLN77),.WL(WL2));
sram_cell_6t_5 inst_cell_2_78 (.BL(BL78),.BLN(BLN78),.WL(WL2));
sram_cell_6t_5 inst_cell_2_79 (.BL(BL79),.BLN(BLN79),.WL(WL2));
sram_cell_6t_5 inst_cell_2_80 (.BL(BL80),.BLN(BLN80),.WL(WL2));
sram_cell_6t_5 inst_cell_2_81 (.BL(BL81),.BLN(BLN81),.WL(WL2));
sram_cell_6t_5 inst_cell_2_82 (.BL(BL82),.BLN(BLN82),.WL(WL2));
sram_cell_6t_5 inst_cell_2_83 (.BL(BL83),.BLN(BLN83),.WL(WL2));
sram_cell_6t_5 inst_cell_2_84 (.BL(BL84),.BLN(BLN84),.WL(WL2));
sram_cell_6t_5 inst_cell_2_85 (.BL(BL85),.BLN(BLN85),.WL(WL2));
sram_cell_6t_5 inst_cell_2_86 (.BL(BL86),.BLN(BLN86),.WL(WL2));
sram_cell_6t_5 inst_cell_2_87 (.BL(BL87),.BLN(BLN87),.WL(WL2));
sram_cell_6t_5 inst_cell_2_88 (.BL(BL88),.BLN(BLN88),.WL(WL2));
sram_cell_6t_5 inst_cell_2_89 (.BL(BL89),.BLN(BLN89),.WL(WL2));
sram_cell_6t_5 inst_cell_2_90 (.BL(BL90),.BLN(BLN90),.WL(WL2));
sram_cell_6t_5 inst_cell_2_91 (.BL(BL91),.BLN(BLN91),.WL(WL2));
sram_cell_6t_5 inst_cell_2_92 (.BL(BL92),.BLN(BLN92),.WL(WL2));
sram_cell_6t_5 inst_cell_2_93 (.BL(BL93),.BLN(BLN93),.WL(WL2));
sram_cell_6t_5 inst_cell_2_94 (.BL(BL94),.BLN(BLN94),.WL(WL2));
sram_cell_6t_5 inst_cell_2_95 (.BL(BL95),.BLN(BLN95),.WL(WL2));
sram_cell_6t_5 inst_cell_2_96 (.BL(BL96),.BLN(BLN96),.WL(WL2));
sram_cell_6t_5 inst_cell_2_97 (.BL(BL97),.BLN(BLN97),.WL(WL2));
sram_cell_6t_5 inst_cell_2_98 (.BL(BL98),.BLN(BLN98),.WL(WL2));
sram_cell_6t_5 inst_cell_2_99 (.BL(BL99),.BLN(BLN99),.WL(WL2));
sram_cell_6t_5 inst_cell_2_100 (.BL(BL100),.BLN(BLN100),.WL(WL2));
sram_cell_6t_5 inst_cell_2_101 (.BL(BL101),.BLN(BLN101),.WL(WL2));
sram_cell_6t_5 inst_cell_2_102 (.BL(BL102),.BLN(BLN102),.WL(WL2));
sram_cell_6t_5 inst_cell_2_103 (.BL(BL103),.BLN(BLN103),.WL(WL2));
sram_cell_6t_5 inst_cell_2_104 (.BL(BL104),.BLN(BLN104),.WL(WL2));
sram_cell_6t_5 inst_cell_2_105 (.BL(BL105),.BLN(BLN105),.WL(WL2));
sram_cell_6t_5 inst_cell_2_106 (.BL(BL106),.BLN(BLN106),.WL(WL2));
sram_cell_6t_5 inst_cell_2_107 (.BL(BL107),.BLN(BLN107),.WL(WL2));
sram_cell_6t_5 inst_cell_2_108 (.BL(BL108),.BLN(BLN108),.WL(WL2));
sram_cell_6t_5 inst_cell_2_109 (.BL(BL109),.BLN(BLN109),.WL(WL2));
sram_cell_6t_5 inst_cell_2_110 (.BL(BL110),.BLN(BLN110),.WL(WL2));
sram_cell_6t_5 inst_cell_2_111 (.BL(BL111),.BLN(BLN111),.WL(WL2));
sram_cell_6t_5 inst_cell_2_112 (.BL(BL112),.BLN(BLN112),.WL(WL2));
sram_cell_6t_5 inst_cell_2_113 (.BL(BL113),.BLN(BLN113),.WL(WL2));
sram_cell_6t_5 inst_cell_2_114 (.BL(BL114),.BLN(BLN114),.WL(WL2));
sram_cell_6t_5 inst_cell_2_115 (.BL(BL115),.BLN(BLN115),.WL(WL2));
sram_cell_6t_5 inst_cell_2_116 (.BL(BL116),.BLN(BLN116),.WL(WL2));
sram_cell_6t_5 inst_cell_2_117 (.BL(BL117),.BLN(BLN117),.WL(WL2));
sram_cell_6t_5 inst_cell_2_118 (.BL(BL118),.BLN(BLN118),.WL(WL2));
sram_cell_6t_5 inst_cell_2_119 (.BL(BL119),.BLN(BLN119),.WL(WL2));
sram_cell_6t_5 inst_cell_2_120 (.BL(BL120),.BLN(BLN120),.WL(WL2));
sram_cell_6t_5 inst_cell_2_121 (.BL(BL121),.BLN(BLN121),.WL(WL2));
sram_cell_6t_5 inst_cell_2_122 (.BL(BL122),.BLN(BLN122),.WL(WL2));
sram_cell_6t_5 inst_cell_2_123 (.BL(BL123),.BLN(BLN123),.WL(WL2));
sram_cell_6t_5 inst_cell_2_124 (.BL(BL124),.BLN(BLN124),.WL(WL2));
sram_cell_6t_5 inst_cell_2_125 (.BL(BL125),.BLN(BLN125),.WL(WL2));
sram_cell_6t_5 inst_cell_2_126 (.BL(BL126),.BLN(BLN126),.WL(WL2));
sram_cell_6t_5 inst_cell_2_127 (.BL(BL127),.BLN(BLN127),.WL(WL2));
sram_cell_6t_5 inst_cell_3_0 (.BL(BL0),.BLN(BLN0),.WL(WL3));
sram_cell_6t_5 inst_cell_3_1 (.BL(BL1),.BLN(BLN1),.WL(WL3));
sram_cell_6t_5 inst_cell_3_2 (.BL(BL2),.BLN(BLN2),.WL(WL3));
sram_cell_6t_5 inst_cell_3_3 (.BL(BL3),.BLN(BLN3),.WL(WL3));
sram_cell_6t_5 inst_cell_3_4 (.BL(BL4),.BLN(BLN4),.WL(WL3));
sram_cell_6t_5 inst_cell_3_5 (.BL(BL5),.BLN(BLN5),.WL(WL3));
sram_cell_6t_5 inst_cell_3_6 (.BL(BL6),.BLN(BLN6),.WL(WL3));
sram_cell_6t_5 inst_cell_3_7 (.BL(BL7),.BLN(BLN7),.WL(WL3));
sram_cell_6t_5 inst_cell_3_8 (.BL(BL8),.BLN(BLN8),.WL(WL3));
sram_cell_6t_5 inst_cell_3_9 (.BL(BL9),.BLN(BLN9),.WL(WL3));
sram_cell_6t_5 inst_cell_3_10 (.BL(BL10),.BLN(BLN10),.WL(WL3));
sram_cell_6t_5 inst_cell_3_11 (.BL(BL11),.BLN(BLN11),.WL(WL3));
sram_cell_6t_5 inst_cell_3_12 (.BL(BL12),.BLN(BLN12),.WL(WL3));
sram_cell_6t_5 inst_cell_3_13 (.BL(BL13),.BLN(BLN13),.WL(WL3));
sram_cell_6t_5 inst_cell_3_14 (.BL(BL14),.BLN(BLN14),.WL(WL3));
sram_cell_6t_5 inst_cell_3_15 (.BL(BL15),.BLN(BLN15),.WL(WL3));
sram_cell_6t_5 inst_cell_3_16 (.BL(BL16),.BLN(BLN16),.WL(WL3));
sram_cell_6t_5 inst_cell_3_17 (.BL(BL17),.BLN(BLN17),.WL(WL3));
sram_cell_6t_5 inst_cell_3_18 (.BL(BL18),.BLN(BLN18),.WL(WL3));
sram_cell_6t_5 inst_cell_3_19 (.BL(BL19),.BLN(BLN19),.WL(WL3));
sram_cell_6t_5 inst_cell_3_20 (.BL(BL20),.BLN(BLN20),.WL(WL3));
sram_cell_6t_5 inst_cell_3_21 (.BL(BL21),.BLN(BLN21),.WL(WL3));
sram_cell_6t_5 inst_cell_3_22 (.BL(BL22),.BLN(BLN22),.WL(WL3));
sram_cell_6t_5 inst_cell_3_23 (.BL(BL23),.BLN(BLN23),.WL(WL3));
sram_cell_6t_5 inst_cell_3_24 (.BL(BL24),.BLN(BLN24),.WL(WL3));
sram_cell_6t_5 inst_cell_3_25 (.BL(BL25),.BLN(BLN25),.WL(WL3));
sram_cell_6t_5 inst_cell_3_26 (.BL(BL26),.BLN(BLN26),.WL(WL3));
sram_cell_6t_5 inst_cell_3_27 (.BL(BL27),.BLN(BLN27),.WL(WL3));
sram_cell_6t_5 inst_cell_3_28 (.BL(BL28),.BLN(BLN28),.WL(WL3));
sram_cell_6t_5 inst_cell_3_29 (.BL(BL29),.BLN(BLN29),.WL(WL3));
sram_cell_6t_5 inst_cell_3_30 (.BL(BL30),.BLN(BLN30),.WL(WL3));
sram_cell_6t_5 inst_cell_3_31 (.BL(BL31),.BLN(BLN31),.WL(WL3));
sram_cell_6t_5 inst_cell_3_32 (.BL(BL32),.BLN(BLN32),.WL(WL3));
sram_cell_6t_5 inst_cell_3_33 (.BL(BL33),.BLN(BLN33),.WL(WL3));
sram_cell_6t_5 inst_cell_3_34 (.BL(BL34),.BLN(BLN34),.WL(WL3));
sram_cell_6t_5 inst_cell_3_35 (.BL(BL35),.BLN(BLN35),.WL(WL3));
sram_cell_6t_5 inst_cell_3_36 (.BL(BL36),.BLN(BLN36),.WL(WL3));
sram_cell_6t_5 inst_cell_3_37 (.BL(BL37),.BLN(BLN37),.WL(WL3));
sram_cell_6t_5 inst_cell_3_38 (.BL(BL38),.BLN(BLN38),.WL(WL3));
sram_cell_6t_5 inst_cell_3_39 (.BL(BL39),.BLN(BLN39),.WL(WL3));
sram_cell_6t_5 inst_cell_3_40 (.BL(BL40),.BLN(BLN40),.WL(WL3));
sram_cell_6t_5 inst_cell_3_41 (.BL(BL41),.BLN(BLN41),.WL(WL3));
sram_cell_6t_5 inst_cell_3_42 (.BL(BL42),.BLN(BLN42),.WL(WL3));
sram_cell_6t_5 inst_cell_3_43 (.BL(BL43),.BLN(BLN43),.WL(WL3));
sram_cell_6t_5 inst_cell_3_44 (.BL(BL44),.BLN(BLN44),.WL(WL3));
sram_cell_6t_5 inst_cell_3_45 (.BL(BL45),.BLN(BLN45),.WL(WL3));
sram_cell_6t_5 inst_cell_3_46 (.BL(BL46),.BLN(BLN46),.WL(WL3));
sram_cell_6t_5 inst_cell_3_47 (.BL(BL47),.BLN(BLN47),.WL(WL3));
sram_cell_6t_5 inst_cell_3_48 (.BL(BL48),.BLN(BLN48),.WL(WL3));
sram_cell_6t_5 inst_cell_3_49 (.BL(BL49),.BLN(BLN49),.WL(WL3));
sram_cell_6t_5 inst_cell_3_50 (.BL(BL50),.BLN(BLN50),.WL(WL3));
sram_cell_6t_5 inst_cell_3_51 (.BL(BL51),.BLN(BLN51),.WL(WL3));
sram_cell_6t_5 inst_cell_3_52 (.BL(BL52),.BLN(BLN52),.WL(WL3));
sram_cell_6t_5 inst_cell_3_53 (.BL(BL53),.BLN(BLN53),.WL(WL3));
sram_cell_6t_5 inst_cell_3_54 (.BL(BL54),.BLN(BLN54),.WL(WL3));
sram_cell_6t_5 inst_cell_3_55 (.BL(BL55),.BLN(BLN55),.WL(WL3));
sram_cell_6t_5 inst_cell_3_56 (.BL(BL56),.BLN(BLN56),.WL(WL3));
sram_cell_6t_5 inst_cell_3_57 (.BL(BL57),.BLN(BLN57),.WL(WL3));
sram_cell_6t_5 inst_cell_3_58 (.BL(BL58),.BLN(BLN58),.WL(WL3));
sram_cell_6t_5 inst_cell_3_59 (.BL(BL59),.BLN(BLN59),.WL(WL3));
sram_cell_6t_5 inst_cell_3_60 (.BL(BL60),.BLN(BLN60),.WL(WL3));
sram_cell_6t_5 inst_cell_3_61 (.BL(BL61),.BLN(BLN61),.WL(WL3));
sram_cell_6t_5 inst_cell_3_62 (.BL(BL62),.BLN(BLN62),.WL(WL3));
sram_cell_6t_5 inst_cell_3_63 (.BL(BL63),.BLN(BLN63),.WL(WL3));
sram_cell_6t_5 inst_cell_3_64 (.BL(BL64),.BLN(BLN64),.WL(WL3));
sram_cell_6t_5 inst_cell_3_65 (.BL(BL65),.BLN(BLN65),.WL(WL3));
sram_cell_6t_5 inst_cell_3_66 (.BL(BL66),.BLN(BLN66),.WL(WL3));
sram_cell_6t_5 inst_cell_3_67 (.BL(BL67),.BLN(BLN67),.WL(WL3));
sram_cell_6t_5 inst_cell_3_68 (.BL(BL68),.BLN(BLN68),.WL(WL3));
sram_cell_6t_5 inst_cell_3_69 (.BL(BL69),.BLN(BLN69),.WL(WL3));
sram_cell_6t_5 inst_cell_3_70 (.BL(BL70),.BLN(BLN70),.WL(WL3));
sram_cell_6t_5 inst_cell_3_71 (.BL(BL71),.BLN(BLN71),.WL(WL3));
sram_cell_6t_5 inst_cell_3_72 (.BL(BL72),.BLN(BLN72),.WL(WL3));
sram_cell_6t_5 inst_cell_3_73 (.BL(BL73),.BLN(BLN73),.WL(WL3));
sram_cell_6t_5 inst_cell_3_74 (.BL(BL74),.BLN(BLN74),.WL(WL3));
sram_cell_6t_5 inst_cell_3_75 (.BL(BL75),.BLN(BLN75),.WL(WL3));
sram_cell_6t_5 inst_cell_3_76 (.BL(BL76),.BLN(BLN76),.WL(WL3));
sram_cell_6t_5 inst_cell_3_77 (.BL(BL77),.BLN(BLN77),.WL(WL3));
sram_cell_6t_5 inst_cell_3_78 (.BL(BL78),.BLN(BLN78),.WL(WL3));
sram_cell_6t_5 inst_cell_3_79 (.BL(BL79),.BLN(BLN79),.WL(WL3));
sram_cell_6t_5 inst_cell_3_80 (.BL(BL80),.BLN(BLN80),.WL(WL3));
sram_cell_6t_5 inst_cell_3_81 (.BL(BL81),.BLN(BLN81),.WL(WL3));
sram_cell_6t_5 inst_cell_3_82 (.BL(BL82),.BLN(BLN82),.WL(WL3));
sram_cell_6t_5 inst_cell_3_83 (.BL(BL83),.BLN(BLN83),.WL(WL3));
sram_cell_6t_5 inst_cell_3_84 (.BL(BL84),.BLN(BLN84),.WL(WL3));
sram_cell_6t_5 inst_cell_3_85 (.BL(BL85),.BLN(BLN85),.WL(WL3));
sram_cell_6t_5 inst_cell_3_86 (.BL(BL86),.BLN(BLN86),.WL(WL3));
sram_cell_6t_5 inst_cell_3_87 (.BL(BL87),.BLN(BLN87),.WL(WL3));
sram_cell_6t_5 inst_cell_3_88 (.BL(BL88),.BLN(BLN88),.WL(WL3));
sram_cell_6t_5 inst_cell_3_89 (.BL(BL89),.BLN(BLN89),.WL(WL3));
sram_cell_6t_5 inst_cell_3_90 (.BL(BL90),.BLN(BLN90),.WL(WL3));
sram_cell_6t_5 inst_cell_3_91 (.BL(BL91),.BLN(BLN91),.WL(WL3));
sram_cell_6t_5 inst_cell_3_92 (.BL(BL92),.BLN(BLN92),.WL(WL3));
sram_cell_6t_5 inst_cell_3_93 (.BL(BL93),.BLN(BLN93),.WL(WL3));
sram_cell_6t_5 inst_cell_3_94 (.BL(BL94),.BLN(BLN94),.WL(WL3));
sram_cell_6t_5 inst_cell_3_95 (.BL(BL95),.BLN(BLN95),.WL(WL3));
sram_cell_6t_5 inst_cell_3_96 (.BL(BL96),.BLN(BLN96),.WL(WL3));
sram_cell_6t_5 inst_cell_3_97 (.BL(BL97),.BLN(BLN97),.WL(WL3));
sram_cell_6t_5 inst_cell_3_98 (.BL(BL98),.BLN(BLN98),.WL(WL3));
sram_cell_6t_5 inst_cell_3_99 (.BL(BL99),.BLN(BLN99),.WL(WL3));
sram_cell_6t_5 inst_cell_3_100 (.BL(BL100),.BLN(BLN100),.WL(WL3));
sram_cell_6t_5 inst_cell_3_101 (.BL(BL101),.BLN(BLN101),.WL(WL3));
sram_cell_6t_5 inst_cell_3_102 (.BL(BL102),.BLN(BLN102),.WL(WL3));
sram_cell_6t_5 inst_cell_3_103 (.BL(BL103),.BLN(BLN103),.WL(WL3));
sram_cell_6t_5 inst_cell_3_104 (.BL(BL104),.BLN(BLN104),.WL(WL3));
sram_cell_6t_5 inst_cell_3_105 (.BL(BL105),.BLN(BLN105),.WL(WL3));
sram_cell_6t_5 inst_cell_3_106 (.BL(BL106),.BLN(BLN106),.WL(WL3));
sram_cell_6t_5 inst_cell_3_107 (.BL(BL107),.BLN(BLN107),.WL(WL3));
sram_cell_6t_5 inst_cell_3_108 (.BL(BL108),.BLN(BLN108),.WL(WL3));
sram_cell_6t_5 inst_cell_3_109 (.BL(BL109),.BLN(BLN109),.WL(WL3));
sram_cell_6t_5 inst_cell_3_110 (.BL(BL110),.BLN(BLN110),.WL(WL3));
sram_cell_6t_5 inst_cell_3_111 (.BL(BL111),.BLN(BLN111),.WL(WL3));
sram_cell_6t_5 inst_cell_3_112 (.BL(BL112),.BLN(BLN112),.WL(WL3));
sram_cell_6t_5 inst_cell_3_113 (.BL(BL113),.BLN(BLN113),.WL(WL3));
sram_cell_6t_5 inst_cell_3_114 (.BL(BL114),.BLN(BLN114),.WL(WL3));
sram_cell_6t_5 inst_cell_3_115 (.BL(BL115),.BLN(BLN115),.WL(WL3));
sram_cell_6t_5 inst_cell_3_116 (.BL(BL116),.BLN(BLN116),.WL(WL3));
sram_cell_6t_5 inst_cell_3_117 (.BL(BL117),.BLN(BLN117),.WL(WL3));
sram_cell_6t_5 inst_cell_3_118 (.BL(BL118),.BLN(BLN118),.WL(WL3));
sram_cell_6t_5 inst_cell_3_119 (.BL(BL119),.BLN(BLN119),.WL(WL3));
sram_cell_6t_5 inst_cell_3_120 (.BL(BL120),.BLN(BLN120),.WL(WL3));
sram_cell_6t_5 inst_cell_3_121 (.BL(BL121),.BLN(BLN121),.WL(WL3));
sram_cell_6t_5 inst_cell_3_122 (.BL(BL122),.BLN(BLN122),.WL(WL3));
sram_cell_6t_5 inst_cell_3_123 (.BL(BL123),.BLN(BLN123),.WL(WL3));
sram_cell_6t_5 inst_cell_3_124 (.BL(BL124),.BLN(BLN124),.WL(WL3));
sram_cell_6t_5 inst_cell_3_125 (.BL(BL125),.BLN(BLN125),.WL(WL3));
sram_cell_6t_5 inst_cell_3_126 (.BL(BL126),.BLN(BLN126),.WL(WL3));
sram_cell_6t_5 inst_cell_3_127 (.BL(BL127),.BLN(BLN127),.WL(WL3));
sram_cell_6t_5 inst_cell_4_0 (.BL(BL0),.BLN(BLN0),.WL(WL4));
sram_cell_6t_5 inst_cell_4_1 (.BL(BL1),.BLN(BLN1),.WL(WL4));
sram_cell_6t_5 inst_cell_4_2 (.BL(BL2),.BLN(BLN2),.WL(WL4));
sram_cell_6t_5 inst_cell_4_3 (.BL(BL3),.BLN(BLN3),.WL(WL4));
sram_cell_6t_5 inst_cell_4_4 (.BL(BL4),.BLN(BLN4),.WL(WL4));
sram_cell_6t_5 inst_cell_4_5 (.BL(BL5),.BLN(BLN5),.WL(WL4));
sram_cell_6t_5 inst_cell_4_6 (.BL(BL6),.BLN(BLN6),.WL(WL4));
sram_cell_6t_5 inst_cell_4_7 (.BL(BL7),.BLN(BLN7),.WL(WL4));
sram_cell_6t_5 inst_cell_4_8 (.BL(BL8),.BLN(BLN8),.WL(WL4));
sram_cell_6t_5 inst_cell_4_9 (.BL(BL9),.BLN(BLN9),.WL(WL4));
sram_cell_6t_5 inst_cell_4_10 (.BL(BL10),.BLN(BLN10),.WL(WL4));
sram_cell_6t_5 inst_cell_4_11 (.BL(BL11),.BLN(BLN11),.WL(WL4));
sram_cell_6t_5 inst_cell_4_12 (.BL(BL12),.BLN(BLN12),.WL(WL4));
sram_cell_6t_5 inst_cell_4_13 (.BL(BL13),.BLN(BLN13),.WL(WL4));
sram_cell_6t_5 inst_cell_4_14 (.BL(BL14),.BLN(BLN14),.WL(WL4));
sram_cell_6t_5 inst_cell_4_15 (.BL(BL15),.BLN(BLN15),.WL(WL4));
sram_cell_6t_5 inst_cell_4_16 (.BL(BL16),.BLN(BLN16),.WL(WL4));
sram_cell_6t_5 inst_cell_4_17 (.BL(BL17),.BLN(BLN17),.WL(WL4));
sram_cell_6t_5 inst_cell_4_18 (.BL(BL18),.BLN(BLN18),.WL(WL4));
sram_cell_6t_5 inst_cell_4_19 (.BL(BL19),.BLN(BLN19),.WL(WL4));
sram_cell_6t_5 inst_cell_4_20 (.BL(BL20),.BLN(BLN20),.WL(WL4));
sram_cell_6t_5 inst_cell_4_21 (.BL(BL21),.BLN(BLN21),.WL(WL4));
sram_cell_6t_5 inst_cell_4_22 (.BL(BL22),.BLN(BLN22),.WL(WL4));
sram_cell_6t_5 inst_cell_4_23 (.BL(BL23),.BLN(BLN23),.WL(WL4));
sram_cell_6t_5 inst_cell_4_24 (.BL(BL24),.BLN(BLN24),.WL(WL4));
sram_cell_6t_5 inst_cell_4_25 (.BL(BL25),.BLN(BLN25),.WL(WL4));
sram_cell_6t_5 inst_cell_4_26 (.BL(BL26),.BLN(BLN26),.WL(WL4));
sram_cell_6t_5 inst_cell_4_27 (.BL(BL27),.BLN(BLN27),.WL(WL4));
sram_cell_6t_5 inst_cell_4_28 (.BL(BL28),.BLN(BLN28),.WL(WL4));
sram_cell_6t_5 inst_cell_4_29 (.BL(BL29),.BLN(BLN29),.WL(WL4));
sram_cell_6t_5 inst_cell_4_30 (.BL(BL30),.BLN(BLN30),.WL(WL4));
sram_cell_6t_5 inst_cell_4_31 (.BL(BL31),.BLN(BLN31),.WL(WL4));
sram_cell_6t_5 inst_cell_4_32 (.BL(BL32),.BLN(BLN32),.WL(WL4));
sram_cell_6t_5 inst_cell_4_33 (.BL(BL33),.BLN(BLN33),.WL(WL4));
sram_cell_6t_5 inst_cell_4_34 (.BL(BL34),.BLN(BLN34),.WL(WL4));
sram_cell_6t_5 inst_cell_4_35 (.BL(BL35),.BLN(BLN35),.WL(WL4));
sram_cell_6t_5 inst_cell_4_36 (.BL(BL36),.BLN(BLN36),.WL(WL4));
sram_cell_6t_5 inst_cell_4_37 (.BL(BL37),.BLN(BLN37),.WL(WL4));
sram_cell_6t_5 inst_cell_4_38 (.BL(BL38),.BLN(BLN38),.WL(WL4));
sram_cell_6t_5 inst_cell_4_39 (.BL(BL39),.BLN(BLN39),.WL(WL4));
sram_cell_6t_5 inst_cell_4_40 (.BL(BL40),.BLN(BLN40),.WL(WL4));
sram_cell_6t_5 inst_cell_4_41 (.BL(BL41),.BLN(BLN41),.WL(WL4));
sram_cell_6t_5 inst_cell_4_42 (.BL(BL42),.BLN(BLN42),.WL(WL4));
sram_cell_6t_5 inst_cell_4_43 (.BL(BL43),.BLN(BLN43),.WL(WL4));
sram_cell_6t_5 inst_cell_4_44 (.BL(BL44),.BLN(BLN44),.WL(WL4));
sram_cell_6t_5 inst_cell_4_45 (.BL(BL45),.BLN(BLN45),.WL(WL4));
sram_cell_6t_5 inst_cell_4_46 (.BL(BL46),.BLN(BLN46),.WL(WL4));
sram_cell_6t_5 inst_cell_4_47 (.BL(BL47),.BLN(BLN47),.WL(WL4));
sram_cell_6t_5 inst_cell_4_48 (.BL(BL48),.BLN(BLN48),.WL(WL4));
sram_cell_6t_5 inst_cell_4_49 (.BL(BL49),.BLN(BLN49),.WL(WL4));
sram_cell_6t_5 inst_cell_4_50 (.BL(BL50),.BLN(BLN50),.WL(WL4));
sram_cell_6t_5 inst_cell_4_51 (.BL(BL51),.BLN(BLN51),.WL(WL4));
sram_cell_6t_5 inst_cell_4_52 (.BL(BL52),.BLN(BLN52),.WL(WL4));
sram_cell_6t_5 inst_cell_4_53 (.BL(BL53),.BLN(BLN53),.WL(WL4));
sram_cell_6t_5 inst_cell_4_54 (.BL(BL54),.BLN(BLN54),.WL(WL4));
sram_cell_6t_5 inst_cell_4_55 (.BL(BL55),.BLN(BLN55),.WL(WL4));
sram_cell_6t_5 inst_cell_4_56 (.BL(BL56),.BLN(BLN56),.WL(WL4));
sram_cell_6t_5 inst_cell_4_57 (.BL(BL57),.BLN(BLN57),.WL(WL4));
sram_cell_6t_5 inst_cell_4_58 (.BL(BL58),.BLN(BLN58),.WL(WL4));
sram_cell_6t_5 inst_cell_4_59 (.BL(BL59),.BLN(BLN59),.WL(WL4));
sram_cell_6t_5 inst_cell_4_60 (.BL(BL60),.BLN(BLN60),.WL(WL4));
sram_cell_6t_5 inst_cell_4_61 (.BL(BL61),.BLN(BLN61),.WL(WL4));
sram_cell_6t_5 inst_cell_4_62 (.BL(BL62),.BLN(BLN62),.WL(WL4));
sram_cell_6t_5 inst_cell_4_63 (.BL(BL63),.BLN(BLN63),.WL(WL4));
sram_cell_6t_5 inst_cell_4_64 (.BL(BL64),.BLN(BLN64),.WL(WL4));
sram_cell_6t_5 inst_cell_4_65 (.BL(BL65),.BLN(BLN65),.WL(WL4));
sram_cell_6t_5 inst_cell_4_66 (.BL(BL66),.BLN(BLN66),.WL(WL4));
sram_cell_6t_5 inst_cell_4_67 (.BL(BL67),.BLN(BLN67),.WL(WL4));
sram_cell_6t_5 inst_cell_4_68 (.BL(BL68),.BLN(BLN68),.WL(WL4));
sram_cell_6t_5 inst_cell_4_69 (.BL(BL69),.BLN(BLN69),.WL(WL4));
sram_cell_6t_5 inst_cell_4_70 (.BL(BL70),.BLN(BLN70),.WL(WL4));
sram_cell_6t_5 inst_cell_4_71 (.BL(BL71),.BLN(BLN71),.WL(WL4));
sram_cell_6t_5 inst_cell_4_72 (.BL(BL72),.BLN(BLN72),.WL(WL4));
sram_cell_6t_5 inst_cell_4_73 (.BL(BL73),.BLN(BLN73),.WL(WL4));
sram_cell_6t_5 inst_cell_4_74 (.BL(BL74),.BLN(BLN74),.WL(WL4));
sram_cell_6t_5 inst_cell_4_75 (.BL(BL75),.BLN(BLN75),.WL(WL4));
sram_cell_6t_5 inst_cell_4_76 (.BL(BL76),.BLN(BLN76),.WL(WL4));
sram_cell_6t_5 inst_cell_4_77 (.BL(BL77),.BLN(BLN77),.WL(WL4));
sram_cell_6t_5 inst_cell_4_78 (.BL(BL78),.BLN(BLN78),.WL(WL4));
sram_cell_6t_5 inst_cell_4_79 (.BL(BL79),.BLN(BLN79),.WL(WL4));
sram_cell_6t_5 inst_cell_4_80 (.BL(BL80),.BLN(BLN80),.WL(WL4));
sram_cell_6t_5 inst_cell_4_81 (.BL(BL81),.BLN(BLN81),.WL(WL4));
sram_cell_6t_5 inst_cell_4_82 (.BL(BL82),.BLN(BLN82),.WL(WL4));
sram_cell_6t_5 inst_cell_4_83 (.BL(BL83),.BLN(BLN83),.WL(WL4));
sram_cell_6t_5 inst_cell_4_84 (.BL(BL84),.BLN(BLN84),.WL(WL4));
sram_cell_6t_5 inst_cell_4_85 (.BL(BL85),.BLN(BLN85),.WL(WL4));
sram_cell_6t_5 inst_cell_4_86 (.BL(BL86),.BLN(BLN86),.WL(WL4));
sram_cell_6t_5 inst_cell_4_87 (.BL(BL87),.BLN(BLN87),.WL(WL4));
sram_cell_6t_5 inst_cell_4_88 (.BL(BL88),.BLN(BLN88),.WL(WL4));
sram_cell_6t_5 inst_cell_4_89 (.BL(BL89),.BLN(BLN89),.WL(WL4));
sram_cell_6t_5 inst_cell_4_90 (.BL(BL90),.BLN(BLN90),.WL(WL4));
sram_cell_6t_5 inst_cell_4_91 (.BL(BL91),.BLN(BLN91),.WL(WL4));
sram_cell_6t_5 inst_cell_4_92 (.BL(BL92),.BLN(BLN92),.WL(WL4));
sram_cell_6t_5 inst_cell_4_93 (.BL(BL93),.BLN(BLN93),.WL(WL4));
sram_cell_6t_5 inst_cell_4_94 (.BL(BL94),.BLN(BLN94),.WL(WL4));
sram_cell_6t_5 inst_cell_4_95 (.BL(BL95),.BLN(BLN95),.WL(WL4));
sram_cell_6t_5 inst_cell_4_96 (.BL(BL96),.BLN(BLN96),.WL(WL4));
sram_cell_6t_5 inst_cell_4_97 (.BL(BL97),.BLN(BLN97),.WL(WL4));
sram_cell_6t_5 inst_cell_4_98 (.BL(BL98),.BLN(BLN98),.WL(WL4));
sram_cell_6t_5 inst_cell_4_99 (.BL(BL99),.BLN(BLN99),.WL(WL4));
sram_cell_6t_5 inst_cell_4_100 (.BL(BL100),.BLN(BLN100),.WL(WL4));
sram_cell_6t_5 inst_cell_4_101 (.BL(BL101),.BLN(BLN101),.WL(WL4));
sram_cell_6t_5 inst_cell_4_102 (.BL(BL102),.BLN(BLN102),.WL(WL4));
sram_cell_6t_5 inst_cell_4_103 (.BL(BL103),.BLN(BLN103),.WL(WL4));
sram_cell_6t_5 inst_cell_4_104 (.BL(BL104),.BLN(BLN104),.WL(WL4));
sram_cell_6t_5 inst_cell_4_105 (.BL(BL105),.BLN(BLN105),.WL(WL4));
sram_cell_6t_5 inst_cell_4_106 (.BL(BL106),.BLN(BLN106),.WL(WL4));
sram_cell_6t_5 inst_cell_4_107 (.BL(BL107),.BLN(BLN107),.WL(WL4));
sram_cell_6t_5 inst_cell_4_108 (.BL(BL108),.BLN(BLN108),.WL(WL4));
sram_cell_6t_5 inst_cell_4_109 (.BL(BL109),.BLN(BLN109),.WL(WL4));
sram_cell_6t_5 inst_cell_4_110 (.BL(BL110),.BLN(BLN110),.WL(WL4));
sram_cell_6t_5 inst_cell_4_111 (.BL(BL111),.BLN(BLN111),.WL(WL4));
sram_cell_6t_5 inst_cell_4_112 (.BL(BL112),.BLN(BLN112),.WL(WL4));
sram_cell_6t_5 inst_cell_4_113 (.BL(BL113),.BLN(BLN113),.WL(WL4));
sram_cell_6t_5 inst_cell_4_114 (.BL(BL114),.BLN(BLN114),.WL(WL4));
sram_cell_6t_5 inst_cell_4_115 (.BL(BL115),.BLN(BLN115),.WL(WL4));
sram_cell_6t_5 inst_cell_4_116 (.BL(BL116),.BLN(BLN116),.WL(WL4));
sram_cell_6t_5 inst_cell_4_117 (.BL(BL117),.BLN(BLN117),.WL(WL4));
sram_cell_6t_5 inst_cell_4_118 (.BL(BL118),.BLN(BLN118),.WL(WL4));
sram_cell_6t_5 inst_cell_4_119 (.BL(BL119),.BLN(BLN119),.WL(WL4));
sram_cell_6t_5 inst_cell_4_120 (.BL(BL120),.BLN(BLN120),.WL(WL4));
sram_cell_6t_5 inst_cell_4_121 (.BL(BL121),.BLN(BLN121),.WL(WL4));
sram_cell_6t_5 inst_cell_4_122 (.BL(BL122),.BLN(BLN122),.WL(WL4));
sram_cell_6t_5 inst_cell_4_123 (.BL(BL123),.BLN(BLN123),.WL(WL4));
sram_cell_6t_5 inst_cell_4_124 (.BL(BL124),.BLN(BLN124),.WL(WL4));
sram_cell_6t_5 inst_cell_4_125 (.BL(BL125),.BLN(BLN125),.WL(WL4));
sram_cell_6t_5 inst_cell_4_126 (.BL(BL126),.BLN(BLN126),.WL(WL4));
sram_cell_6t_5 inst_cell_4_127 (.BL(BL127),.BLN(BLN127),.WL(WL4));
sram_cell_6t_5 inst_cell_5_0 (.BL(BL0),.BLN(BLN0),.WL(WL5));
sram_cell_6t_5 inst_cell_5_1 (.BL(BL1),.BLN(BLN1),.WL(WL5));
sram_cell_6t_5 inst_cell_5_2 (.BL(BL2),.BLN(BLN2),.WL(WL5));
sram_cell_6t_5 inst_cell_5_3 (.BL(BL3),.BLN(BLN3),.WL(WL5));
sram_cell_6t_5 inst_cell_5_4 (.BL(BL4),.BLN(BLN4),.WL(WL5));
sram_cell_6t_5 inst_cell_5_5 (.BL(BL5),.BLN(BLN5),.WL(WL5));
sram_cell_6t_5 inst_cell_5_6 (.BL(BL6),.BLN(BLN6),.WL(WL5));
sram_cell_6t_5 inst_cell_5_7 (.BL(BL7),.BLN(BLN7),.WL(WL5));
sram_cell_6t_5 inst_cell_5_8 (.BL(BL8),.BLN(BLN8),.WL(WL5));
sram_cell_6t_5 inst_cell_5_9 (.BL(BL9),.BLN(BLN9),.WL(WL5));
sram_cell_6t_5 inst_cell_5_10 (.BL(BL10),.BLN(BLN10),.WL(WL5));
sram_cell_6t_5 inst_cell_5_11 (.BL(BL11),.BLN(BLN11),.WL(WL5));
sram_cell_6t_5 inst_cell_5_12 (.BL(BL12),.BLN(BLN12),.WL(WL5));
sram_cell_6t_5 inst_cell_5_13 (.BL(BL13),.BLN(BLN13),.WL(WL5));
sram_cell_6t_5 inst_cell_5_14 (.BL(BL14),.BLN(BLN14),.WL(WL5));
sram_cell_6t_5 inst_cell_5_15 (.BL(BL15),.BLN(BLN15),.WL(WL5));
sram_cell_6t_5 inst_cell_5_16 (.BL(BL16),.BLN(BLN16),.WL(WL5));
sram_cell_6t_5 inst_cell_5_17 (.BL(BL17),.BLN(BLN17),.WL(WL5));
sram_cell_6t_5 inst_cell_5_18 (.BL(BL18),.BLN(BLN18),.WL(WL5));
sram_cell_6t_5 inst_cell_5_19 (.BL(BL19),.BLN(BLN19),.WL(WL5));
sram_cell_6t_5 inst_cell_5_20 (.BL(BL20),.BLN(BLN20),.WL(WL5));
sram_cell_6t_5 inst_cell_5_21 (.BL(BL21),.BLN(BLN21),.WL(WL5));
sram_cell_6t_5 inst_cell_5_22 (.BL(BL22),.BLN(BLN22),.WL(WL5));
sram_cell_6t_5 inst_cell_5_23 (.BL(BL23),.BLN(BLN23),.WL(WL5));
sram_cell_6t_5 inst_cell_5_24 (.BL(BL24),.BLN(BLN24),.WL(WL5));
sram_cell_6t_5 inst_cell_5_25 (.BL(BL25),.BLN(BLN25),.WL(WL5));
sram_cell_6t_5 inst_cell_5_26 (.BL(BL26),.BLN(BLN26),.WL(WL5));
sram_cell_6t_5 inst_cell_5_27 (.BL(BL27),.BLN(BLN27),.WL(WL5));
sram_cell_6t_5 inst_cell_5_28 (.BL(BL28),.BLN(BLN28),.WL(WL5));
sram_cell_6t_5 inst_cell_5_29 (.BL(BL29),.BLN(BLN29),.WL(WL5));
sram_cell_6t_5 inst_cell_5_30 (.BL(BL30),.BLN(BLN30),.WL(WL5));
sram_cell_6t_5 inst_cell_5_31 (.BL(BL31),.BLN(BLN31),.WL(WL5));
sram_cell_6t_5 inst_cell_5_32 (.BL(BL32),.BLN(BLN32),.WL(WL5));
sram_cell_6t_5 inst_cell_5_33 (.BL(BL33),.BLN(BLN33),.WL(WL5));
sram_cell_6t_5 inst_cell_5_34 (.BL(BL34),.BLN(BLN34),.WL(WL5));
sram_cell_6t_5 inst_cell_5_35 (.BL(BL35),.BLN(BLN35),.WL(WL5));
sram_cell_6t_5 inst_cell_5_36 (.BL(BL36),.BLN(BLN36),.WL(WL5));
sram_cell_6t_5 inst_cell_5_37 (.BL(BL37),.BLN(BLN37),.WL(WL5));
sram_cell_6t_5 inst_cell_5_38 (.BL(BL38),.BLN(BLN38),.WL(WL5));
sram_cell_6t_5 inst_cell_5_39 (.BL(BL39),.BLN(BLN39),.WL(WL5));
sram_cell_6t_5 inst_cell_5_40 (.BL(BL40),.BLN(BLN40),.WL(WL5));
sram_cell_6t_5 inst_cell_5_41 (.BL(BL41),.BLN(BLN41),.WL(WL5));
sram_cell_6t_5 inst_cell_5_42 (.BL(BL42),.BLN(BLN42),.WL(WL5));
sram_cell_6t_5 inst_cell_5_43 (.BL(BL43),.BLN(BLN43),.WL(WL5));
sram_cell_6t_5 inst_cell_5_44 (.BL(BL44),.BLN(BLN44),.WL(WL5));
sram_cell_6t_5 inst_cell_5_45 (.BL(BL45),.BLN(BLN45),.WL(WL5));
sram_cell_6t_5 inst_cell_5_46 (.BL(BL46),.BLN(BLN46),.WL(WL5));
sram_cell_6t_5 inst_cell_5_47 (.BL(BL47),.BLN(BLN47),.WL(WL5));
sram_cell_6t_5 inst_cell_5_48 (.BL(BL48),.BLN(BLN48),.WL(WL5));
sram_cell_6t_5 inst_cell_5_49 (.BL(BL49),.BLN(BLN49),.WL(WL5));
sram_cell_6t_5 inst_cell_5_50 (.BL(BL50),.BLN(BLN50),.WL(WL5));
sram_cell_6t_5 inst_cell_5_51 (.BL(BL51),.BLN(BLN51),.WL(WL5));
sram_cell_6t_5 inst_cell_5_52 (.BL(BL52),.BLN(BLN52),.WL(WL5));
sram_cell_6t_5 inst_cell_5_53 (.BL(BL53),.BLN(BLN53),.WL(WL5));
sram_cell_6t_5 inst_cell_5_54 (.BL(BL54),.BLN(BLN54),.WL(WL5));
sram_cell_6t_5 inst_cell_5_55 (.BL(BL55),.BLN(BLN55),.WL(WL5));
sram_cell_6t_5 inst_cell_5_56 (.BL(BL56),.BLN(BLN56),.WL(WL5));
sram_cell_6t_5 inst_cell_5_57 (.BL(BL57),.BLN(BLN57),.WL(WL5));
sram_cell_6t_5 inst_cell_5_58 (.BL(BL58),.BLN(BLN58),.WL(WL5));
sram_cell_6t_5 inst_cell_5_59 (.BL(BL59),.BLN(BLN59),.WL(WL5));
sram_cell_6t_5 inst_cell_5_60 (.BL(BL60),.BLN(BLN60),.WL(WL5));
sram_cell_6t_5 inst_cell_5_61 (.BL(BL61),.BLN(BLN61),.WL(WL5));
sram_cell_6t_5 inst_cell_5_62 (.BL(BL62),.BLN(BLN62),.WL(WL5));
sram_cell_6t_5 inst_cell_5_63 (.BL(BL63),.BLN(BLN63),.WL(WL5));
sram_cell_6t_5 inst_cell_5_64 (.BL(BL64),.BLN(BLN64),.WL(WL5));
sram_cell_6t_5 inst_cell_5_65 (.BL(BL65),.BLN(BLN65),.WL(WL5));
sram_cell_6t_5 inst_cell_5_66 (.BL(BL66),.BLN(BLN66),.WL(WL5));
sram_cell_6t_5 inst_cell_5_67 (.BL(BL67),.BLN(BLN67),.WL(WL5));
sram_cell_6t_5 inst_cell_5_68 (.BL(BL68),.BLN(BLN68),.WL(WL5));
sram_cell_6t_5 inst_cell_5_69 (.BL(BL69),.BLN(BLN69),.WL(WL5));
sram_cell_6t_5 inst_cell_5_70 (.BL(BL70),.BLN(BLN70),.WL(WL5));
sram_cell_6t_5 inst_cell_5_71 (.BL(BL71),.BLN(BLN71),.WL(WL5));
sram_cell_6t_5 inst_cell_5_72 (.BL(BL72),.BLN(BLN72),.WL(WL5));
sram_cell_6t_5 inst_cell_5_73 (.BL(BL73),.BLN(BLN73),.WL(WL5));
sram_cell_6t_5 inst_cell_5_74 (.BL(BL74),.BLN(BLN74),.WL(WL5));
sram_cell_6t_5 inst_cell_5_75 (.BL(BL75),.BLN(BLN75),.WL(WL5));
sram_cell_6t_5 inst_cell_5_76 (.BL(BL76),.BLN(BLN76),.WL(WL5));
sram_cell_6t_5 inst_cell_5_77 (.BL(BL77),.BLN(BLN77),.WL(WL5));
sram_cell_6t_5 inst_cell_5_78 (.BL(BL78),.BLN(BLN78),.WL(WL5));
sram_cell_6t_5 inst_cell_5_79 (.BL(BL79),.BLN(BLN79),.WL(WL5));
sram_cell_6t_5 inst_cell_5_80 (.BL(BL80),.BLN(BLN80),.WL(WL5));
sram_cell_6t_5 inst_cell_5_81 (.BL(BL81),.BLN(BLN81),.WL(WL5));
sram_cell_6t_5 inst_cell_5_82 (.BL(BL82),.BLN(BLN82),.WL(WL5));
sram_cell_6t_5 inst_cell_5_83 (.BL(BL83),.BLN(BLN83),.WL(WL5));
sram_cell_6t_5 inst_cell_5_84 (.BL(BL84),.BLN(BLN84),.WL(WL5));
sram_cell_6t_5 inst_cell_5_85 (.BL(BL85),.BLN(BLN85),.WL(WL5));
sram_cell_6t_5 inst_cell_5_86 (.BL(BL86),.BLN(BLN86),.WL(WL5));
sram_cell_6t_5 inst_cell_5_87 (.BL(BL87),.BLN(BLN87),.WL(WL5));
sram_cell_6t_5 inst_cell_5_88 (.BL(BL88),.BLN(BLN88),.WL(WL5));
sram_cell_6t_5 inst_cell_5_89 (.BL(BL89),.BLN(BLN89),.WL(WL5));
sram_cell_6t_5 inst_cell_5_90 (.BL(BL90),.BLN(BLN90),.WL(WL5));
sram_cell_6t_5 inst_cell_5_91 (.BL(BL91),.BLN(BLN91),.WL(WL5));
sram_cell_6t_5 inst_cell_5_92 (.BL(BL92),.BLN(BLN92),.WL(WL5));
sram_cell_6t_5 inst_cell_5_93 (.BL(BL93),.BLN(BLN93),.WL(WL5));
sram_cell_6t_5 inst_cell_5_94 (.BL(BL94),.BLN(BLN94),.WL(WL5));
sram_cell_6t_5 inst_cell_5_95 (.BL(BL95),.BLN(BLN95),.WL(WL5));
sram_cell_6t_5 inst_cell_5_96 (.BL(BL96),.BLN(BLN96),.WL(WL5));
sram_cell_6t_5 inst_cell_5_97 (.BL(BL97),.BLN(BLN97),.WL(WL5));
sram_cell_6t_5 inst_cell_5_98 (.BL(BL98),.BLN(BLN98),.WL(WL5));
sram_cell_6t_5 inst_cell_5_99 (.BL(BL99),.BLN(BLN99),.WL(WL5));
sram_cell_6t_5 inst_cell_5_100 (.BL(BL100),.BLN(BLN100),.WL(WL5));
sram_cell_6t_5 inst_cell_5_101 (.BL(BL101),.BLN(BLN101),.WL(WL5));
sram_cell_6t_5 inst_cell_5_102 (.BL(BL102),.BLN(BLN102),.WL(WL5));
sram_cell_6t_5 inst_cell_5_103 (.BL(BL103),.BLN(BLN103),.WL(WL5));
sram_cell_6t_5 inst_cell_5_104 (.BL(BL104),.BLN(BLN104),.WL(WL5));
sram_cell_6t_5 inst_cell_5_105 (.BL(BL105),.BLN(BLN105),.WL(WL5));
sram_cell_6t_5 inst_cell_5_106 (.BL(BL106),.BLN(BLN106),.WL(WL5));
sram_cell_6t_5 inst_cell_5_107 (.BL(BL107),.BLN(BLN107),.WL(WL5));
sram_cell_6t_5 inst_cell_5_108 (.BL(BL108),.BLN(BLN108),.WL(WL5));
sram_cell_6t_5 inst_cell_5_109 (.BL(BL109),.BLN(BLN109),.WL(WL5));
sram_cell_6t_5 inst_cell_5_110 (.BL(BL110),.BLN(BLN110),.WL(WL5));
sram_cell_6t_5 inst_cell_5_111 (.BL(BL111),.BLN(BLN111),.WL(WL5));
sram_cell_6t_5 inst_cell_5_112 (.BL(BL112),.BLN(BLN112),.WL(WL5));
sram_cell_6t_5 inst_cell_5_113 (.BL(BL113),.BLN(BLN113),.WL(WL5));
sram_cell_6t_5 inst_cell_5_114 (.BL(BL114),.BLN(BLN114),.WL(WL5));
sram_cell_6t_5 inst_cell_5_115 (.BL(BL115),.BLN(BLN115),.WL(WL5));
sram_cell_6t_5 inst_cell_5_116 (.BL(BL116),.BLN(BLN116),.WL(WL5));
sram_cell_6t_5 inst_cell_5_117 (.BL(BL117),.BLN(BLN117),.WL(WL5));
sram_cell_6t_5 inst_cell_5_118 (.BL(BL118),.BLN(BLN118),.WL(WL5));
sram_cell_6t_5 inst_cell_5_119 (.BL(BL119),.BLN(BLN119),.WL(WL5));
sram_cell_6t_5 inst_cell_5_120 (.BL(BL120),.BLN(BLN120),.WL(WL5));
sram_cell_6t_5 inst_cell_5_121 (.BL(BL121),.BLN(BLN121),.WL(WL5));
sram_cell_6t_5 inst_cell_5_122 (.BL(BL122),.BLN(BLN122),.WL(WL5));
sram_cell_6t_5 inst_cell_5_123 (.BL(BL123),.BLN(BLN123),.WL(WL5));
sram_cell_6t_5 inst_cell_5_124 (.BL(BL124),.BLN(BLN124),.WL(WL5));
sram_cell_6t_5 inst_cell_5_125 (.BL(BL125),.BLN(BLN125),.WL(WL5));
sram_cell_6t_5 inst_cell_5_126 (.BL(BL126),.BLN(BLN126),.WL(WL5));
sram_cell_6t_5 inst_cell_5_127 (.BL(BL127),.BLN(BLN127),.WL(WL5));
sram_cell_6t_5 inst_cell_6_0 (.BL(BL0),.BLN(BLN0),.WL(WL6));
sram_cell_6t_5 inst_cell_6_1 (.BL(BL1),.BLN(BLN1),.WL(WL6));
sram_cell_6t_5 inst_cell_6_2 (.BL(BL2),.BLN(BLN2),.WL(WL6));
sram_cell_6t_5 inst_cell_6_3 (.BL(BL3),.BLN(BLN3),.WL(WL6));
sram_cell_6t_5 inst_cell_6_4 (.BL(BL4),.BLN(BLN4),.WL(WL6));
sram_cell_6t_5 inst_cell_6_5 (.BL(BL5),.BLN(BLN5),.WL(WL6));
sram_cell_6t_5 inst_cell_6_6 (.BL(BL6),.BLN(BLN6),.WL(WL6));
sram_cell_6t_5 inst_cell_6_7 (.BL(BL7),.BLN(BLN7),.WL(WL6));
sram_cell_6t_5 inst_cell_6_8 (.BL(BL8),.BLN(BLN8),.WL(WL6));
sram_cell_6t_5 inst_cell_6_9 (.BL(BL9),.BLN(BLN9),.WL(WL6));
sram_cell_6t_5 inst_cell_6_10 (.BL(BL10),.BLN(BLN10),.WL(WL6));
sram_cell_6t_5 inst_cell_6_11 (.BL(BL11),.BLN(BLN11),.WL(WL6));
sram_cell_6t_5 inst_cell_6_12 (.BL(BL12),.BLN(BLN12),.WL(WL6));
sram_cell_6t_5 inst_cell_6_13 (.BL(BL13),.BLN(BLN13),.WL(WL6));
sram_cell_6t_5 inst_cell_6_14 (.BL(BL14),.BLN(BLN14),.WL(WL6));
sram_cell_6t_5 inst_cell_6_15 (.BL(BL15),.BLN(BLN15),.WL(WL6));
sram_cell_6t_5 inst_cell_6_16 (.BL(BL16),.BLN(BLN16),.WL(WL6));
sram_cell_6t_5 inst_cell_6_17 (.BL(BL17),.BLN(BLN17),.WL(WL6));
sram_cell_6t_5 inst_cell_6_18 (.BL(BL18),.BLN(BLN18),.WL(WL6));
sram_cell_6t_5 inst_cell_6_19 (.BL(BL19),.BLN(BLN19),.WL(WL6));
sram_cell_6t_5 inst_cell_6_20 (.BL(BL20),.BLN(BLN20),.WL(WL6));
sram_cell_6t_5 inst_cell_6_21 (.BL(BL21),.BLN(BLN21),.WL(WL6));
sram_cell_6t_5 inst_cell_6_22 (.BL(BL22),.BLN(BLN22),.WL(WL6));
sram_cell_6t_5 inst_cell_6_23 (.BL(BL23),.BLN(BLN23),.WL(WL6));
sram_cell_6t_5 inst_cell_6_24 (.BL(BL24),.BLN(BLN24),.WL(WL6));
sram_cell_6t_5 inst_cell_6_25 (.BL(BL25),.BLN(BLN25),.WL(WL6));
sram_cell_6t_5 inst_cell_6_26 (.BL(BL26),.BLN(BLN26),.WL(WL6));
sram_cell_6t_5 inst_cell_6_27 (.BL(BL27),.BLN(BLN27),.WL(WL6));
sram_cell_6t_5 inst_cell_6_28 (.BL(BL28),.BLN(BLN28),.WL(WL6));
sram_cell_6t_5 inst_cell_6_29 (.BL(BL29),.BLN(BLN29),.WL(WL6));
sram_cell_6t_5 inst_cell_6_30 (.BL(BL30),.BLN(BLN30),.WL(WL6));
sram_cell_6t_5 inst_cell_6_31 (.BL(BL31),.BLN(BLN31),.WL(WL6));
sram_cell_6t_5 inst_cell_6_32 (.BL(BL32),.BLN(BLN32),.WL(WL6));
sram_cell_6t_5 inst_cell_6_33 (.BL(BL33),.BLN(BLN33),.WL(WL6));
sram_cell_6t_5 inst_cell_6_34 (.BL(BL34),.BLN(BLN34),.WL(WL6));
sram_cell_6t_5 inst_cell_6_35 (.BL(BL35),.BLN(BLN35),.WL(WL6));
sram_cell_6t_5 inst_cell_6_36 (.BL(BL36),.BLN(BLN36),.WL(WL6));
sram_cell_6t_5 inst_cell_6_37 (.BL(BL37),.BLN(BLN37),.WL(WL6));
sram_cell_6t_5 inst_cell_6_38 (.BL(BL38),.BLN(BLN38),.WL(WL6));
sram_cell_6t_5 inst_cell_6_39 (.BL(BL39),.BLN(BLN39),.WL(WL6));
sram_cell_6t_5 inst_cell_6_40 (.BL(BL40),.BLN(BLN40),.WL(WL6));
sram_cell_6t_5 inst_cell_6_41 (.BL(BL41),.BLN(BLN41),.WL(WL6));
sram_cell_6t_5 inst_cell_6_42 (.BL(BL42),.BLN(BLN42),.WL(WL6));
sram_cell_6t_5 inst_cell_6_43 (.BL(BL43),.BLN(BLN43),.WL(WL6));
sram_cell_6t_5 inst_cell_6_44 (.BL(BL44),.BLN(BLN44),.WL(WL6));
sram_cell_6t_5 inst_cell_6_45 (.BL(BL45),.BLN(BLN45),.WL(WL6));
sram_cell_6t_5 inst_cell_6_46 (.BL(BL46),.BLN(BLN46),.WL(WL6));
sram_cell_6t_5 inst_cell_6_47 (.BL(BL47),.BLN(BLN47),.WL(WL6));
sram_cell_6t_5 inst_cell_6_48 (.BL(BL48),.BLN(BLN48),.WL(WL6));
sram_cell_6t_5 inst_cell_6_49 (.BL(BL49),.BLN(BLN49),.WL(WL6));
sram_cell_6t_5 inst_cell_6_50 (.BL(BL50),.BLN(BLN50),.WL(WL6));
sram_cell_6t_5 inst_cell_6_51 (.BL(BL51),.BLN(BLN51),.WL(WL6));
sram_cell_6t_5 inst_cell_6_52 (.BL(BL52),.BLN(BLN52),.WL(WL6));
sram_cell_6t_5 inst_cell_6_53 (.BL(BL53),.BLN(BLN53),.WL(WL6));
sram_cell_6t_5 inst_cell_6_54 (.BL(BL54),.BLN(BLN54),.WL(WL6));
sram_cell_6t_5 inst_cell_6_55 (.BL(BL55),.BLN(BLN55),.WL(WL6));
sram_cell_6t_5 inst_cell_6_56 (.BL(BL56),.BLN(BLN56),.WL(WL6));
sram_cell_6t_5 inst_cell_6_57 (.BL(BL57),.BLN(BLN57),.WL(WL6));
sram_cell_6t_5 inst_cell_6_58 (.BL(BL58),.BLN(BLN58),.WL(WL6));
sram_cell_6t_5 inst_cell_6_59 (.BL(BL59),.BLN(BLN59),.WL(WL6));
sram_cell_6t_5 inst_cell_6_60 (.BL(BL60),.BLN(BLN60),.WL(WL6));
sram_cell_6t_5 inst_cell_6_61 (.BL(BL61),.BLN(BLN61),.WL(WL6));
sram_cell_6t_5 inst_cell_6_62 (.BL(BL62),.BLN(BLN62),.WL(WL6));
sram_cell_6t_5 inst_cell_6_63 (.BL(BL63),.BLN(BLN63),.WL(WL6));
sram_cell_6t_5 inst_cell_6_64 (.BL(BL64),.BLN(BLN64),.WL(WL6));
sram_cell_6t_5 inst_cell_6_65 (.BL(BL65),.BLN(BLN65),.WL(WL6));
sram_cell_6t_5 inst_cell_6_66 (.BL(BL66),.BLN(BLN66),.WL(WL6));
sram_cell_6t_5 inst_cell_6_67 (.BL(BL67),.BLN(BLN67),.WL(WL6));
sram_cell_6t_5 inst_cell_6_68 (.BL(BL68),.BLN(BLN68),.WL(WL6));
sram_cell_6t_5 inst_cell_6_69 (.BL(BL69),.BLN(BLN69),.WL(WL6));
sram_cell_6t_5 inst_cell_6_70 (.BL(BL70),.BLN(BLN70),.WL(WL6));
sram_cell_6t_5 inst_cell_6_71 (.BL(BL71),.BLN(BLN71),.WL(WL6));
sram_cell_6t_5 inst_cell_6_72 (.BL(BL72),.BLN(BLN72),.WL(WL6));
sram_cell_6t_5 inst_cell_6_73 (.BL(BL73),.BLN(BLN73),.WL(WL6));
sram_cell_6t_5 inst_cell_6_74 (.BL(BL74),.BLN(BLN74),.WL(WL6));
sram_cell_6t_5 inst_cell_6_75 (.BL(BL75),.BLN(BLN75),.WL(WL6));
sram_cell_6t_5 inst_cell_6_76 (.BL(BL76),.BLN(BLN76),.WL(WL6));
sram_cell_6t_5 inst_cell_6_77 (.BL(BL77),.BLN(BLN77),.WL(WL6));
sram_cell_6t_5 inst_cell_6_78 (.BL(BL78),.BLN(BLN78),.WL(WL6));
sram_cell_6t_5 inst_cell_6_79 (.BL(BL79),.BLN(BLN79),.WL(WL6));
sram_cell_6t_5 inst_cell_6_80 (.BL(BL80),.BLN(BLN80),.WL(WL6));
sram_cell_6t_5 inst_cell_6_81 (.BL(BL81),.BLN(BLN81),.WL(WL6));
sram_cell_6t_5 inst_cell_6_82 (.BL(BL82),.BLN(BLN82),.WL(WL6));
sram_cell_6t_5 inst_cell_6_83 (.BL(BL83),.BLN(BLN83),.WL(WL6));
sram_cell_6t_5 inst_cell_6_84 (.BL(BL84),.BLN(BLN84),.WL(WL6));
sram_cell_6t_5 inst_cell_6_85 (.BL(BL85),.BLN(BLN85),.WL(WL6));
sram_cell_6t_5 inst_cell_6_86 (.BL(BL86),.BLN(BLN86),.WL(WL6));
sram_cell_6t_5 inst_cell_6_87 (.BL(BL87),.BLN(BLN87),.WL(WL6));
sram_cell_6t_5 inst_cell_6_88 (.BL(BL88),.BLN(BLN88),.WL(WL6));
sram_cell_6t_5 inst_cell_6_89 (.BL(BL89),.BLN(BLN89),.WL(WL6));
sram_cell_6t_5 inst_cell_6_90 (.BL(BL90),.BLN(BLN90),.WL(WL6));
sram_cell_6t_5 inst_cell_6_91 (.BL(BL91),.BLN(BLN91),.WL(WL6));
sram_cell_6t_5 inst_cell_6_92 (.BL(BL92),.BLN(BLN92),.WL(WL6));
sram_cell_6t_5 inst_cell_6_93 (.BL(BL93),.BLN(BLN93),.WL(WL6));
sram_cell_6t_5 inst_cell_6_94 (.BL(BL94),.BLN(BLN94),.WL(WL6));
sram_cell_6t_5 inst_cell_6_95 (.BL(BL95),.BLN(BLN95),.WL(WL6));
sram_cell_6t_5 inst_cell_6_96 (.BL(BL96),.BLN(BLN96),.WL(WL6));
sram_cell_6t_5 inst_cell_6_97 (.BL(BL97),.BLN(BLN97),.WL(WL6));
sram_cell_6t_5 inst_cell_6_98 (.BL(BL98),.BLN(BLN98),.WL(WL6));
sram_cell_6t_5 inst_cell_6_99 (.BL(BL99),.BLN(BLN99),.WL(WL6));
sram_cell_6t_5 inst_cell_6_100 (.BL(BL100),.BLN(BLN100),.WL(WL6));
sram_cell_6t_5 inst_cell_6_101 (.BL(BL101),.BLN(BLN101),.WL(WL6));
sram_cell_6t_5 inst_cell_6_102 (.BL(BL102),.BLN(BLN102),.WL(WL6));
sram_cell_6t_5 inst_cell_6_103 (.BL(BL103),.BLN(BLN103),.WL(WL6));
sram_cell_6t_5 inst_cell_6_104 (.BL(BL104),.BLN(BLN104),.WL(WL6));
sram_cell_6t_5 inst_cell_6_105 (.BL(BL105),.BLN(BLN105),.WL(WL6));
sram_cell_6t_5 inst_cell_6_106 (.BL(BL106),.BLN(BLN106),.WL(WL6));
sram_cell_6t_5 inst_cell_6_107 (.BL(BL107),.BLN(BLN107),.WL(WL6));
sram_cell_6t_5 inst_cell_6_108 (.BL(BL108),.BLN(BLN108),.WL(WL6));
sram_cell_6t_5 inst_cell_6_109 (.BL(BL109),.BLN(BLN109),.WL(WL6));
sram_cell_6t_5 inst_cell_6_110 (.BL(BL110),.BLN(BLN110),.WL(WL6));
sram_cell_6t_5 inst_cell_6_111 (.BL(BL111),.BLN(BLN111),.WL(WL6));
sram_cell_6t_5 inst_cell_6_112 (.BL(BL112),.BLN(BLN112),.WL(WL6));
sram_cell_6t_5 inst_cell_6_113 (.BL(BL113),.BLN(BLN113),.WL(WL6));
sram_cell_6t_5 inst_cell_6_114 (.BL(BL114),.BLN(BLN114),.WL(WL6));
sram_cell_6t_5 inst_cell_6_115 (.BL(BL115),.BLN(BLN115),.WL(WL6));
sram_cell_6t_5 inst_cell_6_116 (.BL(BL116),.BLN(BLN116),.WL(WL6));
sram_cell_6t_5 inst_cell_6_117 (.BL(BL117),.BLN(BLN117),.WL(WL6));
sram_cell_6t_5 inst_cell_6_118 (.BL(BL118),.BLN(BLN118),.WL(WL6));
sram_cell_6t_5 inst_cell_6_119 (.BL(BL119),.BLN(BLN119),.WL(WL6));
sram_cell_6t_5 inst_cell_6_120 (.BL(BL120),.BLN(BLN120),.WL(WL6));
sram_cell_6t_5 inst_cell_6_121 (.BL(BL121),.BLN(BLN121),.WL(WL6));
sram_cell_6t_5 inst_cell_6_122 (.BL(BL122),.BLN(BLN122),.WL(WL6));
sram_cell_6t_5 inst_cell_6_123 (.BL(BL123),.BLN(BLN123),.WL(WL6));
sram_cell_6t_5 inst_cell_6_124 (.BL(BL124),.BLN(BLN124),.WL(WL6));
sram_cell_6t_5 inst_cell_6_125 (.BL(BL125),.BLN(BLN125),.WL(WL6));
sram_cell_6t_5 inst_cell_6_126 (.BL(BL126),.BLN(BLN126),.WL(WL6));
sram_cell_6t_5 inst_cell_6_127 (.BL(BL127),.BLN(BLN127),.WL(WL6));
sram_cell_6t_5 inst_cell_7_0 (.BL(BL0),.BLN(BLN0),.WL(WL7));
sram_cell_6t_5 inst_cell_7_1 (.BL(BL1),.BLN(BLN1),.WL(WL7));
sram_cell_6t_5 inst_cell_7_2 (.BL(BL2),.BLN(BLN2),.WL(WL7));
sram_cell_6t_5 inst_cell_7_3 (.BL(BL3),.BLN(BLN3),.WL(WL7));
sram_cell_6t_5 inst_cell_7_4 (.BL(BL4),.BLN(BLN4),.WL(WL7));
sram_cell_6t_5 inst_cell_7_5 (.BL(BL5),.BLN(BLN5),.WL(WL7));
sram_cell_6t_5 inst_cell_7_6 (.BL(BL6),.BLN(BLN6),.WL(WL7));
sram_cell_6t_5 inst_cell_7_7 (.BL(BL7),.BLN(BLN7),.WL(WL7));
sram_cell_6t_5 inst_cell_7_8 (.BL(BL8),.BLN(BLN8),.WL(WL7));
sram_cell_6t_5 inst_cell_7_9 (.BL(BL9),.BLN(BLN9),.WL(WL7));
sram_cell_6t_5 inst_cell_7_10 (.BL(BL10),.BLN(BLN10),.WL(WL7));
sram_cell_6t_5 inst_cell_7_11 (.BL(BL11),.BLN(BLN11),.WL(WL7));
sram_cell_6t_5 inst_cell_7_12 (.BL(BL12),.BLN(BLN12),.WL(WL7));
sram_cell_6t_5 inst_cell_7_13 (.BL(BL13),.BLN(BLN13),.WL(WL7));
sram_cell_6t_5 inst_cell_7_14 (.BL(BL14),.BLN(BLN14),.WL(WL7));
sram_cell_6t_5 inst_cell_7_15 (.BL(BL15),.BLN(BLN15),.WL(WL7));
sram_cell_6t_5 inst_cell_7_16 (.BL(BL16),.BLN(BLN16),.WL(WL7));
sram_cell_6t_5 inst_cell_7_17 (.BL(BL17),.BLN(BLN17),.WL(WL7));
sram_cell_6t_5 inst_cell_7_18 (.BL(BL18),.BLN(BLN18),.WL(WL7));
sram_cell_6t_5 inst_cell_7_19 (.BL(BL19),.BLN(BLN19),.WL(WL7));
sram_cell_6t_5 inst_cell_7_20 (.BL(BL20),.BLN(BLN20),.WL(WL7));
sram_cell_6t_5 inst_cell_7_21 (.BL(BL21),.BLN(BLN21),.WL(WL7));
sram_cell_6t_5 inst_cell_7_22 (.BL(BL22),.BLN(BLN22),.WL(WL7));
sram_cell_6t_5 inst_cell_7_23 (.BL(BL23),.BLN(BLN23),.WL(WL7));
sram_cell_6t_5 inst_cell_7_24 (.BL(BL24),.BLN(BLN24),.WL(WL7));
sram_cell_6t_5 inst_cell_7_25 (.BL(BL25),.BLN(BLN25),.WL(WL7));
sram_cell_6t_5 inst_cell_7_26 (.BL(BL26),.BLN(BLN26),.WL(WL7));
sram_cell_6t_5 inst_cell_7_27 (.BL(BL27),.BLN(BLN27),.WL(WL7));
sram_cell_6t_5 inst_cell_7_28 (.BL(BL28),.BLN(BLN28),.WL(WL7));
sram_cell_6t_5 inst_cell_7_29 (.BL(BL29),.BLN(BLN29),.WL(WL7));
sram_cell_6t_5 inst_cell_7_30 (.BL(BL30),.BLN(BLN30),.WL(WL7));
sram_cell_6t_5 inst_cell_7_31 (.BL(BL31),.BLN(BLN31),.WL(WL7));
sram_cell_6t_5 inst_cell_7_32 (.BL(BL32),.BLN(BLN32),.WL(WL7));
sram_cell_6t_5 inst_cell_7_33 (.BL(BL33),.BLN(BLN33),.WL(WL7));
sram_cell_6t_5 inst_cell_7_34 (.BL(BL34),.BLN(BLN34),.WL(WL7));
sram_cell_6t_5 inst_cell_7_35 (.BL(BL35),.BLN(BLN35),.WL(WL7));
sram_cell_6t_5 inst_cell_7_36 (.BL(BL36),.BLN(BLN36),.WL(WL7));
sram_cell_6t_5 inst_cell_7_37 (.BL(BL37),.BLN(BLN37),.WL(WL7));
sram_cell_6t_5 inst_cell_7_38 (.BL(BL38),.BLN(BLN38),.WL(WL7));
sram_cell_6t_5 inst_cell_7_39 (.BL(BL39),.BLN(BLN39),.WL(WL7));
sram_cell_6t_5 inst_cell_7_40 (.BL(BL40),.BLN(BLN40),.WL(WL7));
sram_cell_6t_5 inst_cell_7_41 (.BL(BL41),.BLN(BLN41),.WL(WL7));
sram_cell_6t_5 inst_cell_7_42 (.BL(BL42),.BLN(BLN42),.WL(WL7));
sram_cell_6t_5 inst_cell_7_43 (.BL(BL43),.BLN(BLN43),.WL(WL7));
sram_cell_6t_5 inst_cell_7_44 (.BL(BL44),.BLN(BLN44),.WL(WL7));
sram_cell_6t_5 inst_cell_7_45 (.BL(BL45),.BLN(BLN45),.WL(WL7));
sram_cell_6t_5 inst_cell_7_46 (.BL(BL46),.BLN(BLN46),.WL(WL7));
sram_cell_6t_5 inst_cell_7_47 (.BL(BL47),.BLN(BLN47),.WL(WL7));
sram_cell_6t_5 inst_cell_7_48 (.BL(BL48),.BLN(BLN48),.WL(WL7));
sram_cell_6t_5 inst_cell_7_49 (.BL(BL49),.BLN(BLN49),.WL(WL7));
sram_cell_6t_5 inst_cell_7_50 (.BL(BL50),.BLN(BLN50),.WL(WL7));
sram_cell_6t_5 inst_cell_7_51 (.BL(BL51),.BLN(BLN51),.WL(WL7));
sram_cell_6t_5 inst_cell_7_52 (.BL(BL52),.BLN(BLN52),.WL(WL7));
sram_cell_6t_5 inst_cell_7_53 (.BL(BL53),.BLN(BLN53),.WL(WL7));
sram_cell_6t_5 inst_cell_7_54 (.BL(BL54),.BLN(BLN54),.WL(WL7));
sram_cell_6t_5 inst_cell_7_55 (.BL(BL55),.BLN(BLN55),.WL(WL7));
sram_cell_6t_5 inst_cell_7_56 (.BL(BL56),.BLN(BLN56),.WL(WL7));
sram_cell_6t_5 inst_cell_7_57 (.BL(BL57),.BLN(BLN57),.WL(WL7));
sram_cell_6t_5 inst_cell_7_58 (.BL(BL58),.BLN(BLN58),.WL(WL7));
sram_cell_6t_5 inst_cell_7_59 (.BL(BL59),.BLN(BLN59),.WL(WL7));
sram_cell_6t_5 inst_cell_7_60 (.BL(BL60),.BLN(BLN60),.WL(WL7));
sram_cell_6t_5 inst_cell_7_61 (.BL(BL61),.BLN(BLN61),.WL(WL7));
sram_cell_6t_5 inst_cell_7_62 (.BL(BL62),.BLN(BLN62),.WL(WL7));
sram_cell_6t_5 inst_cell_7_63 (.BL(BL63),.BLN(BLN63),.WL(WL7));
sram_cell_6t_5 inst_cell_7_64 (.BL(BL64),.BLN(BLN64),.WL(WL7));
sram_cell_6t_5 inst_cell_7_65 (.BL(BL65),.BLN(BLN65),.WL(WL7));
sram_cell_6t_5 inst_cell_7_66 (.BL(BL66),.BLN(BLN66),.WL(WL7));
sram_cell_6t_5 inst_cell_7_67 (.BL(BL67),.BLN(BLN67),.WL(WL7));
sram_cell_6t_5 inst_cell_7_68 (.BL(BL68),.BLN(BLN68),.WL(WL7));
sram_cell_6t_5 inst_cell_7_69 (.BL(BL69),.BLN(BLN69),.WL(WL7));
sram_cell_6t_5 inst_cell_7_70 (.BL(BL70),.BLN(BLN70),.WL(WL7));
sram_cell_6t_5 inst_cell_7_71 (.BL(BL71),.BLN(BLN71),.WL(WL7));
sram_cell_6t_5 inst_cell_7_72 (.BL(BL72),.BLN(BLN72),.WL(WL7));
sram_cell_6t_5 inst_cell_7_73 (.BL(BL73),.BLN(BLN73),.WL(WL7));
sram_cell_6t_5 inst_cell_7_74 (.BL(BL74),.BLN(BLN74),.WL(WL7));
sram_cell_6t_5 inst_cell_7_75 (.BL(BL75),.BLN(BLN75),.WL(WL7));
sram_cell_6t_5 inst_cell_7_76 (.BL(BL76),.BLN(BLN76),.WL(WL7));
sram_cell_6t_5 inst_cell_7_77 (.BL(BL77),.BLN(BLN77),.WL(WL7));
sram_cell_6t_5 inst_cell_7_78 (.BL(BL78),.BLN(BLN78),.WL(WL7));
sram_cell_6t_5 inst_cell_7_79 (.BL(BL79),.BLN(BLN79),.WL(WL7));
sram_cell_6t_5 inst_cell_7_80 (.BL(BL80),.BLN(BLN80),.WL(WL7));
sram_cell_6t_5 inst_cell_7_81 (.BL(BL81),.BLN(BLN81),.WL(WL7));
sram_cell_6t_5 inst_cell_7_82 (.BL(BL82),.BLN(BLN82),.WL(WL7));
sram_cell_6t_5 inst_cell_7_83 (.BL(BL83),.BLN(BLN83),.WL(WL7));
sram_cell_6t_5 inst_cell_7_84 (.BL(BL84),.BLN(BLN84),.WL(WL7));
sram_cell_6t_5 inst_cell_7_85 (.BL(BL85),.BLN(BLN85),.WL(WL7));
sram_cell_6t_5 inst_cell_7_86 (.BL(BL86),.BLN(BLN86),.WL(WL7));
sram_cell_6t_5 inst_cell_7_87 (.BL(BL87),.BLN(BLN87),.WL(WL7));
sram_cell_6t_5 inst_cell_7_88 (.BL(BL88),.BLN(BLN88),.WL(WL7));
sram_cell_6t_5 inst_cell_7_89 (.BL(BL89),.BLN(BLN89),.WL(WL7));
sram_cell_6t_5 inst_cell_7_90 (.BL(BL90),.BLN(BLN90),.WL(WL7));
sram_cell_6t_5 inst_cell_7_91 (.BL(BL91),.BLN(BLN91),.WL(WL7));
sram_cell_6t_5 inst_cell_7_92 (.BL(BL92),.BLN(BLN92),.WL(WL7));
sram_cell_6t_5 inst_cell_7_93 (.BL(BL93),.BLN(BLN93),.WL(WL7));
sram_cell_6t_5 inst_cell_7_94 (.BL(BL94),.BLN(BLN94),.WL(WL7));
sram_cell_6t_5 inst_cell_7_95 (.BL(BL95),.BLN(BLN95),.WL(WL7));
sram_cell_6t_5 inst_cell_7_96 (.BL(BL96),.BLN(BLN96),.WL(WL7));
sram_cell_6t_5 inst_cell_7_97 (.BL(BL97),.BLN(BLN97),.WL(WL7));
sram_cell_6t_5 inst_cell_7_98 (.BL(BL98),.BLN(BLN98),.WL(WL7));
sram_cell_6t_5 inst_cell_7_99 (.BL(BL99),.BLN(BLN99),.WL(WL7));
sram_cell_6t_5 inst_cell_7_100 (.BL(BL100),.BLN(BLN100),.WL(WL7));
sram_cell_6t_5 inst_cell_7_101 (.BL(BL101),.BLN(BLN101),.WL(WL7));
sram_cell_6t_5 inst_cell_7_102 (.BL(BL102),.BLN(BLN102),.WL(WL7));
sram_cell_6t_5 inst_cell_7_103 (.BL(BL103),.BLN(BLN103),.WL(WL7));
sram_cell_6t_5 inst_cell_7_104 (.BL(BL104),.BLN(BLN104),.WL(WL7));
sram_cell_6t_5 inst_cell_7_105 (.BL(BL105),.BLN(BLN105),.WL(WL7));
sram_cell_6t_5 inst_cell_7_106 (.BL(BL106),.BLN(BLN106),.WL(WL7));
sram_cell_6t_5 inst_cell_7_107 (.BL(BL107),.BLN(BLN107),.WL(WL7));
sram_cell_6t_5 inst_cell_7_108 (.BL(BL108),.BLN(BLN108),.WL(WL7));
sram_cell_6t_5 inst_cell_7_109 (.BL(BL109),.BLN(BLN109),.WL(WL7));
sram_cell_6t_5 inst_cell_7_110 (.BL(BL110),.BLN(BLN110),.WL(WL7));
sram_cell_6t_5 inst_cell_7_111 (.BL(BL111),.BLN(BLN111),.WL(WL7));
sram_cell_6t_5 inst_cell_7_112 (.BL(BL112),.BLN(BLN112),.WL(WL7));
sram_cell_6t_5 inst_cell_7_113 (.BL(BL113),.BLN(BLN113),.WL(WL7));
sram_cell_6t_5 inst_cell_7_114 (.BL(BL114),.BLN(BLN114),.WL(WL7));
sram_cell_6t_5 inst_cell_7_115 (.BL(BL115),.BLN(BLN115),.WL(WL7));
sram_cell_6t_5 inst_cell_7_116 (.BL(BL116),.BLN(BLN116),.WL(WL7));
sram_cell_6t_5 inst_cell_7_117 (.BL(BL117),.BLN(BLN117),.WL(WL7));
sram_cell_6t_5 inst_cell_7_118 (.BL(BL118),.BLN(BLN118),.WL(WL7));
sram_cell_6t_5 inst_cell_7_119 (.BL(BL119),.BLN(BLN119),.WL(WL7));
sram_cell_6t_5 inst_cell_7_120 (.BL(BL120),.BLN(BLN120),.WL(WL7));
sram_cell_6t_5 inst_cell_7_121 (.BL(BL121),.BLN(BLN121),.WL(WL7));
sram_cell_6t_5 inst_cell_7_122 (.BL(BL122),.BLN(BLN122),.WL(WL7));
sram_cell_6t_5 inst_cell_7_123 (.BL(BL123),.BLN(BLN123),.WL(WL7));
sram_cell_6t_5 inst_cell_7_124 (.BL(BL124),.BLN(BLN124),.WL(WL7));
sram_cell_6t_5 inst_cell_7_125 (.BL(BL125),.BLN(BLN125),.WL(WL7));
sram_cell_6t_5 inst_cell_7_126 (.BL(BL126),.BLN(BLN126),.WL(WL7));
sram_cell_6t_5 inst_cell_7_127 (.BL(BL127),.BLN(BLN127),.WL(WL7));
sram_cell_6t_5 inst_cell_8_0 (.BL(BL0),.BLN(BLN0),.WL(WL8));
sram_cell_6t_5 inst_cell_8_1 (.BL(BL1),.BLN(BLN1),.WL(WL8));
sram_cell_6t_5 inst_cell_8_2 (.BL(BL2),.BLN(BLN2),.WL(WL8));
sram_cell_6t_5 inst_cell_8_3 (.BL(BL3),.BLN(BLN3),.WL(WL8));
sram_cell_6t_5 inst_cell_8_4 (.BL(BL4),.BLN(BLN4),.WL(WL8));
sram_cell_6t_5 inst_cell_8_5 (.BL(BL5),.BLN(BLN5),.WL(WL8));
sram_cell_6t_5 inst_cell_8_6 (.BL(BL6),.BLN(BLN6),.WL(WL8));
sram_cell_6t_5 inst_cell_8_7 (.BL(BL7),.BLN(BLN7),.WL(WL8));
sram_cell_6t_5 inst_cell_8_8 (.BL(BL8),.BLN(BLN8),.WL(WL8));
sram_cell_6t_5 inst_cell_8_9 (.BL(BL9),.BLN(BLN9),.WL(WL8));
sram_cell_6t_5 inst_cell_8_10 (.BL(BL10),.BLN(BLN10),.WL(WL8));
sram_cell_6t_5 inst_cell_8_11 (.BL(BL11),.BLN(BLN11),.WL(WL8));
sram_cell_6t_5 inst_cell_8_12 (.BL(BL12),.BLN(BLN12),.WL(WL8));
sram_cell_6t_5 inst_cell_8_13 (.BL(BL13),.BLN(BLN13),.WL(WL8));
sram_cell_6t_5 inst_cell_8_14 (.BL(BL14),.BLN(BLN14),.WL(WL8));
sram_cell_6t_5 inst_cell_8_15 (.BL(BL15),.BLN(BLN15),.WL(WL8));
sram_cell_6t_5 inst_cell_8_16 (.BL(BL16),.BLN(BLN16),.WL(WL8));
sram_cell_6t_5 inst_cell_8_17 (.BL(BL17),.BLN(BLN17),.WL(WL8));
sram_cell_6t_5 inst_cell_8_18 (.BL(BL18),.BLN(BLN18),.WL(WL8));
sram_cell_6t_5 inst_cell_8_19 (.BL(BL19),.BLN(BLN19),.WL(WL8));
sram_cell_6t_5 inst_cell_8_20 (.BL(BL20),.BLN(BLN20),.WL(WL8));
sram_cell_6t_5 inst_cell_8_21 (.BL(BL21),.BLN(BLN21),.WL(WL8));
sram_cell_6t_5 inst_cell_8_22 (.BL(BL22),.BLN(BLN22),.WL(WL8));
sram_cell_6t_5 inst_cell_8_23 (.BL(BL23),.BLN(BLN23),.WL(WL8));
sram_cell_6t_5 inst_cell_8_24 (.BL(BL24),.BLN(BLN24),.WL(WL8));
sram_cell_6t_5 inst_cell_8_25 (.BL(BL25),.BLN(BLN25),.WL(WL8));
sram_cell_6t_5 inst_cell_8_26 (.BL(BL26),.BLN(BLN26),.WL(WL8));
sram_cell_6t_5 inst_cell_8_27 (.BL(BL27),.BLN(BLN27),.WL(WL8));
sram_cell_6t_5 inst_cell_8_28 (.BL(BL28),.BLN(BLN28),.WL(WL8));
sram_cell_6t_5 inst_cell_8_29 (.BL(BL29),.BLN(BLN29),.WL(WL8));
sram_cell_6t_5 inst_cell_8_30 (.BL(BL30),.BLN(BLN30),.WL(WL8));
sram_cell_6t_5 inst_cell_8_31 (.BL(BL31),.BLN(BLN31),.WL(WL8));
sram_cell_6t_5 inst_cell_8_32 (.BL(BL32),.BLN(BLN32),.WL(WL8));
sram_cell_6t_5 inst_cell_8_33 (.BL(BL33),.BLN(BLN33),.WL(WL8));
sram_cell_6t_5 inst_cell_8_34 (.BL(BL34),.BLN(BLN34),.WL(WL8));
sram_cell_6t_5 inst_cell_8_35 (.BL(BL35),.BLN(BLN35),.WL(WL8));
sram_cell_6t_5 inst_cell_8_36 (.BL(BL36),.BLN(BLN36),.WL(WL8));
sram_cell_6t_5 inst_cell_8_37 (.BL(BL37),.BLN(BLN37),.WL(WL8));
sram_cell_6t_5 inst_cell_8_38 (.BL(BL38),.BLN(BLN38),.WL(WL8));
sram_cell_6t_5 inst_cell_8_39 (.BL(BL39),.BLN(BLN39),.WL(WL8));
sram_cell_6t_5 inst_cell_8_40 (.BL(BL40),.BLN(BLN40),.WL(WL8));
sram_cell_6t_5 inst_cell_8_41 (.BL(BL41),.BLN(BLN41),.WL(WL8));
sram_cell_6t_5 inst_cell_8_42 (.BL(BL42),.BLN(BLN42),.WL(WL8));
sram_cell_6t_5 inst_cell_8_43 (.BL(BL43),.BLN(BLN43),.WL(WL8));
sram_cell_6t_5 inst_cell_8_44 (.BL(BL44),.BLN(BLN44),.WL(WL8));
sram_cell_6t_5 inst_cell_8_45 (.BL(BL45),.BLN(BLN45),.WL(WL8));
sram_cell_6t_5 inst_cell_8_46 (.BL(BL46),.BLN(BLN46),.WL(WL8));
sram_cell_6t_5 inst_cell_8_47 (.BL(BL47),.BLN(BLN47),.WL(WL8));
sram_cell_6t_5 inst_cell_8_48 (.BL(BL48),.BLN(BLN48),.WL(WL8));
sram_cell_6t_5 inst_cell_8_49 (.BL(BL49),.BLN(BLN49),.WL(WL8));
sram_cell_6t_5 inst_cell_8_50 (.BL(BL50),.BLN(BLN50),.WL(WL8));
sram_cell_6t_5 inst_cell_8_51 (.BL(BL51),.BLN(BLN51),.WL(WL8));
sram_cell_6t_5 inst_cell_8_52 (.BL(BL52),.BLN(BLN52),.WL(WL8));
sram_cell_6t_5 inst_cell_8_53 (.BL(BL53),.BLN(BLN53),.WL(WL8));
sram_cell_6t_5 inst_cell_8_54 (.BL(BL54),.BLN(BLN54),.WL(WL8));
sram_cell_6t_5 inst_cell_8_55 (.BL(BL55),.BLN(BLN55),.WL(WL8));
sram_cell_6t_5 inst_cell_8_56 (.BL(BL56),.BLN(BLN56),.WL(WL8));
sram_cell_6t_5 inst_cell_8_57 (.BL(BL57),.BLN(BLN57),.WL(WL8));
sram_cell_6t_5 inst_cell_8_58 (.BL(BL58),.BLN(BLN58),.WL(WL8));
sram_cell_6t_5 inst_cell_8_59 (.BL(BL59),.BLN(BLN59),.WL(WL8));
sram_cell_6t_5 inst_cell_8_60 (.BL(BL60),.BLN(BLN60),.WL(WL8));
sram_cell_6t_5 inst_cell_8_61 (.BL(BL61),.BLN(BLN61),.WL(WL8));
sram_cell_6t_5 inst_cell_8_62 (.BL(BL62),.BLN(BLN62),.WL(WL8));
sram_cell_6t_5 inst_cell_8_63 (.BL(BL63),.BLN(BLN63),.WL(WL8));
sram_cell_6t_5 inst_cell_8_64 (.BL(BL64),.BLN(BLN64),.WL(WL8));
sram_cell_6t_5 inst_cell_8_65 (.BL(BL65),.BLN(BLN65),.WL(WL8));
sram_cell_6t_5 inst_cell_8_66 (.BL(BL66),.BLN(BLN66),.WL(WL8));
sram_cell_6t_5 inst_cell_8_67 (.BL(BL67),.BLN(BLN67),.WL(WL8));
sram_cell_6t_5 inst_cell_8_68 (.BL(BL68),.BLN(BLN68),.WL(WL8));
sram_cell_6t_5 inst_cell_8_69 (.BL(BL69),.BLN(BLN69),.WL(WL8));
sram_cell_6t_5 inst_cell_8_70 (.BL(BL70),.BLN(BLN70),.WL(WL8));
sram_cell_6t_5 inst_cell_8_71 (.BL(BL71),.BLN(BLN71),.WL(WL8));
sram_cell_6t_5 inst_cell_8_72 (.BL(BL72),.BLN(BLN72),.WL(WL8));
sram_cell_6t_5 inst_cell_8_73 (.BL(BL73),.BLN(BLN73),.WL(WL8));
sram_cell_6t_5 inst_cell_8_74 (.BL(BL74),.BLN(BLN74),.WL(WL8));
sram_cell_6t_5 inst_cell_8_75 (.BL(BL75),.BLN(BLN75),.WL(WL8));
sram_cell_6t_5 inst_cell_8_76 (.BL(BL76),.BLN(BLN76),.WL(WL8));
sram_cell_6t_5 inst_cell_8_77 (.BL(BL77),.BLN(BLN77),.WL(WL8));
sram_cell_6t_5 inst_cell_8_78 (.BL(BL78),.BLN(BLN78),.WL(WL8));
sram_cell_6t_5 inst_cell_8_79 (.BL(BL79),.BLN(BLN79),.WL(WL8));
sram_cell_6t_5 inst_cell_8_80 (.BL(BL80),.BLN(BLN80),.WL(WL8));
sram_cell_6t_5 inst_cell_8_81 (.BL(BL81),.BLN(BLN81),.WL(WL8));
sram_cell_6t_5 inst_cell_8_82 (.BL(BL82),.BLN(BLN82),.WL(WL8));
sram_cell_6t_5 inst_cell_8_83 (.BL(BL83),.BLN(BLN83),.WL(WL8));
sram_cell_6t_5 inst_cell_8_84 (.BL(BL84),.BLN(BLN84),.WL(WL8));
sram_cell_6t_5 inst_cell_8_85 (.BL(BL85),.BLN(BLN85),.WL(WL8));
sram_cell_6t_5 inst_cell_8_86 (.BL(BL86),.BLN(BLN86),.WL(WL8));
sram_cell_6t_5 inst_cell_8_87 (.BL(BL87),.BLN(BLN87),.WL(WL8));
sram_cell_6t_5 inst_cell_8_88 (.BL(BL88),.BLN(BLN88),.WL(WL8));
sram_cell_6t_5 inst_cell_8_89 (.BL(BL89),.BLN(BLN89),.WL(WL8));
sram_cell_6t_5 inst_cell_8_90 (.BL(BL90),.BLN(BLN90),.WL(WL8));
sram_cell_6t_5 inst_cell_8_91 (.BL(BL91),.BLN(BLN91),.WL(WL8));
sram_cell_6t_5 inst_cell_8_92 (.BL(BL92),.BLN(BLN92),.WL(WL8));
sram_cell_6t_5 inst_cell_8_93 (.BL(BL93),.BLN(BLN93),.WL(WL8));
sram_cell_6t_5 inst_cell_8_94 (.BL(BL94),.BLN(BLN94),.WL(WL8));
sram_cell_6t_5 inst_cell_8_95 (.BL(BL95),.BLN(BLN95),.WL(WL8));
sram_cell_6t_5 inst_cell_8_96 (.BL(BL96),.BLN(BLN96),.WL(WL8));
sram_cell_6t_5 inst_cell_8_97 (.BL(BL97),.BLN(BLN97),.WL(WL8));
sram_cell_6t_5 inst_cell_8_98 (.BL(BL98),.BLN(BLN98),.WL(WL8));
sram_cell_6t_5 inst_cell_8_99 (.BL(BL99),.BLN(BLN99),.WL(WL8));
sram_cell_6t_5 inst_cell_8_100 (.BL(BL100),.BLN(BLN100),.WL(WL8));
sram_cell_6t_5 inst_cell_8_101 (.BL(BL101),.BLN(BLN101),.WL(WL8));
sram_cell_6t_5 inst_cell_8_102 (.BL(BL102),.BLN(BLN102),.WL(WL8));
sram_cell_6t_5 inst_cell_8_103 (.BL(BL103),.BLN(BLN103),.WL(WL8));
sram_cell_6t_5 inst_cell_8_104 (.BL(BL104),.BLN(BLN104),.WL(WL8));
sram_cell_6t_5 inst_cell_8_105 (.BL(BL105),.BLN(BLN105),.WL(WL8));
sram_cell_6t_5 inst_cell_8_106 (.BL(BL106),.BLN(BLN106),.WL(WL8));
sram_cell_6t_5 inst_cell_8_107 (.BL(BL107),.BLN(BLN107),.WL(WL8));
sram_cell_6t_5 inst_cell_8_108 (.BL(BL108),.BLN(BLN108),.WL(WL8));
sram_cell_6t_5 inst_cell_8_109 (.BL(BL109),.BLN(BLN109),.WL(WL8));
sram_cell_6t_5 inst_cell_8_110 (.BL(BL110),.BLN(BLN110),.WL(WL8));
sram_cell_6t_5 inst_cell_8_111 (.BL(BL111),.BLN(BLN111),.WL(WL8));
sram_cell_6t_5 inst_cell_8_112 (.BL(BL112),.BLN(BLN112),.WL(WL8));
sram_cell_6t_5 inst_cell_8_113 (.BL(BL113),.BLN(BLN113),.WL(WL8));
sram_cell_6t_5 inst_cell_8_114 (.BL(BL114),.BLN(BLN114),.WL(WL8));
sram_cell_6t_5 inst_cell_8_115 (.BL(BL115),.BLN(BLN115),.WL(WL8));
sram_cell_6t_5 inst_cell_8_116 (.BL(BL116),.BLN(BLN116),.WL(WL8));
sram_cell_6t_5 inst_cell_8_117 (.BL(BL117),.BLN(BLN117),.WL(WL8));
sram_cell_6t_5 inst_cell_8_118 (.BL(BL118),.BLN(BLN118),.WL(WL8));
sram_cell_6t_5 inst_cell_8_119 (.BL(BL119),.BLN(BLN119),.WL(WL8));
sram_cell_6t_5 inst_cell_8_120 (.BL(BL120),.BLN(BLN120),.WL(WL8));
sram_cell_6t_5 inst_cell_8_121 (.BL(BL121),.BLN(BLN121),.WL(WL8));
sram_cell_6t_5 inst_cell_8_122 (.BL(BL122),.BLN(BLN122),.WL(WL8));
sram_cell_6t_5 inst_cell_8_123 (.BL(BL123),.BLN(BLN123),.WL(WL8));
sram_cell_6t_5 inst_cell_8_124 (.BL(BL124),.BLN(BLN124),.WL(WL8));
sram_cell_6t_5 inst_cell_8_125 (.BL(BL125),.BLN(BLN125),.WL(WL8));
sram_cell_6t_5 inst_cell_8_126 (.BL(BL126),.BLN(BLN126),.WL(WL8));
sram_cell_6t_5 inst_cell_8_127 (.BL(BL127),.BLN(BLN127),.WL(WL8));
sram_cell_6t_5 inst_cell_9_0 (.BL(BL0),.BLN(BLN0),.WL(WL9));
sram_cell_6t_5 inst_cell_9_1 (.BL(BL1),.BLN(BLN1),.WL(WL9));
sram_cell_6t_5 inst_cell_9_2 (.BL(BL2),.BLN(BLN2),.WL(WL9));
sram_cell_6t_5 inst_cell_9_3 (.BL(BL3),.BLN(BLN3),.WL(WL9));
sram_cell_6t_5 inst_cell_9_4 (.BL(BL4),.BLN(BLN4),.WL(WL9));
sram_cell_6t_5 inst_cell_9_5 (.BL(BL5),.BLN(BLN5),.WL(WL9));
sram_cell_6t_5 inst_cell_9_6 (.BL(BL6),.BLN(BLN6),.WL(WL9));
sram_cell_6t_5 inst_cell_9_7 (.BL(BL7),.BLN(BLN7),.WL(WL9));
sram_cell_6t_5 inst_cell_9_8 (.BL(BL8),.BLN(BLN8),.WL(WL9));
sram_cell_6t_5 inst_cell_9_9 (.BL(BL9),.BLN(BLN9),.WL(WL9));
sram_cell_6t_5 inst_cell_9_10 (.BL(BL10),.BLN(BLN10),.WL(WL9));
sram_cell_6t_5 inst_cell_9_11 (.BL(BL11),.BLN(BLN11),.WL(WL9));
sram_cell_6t_5 inst_cell_9_12 (.BL(BL12),.BLN(BLN12),.WL(WL9));
sram_cell_6t_5 inst_cell_9_13 (.BL(BL13),.BLN(BLN13),.WL(WL9));
sram_cell_6t_5 inst_cell_9_14 (.BL(BL14),.BLN(BLN14),.WL(WL9));
sram_cell_6t_5 inst_cell_9_15 (.BL(BL15),.BLN(BLN15),.WL(WL9));
sram_cell_6t_5 inst_cell_9_16 (.BL(BL16),.BLN(BLN16),.WL(WL9));
sram_cell_6t_5 inst_cell_9_17 (.BL(BL17),.BLN(BLN17),.WL(WL9));
sram_cell_6t_5 inst_cell_9_18 (.BL(BL18),.BLN(BLN18),.WL(WL9));
sram_cell_6t_5 inst_cell_9_19 (.BL(BL19),.BLN(BLN19),.WL(WL9));
sram_cell_6t_5 inst_cell_9_20 (.BL(BL20),.BLN(BLN20),.WL(WL9));
sram_cell_6t_5 inst_cell_9_21 (.BL(BL21),.BLN(BLN21),.WL(WL9));
sram_cell_6t_5 inst_cell_9_22 (.BL(BL22),.BLN(BLN22),.WL(WL9));
sram_cell_6t_5 inst_cell_9_23 (.BL(BL23),.BLN(BLN23),.WL(WL9));
sram_cell_6t_5 inst_cell_9_24 (.BL(BL24),.BLN(BLN24),.WL(WL9));
sram_cell_6t_5 inst_cell_9_25 (.BL(BL25),.BLN(BLN25),.WL(WL9));
sram_cell_6t_5 inst_cell_9_26 (.BL(BL26),.BLN(BLN26),.WL(WL9));
sram_cell_6t_5 inst_cell_9_27 (.BL(BL27),.BLN(BLN27),.WL(WL9));
sram_cell_6t_5 inst_cell_9_28 (.BL(BL28),.BLN(BLN28),.WL(WL9));
sram_cell_6t_5 inst_cell_9_29 (.BL(BL29),.BLN(BLN29),.WL(WL9));
sram_cell_6t_5 inst_cell_9_30 (.BL(BL30),.BLN(BLN30),.WL(WL9));
sram_cell_6t_5 inst_cell_9_31 (.BL(BL31),.BLN(BLN31),.WL(WL9));
sram_cell_6t_5 inst_cell_9_32 (.BL(BL32),.BLN(BLN32),.WL(WL9));
sram_cell_6t_5 inst_cell_9_33 (.BL(BL33),.BLN(BLN33),.WL(WL9));
sram_cell_6t_5 inst_cell_9_34 (.BL(BL34),.BLN(BLN34),.WL(WL9));
sram_cell_6t_5 inst_cell_9_35 (.BL(BL35),.BLN(BLN35),.WL(WL9));
sram_cell_6t_5 inst_cell_9_36 (.BL(BL36),.BLN(BLN36),.WL(WL9));
sram_cell_6t_5 inst_cell_9_37 (.BL(BL37),.BLN(BLN37),.WL(WL9));
sram_cell_6t_5 inst_cell_9_38 (.BL(BL38),.BLN(BLN38),.WL(WL9));
sram_cell_6t_5 inst_cell_9_39 (.BL(BL39),.BLN(BLN39),.WL(WL9));
sram_cell_6t_5 inst_cell_9_40 (.BL(BL40),.BLN(BLN40),.WL(WL9));
sram_cell_6t_5 inst_cell_9_41 (.BL(BL41),.BLN(BLN41),.WL(WL9));
sram_cell_6t_5 inst_cell_9_42 (.BL(BL42),.BLN(BLN42),.WL(WL9));
sram_cell_6t_5 inst_cell_9_43 (.BL(BL43),.BLN(BLN43),.WL(WL9));
sram_cell_6t_5 inst_cell_9_44 (.BL(BL44),.BLN(BLN44),.WL(WL9));
sram_cell_6t_5 inst_cell_9_45 (.BL(BL45),.BLN(BLN45),.WL(WL9));
sram_cell_6t_5 inst_cell_9_46 (.BL(BL46),.BLN(BLN46),.WL(WL9));
sram_cell_6t_5 inst_cell_9_47 (.BL(BL47),.BLN(BLN47),.WL(WL9));
sram_cell_6t_5 inst_cell_9_48 (.BL(BL48),.BLN(BLN48),.WL(WL9));
sram_cell_6t_5 inst_cell_9_49 (.BL(BL49),.BLN(BLN49),.WL(WL9));
sram_cell_6t_5 inst_cell_9_50 (.BL(BL50),.BLN(BLN50),.WL(WL9));
sram_cell_6t_5 inst_cell_9_51 (.BL(BL51),.BLN(BLN51),.WL(WL9));
sram_cell_6t_5 inst_cell_9_52 (.BL(BL52),.BLN(BLN52),.WL(WL9));
sram_cell_6t_5 inst_cell_9_53 (.BL(BL53),.BLN(BLN53),.WL(WL9));
sram_cell_6t_5 inst_cell_9_54 (.BL(BL54),.BLN(BLN54),.WL(WL9));
sram_cell_6t_5 inst_cell_9_55 (.BL(BL55),.BLN(BLN55),.WL(WL9));
sram_cell_6t_5 inst_cell_9_56 (.BL(BL56),.BLN(BLN56),.WL(WL9));
sram_cell_6t_5 inst_cell_9_57 (.BL(BL57),.BLN(BLN57),.WL(WL9));
sram_cell_6t_5 inst_cell_9_58 (.BL(BL58),.BLN(BLN58),.WL(WL9));
sram_cell_6t_5 inst_cell_9_59 (.BL(BL59),.BLN(BLN59),.WL(WL9));
sram_cell_6t_5 inst_cell_9_60 (.BL(BL60),.BLN(BLN60),.WL(WL9));
sram_cell_6t_5 inst_cell_9_61 (.BL(BL61),.BLN(BLN61),.WL(WL9));
sram_cell_6t_5 inst_cell_9_62 (.BL(BL62),.BLN(BLN62),.WL(WL9));
sram_cell_6t_5 inst_cell_9_63 (.BL(BL63),.BLN(BLN63),.WL(WL9));
sram_cell_6t_5 inst_cell_9_64 (.BL(BL64),.BLN(BLN64),.WL(WL9));
sram_cell_6t_5 inst_cell_9_65 (.BL(BL65),.BLN(BLN65),.WL(WL9));
sram_cell_6t_5 inst_cell_9_66 (.BL(BL66),.BLN(BLN66),.WL(WL9));
sram_cell_6t_5 inst_cell_9_67 (.BL(BL67),.BLN(BLN67),.WL(WL9));
sram_cell_6t_5 inst_cell_9_68 (.BL(BL68),.BLN(BLN68),.WL(WL9));
sram_cell_6t_5 inst_cell_9_69 (.BL(BL69),.BLN(BLN69),.WL(WL9));
sram_cell_6t_5 inst_cell_9_70 (.BL(BL70),.BLN(BLN70),.WL(WL9));
sram_cell_6t_5 inst_cell_9_71 (.BL(BL71),.BLN(BLN71),.WL(WL9));
sram_cell_6t_5 inst_cell_9_72 (.BL(BL72),.BLN(BLN72),.WL(WL9));
sram_cell_6t_5 inst_cell_9_73 (.BL(BL73),.BLN(BLN73),.WL(WL9));
sram_cell_6t_5 inst_cell_9_74 (.BL(BL74),.BLN(BLN74),.WL(WL9));
sram_cell_6t_5 inst_cell_9_75 (.BL(BL75),.BLN(BLN75),.WL(WL9));
sram_cell_6t_5 inst_cell_9_76 (.BL(BL76),.BLN(BLN76),.WL(WL9));
sram_cell_6t_5 inst_cell_9_77 (.BL(BL77),.BLN(BLN77),.WL(WL9));
sram_cell_6t_5 inst_cell_9_78 (.BL(BL78),.BLN(BLN78),.WL(WL9));
sram_cell_6t_5 inst_cell_9_79 (.BL(BL79),.BLN(BLN79),.WL(WL9));
sram_cell_6t_5 inst_cell_9_80 (.BL(BL80),.BLN(BLN80),.WL(WL9));
sram_cell_6t_5 inst_cell_9_81 (.BL(BL81),.BLN(BLN81),.WL(WL9));
sram_cell_6t_5 inst_cell_9_82 (.BL(BL82),.BLN(BLN82),.WL(WL9));
sram_cell_6t_5 inst_cell_9_83 (.BL(BL83),.BLN(BLN83),.WL(WL9));
sram_cell_6t_5 inst_cell_9_84 (.BL(BL84),.BLN(BLN84),.WL(WL9));
sram_cell_6t_5 inst_cell_9_85 (.BL(BL85),.BLN(BLN85),.WL(WL9));
sram_cell_6t_5 inst_cell_9_86 (.BL(BL86),.BLN(BLN86),.WL(WL9));
sram_cell_6t_5 inst_cell_9_87 (.BL(BL87),.BLN(BLN87),.WL(WL9));
sram_cell_6t_5 inst_cell_9_88 (.BL(BL88),.BLN(BLN88),.WL(WL9));
sram_cell_6t_5 inst_cell_9_89 (.BL(BL89),.BLN(BLN89),.WL(WL9));
sram_cell_6t_5 inst_cell_9_90 (.BL(BL90),.BLN(BLN90),.WL(WL9));
sram_cell_6t_5 inst_cell_9_91 (.BL(BL91),.BLN(BLN91),.WL(WL9));
sram_cell_6t_5 inst_cell_9_92 (.BL(BL92),.BLN(BLN92),.WL(WL9));
sram_cell_6t_5 inst_cell_9_93 (.BL(BL93),.BLN(BLN93),.WL(WL9));
sram_cell_6t_5 inst_cell_9_94 (.BL(BL94),.BLN(BLN94),.WL(WL9));
sram_cell_6t_5 inst_cell_9_95 (.BL(BL95),.BLN(BLN95),.WL(WL9));
sram_cell_6t_5 inst_cell_9_96 (.BL(BL96),.BLN(BLN96),.WL(WL9));
sram_cell_6t_5 inst_cell_9_97 (.BL(BL97),.BLN(BLN97),.WL(WL9));
sram_cell_6t_5 inst_cell_9_98 (.BL(BL98),.BLN(BLN98),.WL(WL9));
sram_cell_6t_5 inst_cell_9_99 (.BL(BL99),.BLN(BLN99),.WL(WL9));
sram_cell_6t_5 inst_cell_9_100 (.BL(BL100),.BLN(BLN100),.WL(WL9));
sram_cell_6t_5 inst_cell_9_101 (.BL(BL101),.BLN(BLN101),.WL(WL9));
sram_cell_6t_5 inst_cell_9_102 (.BL(BL102),.BLN(BLN102),.WL(WL9));
sram_cell_6t_5 inst_cell_9_103 (.BL(BL103),.BLN(BLN103),.WL(WL9));
sram_cell_6t_5 inst_cell_9_104 (.BL(BL104),.BLN(BLN104),.WL(WL9));
sram_cell_6t_5 inst_cell_9_105 (.BL(BL105),.BLN(BLN105),.WL(WL9));
sram_cell_6t_5 inst_cell_9_106 (.BL(BL106),.BLN(BLN106),.WL(WL9));
sram_cell_6t_5 inst_cell_9_107 (.BL(BL107),.BLN(BLN107),.WL(WL9));
sram_cell_6t_5 inst_cell_9_108 (.BL(BL108),.BLN(BLN108),.WL(WL9));
sram_cell_6t_5 inst_cell_9_109 (.BL(BL109),.BLN(BLN109),.WL(WL9));
sram_cell_6t_5 inst_cell_9_110 (.BL(BL110),.BLN(BLN110),.WL(WL9));
sram_cell_6t_5 inst_cell_9_111 (.BL(BL111),.BLN(BLN111),.WL(WL9));
sram_cell_6t_5 inst_cell_9_112 (.BL(BL112),.BLN(BLN112),.WL(WL9));
sram_cell_6t_5 inst_cell_9_113 (.BL(BL113),.BLN(BLN113),.WL(WL9));
sram_cell_6t_5 inst_cell_9_114 (.BL(BL114),.BLN(BLN114),.WL(WL9));
sram_cell_6t_5 inst_cell_9_115 (.BL(BL115),.BLN(BLN115),.WL(WL9));
sram_cell_6t_5 inst_cell_9_116 (.BL(BL116),.BLN(BLN116),.WL(WL9));
sram_cell_6t_5 inst_cell_9_117 (.BL(BL117),.BLN(BLN117),.WL(WL9));
sram_cell_6t_5 inst_cell_9_118 (.BL(BL118),.BLN(BLN118),.WL(WL9));
sram_cell_6t_5 inst_cell_9_119 (.BL(BL119),.BLN(BLN119),.WL(WL9));
sram_cell_6t_5 inst_cell_9_120 (.BL(BL120),.BLN(BLN120),.WL(WL9));
sram_cell_6t_5 inst_cell_9_121 (.BL(BL121),.BLN(BLN121),.WL(WL9));
sram_cell_6t_5 inst_cell_9_122 (.BL(BL122),.BLN(BLN122),.WL(WL9));
sram_cell_6t_5 inst_cell_9_123 (.BL(BL123),.BLN(BLN123),.WL(WL9));
sram_cell_6t_5 inst_cell_9_124 (.BL(BL124),.BLN(BLN124),.WL(WL9));
sram_cell_6t_5 inst_cell_9_125 (.BL(BL125),.BLN(BLN125),.WL(WL9));
sram_cell_6t_5 inst_cell_9_126 (.BL(BL126),.BLN(BLN126),.WL(WL9));
sram_cell_6t_5 inst_cell_9_127 (.BL(BL127),.BLN(BLN127),.WL(WL9));
sram_cell_6t_5 inst_cell_10_0 (.BL(BL0),.BLN(BLN0),.WL(WL10));
sram_cell_6t_5 inst_cell_10_1 (.BL(BL1),.BLN(BLN1),.WL(WL10));
sram_cell_6t_5 inst_cell_10_2 (.BL(BL2),.BLN(BLN2),.WL(WL10));
sram_cell_6t_5 inst_cell_10_3 (.BL(BL3),.BLN(BLN3),.WL(WL10));
sram_cell_6t_5 inst_cell_10_4 (.BL(BL4),.BLN(BLN4),.WL(WL10));
sram_cell_6t_5 inst_cell_10_5 (.BL(BL5),.BLN(BLN5),.WL(WL10));
sram_cell_6t_5 inst_cell_10_6 (.BL(BL6),.BLN(BLN6),.WL(WL10));
sram_cell_6t_5 inst_cell_10_7 (.BL(BL7),.BLN(BLN7),.WL(WL10));
sram_cell_6t_5 inst_cell_10_8 (.BL(BL8),.BLN(BLN8),.WL(WL10));
sram_cell_6t_5 inst_cell_10_9 (.BL(BL9),.BLN(BLN9),.WL(WL10));
sram_cell_6t_5 inst_cell_10_10 (.BL(BL10),.BLN(BLN10),.WL(WL10));
sram_cell_6t_5 inst_cell_10_11 (.BL(BL11),.BLN(BLN11),.WL(WL10));
sram_cell_6t_5 inst_cell_10_12 (.BL(BL12),.BLN(BLN12),.WL(WL10));
sram_cell_6t_5 inst_cell_10_13 (.BL(BL13),.BLN(BLN13),.WL(WL10));
sram_cell_6t_5 inst_cell_10_14 (.BL(BL14),.BLN(BLN14),.WL(WL10));
sram_cell_6t_5 inst_cell_10_15 (.BL(BL15),.BLN(BLN15),.WL(WL10));
sram_cell_6t_5 inst_cell_10_16 (.BL(BL16),.BLN(BLN16),.WL(WL10));
sram_cell_6t_5 inst_cell_10_17 (.BL(BL17),.BLN(BLN17),.WL(WL10));
sram_cell_6t_5 inst_cell_10_18 (.BL(BL18),.BLN(BLN18),.WL(WL10));
sram_cell_6t_5 inst_cell_10_19 (.BL(BL19),.BLN(BLN19),.WL(WL10));
sram_cell_6t_5 inst_cell_10_20 (.BL(BL20),.BLN(BLN20),.WL(WL10));
sram_cell_6t_5 inst_cell_10_21 (.BL(BL21),.BLN(BLN21),.WL(WL10));
sram_cell_6t_5 inst_cell_10_22 (.BL(BL22),.BLN(BLN22),.WL(WL10));
sram_cell_6t_5 inst_cell_10_23 (.BL(BL23),.BLN(BLN23),.WL(WL10));
sram_cell_6t_5 inst_cell_10_24 (.BL(BL24),.BLN(BLN24),.WL(WL10));
sram_cell_6t_5 inst_cell_10_25 (.BL(BL25),.BLN(BLN25),.WL(WL10));
sram_cell_6t_5 inst_cell_10_26 (.BL(BL26),.BLN(BLN26),.WL(WL10));
sram_cell_6t_5 inst_cell_10_27 (.BL(BL27),.BLN(BLN27),.WL(WL10));
sram_cell_6t_5 inst_cell_10_28 (.BL(BL28),.BLN(BLN28),.WL(WL10));
sram_cell_6t_5 inst_cell_10_29 (.BL(BL29),.BLN(BLN29),.WL(WL10));
sram_cell_6t_5 inst_cell_10_30 (.BL(BL30),.BLN(BLN30),.WL(WL10));
sram_cell_6t_5 inst_cell_10_31 (.BL(BL31),.BLN(BLN31),.WL(WL10));
sram_cell_6t_5 inst_cell_10_32 (.BL(BL32),.BLN(BLN32),.WL(WL10));
sram_cell_6t_5 inst_cell_10_33 (.BL(BL33),.BLN(BLN33),.WL(WL10));
sram_cell_6t_5 inst_cell_10_34 (.BL(BL34),.BLN(BLN34),.WL(WL10));
sram_cell_6t_5 inst_cell_10_35 (.BL(BL35),.BLN(BLN35),.WL(WL10));
sram_cell_6t_5 inst_cell_10_36 (.BL(BL36),.BLN(BLN36),.WL(WL10));
sram_cell_6t_5 inst_cell_10_37 (.BL(BL37),.BLN(BLN37),.WL(WL10));
sram_cell_6t_5 inst_cell_10_38 (.BL(BL38),.BLN(BLN38),.WL(WL10));
sram_cell_6t_5 inst_cell_10_39 (.BL(BL39),.BLN(BLN39),.WL(WL10));
sram_cell_6t_5 inst_cell_10_40 (.BL(BL40),.BLN(BLN40),.WL(WL10));
sram_cell_6t_5 inst_cell_10_41 (.BL(BL41),.BLN(BLN41),.WL(WL10));
sram_cell_6t_5 inst_cell_10_42 (.BL(BL42),.BLN(BLN42),.WL(WL10));
sram_cell_6t_5 inst_cell_10_43 (.BL(BL43),.BLN(BLN43),.WL(WL10));
sram_cell_6t_5 inst_cell_10_44 (.BL(BL44),.BLN(BLN44),.WL(WL10));
sram_cell_6t_5 inst_cell_10_45 (.BL(BL45),.BLN(BLN45),.WL(WL10));
sram_cell_6t_5 inst_cell_10_46 (.BL(BL46),.BLN(BLN46),.WL(WL10));
sram_cell_6t_5 inst_cell_10_47 (.BL(BL47),.BLN(BLN47),.WL(WL10));
sram_cell_6t_5 inst_cell_10_48 (.BL(BL48),.BLN(BLN48),.WL(WL10));
sram_cell_6t_5 inst_cell_10_49 (.BL(BL49),.BLN(BLN49),.WL(WL10));
sram_cell_6t_5 inst_cell_10_50 (.BL(BL50),.BLN(BLN50),.WL(WL10));
sram_cell_6t_5 inst_cell_10_51 (.BL(BL51),.BLN(BLN51),.WL(WL10));
sram_cell_6t_5 inst_cell_10_52 (.BL(BL52),.BLN(BLN52),.WL(WL10));
sram_cell_6t_5 inst_cell_10_53 (.BL(BL53),.BLN(BLN53),.WL(WL10));
sram_cell_6t_5 inst_cell_10_54 (.BL(BL54),.BLN(BLN54),.WL(WL10));
sram_cell_6t_5 inst_cell_10_55 (.BL(BL55),.BLN(BLN55),.WL(WL10));
sram_cell_6t_5 inst_cell_10_56 (.BL(BL56),.BLN(BLN56),.WL(WL10));
sram_cell_6t_5 inst_cell_10_57 (.BL(BL57),.BLN(BLN57),.WL(WL10));
sram_cell_6t_5 inst_cell_10_58 (.BL(BL58),.BLN(BLN58),.WL(WL10));
sram_cell_6t_5 inst_cell_10_59 (.BL(BL59),.BLN(BLN59),.WL(WL10));
sram_cell_6t_5 inst_cell_10_60 (.BL(BL60),.BLN(BLN60),.WL(WL10));
sram_cell_6t_5 inst_cell_10_61 (.BL(BL61),.BLN(BLN61),.WL(WL10));
sram_cell_6t_5 inst_cell_10_62 (.BL(BL62),.BLN(BLN62),.WL(WL10));
sram_cell_6t_5 inst_cell_10_63 (.BL(BL63),.BLN(BLN63),.WL(WL10));
sram_cell_6t_5 inst_cell_10_64 (.BL(BL64),.BLN(BLN64),.WL(WL10));
sram_cell_6t_5 inst_cell_10_65 (.BL(BL65),.BLN(BLN65),.WL(WL10));
sram_cell_6t_5 inst_cell_10_66 (.BL(BL66),.BLN(BLN66),.WL(WL10));
sram_cell_6t_5 inst_cell_10_67 (.BL(BL67),.BLN(BLN67),.WL(WL10));
sram_cell_6t_5 inst_cell_10_68 (.BL(BL68),.BLN(BLN68),.WL(WL10));
sram_cell_6t_5 inst_cell_10_69 (.BL(BL69),.BLN(BLN69),.WL(WL10));
sram_cell_6t_5 inst_cell_10_70 (.BL(BL70),.BLN(BLN70),.WL(WL10));
sram_cell_6t_5 inst_cell_10_71 (.BL(BL71),.BLN(BLN71),.WL(WL10));
sram_cell_6t_5 inst_cell_10_72 (.BL(BL72),.BLN(BLN72),.WL(WL10));
sram_cell_6t_5 inst_cell_10_73 (.BL(BL73),.BLN(BLN73),.WL(WL10));
sram_cell_6t_5 inst_cell_10_74 (.BL(BL74),.BLN(BLN74),.WL(WL10));
sram_cell_6t_5 inst_cell_10_75 (.BL(BL75),.BLN(BLN75),.WL(WL10));
sram_cell_6t_5 inst_cell_10_76 (.BL(BL76),.BLN(BLN76),.WL(WL10));
sram_cell_6t_5 inst_cell_10_77 (.BL(BL77),.BLN(BLN77),.WL(WL10));
sram_cell_6t_5 inst_cell_10_78 (.BL(BL78),.BLN(BLN78),.WL(WL10));
sram_cell_6t_5 inst_cell_10_79 (.BL(BL79),.BLN(BLN79),.WL(WL10));
sram_cell_6t_5 inst_cell_10_80 (.BL(BL80),.BLN(BLN80),.WL(WL10));
sram_cell_6t_5 inst_cell_10_81 (.BL(BL81),.BLN(BLN81),.WL(WL10));
sram_cell_6t_5 inst_cell_10_82 (.BL(BL82),.BLN(BLN82),.WL(WL10));
sram_cell_6t_5 inst_cell_10_83 (.BL(BL83),.BLN(BLN83),.WL(WL10));
sram_cell_6t_5 inst_cell_10_84 (.BL(BL84),.BLN(BLN84),.WL(WL10));
sram_cell_6t_5 inst_cell_10_85 (.BL(BL85),.BLN(BLN85),.WL(WL10));
sram_cell_6t_5 inst_cell_10_86 (.BL(BL86),.BLN(BLN86),.WL(WL10));
sram_cell_6t_5 inst_cell_10_87 (.BL(BL87),.BLN(BLN87),.WL(WL10));
sram_cell_6t_5 inst_cell_10_88 (.BL(BL88),.BLN(BLN88),.WL(WL10));
sram_cell_6t_5 inst_cell_10_89 (.BL(BL89),.BLN(BLN89),.WL(WL10));
sram_cell_6t_5 inst_cell_10_90 (.BL(BL90),.BLN(BLN90),.WL(WL10));
sram_cell_6t_5 inst_cell_10_91 (.BL(BL91),.BLN(BLN91),.WL(WL10));
sram_cell_6t_5 inst_cell_10_92 (.BL(BL92),.BLN(BLN92),.WL(WL10));
sram_cell_6t_5 inst_cell_10_93 (.BL(BL93),.BLN(BLN93),.WL(WL10));
sram_cell_6t_5 inst_cell_10_94 (.BL(BL94),.BLN(BLN94),.WL(WL10));
sram_cell_6t_5 inst_cell_10_95 (.BL(BL95),.BLN(BLN95),.WL(WL10));
sram_cell_6t_5 inst_cell_10_96 (.BL(BL96),.BLN(BLN96),.WL(WL10));
sram_cell_6t_5 inst_cell_10_97 (.BL(BL97),.BLN(BLN97),.WL(WL10));
sram_cell_6t_5 inst_cell_10_98 (.BL(BL98),.BLN(BLN98),.WL(WL10));
sram_cell_6t_5 inst_cell_10_99 (.BL(BL99),.BLN(BLN99),.WL(WL10));
sram_cell_6t_5 inst_cell_10_100 (.BL(BL100),.BLN(BLN100),.WL(WL10));
sram_cell_6t_5 inst_cell_10_101 (.BL(BL101),.BLN(BLN101),.WL(WL10));
sram_cell_6t_5 inst_cell_10_102 (.BL(BL102),.BLN(BLN102),.WL(WL10));
sram_cell_6t_5 inst_cell_10_103 (.BL(BL103),.BLN(BLN103),.WL(WL10));
sram_cell_6t_5 inst_cell_10_104 (.BL(BL104),.BLN(BLN104),.WL(WL10));
sram_cell_6t_5 inst_cell_10_105 (.BL(BL105),.BLN(BLN105),.WL(WL10));
sram_cell_6t_5 inst_cell_10_106 (.BL(BL106),.BLN(BLN106),.WL(WL10));
sram_cell_6t_5 inst_cell_10_107 (.BL(BL107),.BLN(BLN107),.WL(WL10));
sram_cell_6t_5 inst_cell_10_108 (.BL(BL108),.BLN(BLN108),.WL(WL10));
sram_cell_6t_5 inst_cell_10_109 (.BL(BL109),.BLN(BLN109),.WL(WL10));
sram_cell_6t_5 inst_cell_10_110 (.BL(BL110),.BLN(BLN110),.WL(WL10));
sram_cell_6t_5 inst_cell_10_111 (.BL(BL111),.BLN(BLN111),.WL(WL10));
sram_cell_6t_5 inst_cell_10_112 (.BL(BL112),.BLN(BLN112),.WL(WL10));
sram_cell_6t_5 inst_cell_10_113 (.BL(BL113),.BLN(BLN113),.WL(WL10));
sram_cell_6t_5 inst_cell_10_114 (.BL(BL114),.BLN(BLN114),.WL(WL10));
sram_cell_6t_5 inst_cell_10_115 (.BL(BL115),.BLN(BLN115),.WL(WL10));
sram_cell_6t_5 inst_cell_10_116 (.BL(BL116),.BLN(BLN116),.WL(WL10));
sram_cell_6t_5 inst_cell_10_117 (.BL(BL117),.BLN(BLN117),.WL(WL10));
sram_cell_6t_5 inst_cell_10_118 (.BL(BL118),.BLN(BLN118),.WL(WL10));
sram_cell_6t_5 inst_cell_10_119 (.BL(BL119),.BLN(BLN119),.WL(WL10));
sram_cell_6t_5 inst_cell_10_120 (.BL(BL120),.BLN(BLN120),.WL(WL10));
sram_cell_6t_5 inst_cell_10_121 (.BL(BL121),.BLN(BLN121),.WL(WL10));
sram_cell_6t_5 inst_cell_10_122 (.BL(BL122),.BLN(BLN122),.WL(WL10));
sram_cell_6t_5 inst_cell_10_123 (.BL(BL123),.BLN(BLN123),.WL(WL10));
sram_cell_6t_5 inst_cell_10_124 (.BL(BL124),.BLN(BLN124),.WL(WL10));
sram_cell_6t_5 inst_cell_10_125 (.BL(BL125),.BLN(BLN125),.WL(WL10));
sram_cell_6t_5 inst_cell_10_126 (.BL(BL126),.BLN(BLN126),.WL(WL10));
sram_cell_6t_5 inst_cell_10_127 (.BL(BL127),.BLN(BLN127),.WL(WL10));
sram_cell_6t_5 inst_cell_11_0 (.BL(BL0),.BLN(BLN0),.WL(WL11));
sram_cell_6t_5 inst_cell_11_1 (.BL(BL1),.BLN(BLN1),.WL(WL11));
sram_cell_6t_5 inst_cell_11_2 (.BL(BL2),.BLN(BLN2),.WL(WL11));
sram_cell_6t_5 inst_cell_11_3 (.BL(BL3),.BLN(BLN3),.WL(WL11));
sram_cell_6t_5 inst_cell_11_4 (.BL(BL4),.BLN(BLN4),.WL(WL11));
sram_cell_6t_5 inst_cell_11_5 (.BL(BL5),.BLN(BLN5),.WL(WL11));
sram_cell_6t_5 inst_cell_11_6 (.BL(BL6),.BLN(BLN6),.WL(WL11));
sram_cell_6t_5 inst_cell_11_7 (.BL(BL7),.BLN(BLN7),.WL(WL11));
sram_cell_6t_5 inst_cell_11_8 (.BL(BL8),.BLN(BLN8),.WL(WL11));
sram_cell_6t_5 inst_cell_11_9 (.BL(BL9),.BLN(BLN9),.WL(WL11));
sram_cell_6t_5 inst_cell_11_10 (.BL(BL10),.BLN(BLN10),.WL(WL11));
sram_cell_6t_5 inst_cell_11_11 (.BL(BL11),.BLN(BLN11),.WL(WL11));
sram_cell_6t_5 inst_cell_11_12 (.BL(BL12),.BLN(BLN12),.WL(WL11));
sram_cell_6t_5 inst_cell_11_13 (.BL(BL13),.BLN(BLN13),.WL(WL11));
sram_cell_6t_5 inst_cell_11_14 (.BL(BL14),.BLN(BLN14),.WL(WL11));
sram_cell_6t_5 inst_cell_11_15 (.BL(BL15),.BLN(BLN15),.WL(WL11));
sram_cell_6t_5 inst_cell_11_16 (.BL(BL16),.BLN(BLN16),.WL(WL11));
sram_cell_6t_5 inst_cell_11_17 (.BL(BL17),.BLN(BLN17),.WL(WL11));
sram_cell_6t_5 inst_cell_11_18 (.BL(BL18),.BLN(BLN18),.WL(WL11));
sram_cell_6t_5 inst_cell_11_19 (.BL(BL19),.BLN(BLN19),.WL(WL11));
sram_cell_6t_5 inst_cell_11_20 (.BL(BL20),.BLN(BLN20),.WL(WL11));
sram_cell_6t_5 inst_cell_11_21 (.BL(BL21),.BLN(BLN21),.WL(WL11));
sram_cell_6t_5 inst_cell_11_22 (.BL(BL22),.BLN(BLN22),.WL(WL11));
sram_cell_6t_5 inst_cell_11_23 (.BL(BL23),.BLN(BLN23),.WL(WL11));
sram_cell_6t_5 inst_cell_11_24 (.BL(BL24),.BLN(BLN24),.WL(WL11));
sram_cell_6t_5 inst_cell_11_25 (.BL(BL25),.BLN(BLN25),.WL(WL11));
sram_cell_6t_5 inst_cell_11_26 (.BL(BL26),.BLN(BLN26),.WL(WL11));
sram_cell_6t_5 inst_cell_11_27 (.BL(BL27),.BLN(BLN27),.WL(WL11));
sram_cell_6t_5 inst_cell_11_28 (.BL(BL28),.BLN(BLN28),.WL(WL11));
sram_cell_6t_5 inst_cell_11_29 (.BL(BL29),.BLN(BLN29),.WL(WL11));
sram_cell_6t_5 inst_cell_11_30 (.BL(BL30),.BLN(BLN30),.WL(WL11));
sram_cell_6t_5 inst_cell_11_31 (.BL(BL31),.BLN(BLN31),.WL(WL11));
sram_cell_6t_5 inst_cell_11_32 (.BL(BL32),.BLN(BLN32),.WL(WL11));
sram_cell_6t_5 inst_cell_11_33 (.BL(BL33),.BLN(BLN33),.WL(WL11));
sram_cell_6t_5 inst_cell_11_34 (.BL(BL34),.BLN(BLN34),.WL(WL11));
sram_cell_6t_5 inst_cell_11_35 (.BL(BL35),.BLN(BLN35),.WL(WL11));
sram_cell_6t_5 inst_cell_11_36 (.BL(BL36),.BLN(BLN36),.WL(WL11));
sram_cell_6t_5 inst_cell_11_37 (.BL(BL37),.BLN(BLN37),.WL(WL11));
sram_cell_6t_5 inst_cell_11_38 (.BL(BL38),.BLN(BLN38),.WL(WL11));
sram_cell_6t_5 inst_cell_11_39 (.BL(BL39),.BLN(BLN39),.WL(WL11));
sram_cell_6t_5 inst_cell_11_40 (.BL(BL40),.BLN(BLN40),.WL(WL11));
sram_cell_6t_5 inst_cell_11_41 (.BL(BL41),.BLN(BLN41),.WL(WL11));
sram_cell_6t_5 inst_cell_11_42 (.BL(BL42),.BLN(BLN42),.WL(WL11));
sram_cell_6t_5 inst_cell_11_43 (.BL(BL43),.BLN(BLN43),.WL(WL11));
sram_cell_6t_5 inst_cell_11_44 (.BL(BL44),.BLN(BLN44),.WL(WL11));
sram_cell_6t_5 inst_cell_11_45 (.BL(BL45),.BLN(BLN45),.WL(WL11));
sram_cell_6t_5 inst_cell_11_46 (.BL(BL46),.BLN(BLN46),.WL(WL11));
sram_cell_6t_5 inst_cell_11_47 (.BL(BL47),.BLN(BLN47),.WL(WL11));
sram_cell_6t_5 inst_cell_11_48 (.BL(BL48),.BLN(BLN48),.WL(WL11));
sram_cell_6t_5 inst_cell_11_49 (.BL(BL49),.BLN(BLN49),.WL(WL11));
sram_cell_6t_5 inst_cell_11_50 (.BL(BL50),.BLN(BLN50),.WL(WL11));
sram_cell_6t_5 inst_cell_11_51 (.BL(BL51),.BLN(BLN51),.WL(WL11));
sram_cell_6t_5 inst_cell_11_52 (.BL(BL52),.BLN(BLN52),.WL(WL11));
sram_cell_6t_5 inst_cell_11_53 (.BL(BL53),.BLN(BLN53),.WL(WL11));
sram_cell_6t_5 inst_cell_11_54 (.BL(BL54),.BLN(BLN54),.WL(WL11));
sram_cell_6t_5 inst_cell_11_55 (.BL(BL55),.BLN(BLN55),.WL(WL11));
sram_cell_6t_5 inst_cell_11_56 (.BL(BL56),.BLN(BLN56),.WL(WL11));
sram_cell_6t_5 inst_cell_11_57 (.BL(BL57),.BLN(BLN57),.WL(WL11));
sram_cell_6t_5 inst_cell_11_58 (.BL(BL58),.BLN(BLN58),.WL(WL11));
sram_cell_6t_5 inst_cell_11_59 (.BL(BL59),.BLN(BLN59),.WL(WL11));
sram_cell_6t_5 inst_cell_11_60 (.BL(BL60),.BLN(BLN60),.WL(WL11));
sram_cell_6t_5 inst_cell_11_61 (.BL(BL61),.BLN(BLN61),.WL(WL11));
sram_cell_6t_5 inst_cell_11_62 (.BL(BL62),.BLN(BLN62),.WL(WL11));
sram_cell_6t_5 inst_cell_11_63 (.BL(BL63),.BLN(BLN63),.WL(WL11));
sram_cell_6t_5 inst_cell_11_64 (.BL(BL64),.BLN(BLN64),.WL(WL11));
sram_cell_6t_5 inst_cell_11_65 (.BL(BL65),.BLN(BLN65),.WL(WL11));
sram_cell_6t_5 inst_cell_11_66 (.BL(BL66),.BLN(BLN66),.WL(WL11));
sram_cell_6t_5 inst_cell_11_67 (.BL(BL67),.BLN(BLN67),.WL(WL11));
sram_cell_6t_5 inst_cell_11_68 (.BL(BL68),.BLN(BLN68),.WL(WL11));
sram_cell_6t_5 inst_cell_11_69 (.BL(BL69),.BLN(BLN69),.WL(WL11));
sram_cell_6t_5 inst_cell_11_70 (.BL(BL70),.BLN(BLN70),.WL(WL11));
sram_cell_6t_5 inst_cell_11_71 (.BL(BL71),.BLN(BLN71),.WL(WL11));
sram_cell_6t_5 inst_cell_11_72 (.BL(BL72),.BLN(BLN72),.WL(WL11));
sram_cell_6t_5 inst_cell_11_73 (.BL(BL73),.BLN(BLN73),.WL(WL11));
sram_cell_6t_5 inst_cell_11_74 (.BL(BL74),.BLN(BLN74),.WL(WL11));
sram_cell_6t_5 inst_cell_11_75 (.BL(BL75),.BLN(BLN75),.WL(WL11));
sram_cell_6t_5 inst_cell_11_76 (.BL(BL76),.BLN(BLN76),.WL(WL11));
sram_cell_6t_5 inst_cell_11_77 (.BL(BL77),.BLN(BLN77),.WL(WL11));
sram_cell_6t_5 inst_cell_11_78 (.BL(BL78),.BLN(BLN78),.WL(WL11));
sram_cell_6t_5 inst_cell_11_79 (.BL(BL79),.BLN(BLN79),.WL(WL11));
sram_cell_6t_5 inst_cell_11_80 (.BL(BL80),.BLN(BLN80),.WL(WL11));
sram_cell_6t_5 inst_cell_11_81 (.BL(BL81),.BLN(BLN81),.WL(WL11));
sram_cell_6t_5 inst_cell_11_82 (.BL(BL82),.BLN(BLN82),.WL(WL11));
sram_cell_6t_5 inst_cell_11_83 (.BL(BL83),.BLN(BLN83),.WL(WL11));
sram_cell_6t_5 inst_cell_11_84 (.BL(BL84),.BLN(BLN84),.WL(WL11));
sram_cell_6t_5 inst_cell_11_85 (.BL(BL85),.BLN(BLN85),.WL(WL11));
sram_cell_6t_5 inst_cell_11_86 (.BL(BL86),.BLN(BLN86),.WL(WL11));
sram_cell_6t_5 inst_cell_11_87 (.BL(BL87),.BLN(BLN87),.WL(WL11));
sram_cell_6t_5 inst_cell_11_88 (.BL(BL88),.BLN(BLN88),.WL(WL11));
sram_cell_6t_5 inst_cell_11_89 (.BL(BL89),.BLN(BLN89),.WL(WL11));
sram_cell_6t_5 inst_cell_11_90 (.BL(BL90),.BLN(BLN90),.WL(WL11));
sram_cell_6t_5 inst_cell_11_91 (.BL(BL91),.BLN(BLN91),.WL(WL11));
sram_cell_6t_5 inst_cell_11_92 (.BL(BL92),.BLN(BLN92),.WL(WL11));
sram_cell_6t_5 inst_cell_11_93 (.BL(BL93),.BLN(BLN93),.WL(WL11));
sram_cell_6t_5 inst_cell_11_94 (.BL(BL94),.BLN(BLN94),.WL(WL11));
sram_cell_6t_5 inst_cell_11_95 (.BL(BL95),.BLN(BLN95),.WL(WL11));
sram_cell_6t_5 inst_cell_11_96 (.BL(BL96),.BLN(BLN96),.WL(WL11));
sram_cell_6t_5 inst_cell_11_97 (.BL(BL97),.BLN(BLN97),.WL(WL11));
sram_cell_6t_5 inst_cell_11_98 (.BL(BL98),.BLN(BLN98),.WL(WL11));
sram_cell_6t_5 inst_cell_11_99 (.BL(BL99),.BLN(BLN99),.WL(WL11));
sram_cell_6t_5 inst_cell_11_100 (.BL(BL100),.BLN(BLN100),.WL(WL11));
sram_cell_6t_5 inst_cell_11_101 (.BL(BL101),.BLN(BLN101),.WL(WL11));
sram_cell_6t_5 inst_cell_11_102 (.BL(BL102),.BLN(BLN102),.WL(WL11));
sram_cell_6t_5 inst_cell_11_103 (.BL(BL103),.BLN(BLN103),.WL(WL11));
sram_cell_6t_5 inst_cell_11_104 (.BL(BL104),.BLN(BLN104),.WL(WL11));
sram_cell_6t_5 inst_cell_11_105 (.BL(BL105),.BLN(BLN105),.WL(WL11));
sram_cell_6t_5 inst_cell_11_106 (.BL(BL106),.BLN(BLN106),.WL(WL11));
sram_cell_6t_5 inst_cell_11_107 (.BL(BL107),.BLN(BLN107),.WL(WL11));
sram_cell_6t_5 inst_cell_11_108 (.BL(BL108),.BLN(BLN108),.WL(WL11));
sram_cell_6t_5 inst_cell_11_109 (.BL(BL109),.BLN(BLN109),.WL(WL11));
sram_cell_6t_5 inst_cell_11_110 (.BL(BL110),.BLN(BLN110),.WL(WL11));
sram_cell_6t_5 inst_cell_11_111 (.BL(BL111),.BLN(BLN111),.WL(WL11));
sram_cell_6t_5 inst_cell_11_112 (.BL(BL112),.BLN(BLN112),.WL(WL11));
sram_cell_6t_5 inst_cell_11_113 (.BL(BL113),.BLN(BLN113),.WL(WL11));
sram_cell_6t_5 inst_cell_11_114 (.BL(BL114),.BLN(BLN114),.WL(WL11));
sram_cell_6t_5 inst_cell_11_115 (.BL(BL115),.BLN(BLN115),.WL(WL11));
sram_cell_6t_5 inst_cell_11_116 (.BL(BL116),.BLN(BLN116),.WL(WL11));
sram_cell_6t_5 inst_cell_11_117 (.BL(BL117),.BLN(BLN117),.WL(WL11));
sram_cell_6t_5 inst_cell_11_118 (.BL(BL118),.BLN(BLN118),.WL(WL11));
sram_cell_6t_5 inst_cell_11_119 (.BL(BL119),.BLN(BLN119),.WL(WL11));
sram_cell_6t_5 inst_cell_11_120 (.BL(BL120),.BLN(BLN120),.WL(WL11));
sram_cell_6t_5 inst_cell_11_121 (.BL(BL121),.BLN(BLN121),.WL(WL11));
sram_cell_6t_5 inst_cell_11_122 (.BL(BL122),.BLN(BLN122),.WL(WL11));
sram_cell_6t_5 inst_cell_11_123 (.BL(BL123),.BLN(BLN123),.WL(WL11));
sram_cell_6t_5 inst_cell_11_124 (.BL(BL124),.BLN(BLN124),.WL(WL11));
sram_cell_6t_5 inst_cell_11_125 (.BL(BL125),.BLN(BLN125),.WL(WL11));
sram_cell_6t_5 inst_cell_11_126 (.BL(BL126),.BLN(BLN126),.WL(WL11));
sram_cell_6t_5 inst_cell_11_127 (.BL(BL127),.BLN(BLN127),.WL(WL11));
sram_cell_6t_5 inst_cell_12_0 (.BL(BL0),.BLN(BLN0),.WL(WL12));
sram_cell_6t_5 inst_cell_12_1 (.BL(BL1),.BLN(BLN1),.WL(WL12));
sram_cell_6t_5 inst_cell_12_2 (.BL(BL2),.BLN(BLN2),.WL(WL12));
sram_cell_6t_5 inst_cell_12_3 (.BL(BL3),.BLN(BLN3),.WL(WL12));
sram_cell_6t_5 inst_cell_12_4 (.BL(BL4),.BLN(BLN4),.WL(WL12));
sram_cell_6t_5 inst_cell_12_5 (.BL(BL5),.BLN(BLN5),.WL(WL12));
sram_cell_6t_5 inst_cell_12_6 (.BL(BL6),.BLN(BLN6),.WL(WL12));
sram_cell_6t_5 inst_cell_12_7 (.BL(BL7),.BLN(BLN7),.WL(WL12));
sram_cell_6t_5 inst_cell_12_8 (.BL(BL8),.BLN(BLN8),.WL(WL12));
sram_cell_6t_5 inst_cell_12_9 (.BL(BL9),.BLN(BLN9),.WL(WL12));
sram_cell_6t_5 inst_cell_12_10 (.BL(BL10),.BLN(BLN10),.WL(WL12));
sram_cell_6t_5 inst_cell_12_11 (.BL(BL11),.BLN(BLN11),.WL(WL12));
sram_cell_6t_5 inst_cell_12_12 (.BL(BL12),.BLN(BLN12),.WL(WL12));
sram_cell_6t_5 inst_cell_12_13 (.BL(BL13),.BLN(BLN13),.WL(WL12));
sram_cell_6t_5 inst_cell_12_14 (.BL(BL14),.BLN(BLN14),.WL(WL12));
sram_cell_6t_5 inst_cell_12_15 (.BL(BL15),.BLN(BLN15),.WL(WL12));
sram_cell_6t_5 inst_cell_12_16 (.BL(BL16),.BLN(BLN16),.WL(WL12));
sram_cell_6t_5 inst_cell_12_17 (.BL(BL17),.BLN(BLN17),.WL(WL12));
sram_cell_6t_5 inst_cell_12_18 (.BL(BL18),.BLN(BLN18),.WL(WL12));
sram_cell_6t_5 inst_cell_12_19 (.BL(BL19),.BLN(BLN19),.WL(WL12));
sram_cell_6t_5 inst_cell_12_20 (.BL(BL20),.BLN(BLN20),.WL(WL12));
sram_cell_6t_5 inst_cell_12_21 (.BL(BL21),.BLN(BLN21),.WL(WL12));
sram_cell_6t_5 inst_cell_12_22 (.BL(BL22),.BLN(BLN22),.WL(WL12));
sram_cell_6t_5 inst_cell_12_23 (.BL(BL23),.BLN(BLN23),.WL(WL12));
sram_cell_6t_5 inst_cell_12_24 (.BL(BL24),.BLN(BLN24),.WL(WL12));
sram_cell_6t_5 inst_cell_12_25 (.BL(BL25),.BLN(BLN25),.WL(WL12));
sram_cell_6t_5 inst_cell_12_26 (.BL(BL26),.BLN(BLN26),.WL(WL12));
sram_cell_6t_5 inst_cell_12_27 (.BL(BL27),.BLN(BLN27),.WL(WL12));
sram_cell_6t_5 inst_cell_12_28 (.BL(BL28),.BLN(BLN28),.WL(WL12));
sram_cell_6t_5 inst_cell_12_29 (.BL(BL29),.BLN(BLN29),.WL(WL12));
sram_cell_6t_5 inst_cell_12_30 (.BL(BL30),.BLN(BLN30),.WL(WL12));
sram_cell_6t_5 inst_cell_12_31 (.BL(BL31),.BLN(BLN31),.WL(WL12));
sram_cell_6t_5 inst_cell_12_32 (.BL(BL32),.BLN(BLN32),.WL(WL12));
sram_cell_6t_5 inst_cell_12_33 (.BL(BL33),.BLN(BLN33),.WL(WL12));
sram_cell_6t_5 inst_cell_12_34 (.BL(BL34),.BLN(BLN34),.WL(WL12));
sram_cell_6t_5 inst_cell_12_35 (.BL(BL35),.BLN(BLN35),.WL(WL12));
sram_cell_6t_5 inst_cell_12_36 (.BL(BL36),.BLN(BLN36),.WL(WL12));
sram_cell_6t_5 inst_cell_12_37 (.BL(BL37),.BLN(BLN37),.WL(WL12));
sram_cell_6t_5 inst_cell_12_38 (.BL(BL38),.BLN(BLN38),.WL(WL12));
sram_cell_6t_5 inst_cell_12_39 (.BL(BL39),.BLN(BLN39),.WL(WL12));
sram_cell_6t_5 inst_cell_12_40 (.BL(BL40),.BLN(BLN40),.WL(WL12));
sram_cell_6t_5 inst_cell_12_41 (.BL(BL41),.BLN(BLN41),.WL(WL12));
sram_cell_6t_5 inst_cell_12_42 (.BL(BL42),.BLN(BLN42),.WL(WL12));
sram_cell_6t_5 inst_cell_12_43 (.BL(BL43),.BLN(BLN43),.WL(WL12));
sram_cell_6t_5 inst_cell_12_44 (.BL(BL44),.BLN(BLN44),.WL(WL12));
sram_cell_6t_5 inst_cell_12_45 (.BL(BL45),.BLN(BLN45),.WL(WL12));
sram_cell_6t_5 inst_cell_12_46 (.BL(BL46),.BLN(BLN46),.WL(WL12));
sram_cell_6t_5 inst_cell_12_47 (.BL(BL47),.BLN(BLN47),.WL(WL12));
sram_cell_6t_5 inst_cell_12_48 (.BL(BL48),.BLN(BLN48),.WL(WL12));
sram_cell_6t_5 inst_cell_12_49 (.BL(BL49),.BLN(BLN49),.WL(WL12));
sram_cell_6t_5 inst_cell_12_50 (.BL(BL50),.BLN(BLN50),.WL(WL12));
sram_cell_6t_5 inst_cell_12_51 (.BL(BL51),.BLN(BLN51),.WL(WL12));
sram_cell_6t_5 inst_cell_12_52 (.BL(BL52),.BLN(BLN52),.WL(WL12));
sram_cell_6t_5 inst_cell_12_53 (.BL(BL53),.BLN(BLN53),.WL(WL12));
sram_cell_6t_5 inst_cell_12_54 (.BL(BL54),.BLN(BLN54),.WL(WL12));
sram_cell_6t_5 inst_cell_12_55 (.BL(BL55),.BLN(BLN55),.WL(WL12));
sram_cell_6t_5 inst_cell_12_56 (.BL(BL56),.BLN(BLN56),.WL(WL12));
sram_cell_6t_5 inst_cell_12_57 (.BL(BL57),.BLN(BLN57),.WL(WL12));
sram_cell_6t_5 inst_cell_12_58 (.BL(BL58),.BLN(BLN58),.WL(WL12));
sram_cell_6t_5 inst_cell_12_59 (.BL(BL59),.BLN(BLN59),.WL(WL12));
sram_cell_6t_5 inst_cell_12_60 (.BL(BL60),.BLN(BLN60),.WL(WL12));
sram_cell_6t_5 inst_cell_12_61 (.BL(BL61),.BLN(BLN61),.WL(WL12));
sram_cell_6t_5 inst_cell_12_62 (.BL(BL62),.BLN(BLN62),.WL(WL12));
sram_cell_6t_5 inst_cell_12_63 (.BL(BL63),.BLN(BLN63),.WL(WL12));
sram_cell_6t_5 inst_cell_12_64 (.BL(BL64),.BLN(BLN64),.WL(WL12));
sram_cell_6t_5 inst_cell_12_65 (.BL(BL65),.BLN(BLN65),.WL(WL12));
sram_cell_6t_5 inst_cell_12_66 (.BL(BL66),.BLN(BLN66),.WL(WL12));
sram_cell_6t_5 inst_cell_12_67 (.BL(BL67),.BLN(BLN67),.WL(WL12));
sram_cell_6t_5 inst_cell_12_68 (.BL(BL68),.BLN(BLN68),.WL(WL12));
sram_cell_6t_5 inst_cell_12_69 (.BL(BL69),.BLN(BLN69),.WL(WL12));
sram_cell_6t_5 inst_cell_12_70 (.BL(BL70),.BLN(BLN70),.WL(WL12));
sram_cell_6t_5 inst_cell_12_71 (.BL(BL71),.BLN(BLN71),.WL(WL12));
sram_cell_6t_5 inst_cell_12_72 (.BL(BL72),.BLN(BLN72),.WL(WL12));
sram_cell_6t_5 inst_cell_12_73 (.BL(BL73),.BLN(BLN73),.WL(WL12));
sram_cell_6t_5 inst_cell_12_74 (.BL(BL74),.BLN(BLN74),.WL(WL12));
sram_cell_6t_5 inst_cell_12_75 (.BL(BL75),.BLN(BLN75),.WL(WL12));
sram_cell_6t_5 inst_cell_12_76 (.BL(BL76),.BLN(BLN76),.WL(WL12));
sram_cell_6t_5 inst_cell_12_77 (.BL(BL77),.BLN(BLN77),.WL(WL12));
sram_cell_6t_5 inst_cell_12_78 (.BL(BL78),.BLN(BLN78),.WL(WL12));
sram_cell_6t_5 inst_cell_12_79 (.BL(BL79),.BLN(BLN79),.WL(WL12));
sram_cell_6t_5 inst_cell_12_80 (.BL(BL80),.BLN(BLN80),.WL(WL12));
sram_cell_6t_5 inst_cell_12_81 (.BL(BL81),.BLN(BLN81),.WL(WL12));
sram_cell_6t_5 inst_cell_12_82 (.BL(BL82),.BLN(BLN82),.WL(WL12));
sram_cell_6t_5 inst_cell_12_83 (.BL(BL83),.BLN(BLN83),.WL(WL12));
sram_cell_6t_5 inst_cell_12_84 (.BL(BL84),.BLN(BLN84),.WL(WL12));
sram_cell_6t_5 inst_cell_12_85 (.BL(BL85),.BLN(BLN85),.WL(WL12));
sram_cell_6t_5 inst_cell_12_86 (.BL(BL86),.BLN(BLN86),.WL(WL12));
sram_cell_6t_5 inst_cell_12_87 (.BL(BL87),.BLN(BLN87),.WL(WL12));
sram_cell_6t_5 inst_cell_12_88 (.BL(BL88),.BLN(BLN88),.WL(WL12));
sram_cell_6t_5 inst_cell_12_89 (.BL(BL89),.BLN(BLN89),.WL(WL12));
sram_cell_6t_5 inst_cell_12_90 (.BL(BL90),.BLN(BLN90),.WL(WL12));
sram_cell_6t_5 inst_cell_12_91 (.BL(BL91),.BLN(BLN91),.WL(WL12));
sram_cell_6t_5 inst_cell_12_92 (.BL(BL92),.BLN(BLN92),.WL(WL12));
sram_cell_6t_5 inst_cell_12_93 (.BL(BL93),.BLN(BLN93),.WL(WL12));
sram_cell_6t_5 inst_cell_12_94 (.BL(BL94),.BLN(BLN94),.WL(WL12));
sram_cell_6t_5 inst_cell_12_95 (.BL(BL95),.BLN(BLN95),.WL(WL12));
sram_cell_6t_5 inst_cell_12_96 (.BL(BL96),.BLN(BLN96),.WL(WL12));
sram_cell_6t_5 inst_cell_12_97 (.BL(BL97),.BLN(BLN97),.WL(WL12));
sram_cell_6t_5 inst_cell_12_98 (.BL(BL98),.BLN(BLN98),.WL(WL12));
sram_cell_6t_5 inst_cell_12_99 (.BL(BL99),.BLN(BLN99),.WL(WL12));
sram_cell_6t_5 inst_cell_12_100 (.BL(BL100),.BLN(BLN100),.WL(WL12));
sram_cell_6t_5 inst_cell_12_101 (.BL(BL101),.BLN(BLN101),.WL(WL12));
sram_cell_6t_5 inst_cell_12_102 (.BL(BL102),.BLN(BLN102),.WL(WL12));
sram_cell_6t_5 inst_cell_12_103 (.BL(BL103),.BLN(BLN103),.WL(WL12));
sram_cell_6t_5 inst_cell_12_104 (.BL(BL104),.BLN(BLN104),.WL(WL12));
sram_cell_6t_5 inst_cell_12_105 (.BL(BL105),.BLN(BLN105),.WL(WL12));
sram_cell_6t_5 inst_cell_12_106 (.BL(BL106),.BLN(BLN106),.WL(WL12));
sram_cell_6t_5 inst_cell_12_107 (.BL(BL107),.BLN(BLN107),.WL(WL12));
sram_cell_6t_5 inst_cell_12_108 (.BL(BL108),.BLN(BLN108),.WL(WL12));
sram_cell_6t_5 inst_cell_12_109 (.BL(BL109),.BLN(BLN109),.WL(WL12));
sram_cell_6t_5 inst_cell_12_110 (.BL(BL110),.BLN(BLN110),.WL(WL12));
sram_cell_6t_5 inst_cell_12_111 (.BL(BL111),.BLN(BLN111),.WL(WL12));
sram_cell_6t_5 inst_cell_12_112 (.BL(BL112),.BLN(BLN112),.WL(WL12));
sram_cell_6t_5 inst_cell_12_113 (.BL(BL113),.BLN(BLN113),.WL(WL12));
sram_cell_6t_5 inst_cell_12_114 (.BL(BL114),.BLN(BLN114),.WL(WL12));
sram_cell_6t_5 inst_cell_12_115 (.BL(BL115),.BLN(BLN115),.WL(WL12));
sram_cell_6t_5 inst_cell_12_116 (.BL(BL116),.BLN(BLN116),.WL(WL12));
sram_cell_6t_5 inst_cell_12_117 (.BL(BL117),.BLN(BLN117),.WL(WL12));
sram_cell_6t_5 inst_cell_12_118 (.BL(BL118),.BLN(BLN118),.WL(WL12));
sram_cell_6t_5 inst_cell_12_119 (.BL(BL119),.BLN(BLN119),.WL(WL12));
sram_cell_6t_5 inst_cell_12_120 (.BL(BL120),.BLN(BLN120),.WL(WL12));
sram_cell_6t_5 inst_cell_12_121 (.BL(BL121),.BLN(BLN121),.WL(WL12));
sram_cell_6t_5 inst_cell_12_122 (.BL(BL122),.BLN(BLN122),.WL(WL12));
sram_cell_6t_5 inst_cell_12_123 (.BL(BL123),.BLN(BLN123),.WL(WL12));
sram_cell_6t_5 inst_cell_12_124 (.BL(BL124),.BLN(BLN124),.WL(WL12));
sram_cell_6t_5 inst_cell_12_125 (.BL(BL125),.BLN(BLN125),.WL(WL12));
sram_cell_6t_5 inst_cell_12_126 (.BL(BL126),.BLN(BLN126),.WL(WL12));
sram_cell_6t_5 inst_cell_12_127 (.BL(BL127),.BLN(BLN127),.WL(WL12));
sram_cell_6t_5 inst_cell_13_0 (.BL(BL0),.BLN(BLN0),.WL(WL13));
sram_cell_6t_5 inst_cell_13_1 (.BL(BL1),.BLN(BLN1),.WL(WL13));
sram_cell_6t_5 inst_cell_13_2 (.BL(BL2),.BLN(BLN2),.WL(WL13));
sram_cell_6t_5 inst_cell_13_3 (.BL(BL3),.BLN(BLN3),.WL(WL13));
sram_cell_6t_5 inst_cell_13_4 (.BL(BL4),.BLN(BLN4),.WL(WL13));
sram_cell_6t_5 inst_cell_13_5 (.BL(BL5),.BLN(BLN5),.WL(WL13));
sram_cell_6t_5 inst_cell_13_6 (.BL(BL6),.BLN(BLN6),.WL(WL13));
sram_cell_6t_5 inst_cell_13_7 (.BL(BL7),.BLN(BLN7),.WL(WL13));
sram_cell_6t_5 inst_cell_13_8 (.BL(BL8),.BLN(BLN8),.WL(WL13));
sram_cell_6t_5 inst_cell_13_9 (.BL(BL9),.BLN(BLN9),.WL(WL13));
sram_cell_6t_5 inst_cell_13_10 (.BL(BL10),.BLN(BLN10),.WL(WL13));
sram_cell_6t_5 inst_cell_13_11 (.BL(BL11),.BLN(BLN11),.WL(WL13));
sram_cell_6t_5 inst_cell_13_12 (.BL(BL12),.BLN(BLN12),.WL(WL13));
sram_cell_6t_5 inst_cell_13_13 (.BL(BL13),.BLN(BLN13),.WL(WL13));
sram_cell_6t_5 inst_cell_13_14 (.BL(BL14),.BLN(BLN14),.WL(WL13));
sram_cell_6t_5 inst_cell_13_15 (.BL(BL15),.BLN(BLN15),.WL(WL13));
sram_cell_6t_5 inst_cell_13_16 (.BL(BL16),.BLN(BLN16),.WL(WL13));
sram_cell_6t_5 inst_cell_13_17 (.BL(BL17),.BLN(BLN17),.WL(WL13));
sram_cell_6t_5 inst_cell_13_18 (.BL(BL18),.BLN(BLN18),.WL(WL13));
sram_cell_6t_5 inst_cell_13_19 (.BL(BL19),.BLN(BLN19),.WL(WL13));
sram_cell_6t_5 inst_cell_13_20 (.BL(BL20),.BLN(BLN20),.WL(WL13));
sram_cell_6t_5 inst_cell_13_21 (.BL(BL21),.BLN(BLN21),.WL(WL13));
sram_cell_6t_5 inst_cell_13_22 (.BL(BL22),.BLN(BLN22),.WL(WL13));
sram_cell_6t_5 inst_cell_13_23 (.BL(BL23),.BLN(BLN23),.WL(WL13));
sram_cell_6t_5 inst_cell_13_24 (.BL(BL24),.BLN(BLN24),.WL(WL13));
sram_cell_6t_5 inst_cell_13_25 (.BL(BL25),.BLN(BLN25),.WL(WL13));
sram_cell_6t_5 inst_cell_13_26 (.BL(BL26),.BLN(BLN26),.WL(WL13));
sram_cell_6t_5 inst_cell_13_27 (.BL(BL27),.BLN(BLN27),.WL(WL13));
sram_cell_6t_5 inst_cell_13_28 (.BL(BL28),.BLN(BLN28),.WL(WL13));
sram_cell_6t_5 inst_cell_13_29 (.BL(BL29),.BLN(BLN29),.WL(WL13));
sram_cell_6t_5 inst_cell_13_30 (.BL(BL30),.BLN(BLN30),.WL(WL13));
sram_cell_6t_5 inst_cell_13_31 (.BL(BL31),.BLN(BLN31),.WL(WL13));
sram_cell_6t_5 inst_cell_13_32 (.BL(BL32),.BLN(BLN32),.WL(WL13));
sram_cell_6t_5 inst_cell_13_33 (.BL(BL33),.BLN(BLN33),.WL(WL13));
sram_cell_6t_5 inst_cell_13_34 (.BL(BL34),.BLN(BLN34),.WL(WL13));
sram_cell_6t_5 inst_cell_13_35 (.BL(BL35),.BLN(BLN35),.WL(WL13));
sram_cell_6t_5 inst_cell_13_36 (.BL(BL36),.BLN(BLN36),.WL(WL13));
sram_cell_6t_5 inst_cell_13_37 (.BL(BL37),.BLN(BLN37),.WL(WL13));
sram_cell_6t_5 inst_cell_13_38 (.BL(BL38),.BLN(BLN38),.WL(WL13));
sram_cell_6t_5 inst_cell_13_39 (.BL(BL39),.BLN(BLN39),.WL(WL13));
sram_cell_6t_5 inst_cell_13_40 (.BL(BL40),.BLN(BLN40),.WL(WL13));
sram_cell_6t_5 inst_cell_13_41 (.BL(BL41),.BLN(BLN41),.WL(WL13));
sram_cell_6t_5 inst_cell_13_42 (.BL(BL42),.BLN(BLN42),.WL(WL13));
sram_cell_6t_5 inst_cell_13_43 (.BL(BL43),.BLN(BLN43),.WL(WL13));
sram_cell_6t_5 inst_cell_13_44 (.BL(BL44),.BLN(BLN44),.WL(WL13));
sram_cell_6t_5 inst_cell_13_45 (.BL(BL45),.BLN(BLN45),.WL(WL13));
sram_cell_6t_5 inst_cell_13_46 (.BL(BL46),.BLN(BLN46),.WL(WL13));
sram_cell_6t_5 inst_cell_13_47 (.BL(BL47),.BLN(BLN47),.WL(WL13));
sram_cell_6t_5 inst_cell_13_48 (.BL(BL48),.BLN(BLN48),.WL(WL13));
sram_cell_6t_5 inst_cell_13_49 (.BL(BL49),.BLN(BLN49),.WL(WL13));
sram_cell_6t_5 inst_cell_13_50 (.BL(BL50),.BLN(BLN50),.WL(WL13));
sram_cell_6t_5 inst_cell_13_51 (.BL(BL51),.BLN(BLN51),.WL(WL13));
sram_cell_6t_5 inst_cell_13_52 (.BL(BL52),.BLN(BLN52),.WL(WL13));
sram_cell_6t_5 inst_cell_13_53 (.BL(BL53),.BLN(BLN53),.WL(WL13));
sram_cell_6t_5 inst_cell_13_54 (.BL(BL54),.BLN(BLN54),.WL(WL13));
sram_cell_6t_5 inst_cell_13_55 (.BL(BL55),.BLN(BLN55),.WL(WL13));
sram_cell_6t_5 inst_cell_13_56 (.BL(BL56),.BLN(BLN56),.WL(WL13));
sram_cell_6t_5 inst_cell_13_57 (.BL(BL57),.BLN(BLN57),.WL(WL13));
sram_cell_6t_5 inst_cell_13_58 (.BL(BL58),.BLN(BLN58),.WL(WL13));
sram_cell_6t_5 inst_cell_13_59 (.BL(BL59),.BLN(BLN59),.WL(WL13));
sram_cell_6t_5 inst_cell_13_60 (.BL(BL60),.BLN(BLN60),.WL(WL13));
sram_cell_6t_5 inst_cell_13_61 (.BL(BL61),.BLN(BLN61),.WL(WL13));
sram_cell_6t_5 inst_cell_13_62 (.BL(BL62),.BLN(BLN62),.WL(WL13));
sram_cell_6t_5 inst_cell_13_63 (.BL(BL63),.BLN(BLN63),.WL(WL13));
sram_cell_6t_5 inst_cell_13_64 (.BL(BL64),.BLN(BLN64),.WL(WL13));
sram_cell_6t_5 inst_cell_13_65 (.BL(BL65),.BLN(BLN65),.WL(WL13));
sram_cell_6t_5 inst_cell_13_66 (.BL(BL66),.BLN(BLN66),.WL(WL13));
sram_cell_6t_5 inst_cell_13_67 (.BL(BL67),.BLN(BLN67),.WL(WL13));
sram_cell_6t_5 inst_cell_13_68 (.BL(BL68),.BLN(BLN68),.WL(WL13));
sram_cell_6t_5 inst_cell_13_69 (.BL(BL69),.BLN(BLN69),.WL(WL13));
sram_cell_6t_5 inst_cell_13_70 (.BL(BL70),.BLN(BLN70),.WL(WL13));
sram_cell_6t_5 inst_cell_13_71 (.BL(BL71),.BLN(BLN71),.WL(WL13));
sram_cell_6t_5 inst_cell_13_72 (.BL(BL72),.BLN(BLN72),.WL(WL13));
sram_cell_6t_5 inst_cell_13_73 (.BL(BL73),.BLN(BLN73),.WL(WL13));
sram_cell_6t_5 inst_cell_13_74 (.BL(BL74),.BLN(BLN74),.WL(WL13));
sram_cell_6t_5 inst_cell_13_75 (.BL(BL75),.BLN(BLN75),.WL(WL13));
sram_cell_6t_5 inst_cell_13_76 (.BL(BL76),.BLN(BLN76),.WL(WL13));
sram_cell_6t_5 inst_cell_13_77 (.BL(BL77),.BLN(BLN77),.WL(WL13));
sram_cell_6t_5 inst_cell_13_78 (.BL(BL78),.BLN(BLN78),.WL(WL13));
sram_cell_6t_5 inst_cell_13_79 (.BL(BL79),.BLN(BLN79),.WL(WL13));
sram_cell_6t_5 inst_cell_13_80 (.BL(BL80),.BLN(BLN80),.WL(WL13));
sram_cell_6t_5 inst_cell_13_81 (.BL(BL81),.BLN(BLN81),.WL(WL13));
sram_cell_6t_5 inst_cell_13_82 (.BL(BL82),.BLN(BLN82),.WL(WL13));
sram_cell_6t_5 inst_cell_13_83 (.BL(BL83),.BLN(BLN83),.WL(WL13));
sram_cell_6t_5 inst_cell_13_84 (.BL(BL84),.BLN(BLN84),.WL(WL13));
sram_cell_6t_5 inst_cell_13_85 (.BL(BL85),.BLN(BLN85),.WL(WL13));
sram_cell_6t_5 inst_cell_13_86 (.BL(BL86),.BLN(BLN86),.WL(WL13));
sram_cell_6t_5 inst_cell_13_87 (.BL(BL87),.BLN(BLN87),.WL(WL13));
sram_cell_6t_5 inst_cell_13_88 (.BL(BL88),.BLN(BLN88),.WL(WL13));
sram_cell_6t_5 inst_cell_13_89 (.BL(BL89),.BLN(BLN89),.WL(WL13));
sram_cell_6t_5 inst_cell_13_90 (.BL(BL90),.BLN(BLN90),.WL(WL13));
sram_cell_6t_5 inst_cell_13_91 (.BL(BL91),.BLN(BLN91),.WL(WL13));
sram_cell_6t_5 inst_cell_13_92 (.BL(BL92),.BLN(BLN92),.WL(WL13));
sram_cell_6t_5 inst_cell_13_93 (.BL(BL93),.BLN(BLN93),.WL(WL13));
sram_cell_6t_5 inst_cell_13_94 (.BL(BL94),.BLN(BLN94),.WL(WL13));
sram_cell_6t_5 inst_cell_13_95 (.BL(BL95),.BLN(BLN95),.WL(WL13));
sram_cell_6t_5 inst_cell_13_96 (.BL(BL96),.BLN(BLN96),.WL(WL13));
sram_cell_6t_5 inst_cell_13_97 (.BL(BL97),.BLN(BLN97),.WL(WL13));
sram_cell_6t_5 inst_cell_13_98 (.BL(BL98),.BLN(BLN98),.WL(WL13));
sram_cell_6t_5 inst_cell_13_99 (.BL(BL99),.BLN(BLN99),.WL(WL13));
sram_cell_6t_5 inst_cell_13_100 (.BL(BL100),.BLN(BLN100),.WL(WL13));
sram_cell_6t_5 inst_cell_13_101 (.BL(BL101),.BLN(BLN101),.WL(WL13));
sram_cell_6t_5 inst_cell_13_102 (.BL(BL102),.BLN(BLN102),.WL(WL13));
sram_cell_6t_5 inst_cell_13_103 (.BL(BL103),.BLN(BLN103),.WL(WL13));
sram_cell_6t_5 inst_cell_13_104 (.BL(BL104),.BLN(BLN104),.WL(WL13));
sram_cell_6t_5 inst_cell_13_105 (.BL(BL105),.BLN(BLN105),.WL(WL13));
sram_cell_6t_5 inst_cell_13_106 (.BL(BL106),.BLN(BLN106),.WL(WL13));
sram_cell_6t_5 inst_cell_13_107 (.BL(BL107),.BLN(BLN107),.WL(WL13));
sram_cell_6t_5 inst_cell_13_108 (.BL(BL108),.BLN(BLN108),.WL(WL13));
sram_cell_6t_5 inst_cell_13_109 (.BL(BL109),.BLN(BLN109),.WL(WL13));
sram_cell_6t_5 inst_cell_13_110 (.BL(BL110),.BLN(BLN110),.WL(WL13));
sram_cell_6t_5 inst_cell_13_111 (.BL(BL111),.BLN(BLN111),.WL(WL13));
sram_cell_6t_5 inst_cell_13_112 (.BL(BL112),.BLN(BLN112),.WL(WL13));
sram_cell_6t_5 inst_cell_13_113 (.BL(BL113),.BLN(BLN113),.WL(WL13));
sram_cell_6t_5 inst_cell_13_114 (.BL(BL114),.BLN(BLN114),.WL(WL13));
sram_cell_6t_5 inst_cell_13_115 (.BL(BL115),.BLN(BLN115),.WL(WL13));
sram_cell_6t_5 inst_cell_13_116 (.BL(BL116),.BLN(BLN116),.WL(WL13));
sram_cell_6t_5 inst_cell_13_117 (.BL(BL117),.BLN(BLN117),.WL(WL13));
sram_cell_6t_5 inst_cell_13_118 (.BL(BL118),.BLN(BLN118),.WL(WL13));
sram_cell_6t_5 inst_cell_13_119 (.BL(BL119),.BLN(BLN119),.WL(WL13));
sram_cell_6t_5 inst_cell_13_120 (.BL(BL120),.BLN(BLN120),.WL(WL13));
sram_cell_6t_5 inst_cell_13_121 (.BL(BL121),.BLN(BLN121),.WL(WL13));
sram_cell_6t_5 inst_cell_13_122 (.BL(BL122),.BLN(BLN122),.WL(WL13));
sram_cell_6t_5 inst_cell_13_123 (.BL(BL123),.BLN(BLN123),.WL(WL13));
sram_cell_6t_5 inst_cell_13_124 (.BL(BL124),.BLN(BLN124),.WL(WL13));
sram_cell_6t_5 inst_cell_13_125 (.BL(BL125),.BLN(BLN125),.WL(WL13));
sram_cell_6t_5 inst_cell_13_126 (.BL(BL126),.BLN(BLN126),.WL(WL13));
sram_cell_6t_5 inst_cell_13_127 (.BL(BL127),.BLN(BLN127),.WL(WL13));
sram_cell_6t_5 inst_cell_14_0 (.BL(BL0),.BLN(BLN0),.WL(WL14));
sram_cell_6t_5 inst_cell_14_1 (.BL(BL1),.BLN(BLN1),.WL(WL14));
sram_cell_6t_5 inst_cell_14_2 (.BL(BL2),.BLN(BLN2),.WL(WL14));
sram_cell_6t_5 inst_cell_14_3 (.BL(BL3),.BLN(BLN3),.WL(WL14));
sram_cell_6t_5 inst_cell_14_4 (.BL(BL4),.BLN(BLN4),.WL(WL14));
sram_cell_6t_5 inst_cell_14_5 (.BL(BL5),.BLN(BLN5),.WL(WL14));
sram_cell_6t_5 inst_cell_14_6 (.BL(BL6),.BLN(BLN6),.WL(WL14));
sram_cell_6t_5 inst_cell_14_7 (.BL(BL7),.BLN(BLN7),.WL(WL14));
sram_cell_6t_5 inst_cell_14_8 (.BL(BL8),.BLN(BLN8),.WL(WL14));
sram_cell_6t_5 inst_cell_14_9 (.BL(BL9),.BLN(BLN9),.WL(WL14));
sram_cell_6t_5 inst_cell_14_10 (.BL(BL10),.BLN(BLN10),.WL(WL14));
sram_cell_6t_5 inst_cell_14_11 (.BL(BL11),.BLN(BLN11),.WL(WL14));
sram_cell_6t_5 inst_cell_14_12 (.BL(BL12),.BLN(BLN12),.WL(WL14));
sram_cell_6t_5 inst_cell_14_13 (.BL(BL13),.BLN(BLN13),.WL(WL14));
sram_cell_6t_5 inst_cell_14_14 (.BL(BL14),.BLN(BLN14),.WL(WL14));
sram_cell_6t_5 inst_cell_14_15 (.BL(BL15),.BLN(BLN15),.WL(WL14));
sram_cell_6t_5 inst_cell_14_16 (.BL(BL16),.BLN(BLN16),.WL(WL14));
sram_cell_6t_5 inst_cell_14_17 (.BL(BL17),.BLN(BLN17),.WL(WL14));
sram_cell_6t_5 inst_cell_14_18 (.BL(BL18),.BLN(BLN18),.WL(WL14));
sram_cell_6t_5 inst_cell_14_19 (.BL(BL19),.BLN(BLN19),.WL(WL14));
sram_cell_6t_5 inst_cell_14_20 (.BL(BL20),.BLN(BLN20),.WL(WL14));
sram_cell_6t_5 inst_cell_14_21 (.BL(BL21),.BLN(BLN21),.WL(WL14));
sram_cell_6t_5 inst_cell_14_22 (.BL(BL22),.BLN(BLN22),.WL(WL14));
sram_cell_6t_5 inst_cell_14_23 (.BL(BL23),.BLN(BLN23),.WL(WL14));
sram_cell_6t_5 inst_cell_14_24 (.BL(BL24),.BLN(BLN24),.WL(WL14));
sram_cell_6t_5 inst_cell_14_25 (.BL(BL25),.BLN(BLN25),.WL(WL14));
sram_cell_6t_5 inst_cell_14_26 (.BL(BL26),.BLN(BLN26),.WL(WL14));
sram_cell_6t_5 inst_cell_14_27 (.BL(BL27),.BLN(BLN27),.WL(WL14));
sram_cell_6t_5 inst_cell_14_28 (.BL(BL28),.BLN(BLN28),.WL(WL14));
sram_cell_6t_5 inst_cell_14_29 (.BL(BL29),.BLN(BLN29),.WL(WL14));
sram_cell_6t_5 inst_cell_14_30 (.BL(BL30),.BLN(BLN30),.WL(WL14));
sram_cell_6t_5 inst_cell_14_31 (.BL(BL31),.BLN(BLN31),.WL(WL14));
sram_cell_6t_5 inst_cell_14_32 (.BL(BL32),.BLN(BLN32),.WL(WL14));
sram_cell_6t_5 inst_cell_14_33 (.BL(BL33),.BLN(BLN33),.WL(WL14));
sram_cell_6t_5 inst_cell_14_34 (.BL(BL34),.BLN(BLN34),.WL(WL14));
sram_cell_6t_5 inst_cell_14_35 (.BL(BL35),.BLN(BLN35),.WL(WL14));
sram_cell_6t_5 inst_cell_14_36 (.BL(BL36),.BLN(BLN36),.WL(WL14));
sram_cell_6t_5 inst_cell_14_37 (.BL(BL37),.BLN(BLN37),.WL(WL14));
sram_cell_6t_5 inst_cell_14_38 (.BL(BL38),.BLN(BLN38),.WL(WL14));
sram_cell_6t_5 inst_cell_14_39 (.BL(BL39),.BLN(BLN39),.WL(WL14));
sram_cell_6t_5 inst_cell_14_40 (.BL(BL40),.BLN(BLN40),.WL(WL14));
sram_cell_6t_5 inst_cell_14_41 (.BL(BL41),.BLN(BLN41),.WL(WL14));
sram_cell_6t_5 inst_cell_14_42 (.BL(BL42),.BLN(BLN42),.WL(WL14));
sram_cell_6t_5 inst_cell_14_43 (.BL(BL43),.BLN(BLN43),.WL(WL14));
sram_cell_6t_5 inst_cell_14_44 (.BL(BL44),.BLN(BLN44),.WL(WL14));
sram_cell_6t_5 inst_cell_14_45 (.BL(BL45),.BLN(BLN45),.WL(WL14));
sram_cell_6t_5 inst_cell_14_46 (.BL(BL46),.BLN(BLN46),.WL(WL14));
sram_cell_6t_5 inst_cell_14_47 (.BL(BL47),.BLN(BLN47),.WL(WL14));
sram_cell_6t_5 inst_cell_14_48 (.BL(BL48),.BLN(BLN48),.WL(WL14));
sram_cell_6t_5 inst_cell_14_49 (.BL(BL49),.BLN(BLN49),.WL(WL14));
sram_cell_6t_5 inst_cell_14_50 (.BL(BL50),.BLN(BLN50),.WL(WL14));
sram_cell_6t_5 inst_cell_14_51 (.BL(BL51),.BLN(BLN51),.WL(WL14));
sram_cell_6t_5 inst_cell_14_52 (.BL(BL52),.BLN(BLN52),.WL(WL14));
sram_cell_6t_5 inst_cell_14_53 (.BL(BL53),.BLN(BLN53),.WL(WL14));
sram_cell_6t_5 inst_cell_14_54 (.BL(BL54),.BLN(BLN54),.WL(WL14));
sram_cell_6t_5 inst_cell_14_55 (.BL(BL55),.BLN(BLN55),.WL(WL14));
sram_cell_6t_5 inst_cell_14_56 (.BL(BL56),.BLN(BLN56),.WL(WL14));
sram_cell_6t_5 inst_cell_14_57 (.BL(BL57),.BLN(BLN57),.WL(WL14));
sram_cell_6t_5 inst_cell_14_58 (.BL(BL58),.BLN(BLN58),.WL(WL14));
sram_cell_6t_5 inst_cell_14_59 (.BL(BL59),.BLN(BLN59),.WL(WL14));
sram_cell_6t_5 inst_cell_14_60 (.BL(BL60),.BLN(BLN60),.WL(WL14));
sram_cell_6t_5 inst_cell_14_61 (.BL(BL61),.BLN(BLN61),.WL(WL14));
sram_cell_6t_5 inst_cell_14_62 (.BL(BL62),.BLN(BLN62),.WL(WL14));
sram_cell_6t_5 inst_cell_14_63 (.BL(BL63),.BLN(BLN63),.WL(WL14));
sram_cell_6t_5 inst_cell_14_64 (.BL(BL64),.BLN(BLN64),.WL(WL14));
sram_cell_6t_5 inst_cell_14_65 (.BL(BL65),.BLN(BLN65),.WL(WL14));
sram_cell_6t_5 inst_cell_14_66 (.BL(BL66),.BLN(BLN66),.WL(WL14));
sram_cell_6t_5 inst_cell_14_67 (.BL(BL67),.BLN(BLN67),.WL(WL14));
sram_cell_6t_5 inst_cell_14_68 (.BL(BL68),.BLN(BLN68),.WL(WL14));
sram_cell_6t_5 inst_cell_14_69 (.BL(BL69),.BLN(BLN69),.WL(WL14));
sram_cell_6t_5 inst_cell_14_70 (.BL(BL70),.BLN(BLN70),.WL(WL14));
sram_cell_6t_5 inst_cell_14_71 (.BL(BL71),.BLN(BLN71),.WL(WL14));
sram_cell_6t_5 inst_cell_14_72 (.BL(BL72),.BLN(BLN72),.WL(WL14));
sram_cell_6t_5 inst_cell_14_73 (.BL(BL73),.BLN(BLN73),.WL(WL14));
sram_cell_6t_5 inst_cell_14_74 (.BL(BL74),.BLN(BLN74),.WL(WL14));
sram_cell_6t_5 inst_cell_14_75 (.BL(BL75),.BLN(BLN75),.WL(WL14));
sram_cell_6t_5 inst_cell_14_76 (.BL(BL76),.BLN(BLN76),.WL(WL14));
sram_cell_6t_5 inst_cell_14_77 (.BL(BL77),.BLN(BLN77),.WL(WL14));
sram_cell_6t_5 inst_cell_14_78 (.BL(BL78),.BLN(BLN78),.WL(WL14));
sram_cell_6t_5 inst_cell_14_79 (.BL(BL79),.BLN(BLN79),.WL(WL14));
sram_cell_6t_5 inst_cell_14_80 (.BL(BL80),.BLN(BLN80),.WL(WL14));
sram_cell_6t_5 inst_cell_14_81 (.BL(BL81),.BLN(BLN81),.WL(WL14));
sram_cell_6t_5 inst_cell_14_82 (.BL(BL82),.BLN(BLN82),.WL(WL14));
sram_cell_6t_5 inst_cell_14_83 (.BL(BL83),.BLN(BLN83),.WL(WL14));
sram_cell_6t_5 inst_cell_14_84 (.BL(BL84),.BLN(BLN84),.WL(WL14));
sram_cell_6t_5 inst_cell_14_85 (.BL(BL85),.BLN(BLN85),.WL(WL14));
sram_cell_6t_5 inst_cell_14_86 (.BL(BL86),.BLN(BLN86),.WL(WL14));
sram_cell_6t_5 inst_cell_14_87 (.BL(BL87),.BLN(BLN87),.WL(WL14));
sram_cell_6t_5 inst_cell_14_88 (.BL(BL88),.BLN(BLN88),.WL(WL14));
sram_cell_6t_5 inst_cell_14_89 (.BL(BL89),.BLN(BLN89),.WL(WL14));
sram_cell_6t_5 inst_cell_14_90 (.BL(BL90),.BLN(BLN90),.WL(WL14));
sram_cell_6t_5 inst_cell_14_91 (.BL(BL91),.BLN(BLN91),.WL(WL14));
sram_cell_6t_5 inst_cell_14_92 (.BL(BL92),.BLN(BLN92),.WL(WL14));
sram_cell_6t_5 inst_cell_14_93 (.BL(BL93),.BLN(BLN93),.WL(WL14));
sram_cell_6t_5 inst_cell_14_94 (.BL(BL94),.BLN(BLN94),.WL(WL14));
sram_cell_6t_5 inst_cell_14_95 (.BL(BL95),.BLN(BLN95),.WL(WL14));
sram_cell_6t_5 inst_cell_14_96 (.BL(BL96),.BLN(BLN96),.WL(WL14));
sram_cell_6t_5 inst_cell_14_97 (.BL(BL97),.BLN(BLN97),.WL(WL14));
sram_cell_6t_5 inst_cell_14_98 (.BL(BL98),.BLN(BLN98),.WL(WL14));
sram_cell_6t_5 inst_cell_14_99 (.BL(BL99),.BLN(BLN99),.WL(WL14));
sram_cell_6t_5 inst_cell_14_100 (.BL(BL100),.BLN(BLN100),.WL(WL14));
sram_cell_6t_5 inst_cell_14_101 (.BL(BL101),.BLN(BLN101),.WL(WL14));
sram_cell_6t_5 inst_cell_14_102 (.BL(BL102),.BLN(BLN102),.WL(WL14));
sram_cell_6t_5 inst_cell_14_103 (.BL(BL103),.BLN(BLN103),.WL(WL14));
sram_cell_6t_5 inst_cell_14_104 (.BL(BL104),.BLN(BLN104),.WL(WL14));
sram_cell_6t_5 inst_cell_14_105 (.BL(BL105),.BLN(BLN105),.WL(WL14));
sram_cell_6t_5 inst_cell_14_106 (.BL(BL106),.BLN(BLN106),.WL(WL14));
sram_cell_6t_5 inst_cell_14_107 (.BL(BL107),.BLN(BLN107),.WL(WL14));
sram_cell_6t_5 inst_cell_14_108 (.BL(BL108),.BLN(BLN108),.WL(WL14));
sram_cell_6t_5 inst_cell_14_109 (.BL(BL109),.BLN(BLN109),.WL(WL14));
sram_cell_6t_5 inst_cell_14_110 (.BL(BL110),.BLN(BLN110),.WL(WL14));
sram_cell_6t_5 inst_cell_14_111 (.BL(BL111),.BLN(BLN111),.WL(WL14));
sram_cell_6t_5 inst_cell_14_112 (.BL(BL112),.BLN(BLN112),.WL(WL14));
sram_cell_6t_5 inst_cell_14_113 (.BL(BL113),.BLN(BLN113),.WL(WL14));
sram_cell_6t_5 inst_cell_14_114 (.BL(BL114),.BLN(BLN114),.WL(WL14));
sram_cell_6t_5 inst_cell_14_115 (.BL(BL115),.BLN(BLN115),.WL(WL14));
sram_cell_6t_5 inst_cell_14_116 (.BL(BL116),.BLN(BLN116),.WL(WL14));
sram_cell_6t_5 inst_cell_14_117 (.BL(BL117),.BLN(BLN117),.WL(WL14));
sram_cell_6t_5 inst_cell_14_118 (.BL(BL118),.BLN(BLN118),.WL(WL14));
sram_cell_6t_5 inst_cell_14_119 (.BL(BL119),.BLN(BLN119),.WL(WL14));
sram_cell_6t_5 inst_cell_14_120 (.BL(BL120),.BLN(BLN120),.WL(WL14));
sram_cell_6t_5 inst_cell_14_121 (.BL(BL121),.BLN(BLN121),.WL(WL14));
sram_cell_6t_5 inst_cell_14_122 (.BL(BL122),.BLN(BLN122),.WL(WL14));
sram_cell_6t_5 inst_cell_14_123 (.BL(BL123),.BLN(BLN123),.WL(WL14));
sram_cell_6t_5 inst_cell_14_124 (.BL(BL124),.BLN(BLN124),.WL(WL14));
sram_cell_6t_5 inst_cell_14_125 (.BL(BL125),.BLN(BLN125),.WL(WL14));
sram_cell_6t_5 inst_cell_14_126 (.BL(BL126),.BLN(BLN126),.WL(WL14));
sram_cell_6t_5 inst_cell_14_127 (.BL(BL127),.BLN(BLN127),.WL(WL14));
sram_cell_6t_5 inst_cell_15_0 (.BL(BL0),.BLN(BLN0),.WL(WL15));
sram_cell_6t_5 inst_cell_15_1 (.BL(BL1),.BLN(BLN1),.WL(WL15));
sram_cell_6t_5 inst_cell_15_2 (.BL(BL2),.BLN(BLN2),.WL(WL15));
sram_cell_6t_5 inst_cell_15_3 (.BL(BL3),.BLN(BLN3),.WL(WL15));
sram_cell_6t_5 inst_cell_15_4 (.BL(BL4),.BLN(BLN4),.WL(WL15));
sram_cell_6t_5 inst_cell_15_5 (.BL(BL5),.BLN(BLN5),.WL(WL15));
sram_cell_6t_5 inst_cell_15_6 (.BL(BL6),.BLN(BLN6),.WL(WL15));
sram_cell_6t_5 inst_cell_15_7 (.BL(BL7),.BLN(BLN7),.WL(WL15));
sram_cell_6t_5 inst_cell_15_8 (.BL(BL8),.BLN(BLN8),.WL(WL15));
sram_cell_6t_5 inst_cell_15_9 (.BL(BL9),.BLN(BLN9),.WL(WL15));
sram_cell_6t_5 inst_cell_15_10 (.BL(BL10),.BLN(BLN10),.WL(WL15));
sram_cell_6t_5 inst_cell_15_11 (.BL(BL11),.BLN(BLN11),.WL(WL15));
sram_cell_6t_5 inst_cell_15_12 (.BL(BL12),.BLN(BLN12),.WL(WL15));
sram_cell_6t_5 inst_cell_15_13 (.BL(BL13),.BLN(BLN13),.WL(WL15));
sram_cell_6t_5 inst_cell_15_14 (.BL(BL14),.BLN(BLN14),.WL(WL15));
sram_cell_6t_5 inst_cell_15_15 (.BL(BL15),.BLN(BLN15),.WL(WL15));
sram_cell_6t_5 inst_cell_15_16 (.BL(BL16),.BLN(BLN16),.WL(WL15));
sram_cell_6t_5 inst_cell_15_17 (.BL(BL17),.BLN(BLN17),.WL(WL15));
sram_cell_6t_5 inst_cell_15_18 (.BL(BL18),.BLN(BLN18),.WL(WL15));
sram_cell_6t_5 inst_cell_15_19 (.BL(BL19),.BLN(BLN19),.WL(WL15));
sram_cell_6t_5 inst_cell_15_20 (.BL(BL20),.BLN(BLN20),.WL(WL15));
sram_cell_6t_5 inst_cell_15_21 (.BL(BL21),.BLN(BLN21),.WL(WL15));
sram_cell_6t_5 inst_cell_15_22 (.BL(BL22),.BLN(BLN22),.WL(WL15));
sram_cell_6t_5 inst_cell_15_23 (.BL(BL23),.BLN(BLN23),.WL(WL15));
sram_cell_6t_5 inst_cell_15_24 (.BL(BL24),.BLN(BLN24),.WL(WL15));
sram_cell_6t_5 inst_cell_15_25 (.BL(BL25),.BLN(BLN25),.WL(WL15));
sram_cell_6t_5 inst_cell_15_26 (.BL(BL26),.BLN(BLN26),.WL(WL15));
sram_cell_6t_5 inst_cell_15_27 (.BL(BL27),.BLN(BLN27),.WL(WL15));
sram_cell_6t_5 inst_cell_15_28 (.BL(BL28),.BLN(BLN28),.WL(WL15));
sram_cell_6t_5 inst_cell_15_29 (.BL(BL29),.BLN(BLN29),.WL(WL15));
sram_cell_6t_5 inst_cell_15_30 (.BL(BL30),.BLN(BLN30),.WL(WL15));
sram_cell_6t_5 inst_cell_15_31 (.BL(BL31),.BLN(BLN31),.WL(WL15));
sram_cell_6t_5 inst_cell_15_32 (.BL(BL32),.BLN(BLN32),.WL(WL15));
sram_cell_6t_5 inst_cell_15_33 (.BL(BL33),.BLN(BLN33),.WL(WL15));
sram_cell_6t_5 inst_cell_15_34 (.BL(BL34),.BLN(BLN34),.WL(WL15));
sram_cell_6t_5 inst_cell_15_35 (.BL(BL35),.BLN(BLN35),.WL(WL15));
sram_cell_6t_5 inst_cell_15_36 (.BL(BL36),.BLN(BLN36),.WL(WL15));
sram_cell_6t_5 inst_cell_15_37 (.BL(BL37),.BLN(BLN37),.WL(WL15));
sram_cell_6t_5 inst_cell_15_38 (.BL(BL38),.BLN(BLN38),.WL(WL15));
sram_cell_6t_5 inst_cell_15_39 (.BL(BL39),.BLN(BLN39),.WL(WL15));
sram_cell_6t_5 inst_cell_15_40 (.BL(BL40),.BLN(BLN40),.WL(WL15));
sram_cell_6t_5 inst_cell_15_41 (.BL(BL41),.BLN(BLN41),.WL(WL15));
sram_cell_6t_5 inst_cell_15_42 (.BL(BL42),.BLN(BLN42),.WL(WL15));
sram_cell_6t_5 inst_cell_15_43 (.BL(BL43),.BLN(BLN43),.WL(WL15));
sram_cell_6t_5 inst_cell_15_44 (.BL(BL44),.BLN(BLN44),.WL(WL15));
sram_cell_6t_5 inst_cell_15_45 (.BL(BL45),.BLN(BLN45),.WL(WL15));
sram_cell_6t_5 inst_cell_15_46 (.BL(BL46),.BLN(BLN46),.WL(WL15));
sram_cell_6t_5 inst_cell_15_47 (.BL(BL47),.BLN(BLN47),.WL(WL15));
sram_cell_6t_5 inst_cell_15_48 (.BL(BL48),.BLN(BLN48),.WL(WL15));
sram_cell_6t_5 inst_cell_15_49 (.BL(BL49),.BLN(BLN49),.WL(WL15));
sram_cell_6t_5 inst_cell_15_50 (.BL(BL50),.BLN(BLN50),.WL(WL15));
sram_cell_6t_5 inst_cell_15_51 (.BL(BL51),.BLN(BLN51),.WL(WL15));
sram_cell_6t_5 inst_cell_15_52 (.BL(BL52),.BLN(BLN52),.WL(WL15));
sram_cell_6t_5 inst_cell_15_53 (.BL(BL53),.BLN(BLN53),.WL(WL15));
sram_cell_6t_5 inst_cell_15_54 (.BL(BL54),.BLN(BLN54),.WL(WL15));
sram_cell_6t_5 inst_cell_15_55 (.BL(BL55),.BLN(BLN55),.WL(WL15));
sram_cell_6t_5 inst_cell_15_56 (.BL(BL56),.BLN(BLN56),.WL(WL15));
sram_cell_6t_5 inst_cell_15_57 (.BL(BL57),.BLN(BLN57),.WL(WL15));
sram_cell_6t_5 inst_cell_15_58 (.BL(BL58),.BLN(BLN58),.WL(WL15));
sram_cell_6t_5 inst_cell_15_59 (.BL(BL59),.BLN(BLN59),.WL(WL15));
sram_cell_6t_5 inst_cell_15_60 (.BL(BL60),.BLN(BLN60),.WL(WL15));
sram_cell_6t_5 inst_cell_15_61 (.BL(BL61),.BLN(BLN61),.WL(WL15));
sram_cell_6t_5 inst_cell_15_62 (.BL(BL62),.BLN(BLN62),.WL(WL15));
sram_cell_6t_5 inst_cell_15_63 (.BL(BL63),.BLN(BLN63),.WL(WL15));
sram_cell_6t_5 inst_cell_15_64 (.BL(BL64),.BLN(BLN64),.WL(WL15));
sram_cell_6t_5 inst_cell_15_65 (.BL(BL65),.BLN(BLN65),.WL(WL15));
sram_cell_6t_5 inst_cell_15_66 (.BL(BL66),.BLN(BLN66),.WL(WL15));
sram_cell_6t_5 inst_cell_15_67 (.BL(BL67),.BLN(BLN67),.WL(WL15));
sram_cell_6t_5 inst_cell_15_68 (.BL(BL68),.BLN(BLN68),.WL(WL15));
sram_cell_6t_5 inst_cell_15_69 (.BL(BL69),.BLN(BLN69),.WL(WL15));
sram_cell_6t_5 inst_cell_15_70 (.BL(BL70),.BLN(BLN70),.WL(WL15));
sram_cell_6t_5 inst_cell_15_71 (.BL(BL71),.BLN(BLN71),.WL(WL15));
sram_cell_6t_5 inst_cell_15_72 (.BL(BL72),.BLN(BLN72),.WL(WL15));
sram_cell_6t_5 inst_cell_15_73 (.BL(BL73),.BLN(BLN73),.WL(WL15));
sram_cell_6t_5 inst_cell_15_74 (.BL(BL74),.BLN(BLN74),.WL(WL15));
sram_cell_6t_5 inst_cell_15_75 (.BL(BL75),.BLN(BLN75),.WL(WL15));
sram_cell_6t_5 inst_cell_15_76 (.BL(BL76),.BLN(BLN76),.WL(WL15));
sram_cell_6t_5 inst_cell_15_77 (.BL(BL77),.BLN(BLN77),.WL(WL15));
sram_cell_6t_5 inst_cell_15_78 (.BL(BL78),.BLN(BLN78),.WL(WL15));
sram_cell_6t_5 inst_cell_15_79 (.BL(BL79),.BLN(BLN79),.WL(WL15));
sram_cell_6t_5 inst_cell_15_80 (.BL(BL80),.BLN(BLN80),.WL(WL15));
sram_cell_6t_5 inst_cell_15_81 (.BL(BL81),.BLN(BLN81),.WL(WL15));
sram_cell_6t_5 inst_cell_15_82 (.BL(BL82),.BLN(BLN82),.WL(WL15));
sram_cell_6t_5 inst_cell_15_83 (.BL(BL83),.BLN(BLN83),.WL(WL15));
sram_cell_6t_5 inst_cell_15_84 (.BL(BL84),.BLN(BLN84),.WL(WL15));
sram_cell_6t_5 inst_cell_15_85 (.BL(BL85),.BLN(BLN85),.WL(WL15));
sram_cell_6t_5 inst_cell_15_86 (.BL(BL86),.BLN(BLN86),.WL(WL15));
sram_cell_6t_5 inst_cell_15_87 (.BL(BL87),.BLN(BLN87),.WL(WL15));
sram_cell_6t_5 inst_cell_15_88 (.BL(BL88),.BLN(BLN88),.WL(WL15));
sram_cell_6t_5 inst_cell_15_89 (.BL(BL89),.BLN(BLN89),.WL(WL15));
sram_cell_6t_5 inst_cell_15_90 (.BL(BL90),.BLN(BLN90),.WL(WL15));
sram_cell_6t_5 inst_cell_15_91 (.BL(BL91),.BLN(BLN91),.WL(WL15));
sram_cell_6t_5 inst_cell_15_92 (.BL(BL92),.BLN(BLN92),.WL(WL15));
sram_cell_6t_5 inst_cell_15_93 (.BL(BL93),.BLN(BLN93),.WL(WL15));
sram_cell_6t_5 inst_cell_15_94 (.BL(BL94),.BLN(BLN94),.WL(WL15));
sram_cell_6t_5 inst_cell_15_95 (.BL(BL95),.BLN(BLN95),.WL(WL15));
sram_cell_6t_5 inst_cell_15_96 (.BL(BL96),.BLN(BLN96),.WL(WL15));
sram_cell_6t_5 inst_cell_15_97 (.BL(BL97),.BLN(BLN97),.WL(WL15));
sram_cell_6t_5 inst_cell_15_98 (.BL(BL98),.BLN(BLN98),.WL(WL15));
sram_cell_6t_5 inst_cell_15_99 (.BL(BL99),.BLN(BLN99),.WL(WL15));
sram_cell_6t_5 inst_cell_15_100 (.BL(BL100),.BLN(BLN100),.WL(WL15));
sram_cell_6t_5 inst_cell_15_101 (.BL(BL101),.BLN(BLN101),.WL(WL15));
sram_cell_6t_5 inst_cell_15_102 (.BL(BL102),.BLN(BLN102),.WL(WL15));
sram_cell_6t_5 inst_cell_15_103 (.BL(BL103),.BLN(BLN103),.WL(WL15));
sram_cell_6t_5 inst_cell_15_104 (.BL(BL104),.BLN(BLN104),.WL(WL15));
sram_cell_6t_5 inst_cell_15_105 (.BL(BL105),.BLN(BLN105),.WL(WL15));
sram_cell_6t_5 inst_cell_15_106 (.BL(BL106),.BLN(BLN106),.WL(WL15));
sram_cell_6t_5 inst_cell_15_107 (.BL(BL107),.BLN(BLN107),.WL(WL15));
sram_cell_6t_5 inst_cell_15_108 (.BL(BL108),.BLN(BLN108),.WL(WL15));
sram_cell_6t_5 inst_cell_15_109 (.BL(BL109),.BLN(BLN109),.WL(WL15));
sram_cell_6t_5 inst_cell_15_110 (.BL(BL110),.BLN(BLN110),.WL(WL15));
sram_cell_6t_5 inst_cell_15_111 (.BL(BL111),.BLN(BLN111),.WL(WL15));
sram_cell_6t_5 inst_cell_15_112 (.BL(BL112),.BLN(BLN112),.WL(WL15));
sram_cell_6t_5 inst_cell_15_113 (.BL(BL113),.BLN(BLN113),.WL(WL15));
sram_cell_6t_5 inst_cell_15_114 (.BL(BL114),.BLN(BLN114),.WL(WL15));
sram_cell_6t_5 inst_cell_15_115 (.BL(BL115),.BLN(BLN115),.WL(WL15));
sram_cell_6t_5 inst_cell_15_116 (.BL(BL116),.BLN(BLN116),.WL(WL15));
sram_cell_6t_5 inst_cell_15_117 (.BL(BL117),.BLN(BLN117),.WL(WL15));
sram_cell_6t_5 inst_cell_15_118 (.BL(BL118),.BLN(BLN118),.WL(WL15));
sram_cell_6t_5 inst_cell_15_119 (.BL(BL119),.BLN(BLN119),.WL(WL15));
sram_cell_6t_5 inst_cell_15_120 (.BL(BL120),.BLN(BLN120),.WL(WL15));
sram_cell_6t_5 inst_cell_15_121 (.BL(BL121),.BLN(BLN121),.WL(WL15));
sram_cell_6t_5 inst_cell_15_122 (.BL(BL122),.BLN(BLN122),.WL(WL15));
sram_cell_6t_5 inst_cell_15_123 (.BL(BL123),.BLN(BLN123),.WL(WL15));
sram_cell_6t_5 inst_cell_15_124 (.BL(BL124),.BLN(BLN124),.WL(WL15));
sram_cell_6t_5 inst_cell_15_125 (.BL(BL125),.BLN(BLN125),.WL(WL15));
sram_cell_6t_5 inst_cell_15_126 (.BL(BL126),.BLN(BLN126),.WL(WL15));
sram_cell_6t_5 inst_cell_15_127 (.BL(BL127),.BLN(BLN127),.WL(WL15));
sram_cell_6t_5 inst_cell_16_0 (.BL(BL0),.BLN(BLN0),.WL(WL16));
sram_cell_6t_5 inst_cell_16_1 (.BL(BL1),.BLN(BLN1),.WL(WL16));
sram_cell_6t_5 inst_cell_16_2 (.BL(BL2),.BLN(BLN2),.WL(WL16));
sram_cell_6t_5 inst_cell_16_3 (.BL(BL3),.BLN(BLN3),.WL(WL16));
sram_cell_6t_5 inst_cell_16_4 (.BL(BL4),.BLN(BLN4),.WL(WL16));
sram_cell_6t_5 inst_cell_16_5 (.BL(BL5),.BLN(BLN5),.WL(WL16));
sram_cell_6t_5 inst_cell_16_6 (.BL(BL6),.BLN(BLN6),.WL(WL16));
sram_cell_6t_5 inst_cell_16_7 (.BL(BL7),.BLN(BLN7),.WL(WL16));
sram_cell_6t_5 inst_cell_16_8 (.BL(BL8),.BLN(BLN8),.WL(WL16));
sram_cell_6t_5 inst_cell_16_9 (.BL(BL9),.BLN(BLN9),.WL(WL16));
sram_cell_6t_5 inst_cell_16_10 (.BL(BL10),.BLN(BLN10),.WL(WL16));
sram_cell_6t_5 inst_cell_16_11 (.BL(BL11),.BLN(BLN11),.WL(WL16));
sram_cell_6t_5 inst_cell_16_12 (.BL(BL12),.BLN(BLN12),.WL(WL16));
sram_cell_6t_5 inst_cell_16_13 (.BL(BL13),.BLN(BLN13),.WL(WL16));
sram_cell_6t_5 inst_cell_16_14 (.BL(BL14),.BLN(BLN14),.WL(WL16));
sram_cell_6t_5 inst_cell_16_15 (.BL(BL15),.BLN(BLN15),.WL(WL16));
sram_cell_6t_5 inst_cell_16_16 (.BL(BL16),.BLN(BLN16),.WL(WL16));
sram_cell_6t_5 inst_cell_16_17 (.BL(BL17),.BLN(BLN17),.WL(WL16));
sram_cell_6t_5 inst_cell_16_18 (.BL(BL18),.BLN(BLN18),.WL(WL16));
sram_cell_6t_5 inst_cell_16_19 (.BL(BL19),.BLN(BLN19),.WL(WL16));
sram_cell_6t_5 inst_cell_16_20 (.BL(BL20),.BLN(BLN20),.WL(WL16));
sram_cell_6t_5 inst_cell_16_21 (.BL(BL21),.BLN(BLN21),.WL(WL16));
sram_cell_6t_5 inst_cell_16_22 (.BL(BL22),.BLN(BLN22),.WL(WL16));
sram_cell_6t_5 inst_cell_16_23 (.BL(BL23),.BLN(BLN23),.WL(WL16));
sram_cell_6t_5 inst_cell_16_24 (.BL(BL24),.BLN(BLN24),.WL(WL16));
sram_cell_6t_5 inst_cell_16_25 (.BL(BL25),.BLN(BLN25),.WL(WL16));
sram_cell_6t_5 inst_cell_16_26 (.BL(BL26),.BLN(BLN26),.WL(WL16));
sram_cell_6t_5 inst_cell_16_27 (.BL(BL27),.BLN(BLN27),.WL(WL16));
sram_cell_6t_5 inst_cell_16_28 (.BL(BL28),.BLN(BLN28),.WL(WL16));
sram_cell_6t_5 inst_cell_16_29 (.BL(BL29),.BLN(BLN29),.WL(WL16));
sram_cell_6t_5 inst_cell_16_30 (.BL(BL30),.BLN(BLN30),.WL(WL16));
sram_cell_6t_5 inst_cell_16_31 (.BL(BL31),.BLN(BLN31),.WL(WL16));
sram_cell_6t_5 inst_cell_16_32 (.BL(BL32),.BLN(BLN32),.WL(WL16));
sram_cell_6t_5 inst_cell_16_33 (.BL(BL33),.BLN(BLN33),.WL(WL16));
sram_cell_6t_5 inst_cell_16_34 (.BL(BL34),.BLN(BLN34),.WL(WL16));
sram_cell_6t_5 inst_cell_16_35 (.BL(BL35),.BLN(BLN35),.WL(WL16));
sram_cell_6t_5 inst_cell_16_36 (.BL(BL36),.BLN(BLN36),.WL(WL16));
sram_cell_6t_5 inst_cell_16_37 (.BL(BL37),.BLN(BLN37),.WL(WL16));
sram_cell_6t_5 inst_cell_16_38 (.BL(BL38),.BLN(BLN38),.WL(WL16));
sram_cell_6t_5 inst_cell_16_39 (.BL(BL39),.BLN(BLN39),.WL(WL16));
sram_cell_6t_5 inst_cell_16_40 (.BL(BL40),.BLN(BLN40),.WL(WL16));
sram_cell_6t_5 inst_cell_16_41 (.BL(BL41),.BLN(BLN41),.WL(WL16));
sram_cell_6t_5 inst_cell_16_42 (.BL(BL42),.BLN(BLN42),.WL(WL16));
sram_cell_6t_5 inst_cell_16_43 (.BL(BL43),.BLN(BLN43),.WL(WL16));
sram_cell_6t_5 inst_cell_16_44 (.BL(BL44),.BLN(BLN44),.WL(WL16));
sram_cell_6t_5 inst_cell_16_45 (.BL(BL45),.BLN(BLN45),.WL(WL16));
sram_cell_6t_5 inst_cell_16_46 (.BL(BL46),.BLN(BLN46),.WL(WL16));
sram_cell_6t_5 inst_cell_16_47 (.BL(BL47),.BLN(BLN47),.WL(WL16));
sram_cell_6t_5 inst_cell_16_48 (.BL(BL48),.BLN(BLN48),.WL(WL16));
sram_cell_6t_5 inst_cell_16_49 (.BL(BL49),.BLN(BLN49),.WL(WL16));
sram_cell_6t_5 inst_cell_16_50 (.BL(BL50),.BLN(BLN50),.WL(WL16));
sram_cell_6t_5 inst_cell_16_51 (.BL(BL51),.BLN(BLN51),.WL(WL16));
sram_cell_6t_5 inst_cell_16_52 (.BL(BL52),.BLN(BLN52),.WL(WL16));
sram_cell_6t_5 inst_cell_16_53 (.BL(BL53),.BLN(BLN53),.WL(WL16));
sram_cell_6t_5 inst_cell_16_54 (.BL(BL54),.BLN(BLN54),.WL(WL16));
sram_cell_6t_5 inst_cell_16_55 (.BL(BL55),.BLN(BLN55),.WL(WL16));
sram_cell_6t_5 inst_cell_16_56 (.BL(BL56),.BLN(BLN56),.WL(WL16));
sram_cell_6t_5 inst_cell_16_57 (.BL(BL57),.BLN(BLN57),.WL(WL16));
sram_cell_6t_5 inst_cell_16_58 (.BL(BL58),.BLN(BLN58),.WL(WL16));
sram_cell_6t_5 inst_cell_16_59 (.BL(BL59),.BLN(BLN59),.WL(WL16));
sram_cell_6t_5 inst_cell_16_60 (.BL(BL60),.BLN(BLN60),.WL(WL16));
sram_cell_6t_5 inst_cell_16_61 (.BL(BL61),.BLN(BLN61),.WL(WL16));
sram_cell_6t_5 inst_cell_16_62 (.BL(BL62),.BLN(BLN62),.WL(WL16));
sram_cell_6t_5 inst_cell_16_63 (.BL(BL63),.BLN(BLN63),.WL(WL16));
sram_cell_6t_5 inst_cell_16_64 (.BL(BL64),.BLN(BLN64),.WL(WL16));
sram_cell_6t_5 inst_cell_16_65 (.BL(BL65),.BLN(BLN65),.WL(WL16));
sram_cell_6t_5 inst_cell_16_66 (.BL(BL66),.BLN(BLN66),.WL(WL16));
sram_cell_6t_5 inst_cell_16_67 (.BL(BL67),.BLN(BLN67),.WL(WL16));
sram_cell_6t_5 inst_cell_16_68 (.BL(BL68),.BLN(BLN68),.WL(WL16));
sram_cell_6t_5 inst_cell_16_69 (.BL(BL69),.BLN(BLN69),.WL(WL16));
sram_cell_6t_5 inst_cell_16_70 (.BL(BL70),.BLN(BLN70),.WL(WL16));
sram_cell_6t_5 inst_cell_16_71 (.BL(BL71),.BLN(BLN71),.WL(WL16));
sram_cell_6t_5 inst_cell_16_72 (.BL(BL72),.BLN(BLN72),.WL(WL16));
sram_cell_6t_5 inst_cell_16_73 (.BL(BL73),.BLN(BLN73),.WL(WL16));
sram_cell_6t_5 inst_cell_16_74 (.BL(BL74),.BLN(BLN74),.WL(WL16));
sram_cell_6t_5 inst_cell_16_75 (.BL(BL75),.BLN(BLN75),.WL(WL16));
sram_cell_6t_5 inst_cell_16_76 (.BL(BL76),.BLN(BLN76),.WL(WL16));
sram_cell_6t_5 inst_cell_16_77 (.BL(BL77),.BLN(BLN77),.WL(WL16));
sram_cell_6t_5 inst_cell_16_78 (.BL(BL78),.BLN(BLN78),.WL(WL16));
sram_cell_6t_5 inst_cell_16_79 (.BL(BL79),.BLN(BLN79),.WL(WL16));
sram_cell_6t_5 inst_cell_16_80 (.BL(BL80),.BLN(BLN80),.WL(WL16));
sram_cell_6t_5 inst_cell_16_81 (.BL(BL81),.BLN(BLN81),.WL(WL16));
sram_cell_6t_5 inst_cell_16_82 (.BL(BL82),.BLN(BLN82),.WL(WL16));
sram_cell_6t_5 inst_cell_16_83 (.BL(BL83),.BLN(BLN83),.WL(WL16));
sram_cell_6t_5 inst_cell_16_84 (.BL(BL84),.BLN(BLN84),.WL(WL16));
sram_cell_6t_5 inst_cell_16_85 (.BL(BL85),.BLN(BLN85),.WL(WL16));
sram_cell_6t_5 inst_cell_16_86 (.BL(BL86),.BLN(BLN86),.WL(WL16));
sram_cell_6t_5 inst_cell_16_87 (.BL(BL87),.BLN(BLN87),.WL(WL16));
sram_cell_6t_5 inst_cell_16_88 (.BL(BL88),.BLN(BLN88),.WL(WL16));
sram_cell_6t_5 inst_cell_16_89 (.BL(BL89),.BLN(BLN89),.WL(WL16));
sram_cell_6t_5 inst_cell_16_90 (.BL(BL90),.BLN(BLN90),.WL(WL16));
sram_cell_6t_5 inst_cell_16_91 (.BL(BL91),.BLN(BLN91),.WL(WL16));
sram_cell_6t_5 inst_cell_16_92 (.BL(BL92),.BLN(BLN92),.WL(WL16));
sram_cell_6t_5 inst_cell_16_93 (.BL(BL93),.BLN(BLN93),.WL(WL16));
sram_cell_6t_5 inst_cell_16_94 (.BL(BL94),.BLN(BLN94),.WL(WL16));
sram_cell_6t_5 inst_cell_16_95 (.BL(BL95),.BLN(BLN95),.WL(WL16));
sram_cell_6t_5 inst_cell_16_96 (.BL(BL96),.BLN(BLN96),.WL(WL16));
sram_cell_6t_5 inst_cell_16_97 (.BL(BL97),.BLN(BLN97),.WL(WL16));
sram_cell_6t_5 inst_cell_16_98 (.BL(BL98),.BLN(BLN98),.WL(WL16));
sram_cell_6t_5 inst_cell_16_99 (.BL(BL99),.BLN(BLN99),.WL(WL16));
sram_cell_6t_5 inst_cell_16_100 (.BL(BL100),.BLN(BLN100),.WL(WL16));
sram_cell_6t_5 inst_cell_16_101 (.BL(BL101),.BLN(BLN101),.WL(WL16));
sram_cell_6t_5 inst_cell_16_102 (.BL(BL102),.BLN(BLN102),.WL(WL16));
sram_cell_6t_5 inst_cell_16_103 (.BL(BL103),.BLN(BLN103),.WL(WL16));
sram_cell_6t_5 inst_cell_16_104 (.BL(BL104),.BLN(BLN104),.WL(WL16));
sram_cell_6t_5 inst_cell_16_105 (.BL(BL105),.BLN(BLN105),.WL(WL16));
sram_cell_6t_5 inst_cell_16_106 (.BL(BL106),.BLN(BLN106),.WL(WL16));
sram_cell_6t_5 inst_cell_16_107 (.BL(BL107),.BLN(BLN107),.WL(WL16));
sram_cell_6t_5 inst_cell_16_108 (.BL(BL108),.BLN(BLN108),.WL(WL16));
sram_cell_6t_5 inst_cell_16_109 (.BL(BL109),.BLN(BLN109),.WL(WL16));
sram_cell_6t_5 inst_cell_16_110 (.BL(BL110),.BLN(BLN110),.WL(WL16));
sram_cell_6t_5 inst_cell_16_111 (.BL(BL111),.BLN(BLN111),.WL(WL16));
sram_cell_6t_5 inst_cell_16_112 (.BL(BL112),.BLN(BLN112),.WL(WL16));
sram_cell_6t_5 inst_cell_16_113 (.BL(BL113),.BLN(BLN113),.WL(WL16));
sram_cell_6t_5 inst_cell_16_114 (.BL(BL114),.BLN(BLN114),.WL(WL16));
sram_cell_6t_5 inst_cell_16_115 (.BL(BL115),.BLN(BLN115),.WL(WL16));
sram_cell_6t_5 inst_cell_16_116 (.BL(BL116),.BLN(BLN116),.WL(WL16));
sram_cell_6t_5 inst_cell_16_117 (.BL(BL117),.BLN(BLN117),.WL(WL16));
sram_cell_6t_5 inst_cell_16_118 (.BL(BL118),.BLN(BLN118),.WL(WL16));
sram_cell_6t_5 inst_cell_16_119 (.BL(BL119),.BLN(BLN119),.WL(WL16));
sram_cell_6t_5 inst_cell_16_120 (.BL(BL120),.BLN(BLN120),.WL(WL16));
sram_cell_6t_5 inst_cell_16_121 (.BL(BL121),.BLN(BLN121),.WL(WL16));
sram_cell_6t_5 inst_cell_16_122 (.BL(BL122),.BLN(BLN122),.WL(WL16));
sram_cell_6t_5 inst_cell_16_123 (.BL(BL123),.BLN(BLN123),.WL(WL16));
sram_cell_6t_5 inst_cell_16_124 (.BL(BL124),.BLN(BLN124),.WL(WL16));
sram_cell_6t_5 inst_cell_16_125 (.BL(BL125),.BLN(BLN125),.WL(WL16));
sram_cell_6t_5 inst_cell_16_126 (.BL(BL126),.BLN(BLN126),.WL(WL16));
sram_cell_6t_5 inst_cell_16_127 (.BL(BL127),.BLN(BLN127),.WL(WL16));
sram_cell_6t_5 inst_cell_17_0 (.BL(BL0),.BLN(BLN0),.WL(WL17));
sram_cell_6t_5 inst_cell_17_1 (.BL(BL1),.BLN(BLN1),.WL(WL17));
sram_cell_6t_5 inst_cell_17_2 (.BL(BL2),.BLN(BLN2),.WL(WL17));
sram_cell_6t_5 inst_cell_17_3 (.BL(BL3),.BLN(BLN3),.WL(WL17));
sram_cell_6t_5 inst_cell_17_4 (.BL(BL4),.BLN(BLN4),.WL(WL17));
sram_cell_6t_5 inst_cell_17_5 (.BL(BL5),.BLN(BLN5),.WL(WL17));
sram_cell_6t_5 inst_cell_17_6 (.BL(BL6),.BLN(BLN6),.WL(WL17));
sram_cell_6t_5 inst_cell_17_7 (.BL(BL7),.BLN(BLN7),.WL(WL17));
sram_cell_6t_5 inst_cell_17_8 (.BL(BL8),.BLN(BLN8),.WL(WL17));
sram_cell_6t_5 inst_cell_17_9 (.BL(BL9),.BLN(BLN9),.WL(WL17));
sram_cell_6t_5 inst_cell_17_10 (.BL(BL10),.BLN(BLN10),.WL(WL17));
sram_cell_6t_5 inst_cell_17_11 (.BL(BL11),.BLN(BLN11),.WL(WL17));
sram_cell_6t_5 inst_cell_17_12 (.BL(BL12),.BLN(BLN12),.WL(WL17));
sram_cell_6t_5 inst_cell_17_13 (.BL(BL13),.BLN(BLN13),.WL(WL17));
sram_cell_6t_5 inst_cell_17_14 (.BL(BL14),.BLN(BLN14),.WL(WL17));
sram_cell_6t_5 inst_cell_17_15 (.BL(BL15),.BLN(BLN15),.WL(WL17));
sram_cell_6t_5 inst_cell_17_16 (.BL(BL16),.BLN(BLN16),.WL(WL17));
sram_cell_6t_5 inst_cell_17_17 (.BL(BL17),.BLN(BLN17),.WL(WL17));
sram_cell_6t_5 inst_cell_17_18 (.BL(BL18),.BLN(BLN18),.WL(WL17));
sram_cell_6t_5 inst_cell_17_19 (.BL(BL19),.BLN(BLN19),.WL(WL17));
sram_cell_6t_5 inst_cell_17_20 (.BL(BL20),.BLN(BLN20),.WL(WL17));
sram_cell_6t_5 inst_cell_17_21 (.BL(BL21),.BLN(BLN21),.WL(WL17));
sram_cell_6t_5 inst_cell_17_22 (.BL(BL22),.BLN(BLN22),.WL(WL17));
sram_cell_6t_5 inst_cell_17_23 (.BL(BL23),.BLN(BLN23),.WL(WL17));
sram_cell_6t_5 inst_cell_17_24 (.BL(BL24),.BLN(BLN24),.WL(WL17));
sram_cell_6t_5 inst_cell_17_25 (.BL(BL25),.BLN(BLN25),.WL(WL17));
sram_cell_6t_5 inst_cell_17_26 (.BL(BL26),.BLN(BLN26),.WL(WL17));
sram_cell_6t_5 inst_cell_17_27 (.BL(BL27),.BLN(BLN27),.WL(WL17));
sram_cell_6t_5 inst_cell_17_28 (.BL(BL28),.BLN(BLN28),.WL(WL17));
sram_cell_6t_5 inst_cell_17_29 (.BL(BL29),.BLN(BLN29),.WL(WL17));
sram_cell_6t_5 inst_cell_17_30 (.BL(BL30),.BLN(BLN30),.WL(WL17));
sram_cell_6t_5 inst_cell_17_31 (.BL(BL31),.BLN(BLN31),.WL(WL17));
sram_cell_6t_5 inst_cell_17_32 (.BL(BL32),.BLN(BLN32),.WL(WL17));
sram_cell_6t_5 inst_cell_17_33 (.BL(BL33),.BLN(BLN33),.WL(WL17));
sram_cell_6t_5 inst_cell_17_34 (.BL(BL34),.BLN(BLN34),.WL(WL17));
sram_cell_6t_5 inst_cell_17_35 (.BL(BL35),.BLN(BLN35),.WL(WL17));
sram_cell_6t_5 inst_cell_17_36 (.BL(BL36),.BLN(BLN36),.WL(WL17));
sram_cell_6t_5 inst_cell_17_37 (.BL(BL37),.BLN(BLN37),.WL(WL17));
sram_cell_6t_5 inst_cell_17_38 (.BL(BL38),.BLN(BLN38),.WL(WL17));
sram_cell_6t_5 inst_cell_17_39 (.BL(BL39),.BLN(BLN39),.WL(WL17));
sram_cell_6t_5 inst_cell_17_40 (.BL(BL40),.BLN(BLN40),.WL(WL17));
sram_cell_6t_5 inst_cell_17_41 (.BL(BL41),.BLN(BLN41),.WL(WL17));
sram_cell_6t_5 inst_cell_17_42 (.BL(BL42),.BLN(BLN42),.WL(WL17));
sram_cell_6t_5 inst_cell_17_43 (.BL(BL43),.BLN(BLN43),.WL(WL17));
sram_cell_6t_5 inst_cell_17_44 (.BL(BL44),.BLN(BLN44),.WL(WL17));
sram_cell_6t_5 inst_cell_17_45 (.BL(BL45),.BLN(BLN45),.WL(WL17));
sram_cell_6t_5 inst_cell_17_46 (.BL(BL46),.BLN(BLN46),.WL(WL17));
sram_cell_6t_5 inst_cell_17_47 (.BL(BL47),.BLN(BLN47),.WL(WL17));
sram_cell_6t_5 inst_cell_17_48 (.BL(BL48),.BLN(BLN48),.WL(WL17));
sram_cell_6t_5 inst_cell_17_49 (.BL(BL49),.BLN(BLN49),.WL(WL17));
sram_cell_6t_5 inst_cell_17_50 (.BL(BL50),.BLN(BLN50),.WL(WL17));
sram_cell_6t_5 inst_cell_17_51 (.BL(BL51),.BLN(BLN51),.WL(WL17));
sram_cell_6t_5 inst_cell_17_52 (.BL(BL52),.BLN(BLN52),.WL(WL17));
sram_cell_6t_5 inst_cell_17_53 (.BL(BL53),.BLN(BLN53),.WL(WL17));
sram_cell_6t_5 inst_cell_17_54 (.BL(BL54),.BLN(BLN54),.WL(WL17));
sram_cell_6t_5 inst_cell_17_55 (.BL(BL55),.BLN(BLN55),.WL(WL17));
sram_cell_6t_5 inst_cell_17_56 (.BL(BL56),.BLN(BLN56),.WL(WL17));
sram_cell_6t_5 inst_cell_17_57 (.BL(BL57),.BLN(BLN57),.WL(WL17));
sram_cell_6t_5 inst_cell_17_58 (.BL(BL58),.BLN(BLN58),.WL(WL17));
sram_cell_6t_5 inst_cell_17_59 (.BL(BL59),.BLN(BLN59),.WL(WL17));
sram_cell_6t_5 inst_cell_17_60 (.BL(BL60),.BLN(BLN60),.WL(WL17));
sram_cell_6t_5 inst_cell_17_61 (.BL(BL61),.BLN(BLN61),.WL(WL17));
sram_cell_6t_5 inst_cell_17_62 (.BL(BL62),.BLN(BLN62),.WL(WL17));
sram_cell_6t_5 inst_cell_17_63 (.BL(BL63),.BLN(BLN63),.WL(WL17));
sram_cell_6t_5 inst_cell_17_64 (.BL(BL64),.BLN(BLN64),.WL(WL17));
sram_cell_6t_5 inst_cell_17_65 (.BL(BL65),.BLN(BLN65),.WL(WL17));
sram_cell_6t_5 inst_cell_17_66 (.BL(BL66),.BLN(BLN66),.WL(WL17));
sram_cell_6t_5 inst_cell_17_67 (.BL(BL67),.BLN(BLN67),.WL(WL17));
sram_cell_6t_5 inst_cell_17_68 (.BL(BL68),.BLN(BLN68),.WL(WL17));
sram_cell_6t_5 inst_cell_17_69 (.BL(BL69),.BLN(BLN69),.WL(WL17));
sram_cell_6t_5 inst_cell_17_70 (.BL(BL70),.BLN(BLN70),.WL(WL17));
sram_cell_6t_5 inst_cell_17_71 (.BL(BL71),.BLN(BLN71),.WL(WL17));
sram_cell_6t_5 inst_cell_17_72 (.BL(BL72),.BLN(BLN72),.WL(WL17));
sram_cell_6t_5 inst_cell_17_73 (.BL(BL73),.BLN(BLN73),.WL(WL17));
sram_cell_6t_5 inst_cell_17_74 (.BL(BL74),.BLN(BLN74),.WL(WL17));
sram_cell_6t_5 inst_cell_17_75 (.BL(BL75),.BLN(BLN75),.WL(WL17));
sram_cell_6t_5 inst_cell_17_76 (.BL(BL76),.BLN(BLN76),.WL(WL17));
sram_cell_6t_5 inst_cell_17_77 (.BL(BL77),.BLN(BLN77),.WL(WL17));
sram_cell_6t_5 inst_cell_17_78 (.BL(BL78),.BLN(BLN78),.WL(WL17));
sram_cell_6t_5 inst_cell_17_79 (.BL(BL79),.BLN(BLN79),.WL(WL17));
sram_cell_6t_5 inst_cell_17_80 (.BL(BL80),.BLN(BLN80),.WL(WL17));
sram_cell_6t_5 inst_cell_17_81 (.BL(BL81),.BLN(BLN81),.WL(WL17));
sram_cell_6t_5 inst_cell_17_82 (.BL(BL82),.BLN(BLN82),.WL(WL17));
sram_cell_6t_5 inst_cell_17_83 (.BL(BL83),.BLN(BLN83),.WL(WL17));
sram_cell_6t_5 inst_cell_17_84 (.BL(BL84),.BLN(BLN84),.WL(WL17));
sram_cell_6t_5 inst_cell_17_85 (.BL(BL85),.BLN(BLN85),.WL(WL17));
sram_cell_6t_5 inst_cell_17_86 (.BL(BL86),.BLN(BLN86),.WL(WL17));
sram_cell_6t_5 inst_cell_17_87 (.BL(BL87),.BLN(BLN87),.WL(WL17));
sram_cell_6t_5 inst_cell_17_88 (.BL(BL88),.BLN(BLN88),.WL(WL17));
sram_cell_6t_5 inst_cell_17_89 (.BL(BL89),.BLN(BLN89),.WL(WL17));
sram_cell_6t_5 inst_cell_17_90 (.BL(BL90),.BLN(BLN90),.WL(WL17));
sram_cell_6t_5 inst_cell_17_91 (.BL(BL91),.BLN(BLN91),.WL(WL17));
sram_cell_6t_5 inst_cell_17_92 (.BL(BL92),.BLN(BLN92),.WL(WL17));
sram_cell_6t_5 inst_cell_17_93 (.BL(BL93),.BLN(BLN93),.WL(WL17));
sram_cell_6t_5 inst_cell_17_94 (.BL(BL94),.BLN(BLN94),.WL(WL17));
sram_cell_6t_5 inst_cell_17_95 (.BL(BL95),.BLN(BLN95),.WL(WL17));
sram_cell_6t_5 inst_cell_17_96 (.BL(BL96),.BLN(BLN96),.WL(WL17));
sram_cell_6t_5 inst_cell_17_97 (.BL(BL97),.BLN(BLN97),.WL(WL17));
sram_cell_6t_5 inst_cell_17_98 (.BL(BL98),.BLN(BLN98),.WL(WL17));
sram_cell_6t_5 inst_cell_17_99 (.BL(BL99),.BLN(BLN99),.WL(WL17));
sram_cell_6t_5 inst_cell_17_100 (.BL(BL100),.BLN(BLN100),.WL(WL17));
sram_cell_6t_5 inst_cell_17_101 (.BL(BL101),.BLN(BLN101),.WL(WL17));
sram_cell_6t_5 inst_cell_17_102 (.BL(BL102),.BLN(BLN102),.WL(WL17));
sram_cell_6t_5 inst_cell_17_103 (.BL(BL103),.BLN(BLN103),.WL(WL17));
sram_cell_6t_5 inst_cell_17_104 (.BL(BL104),.BLN(BLN104),.WL(WL17));
sram_cell_6t_5 inst_cell_17_105 (.BL(BL105),.BLN(BLN105),.WL(WL17));
sram_cell_6t_5 inst_cell_17_106 (.BL(BL106),.BLN(BLN106),.WL(WL17));
sram_cell_6t_5 inst_cell_17_107 (.BL(BL107),.BLN(BLN107),.WL(WL17));
sram_cell_6t_5 inst_cell_17_108 (.BL(BL108),.BLN(BLN108),.WL(WL17));
sram_cell_6t_5 inst_cell_17_109 (.BL(BL109),.BLN(BLN109),.WL(WL17));
sram_cell_6t_5 inst_cell_17_110 (.BL(BL110),.BLN(BLN110),.WL(WL17));
sram_cell_6t_5 inst_cell_17_111 (.BL(BL111),.BLN(BLN111),.WL(WL17));
sram_cell_6t_5 inst_cell_17_112 (.BL(BL112),.BLN(BLN112),.WL(WL17));
sram_cell_6t_5 inst_cell_17_113 (.BL(BL113),.BLN(BLN113),.WL(WL17));
sram_cell_6t_5 inst_cell_17_114 (.BL(BL114),.BLN(BLN114),.WL(WL17));
sram_cell_6t_5 inst_cell_17_115 (.BL(BL115),.BLN(BLN115),.WL(WL17));
sram_cell_6t_5 inst_cell_17_116 (.BL(BL116),.BLN(BLN116),.WL(WL17));
sram_cell_6t_5 inst_cell_17_117 (.BL(BL117),.BLN(BLN117),.WL(WL17));
sram_cell_6t_5 inst_cell_17_118 (.BL(BL118),.BLN(BLN118),.WL(WL17));
sram_cell_6t_5 inst_cell_17_119 (.BL(BL119),.BLN(BLN119),.WL(WL17));
sram_cell_6t_5 inst_cell_17_120 (.BL(BL120),.BLN(BLN120),.WL(WL17));
sram_cell_6t_5 inst_cell_17_121 (.BL(BL121),.BLN(BLN121),.WL(WL17));
sram_cell_6t_5 inst_cell_17_122 (.BL(BL122),.BLN(BLN122),.WL(WL17));
sram_cell_6t_5 inst_cell_17_123 (.BL(BL123),.BLN(BLN123),.WL(WL17));
sram_cell_6t_5 inst_cell_17_124 (.BL(BL124),.BLN(BLN124),.WL(WL17));
sram_cell_6t_5 inst_cell_17_125 (.BL(BL125),.BLN(BLN125),.WL(WL17));
sram_cell_6t_5 inst_cell_17_126 (.BL(BL126),.BLN(BLN126),.WL(WL17));
sram_cell_6t_5 inst_cell_17_127 (.BL(BL127),.BLN(BLN127),.WL(WL17));
sram_cell_6t_5 inst_cell_18_0 (.BL(BL0),.BLN(BLN0),.WL(WL18));
sram_cell_6t_5 inst_cell_18_1 (.BL(BL1),.BLN(BLN1),.WL(WL18));
sram_cell_6t_5 inst_cell_18_2 (.BL(BL2),.BLN(BLN2),.WL(WL18));
sram_cell_6t_5 inst_cell_18_3 (.BL(BL3),.BLN(BLN3),.WL(WL18));
sram_cell_6t_5 inst_cell_18_4 (.BL(BL4),.BLN(BLN4),.WL(WL18));
sram_cell_6t_5 inst_cell_18_5 (.BL(BL5),.BLN(BLN5),.WL(WL18));
sram_cell_6t_5 inst_cell_18_6 (.BL(BL6),.BLN(BLN6),.WL(WL18));
sram_cell_6t_5 inst_cell_18_7 (.BL(BL7),.BLN(BLN7),.WL(WL18));
sram_cell_6t_5 inst_cell_18_8 (.BL(BL8),.BLN(BLN8),.WL(WL18));
sram_cell_6t_5 inst_cell_18_9 (.BL(BL9),.BLN(BLN9),.WL(WL18));
sram_cell_6t_5 inst_cell_18_10 (.BL(BL10),.BLN(BLN10),.WL(WL18));
sram_cell_6t_5 inst_cell_18_11 (.BL(BL11),.BLN(BLN11),.WL(WL18));
sram_cell_6t_5 inst_cell_18_12 (.BL(BL12),.BLN(BLN12),.WL(WL18));
sram_cell_6t_5 inst_cell_18_13 (.BL(BL13),.BLN(BLN13),.WL(WL18));
sram_cell_6t_5 inst_cell_18_14 (.BL(BL14),.BLN(BLN14),.WL(WL18));
sram_cell_6t_5 inst_cell_18_15 (.BL(BL15),.BLN(BLN15),.WL(WL18));
sram_cell_6t_5 inst_cell_18_16 (.BL(BL16),.BLN(BLN16),.WL(WL18));
sram_cell_6t_5 inst_cell_18_17 (.BL(BL17),.BLN(BLN17),.WL(WL18));
sram_cell_6t_5 inst_cell_18_18 (.BL(BL18),.BLN(BLN18),.WL(WL18));
sram_cell_6t_5 inst_cell_18_19 (.BL(BL19),.BLN(BLN19),.WL(WL18));
sram_cell_6t_5 inst_cell_18_20 (.BL(BL20),.BLN(BLN20),.WL(WL18));
sram_cell_6t_5 inst_cell_18_21 (.BL(BL21),.BLN(BLN21),.WL(WL18));
sram_cell_6t_5 inst_cell_18_22 (.BL(BL22),.BLN(BLN22),.WL(WL18));
sram_cell_6t_5 inst_cell_18_23 (.BL(BL23),.BLN(BLN23),.WL(WL18));
sram_cell_6t_5 inst_cell_18_24 (.BL(BL24),.BLN(BLN24),.WL(WL18));
sram_cell_6t_5 inst_cell_18_25 (.BL(BL25),.BLN(BLN25),.WL(WL18));
sram_cell_6t_5 inst_cell_18_26 (.BL(BL26),.BLN(BLN26),.WL(WL18));
sram_cell_6t_5 inst_cell_18_27 (.BL(BL27),.BLN(BLN27),.WL(WL18));
sram_cell_6t_5 inst_cell_18_28 (.BL(BL28),.BLN(BLN28),.WL(WL18));
sram_cell_6t_5 inst_cell_18_29 (.BL(BL29),.BLN(BLN29),.WL(WL18));
sram_cell_6t_5 inst_cell_18_30 (.BL(BL30),.BLN(BLN30),.WL(WL18));
sram_cell_6t_5 inst_cell_18_31 (.BL(BL31),.BLN(BLN31),.WL(WL18));
sram_cell_6t_5 inst_cell_18_32 (.BL(BL32),.BLN(BLN32),.WL(WL18));
sram_cell_6t_5 inst_cell_18_33 (.BL(BL33),.BLN(BLN33),.WL(WL18));
sram_cell_6t_5 inst_cell_18_34 (.BL(BL34),.BLN(BLN34),.WL(WL18));
sram_cell_6t_5 inst_cell_18_35 (.BL(BL35),.BLN(BLN35),.WL(WL18));
sram_cell_6t_5 inst_cell_18_36 (.BL(BL36),.BLN(BLN36),.WL(WL18));
sram_cell_6t_5 inst_cell_18_37 (.BL(BL37),.BLN(BLN37),.WL(WL18));
sram_cell_6t_5 inst_cell_18_38 (.BL(BL38),.BLN(BLN38),.WL(WL18));
sram_cell_6t_5 inst_cell_18_39 (.BL(BL39),.BLN(BLN39),.WL(WL18));
sram_cell_6t_5 inst_cell_18_40 (.BL(BL40),.BLN(BLN40),.WL(WL18));
sram_cell_6t_5 inst_cell_18_41 (.BL(BL41),.BLN(BLN41),.WL(WL18));
sram_cell_6t_5 inst_cell_18_42 (.BL(BL42),.BLN(BLN42),.WL(WL18));
sram_cell_6t_5 inst_cell_18_43 (.BL(BL43),.BLN(BLN43),.WL(WL18));
sram_cell_6t_5 inst_cell_18_44 (.BL(BL44),.BLN(BLN44),.WL(WL18));
sram_cell_6t_5 inst_cell_18_45 (.BL(BL45),.BLN(BLN45),.WL(WL18));
sram_cell_6t_5 inst_cell_18_46 (.BL(BL46),.BLN(BLN46),.WL(WL18));
sram_cell_6t_5 inst_cell_18_47 (.BL(BL47),.BLN(BLN47),.WL(WL18));
sram_cell_6t_5 inst_cell_18_48 (.BL(BL48),.BLN(BLN48),.WL(WL18));
sram_cell_6t_5 inst_cell_18_49 (.BL(BL49),.BLN(BLN49),.WL(WL18));
sram_cell_6t_5 inst_cell_18_50 (.BL(BL50),.BLN(BLN50),.WL(WL18));
sram_cell_6t_5 inst_cell_18_51 (.BL(BL51),.BLN(BLN51),.WL(WL18));
sram_cell_6t_5 inst_cell_18_52 (.BL(BL52),.BLN(BLN52),.WL(WL18));
sram_cell_6t_5 inst_cell_18_53 (.BL(BL53),.BLN(BLN53),.WL(WL18));
sram_cell_6t_5 inst_cell_18_54 (.BL(BL54),.BLN(BLN54),.WL(WL18));
sram_cell_6t_5 inst_cell_18_55 (.BL(BL55),.BLN(BLN55),.WL(WL18));
sram_cell_6t_5 inst_cell_18_56 (.BL(BL56),.BLN(BLN56),.WL(WL18));
sram_cell_6t_5 inst_cell_18_57 (.BL(BL57),.BLN(BLN57),.WL(WL18));
sram_cell_6t_5 inst_cell_18_58 (.BL(BL58),.BLN(BLN58),.WL(WL18));
sram_cell_6t_5 inst_cell_18_59 (.BL(BL59),.BLN(BLN59),.WL(WL18));
sram_cell_6t_5 inst_cell_18_60 (.BL(BL60),.BLN(BLN60),.WL(WL18));
sram_cell_6t_5 inst_cell_18_61 (.BL(BL61),.BLN(BLN61),.WL(WL18));
sram_cell_6t_5 inst_cell_18_62 (.BL(BL62),.BLN(BLN62),.WL(WL18));
sram_cell_6t_5 inst_cell_18_63 (.BL(BL63),.BLN(BLN63),.WL(WL18));
sram_cell_6t_5 inst_cell_18_64 (.BL(BL64),.BLN(BLN64),.WL(WL18));
sram_cell_6t_5 inst_cell_18_65 (.BL(BL65),.BLN(BLN65),.WL(WL18));
sram_cell_6t_5 inst_cell_18_66 (.BL(BL66),.BLN(BLN66),.WL(WL18));
sram_cell_6t_5 inst_cell_18_67 (.BL(BL67),.BLN(BLN67),.WL(WL18));
sram_cell_6t_5 inst_cell_18_68 (.BL(BL68),.BLN(BLN68),.WL(WL18));
sram_cell_6t_5 inst_cell_18_69 (.BL(BL69),.BLN(BLN69),.WL(WL18));
sram_cell_6t_5 inst_cell_18_70 (.BL(BL70),.BLN(BLN70),.WL(WL18));
sram_cell_6t_5 inst_cell_18_71 (.BL(BL71),.BLN(BLN71),.WL(WL18));
sram_cell_6t_5 inst_cell_18_72 (.BL(BL72),.BLN(BLN72),.WL(WL18));
sram_cell_6t_5 inst_cell_18_73 (.BL(BL73),.BLN(BLN73),.WL(WL18));
sram_cell_6t_5 inst_cell_18_74 (.BL(BL74),.BLN(BLN74),.WL(WL18));
sram_cell_6t_5 inst_cell_18_75 (.BL(BL75),.BLN(BLN75),.WL(WL18));
sram_cell_6t_5 inst_cell_18_76 (.BL(BL76),.BLN(BLN76),.WL(WL18));
sram_cell_6t_5 inst_cell_18_77 (.BL(BL77),.BLN(BLN77),.WL(WL18));
sram_cell_6t_5 inst_cell_18_78 (.BL(BL78),.BLN(BLN78),.WL(WL18));
sram_cell_6t_5 inst_cell_18_79 (.BL(BL79),.BLN(BLN79),.WL(WL18));
sram_cell_6t_5 inst_cell_18_80 (.BL(BL80),.BLN(BLN80),.WL(WL18));
sram_cell_6t_5 inst_cell_18_81 (.BL(BL81),.BLN(BLN81),.WL(WL18));
sram_cell_6t_5 inst_cell_18_82 (.BL(BL82),.BLN(BLN82),.WL(WL18));
sram_cell_6t_5 inst_cell_18_83 (.BL(BL83),.BLN(BLN83),.WL(WL18));
sram_cell_6t_5 inst_cell_18_84 (.BL(BL84),.BLN(BLN84),.WL(WL18));
sram_cell_6t_5 inst_cell_18_85 (.BL(BL85),.BLN(BLN85),.WL(WL18));
sram_cell_6t_5 inst_cell_18_86 (.BL(BL86),.BLN(BLN86),.WL(WL18));
sram_cell_6t_5 inst_cell_18_87 (.BL(BL87),.BLN(BLN87),.WL(WL18));
sram_cell_6t_5 inst_cell_18_88 (.BL(BL88),.BLN(BLN88),.WL(WL18));
sram_cell_6t_5 inst_cell_18_89 (.BL(BL89),.BLN(BLN89),.WL(WL18));
sram_cell_6t_5 inst_cell_18_90 (.BL(BL90),.BLN(BLN90),.WL(WL18));
sram_cell_6t_5 inst_cell_18_91 (.BL(BL91),.BLN(BLN91),.WL(WL18));
sram_cell_6t_5 inst_cell_18_92 (.BL(BL92),.BLN(BLN92),.WL(WL18));
sram_cell_6t_5 inst_cell_18_93 (.BL(BL93),.BLN(BLN93),.WL(WL18));
sram_cell_6t_5 inst_cell_18_94 (.BL(BL94),.BLN(BLN94),.WL(WL18));
sram_cell_6t_5 inst_cell_18_95 (.BL(BL95),.BLN(BLN95),.WL(WL18));
sram_cell_6t_5 inst_cell_18_96 (.BL(BL96),.BLN(BLN96),.WL(WL18));
sram_cell_6t_5 inst_cell_18_97 (.BL(BL97),.BLN(BLN97),.WL(WL18));
sram_cell_6t_5 inst_cell_18_98 (.BL(BL98),.BLN(BLN98),.WL(WL18));
sram_cell_6t_5 inst_cell_18_99 (.BL(BL99),.BLN(BLN99),.WL(WL18));
sram_cell_6t_5 inst_cell_18_100 (.BL(BL100),.BLN(BLN100),.WL(WL18));
sram_cell_6t_5 inst_cell_18_101 (.BL(BL101),.BLN(BLN101),.WL(WL18));
sram_cell_6t_5 inst_cell_18_102 (.BL(BL102),.BLN(BLN102),.WL(WL18));
sram_cell_6t_5 inst_cell_18_103 (.BL(BL103),.BLN(BLN103),.WL(WL18));
sram_cell_6t_5 inst_cell_18_104 (.BL(BL104),.BLN(BLN104),.WL(WL18));
sram_cell_6t_5 inst_cell_18_105 (.BL(BL105),.BLN(BLN105),.WL(WL18));
sram_cell_6t_5 inst_cell_18_106 (.BL(BL106),.BLN(BLN106),.WL(WL18));
sram_cell_6t_5 inst_cell_18_107 (.BL(BL107),.BLN(BLN107),.WL(WL18));
sram_cell_6t_5 inst_cell_18_108 (.BL(BL108),.BLN(BLN108),.WL(WL18));
sram_cell_6t_5 inst_cell_18_109 (.BL(BL109),.BLN(BLN109),.WL(WL18));
sram_cell_6t_5 inst_cell_18_110 (.BL(BL110),.BLN(BLN110),.WL(WL18));
sram_cell_6t_5 inst_cell_18_111 (.BL(BL111),.BLN(BLN111),.WL(WL18));
sram_cell_6t_5 inst_cell_18_112 (.BL(BL112),.BLN(BLN112),.WL(WL18));
sram_cell_6t_5 inst_cell_18_113 (.BL(BL113),.BLN(BLN113),.WL(WL18));
sram_cell_6t_5 inst_cell_18_114 (.BL(BL114),.BLN(BLN114),.WL(WL18));
sram_cell_6t_5 inst_cell_18_115 (.BL(BL115),.BLN(BLN115),.WL(WL18));
sram_cell_6t_5 inst_cell_18_116 (.BL(BL116),.BLN(BLN116),.WL(WL18));
sram_cell_6t_5 inst_cell_18_117 (.BL(BL117),.BLN(BLN117),.WL(WL18));
sram_cell_6t_5 inst_cell_18_118 (.BL(BL118),.BLN(BLN118),.WL(WL18));
sram_cell_6t_5 inst_cell_18_119 (.BL(BL119),.BLN(BLN119),.WL(WL18));
sram_cell_6t_5 inst_cell_18_120 (.BL(BL120),.BLN(BLN120),.WL(WL18));
sram_cell_6t_5 inst_cell_18_121 (.BL(BL121),.BLN(BLN121),.WL(WL18));
sram_cell_6t_5 inst_cell_18_122 (.BL(BL122),.BLN(BLN122),.WL(WL18));
sram_cell_6t_5 inst_cell_18_123 (.BL(BL123),.BLN(BLN123),.WL(WL18));
sram_cell_6t_5 inst_cell_18_124 (.BL(BL124),.BLN(BLN124),.WL(WL18));
sram_cell_6t_5 inst_cell_18_125 (.BL(BL125),.BLN(BLN125),.WL(WL18));
sram_cell_6t_5 inst_cell_18_126 (.BL(BL126),.BLN(BLN126),.WL(WL18));
sram_cell_6t_5 inst_cell_18_127 (.BL(BL127),.BLN(BLN127),.WL(WL18));
sram_cell_6t_5 inst_cell_19_0 (.BL(BL0),.BLN(BLN0),.WL(WL19));
sram_cell_6t_5 inst_cell_19_1 (.BL(BL1),.BLN(BLN1),.WL(WL19));
sram_cell_6t_5 inst_cell_19_2 (.BL(BL2),.BLN(BLN2),.WL(WL19));
sram_cell_6t_5 inst_cell_19_3 (.BL(BL3),.BLN(BLN3),.WL(WL19));
sram_cell_6t_5 inst_cell_19_4 (.BL(BL4),.BLN(BLN4),.WL(WL19));
sram_cell_6t_5 inst_cell_19_5 (.BL(BL5),.BLN(BLN5),.WL(WL19));
sram_cell_6t_5 inst_cell_19_6 (.BL(BL6),.BLN(BLN6),.WL(WL19));
sram_cell_6t_5 inst_cell_19_7 (.BL(BL7),.BLN(BLN7),.WL(WL19));
sram_cell_6t_5 inst_cell_19_8 (.BL(BL8),.BLN(BLN8),.WL(WL19));
sram_cell_6t_5 inst_cell_19_9 (.BL(BL9),.BLN(BLN9),.WL(WL19));
sram_cell_6t_5 inst_cell_19_10 (.BL(BL10),.BLN(BLN10),.WL(WL19));
sram_cell_6t_5 inst_cell_19_11 (.BL(BL11),.BLN(BLN11),.WL(WL19));
sram_cell_6t_5 inst_cell_19_12 (.BL(BL12),.BLN(BLN12),.WL(WL19));
sram_cell_6t_5 inst_cell_19_13 (.BL(BL13),.BLN(BLN13),.WL(WL19));
sram_cell_6t_5 inst_cell_19_14 (.BL(BL14),.BLN(BLN14),.WL(WL19));
sram_cell_6t_5 inst_cell_19_15 (.BL(BL15),.BLN(BLN15),.WL(WL19));
sram_cell_6t_5 inst_cell_19_16 (.BL(BL16),.BLN(BLN16),.WL(WL19));
sram_cell_6t_5 inst_cell_19_17 (.BL(BL17),.BLN(BLN17),.WL(WL19));
sram_cell_6t_5 inst_cell_19_18 (.BL(BL18),.BLN(BLN18),.WL(WL19));
sram_cell_6t_5 inst_cell_19_19 (.BL(BL19),.BLN(BLN19),.WL(WL19));
sram_cell_6t_5 inst_cell_19_20 (.BL(BL20),.BLN(BLN20),.WL(WL19));
sram_cell_6t_5 inst_cell_19_21 (.BL(BL21),.BLN(BLN21),.WL(WL19));
sram_cell_6t_5 inst_cell_19_22 (.BL(BL22),.BLN(BLN22),.WL(WL19));
sram_cell_6t_5 inst_cell_19_23 (.BL(BL23),.BLN(BLN23),.WL(WL19));
sram_cell_6t_5 inst_cell_19_24 (.BL(BL24),.BLN(BLN24),.WL(WL19));
sram_cell_6t_5 inst_cell_19_25 (.BL(BL25),.BLN(BLN25),.WL(WL19));
sram_cell_6t_5 inst_cell_19_26 (.BL(BL26),.BLN(BLN26),.WL(WL19));
sram_cell_6t_5 inst_cell_19_27 (.BL(BL27),.BLN(BLN27),.WL(WL19));
sram_cell_6t_5 inst_cell_19_28 (.BL(BL28),.BLN(BLN28),.WL(WL19));
sram_cell_6t_5 inst_cell_19_29 (.BL(BL29),.BLN(BLN29),.WL(WL19));
sram_cell_6t_5 inst_cell_19_30 (.BL(BL30),.BLN(BLN30),.WL(WL19));
sram_cell_6t_5 inst_cell_19_31 (.BL(BL31),.BLN(BLN31),.WL(WL19));
sram_cell_6t_5 inst_cell_19_32 (.BL(BL32),.BLN(BLN32),.WL(WL19));
sram_cell_6t_5 inst_cell_19_33 (.BL(BL33),.BLN(BLN33),.WL(WL19));
sram_cell_6t_5 inst_cell_19_34 (.BL(BL34),.BLN(BLN34),.WL(WL19));
sram_cell_6t_5 inst_cell_19_35 (.BL(BL35),.BLN(BLN35),.WL(WL19));
sram_cell_6t_5 inst_cell_19_36 (.BL(BL36),.BLN(BLN36),.WL(WL19));
sram_cell_6t_5 inst_cell_19_37 (.BL(BL37),.BLN(BLN37),.WL(WL19));
sram_cell_6t_5 inst_cell_19_38 (.BL(BL38),.BLN(BLN38),.WL(WL19));
sram_cell_6t_5 inst_cell_19_39 (.BL(BL39),.BLN(BLN39),.WL(WL19));
sram_cell_6t_5 inst_cell_19_40 (.BL(BL40),.BLN(BLN40),.WL(WL19));
sram_cell_6t_5 inst_cell_19_41 (.BL(BL41),.BLN(BLN41),.WL(WL19));
sram_cell_6t_5 inst_cell_19_42 (.BL(BL42),.BLN(BLN42),.WL(WL19));
sram_cell_6t_5 inst_cell_19_43 (.BL(BL43),.BLN(BLN43),.WL(WL19));
sram_cell_6t_5 inst_cell_19_44 (.BL(BL44),.BLN(BLN44),.WL(WL19));
sram_cell_6t_5 inst_cell_19_45 (.BL(BL45),.BLN(BLN45),.WL(WL19));
sram_cell_6t_5 inst_cell_19_46 (.BL(BL46),.BLN(BLN46),.WL(WL19));
sram_cell_6t_5 inst_cell_19_47 (.BL(BL47),.BLN(BLN47),.WL(WL19));
sram_cell_6t_5 inst_cell_19_48 (.BL(BL48),.BLN(BLN48),.WL(WL19));
sram_cell_6t_5 inst_cell_19_49 (.BL(BL49),.BLN(BLN49),.WL(WL19));
sram_cell_6t_5 inst_cell_19_50 (.BL(BL50),.BLN(BLN50),.WL(WL19));
sram_cell_6t_5 inst_cell_19_51 (.BL(BL51),.BLN(BLN51),.WL(WL19));
sram_cell_6t_5 inst_cell_19_52 (.BL(BL52),.BLN(BLN52),.WL(WL19));
sram_cell_6t_5 inst_cell_19_53 (.BL(BL53),.BLN(BLN53),.WL(WL19));
sram_cell_6t_5 inst_cell_19_54 (.BL(BL54),.BLN(BLN54),.WL(WL19));
sram_cell_6t_5 inst_cell_19_55 (.BL(BL55),.BLN(BLN55),.WL(WL19));
sram_cell_6t_5 inst_cell_19_56 (.BL(BL56),.BLN(BLN56),.WL(WL19));
sram_cell_6t_5 inst_cell_19_57 (.BL(BL57),.BLN(BLN57),.WL(WL19));
sram_cell_6t_5 inst_cell_19_58 (.BL(BL58),.BLN(BLN58),.WL(WL19));
sram_cell_6t_5 inst_cell_19_59 (.BL(BL59),.BLN(BLN59),.WL(WL19));
sram_cell_6t_5 inst_cell_19_60 (.BL(BL60),.BLN(BLN60),.WL(WL19));
sram_cell_6t_5 inst_cell_19_61 (.BL(BL61),.BLN(BLN61),.WL(WL19));
sram_cell_6t_5 inst_cell_19_62 (.BL(BL62),.BLN(BLN62),.WL(WL19));
sram_cell_6t_5 inst_cell_19_63 (.BL(BL63),.BLN(BLN63),.WL(WL19));
sram_cell_6t_5 inst_cell_19_64 (.BL(BL64),.BLN(BLN64),.WL(WL19));
sram_cell_6t_5 inst_cell_19_65 (.BL(BL65),.BLN(BLN65),.WL(WL19));
sram_cell_6t_5 inst_cell_19_66 (.BL(BL66),.BLN(BLN66),.WL(WL19));
sram_cell_6t_5 inst_cell_19_67 (.BL(BL67),.BLN(BLN67),.WL(WL19));
sram_cell_6t_5 inst_cell_19_68 (.BL(BL68),.BLN(BLN68),.WL(WL19));
sram_cell_6t_5 inst_cell_19_69 (.BL(BL69),.BLN(BLN69),.WL(WL19));
sram_cell_6t_5 inst_cell_19_70 (.BL(BL70),.BLN(BLN70),.WL(WL19));
sram_cell_6t_5 inst_cell_19_71 (.BL(BL71),.BLN(BLN71),.WL(WL19));
sram_cell_6t_5 inst_cell_19_72 (.BL(BL72),.BLN(BLN72),.WL(WL19));
sram_cell_6t_5 inst_cell_19_73 (.BL(BL73),.BLN(BLN73),.WL(WL19));
sram_cell_6t_5 inst_cell_19_74 (.BL(BL74),.BLN(BLN74),.WL(WL19));
sram_cell_6t_5 inst_cell_19_75 (.BL(BL75),.BLN(BLN75),.WL(WL19));
sram_cell_6t_5 inst_cell_19_76 (.BL(BL76),.BLN(BLN76),.WL(WL19));
sram_cell_6t_5 inst_cell_19_77 (.BL(BL77),.BLN(BLN77),.WL(WL19));
sram_cell_6t_5 inst_cell_19_78 (.BL(BL78),.BLN(BLN78),.WL(WL19));
sram_cell_6t_5 inst_cell_19_79 (.BL(BL79),.BLN(BLN79),.WL(WL19));
sram_cell_6t_5 inst_cell_19_80 (.BL(BL80),.BLN(BLN80),.WL(WL19));
sram_cell_6t_5 inst_cell_19_81 (.BL(BL81),.BLN(BLN81),.WL(WL19));
sram_cell_6t_5 inst_cell_19_82 (.BL(BL82),.BLN(BLN82),.WL(WL19));
sram_cell_6t_5 inst_cell_19_83 (.BL(BL83),.BLN(BLN83),.WL(WL19));
sram_cell_6t_5 inst_cell_19_84 (.BL(BL84),.BLN(BLN84),.WL(WL19));
sram_cell_6t_5 inst_cell_19_85 (.BL(BL85),.BLN(BLN85),.WL(WL19));
sram_cell_6t_5 inst_cell_19_86 (.BL(BL86),.BLN(BLN86),.WL(WL19));
sram_cell_6t_5 inst_cell_19_87 (.BL(BL87),.BLN(BLN87),.WL(WL19));
sram_cell_6t_5 inst_cell_19_88 (.BL(BL88),.BLN(BLN88),.WL(WL19));
sram_cell_6t_5 inst_cell_19_89 (.BL(BL89),.BLN(BLN89),.WL(WL19));
sram_cell_6t_5 inst_cell_19_90 (.BL(BL90),.BLN(BLN90),.WL(WL19));
sram_cell_6t_5 inst_cell_19_91 (.BL(BL91),.BLN(BLN91),.WL(WL19));
sram_cell_6t_5 inst_cell_19_92 (.BL(BL92),.BLN(BLN92),.WL(WL19));
sram_cell_6t_5 inst_cell_19_93 (.BL(BL93),.BLN(BLN93),.WL(WL19));
sram_cell_6t_5 inst_cell_19_94 (.BL(BL94),.BLN(BLN94),.WL(WL19));
sram_cell_6t_5 inst_cell_19_95 (.BL(BL95),.BLN(BLN95),.WL(WL19));
sram_cell_6t_5 inst_cell_19_96 (.BL(BL96),.BLN(BLN96),.WL(WL19));
sram_cell_6t_5 inst_cell_19_97 (.BL(BL97),.BLN(BLN97),.WL(WL19));
sram_cell_6t_5 inst_cell_19_98 (.BL(BL98),.BLN(BLN98),.WL(WL19));
sram_cell_6t_5 inst_cell_19_99 (.BL(BL99),.BLN(BLN99),.WL(WL19));
sram_cell_6t_5 inst_cell_19_100 (.BL(BL100),.BLN(BLN100),.WL(WL19));
sram_cell_6t_5 inst_cell_19_101 (.BL(BL101),.BLN(BLN101),.WL(WL19));
sram_cell_6t_5 inst_cell_19_102 (.BL(BL102),.BLN(BLN102),.WL(WL19));
sram_cell_6t_5 inst_cell_19_103 (.BL(BL103),.BLN(BLN103),.WL(WL19));
sram_cell_6t_5 inst_cell_19_104 (.BL(BL104),.BLN(BLN104),.WL(WL19));
sram_cell_6t_5 inst_cell_19_105 (.BL(BL105),.BLN(BLN105),.WL(WL19));
sram_cell_6t_5 inst_cell_19_106 (.BL(BL106),.BLN(BLN106),.WL(WL19));
sram_cell_6t_5 inst_cell_19_107 (.BL(BL107),.BLN(BLN107),.WL(WL19));
sram_cell_6t_5 inst_cell_19_108 (.BL(BL108),.BLN(BLN108),.WL(WL19));
sram_cell_6t_5 inst_cell_19_109 (.BL(BL109),.BLN(BLN109),.WL(WL19));
sram_cell_6t_5 inst_cell_19_110 (.BL(BL110),.BLN(BLN110),.WL(WL19));
sram_cell_6t_5 inst_cell_19_111 (.BL(BL111),.BLN(BLN111),.WL(WL19));
sram_cell_6t_5 inst_cell_19_112 (.BL(BL112),.BLN(BLN112),.WL(WL19));
sram_cell_6t_5 inst_cell_19_113 (.BL(BL113),.BLN(BLN113),.WL(WL19));
sram_cell_6t_5 inst_cell_19_114 (.BL(BL114),.BLN(BLN114),.WL(WL19));
sram_cell_6t_5 inst_cell_19_115 (.BL(BL115),.BLN(BLN115),.WL(WL19));
sram_cell_6t_5 inst_cell_19_116 (.BL(BL116),.BLN(BLN116),.WL(WL19));
sram_cell_6t_5 inst_cell_19_117 (.BL(BL117),.BLN(BLN117),.WL(WL19));
sram_cell_6t_5 inst_cell_19_118 (.BL(BL118),.BLN(BLN118),.WL(WL19));
sram_cell_6t_5 inst_cell_19_119 (.BL(BL119),.BLN(BLN119),.WL(WL19));
sram_cell_6t_5 inst_cell_19_120 (.BL(BL120),.BLN(BLN120),.WL(WL19));
sram_cell_6t_5 inst_cell_19_121 (.BL(BL121),.BLN(BLN121),.WL(WL19));
sram_cell_6t_5 inst_cell_19_122 (.BL(BL122),.BLN(BLN122),.WL(WL19));
sram_cell_6t_5 inst_cell_19_123 (.BL(BL123),.BLN(BLN123),.WL(WL19));
sram_cell_6t_5 inst_cell_19_124 (.BL(BL124),.BLN(BLN124),.WL(WL19));
sram_cell_6t_5 inst_cell_19_125 (.BL(BL125),.BLN(BLN125),.WL(WL19));
sram_cell_6t_5 inst_cell_19_126 (.BL(BL126),.BLN(BLN126),.WL(WL19));
sram_cell_6t_5 inst_cell_19_127 (.BL(BL127),.BLN(BLN127),.WL(WL19));
sram_cell_6t_5 inst_cell_20_0 (.BL(BL0),.BLN(BLN0),.WL(WL20));
sram_cell_6t_5 inst_cell_20_1 (.BL(BL1),.BLN(BLN1),.WL(WL20));
sram_cell_6t_5 inst_cell_20_2 (.BL(BL2),.BLN(BLN2),.WL(WL20));
sram_cell_6t_5 inst_cell_20_3 (.BL(BL3),.BLN(BLN3),.WL(WL20));
sram_cell_6t_5 inst_cell_20_4 (.BL(BL4),.BLN(BLN4),.WL(WL20));
sram_cell_6t_5 inst_cell_20_5 (.BL(BL5),.BLN(BLN5),.WL(WL20));
sram_cell_6t_5 inst_cell_20_6 (.BL(BL6),.BLN(BLN6),.WL(WL20));
sram_cell_6t_5 inst_cell_20_7 (.BL(BL7),.BLN(BLN7),.WL(WL20));
sram_cell_6t_5 inst_cell_20_8 (.BL(BL8),.BLN(BLN8),.WL(WL20));
sram_cell_6t_5 inst_cell_20_9 (.BL(BL9),.BLN(BLN9),.WL(WL20));
sram_cell_6t_5 inst_cell_20_10 (.BL(BL10),.BLN(BLN10),.WL(WL20));
sram_cell_6t_5 inst_cell_20_11 (.BL(BL11),.BLN(BLN11),.WL(WL20));
sram_cell_6t_5 inst_cell_20_12 (.BL(BL12),.BLN(BLN12),.WL(WL20));
sram_cell_6t_5 inst_cell_20_13 (.BL(BL13),.BLN(BLN13),.WL(WL20));
sram_cell_6t_5 inst_cell_20_14 (.BL(BL14),.BLN(BLN14),.WL(WL20));
sram_cell_6t_5 inst_cell_20_15 (.BL(BL15),.BLN(BLN15),.WL(WL20));
sram_cell_6t_5 inst_cell_20_16 (.BL(BL16),.BLN(BLN16),.WL(WL20));
sram_cell_6t_5 inst_cell_20_17 (.BL(BL17),.BLN(BLN17),.WL(WL20));
sram_cell_6t_5 inst_cell_20_18 (.BL(BL18),.BLN(BLN18),.WL(WL20));
sram_cell_6t_5 inst_cell_20_19 (.BL(BL19),.BLN(BLN19),.WL(WL20));
sram_cell_6t_5 inst_cell_20_20 (.BL(BL20),.BLN(BLN20),.WL(WL20));
sram_cell_6t_5 inst_cell_20_21 (.BL(BL21),.BLN(BLN21),.WL(WL20));
sram_cell_6t_5 inst_cell_20_22 (.BL(BL22),.BLN(BLN22),.WL(WL20));
sram_cell_6t_5 inst_cell_20_23 (.BL(BL23),.BLN(BLN23),.WL(WL20));
sram_cell_6t_5 inst_cell_20_24 (.BL(BL24),.BLN(BLN24),.WL(WL20));
sram_cell_6t_5 inst_cell_20_25 (.BL(BL25),.BLN(BLN25),.WL(WL20));
sram_cell_6t_5 inst_cell_20_26 (.BL(BL26),.BLN(BLN26),.WL(WL20));
sram_cell_6t_5 inst_cell_20_27 (.BL(BL27),.BLN(BLN27),.WL(WL20));
sram_cell_6t_5 inst_cell_20_28 (.BL(BL28),.BLN(BLN28),.WL(WL20));
sram_cell_6t_5 inst_cell_20_29 (.BL(BL29),.BLN(BLN29),.WL(WL20));
sram_cell_6t_5 inst_cell_20_30 (.BL(BL30),.BLN(BLN30),.WL(WL20));
sram_cell_6t_5 inst_cell_20_31 (.BL(BL31),.BLN(BLN31),.WL(WL20));
sram_cell_6t_5 inst_cell_20_32 (.BL(BL32),.BLN(BLN32),.WL(WL20));
sram_cell_6t_5 inst_cell_20_33 (.BL(BL33),.BLN(BLN33),.WL(WL20));
sram_cell_6t_5 inst_cell_20_34 (.BL(BL34),.BLN(BLN34),.WL(WL20));
sram_cell_6t_5 inst_cell_20_35 (.BL(BL35),.BLN(BLN35),.WL(WL20));
sram_cell_6t_5 inst_cell_20_36 (.BL(BL36),.BLN(BLN36),.WL(WL20));
sram_cell_6t_5 inst_cell_20_37 (.BL(BL37),.BLN(BLN37),.WL(WL20));
sram_cell_6t_5 inst_cell_20_38 (.BL(BL38),.BLN(BLN38),.WL(WL20));
sram_cell_6t_5 inst_cell_20_39 (.BL(BL39),.BLN(BLN39),.WL(WL20));
sram_cell_6t_5 inst_cell_20_40 (.BL(BL40),.BLN(BLN40),.WL(WL20));
sram_cell_6t_5 inst_cell_20_41 (.BL(BL41),.BLN(BLN41),.WL(WL20));
sram_cell_6t_5 inst_cell_20_42 (.BL(BL42),.BLN(BLN42),.WL(WL20));
sram_cell_6t_5 inst_cell_20_43 (.BL(BL43),.BLN(BLN43),.WL(WL20));
sram_cell_6t_5 inst_cell_20_44 (.BL(BL44),.BLN(BLN44),.WL(WL20));
sram_cell_6t_5 inst_cell_20_45 (.BL(BL45),.BLN(BLN45),.WL(WL20));
sram_cell_6t_5 inst_cell_20_46 (.BL(BL46),.BLN(BLN46),.WL(WL20));
sram_cell_6t_5 inst_cell_20_47 (.BL(BL47),.BLN(BLN47),.WL(WL20));
sram_cell_6t_5 inst_cell_20_48 (.BL(BL48),.BLN(BLN48),.WL(WL20));
sram_cell_6t_5 inst_cell_20_49 (.BL(BL49),.BLN(BLN49),.WL(WL20));
sram_cell_6t_5 inst_cell_20_50 (.BL(BL50),.BLN(BLN50),.WL(WL20));
sram_cell_6t_5 inst_cell_20_51 (.BL(BL51),.BLN(BLN51),.WL(WL20));
sram_cell_6t_5 inst_cell_20_52 (.BL(BL52),.BLN(BLN52),.WL(WL20));
sram_cell_6t_5 inst_cell_20_53 (.BL(BL53),.BLN(BLN53),.WL(WL20));
sram_cell_6t_5 inst_cell_20_54 (.BL(BL54),.BLN(BLN54),.WL(WL20));
sram_cell_6t_5 inst_cell_20_55 (.BL(BL55),.BLN(BLN55),.WL(WL20));
sram_cell_6t_5 inst_cell_20_56 (.BL(BL56),.BLN(BLN56),.WL(WL20));
sram_cell_6t_5 inst_cell_20_57 (.BL(BL57),.BLN(BLN57),.WL(WL20));
sram_cell_6t_5 inst_cell_20_58 (.BL(BL58),.BLN(BLN58),.WL(WL20));
sram_cell_6t_5 inst_cell_20_59 (.BL(BL59),.BLN(BLN59),.WL(WL20));
sram_cell_6t_5 inst_cell_20_60 (.BL(BL60),.BLN(BLN60),.WL(WL20));
sram_cell_6t_5 inst_cell_20_61 (.BL(BL61),.BLN(BLN61),.WL(WL20));
sram_cell_6t_5 inst_cell_20_62 (.BL(BL62),.BLN(BLN62),.WL(WL20));
sram_cell_6t_5 inst_cell_20_63 (.BL(BL63),.BLN(BLN63),.WL(WL20));
sram_cell_6t_5 inst_cell_20_64 (.BL(BL64),.BLN(BLN64),.WL(WL20));
sram_cell_6t_5 inst_cell_20_65 (.BL(BL65),.BLN(BLN65),.WL(WL20));
sram_cell_6t_5 inst_cell_20_66 (.BL(BL66),.BLN(BLN66),.WL(WL20));
sram_cell_6t_5 inst_cell_20_67 (.BL(BL67),.BLN(BLN67),.WL(WL20));
sram_cell_6t_5 inst_cell_20_68 (.BL(BL68),.BLN(BLN68),.WL(WL20));
sram_cell_6t_5 inst_cell_20_69 (.BL(BL69),.BLN(BLN69),.WL(WL20));
sram_cell_6t_5 inst_cell_20_70 (.BL(BL70),.BLN(BLN70),.WL(WL20));
sram_cell_6t_5 inst_cell_20_71 (.BL(BL71),.BLN(BLN71),.WL(WL20));
sram_cell_6t_5 inst_cell_20_72 (.BL(BL72),.BLN(BLN72),.WL(WL20));
sram_cell_6t_5 inst_cell_20_73 (.BL(BL73),.BLN(BLN73),.WL(WL20));
sram_cell_6t_5 inst_cell_20_74 (.BL(BL74),.BLN(BLN74),.WL(WL20));
sram_cell_6t_5 inst_cell_20_75 (.BL(BL75),.BLN(BLN75),.WL(WL20));
sram_cell_6t_5 inst_cell_20_76 (.BL(BL76),.BLN(BLN76),.WL(WL20));
sram_cell_6t_5 inst_cell_20_77 (.BL(BL77),.BLN(BLN77),.WL(WL20));
sram_cell_6t_5 inst_cell_20_78 (.BL(BL78),.BLN(BLN78),.WL(WL20));
sram_cell_6t_5 inst_cell_20_79 (.BL(BL79),.BLN(BLN79),.WL(WL20));
sram_cell_6t_5 inst_cell_20_80 (.BL(BL80),.BLN(BLN80),.WL(WL20));
sram_cell_6t_5 inst_cell_20_81 (.BL(BL81),.BLN(BLN81),.WL(WL20));
sram_cell_6t_5 inst_cell_20_82 (.BL(BL82),.BLN(BLN82),.WL(WL20));
sram_cell_6t_5 inst_cell_20_83 (.BL(BL83),.BLN(BLN83),.WL(WL20));
sram_cell_6t_5 inst_cell_20_84 (.BL(BL84),.BLN(BLN84),.WL(WL20));
sram_cell_6t_5 inst_cell_20_85 (.BL(BL85),.BLN(BLN85),.WL(WL20));
sram_cell_6t_5 inst_cell_20_86 (.BL(BL86),.BLN(BLN86),.WL(WL20));
sram_cell_6t_5 inst_cell_20_87 (.BL(BL87),.BLN(BLN87),.WL(WL20));
sram_cell_6t_5 inst_cell_20_88 (.BL(BL88),.BLN(BLN88),.WL(WL20));
sram_cell_6t_5 inst_cell_20_89 (.BL(BL89),.BLN(BLN89),.WL(WL20));
sram_cell_6t_5 inst_cell_20_90 (.BL(BL90),.BLN(BLN90),.WL(WL20));
sram_cell_6t_5 inst_cell_20_91 (.BL(BL91),.BLN(BLN91),.WL(WL20));
sram_cell_6t_5 inst_cell_20_92 (.BL(BL92),.BLN(BLN92),.WL(WL20));
sram_cell_6t_5 inst_cell_20_93 (.BL(BL93),.BLN(BLN93),.WL(WL20));
sram_cell_6t_5 inst_cell_20_94 (.BL(BL94),.BLN(BLN94),.WL(WL20));
sram_cell_6t_5 inst_cell_20_95 (.BL(BL95),.BLN(BLN95),.WL(WL20));
sram_cell_6t_5 inst_cell_20_96 (.BL(BL96),.BLN(BLN96),.WL(WL20));
sram_cell_6t_5 inst_cell_20_97 (.BL(BL97),.BLN(BLN97),.WL(WL20));
sram_cell_6t_5 inst_cell_20_98 (.BL(BL98),.BLN(BLN98),.WL(WL20));
sram_cell_6t_5 inst_cell_20_99 (.BL(BL99),.BLN(BLN99),.WL(WL20));
sram_cell_6t_5 inst_cell_20_100 (.BL(BL100),.BLN(BLN100),.WL(WL20));
sram_cell_6t_5 inst_cell_20_101 (.BL(BL101),.BLN(BLN101),.WL(WL20));
sram_cell_6t_5 inst_cell_20_102 (.BL(BL102),.BLN(BLN102),.WL(WL20));
sram_cell_6t_5 inst_cell_20_103 (.BL(BL103),.BLN(BLN103),.WL(WL20));
sram_cell_6t_5 inst_cell_20_104 (.BL(BL104),.BLN(BLN104),.WL(WL20));
sram_cell_6t_5 inst_cell_20_105 (.BL(BL105),.BLN(BLN105),.WL(WL20));
sram_cell_6t_5 inst_cell_20_106 (.BL(BL106),.BLN(BLN106),.WL(WL20));
sram_cell_6t_5 inst_cell_20_107 (.BL(BL107),.BLN(BLN107),.WL(WL20));
sram_cell_6t_5 inst_cell_20_108 (.BL(BL108),.BLN(BLN108),.WL(WL20));
sram_cell_6t_5 inst_cell_20_109 (.BL(BL109),.BLN(BLN109),.WL(WL20));
sram_cell_6t_5 inst_cell_20_110 (.BL(BL110),.BLN(BLN110),.WL(WL20));
sram_cell_6t_5 inst_cell_20_111 (.BL(BL111),.BLN(BLN111),.WL(WL20));
sram_cell_6t_5 inst_cell_20_112 (.BL(BL112),.BLN(BLN112),.WL(WL20));
sram_cell_6t_5 inst_cell_20_113 (.BL(BL113),.BLN(BLN113),.WL(WL20));
sram_cell_6t_5 inst_cell_20_114 (.BL(BL114),.BLN(BLN114),.WL(WL20));
sram_cell_6t_5 inst_cell_20_115 (.BL(BL115),.BLN(BLN115),.WL(WL20));
sram_cell_6t_5 inst_cell_20_116 (.BL(BL116),.BLN(BLN116),.WL(WL20));
sram_cell_6t_5 inst_cell_20_117 (.BL(BL117),.BLN(BLN117),.WL(WL20));
sram_cell_6t_5 inst_cell_20_118 (.BL(BL118),.BLN(BLN118),.WL(WL20));
sram_cell_6t_5 inst_cell_20_119 (.BL(BL119),.BLN(BLN119),.WL(WL20));
sram_cell_6t_5 inst_cell_20_120 (.BL(BL120),.BLN(BLN120),.WL(WL20));
sram_cell_6t_5 inst_cell_20_121 (.BL(BL121),.BLN(BLN121),.WL(WL20));
sram_cell_6t_5 inst_cell_20_122 (.BL(BL122),.BLN(BLN122),.WL(WL20));
sram_cell_6t_5 inst_cell_20_123 (.BL(BL123),.BLN(BLN123),.WL(WL20));
sram_cell_6t_5 inst_cell_20_124 (.BL(BL124),.BLN(BLN124),.WL(WL20));
sram_cell_6t_5 inst_cell_20_125 (.BL(BL125),.BLN(BLN125),.WL(WL20));
sram_cell_6t_5 inst_cell_20_126 (.BL(BL126),.BLN(BLN126),.WL(WL20));
sram_cell_6t_5 inst_cell_20_127 (.BL(BL127),.BLN(BLN127),.WL(WL20));
sram_cell_6t_5 inst_cell_21_0 (.BL(BL0),.BLN(BLN0),.WL(WL21));
sram_cell_6t_5 inst_cell_21_1 (.BL(BL1),.BLN(BLN1),.WL(WL21));
sram_cell_6t_5 inst_cell_21_2 (.BL(BL2),.BLN(BLN2),.WL(WL21));
sram_cell_6t_5 inst_cell_21_3 (.BL(BL3),.BLN(BLN3),.WL(WL21));
sram_cell_6t_5 inst_cell_21_4 (.BL(BL4),.BLN(BLN4),.WL(WL21));
sram_cell_6t_5 inst_cell_21_5 (.BL(BL5),.BLN(BLN5),.WL(WL21));
sram_cell_6t_5 inst_cell_21_6 (.BL(BL6),.BLN(BLN6),.WL(WL21));
sram_cell_6t_5 inst_cell_21_7 (.BL(BL7),.BLN(BLN7),.WL(WL21));
sram_cell_6t_5 inst_cell_21_8 (.BL(BL8),.BLN(BLN8),.WL(WL21));
sram_cell_6t_5 inst_cell_21_9 (.BL(BL9),.BLN(BLN9),.WL(WL21));
sram_cell_6t_5 inst_cell_21_10 (.BL(BL10),.BLN(BLN10),.WL(WL21));
sram_cell_6t_5 inst_cell_21_11 (.BL(BL11),.BLN(BLN11),.WL(WL21));
sram_cell_6t_5 inst_cell_21_12 (.BL(BL12),.BLN(BLN12),.WL(WL21));
sram_cell_6t_5 inst_cell_21_13 (.BL(BL13),.BLN(BLN13),.WL(WL21));
sram_cell_6t_5 inst_cell_21_14 (.BL(BL14),.BLN(BLN14),.WL(WL21));
sram_cell_6t_5 inst_cell_21_15 (.BL(BL15),.BLN(BLN15),.WL(WL21));
sram_cell_6t_5 inst_cell_21_16 (.BL(BL16),.BLN(BLN16),.WL(WL21));
sram_cell_6t_5 inst_cell_21_17 (.BL(BL17),.BLN(BLN17),.WL(WL21));
sram_cell_6t_5 inst_cell_21_18 (.BL(BL18),.BLN(BLN18),.WL(WL21));
sram_cell_6t_5 inst_cell_21_19 (.BL(BL19),.BLN(BLN19),.WL(WL21));
sram_cell_6t_5 inst_cell_21_20 (.BL(BL20),.BLN(BLN20),.WL(WL21));
sram_cell_6t_5 inst_cell_21_21 (.BL(BL21),.BLN(BLN21),.WL(WL21));
sram_cell_6t_5 inst_cell_21_22 (.BL(BL22),.BLN(BLN22),.WL(WL21));
sram_cell_6t_5 inst_cell_21_23 (.BL(BL23),.BLN(BLN23),.WL(WL21));
sram_cell_6t_5 inst_cell_21_24 (.BL(BL24),.BLN(BLN24),.WL(WL21));
sram_cell_6t_5 inst_cell_21_25 (.BL(BL25),.BLN(BLN25),.WL(WL21));
sram_cell_6t_5 inst_cell_21_26 (.BL(BL26),.BLN(BLN26),.WL(WL21));
sram_cell_6t_5 inst_cell_21_27 (.BL(BL27),.BLN(BLN27),.WL(WL21));
sram_cell_6t_5 inst_cell_21_28 (.BL(BL28),.BLN(BLN28),.WL(WL21));
sram_cell_6t_5 inst_cell_21_29 (.BL(BL29),.BLN(BLN29),.WL(WL21));
sram_cell_6t_5 inst_cell_21_30 (.BL(BL30),.BLN(BLN30),.WL(WL21));
sram_cell_6t_5 inst_cell_21_31 (.BL(BL31),.BLN(BLN31),.WL(WL21));
sram_cell_6t_5 inst_cell_21_32 (.BL(BL32),.BLN(BLN32),.WL(WL21));
sram_cell_6t_5 inst_cell_21_33 (.BL(BL33),.BLN(BLN33),.WL(WL21));
sram_cell_6t_5 inst_cell_21_34 (.BL(BL34),.BLN(BLN34),.WL(WL21));
sram_cell_6t_5 inst_cell_21_35 (.BL(BL35),.BLN(BLN35),.WL(WL21));
sram_cell_6t_5 inst_cell_21_36 (.BL(BL36),.BLN(BLN36),.WL(WL21));
sram_cell_6t_5 inst_cell_21_37 (.BL(BL37),.BLN(BLN37),.WL(WL21));
sram_cell_6t_5 inst_cell_21_38 (.BL(BL38),.BLN(BLN38),.WL(WL21));
sram_cell_6t_5 inst_cell_21_39 (.BL(BL39),.BLN(BLN39),.WL(WL21));
sram_cell_6t_5 inst_cell_21_40 (.BL(BL40),.BLN(BLN40),.WL(WL21));
sram_cell_6t_5 inst_cell_21_41 (.BL(BL41),.BLN(BLN41),.WL(WL21));
sram_cell_6t_5 inst_cell_21_42 (.BL(BL42),.BLN(BLN42),.WL(WL21));
sram_cell_6t_5 inst_cell_21_43 (.BL(BL43),.BLN(BLN43),.WL(WL21));
sram_cell_6t_5 inst_cell_21_44 (.BL(BL44),.BLN(BLN44),.WL(WL21));
sram_cell_6t_5 inst_cell_21_45 (.BL(BL45),.BLN(BLN45),.WL(WL21));
sram_cell_6t_5 inst_cell_21_46 (.BL(BL46),.BLN(BLN46),.WL(WL21));
sram_cell_6t_5 inst_cell_21_47 (.BL(BL47),.BLN(BLN47),.WL(WL21));
sram_cell_6t_5 inst_cell_21_48 (.BL(BL48),.BLN(BLN48),.WL(WL21));
sram_cell_6t_5 inst_cell_21_49 (.BL(BL49),.BLN(BLN49),.WL(WL21));
sram_cell_6t_5 inst_cell_21_50 (.BL(BL50),.BLN(BLN50),.WL(WL21));
sram_cell_6t_5 inst_cell_21_51 (.BL(BL51),.BLN(BLN51),.WL(WL21));
sram_cell_6t_5 inst_cell_21_52 (.BL(BL52),.BLN(BLN52),.WL(WL21));
sram_cell_6t_5 inst_cell_21_53 (.BL(BL53),.BLN(BLN53),.WL(WL21));
sram_cell_6t_5 inst_cell_21_54 (.BL(BL54),.BLN(BLN54),.WL(WL21));
sram_cell_6t_5 inst_cell_21_55 (.BL(BL55),.BLN(BLN55),.WL(WL21));
sram_cell_6t_5 inst_cell_21_56 (.BL(BL56),.BLN(BLN56),.WL(WL21));
sram_cell_6t_5 inst_cell_21_57 (.BL(BL57),.BLN(BLN57),.WL(WL21));
sram_cell_6t_5 inst_cell_21_58 (.BL(BL58),.BLN(BLN58),.WL(WL21));
sram_cell_6t_5 inst_cell_21_59 (.BL(BL59),.BLN(BLN59),.WL(WL21));
sram_cell_6t_5 inst_cell_21_60 (.BL(BL60),.BLN(BLN60),.WL(WL21));
sram_cell_6t_5 inst_cell_21_61 (.BL(BL61),.BLN(BLN61),.WL(WL21));
sram_cell_6t_5 inst_cell_21_62 (.BL(BL62),.BLN(BLN62),.WL(WL21));
sram_cell_6t_5 inst_cell_21_63 (.BL(BL63),.BLN(BLN63),.WL(WL21));
sram_cell_6t_5 inst_cell_21_64 (.BL(BL64),.BLN(BLN64),.WL(WL21));
sram_cell_6t_5 inst_cell_21_65 (.BL(BL65),.BLN(BLN65),.WL(WL21));
sram_cell_6t_5 inst_cell_21_66 (.BL(BL66),.BLN(BLN66),.WL(WL21));
sram_cell_6t_5 inst_cell_21_67 (.BL(BL67),.BLN(BLN67),.WL(WL21));
sram_cell_6t_5 inst_cell_21_68 (.BL(BL68),.BLN(BLN68),.WL(WL21));
sram_cell_6t_5 inst_cell_21_69 (.BL(BL69),.BLN(BLN69),.WL(WL21));
sram_cell_6t_5 inst_cell_21_70 (.BL(BL70),.BLN(BLN70),.WL(WL21));
sram_cell_6t_5 inst_cell_21_71 (.BL(BL71),.BLN(BLN71),.WL(WL21));
sram_cell_6t_5 inst_cell_21_72 (.BL(BL72),.BLN(BLN72),.WL(WL21));
sram_cell_6t_5 inst_cell_21_73 (.BL(BL73),.BLN(BLN73),.WL(WL21));
sram_cell_6t_5 inst_cell_21_74 (.BL(BL74),.BLN(BLN74),.WL(WL21));
sram_cell_6t_5 inst_cell_21_75 (.BL(BL75),.BLN(BLN75),.WL(WL21));
sram_cell_6t_5 inst_cell_21_76 (.BL(BL76),.BLN(BLN76),.WL(WL21));
sram_cell_6t_5 inst_cell_21_77 (.BL(BL77),.BLN(BLN77),.WL(WL21));
sram_cell_6t_5 inst_cell_21_78 (.BL(BL78),.BLN(BLN78),.WL(WL21));
sram_cell_6t_5 inst_cell_21_79 (.BL(BL79),.BLN(BLN79),.WL(WL21));
sram_cell_6t_5 inst_cell_21_80 (.BL(BL80),.BLN(BLN80),.WL(WL21));
sram_cell_6t_5 inst_cell_21_81 (.BL(BL81),.BLN(BLN81),.WL(WL21));
sram_cell_6t_5 inst_cell_21_82 (.BL(BL82),.BLN(BLN82),.WL(WL21));
sram_cell_6t_5 inst_cell_21_83 (.BL(BL83),.BLN(BLN83),.WL(WL21));
sram_cell_6t_5 inst_cell_21_84 (.BL(BL84),.BLN(BLN84),.WL(WL21));
sram_cell_6t_5 inst_cell_21_85 (.BL(BL85),.BLN(BLN85),.WL(WL21));
sram_cell_6t_5 inst_cell_21_86 (.BL(BL86),.BLN(BLN86),.WL(WL21));
sram_cell_6t_5 inst_cell_21_87 (.BL(BL87),.BLN(BLN87),.WL(WL21));
sram_cell_6t_5 inst_cell_21_88 (.BL(BL88),.BLN(BLN88),.WL(WL21));
sram_cell_6t_5 inst_cell_21_89 (.BL(BL89),.BLN(BLN89),.WL(WL21));
sram_cell_6t_5 inst_cell_21_90 (.BL(BL90),.BLN(BLN90),.WL(WL21));
sram_cell_6t_5 inst_cell_21_91 (.BL(BL91),.BLN(BLN91),.WL(WL21));
sram_cell_6t_5 inst_cell_21_92 (.BL(BL92),.BLN(BLN92),.WL(WL21));
sram_cell_6t_5 inst_cell_21_93 (.BL(BL93),.BLN(BLN93),.WL(WL21));
sram_cell_6t_5 inst_cell_21_94 (.BL(BL94),.BLN(BLN94),.WL(WL21));
sram_cell_6t_5 inst_cell_21_95 (.BL(BL95),.BLN(BLN95),.WL(WL21));
sram_cell_6t_5 inst_cell_21_96 (.BL(BL96),.BLN(BLN96),.WL(WL21));
sram_cell_6t_5 inst_cell_21_97 (.BL(BL97),.BLN(BLN97),.WL(WL21));
sram_cell_6t_5 inst_cell_21_98 (.BL(BL98),.BLN(BLN98),.WL(WL21));
sram_cell_6t_5 inst_cell_21_99 (.BL(BL99),.BLN(BLN99),.WL(WL21));
sram_cell_6t_5 inst_cell_21_100 (.BL(BL100),.BLN(BLN100),.WL(WL21));
sram_cell_6t_5 inst_cell_21_101 (.BL(BL101),.BLN(BLN101),.WL(WL21));
sram_cell_6t_5 inst_cell_21_102 (.BL(BL102),.BLN(BLN102),.WL(WL21));
sram_cell_6t_5 inst_cell_21_103 (.BL(BL103),.BLN(BLN103),.WL(WL21));
sram_cell_6t_5 inst_cell_21_104 (.BL(BL104),.BLN(BLN104),.WL(WL21));
sram_cell_6t_5 inst_cell_21_105 (.BL(BL105),.BLN(BLN105),.WL(WL21));
sram_cell_6t_5 inst_cell_21_106 (.BL(BL106),.BLN(BLN106),.WL(WL21));
sram_cell_6t_5 inst_cell_21_107 (.BL(BL107),.BLN(BLN107),.WL(WL21));
sram_cell_6t_5 inst_cell_21_108 (.BL(BL108),.BLN(BLN108),.WL(WL21));
sram_cell_6t_5 inst_cell_21_109 (.BL(BL109),.BLN(BLN109),.WL(WL21));
sram_cell_6t_5 inst_cell_21_110 (.BL(BL110),.BLN(BLN110),.WL(WL21));
sram_cell_6t_5 inst_cell_21_111 (.BL(BL111),.BLN(BLN111),.WL(WL21));
sram_cell_6t_5 inst_cell_21_112 (.BL(BL112),.BLN(BLN112),.WL(WL21));
sram_cell_6t_5 inst_cell_21_113 (.BL(BL113),.BLN(BLN113),.WL(WL21));
sram_cell_6t_5 inst_cell_21_114 (.BL(BL114),.BLN(BLN114),.WL(WL21));
sram_cell_6t_5 inst_cell_21_115 (.BL(BL115),.BLN(BLN115),.WL(WL21));
sram_cell_6t_5 inst_cell_21_116 (.BL(BL116),.BLN(BLN116),.WL(WL21));
sram_cell_6t_5 inst_cell_21_117 (.BL(BL117),.BLN(BLN117),.WL(WL21));
sram_cell_6t_5 inst_cell_21_118 (.BL(BL118),.BLN(BLN118),.WL(WL21));
sram_cell_6t_5 inst_cell_21_119 (.BL(BL119),.BLN(BLN119),.WL(WL21));
sram_cell_6t_5 inst_cell_21_120 (.BL(BL120),.BLN(BLN120),.WL(WL21));
sram_cell_6t_5 inst_cell_21_121 (.BL(BL121),.BLN(BLN121),.WL(WL21));
sram_cell_6t_5 inst_cell_21_122 (.BL(BL122),.BLN(BLN122),.WL(WL21));
sram_cell_6t_5 inst_cell_21_123 (.BL(BL123),.BLN(BLN123),.WL(WL21));
sram_cell_6t_5 inst_cell_21_124 (.BL(BL124),.BLN(BLN124),.WL(WL21));
sram_cell_6t_5 inst_cell_21_125 (.BL(BL125),.BLN(BLN125),.WL(WL21));
sram_cell_6t_5 inst_cell_21_126 (.BL(BL126),.BLN(BLN126),.WL(WL21));
sram_cell_6t_5 inst_cell_21_127 (.BL(BL127),.BLN(BLN127),.WL(WL21));
sram_cell_6t_5 inst_cell_22_0 (.BL(BL0),.BLN(BLN0),.WL(WL22));
sram_cell_6t_5 inst_cell_22_1 (.BL(BL1),.BLN(BLN1),.WL(WL22));
sram_cell_6t_5 inst_cell_22_2 (.BL(BL2),.BLN(BLN2),.WL(WL22));
sram_cell_6t_5 inst_cell_22_3 (.BL(BL3),.BLN(BLN3),.WL(WL22));
sram_cell_6t_5 inst_cell_22_4 (.BL(BL4),.BLN(BLN4),.WL(WL22));
sram_cell_6t_5 inst_cell_22_5 (.BL(BL5),.BLN(BLN5),.WL(WL22));
sram_cell_6t_5 inst_cell_22_6 (.BL(BL6),.BLN(BLN6),.WL(WL22));
sram_cell_6t_5 inst_cell_22_7 (.BL(BL7),.BLN(BLN7),.WL(WL22));
sram_cell_6t_5 inst_cell_22_8 (.BL(BL8),.BLN(BLN8),.WL(WL22));
sram_cell_6t_5 inst_cell_22_9 (.BL(BL9),.BLN(BLN9),.WL(WL22));
sram_cell_6t_5 inst_cell_22_10 (.BL(BL10),.BLN(BLN10),.WL(WL22));
sram_cell_6t_5 inst_cell_22_11 (.BL(BL11),.BLN(BLN11),.WL(WL22));
sram_cell_6t_5 inst_cell_22_12 (.BL(BL12),.BLN(BLN12),.WL(WL22));
sram_cell_6t_5 inst_cell_22_13 (.BL(BL13),.BLN(BLN13),.WL(WL22));
sram_cell_6t_5 inst_cell_22_14 (.BL(BL14),.BLN(BLN14),.WL(WL22));
sram_cell_6t_5 inst_cell_22_15 (.BL(BL15),.BLN(BLN15),.WL(WL22));
sram_cell_6t_5 inst_cell_22_16 (.BL(BL16),.BLN(BLN16),.WL(WL22));
sram_cell_6t_5 inst_cell_22_17 (.BL(BL17),.BLN(BLN17),.WL(WL22));
sram_cell_6t_5 inst_cell_22_18 (.BL(BL18),.BLN(BLN18),.WL(WL22));
sram_cell_6t_5 inst_cell_22_19 (.BL(BL19),.BLN(BLN19),.WL(WL22));
sram_cell_6t_5 inst_cell_22_20 (.BL(BL20),.BLN(BLN20),.WL(WL22));
sram_cell_6t_5 inst_cell_22_21 (.BL(BL21),.BLN(BLN21),.WL(WL22));
sram_cell_6t_5 inst_cell_22_22 (.BL(BL22),.BLN(BLN22),.WL(WL22));
sram_cell_6t_5 inst_cell_22_23 (.BL(BL23),.BLN(BLN23),.WL(WL22));
sram_cell_6t_5 inst_cell_22_24 (.BL(BL24),.BLN(BLN24),.WL(WL22));
sram_cell_6t_5 inst_cell_22_25 (.BL(BL25),.BLN(BLN25),.WL(WL22));
sram_cell_6t_5 inst_cell_22_26 (.BL(BL26),.BLN(BLN26),.WL(WL22));
sram_cell_6t_5 inst_cell_22_27 (.BL(BL27),.BLN(BLN27),.WL(WL22));
sram_cell_6t_5 inst_cell_22_28 (.BL(BL28),.BLN(BLN28),.WL(WL22));
sram_cell_6t_5 inst_cell_22_29 (.BL(BL29),.BLN(BLN29),.WL(WL22));
sram_cell_6t_5 inst_cell_22_30 (.BL(BL30),.BLN(BLN30),.WL(WL22));
sram_cell_6t_5 inst_cell_22_31 (.BL(BL31),.BLN(BLN31),.WL(WL22));
sram_cell_6t_5 inst_cell_22_32 (.BL(BL32),.BLN(BLN32),.WL(WL22));
sram_cell_6t_5 inst_cell_22_33 (.BL(BL33),.BLN(BLN33),.WL(WL22));
sram_cell_6t_5 inst_cell_22_34 (.BL(BL34),.BLN(BLN34),.WL(WL22));
sram_cell_6t_5 inst_cell_22_35 (.BL(BL35),.BLN(BLN35),.WL(WL22));
sram_cell_6t_5 inst_cell_22_36 (.BL(BL36),.BLN(BLN36),.WL(WL22));
sram_cell_6t_5 inst_cell_22_37 (.BL(BL37),.BLN(BLN37),.WL(WL22));
sram_cell_6t_5 inst_cell_22_38 (.BL(BL38),.BLN(BLN38),.WL(WL22));
sram_cell_6t_5 inst_cell_22_39 (.BL(BL39),.BLN(BLN39),.WL(WL22));
sram_cell_6t_5 inst_cell_22_40 (.BL(BL40),.BLN(BLN40),.WL(WL22));
sram_cell_6t_5 inst_cell_22_41 (.BL(BL41),.BLN(BLN41),.WL(WL22));
sram_cell_6t_5 inst_cell_22_42 (.BL(BL42),.BLN(BLN42),.WL(WL22));
sram_cell_6t_5 inst_cell_22_43 (.BL(BL43),.BLN(BLN43),.WL(WL22));
sram_cell_6t_5 inst_cell_22_44 (.BL(BL44),.BLN(BLN44),.WL(WL22));
sram_cell_6t_5 inst_cell_22_45 (.BL(BL45),.BLN(BLN45),.WL(WL22));
sram_cell_6t_5 inst_cell_22_46 (.BL(BL46),.BLN(BLN46),.WL(WL22));
sram_cell_6t_5 inst_cell_22_47 (.BL(BL47),.BLN(BLN47),.WL(WL22));
sram_cell_6t_5 inst_cell_22_48 (.BL(BL48),.BLN(BLN48),.WL(WL22));
sram_cell_6t_5 inst_cell_22_49 (.BL(BL49),.BLN(BLN49),.WL(WL22));
sram_cell_6t_5 inst_cell_22_50 (.BL(BL50),.BLN(BLN50),.WL(WL22));
sram_cell_6t_5 inst_cell_22_51 (.BL(BL51),.BLN(BLN51),.WL(WL22));
sram_cell_6t_5 inst_cell_22_52 (.BL(BL52),.BLN(BLN52),.WL(WL22));
sram_cell_6t_5 inst_cell_22_53 (.BL(BL53),.BLN(BLN53),.WL(WL22));
sram_cell_6t_5 inst_cell_22_54 (.BL(BL54),.BLN(BLN54),.WL(WL22));
sram_cell_6t_5 inst_cell_22_55 (.BL(BL55),.BLN(BLN55),.WL(WL22));
sram_cell_6t_5 inst_cell_22_56 (.BL(BL56),.BLN(BLN56),.WL(WL22));
sram_cell_6t_5 inst_cell_22_57 (.BL(BL57),.BLN(BLN57),.WL(WL22));
sram_cell_6t_5 inst_cell_22_58 (.BL(BL58),.BLN(BLN58),.WL(WL22));
sram_cell_6t_5 inst_cell_22_59 (.BL(BL59),.BLN(BLN59),.WL(WL22));
sram_cell_6t_5 inst_cell_22_60 (.BL(BL60),.BLN(BLN60),.WL(WL22));
sram_cell_6t_5 inst_cell_22_61 (.BL(BL61),.BLN(BLN61),.WL(WL22));
sram_cell_6t_5 inst_cell_22_62 (.BL(BL62),.BLN(BLN62),.WL(WL22));
sram_cell_6t_5 inst_cell_22_63 (.BL(BL63),.BLN(BLN63),.WL(WL22));
sram_cell_6t_5 inst_cell_22_64 (.BL(BL64),.BLN(BLN64),.WL(WL22));
sram_cell_6t_5 inst_cell_22_65 (.BL(BL65),.BLN(BLN65),.WL(WL22));
sram_cell_6t_5 inst_cell_22_66 (.BL(BL66),.BLN(BLN66),.WL(WL22));
sram_cell_6t_5 inst_cell_22_67 (.BL(BL67),.BLN(BLN67),.WL(WL22));
sram_cell_6t_5 inst_cell_22_68 (.BL(BL68),.BLN(BLN68),.WL(WL22));
sram_cell_6t_5 inst_cell_22_69 (.BL(BL69),.BLN(BLN69),.WL(WL22));
sram_cell_6t_5 inst_cell_22_70 (.BL(BL70),.BLN(BLN70),.WL(WL22));
sram_cell_6t_5 inst_cell_22_71 (.BL(BL71),.BLN(BLN71),.WL(WL22));
sram_cell_6t_5 inst_cell_22_72 (.BL(BL72),.BLN(BLN72),.WL(WL22));
sram_cell_6t_5 inst_cell_22_73 (.BL(BL73),.BLN(BLN73),.WL(WL22));
sram_cell_6t_5 inst_cell_22_74 (.BL(BL74),.BLN(BLN74),.WL(WL22));
sram_cell_6t_5 inst_cell_22_75 (.BL(BL75),.BLN(BLN75),.WL(WL22));
sram_cell_6t_5 inst_cell_22_76 (.BL(BL76),.BLN(BLN76),.WL(WL22));
sram_cell_6t_5 inst_cell_22_77 (.BL(BL77),.BLN(BLN77),.WL(WL22));
sram_cell_6t_5 inst_cell_22_78 (.BL(BL78),.BLN(BLN78),.WL(WL22));
sram_cell_6t_5 inst_cell_22_79 (.BL(BL79),.BLN(BLN79),.WL(WL22));
sram_cell_6t_5 inst_cell_22_80 (.BL(BL80),.BLN(BLN80),.WL(WL22));
sram_cell_6t_5 inst_cell_22_81 (.BL(BL81),.BLN(BLN81),.WL(WL22));
sram_cell_6t_5 inst_cell_22_82 (.BL(BL82),.BLN(BLN82),.WL(WL22));
sram_cell_6t_5 inst_cell_22_83 (.BL(BL83),.BLN(BLN83),.WL(WL22));
sram_cell_6t_5 inst_cell_22_84 (.BL(BL84),.BLN(BLN84),.WL(WL22));
sram_cell_6t_5 inst_cell_22_85 (.BL(BL85),.BLN(BLN85),.WL(WL22));
sram_cell_6t_5 inst_cell_22_86 (.BL(BL86),.BLN(BLN86),.WL(WL22));
sram_cell_6t_5 inst_cell_22_87 (.BL(BL87),.BLN(BLN87),.WL(WL22));
sram_cell_6t_5 inst_cell_22_88 (.BL(BL88),.BLN(BLN88),.WL(WL22));
sram_cell_6t_5 inst_cell_22_89 (.BL(BL89),.BLN(BLN89),.WL(WL22));
sram_cell_6t_5 inst_cell_22_90 (.BL(BL90),.BLN(BLN90),.WL(WL22));
sram_cell_6t_5 inst_cell_22_91 (.BL(BL91),.BLN(BLN91),.WL(WL22));
sram_cell_6t_5 inst_cell_22_92 (.BL(BL92),.BLN(BLN92),.WL(WL22));
sram_cell_6t_5 inst_cell_22_93 (.BL(BL93),.BLN(BLN93),.WL(WL22));
sram_cell_6t_5 inst_cell_22_94 (.BL(BL94),.BLN(BLN94),.WL(WL22));
sram_cell_6t_5 inst_cell_22_95 (.BL(BL95),.BLN(BLN95),.WL(WL22));
sram_cell_6t_5 inst_cell_22_96 (.BL(BL96),.BLN(BLN96),.WL(WL22));
sram_cell_6t_5 inst_cell_22_97 (.BL(BL97),.BLN(BLN97),.WL(WL22));
sram_cell_6t_5 inst_cell_22_98 (.BL(BL98),.BLN(BLN98),.WL(WL22));
sram_cell_6t_5 inst_cell_22_99 (.BL(BL99),.BLN(BLN99),.WL(WL22));
sram_cell_6t_5 inst_cell_22_100 (.BL(BL100),.BLN(BLN100),.WL(WL22));
sram_cell_6t_5 inst_cell_22_101 (.BL(BL101),.BLN(BLN101),.WL(WL22));
sram_cell_6t_5 inst_cell_22_102 (.BL(BL102),.BLN(BLN102),.WL(WL22));
sram_cell_6t_5 inst_cell_22_103 (.BL(BL103),.BLN(BLN103),.WL(WL22));
sram_cell_6t_5 inst_cell_22_104 (.BL(BL104),.BLN(BLN104),.WL(WL22));
sram_cell_6t_5 inst_cell_22_105 (.BL(BL105),.BLN(BLN105),.WL(WL22));
sram_cell_6t_5 inst_cell_22_106 (.BL(BL106),.BLN(BLN106),.WL(WL22));
sram_cell_6t_5 inst_cell_22_107 (.BL(BL107),.BLN(BLN107),.WL(WL22));
sram_cell_6t_5 inst_cell_22_108 (.BL(BL108),.BLN(BLN108),.WL(WL22));
sram_cell_6t_5 inst_cell_22_109 (.BL(BL109),.BLN(BLN109),.WL(WL22));
sram_cell_6t_5 inst_cell_22_110 (.BL(BL110),.BLN(BLN110),.WL(WL22));
sram_cell_6t_5 inst_cell_22_111 (.BL(BL111),.BLN(BLN111),.WL(WL22));
sram_cell_6t_5 inst_cell_22_112 (.BL(BL112),.BLN(BLN112),.WL(WL22));
sram_cell_6t_5 inst_cell_22_113 (.BL(BL113),.BLN(BLN113),.WL(WL22));
sram_cell_6t_5 inst_cell_22_114 (.BL(BL114),.BLN(BLN114),.WL(WL22));
sram_cell_6t_5 inst_cell_22_115 (.BL(BL115),.BLN(BLN115),.WL(WL22));
sram_cell_6t_5 inst_cell_22_116 (.BL(BL116),.BLN(BLN116),.WL(WL22));
sram_cell_6t_5 inst_cell_22_117 (.BL(BL117),.BLN(BLN117),.WL(WL22));
sram_cell_6t_5 inst_cell_22_118 (.BL(BL118),.BLN(BLN118),.WL(WL22));
sram_cell_6t_5 inst_cell_22_119 (.BL(BL119),.BLN(BLN119),.WL(WL22));
sram_cell_6t_5 inst_cell_22_120 (.BL(BL120),.BLN(BLN120),.WL(WL22));
sram_cell_6t_5 inst_cell_22_121 (.BL(BL121),.BLN(BLN121),.WL(WL22));
sram_cell_6t_5 inst_cell_22_122 (.BL(BL122),.BLN(BLN122),.WL(WL22));
sram_cell_6t_5 inst_cell_22_123 (.BL(BL123),.BLN(BLN123),.WL(WL22));
sram_cell_6t_5 inst_cell_22_124 (.BL(BL124),.BLN(BLN124),.WL(WL22));
sram_cell_6t_5 inst_cell_22_125 (.BL(BL125),.BLN(BLN125),.WL(WL22));
sram_cell_6t_5 inst_cell_22_126 (.BL(BL126),.BLN(BLN126),.WL(WL22));
sram_cell_6t_5 inst_cell_22_127 (.BL(BL127),.BLN(BLN127),.WL(WL22));
sram_cell_6t_5 inst_cell_23_0 (.BL(BL0),.BLN(BLN0),.WL(WL23));
sram_cell_6t_5 inst_cell_23_1 (.BL(BL1),.BLN(BLN1),.WL(WL23));
sram_cell_6t_5 inst_cell_23_2 (.BL(BL2),.BLN(BLN2),.WL(WL23));
sram_cell_6t_5 inst_cell_23_3 (.BL(BL3),.BLN(BLN3),.WL(WL23));
sram_cell_6t_5 inst_cell_23_4 (.BL(BL4),.BLN(BLN4),.WL(WL23));
sram_cell_6t_5 inst_cell_23_5 (.BL(BL5),.BLN(BLN5),.WL(WL23));
sram_cell_6t_5 inst_cell_23_6 (.BL(BL6),.BLN(BLN6),.WL(WL23));
sram_cell_6t_5 inst_cell_23_7 (.BL(BL7),.BLN(BLN7),.WL(WL23));
sram_cell_6t_5 inst_cell_23_8 (.BL(BL8),.BLN(BLN8),.WL(WL23));
sram_cell_6t_5 inst_cell_23_9 (.BL(BL9),.BLN(BLN9),.WL(WL23));
sram_cell_6t_5 inst_cell_23_10 (.BL(BL10),.BLN(BLN10),.WL(WL23));
sram_cell_6t_5 inst_cell_23_11 (.BL(BL11),.BLN(BLN11),.WL(WL23));
sram_cell_6t_5 inst_cell_23_12 (.BL(BL12),.BLN(BLN12),.WL(WL23));
sram_cell_6t_5 inst_cell_23_13 (.BL(BL13),.BLN(BLN13),.WL(WL23));
sram_cell_6t_5 inst_cell_23_14 (.BL(BL14),.BLN(BLN14),.WL(WL23));
sram_cell_6t_5 inst_cell_23_15 (.BL(BL15),.BLN(BLN15),.WL(WL23));
sram_cell_6t_5 inst_cell_23_16 (.BL(BL16),.BLN(BLN16),.WL(WL23));
sram_cell_6t_5 inst_cell_23_17 (.BL(BL17),.BLN(BLN17),.WL(WL23));
sram_cell_6t_5 inst_cell_23_18 (.BL(BL18),.BLN(BLN18),.WL(WL23));
sram_cell_6t_5 inst_cell_23_19 (.BL(BL19),.BLN(BLN19),.WL(WL23));
sram_cell_6t_5 inst_cell_23_20 (.BL(BL20),.BLN(BLN20),.WL(WL23));
sram_cell_6t_5 inst_cell_23_21 (.BL(BL21),.BLN(BLN21),.WL(WL23));
sram_cell_6t_5 inst_cell_23_22 (.BL(BL22),.BLN(BLN22),.WL(WL23));
sram_cell_6t_5 inst_cell_23_23 (.BL(BL23),.BLN(BLN23),.WL(WL23));
sram_cell_6t_5 inst_cell_23_24 (.BL(BL24),.BLN(BLN24),.WL(WL23));
sram_cell_6t_5 inst_cell_23_25 (.BL(BL25),.BLN(BLN25),.WL(WL23));
sram_cell_6t_5 inst_cell_23_26 (.BL(BL26),.BLN(BLN26),.WL(WL23));
sram_cell_6t_5 inst_cell_23_27 (.BL(BL27),.BLN(BLN27),.WL(WL23));
sram_cell_6t_5 inst_cell_23_28 (.BL(BL28),.BLN(BLN28),.WL(WL23));
sram_cell_6t_5 inst_cell_23_29 (.BL(BL29),.BLN(BLN29),.WL(WL23));
sram_cell_6t_5 inst_cell_23_30 (.BL(BL30),.BLN(BLN30),.WL(WL23));
sram_cell_6t_5 inst_cell_23_31 (.BL(BL31),.BLN(BLN31),.WL(WL23));
sram_cell_6t_5 inst_cell_23_32 (.BL(BL32),.BLN(BLN32),.WL(WL23));
sram_cell_6t_5 inst_cell_23_33 (.BL(BL33),.BLN(BLN33),.WL(WL23));
sram_cell_6t_5 inst_cell_23_34 (.BL(BL34),.BLN(BLN34),.WL(WL23));
sram_cell_6t_5 inst_cell_23_35 (.BL(BL35),.BLN(BLN35),.WL(WL23));
sram_cell_6t_5 inst_cell_23_36 (.BL(BL36),.BLN(BLN36),.WL(WL23));
sram_cell_6t_5 inst_cell_23_37 (.BL(BL37),.BLN(BLN37),.WL(WL23));
sram_cell_6t_5 inst_cell_23_38 (.BL(BL38),.BLN(BLN38),.WL(WL23));
sram_cell_6t_5 inst_cell_23_39 (.BL(BL39),.BLN(BLN39),.WL(WL23));
sram_cell_6t_5 inst_cell_23_40 (.BL(BL40),.BLN(BLN40),.WL(WL23));
sram_cell_6t_5 inst_cell_23_41 (.BL(BL41),.BLN(BLN41),.WL(WL23));
sram_cell_6t_5 inst_cell_23_42 (.BL(BL42),.BLN(BLN42),.WL(WL23));
sram_cell_6t_5 inst_cell_23_43 (.BL(BL43),.BLN(BLN43),.WL(WL23));
sram_cell_6t_5 inst_cell_23_44 (.BL(BL44),.BLN(BLN44),.WL(WL23));
sram_cell_6t_5 inst_cell_23_45 (.BL(BL45),.BLN(BLN45),.WL(WL23));
sram_cell_6t_5 inst_cell_23_46 (.BL(BL46),.BLN(BLN46),.WL(WL23));
sram_cell_6t_5 inst_cell_23_47 (.BL(BL47),.BLN(BLN47),.WL(WL23));
sram_cell_6t_5 inst_cell_23_48 (.BL(BL48),.BLN(BLN48),.WL(WL23));
sram_cell_6t_5 inst_cell_23_49 (.BL(BL49),.BLN(BLN49),.WL(WL23));
sram_cell_6t_5 inst_cell_23_50 (.BL(BL50),.BLN(BLN50),.WL(WL23));
sram_cell_6t_5 inst_cell_23_51 (.BL(BL51),.BLN(BLN51),.WL(WL23));
sram_cell_6t_5 inst_cell_23_52 (.BL(BL52),.BLN(BLN52),.WL(WL23));
sram_cell_6t_5 inst_cell_23_53 (.BL(BL53),.BLN(BLN53),.WL(WL23));
sram_cell_6t_5 inst_cell_23_54 (.BL(BL54),.BLN(BLN54),.WL(WL23));
sram_cell_6t_5 inst_cell_23_55 (.BL(BL55),.BLN(BLN55),.WL(WL23));
sram_cell_6t_5 inst_cell_23_56 (.BL(BL56),.BLN(BLN56),.WL(WL23));
sram_cell_6t_5 inst_cell_23_57 (.BL(BL57),.BLN(BLN57),.WL(WL23));
sram_cell_6t_5 inst_cell_23_58 (.BL(BL58),.BLN(BLN58),.WL(WL23));
sram_cell_6t_5 inst_cell_23_59 (.BL(BL59),.BLN(BLN59),.WL(WL23));
sram_cell_6t_5 inst_cell_23_60 (.BL(BL60),.BLN(BLN60),.WL(WL23));
sram_cell_6t_5 inst_cell_23_61 (.BL(BL61),.BLN(BLN61),.WL(WL23));
sram_cell_6t_5 inst_cell_23_62 (.BL(BL62),.BLN(BLN62),.WL(WL23));
sram_cell_6t_5 inst_cell_23_63 (.BL(BL63),.BLN(BLN63),.WL(WL23));
sram_cell_6t_5 inst_cell_23_64 (.BL(BL64),.BLN(BLN64),.WL(WL23));
sram_cell_6t_5 inst_cell_23_65 (.BL(BL65),.BLN(BLN65),.WL(WL23));
sram_cell_6t_5 inst_cell_23_66 (.BL(BL66),.BLN(BLN66),.WL(WL23));
sram_cell_6t_5 inst_cell_23_67 (.BL(BL67),.BLN(BLN67),.WL(WL23));
sram_cell_6t_5 inst_cell_23_68 (.BL(BL68),.BLN(BLN68),.WL(WL23));
sram_cell_6t_5 inst_cell_23_69 (.BL(BL69),.BLN(BLN69),.WL(WL23));
sram_cell_6t_5 inst_cell_23_70 (.BL(BL70),.BLN(BLN70),.WL(WL23));
sram_cell_6t_5 inst_cell_23_71 (.BL(BL71),.BLN(BLN71),.WL(WL23));
sram_cell_6t_5 inst_cell_23_72 (.BL(BL72),.BLN(BLN72),.WL(WL23));
sram_cell_6t_5 inst_cell_23_73 (.BL(BL73),.BLN(BLN73),.WL(WL23));
sram_cell_6t_5 inst_cell_23_74 (.BL(BL74),.BLN(BLN74),.WL(WL23));
sram_cell_6t_5 inst_cell_23_75 (.BL(BL75),.BLN(BLN75),.WL(WL23));
sram_cell_6t_5 inst_cell_23_76 (.BL(BL76),.BLN(BLN76),.WL(WL23));
sram_cell_6t_5 inst_cell_23_77 (.BL(BL77),.BLN(BLN77),.WL(WL23));
sram_cell_6t_5 inst_cell_23_78 (.BL(BL78),.BLN(BLN78),.WL(WL23));
sram_cell_6t_5 inst_cell_23_79 (.BL(BL79),.BLN(BLN79),.WL(WL23));
sram_cell_6t_5 inst_cell_23_80 (.BL(BL80),.BLN(BLN80),.WL(WL23));
sram_cell_6t_5 inst_cell_23_81 (.BL(BL81),.BLN(BLN81),.WL(WL23));
sram_cell_6t_5 inst_cell_23_82 (.BL(BL82),.BLN(BLN82),.WL(WL23));
sram_cell_6t_5 inst_cell_23_83 (.BL(BL83),.BLN(BLN83),.WL(WL23));
sram_cell_6t_5 inst_cell_23_84 (.BL(BL84),.BLN(BLN84),.WL(WL23));
sram_cell_6t_5 inst_cell_23_85 (.BL(BL85),.BLN(BLN85),.WL(WL23));
sram_cell_6t_5 inst_cell_23_86 (.BL(BL86),.BLN(BLN86),.WL(WL23));
sram_cell_6t_5 inst_cell_23_87 (.BL(BL87),.BLN(BLN87),.WL(WL23));
sram_cell_6t_5 inst_cell_23_88 (.BL(BL88),.BLN(BLN88),.WL(WL23));
sram_cell_6t_5 inst_cell_23_89 (.BL(BL89),.BLN(BLN89),.WL(WL23));
sram_cell_6t_5 inst_cell_23_90 (.BL(BL90),.BLN(BLN90),.WL(WL23));
sram_cell_6t_5 inst_cell_23_91 (.BL(BL91),.BLN(BLN91),.WL(WL23));
sram_cell_6t_5 inst_cell_23_92 (.BL(BL92),.BLN(BLN92),.WL(WL23));
sram_cell_6t_5 inst_cell_23_93 (.BL(BL93),.BLN(BLN93),.WL(WL23));
sram_cell_6t_5 inst_cell_23_94 (.BL(BL94),.BLN(BLN94),.WL(WL23));
sram_cell_6t_5 inst_cell_23_95 (.BL(BL95),.BLN(BLN95),.WL(WL23));
sram_cell_6t_5 inst_cell_23_96 (.BL(BL96),.BLN(BLN96),.WL(WL23));
sram_cell_6t_5 inst_cell_23_97 (.BL(BL97),.BLN(BLN97),.WL(WL23));
sram_cell_6t_5 inst_cell_23_98 (.BL(BL98),.BLN(BLN98),.WL(WL23));
sram_cell_6t_5 inst_cell_23_99 (.BL(BL99),.BLN(BLN99),.WL(WL23));
sram_cell_6t_5 inst_cell_23_100 (.BL(BL100),.BLN(BLN100),.WL(WL23));
sram_cell_6t_5 inst_cell_23_101 (.BL(BL101),.BLN(BLN101),.WL(WL23));
sram_cell_6t_5 inst_cell_23_102 (.BL(BL102),.BLN(BLN102),.WL(WL23));
sram_cell_6t_5 inst_cell_23_103 (.BL(BL103),.BLN(BLN103),.WL(WL23));
sram_cell_6t_5 inst_cell_23_104 (.BL(BL104),.BLN(BLN104),.WL(WL23));
sram_cell_6t_5 inst_cell_23_105 (.BL(BL105),.BLN(BLN105),.WL(WL23));
sram_cell_6t_5 inst_cell_23_106 (.BL(BL106),.BLN(BLN106),.WL(WL23));
sram_cell_6t_5 inst_cell_23_107 (.BL(BL107),.BLN(BLN107),.WL(WL23));
sram_cell_6t_5 inst_cell_23_108 (.BL(BL108),.BLN(BLN108),.WL(WL23));
sram_cell_6t_5 inst_cell_23_109 (.BL(BL109),.BLN(BLN109),.WL(WL23));
sram_cell_6t_5 inst_cell_23_110 (.BL(BL110),.BLN(BLN110),.WL(WL23));
sram_cell_6t_5 inst_cell_23_111 (.BL(BL111),.BLN(BLN111),.WL(WL23));
sram_cell_6t_5 inst_cell_23_112 (.BL(BL112),.BLN(BLN112),.WL(WL23));
sram_cell_6t_5 inst_cell_23_113 (.BL(BL113),.BLN(BLN113),.WL(WL23));
sram_cell_6t_5 inst_cell_23_114 (.BL(BL114),.BLN(BLN114),.WL(WL23));
sram_cell_6t_5 inst_cell_23_115 (.BL(BL115),.BLN(BLN115),.WL(WL23));
sram_cell_6t_5 inst_cell_23_116 (.BL(BL116),.BLN(BLN116),.WL(WL23));
sram_cell_6t_5 inst_cell_23_117 (.BL(BL117),.BLN(BLN117),.WL(WL23));
sram_cell_6t_5 inst_cell_23_118 (.BL(BL118),.BLN(BLN118),.WL(WL23));
sram_cell_6t_5 inst_cell_23_119 (.BL(BL119),.BLN(BLN119),.WL(WL23));
sram_cell_6t_5 inst_cell_23_120 (.BL(BL120),.BLN(BLN120),.WL(WL23));
sram_cell_6t_5 inst_cell_23_121 (.BL(BL121),.BLN(BLN121),.WL(WL23));
sram_cell_6t_5 inst_cell_23_122 (.BL(BL122),.BLN(BLN122),.WL(WL23));
sram_cell_6t_5 inst_cell_23_123 (.BL(BL123),.BLN(BLN123),.WL(WL23));
sram_cell_6t_5 inst_cell_23_124 (.BL(BL124),.BLN(BLN124),.WL(WL23));
sram_cell_6t_5 inst_cell_23_125 (.BL(BL125),.BLN(BLN125),.WL(WL23));
sram_cell_6t_5 inst_cell_23_126 (.BL(BL126),.BLN(BLN126),.WL(WL23));
sram_cell_6t_5 inst_cell_23_127 (.BL(BL127),.BLN(BLN127),.WL(WL23));
sram_cell_6t_5 inst_cell_24_0 (.BL(BL0),.BLN(BLN0),.WL(WL24));
sram_cell_6t_5 inst_cell_24_1 (.BL(BL1),.BLN(BLN1),.WL(WL24));
sram_cell_6t_5 inst_cell_24_2 (.BL(BL2),.BLN(BLN2),.WL(WL24));
sram_cell_6t_5 inst_cell_24_3 (.BL(BL3),.BLN(BLN3),.WL(WL24));
sram_cell_6t_5 inst_cell_24_4 (.BL(BL4),.BLN(BLN4),.WL(WL24));
sram_cell_6t_5 inst_cell_24_5 (.BL(BL5),.BLN(BLN5),.WL(WL24));
sram_cell_6t_5 inst_cell_24_6 (.BL(BL6),.BLN(BLN6),.WL(WL24));
sram_cell_6t_5 inst_cell_24_7 (.BL(BL7),.BLN(BLN7),.WL(WL24));
sram_cell_6t_5 inst_cell_24_8 (.BL(BL8),.BLN(BLN8),.WL(WL24));
sram_cell_6t_5 inst_cell_24_9 (.BL(BL9),.BLN(BLN9),.WL(WL24));
sram_cell_6t_5 inst_cell_24_10 (.BL(BL10),.BLN(BLN10),.WL(WL24));
sram_cell_6t_5 inst_cell_24_11 (.BL(BL11),.BLN(BLN11),.WL(WL24));
sram_cell_6t_5 inst_cell_24_12 (.BL(BL12),.BLN(BLN12),.WL(WL24));
sram_cell_6t_5 inst_cell_24_13 (.BL(BL13),.BLN(BLN13),.WL(WL24));
sram_cell_6t_5 inst_cell_24_14 (.BL(BL14),.BLN(BLN14),.WL(WL24));
sram_cell_6t_5 inst_cell_24_15 (.BL(BL15),.BLN(BLN15),.WL(WL24));
sram_cell_6t_5 inst_cell_24_16 (.BL(BL16),.BLN(BLN16),.WL(WL24));
sram_cell_6t_5 inst_cell_24_17 (.BL(BL17),.BLN(BLN17),.WL(WL24));
sram_cell_6t_5 inst_cell_24_18 (.BL(BL18),.BLN(BLN18),.WL(WL24));
sram_cell_6t_5 inst_cell_24_19 (.BL(BL19),.BLN(BLN19),.WL(WL24));
sram_cell_6t_5 inst_cell_24_20 (.BL(BL20),.BLN(BLN20),.WL(WL24));
sram_cell_6t_5 inst_cell_24_21 (.BL(BL21),.BLN(BLN21),.WL(WL24));
sram_cell_6t_5 inst_cell_24_22 (.BL(BL22),.BLN(BLN22),.WL(WL24));
sram_cell_6t_5 inst_cell_24_23 (.BL(BL23),.BLN(BLN23),.WL(WL24));
sram_cell_6t_5 inst_cell_24_24 (.BL(BL24),.BLN(BLN24),.WL(WL24));
sram_cell_6t_5 inst_cell_24_25 (.BL(BL25),.BLN(BLN25),.WL(WL24));
sram_cell_6t_5 inst_cell_24_26 (.BL(BL26),.BLN(BLN26),.WL(WL24));
sram_cell_6t_5 inst_cell_24_27 (.BL(BL27),.BLN(BLN27),.WL(WL24));
sram_cell_6t_5 inst_cell_24_28 (.BL(BL28),.BLN(BLN28),.WL(WL24));
sram_cell_6t_5 inst_cell_24_29 (.BL(BL29),.BLN(BLN29),.WL(WL24));
sram_cell_6t_5 inst_cell_24_30 (.BL(BL30),.BLN(BLN30),.WL(WL24));
sram_cell_6t_5 inst_cell_24_31 (.BL(BL31),.BLN(BLN31),.WL(WL24));
sram_cell_6t_5 inst_cell_24_32 (.BL(BL32),.BLN(BLN32),.WL(WL24));
sram_cell_6t_5 inst_cell_24_33 (.BL(BL33),.BLN(BLN33),.WL(WL24));
sram_cell_6t_5 inst_cell_24_34 (.BL(BL34),.BLN(BLN34),.WL(WL24));
sram_cell_6t_5 inst_cell_24_35 (.BL(BL35),.BLN(BLN35),.WL(WL24));
sram_cell_6t_5 inst_cell_24_36 (.BL(BL36),.BLN(BLN36),.WL(WL24));
sram_cell_6t_5 inst_cell_24_37 (.BL(BL37),.BLN(BLN37),.WL(WL24));
sram_cell_6t_5 inst_cell_24_38 (.BL(BL38),.BLN(BLN38),.WL(WL24));
sram_cell_6t_5 inst_cell_24_39 (.BL(BL39),.BLN(BLN39),.WL(WL24));
sram_cell_6t_5 inst_cell_24_40 (.BL(BL40),.BLN(BLN40),.WL(WL24));
sram_cell_6t_5 inst_cell_24_41 (.BL(BL41),.BLN(BLN41),.WL(WL24));
sram_cell_6t_5 inst_cell_24_42 (.BL(BL42),.BLN(BLN42),.WL(WL24));
sram_cell_6t_5 inst_cell_24_43 (.BL(BL43),.BLN(BLN43),.WL(WL24));
sram_cell_6t_5 inst_cell_24_44 (.BL(BL44),.BLN(BLN44),.WL(WL24));
sram_cell_6t_5 inst_cell_24_45 (.BL(BL45),.BLN(BLN45),.WL(WL24));
sram_cell_6t_5 inst_cell_24_46 (.BL(BL46),.BLN(BLN46),.WL(WL24));
sram_cell_6t_5 inst_cell_24_47 (.BL(BL47),.BLN(BLN47),.WL(WL24));
sram_cell_6t_5 inst_cell_24_48 (.BL(BL48),.BLN(BLN48),.WL(WL24));
sram_cell_6t_5 inst_cell_24_49 (.BL(BL49),.BLN(BLN49),.WL(WL24));
sram_cell_6t_5 inst_cell_24_50 (.BL(BL50),.BLN(BLN50),.WL(WL24));
sram_cell_6t_5 inst_cell_24_51 (.BL(BL51),.BLN(BLN51),.WL(WL24));
sram_cell_6t_5 inst_cell_24_52 (.BL(BL52),.BLN(BLN52),.WL(WL24));
sram_cell_6t_5 inst_cell_24_53 (.BL(BL53),.BLN(BLN53),.WL(WL24));
sram_cell_6t_5 inst_cell_24_54 (.BL(BL54),.BLN(BLN54),.WL(WL24));
sram_cell_6t_5 inst_cell_24_55 (.BL(BL55),.BLN(BLN55),.WL(WL24));
sram_cell_6t_5 inst_cell_24_56 (.BL(BL56),.BLN(BLN56),.WL(WL24));
sram_cell_6t_5 inst_cell_24_57 (.BL(BL57),.BLN(BLN57),.WL(WL24));
sram_cell_6t_5 inst_cell_24_58 (.BL(BL58),.BLN(BLN58),.WL(WL24));
sram_cell_6t_5 inst_cell_24_59 (.BL(BL59),.BLN(BLN59),.WL(WL24));
sram_cell_6t_5 inst_cell_24_60 (.BL(BL60),.BLN(BLN60),.WL(WL24));
sram_cell_6t_5 inst_cell_24_61 (.BL(BL61),.BLN(BLN61),.WL(WL24));
sram_cell_6t_5 inst_cell_24_62 (.BL(BL62),.BLN(BLN62),.WL(WL24));
sram_cell_6t_5 inst_cell_24_63 (.BL(BL63),.BLN(BLN63),.WL(WL24));
sram_cell_6t_5 inst_cell_24_64 (.BL(BL64),.BLN(BLN64),.WL(WL24));
sram_cell_6t_5 inst_cell_24_65 (.BL(BL65),.BLN(BLN65),.WL(WL24));
sram_cell_6t_5 inst_cell_24_66 (.BL(BL66),.BLN(BLN66),.WL(WL24));
sram_cell_6t_5 inst_cell_24_67 (.BL(BL67),.BLN(BLN67),.WL(WL24));
sram_cell_6t_5 inst_cell_24_68 (.BL(BL68),.BLN(BLN68),.WL(WL24));
sram_cell_6t_5 inst_cell_24_69 (.BL(BL69),.BLN(BLN69),.WL(WL24));
sram_cell_6t_5 inst_cell_24_70 (.BL(BL70),.BLN(BLN70),.WL(WL24));
sram_cell_6t_5 inst_cell_24_71 (.BL(BL71),.BLN(BLN71),.WL(WL24));
sram_cell_6t_5 inst_cell_24_72 (.BL(BL72),.BLN(BLN72),.WL(WL24));
sram_cell_6t_5 inst_cell_24_73 (.BL(BL73),.BLN(BLN73),.WL(WL24));
sram_cell_6t_5 inst_cell_24_74 (.BL(BL74),.BLN(BLN74),.WL(WL24));
sram_cell_6t_5 inst_cell_24_75 (.BL(BL75),.BLN(BLN75),.WL(WL24));
sram_cell_6t_5 inst_cell_24_76 (.BL(BL76),.BLN(BLN76),.WL(WL24));
sram_cell_6t_5 inst_cell_24_77 (.BL(BL77),.BLN(BLN77),.WL(WL24));
sram_cell_6t_5 inst_cell_24_78 (.BL(BL78),.BLN(BLN78),.WL(WL24));
sram_cell_6t_5 inst_cell_24_79 (.BL(BL79),.BLN(BLN79),.WL(WL24));
sram_cell_6t_5 inst_cell_24_80 (.BL(BL80),.BLN(BLN80),.WL(WL24));
sram_cell_6t_5 inst_cell_24_81 (.BL(BL81),.BLN(BLN81),.WL(WL24));
sram_cell_6t_5 inst_cell_24_82 (.BL(BL82),.BLN(BLN82),.WL(WL24));
sram_cell_6t_5 inst_cell_24_83 (.BL(BL83),.BLN(BLN83),.WL(WL24));
sram_cell_6t_5 inst_cell_24_84 (.BL(BL84),.BLN(BLN84),.WL(WL24));
sram_cell_6t_5 inst_cell_24_85 (.BL(BL85),.BLN(BLN85),.WL(WL24));
sram_cell_6t_5 inst_cell_24_86 (.BL(BL86),.BLN(BLN86),.WL(WL24));
sram_cell_6t_5 inst_cell_24_87 (.BL(BL87),.BLN(BLN87),.WL(WL24));
sram_cell_6t_5 inst_cell_24_88 (.BL(BL88),.BLN(BLN88),.WL(WL24));
sram_cell_6t_5 inst_cell_24_89 (.BL(BL89),.BLN(BLN89),.WL(WL24));
sram_cell_6t_5 inst_cell_24_90 (.BL(BL90),.BLN(BLN90),.WL(WL24));
sram_cell_6t_5 inst_cell_24_91 (.BL(BL91),.BLN(BLN91),.WL(WL24));
sram_cell_6t_5 inst_cell_24_92 (.BL(BL92),.BLN(BLN92),.WL(WL24));
sram_cell_6t_5 inst_cell_24_93 (.BL(BL93),.BLN(BLN93),.WL(WL24));
sram_cell_6t_5 inst_cell_24_94 (.BL(BL94),.BLN(BLN94),.WL(WL24));
sram_cell_6t_5 inst_cell_24_95 (.BL(BL95),.BLN(BLN95),.WL(WL24));
sram_cell_6t_5 inst_cell_24_96 (.BL(BL96),.BLN(BLN96),.WL(WL24));
sram_cell_6t_5 inst_cell_24_97 (.BL(BL97),.BLN(BLN97),.WL(WL24));
sram_cell_6t_5 inst_cell_24_98 (.BL(BL98),.BLN(BLN98),.WL(WL24));
sram_cell_6t_5 inst_cell_24_99 (.BL(BL99),.BLN(BLN99),.WL(WL24));
sram_cell_6t_5 inst_cell_24_100 (.BL(BL100),.BLN(BLN100),.WL(WL24));
sram_cell_6t_5 inst_cell_24_101 (.BL(BL101),.BLN(BLN101),.WL(WL24));
sram_cell_6t_5 inst_cell_24_102 (.BL(BL102),.BLN(BLN102),.WL(WL24));
sram_cell_6t_5 inst_cell_24_103 (.BL(BL103),.BLN(BLN103),.WL(WL24));
sram_cell_6t_5 inst_cell_24_104 (.BL(BL104),.BLN(BLN104),.WL(WL24));
sram_cell_6t_5 inst_cell_24_105 (.BL(BL105),.BLN(BLN105),.WL(WL24));
sram_cell_6t_5 inst_cell_24_106 (.BL(BL106),.BLN(BLN106),.WL(WL24));
sram_cell_6t_5 inst_cell_24_107 (.BL(BL107),.BLN(BLN107),.WL(WL24));
sram_cell_6t_5 inst_cell_24_108 (.BL(BL108),.BLN(BLN108),.WL(WL24));
sram_cell_6t_5 inst_cell_24_109 (.BL(BL109),.BLN(BLN109),.WL(WL24));
sram_cell_6t_5 inst_cell_24_110 (.BL(BL110),.BLN(BLN110),.WL(WL24));
sram_cell_6t_5 inst_cell_24_111 (.BL(BL111),.BLN(BLN111),.WL(WL24));
sram_cell_6t_5 inst_cell_24_112 (.BL(BL112),.BLN(BLN112),.WL(WL24));
sram_cell_6t_5 inst_cell_24_113 (.BL(BL113),.BLN(BLN113),.WL(WL24));
sram_cell_6t_5 inst_cell_24_114 (.BL(BL114),.BLN(BLN114),.WL(WL24));
sram_cell_6t_5 inst_cell_24_115 (.BL(BL115),.BLN(BLN115),.WL(WL24));
sram_cell_6t_5 inst_cell_24_116 (.BL(BL116),.BLN(BLN116),.WL(WL24));
sram_cell_6t_5 inst_cell_24_117 (.BL(BL117),.BLN(BLN117),.WL(WL24));
sram_cell_6t_5 inst_cell_24_118 (.BL(BL118),.BLN(BLN118),.WL(WL24));
sram_cell_6t_5 inst_cell_24_119 (.BL(BL119),.BLN(BLN119),.WL(WL24));
sram_cell_6t_5 inst_cell_24_120 (.BL(BL120),.BLN(BLN120),.WL(WL24));
sram_cell_6t_5 inst_cell_24_121 (.BL(BL121),.BLN(BLN121),.WL(WL24));
sram_cell_6t_5 inst_cell_24_122 (.BL(BL122),.BLN(BLN122),.WL(WL24));
sram_cell_6t_5 inst_cell_24_123 (.BL(BL123),.BLN(BLN123),.WL(WL24));
sram_cell_6t_5 inst_cell_24_124 (.BL(BL124),.BLN(BLN124),.WL(WL24));
sram_cell_6t_5 inst_cell_24_125 (.BL(BL125),.BLN(BLN125),.WL(WL24));
sram_cell_6t_5 inst_cell_24_126 (.BL(BL126),.BLN(BLN126),.WL(WL24));
sram_cell_6t_5 inst_cell_24_127 (.BL(BL127),.BLN(BLN127),.WL(WL24));
sram_cell_6t_5 inst_cell_25_0 (.BL(BL0),.BLN(BLN0),.WL(WL25));
sram_cell_6t_5 inst_cell_25_1 (.BL(BL1),.BLN(BLN1),.WL(WL25));
sram_cell_6t_5 inst_cell_25_2 (.BL(BL2),.BLN(BLN2),.WL(WL25));
sram_cell_6t_5 inst_cell_25_3 (.BL(BL3),.BLN(BLN3),.WL(WL25));
sram_cell_6t_5 inst_cell_25_4 (.BL(BL4),.BLN(BLN4),.WL(WL25));
sram_cell_6t_5 inst_cell_25_5 (.BL(BL5),.BLN(BLN5),.WL(WL25));
sram_cell_6t_5 inst_cell_25_6 (.BL(BL6),.BLN(BLN6),.WL(WL25));
sram_cell_6t_5 inst_cell_25_7 (.BL(BL7),.BLN(BLN7),.WL(WL25));
sram_cell_6t_5 inst_cell_25_8 (.BL(BL8),.BLN(BLN8),.WL(WL25));
sram_cell_6t_5 inst_cell_25_9 (.BL(BL9),.BLN(BLN9),.WL(WL25));
sram_cell_6t_5 inst_cell_25_10 (.BL(BL10),.BLN(BLN10),.WL(WL25));
sram_cell_6t_5 inst_cell_25_11 (.BL(BL11),.BLN(BLN11),.WL(WL25));
sram_cell_6t_5 inst_cell_25_12 (.BL(BL12),.BLN(BLN12),.WL(WL25));
sram_cell_6t_5 inst_cell_25_13 (.BL(BL13),.BLN(BLN13),.WL(WL25));
sram_cell_6t_5 inst_cell_25_14 (.BL(BL14),.BLN(BLN14),.WL(WL25));
sram_cell_6t_5 inst_cell_25_15 (.BL(BL15),.BLN(BLN15),.WL(WL25));
sram_cell_6t_5 inst_cell_25_16 (.BL(BL16),.BLN(BLN16),.WL(WL25));
sram_cell_6t_5 inst_cell_25_17 (.BL(BL17),.BLN(BLN17),.WL(WL25));
sram_cell_6t_5 inst_cell_25_18 (.BL(BL18),.BLN(BLN18),.WL(WL25));
sram_cell_6t_5 inst_cell_25_19 (.BL(BL19),.BLN(BLN19),.WL(WL25));
sram_cell_6t_5 inst_cell_25_20 (.BL(BL20),.BLN(BLN20),.WL(WL25));
sram_cell_6t_5 inst_cell_25_21 (.BL(BL21),.BLN(BLN21),.WL(WL25));
sram_cell_6t_5 inst_cell_25_22 (.BL(BL22),.BLN(BLN22),.WL(WL25));
sram_cell_6t_5 inst_cell_25_23 (.BL(BL23),.BLN(BLN23),.WL(WL25));
sram_cell_6t_5 inst_cell_25_24 (.BL(BL24),.BLN(BLN24),.WL(WL25));
sram_cell_6t_5 inst_cell_25_25 (.BL(BL25),.BLN(BLN25),.WL(WL25));
sram_cell_6t_5 inst_cell_25_26 (.BL(BL26),.BLN(BLN26),.WL(WL25));
sram_cell_6t_5 inst_cell_25_27 (.BL(BL27),.BLN(BLN27),.WL(WL25));
sram_cell_6t_5 inst_cell_25_28 (.BL(BL28),.BLN(BLN28),.WL(WL25));
sram_cell_6t_5 inst_cell_25_29 (.BL(BL29),.BLN(BLN29),.WL(WL25));
sram_cell_6t_5 inst_cell_25_30 (.BL(BL30),.BLN(BLN30),.WL(WL25));
sram_cell_6t_5 inst_cell_25_31 (.BL(BL31),.BLN(BLN31),.WL(WL25));
sram_cell_6t_5 inst_cell_25_32 (.BL(BL32),.BLN(BLN32),.WL(WL25));
sram_cell_6t_5 inst_cell_25_33 (.BL(BL33),.BLN(BLN33),.WL(WL25));
sram_cell_6t_5 inst_cell_25_34 (.BL(BL34),.BLN(BLN34),.WL(WL25));
sram_cell_6t_5 inst_cell_25_35 (.BL(BL35),.BLN(BLN35),.WL(WL25));
sram_cell_6t_5 inst_cell_25_36 (.BL(BL36),.BLN(BLN36),.WL(WL25));
sram_cell_6t_5 inst_cell_25_37 (.BL(BL37),.BLN(BLN37),.WL(WL25));
sram_cell_6t_5 inst_cell_25_38 (.BL(BL38),.BLN(BLN38),.WL(WL25));
sram_cell_6t_5 inst_cell_25_39 (.BL(BL39),.BLN(BLN39),.WL(WL25));
sram_cell_6t_5 inst_cell_25_40 (.BL(BL40),.BLN(BLN40),.WL(WL25));
sram_cell_6t_5 inst_cell_25_41 (.BL(BL41),.BLN(BLN41),.WL(WL25));
sram_cell_6t_5 inst_cell_25_42 (.BL(BL42),.BLN(BLN42),.WL(WL25));
sram_cell_6t_5 inst_cell_25_43 (.BL(BL43),.BLN(BLN43),.WL(WL25));
sram_cell_6t_5 inst_cell_25_44 (.BL(BL44),.BLN(BLN44),.WL(WL25));
sram_cell_6t_5 inst_cell_25_45 (.BL(BL45),.BLN(BLN45),.WL(WL25));
sram_cell_6t_5 inst_cell_25_46 (.BL(BL46),.BLN(BLN46),.WL(WL25));
sram_cell_6t_5 inst_cell_25_47 (.BL(BL47),.BLN(BLN47),.WL(WL25));
sram_cell_6t_5 inst_cell_25_48 (.BL(BL48),.BLN(BLN48),.WL(WL25));
sram_cell_6t_5 inst_cell_25_49 (.BL(BL49),.BLN(BLN49),.WL(WL25));
sram_cell_6t_5 inst_cell_25_50 (.BL(BL50),.BLN(BLN50),.WL(WL25));
sram_cell_6t_5 inst_cell_25_51 (.BL(BL51),.BLN(BLN51),.WL(WL25));
sram_cell_6t_5 inst_cell_25_52 (.BL(BL52),.BLN(BLN52),.WL(WL25));
sram_cell_6t_5 inst_cell_25_53 (.BL(BL53),.BLN(BLN53),.WL(WL25));
sram_cell_6t_5 inst_cell_25_54 (.BL(BL54),.BLN(BLN54),.WL(WL25));
sram_cell_6t_5 inst_cell_25_55 (.BL(BL55),.BLN(BLN55),.WL(WL25));
sram_cell_6t_5 inst_cell_25_56 (.BL(BL56),.BLN(BLN56),.WL(WL25));
sram_cell_6t_5 inst_cell_25_57 (.BL(BL57),.BLN(BLN57),.WL(WL25));
sram_cell_6t_5 inst_cell_25_58 (.BL(BL58),.BLN(BLN58),.WL(WL25));
sram_cell_6t_5 inst_cell_25_59 (.BL(BL59),.BLN(BLN59),.WL(WL25));
sram_cell_6t_5 inst_cell_25_60 (.BL(BL60),.BLN(BLN60),.WL(WL25));
sram_cell_6t_5 inst_cell_25_61 (.BL(BL61),.BLN(BLN61),.WL(WL25));
sram_cell_6t_5 inst_cell_25_62 (.BL(BL62),.BLN(BLN62),.WL(WL25));
sram_cell_6t_5 inst_cell_25_63 (.BL(BL63),.BLN(BLN63),.WL(WL25));
sram_cell_6t_5 inst_cell_25_64 (.BL(BL64),.BLN(BLN64),.WL(WL25));
sram_cell_6t_5 inst_cell_25_65 (.BL(BL65),.BLN(BLN65),.WL(WL25));
sram_cell_6t_5 inst_cell_25_66 (.BL(BL66),.BLN(BLN66),.WL(WL25));
sram_cell_6t_5 inst_cell_25_67 (.BL(BL67),.BLN(BLN67),.WL(WL25));
sram_cell_6t_5 inst_cell_25_68 (.BL(BL68),.BLN(BLN68),.WL(WL25));
sram_cell_6t_5 inst_cell_25_69 (.BL(BL69),.BLN(BLN69),.WL(WL25));
sram_cell_6t_5 inst_cell_25_70 (.BL(BL70),.BLN(BLN70),.WL(WL25));
sram_cell_6t_5 inst_cell_25_71 (.BL(BL71),.BLN(BLN71),.WL(WL25));
sram_cell_6t_5 inst_cell_25_72 (.BL(BL72),.BLN(BLN72),.WL(WL25));
sram_cell_6t_5 inst_cell_25_73 (.BL(BL73),.BLN(BLN73),.WL(WL25));
sram_cell_6t_5 inst_cell_25_74 (.BL(BL74),.BLN(BLN74),.WL(WL25));
sram_cell_6t_5 inst_cell_25_75 (.BL(BL75),.BLN(BLN75),.WL(WL25));
sram_cell_6t_5 inst_cell_25_76 (.BL(BL76),.BLN(BLN76),.WL(WL25));
sram_cell_6t_5 inst_cell_25_77 (.BL(BL77),.BLN(BLN77),.WL(WL25));
sram_cell_6t_5 inst_cell_25_78 (.BL(BL78),.BLN(BLN78),.WL(WL25));
sram_cell_6t_5 inst_cell_25_79 (.BL(BL79),.BLN(BLN79),.WL(WL25));
sram_cell_6t_5 inst_cell_25_80 (.BL(BL80),.BLN(BLN80),.WL(WL25));
sram_cell_6t_5 inst_cell_25_81 (.BL(BL81),.BLN(BLN81),.WL(WL25));
sram_cell_6t_5 inst_cell_25_82 (.BL(BL82),.BLN(BLN82),.WL(WL25));
sram_cell_6t_5 inst_cell_25_83 (.BL(BL83),.BLN(BLN83),.WL(WL25));
sram_cell_6t_5 inst_cell_25_84 (.BL(BL84),.BLN(BLN84),.WL(WL25));
sram_cell_6t_5 inst_cell_25_85 (.BL(BL85),.BLN(BLN85),.WL(WL25));
sram_cell_6t_5 inst_cell_25_86 (.BL(BL86),.BLN(BLN86),.WL(WL25));
sram_cell_6t_5 inst_cell_25_87 (.BL(BL87),.BLN(BLN87),.WL(WL25));
sram_cell_6t_5 inst_cell_25_88 (.BL(BL88),.BLN(BLN88),.WL(WL25));
sram_cell_6t_5 inst_cell_25_89 (.BL(BL89),.BLN(BLN89),.WL(WL25));
sram_cell_6t_5 inst_cell_25_90 (.BL(BL90),.BLN(BLN90),.WL(WL25));
sram_cell_6t_5 inst_cell_25_91 (.BL(BL91),.BLN(BLN91),.WL(WL25));
sram_cell_6t_5 inst_cell_25_92 (.BL(BL92),.BLN(BLN92),.WL(WL25));
sram_cell_6t_5 inst_cell_25_93 (.BL(BL93),.BLN(BLN93),.WL(WL25));
sram_cell_6t_5 inst_cell_25_94 (.BL(BL94),.BLN(BLN94),.WL(WL25));
sram_cell_6t_5 inst_cell_25_95 (.BL(BL95),.BLN(BLN95),.WL(WL25));
sram_cell_6t_5 inst_cell_25_96 (.BL(BL96),.BLN(BLN96),.WL(WL25));
sram_cell_6t_5 inst_cell_25_97 (.BL(BL97),.BLN(BLN97),.WL(WL25));
sram_cell_6t_5 inst_cell_25_98 (.BL(BL98),.BLN(BLN98),.WL(WL25));
sram_cell_6t_5 inst_cell_25_99 (.BL(BL99),.BLN(BLN99),.WL(WL25));
sram_cell_6t_5 inst_cell_25_100 (.BL(BL100),.BLN(BLN100),.WL(WL25));
sram_cell_6t_5 inst_cell_25_101 (.BL(BL101),.BLN(BLN101),.WL(WL25));
sram_cell_6t_5 inst_cell_25_102 (.BL(BL102),.BLN(BLN102),.WL(WL25));
sram_cell_6t_5 inst_cell_25_103 (.BL(BL103),.BLN(BLN103),.WL(WL25));
sram_cell_6t_5 inst_cell_25_104 (.BL(BL104),.BLN(BLN104),.WL(WL25));
sram_cell_6t_5 inst_cell_25_105 (.BL(BL105),.BLN(BLN105),.WL(WL25));
sram_cell_6t_5 inst_cell_25_106 (.BL(BL106),.BLN(BLN106),.WL(WL25));
sram_cell_6t_5 inst_cell_25_107 (.BL(BL107),.BLN(BLN107),.WL(WL25));
sram_cell_6t_5 inst_cell_25_108 (.BL(BL108),.BLN(BLN108),.WL(WL25));
sram_cell_6t_5 inst_cell_25_109 (.BL(BL109),.BLN(BLN109),.WL(WL25));
sram_cell_6t_5 inst_cell_25_110 (.BL(BL110),.BLN(BLN110),.WL(WL25));
sram_cell_6t_5 inst_cell_25_111 (.BL(BL111),.BLN(BLN111),.WL(WL25));
sram_cell_6t_5 inst_cell_25_112 (.BL(BL112),.BLN(BLN112),.WL(WL25));
sram_cell_6t_5 inst_cell_25_113 (.BL(BL113),.BLN(BLN113),.WL(WL25));
sram_cell_6t_5 inst_cell_25_114 (.BL(BL114),.BLN(BLN114),.WL(WL25));
sram_cell_6t_5 inst_cell_25_115 (.BL(BL115),.BLN(BLN115),.WL(WL25));
sram_cell_6t_5 inst_cell_25_116 (.BL(BL116),.BLN(BLN116),.WL(WL25));
sram_cell_6t_5 inst_cell_25_117 (.BL(BL117),.BLN(BLN117),.WL(WL25));
sram_cell_6t_5 inst_cell_25_118 (.BL(BL118),.BLN(BLN118),.WL(WL25));
sram_cell_6t_5 inst_cell_25_119 (.BL(BL119),.BLN(BLN119),.WL(WL25));
sram_cell_6t_5 inst_cell_25_120 (.BL(BL120),.BLN(BLN120),.WL(WL25));
sram_cell_6t_5 inst_cell_25_121 (.BL(BL121),.BLN(BLN121),.WL(WL25));
sram_cell_6t_5 inst_cell_25_122 (.BL(BL122),.BLN(BLN122),.WL(WL25));
sram_cell_6t_5 inst_cell_25_123 (.BL(BL123),.BLN(BLN123),.WL(WL25));
sram_cell_6t_5 inst_cell_25_124 (.BL(BL124),.BLN(BLN124),.WL(WL25));
sram_cell_6t_5 inst_cell_25_125 (.BL(BL125),.BLN(BLN125),.WL(WL25));
sram_cell_6t_5 inst_cell_25_126 (.BL(BL126),.BLN(BLN126),.WL(WL25));
sram_cell_6t_5 inst_cell_25_127 (.BL(BL127),.BLN(BLN127),.WL(WL25));
sram_cell_6t_5 inst_cell_26_0 (.BL(BL0),.BLN(BLN0),.WL(WL26));
sram_cell_6t_5 inst_cell_26_1 (.BL(BL1),.BLN(BLN1),.WL(WL26));
sram_cell_6t_5 inst_cell_26_2 (.BL(BL2),.BLN(BLN2),.WL(WL26));
sram_cell_6t_5 inst_cell_26_3 (.BL(BL3),.BLN(BLN3),.WL(WL26));
sram_cell_6t_5 inst_cell_26_4 (.BL(BL4),.BLN(BLN4),.WL(WL26));
sram_cell_6t_5 inst_cell_26_5 (.BL(BL5),.BLN(BLN5),.WL(WL26));
sram_cell_6t_5 inst_cell_26_6 (.BL(BL6),.BLN(BLN6),.WL(WL26));
sram_cell_6t_5 inst_cell_26_7 (.BL(BL7),.BLN(BLN7),.WL(WL26));
sram_cell_6t_5 inst_cell_26_8 (.BL(BL8),.BLN(BLN8),.WL(WL26));
sram_cell_6t_5 inst_cell_26_9 (.BL(BL9),.BLN(BLN9),.WL(WL26));
sram_cell_6t_5 inst_cell_26_10 (.BL(BL10),.BLN(BLN10),.WL(WL26));
sram_cell_6t_5 inst_cell_26_11 (.BL(BL11),.BLN(BLN11),.WL(WL26));
sram_cell_6t_5 inst_cell_26_12 (.BL(BL12),.BLN(BLN12),.WL(WL26));
sram_cell_6t_5 inst_cell_26_13 (.BL(BL13),.BLN(BLN13),.WL(WL26));
sram_cell_6t_5 inst_cell_26_14 (.BL(BL14),.BLN(BLN14),.WL(WL26));
sram_cell_6t_5 inst_cell_26_15 (.BL(BL15),.BLN(BLN15),.WL(WL26));
sram_cell_6t_5 inst_cell_26_16 (.BL(BL16),.BLN(BLN16),.WL(WL26));
sram_cell_6t_5 inst_cell_26_17 (.BL(BL17),.BLN(BLN17),.WL(WL26));
sram_cell_6t_5 inst_cell_26_18 (.BL(BL18),.BLN(BLN18),.WL(WL26));
sram_cell_6t_5 inst_cell_26_19 (.BL(BL19),.BLN(BLN19),.WL(WL26));
sram_cell_6t_5 inst_cell_26_20 (.BL(BL20),.BLN(BLN20),.WL(WL26));
sram_cell_6t_5 inst_cell_26_21 (.BL(BL21),.BLN(BLN21),.WL(WL26));
sram_cell_6t_5 inst_cell_26_22 (.BL(BL22),.BLN(BLN22),.WL(WL26));
sram_cell_6t_5 inst_cell_26_23 (.BL(BL23),.BLN(BLN23),.WL(WL26));
sram_cell_6t_5 inst_cell_26_24 (.BL(BL24),.BLN(BLN24),.WL(WL26));
sram_cell_6t_5 inst_cell_26_25 (.BL(BL25),.BLN(BLN25),.WL(WL26));
sram_cell_6t_5 inst_cell_26_26 (.BL(BL26),.BLN(BLN26),.WL(WL26));
sram_cell_6t_5 inst_cell_26_27 (.BL(BL27),.BLN(BLN27),.WL(WL26));
sram_cell_6t_5 inst_cell_26_28 (.BL(BL28),.BLN(BLN28),.WL(WL26));
sram_cell_6t_5 inst_cell_26_29 (.BL(BL29),.BLN(BLN29),.WL(WL26));
sram_cell_6t_5 inst_cell_26_30 (.BL(BL30),.BLN(BLN30),.WL(WL26));
sram_cell_6t_5 inst_cell_26_31 (.BL(BL31),.BLN(BLN31),.WL(WL26));
sram_cell_6t_5 inst_cell_26_32 (.BL(BL32),.BLN(BLN32),.WL(WL26));
sram_cell_6t_5 inst_cell_26_33 (.BL(BL33),.BLN(BLN33),.WL(WL26));
sram_cell_6t_5 inst_cell_26_34 (.BL(BL34),.BLN(BLN34),.WL(WL26));
sram_cell_6t_5 inst_cell_26_35 (.BL(BL35),.BLN(BLN35),.WL(WL26));
sram_cell_6t_5 inst_cell_26_36 (.BL(BL36),.BLN(BLN36),.WL(WL26));
sram_cell_6t_5 inst_cell_26_37 (.BL(BL37),.BLN(BLN37),.WL(WL26));
sram_cell_6t_5 inst_cell_26_38 (.BL(BL38),.BLN(BLN38),.WL(WL26));
sram_cell_6t_5 inst_cell_26_39 (.BL(BL39),.BLN(BLN39),.WL(WL26));
sram_cell_6t_5 inst_cell_26_40 (.BL(BL40),.BLN(BLN40),.WL(WL26));
sram_cell_6t_5 inst_cell_26_41 (.BL(BL41),.BLN(BLN41),.WL(WL26));
sram_cell_6t_5 inst_cell_26_42 (.BL(BL42),.BLN(BLN42),.WL(WL26));
sram_cell_6t_5 inst_cell_26_43 (.BL(BL43),.BLN(BLN43),.WL(WL26));
sram_cell_6t_5 inst_cell_26_44 (.BL(BL44),.BLN(BLN44),.WL(WL26));
sram_cell_6t_5 inst_cell_26_45 (.BL(BL45),.BLN(BLN45),.WL(WL26));
sram_cell_6t_5 inst_cell_26_46 (.BL(BL46),.BLN(BLN46),.WL(WL26));
sram_cell_6t_5 inst_cell_26_47 (.BL(BL47),.BLN(BLN47),.WL(WL26));
sram_cell_6t_5 inst_cell_26_48 (.BL(BL48),.BLN(BLN48),.WL(WL26));
sram_cell_6t_5 inst_cell_26_49 (.BL(BL49),.BLN(BLN49),.WL(WL26));
sram_cell_6t_5 inst_cell_26_50 (.BL(BL50),.BLN(BLN50),.WL(WL26));
sram_cell_6t_5 inst_cell_26_51 (.BL(BL51),.BLN(BLN51),.WL(WL26));
sram_cell_6t_5 inst_cell_26_52 (.BL(BL52),.BLN(BLN52),.WL(WL26));
sram_cell_6t_5 inst_cell_26_53 (.BL(BL53),.BLN(BLN53),.WL(WL26));
sram_cell_6t_5 inst_cell_26_54 (.BL(BL54),.BLN(BLN54),.WL(WL26));
sram_cell_6t_5 inst_cell_26_55 (.BL(BL55),.BLN(BLN55),.WL(WL26));
sram_cell_6t_5 inst_cell_26_56 (.BL(BL56),.BLN(BLN56),.WL(WL26));
sram_cell_6t_5 inst_cell_26_57 (.BL(BL57),.BLN(BLN57),.WL(WL26));
sram_cell_6t_5 inst_cell_26_58 (.BL(BL58),.BLN(BLN58),.WL(WL26));
sram_cell_6t_5 inst_cell_26_59 (.BL(BL59),.BLN(BLN59),.WL(WL26));
sram_cell_6t_5 inst_cell_26_60 (.BL(BL60),.BLN(BLN60),.WL(WL26));
sram_cell_6t_5 inst_cell_26_61 (.BL(BL61),.BLN(BLN61),.WL(WL26));
sram_cell_6t_5 inst_cell_26_62 (.BL(BL62),.BLN(BLN62),.WL(WL26));
sram_cell_6t_5 inst_cell_26_63 (.BL(BL63),.BLN(BLN63),.WL(WL26));
sram_cell_6t_5 inst_cell_26_64 (.BL(BL64),.BLN(BLN64),.WL(WL26));
sram_cell_6t_5 inst_cell_26_65 (.BL(BL65),.BLN(BLN65),.WL(WL26));
sram_cell_6t_5 inst_cell_26_66 (.BL(BL66),.BLN(BLN66),.WL(WL26));
sram_cell_6t_5 inst_cell_26_67 (.BL(BL67),.BLN(BLN67),.WL(WL26));
sram_cell_6t_5 inst_cell_26_68 (.BL(BL68),.BLN(BLN68),.WL(WL26));
sram_cell_6t_5 inst_cell_26_69 (.BL(BL69),.BLN(BLN69),.WL(WL26));
sram_cell_6t_5 inst_cell_26_70 (.BL(BL70),.BLN(BLN70),.WL(WL26));
sram_cell_6t_5 inst_cell_26_71 (.BL(BL71),.BLN(BLN71),.WL(WL26));
sram_cell_6t_5 inst_cell_26_72 (.BL(BL72),.BLN(BLN72),.WL(WL26));
sram_cell_6t_5 inst_cell_26_73 (.BL(BL73),.BLN(BLN73),.WL(WL26));
sram_cell_6t_5 inst_cell_26_74 (.BL(BL74),.BLN(BLN74),.WL(WL26));
sram_cell_6t_5 inst_cell_26_75 (.BL(BL75),.BLN(BLN75),.WL(WL26));
sram_cell_6t_5 inst_cell_26_76 (.BL(BL76),.BLN(BLN76),.WL(WL26));
sram_cell_6t_5 inst_cell_26_77 (.BL(BL77),.BLN(BLN77),.WL(WL26));
sram_cell_6t_5 inst_cell_26_78 (.BL(BL78),.BLN(BLN78),.WL(WL26));
sram_cell_6t_5 inst_cell_26_79 (.BL(BL79),.BLN(BLN79),.WL(WL26));
sram_cell_6t_5 inst_cell_26_80 (.BL(BL80),.BLN(BLN80),.WL(WL26));
sram_cell_6t_5 inst_cell_26_81 (.BL(BL81),.BLN(BLN81),.WL(WL26));
sram_cell_6t_5 inst_cell_26_82 (.BL(BL82),.BLN(BLN82),.WL(WL26));
sram_cell_6t_5 inst_cell_26_83 (.BL(BL83),.BLN(BLN83),.WL(WL26));
sram_cell_6t_5 inst_cell_26_84 (.BL(BL84),.BLN(BLN84),.WL(WL26));
sram_cell_6t_5 inst_cell_26_85 (.BL(BL85),.BLN(BLN85),.WL(WL26));
sram_cell_6t_5 inst_cell_26_86 (.BL(BL86),.BLN(BLN86),.WL(WL26));
sram_cell_6t_5 inst_cell_26_87 (.BL(BL87),.BLN(BLN87),.WL(WL26));
sram_cell_6t_5 inst_cell_26_88 (.BL(BL88),.BLN(BLN88),.WL(WL26));
sram_cell_6t_5 inst_cell_26_89 (.BL(BL89),.BLN(BLN89),.WL(WL26));
sram_cell_6t_5 inst_cell_26_90 (.BL(BL90),.BLN(BLN90),.WL(WL26));
sram_cell_6t_5 inst_cell_26_91 (.BL(BL91),.BLN(BLN91),.WL(WL26));
sram_cell_6t_5 inst_cell_26_92 (.BL(BL92),.BLN(BLN92),.WL(WL26));
sram_cell_6t_5 inst_cell_26_93 (.BL(BL93),.BLN(BLN93),.WL(WL26));
sram_cell_6t_5 inst_cell_26_94 (.BL(BL94),.BLN(BLN94),.WL(WL26));
sram_cell_6t_5 inst_cell_26_95 (.BL(BL95),.BLN(BLN95),.WL(WL26));
sram_cell_6t_5 inst_cell_26_96 (.BL(BL96),.BLN(BLN96),.WL(WL26));
sram_cell_6t_5 inst_cell_26_97 (.BL(BL97),.BLN(BLN97),.WL(WL26));
sram_cell_6t_5 inst_cell_26_98 (.BL(BL98),.BLN(BLN98),.WL(WL26));
sram_cell_6t_5 inst_cell_26_99 (.BL(BL99),.BLN(BLN99),.WL(WL26));
sram_cell_6t_5 inst_cell_26_100 (.BL(BL100),.BLN(BLN100),.WL(WL26));
sram_cell_6t_5 inst_cell_26_101 (.BL(BL101),.BLN(BLN101),.WL(WL26));
sram_cell_6t_5 inst_cell_26_102 (.BL(BL102),.BLN(BLN102),.WL(WL26));
sram_cell_6t_5 inst_cell_26_103 (.BL(BL103),.BLN(BLN103),.WL(WL26));
sram_cell_6t_5 inst_cell_26_104 (.BL(BL104),.BLN(BLN104),.WL(WL26));
sram_cell_6t_5 inst_cell_26_105 (.BL(BL105),.BLN(BLN105),.WL(WL26));
sram_cell_6t_5 inst_cell_26_106 (.BL(BL106),.BLN(BLN106),.WL(WL26));
sram_cell_6t_5 inst_cell_26_107 (.BL(BL107),.BLN(BLN107),.WL(WL26));
sram_cell_6t_5 inst_cell_26_108 (.BL(BL108),.BLN(BLN108),.WL(WL26));
sram_cell_6t_5 inst_cell_26_109 (.BL(BL109),.BLN(BLN109),.WL(WL26));
sram_cell_6t_5 inst_cell_26_110 (.BL(BL110),.BLN(BLN110),.WL(WL26));
sram_cell_6t_5 inst_cell_26_111 (.BL(BL111),.BLN(BLN111),.WL(WL26));
sram_cell_6t_5 inst_cell_26_112 (.BL(BL112),.BLN(BLN112),.WL(WL26));
sram_cell_6t_5 inst_cell_26_113 (.BL(BL113),.BLN(BLN113),.WL(WL26));
sram_cell_6t_5 inst_cell_26_114 (.BL(BL114),.BLN(BLN114),.WL(WL26));
sram_cell_6t_5 inst_cell_26_115 (.BL(BL115),.BLN(BLN115),.WL(WL26));
sram_cell_6t_5 inst_cell_26_116 (.BL(BL116),.BLN(BLN116),.WL(WL26));
sram_cell_6t_5 inst_cell_26_117 (.BL(BL117),.BLN(BLN117),.WL(WL26));
sram_cell_6t_5 inst_cell_26_118 (.BL(BL118),.BLN(BLN118),.WL(WL26));
sram_cell_6t_5 inst_cell_26_119 (.BL(BL119),.BLN(BLN119),.WL(WL26));
sram_cell_6t_5 inst_cell_26_120 (.BL(BL120),.BLN(BLN120),.WL(WL26));
sram_cell_6t_5 inst_cell_26_121 (.BL(BL121),.BLN(BLN121),.WL(WL26));
sram_cell_6t_5 inst_cell_26_122 (.BL(BL122),.BLN(BLN122),.WL(WL26));
sram_cell_6t_5 inst_cell_26_123 (.BL(BL123),.BLN(BLN123),.WL(WL26));
sram_cell_6t_5 inst_cell_26_124 (.BL(BL124),.BLN(BLN124),.WL(WL26));
sram_cell_6t_5 inst_cell_26_125 (.BL(BL125),.BLN(BLN125),.WL(WL26));
sram_cell_6t_5 inst_cell_26_126 (.BL(BL126),.BLN(BLN126),.WL(WL26));
sram_cell_6t_5 inst_cell_26_127 (.BL(BL127),.BLN(BLN127),.WL(WL26));
sram_cell_6t_5 inst_cell_27_0 (.BL(BL0),.BLN(BLN0),.WL(WL27));
sram_cell_6t_5 inst_cell_27_1 (.BL(BL1),.BLN(BLN1),.WL(WL27));
sram_cell_6t_5 inst_cell_27_2 (.BL(BL2),.BLN(BLN2),.WL(WL27));
sram_cell_6t_5 inst_cell_27_3 (.BL(BL3),.BLN(BLN3),.WL(WL27));
sram_cell_6t_5 inst_cell_27_4 (.BL(BL4),.BLN(BLN4),.WL(WL27));
sram_cell_6t_5 inst_cell_27_5 (.BL(BL5),.BLN(BLN5),.WL(WL27));
sram_cell_6t_5 inst_cell_27_6 (.BL(BL6),.BLN(BLN6),.WL(WL27));
sram_cell_6t_5 inst_cell_27_7 (.BL(BL7),.BLN(BLN7),.WL(WL27));
sram_cell_6t_5 inst_cell_27_8 (.BL(BL8),.BLN(BLN8),.WL(WL27));
sram_cell_6t_5 inst_cell_27_9 (.BL(BL9),.BLN(BLN9),.WL(WL27));
sram_cell_6t_5 inst_cell_27_10 (.BL(BL10),.BLN(BLN10),.WL(WL27));
sram_cell_6t_5 inst_cell_27_11 (.BL(BL11),.BLN(BLN11),.WL(WL27));
sram_cell_6t_5 inst_cell_27_12 (.BL(BL12),.BLN(BLN12),.WL(WL27));
sram_cell_6t_5 inst_cell_27_13 (.BL(BL13),.BLN(BLN13),.WL(WL27));
sram_cell_6t_5 inst_cell_27_14 (.BL(BL14),.BLN(BLN14),.WL(WL27));
sram_cell_6t_5 inst_cell_27_15 (.BL(BL15),.BLN(BLN15),.WL(WL27));
sram_cell_6t_5 inst_cell_27_16 (.BL(BL16),.BLN(BLN16),.WL(WL27));
sram_cell_6t_5 inst_cell_27_17 (.BL(BL17),.BLN(BLN17),.WL(WL27));
sram_cell_6t_5 inst_cell_27_18 (.BL(BL18),.BLN(BLN18),.WL(WL27));
sram_cell_6t_5 inst_cell_27_19 (.BL(BL19),.BLN(BLN19),.WL(WL27));
sram_cell_6t_5 inst_cell_27_20 (.BL(BL20),.BLN(BLN20),.WL(WL27));
sram_cell_6t_5 inst_cell_27_21 (.BL(BL21),.BLN(BLN21),.WL(WL27));
sram_cell_6t_5 inst_cell_27_22 (.BL(BL22),.BLN(BLN22),.WL(WL27));
sram_cell_6t_5 inst_cell_27_23 (.BL(BL23),.BLN(BLN23),.WL(WL27));
sram_cell_6t_5 inst_cell_27_24 (.BL(BL24),.BLN(BLN24),.WL(WL27));
sram_cell_6t_5 inst_cell_27_25 (.BL(BL25),.BLN(BLN25),.WL(WL27));
sram_cell_6t_5 inst_cell_27_26 (.BL(BL26),.BLN(BLN26),.WL(WL27));
sram_cell_6t_5 inst_cell_27_27 (.BL(BL27),.BLN(BLN27),.WL(WL27));
sram_cell_6t_5 inst_cell_27_28 (.BL(BL28),.BLN(BLN28),.WL(WL27));
sram_cell_6t_5 inst_cell_27_29 (.BL(BL29),.BLN(BLN29),.WL(WL27));
sram_cell_6t_5 inst_cell_27_30 (.BL(BL30),.BLN(BLN30),.WL(WL27));
sram_cell_6t_5 inst_cell_27_31 (.BL(BL31),.BLN(BLN31),.WL(WL27));
sram_cell_6t_5 inst_cell_27_32 (.BL(BL32),.BLN(BLN32),.WL(WL27));
sram_cell_6t_5 inst_cell_27_33 (.BL(BL33),.BLN(BLN33),.WL(WL27));
sram_cell_6t_5 inst_cell_27_34 (.BL(BL34),.BLN(BLN34),.WL(WL27));
sram_cell_6t_5 inst_cell_27_35 (.BL(BL35),.BLN(BLN35),.WL(WL27));
sram_cell_6t_5 inst_cell_27_36 (.BL(BL36),.BLN(BLN36),.WL(WL27));
sram_cell_6t_5 inst_cell_27_37 (.BL(BL37),.BLN(BLN37),.WL(WL27));
sram_cell_6t_5 inst_cell_27_38 (.BL(BL38),.BLN(BLN38),.WL(WL27));
sram_cell_6t_5 inst_cell_27_39 (.BL(BL39),.BLN(BLN39),.WL(WL27));
sram_cell_6t_5 inst_cell_27_40 (.BL(BL40),.BLN(BLN40),.WL(WL27));
sram_cell_6t_5 inst_cell_27_41 (.BL(BL41),.BLN(BLN41),.WL(WL27));
sram_cell_6t_5 inst_cell_27_42 (.BL(BL42),.BLN(BLN42),.WL(WL27));
sram_cell_6t_5 inst_cell_27_43 (.BL(BL43),.BLN(BLN43),.WL(WL27));
sram_cell_6t_5 inst_cell_27_44 (.BL(BL44),.BLN(BLN44),.WL(WL27));
sram_cell_6t_5 inst_cell_27_45 (.BL(BL45),.BLN(BLN45),.WL(WL27));
sram_cell_6t_5 inst_cell_27_46 (.BL(BL46),.BLN(BLN46),.WL(WL27));
sram_cell_6t_5 inst_cell_27_47 (.BL(BL47),.BLN(BLN47),.WL(WL27));
sram_cell_6t_5 inst_cell_27_48 (.BL(BL48),.BLN(BLN48),.WL(WL27));
sram_cell_6t_5 inst_cell_27_49 (.BL(BL49),.BLN(BLN49),.WL(WL27));
sram_cell_6t_5 inst_cell_27_50 (.BL(BL50),.BLN(BLN50),.WL(WL27));
sram_cell_6t_5 inst_cell_27_51 (.BL(BL51),.BLN(BLN51),.WL(WL27));
sram_cell_6t_5 inst_cell_27_52 (.BL(BL52),.BLN(BLN52),.WL(WL27));
sram_cell_6t_5 inst_cell_27_53 (.BL(BL53),.BLN(BLN53),.WL(WL27));
sram_cell_6t_5 inst_cell_27_54 (.BL(BL54),.BLN(BLN54),.WL(WL27));
sram_cell_6t_5 inst_cell_27_55 (.BL(BL55),.BLN(BLN55),.WL(WL27));
sram_cell_6t_5 inst_cell_27_56 (.BL(BL56),.BLN(BLN56),.WL(WL27));
sram_cell_6t_5 inst_cell_27_57 (.BL(BL57),.BLN(BLN57),.WL(WL27));
sram_cell_6t_5 inst_cell_27_58 (.BL(BL58),.BLN(BLN58),.WL(WL27));
sram_cell_6t_5 inst_cell_27_59 (.BL(BL59),.BLN(BLN59),.WL(WL27));
sram_cell_6t_5 inst_cell_27_60 (.BL(BL60),.BLN(BLN60),.WL(WL27));
sram_cell_6t_5 inst_cell_27_61 (.BL(BL61),.BLN(BLN61),.WL(WL27));
sram_cell_6t_5 inst_cell_27_62 (.BL(BL62),.BLN(BLN62),.WL(WL27));
sram_cell_6t_5 inst_cell_27_63 (.BL(BL63),.BLN(BLN63),.WL(WL27));
sram_cell_6t_5 inst_cell_27_64 (.BL(BL64),.BLN(BLN64),.WL(WL27));
sram_cell_6t_5 inst_cell_27_65 (.BL(BL65),.BLN(BLN65),.WL(WL27));
sram_cell_6t_5 inst_cell_27_66 (.BL(BL66),.BLN(BLN66),.WL(WL27));
sram_cell_6t_5 inst_cell_27_67 (.BL(BL67),.BLN(BLN67),.WL(WL27));
sram_cell_6t_5 inst_cell_27_68 (.BL(BL68),.BLN(BLN68),.WL(WL27));
sram_cell_6t_5 inst_cell_27_69 (.BL(BL69),.BLN(BLN69),.WL(WL27));
sram_cell_6t_5 inst_cell_27_70 (.BL(BL70),.BLN(BLN70),.WL(WL27));
sram_cell_6t_5 inst_cell_27_71 (.BL(BL71),.BLN(BLN71),.WL(WL27));
sram_cell_6t_5 inst_cell_27_72 (.BL(BL72),.BLN(BLN72),.WL(WL27));
sram_cell_6t_5 inst_cell_27_73 (.BL(BL73),.BLN(BLN73),.WL(WL27));
sram_cell_6t_5 inst_cell_27_74 (.BL(BL74),.BLN(BLN74),.WL(WL27));
sram_cell_6t_5 inst_cell_27_75 (.BL(BL75),.BLN(BLN75),.WL(WL27));
sram_cell_6t_5 inst_cell_27_76 (.BL(BL76),.BLN(BLN76),.WL(WL27));
sram_cell_6t_5 inst_cell_27_77 (.BL(BL77),.BLN(BLN77),.WL(WL27));
sram_cell_6t_5 inst_cell_27_78 (.BL(BL78),.BLN(BLN78),.WL(WL27));
sram_cell_6t_5 inst_cell_27_79 (.BL(BL79),.BLN(BLN79),.WL(WL27));
sram_cell_6t_5 inst_cell_27_80 (.BL(BL80),.BLN(BLN80),.WL(WL27));
sram_cell_6t_5 inst_cell_27_81 (.BL(BL81),.BLN(BLN81),.WL(WL27));
sram_cell_6t_5 inst_cell_27_82 (.BL(BL82),.BLN(BLN82),.WL(WL27));
sram_cell_6t_5 inst_cell_27_83 (.BL(BL83),.BLN(BLN83),.WL(WL27));
sram_cell_6t_5 inst_cell_27_84 (.BL(BL84),.BLN(BLN84),.WL(WL27));
sram_cell_6t_5 inst_cell_27_85 (.BL(BL85),.BLN(BLN85),.WL(WL27));
sram_cell_6t_5 inst_cell_27_86 (.BL(BL86),.BLN(BLN86),.WL(WL27));
sram_cell_6t_5 inst_cell_27_87 (.BL(BL87),.BLN(BLN87),.WL(WL27));
sram_cell_6t_5 inst_cell_27_88 (.BL(BL88),.BLN(BLN88),.WL(WL27));
sram_cell_6t_5 inst_cell_27_89 (.BL(BL89),.BLN(BLN89),.WL(WL27));
sram_cell_6t_5 inst_cell_27_90 (.BL(BL90),.BLN(BLN90),.WL(WL27));
sram_cell_6t_5 inst_cell_27_91 (.BL(BL91),.BLN(BLN91),.WL(WL27));
sram_cell_6t_5 inst_cell_27_92 (.BL(BL92),.BLN(BLN92),.WL(WL27));
sram_cell_6t_5 inst_cell_27_93 (.BL(BL93),.BLN(BLN93),.WL(WL27));
sram_cell_6t_5 inst_cell_27_94 (.BL(BL94),.BLN(BLN94),.WL(WL27));
sram_cell_6t_5 inst_cell_27_95 (.BL(BL95),.BLN(BLN95),.WL(WL27));
sram_cell_6t_5 inst_cell_27_96 (.BL(BL96),.BLN(BLN96),.WL(WL27));
sram_cell_6t_5 inst_cell_27_97 (.BL(BL97),.BLN(BLN97),.WL(WL27));
sram_cell_6t_5 inst_cell_27_98 (.BL(BL98),.BLN(BLN98),.WL(WL27));
sram_cell_6t_5 inst_cell_27_99 (.BL(BL99),.BLN(BLN99),.WL(WL27));
sram_cell_6t_5 inst_cell_27_100 (.BL(BL100),.BLN(BLN100),.WL(WL27));
sram_cell_6t_5 inst_cell_27_101 (.BL(BL101),.BLN(BLN101),.WL(WL27));
sram_cell_6t_5 inst_cell_27_102 (.BL(BL102),.BLN(BLN102),.WL(WL27));
sram_cell_6t_5 inst_cell_27_103 (.BL(BL103),.BLN(BLN103),.WL(WL27));
sram_cell_6t_5 inst_cell_27_104 (.BL(BL104),.BLN(BLN104),.WL(WL27));
sram_cell_6t_5 inst_cell_27_105 (.BL(BL105),.BLN(BLN105),.WL(WL27));
sram_cell_6t_5 inst_cell_27_106 (.BL(BL106),.BLN(BLN106),.WL(WL27));
sram_cell_6t_5 inst_cell_27_107 (.BL(BL107),.BLN(BLN107),.WL(WL27));
sram_cell_6t_5 inst_cell_27_108 (.BL(BL108),.BLN(BLN108),.WL(WL27));
sram_cell_6t_5 inst_cell_27_109 (.BL(BL109),.BLN(BLN109),.WL(WL27));
sram_cell_6t_5 inst_cell_27_110 (.BL(BL110),.BLN(BLN110),.WL(WL27));
sram_cell_6t_5 inst_cell_27_111 (.BL(BL111),.BLN(BLN111),.WL(WL27));
sram_cell_6t_5 inst_cell_27_112 (.BL(BL112),.BLN(BLN112),.WL(WL27));
sram_cell_6t_5 inst_cell_27_113 (.BL(BL113),.BLN(BLN113),.WL(WL27));
sram_cell_6t_5 inst_cell_27_114 (.BL(BL114),.BLN(BLN114),.WL(WL27));
sram_cell_6t_5 inst_cell_27_115 (.BL(BL115),.BLN(BLN115),.WL(WL27));
sram_cell_6t_5 inst_cell_27_116 (.BL(BL116),.BLN(BLN116),.WL(WL27));
sram_cell_6t_5 inst_cell_27_117 (.BL(BL117),.BLN(BLN117),.WL(WL27));
sram_cell_6t_5 inst_cell_27_118 (.BL(BL118),.BLN(BLN118),.WL(WL27));
sram_cell_6t_5 inst_cell_27_119 (.BL(BL119),.BLN(BLN119),.WL(WL27));
sram_cell_6t_5 inst_cell_27_120 (.BL(BL120),.BLN(BLN120),.WL(WL27));
sram_cell_6t_5 inst_cell_27_121 (.BL(BL121),.BLN(BLN121),.WL(WL27));
sram_cell_6t_5 inst_cell_27_122 (.BL(BL122),.BLN(BLN122),.WL(WL27));
sram_cell_6t_5 inst_cell_27_123 (.BL(BL123),.BLN(BLN123),.WL(WL27));
sram_cell_6t_5 inst_cell_27_124 (.BL(BL124),.BLN(BLN124),.WL(WL27));
sram_cell_6t_5 inst_cell_27_125 (.BL(BL125),.BLN(BLN125),.WL(WL27));
sram_cell_6t_5 inst_cell_27_126 (.BL(BL126),.BLN(BLN126),.WL(WL27));
sram_cell_6t_5 inst_cell_27_127 (.BL(BL127),.BLN(BLN127),.WL(WL27));
sram_cell_6t_5 inst_cell_28_0 (.BL(BL0),.BLN(BLN0),.WL(WL28));
sram_cell_6t_5 inst_cell_28_1 (.BL(BL1),.BLN(BLN1),.WL(WL28));
sram_cell_6t_5 inst_cell_28_2 (.BL(BL2),.BLN(BLN2),.WL(WL28));
sram_cell_6t_5 inst_cell_28_3 (.BL(BL3),.BLN(BLN3),.WL(WL28));
sram_cell_6t_5 inst_cell_28_4 (.BL(BL4),.BLN(BLN4),.WL(WL28));
sram_cell_6t_5 inst_cell_28_5 (.BL(BL5),.BLN(BLN5),.WL(WL28));
sram_cell_6t_5 inst_cell_28_6 (.BL(BL6),.BLN(BLN6),.WL(WL28));
sram_cell_6t_5 inst_cell_28_7 (.BL(BL7),.BLN(BLN7),.WL(WL28));
sram_cell_6t_5 inst_cell_28_8 (.BL(BL8),.BLN(BLN8),.WL(WL28));
sram_cell_6t_5 inst_cell_28_9 (.BL(BL9),.BLN(BLN9),.WL(WL28));
sram_cell_6t_5 inst_cell_28_10 (.BL(BL10),.BLN(BLN10),.WL(WL28));
sram_cell_6t_5 inst_cell_28_11 (.BL(BL11),.BLN(BLN11),.WL(WL28));
sram_cell_6t_5 inst_cell_28_12 (.BL(BL12),.BLN(BLN12),.WL(WL28));
sram_cell_6t_5 inst_cell_28_13 (.BL(BL13),.BLN(BLN13),.WL(WL28));
sram_cell_6t_5 inst_cell_28_14 (.BL(BL14),.BLN(BLN14),.WL(WL28));
sram_cell_6t_5 inst_cell_28_15 (.BL(BL15),.BLN(BLN15),.WL(WL28));
sram_cell_6t_5 inst_cell_28_16 (.BL(BL16),.BLN(BLN16),.WL(WL28));
sram_cell_6t_5 inst_cell_28_17 (.BL(BL17),.BLN(BLN17),.WL(WL28));
sram_cell_6t_5 inst_cell_28_18 (.BL(BL18),.BLN(BLN18),.WL(WL28));
sram_cell_6t_5 inst_cell_28_19 (.BL(BL19),.BLN(BLN19),.WL(WL28));
sram_cell_6t_5 inst_cell_28_20 (.BL(BL20),.BLN(BLN20),.WL(WL28));
sram_cell_6t_5 inst_cell_28_21 (.BL(BL21),.BLN(BLN21),.WL(WL28));
sram_cell_6t_5 inst_cell_28_22 (.BL(BL22),.BLN(BLN22),.WL(WL28));
sram_cell_6t_5 inst_cell_28_23 (.BL(BL23),.BLN(BLN23),.WL(WL28));
sram_cell_6t_5 inst_cell_28_24 (.BL(BL24),.BLN(BLN24),.WL(WL28));
sram_cell_6t_5 inst_cell_28_25 (.BL(BL25),.BLN(BLN25),.WL(WL28));
sram_cell_6t_5 inst_cell_28_26 (.BL(BL26),.BLN(BLN26),.WL(WL28));
sram_cell_6t_5 inst_cell_28_27 (.BL(BL27),.BLN(BLN27),.WL(WL28));
sram_cell_6t_5 inst_cell_28_28 (.BL(BL28),.BLN(BLN28),.WL(WL28));
sram_cell_6t_5 inst_cell_28_29 (.BL(BL29),.BLN(BLN29),.WL(WL28));
sram_cell_6t_5 inst_cell_28_30 (.BL(BL30),.BLN(BLN30),.WL(WL28));
sram_cell_6t_5 inst_cell_28_31 (.BL(BL31),.BLN(BLN31),.WL(WL28));
sram_cell_6t_5 inst_cell_28_32 (.BL(BL32),.BLN(BLN32),.WL(WL28));
sram_cell_6t_5 inst_cell_28_33 (.BL(BL33),.BLN(BLN33),.WL(WL28));
sram_cell_6t_5 inst_cell_28_34 (.BL(BL34),.BLN(BLN34),.WL(WL28));
sram_cell_6t_5 inst_cell_28_35 (.BL(BL35),.BLN(BLN35),.WL(WL28));
sram_cell_6t_5 inst_cell_28_36 (.BL(BL36),.BLN(BLN36),.WL(WL28));
sram_cell_6t_5 inst_cell_28_37 (.BL(BL37),.BLN(BLN37),.WL(WL28));
sram_cell_6t_5 inst_cell_28_38 (.BL(BL38),.BLN(BLN38),.WL(WL28));
sram_cell_6t_5 inst_cell_28_39 (.BL(BL39),.BLN(BLN39),.WL(WL28));
sram_cell_6t_5 inst_cell_28_40 (.BL(BL40),.BLN(BLN40),.WL(WL28));
sram_cell_6t_5 inst_cell_28_41 (.BL(BL41),.BLN(BLN41),.WL(WL28));
sram_cell_6t_5 inst_cell_28_42 (.BL(BL42),.BLN(BLN42),.WL(WL28));
sram_cell_6t_5 inst_cell_28_43 (.BL(BL43),.BLN(BLN43),.WL(WL28));
sram_cell_6t_5 inst_cell_28_44 (.BL(BL44),.BLN(BLN44),.WL(WL28));
sram_cell_6t_5 inst_cell_28_45 (.BL(BL45),.BLN(BLN45),.WL(WL28));
sram_cell_6t_5 inst_cell_28_46 (.BL(BL46),.BLN(BLN46),.WL(WL28));
sram_cell_6t_5 inst_cell_28_47 (.BL(BL47),.BLN(BLN47),.WL(WL28));
sram_cell_6t_5 inst_cell_28_48 (.BL(BL48),.BLN(BLN48),.WL(WL28));
sram_cell_6t_5 inst_cell_28_49 (.BL(BL49),.BLN(BLN49),.WL(WL28));
sram_cell_6t_5 inst_cell_28_50 (.BL(BL50),.BLN(BLN50),.WL(WL28));
sram_cell_6t_5 inst_cell_28_51 (.BL(BL51),.BLN(BLN51),.WL(WL28));
sram_cell_6t_5 inst_cell_28_52 (.BL(BL52),.BLN(BLN52),.WL(WL28));
sram_cell_6t_5 inst_cell_28_53 (.BL(BL53),.BLN(BLN53),.WL(WL28));
sram_cell_6t_5 inst_cell_28_54 (.BL(BL54),.BLN(BLN54),.WL(WL28));
sram_cell_6t_5 inst_cell_28_55 (.BL(BL55),.BLN(BLN55),.WL(WL28));
sram_cell_6t_5 inst_cell_28_56 (.BL(BL56),.BLN(BLN56),.WL(WL28));
sram_cell_6t_5 inst_cell_28_57 (.BL(BL57),.BLN(BLN57),.WL(WL28));
sram_cell_6t_5 inst_cell_28_58 (.BL(BL58),.BLN(BLN58),.WL(WL28));
sram_cell_6t_5 inst_cell_28_59 (.BL(BL59),.BLN(BLN59),.WL(WL28));
sram_cell_6t_5 inst_cell_28_60 (.BL(BL60),.BLN(BLN60),.WL(WL28));
sram_cell_6t_5 inst_cell_28_61 (.BL(BL61),.BLN(BLN61),.WL(WL28));
sram_cell_6t_5 inst_cell_28_62 (.BL(BL62),.BLN(BLN62),.WL(WL28));
sram_cell_6t_5 inst_cell_28_63 (.BL(BL63),.BLN(BLN63),.WL(WL28));
sram_cell_6t_5 inst_cell_28_64 (.BL(BL64),.BLN(BLN64),.WL(WL28));
sram_cell_6t_5 inst_cell_28_65 (.BL(BL65),.BLN(BLN65),.WL(WL28));
sram_cell_6t_5 inst_cell_28_66 (.BL(BL66),.BLN(BLN66),.WL(WL28));
sram_cell_6t_5 inst_cell_28_67 (.BL(BL67),.BLN(BLN67),.WL(WL28));
sram_cell_6t_5 inst_cell_28_68 (.BL(BL68),.BLN(BLN68),.WL(WL28));
sram_cell_6t_5 inst_cell_28_69 (.BL(BL69),.BLN(BLN69),.WL(WL28));
sram_cell_6t_5 inst_cell_28_70 (.BL(BL70),.BLN(BLN70),.WL(WL28));
sram_cell_6t_5 inst_cell_28_71 (.BL(BL71),.BLN(BLN71),.WL(WL28));
sram_cell_6t_5 inst_cell_28_72 (.BL(BL72),.BLN(BLN72),.WL(WL28));
sram_cell_6t_5 inst_cell_28_73 (.BL(BL73),.BLN(BLN73),.WL(WL28));
sram_cell_6t_5 inst_cell_28_74 (.BL(BL74),.BLN(BLN74),.WL(WL28));
sram_cell_6t_5 inst_cell_28_75 (.BL(BL75),.BLN(BLN75),.WL(WL28));
sram_cell_6t_5 inst_cell_28_76 (.BL(BL76),.BLN(BLN76),.WL(WL28));
sram_cell_6t_5 inst_cell_28_77 (.BL(BL77),.BLN(BLN77),.WL(WL28));
sram_cell_6t_5 inst_cell_28_78 (.BL(BL78),.BLN(BLN78),.WL(WL28));
sram_cell_6t_5 inst_cell_28_79 (.BL(BL79),.BLN(BLN79),.WL(WL28));
sram_cell_6t_5 inst_cell_28_80 (.BL(BL80),.BLN(BLN80),.WL(WL28));
sram_cell_6t_5 inst_cell_28_81 (.BL(BL81),.BLN(BLN81),.WL(WL28));
sram_cell_6t_5 inst_cell_28_82 (.BL(BL82),.BLN(BLN82),.WL(WL28));
sram_cell_6t_5 inst_cell_28_83 (.BL(BL83),.BLN(BLN83),.WL(WL28));
sram_cell_6t_5 inst_cell_28_84 (.BL(BL84),.BLN(BLN84),.WL(WL28));
sram_cell_6t_5 inst_cell_28_85 (.BL(BL85),.BLN(BLN85),.WL(WL28));
sram_cell_6t_5 inst_cell_28_86 (.BL(BL86),.BLN(BLN86),.WL(WL28));
sram_cell_6t_5 inst_cell_28_87 (.BL(BL87),.BLN(BLN87),.WL(WL28));
sram_cell_6t_5 inst_cell_28_88 (.BL(BL88),.BLN(BLN88),.WL(WL28));
sram_cell_6t_5 inst_cell_28_89 (.BL(BL89),.BLN(BLN89),.WL(WL28));
sram_cell_6t_5 inst_cell_28_90 (.BL(BL90),.BLN(BLN90),.WL(WL28));
sram_cell_6t_5 inst_cell_28_91 (.BL(BL91),.BLN(BLN91),.WL(WL28));
sram_cell_6t_5 inst_cell_28_92 (.BL(BL92),.BLN(BLN92),.WL(WL28));
sram_cell_6t_5 inst_cell_28_93 (.BL(BL93),.BLN(BLN93),.WL(WL28));
sram_cell_6t_5 inst_cell_28_94 (.BL(BL94),.BLN(BLN94),.WL(WL28));
sram_cell_6t_5 inst_cell_28_95 (.BL(BL95),.BLN(BLN95),.WL(WL28));
sram_cell_6t_5 inst_cell_28_96 (.BL(BL96),.BLN(BLN96),.WL(WL28));
sram_cell_6t_5 inst_cell_28_97 (.BL(BL97),.BLN(BLN97),.WL(WL28));
sram_cell_6t_5 inst_cell_28_98 (.BL(BL98),.BLN(BLN98),.WL(WL28));
sram_cell_6t_5 inst_cell_28_99 (.BL(BL99),.BLN(BLN99),.WL(WL28));
sram_cell_6t_5 inst_cell_28_100 (.BL(BL100),.BLN(BLN100),.WL(WL28));
sram_cell_6t_5 inst_cell_28_101 (.BL(BL101),.BLN(BLN101),.WL(WL28));
sram_cell_6t_5 inst_cell_28_102 (.BL(BL102),.BLN(BLN102),.WL(WL28));
sram_cell_6t_5 inst_cell_28_103 (.BL(BL103),.BLN(BLN103),.WL(WL28));
sram_cell_6t_5 inst_cell_28_104 (.BL(BL104),.BLN(BLN104),.WL(WL28));
sram_cell_6t_5 inst_cell_28_105 (.BL(BL105),.BLN(BLN105),.WL(WL28));
sram_cell_6t_5 inst_cell_28_106 (.BL(BL106),.BLN(BLN106),.WL(WL28));
sram_cell_6t_5 inst_cell_28_107 (.BL(BL107),.BLN(BLN107),.WL(WL28));
sram_cell_6t_5 inst_cell_28_108 (.BL(BL108),.BLN(BLN108),.WL(WL28));
sram_cell_6t_5 inst_cell_28_109 (.BL(BL109),.BLN(BLN109),.WL(WL28));
sram_cell_6t_5 inst_cell_28_110 (.BL(BL110),.BLN(BLN110),.WL(WL28));
sram_cell_6t_5 inst_cell_28_111 (.BL(BL111),.BLN(BLN111),.WL(WL28));
sram_cell_6t_5 inst_cell_28_112 (.BL(BL112),.BLN(BLN112),.WL(WL28));
sram_cell_6t_5 inst_cell_28_113 (.BL(BL113),.BLN(BLN113),.WL(WL28));
sram_cell_6t_5 inst_cell_28_114 (.BL(BL114),.BLN(BLN114),.WL(WL28));
sram_cell_6t_5 inst_cell_28_115 (.BL(BL115),.BLN(BLN115),.WL(WL28));
sram_cell_6t_5 inst_cell_28_116 (.BL(BL116),.BLN(BLN116),.WL(WL28));
sram_cell_6t_5 inst_cell_28_117 (.BL(BL117),.BLN(BLN117),.WL(WL28));
sram_cell_6t_5 inst_cell_28_118 (.BL(BL118),.BLN(BLN118),.WL(WL28));
sram_cell_6t_5 inst_cell_28_119 (.BL(BL119),.BLN(BLN119),.WL(WL28));
sram_cell_6t_5 inst_cell_28_120 (.BL(BL120),.BLN(BLN120),.WL(WL28));
sram_cell_6t_5 inst_cell_28_121 (.BL(BL121),.BLN(BLN121),.WL(WL28));
sram_cell_6t_5 inst_cell_28_122 (.BL(BL122),.BLN(BLN122),.WL(WL28));
sram_cell_6t_5 inst_cell_28_123 (.BL(BL123),.BLN(BLN123),.WL(WL28));
sram_cell_6t_5 inst_cell_28_124 (.BL(BL124),.BLN(BLN124),.WL(WL28));
sram_cell_6t_5 inst_cell_28_125 (.BL(BL125),.BLN(BLN125),.WL(WL28));
sram_cell_6t_5 inst_cell_28_126 (.BL(BL126),.BLN(BLN126),.WL(WL28));
sram_cell_6t_5 inst_cell_28_127 (.BL(BL127),.BLN(BLN127),.WL(WL28));
sram_cell_6t_5 inst_cell_29_0 (.BL(BL0),.BLN(BLN0),.WL(WL29));
sram_cell_6t_5 inst_cell_29_1 (.BL(BL1),.BLN(BLN1),.WL(WL29));
sram_cell_6t_5 inst_cell_29_2 (.BL(BL2),.BLN(BLN2),.WL(WL29));
sram_cell_6t_5 inst_cell_29_3 (.BL(BL3),.BLN(BLN3),.WL(WL29));
sram_cell_6t_5 inst_cell_29_4 (.BL(BL4),.BLN(BLN4),.WL(WL29));
sram_cell_6t_5 inst_cell_29_5 (.BL(BL5),.BLN(BLN5),.WL(WL29));
sram_cell_6t_5 inst_cell_29_6 (.BL(BL6),.BLN(BLN6),.WL(WL29));
sram_cell_6t_5 inst_cell_29_7 (.BL(BL7),.BLN(BLN7),.WL(WL29));
sram_cell_6t_5 inst_cell_29_8 (.BL(BL8),.BLN(BLN8),.WL(WL29));
sram_cell_6t_5 inst_cell_29_9 (.BL(BL9),.BLN(BLN9),.WL(WL29));
sram_cell_6t_5 inst_cell_29_10 (.BL(BL10),.BLN(BLN10),.WL(WL29));
sram_cell_6t_5 inst_cell_29_11 (.BL(BL11),.BLN(BLN11),.WL(WL29));
sram_cell_6t_5 inst_cell_29_12 (.BL(BL12),.BLN(BLN12),.WL(WL29));
sram_cell_6t_5 inst_cell_29_13 (.BL(BL13),.BLN(BLN13),.WL(WL29));
sram_cell_6t_5 inst_cell_29_14 (.BL(BL14),.BLN(BLN14),.WL(WL29));
sram_cell_6t_5 inst_cell_29_15 (.BL(BL15),.BLN(BLN15),.WL(WL29));
sram_cell_6t_5 inst_cell_29_16 (.BL(BL16),.BLN(BLN16),.WL(WL29));
sram_cell_6t_5 inst_cell_29_17 (.BL(BL17),.BLN(BLN17),.WL(WL29));
sram_cell_6t_5 inst_cell_29_18 (.BL(BL18),.BLN(BLN18),.WL(WL29));
sram_cell_6t_5 inst_cell_29_19 (.BL(BL19),.BLN(BLN19),.WL(WL29));
sram_cell_6t_5 inst_cell_29_20 (.BL(BL20),.BLN(BLN20),.WL(WL29));
sram_cell_6t_5 inst_cell_29_21 (.BL(BL21),.BLN(BLN21),.WL(WL29));
sram_cell_6t_5 inst_cell_29_22 (.BL(BL22),.BLN(BLN22),.WL(WL29));
sram_cell_6t_5 inst_cell_29_23 (.BL(BL23),.BLN(BLN23),.WL(WL29));
sram_cell_6t_5 inst_cell_29_24 (.BL(BL24),.BLN(BLN24),.WL(WL29));
sram_cell_6t_5 inst_cell_29_25 (.BL(BL25),.BLN(BLN25),.WL(WL29));
sram_cell_6t_5 inst_cell_29_26 (.BL(BL26),.BLN(BLN26),.WL(WL29));
sram_cell_6t_5 inst_cell_29_27 (.BL(BL27),.BLN(BLN27),.WL(WL29));
sram_cell_6t_5 inst_cell_29_28 (.BL(BL28),.BLN(BLN28),.WL(WL29));
sram_cell_6t_5 inst_cell_29_29 (.BL(BL29),.BLN(BLN29),.WL(WL29));
sram_cell_6t_5 inst_cell_29_30 (.BL(BL30),.BLN(BLN30),.WL(WL29));
sram_cell_6t_5 inst_cell_29_31 (.BL(BL31),.BLN(BLN31),.WL(WL29));
sram_cell_6t_5 inst_cell_29_32 (.BL(BL32),.BLN(BLN32),.WL(WL29));
sram_cell_6t_5 inst_cell_29_33 (.BL(BL33),.BLN(BLN33),.WL(WL29));
sram_cell_6t_5 inst_cell_29_34 (.BL(BL34),.BLN(BLN34),.WL(WL29));
sram_cell_6t_5 inst_cell_29_35 (.BL(BL35),.BLN(BLN35),.WL(WL29));
sram_cell_6t_5 inst_cell_29_36 (.BL(BL36),.BLN(BLN36),.WL(WL29));
sram_cell_6t_5 inst_cell_29_37 (.BL(BL37),.BLN(BLN37),.WL(WL29));
sram_cell_6t_5 inst_cell_29_38 (.BL(BL38),.BLN(BLN38),.WL(WL29));
sram_cell_6t_5 inst_cell_29_39 (.BL(BL39),.BLN(BLN39),.WL(WL29));
sram_cell_6t_5 inst_cell_29_40 (.BL(BL40),.BLN(BLN40),.WL(WL29));
sram_cell_6t_5 inst_cell_29_41 (.BL(BL41),.BLN(BLN41),.WL(WL29));
sram_cell_6t_5 inst_cell_29_42 (.BL(BL42),.BLN(BLN42),.WL(WL29));
sram_cell_6t_5 inst_cell_29_43 (.BL(BL43),.BLN(BLN43),.WL(WL29));
sram_cell_6t_5 inst_cell_29_44 (.BL(BL44),.BLN(BLN44),.WL(WL29));
sram_cell_6t_5 inst_cell_29_45 (.BL(BL45),.BLN(BLN45),.WL(WL29));
sram_cell_6t_5 inst_cell_29_46 (.BL(BL46),.BLN(BLN46),.WL(WL29));
sram_cell_6t_5 inst_cell_29_47 (.BL(BL47),.BLN(BLN47),.WL(WL29));
sram_cell_6t_5 inst_cell_29_48 (.BL(BL48),.BLN(BLN48),.WL(WL29));
sram_cell_6t_5 inst_cell_29_49 (.BL(BL49),.BLN(BLN49),.WL(WL29));
sram_cell_6t_5 inst_cell_29_50 (.BL(BL50),.BLN(BLN50),.WL(WL29));
sram_cell_6t_5 inst_cell_29_51 (.BL(BL51),.BLN(BLN51),.WL(WL29));
sram_cell_6t_5 inst_cell_29_52 (.BL(BL52),.BLN(BLN52),.WL(WL29));
sram_cell_6t_5 inst_cell_29_53 (.BL(BL53),.BLN(BLN53),.WL(WL29));
sram_cell_6t_5 inst_cell_29_54 (.BL(BL54),.BLN(BLN54),.WL(WL29));
sram_cell_6t_5 inst_cell_29_55 (.BL(BL55),.BLN(BLN55),.WL(WL29));
sram_cell_6t_5 inst_cell_29_56 (.BL(BL56),.BLN(BLN56),.WL(WL29));
sram_cell_6t_5 inst_cell_29_57 (.BL(BL57),.BLN(BLN57),.WL(WL29));
sram_cell_6t_5 inst_cell_29_58 (.BL(BL58),.BLN(BLN58),.WL(WL29));
sram_cell_6t_5 inst_cell_29_59 (.BL(BL59),.BLN(BLN59),.WL(WL29));
sram_cell_6t_5 inst_cell_29_60 (.BL(BL60),.BLN(BLN60),.WL(WL29));
sram_cell_6t_5 inst_cell_29_61 (.BL(BL61),.BLN(BLN61),.WL(WL29));
sram_cell_6t_5 inst_cell_29_62 (.BL(BL62),.BLN(BLN62),.WL(WL29));
sram_cell_6t_5 inst_cell_29_63 (.BL(BL63),.BLN(BLN63),.WL(WL29));
sram_cell_6t_5 inst_cell_29_64 (.BL(BL64),.BLN(BLN64),.WL(WL29));
sram_cell_6t_5 inst_cell_29_65 (.BL(BL65),.BLN(BLN65),.WL(WL29));
sram_cell_6t_5 inst_cell_29_66 (.BL(BL66),.BLN(BLN66),.WL(WL29));
sram_cell_6t_5 inst_cell_29_67 (.BL(BL67),.BLN(BLN67),.WL(WL29));
sram_cell_6t_5 inst_cell_29_68 (.BL(BL68),.BLN(BLN68),.WL(WL29));
sram_cell_6t_5 inst_cell_29_69 (.BL(BL69),.BLN(BLN69),.WL(WL29));
sram_cell_6t_5 inst_cell_29_70 (.BL(BL70),.BLN(BLN70),.WL(WL29));
sram_cell_6t_5 inst_cell_29_71 (.BL(BL71),.BLN(BLN71),.WL(WL29));
sram_cell_6t_5 inst_cell_29_72 (.BL(BL72),.BLN(BLN72),.WL(WL29));
sram_cell_6t_5 inst_cell_29_73 (.BL(BL73),.BLN(BLN73),.WL(WL29));
sram_cell_6t_5 inst_cell_29_74 (.BL(BL74),.BLN(BLN74),.WL(WL29));
sram_cell_6t_5 inst_cell_29_75 (.BL(BL75),.BLN(BLN75),.WL(WL29));
sram_cell_6t_5 inst_cell_29_76 (.BL(BL76),.BLN(BLN76),.WL(WL29));
sram_cell_6t_5 inst_cell_29_77 (.BL(BL77),.BLN(BLN77),.WL(WL29));
sram_cell_6t_5 inst_cell_29_78 (.BL(BL78),.BLN(BLN78),.WL(WL29));
sram_cell_6t_5 inst_cell_29_79 (.BL(BL79),.BLN(BLN79),.WL(WL29));
sram_cell_6t_5 inst_cell_29_80 (.BL(BL80),.BLN(BLN80),.WL(WL29));
sram_cell_6t_5 inst_cell_29_81 (.BL(BL81),.BLN(BLN81),.WL(WL29));
sram_cell_6t_5 inst_cell_29_82 (.BL(BL82),.BLN(BLN82),.WL(WL29));
sram_cell_6t_5 inst_cell_29_83 (.BL(BL83),.BLN(BLN83),.WL(WL29));
sram_cell_6t_5 inst_cell_29_84 (.BL(BL84),.BLN(BLN84),.WL(WL29));
sram_cell_6t_5 inst_cell_29_85 (.BL(BL85),.BLN(BLN85),.WL(WL29));
sram_cell_6t_5 inst_cell_29_86 (.BL(BL86),.BLN(BLN86),.WL(WL29));
sram_cell_6t_5 inst_cell_29_87 (.BL(BL87),.BLN(BLN87),.WL(WL29));
sram_cell_6t_5 inst_cell_29_88 (.BL(BL88),.BLN(BLN88),.WL(WL29));
sram_cell_6t_5 inst_cell_29_89 (.BL(BL89),.BLN(BLN89),.WL(WL29));
sram_cell_6t_5 inst_cell_29_90 (.BL(BL90),.BLN(BLN90),.WL(WL29));
sram_cell_6t_5 inst_cell_29_91 (.BL(BL91),.BLN(BLN91),.WL(WL29));
sram_cell_6t_5 inst_cell_29_92 (.BL(BL92),.BLN(BLN92),.WL(WL29));
sram_cell_6t_5 inst_cell_29_93 (.BL(BL93),.BLN(BLN93),.WL(WL29));
sram_cell_6t_5 inst_cell_29_94 (.BL(BL94),.BLN(BLN94),.WL(WL29));
sram_cell_6t_5 inst_cell_29_95 (.BL(BL95),.BLN(BLN95),.WL(WL29));
sram_cell_6t_5 inst_cell_29_96 (.BL(BL96),.BLN(BLN96),.WL(WL29));
sram_cell_6t_5 inst_cell_29_97 (.BL(BL97),.BLN(BLN97),.WL(WL29));
sram_cell_6t_5 inst_cell_29_98 (.BL(BL98),.BLN(BLN98),.WL(WL29));
sram_cell_6t_5 inst_cell_29_99 (.BL(BL99),.BLN(BLN99),.WL(WL29));
sram_cell_6t_5 inst_cell_29_100 (.BL(BL100),.BLN(BLN100),.WL(WL29));
sram_cell_6t_5 inst_cell_29_101 (.BL(BL101),.BLN(BLN101),.WL(WL29));
sram_cell_6t_5 inst_cell_29_102 (.BL(BL102),.BLN(BLN102),.WL(WL29));
sram_cell_6t_5 inst_cell_29_103 (.BL(BL103),.BLN(BLN103),.WL(WL29));
sram_cell_6t_5 inst_cell_29_104 (.BL(BL104),.BLN(BLN104),.WL(WL29));
sram_cell_6t_5 inst_cell_29_105 (.BL(BL105),.BLN(BLN105),.WL(WL29));
sram_cell_6t_5 inst_cell_29_106 (.BL(BL106),.BLN(BLN106),.WL(WL29));
sram_cell_6t_5 inst_cell_29_107 (.BL(BL107),.BLN(BLN107),.WL(WL29));
sram_cell_6t_5 inst_cell_29_108 (.BL(BL108),.BLN(BLN108),.WL(WL29));
sram_cell_6t_5 inst_cell_29_109 (.BL(BL109),.BLN(BLN109),.WL(WL29));
sram_cell_6t_5 inst_cell_29_110 (.BL(BL110),.BLN(BLN110),.WL(WL29));
sram_cell_6t_5 inst_cell_29_111 (.BL(BL111),.BLN(BLN111),.WL(WL29));
sram_cell_6t_5 inst_cell_29_112 (.BL(BL112),.BLN(BLN112),.WL(WL29));
sram_cell_6t_5 inst_cell_29_113 (.BL(BL113),.BLN(BLN113),.WL(WL29));
sram_cell_6t_5 inst_cell_29_114 (.BL(BL114),.BLN(BLN114),.WL(WL29));
sram_cell_6t_5 inst_cell_29_115 (.BL(BL115),.BLN(BLN115),.WL(WL29));
sram_cell_6t_5 inst_cell_29_116 (.BL(BL116),.BLN(BLN116),.WL(WL29));
sram_cell_6t_5 inst_cell_29_117 (.BL(BL117),.BLN(BLN117),.WL(WL29));
sram_cell_6t_5 inst_cell_29_118 (.BL(BL118),.BLN(BLN118),.WL(WL29));
sram_cell_6t_5 inst_cell_29_119 (.BL(BL119),.BLN(BLN119),.WL(WL29));
sram_cell_6t_5 inst_cell_29_120 (.BL(BL120),.BLN(BLN120),.WL(WL29));
sram_cell_6t_5 inst_cell_29_121 (.BL(BL121),.BLN(BLN121),.WL(WL29));
sram_cell_6t_5 inst_cell_29_122 (.BL(BL122),.BLN(BLN122),.WL(WL29));
sram_cell_6t_5 inst_cell_29_123 (.BL(BL123),.BLN(BLN123),.WL(WL29));
sram_cell_6t_5 inst_cell_29_124 (.BL(BL124),.BLN(BLN124),.WL(WL29));
sram_cell_6t_5 inst_cell_29_125 (.BL(BL125),.BLN(BLN125),.WL(WL29));
sram_cell_6t_5 inst_cell_29_126 (.BL(BL126),.BLN(BLN126),.WL(WL29));
sram_cell_6t_5 inst_cell_29_127 (.BL(BL127),.BLN(BLN127),.WL(WL29));
sram_cell_6t_5 inst_cell_30_0 (.BL(BL0),.BLN(BLN0),.WL(WL30));
sram_cell_6t_5 inst_cell_30_1 (.BL(BL1),.BLN(BLN1),.WL(WL30));
sram_cell_6t_5 inst_cell_30_2 (.BL(BL2),.BLN(BLN2),.WL(WL30));
sram_cell_6t_5 inst_cell_30_3 (.BL(BL3),.BLN(BLN3),.WL(WL30));
sram_cell_6t_5 inst_cell_30_4 (.BL(BL4),.BLN(BLN4),.WL(WL30));
sram_cell_6t_5 inst_cell_30_5 (.BL(BL5),.BLN(BLN5),.WL(WL30));
sram_cell_6t_5 inst_cell_30_6 (.BL(BL6),.BLN(BLN6),.WL(WL30));
sram_cell_6t_5 inst_cell_30_7 (.BL(BL7),.BLN(BLN7),.WL(WL30));
sram_cell_6t_5 inst_cell_30_8 (.BL(BL8),.BLN(BLN8),.WL(WL30));
sram_cell_6t_5 inst_cell_30_9 (.BL(BL9),.BLN(BLN9),.WL(WL30));
sram_cell_6t_5 inst_cell_30_10 (.BL(BL10),.BLN(BLN10),.WL(WL30));
sram_cell_6t_5 inst_cell_30_11 (.BL(BL11),.BLN(BLN11),.WL(WL30));
sram_cell_6t_5 inst_cell_30_12 (.BL(BL12),.BLN(BLN12),.WL(WL30));
sram_cell_6t_5 inst_cell_30_13 (.BL(BL13),.BLN(BLN13),.WL(WL30));
sram_cell_6t_5 inst_cell_30_14 (.BL(BL14),.BLN(BLN14),.WL(WL30));
sram_cell_6t_5 inst_cell_30_15 (.BL(BL15),.BLN(BLN15),.WL(WL30));
sram_cell_6t_5 inst_cell_30_16 (.BL(BL16),.BLN(BLN16),.WL(WL30));
sram_cell_6t_5 inst_cell_30_17 (.BL(BL17),.BLN(BLN17),.WL(WL30));
sram_cell_6t_5 inst_cell_30_18 (.BL(BL18),.BLN(BLN18),.WL(WL30));
sram_cell_6t_5 inst_cell_30_19 (.BL(BL19),.BLN(BLN19),.WL(WL30));
sram_cell_6t_5 inst_cell_30_20 (.BL(BL20),.BLN(BLN20),.WL(WL30));
sram_cell_6t_5 inst_cell_30_21 (.BL(BL21),.BLN(BLN21),.WL(WL30));
sram_cell_6t_5 inst_cell_30_22 (.BL(BL22),.BLN(BLN22),.WL(WL30));
sram_cell_6t_5 inst_cell_30_23 (.BL(BL23),.BLN(BLN23),.WL(WL30));
sram_cell_6t_5 inst_cell_30_24 (.BL(BL24),.BLN(BLN24),.WL(WL30));
sram_cell_6t_5 inst_cell_30_25 (.BL(BL25),.BLN(BLN25),.WL(WL30));
sram_cell_6t_5 inst_cell_30_26 (.BL(BL26),.BLN(BLN26),.WL(WL30));
sram_cell_6t_5 inst_cell_30_27 (.BL(BL27),.BLN(BLN27),.WL(WL30));
sram_cell_6t_5 inst_cell_30_28 (.BL(BL28),.BLN(BLN28),.WL(WL30));
sram_cell_6t_5 inst_cell_30_29 (.BL(BL29),.BLN(BLN29),.WL(WL30));
sram_cell_6t_5 inst_cell_30_30 (.BL(BL30),.BLN(BLN30),.WL(WL30));
sram_cell_6t_5 inst_cell_30_31 (.BL(BL31),.BLN(BLN31),.WL(WL30));
sram_cell_6t_5 inst_cell_30_32 (.BL(BL32),.BLN(BLN32),.WL(WL30));
sram_cell_6t_5 inst_cell_30_33 (.BL(BL33),.BLN(BLN33),.WL(WL30));
sram_cell_6t_5 inst_cell_30_34 (.BL(BL34),.BLN(BLN34),.WL(WL30));
sram_cell_6t_5 inst_cell_30_35 (.BL(BL35),.BLN(BLN35),.WL(WL30));
sram_cell_6t_5 inst_cell_30_36 (.BL(BL36),.BLN(BLN36),.WL(WL30));
sram_cell_6t_5 inst_cell_30_37 (.BL(BL37),.BLN(BLN37),.WL(WL30));
sram_cell_6t_5 inst_cell_30_38 (.BL(BL38),.BLN(BLN38),.WL(WL30));
sram_cell_6t_5 inst_cell_30_39 (.BL(BL39),.BLN(BLN39),.WL(WL30));
sram_cell_6t_5 inst_cell_30_40 (.BL(BL40),.BLN(BLN40),.WL(WL30));
sram_cell_6t_5 inst_cell_30_41 (.BL(BL41),.BLN(BLN41),.WL(WL30));
sram_cell_6t_5 inst_cell_30_42 (.BL(BL42),.BLN(BLN42),.WL(WL30));
sram_cell_6t_5 inst_cell_30_43 (.BL(BL43),.BLN(BLN43),.WL(WL30));
sram_cell_6t_5 inst_cell_30_44 (.BL(BL44),.BLN(BLN44),.WL(WL30));
sram_cell_6t_5 inst_cell_30_45 (.BL(BL45),.BLN(BLN45),.WL(WL30));
sram_cell_6t_5 inst_cell_30_46 (.BL(BL46),.BLN(BLN46),.WL(WL30));
sram_cell_6t_5 inst_cell_30_47 (.BL(BL47),.BLN(BLN47),.WL(WL30));
sram_cell_6t_5 inst_cell_30_48 (.BL(BL48),.BLN(BLN48),.WL(WL30));
sram_cell_6t_5 inst_cell_30_49 (.BL(BL49),.BLN(BLN49),.WL(WL30));
sram_cell_6t_5 inst_cell_30_50 (.BL(BL50),.BLN(BLN50),.WL(WL30));
sram_cell_6t_5 inst_cell_30_51 (.BL(BL51),.BLN(BLN51),.WL(WL30));
sram_cell_6t_5 inst_cell_30_52 (.BL(BL52),.BLN(BLN52),.WL(WL30));
sram_cell_6t_5 inst_cell_30_53 (.BL(BL53),.BLN(BLN53),.WL(WL30));
sram_cell_6t_5 inst_cell_30_54 (.BL(BL54),.BLN(BLN54),.WL(WL30));
sram_cell_6t_5 inst_cell_30_55 (.BL(BL55),.BLN(BLN55),.WL(WL30));
sram_cell_6t_5 inst_cell_30_56 (.BL(BL56),.BLN(BLN56),.WL(WL30));
sram_cell_6t_5 inst_cell_30_57 (.BL(BL57),.BLN(BLN57),.WL(WL30));
sram_cell_6t_5 inst_cell_30_58 (.BL(BL58),.BLN(BLN58),.WL(WL30));
sram_cell_6t_5 inst_cell_30_59 (.BL(BL59),.BLN(BLN59),.WL(WL30));
sram_cell_6t_5 inst_cell_30_60 (.BL(BL60),.BLN(BLN60),.WL(WL30));
sram_cell_6t_5 inst_cell_30_61 (.BL(BL61),.BLN(BLN61),.WL(WL30));
sram_cell_6t_5 inst_cell_30_62 (.BL(BL62),.BLN(BLN62),.WL(WL30));
sram_cell_6t_5 inst_cell_30_63 (.BL(BL63),.BLN(BLN63),.WL(WL30));
sram_cell_6t_5 inst_cell_30_64 (.BL(BL64),.BLN(BLN64),.WL(WL30));
sram_cell_6t_5 inst_cell_30_65 (.BL(BL65),.BLN(BLN65),.WL(WL30));
sram_cell_6t_5 inst_cell_30_66 (.BL(BL66),.BLN(BLN66),.WL(WL30));
sram_cell_6t_5 inst_cell_30_67 (.BL(BL67),.BLN(BLN67),.WL(WL30));
sram_cell_6t_5 inst_cell_30_68 (.BL(BL68),.BLN(BLN68),.WL(WL30));
sram_cell_6t_5 inst_cell_30_69 (.BL(BL69),.BLN(BLN69),.WL(WL30));
sram_cell_6t_5 inst_cell_30_70 (.BL(BL70),.BLN(BLN70),.WL(WL30));
sram_cell_6t_5 inst_cell_30_71 (.BL(BL71),.BLN(BLN71),.WL(WL30));
sram_cell_6t_5 inst_cell_30_72 (.BL(BL72),.BLN(BLN72),.WL(WL30));
sram_cell_6t_5 inst_cell_30_73 (.BL(BL73),.BLN(BLN73),.WL(WL30));
sram_cell_6t_5 inst_cell_30_74 (.BL(BL74),.BLN(BLN74),.WL(WL30));
sram_cell_6t_5 inst_cell_30_75 (.BL(BL75),.BLN(BLN75),.WL(WL30));
sram_cell_6t_5 inst_cell_30_76 (.BL(BL76),.BLN(BLN76),.WL(WL30));
sram_cell_6t_5 inst_cell_30_77 (.BL(BL77),.BLN(BLN77),.WL(WL30));
sram_cell_6t_5 inst_cell_30_78 (.BL(BL78),.BLN(BLN78),.WL(WL30));
sram_cell_6t_5 inst_cell_30_79 (.BL(BL79),.BLN(BLN79),.WL(WL30));
sram_cell_6t_5 inst_cell_30_80 (.BL(BL80),.BLN(BLN80),.WL(WL30));
sram_cell_6t_5 inst_cell_30_81 (.BL(BL81),.BLN(BLN81),.WL(WL30));
sram_cell_6t_5 inst_cell_30_82 (.BL(BL82),.BLN(BLN82),.WL(WL30));
sram_cell_6t_5 inst_cell_30_83 (.BL(BL83),.BLN(BLN83),.WL(WL30));
sram_cell_6t_5 inst_cell_30_84 (.BL(BL84),.BLN(BLN84),.WL(WL30));
sram_cell_6t_5 inst_cell_30_85 (.BL(BL85),.BLN(BLN85),.WL(WL30));
sram_cell_6t_5 inst_cell_30_86 (.BL(BL86),.BLN(BLN86),.WL(WL30));
sram_cell_6t_5 inst_cell_30_87 (.BL(BL87),.BLN(BLN87),.WL(WL30));
sram_cell_6t_5 inst_cell_30_88 (.BL(BL88),.BLN(BLN88),.WL(WL30));
sram_cell_6t_5 inst_cell_30_89 (.BL(BL89),.BLN(BLN89),.WL(WL30));
sram_cell_6t_5 inst_cell_30_90 (.BL(BL90),.BLN(BLN90),.WL(WL30));
sram_cell_6t_5 inst_cell_30_91 (.BL(BL91),.BLN(BLN91),.WL(WL30));
sram_cell_6t_5 inst_cell_30_92 (.BL(BL92),.BLN(BLN92),.WL(WL30));
sram_cell_6t_5 inst_cell_30_93 (.BL(BL93),.BLN(BLN93),.WL(WL30));
sram_cell_6t_5 inst_cell_30_94 (.BL(BL94),.BLN(BLN94),.WL(WL30));
sram_cell_6t_5 inst_cell_30_95 (.BL(BL95),.BLN(BLN95),.WL(WL30));
sram_cell_6t_5 inst_cell_30_96 (.BL(BL96),.BLN(BLN96),.WL(WL30));
sram_cell_6t_5 inst_cell_30_97 (.BL(BL97),.BLN(BLN97),.WL(WL30));
sram_cell_6t_5 inst_cell_30_98 (.BL(BL98),.BLN(BLN98),.WL(WL30));
sram_cell_6t_5 inst_cell_30_99 (.BL(BL99),.BLN(BLN99),.WL(WL30));
sram_cell_6t_5 inst_cell_30_100 (.BL(BL100),.BLN(BLN100),.WL(WL30));
sram_cell_6t_5 inst_cell_30_101 (.BL(BL101),.BLN(BLN101),.WL(WL30));
sram_cell_6t_5 inst_cell_30_102 (.BL(BL102),.BLN(BLN102),.WL(WL30));
sram_cell_6t_5 inst_cell_30_103 (.BL(BL103),.BLN(BLN103),.WL(WL30));
sram_cell_6t_5 inst_cell_30_104 (.BL(BL104),.BLN(BLN104),.WL(WL30));
sram_cell_6t_5 inst_cell_30_105 (.BL(BL105),.BLN(BLN105),.WL(WL30));
sram_cell_6t_5 inst_cell_30_106 (.BL(BL106),.BLN(BLN106),.WL(WL30));
sram_cell_6t_5 inst_cell_30_107 (.BL(BL107),.BLN(BLN107),.WL(WL30));
sram_cell_6t_5 inst_cell_30_108 (.BL(BL108),.BLN(BLN108),.WL(WL30));
sram_cell_6t_5 inst_cell_30_109 (.BL(BL109),.BLN(BLN109),.WL(WL30));
sram_cell_6t_5 inst_cell_30_110 (.BL(BL110),.BLN(BLN110),.WL(WL30));
sram_cell_6t_5 inst_cell_30_111 (.BL(BL111),.BLN(BLN111),.WL(WL30));
sram_cell_6t_5 inst_cell_30_112 (.BL(BL112),.BLN(BLN112),.WL(WL30));
sram_cell_6t_5 inst_cell_30_113 (.BL(BL113),.BLN(BLN113),.WL(WL30));
sram_cell_6t_5 inst_cell_30_114 (.BL(BL114),.BLN(BLN114),.WL(WL30));
sram_cell_6t_5 inst_cell_30_115 (.BL(BL115),.BLN(BLN115),.WL(WL30));
sram_cell_6t_5 inst_cell_30_116 (.BL(BL116),.BLN(BLN116),.WL(WL30));
sram_cell_6t_5 inst_cell_30_117 (.BL(BL117),.BLN(BLN117),.WL(WL30));
sram_cell_6t_5 inst_cell_30_118 (.BL(BL118),.BLN(BLN118),.WL(WL30));
sram_cell_6t_5 inst_cell_30_119 (.BL(BL119),.BLN(BLN119),.WL(WL30));
sram_cell_6t_5 inst_cell_30_120 (.BL(BL120),.BLN(BLN120),.WL(WL30));
sram_cell_6t_5 inst_cell_30_121 (.BL(BL121),.BLN(BLN121),.WL(WL30));
sram_cell_6t_5 inst_cell_30_122 (.BL(BL122),.BLN(BLN122),.WL(WL30));
sram_cell_6t_5 inst_cell_30_123 (.BL(BL123),.BLN(BLN123),.WL(WL30));
sram_cell_6t_5 inst_cell_30_124 (.BL(BL124),.BLN(BLN124),.WL(WL30));
sram_cell_6t_5 inst_cell_30_125 (.BL(BL125),.BLN(BLN125),.WL(WL30));
sram_cell_6t_5 inst_cell_30_126 (.BL(BL126),.BLN(BLN126),.WL(WL30));
sram_cell_6t_5 inst_cell_30_127 (.BL(BL127),.BLN(BLN127),.WL(WL30));
sram_cell_6t_5 inst_cell_31_0 (.BL(BL0),.BLN(BLN0),.WL(WL31));
sram_cell_6t_5 inst_cell_31_1 (.BL(BL1),.BLN(BLN1),.WL(WL31));
sram_cell_6t_5 inst_cell_31_2 (.BL(BL2),.BLN(BLN2),.WL(WL31));
sram_cell_6t_5 inst_cell_31_3 (.BL(BL3),.BLN(BLN3),.WL(WL31));
sram_cell_6t_5 inst_cell_31_4 (.BL(BL4),.BLN(BLN4),.WL(WL31));
sram_cell_6t_5 inst_cell_31_5 (.BL(BL5),.BLN(BLN5),.WL(WL31));
sram_cell_6t_5 inst_cell_31_6 (.BL(BL6),.BLN(BLN6),.WL(WL31));
sram_cell_6t_5 inst_cell_31_7 (.BL(BL7),.BLN(BLN7),.WL(WL31));
sram_cell_6t_5 inst_cell_31_8 (.BL(BL8),.BLN(BLN8),.WL(WL31));
sram_cell_6t_5 inst_cell_31_9 (.BL(BL9),.BLN(BLN9),.WL(WL31));
sram_cell_6t_5 inst_cell_31_10 (.BL(BL10),.BLN(BLN10),.WL(WL31));
sram_cell_6t_5 inst_cell_31_11 (.BL(BL11),.BLN(BLN11),.WL(WL31));
sram_cell_6t_5 inst_cell_31_12 (.BL(BL12),.BLN(BLN12),.WL(WL31));
sram_cell_6t_5 inst_cell_31_13 (.BL(BL13),.BLN(BLN13),.WL(WL31));
sram_cell_6t_5 inst_cell_31_14 (.BL(BL14),.BLN(BLN14),.WL(WL31));
sram_cell_6t_5 inst_cell_31_15 (.BL(BL15),.BLN(BLN15),.WL(WL31));
sram_cell_6t_5 inst_cell_31_16 (.BL(BL16),.BLN(BLN16),.WL(WL31));
sram_cell_6t_5 inst_cell_31_17 (.BL(BL17),.BLN(BLN17),.WL(WL31));
sram_cell_6t_5 inst_cell_31_18 (.BL(BL18),.BLN(BLN18),.WL(WL31));
sram_cell_6t_5 inst_cell_31_19 (.BL(BL19),.BLN(BLN19),.WL(WL31));
sram_cell_6t_5 inst_cell_31_20 (.BL(BL20),.BLN(BLN20),.WL(WL31));
sram_cell_6t_5 inst_cell_31_21 (.BL(BL21),.BLN(BLN21),.WL(WL31));
sram_cell_6t_5 inst_cell_31_22 (.BL(BL22),.BLN(BLN22),.WL(WL31));
sram_cell_6t_5 inst_cell_31_23 (.BL(BL23),.BLN(BLN23),.WL(WL31));
sram_cell_6t_5 inst_cell_31_24 (.BL(BL24),.BLN(BLN24),.WL(WL31));
sram_cell_6t_5 inst_cell_31_25 (.BL(BL25),.BLN(BLN25),.WL(WL31));
sram_cell_6t_5 inst_cell_31_26 (.BL(BL26),.BLN(BLN26),.WL(WL31));
sram_cell_6t_5 inst_cell_31_27 (.BL(BL27),.BLN(BLN27),.WL(WL31));
sram_cell_6t_5 inst_cell_31_28 (.BL(BL28),.BLN(BLN28),.WL(WL31));
sram_cell_6t_5 inst_cell_31_29 (.BL(BL29),.BLN(BLN29),.WL(WL31));
sram_cell_6t_5 inst_cell_31_30 (.BL(BL30),.BLN(BLN30),.WL(WL31));
sram_cell_6t_5 inst_cell_31_31 (.BL(BL31),.BLN(BLN31),.WL(WL31));
sram_cell_6t_5 inst_cell_31_32 (.BL(BL32),.BLN(BLN32),.WL(WL31));
sram_cell_6t_5 inst_cell_31_33 (.BL(BL33),.BLN(BLN33),.WL(WL31));
sram_cell_6t_5 inst_cell_31_34 (.BL(BL34),.BLN(BLN34),.WL(WL31));
sram_cell_6t_5 inst_cell_31_35 (.BL(BL35),.BLN(BLN35),.WL(WL31));
sram_cell_6t_5 inst_cell_31_36 (.BL(BL36),.BLN(BLN36),.WL(WL31));
sram_cell_6t_5 inst_cell_31_37 (.BL(BL37),.BLN(BLN37),.WL(WL31));
sram_cell_6t_5 inst_cell_31_38 (.BL(BL38),.BLN(BLN38),.WL(WL31));
sram_cell_6t_5 inst_cell_31_39 (.BL(BL39),.BLN(BLN39),.WL(WL31));
sram_cell_6t_5 inst_cell_31_40 (.BL(BL40),.BLN(BLN40),.WL(WL31));
sram_cell_6t_5 inst_cell_31_41 (.BL(BL41),.BLN(BLN41),.WL(WL31));
sram_cell_6t_5 inst_cell_31_42 (.BL(BL42),.BLN(BLN42),.WL(WL31));
sram_cell_6t_5 inst_cell_31_43 (.BL(BL43),.BLN(BLN43),.WL(WL31));
sram_cell_6t_5 inst_cell_31_44 (.BL(BL44),.BLN(BLN44),.WL(WL31));
sram_cell_6t_5 inst_cell_31_45 (.BL(BL45),.BLN(BLN45),.WL(WL31));
sram_cell_6t_5 inst_cell_31_46 (.BL(BL46),.BLN(BLN46),.WL(WL31));
sram_cell_6t_5 inst_cell_31_47 (.BL(BL47),.BLN(BLN47),.WL(WL31));
sram_cell_6t_5 inst_cell_31_48 (.BL(BL48),.BLN(BLN48),.WL(WL31));
sram_cell_6t_5 inst_cell_31_49 (.BL(BL49),.BLN(BLN49),.WL(WL31));
sram_cell_6t_5 inst_cell_31_50 (.BL(BL50),.BLN(BLN50),.WL(WL31));
sram_cell_6t_5 inst_cell_31_51 (.BL(BL51),.BLN(BLN51),.WL(WL31));
sram_cell_6t_5 inst_cell_31_52 (.BL(BL52),.BLN(BLN52),.WL(WL31));
sram_cell_6t_5 inst_cell_31_53 (.BL(BL53),.BLN(BLN53),.WL(WL31));
sram_cell_6t_5 inst_cell_31_54 (.BL(BL54),.BLN(BLN54),.WL(WL31));
sram_cell_6t_5 inst_cell_31_55 (.BL(BL55),.BLN(BLN55),.WL(WL31));
sram_cell_6t_5 inst_cell_31_56 (.BL(BL56),.BLN(BLN56),.WL(WL31));
sram_cell_6t_5 inst_cell_31_57 (.BL(BL57),.BLN(BLN57),.WL(WL31));
sram_cell_6t_5 inst_cell_31_58 (.BL(BL58),.BLN(BLN58),.WL(WL31));
sram_cell_6t_5 inst_cell_31_59 (.BL(BL59),.BLN(BLN59),.WL(WL31));
sram_cell_6t_5 inst_cell_31_60 (.BL(BL60),.BLN(BLN60),.WL(WL31));
sram_cell_6t_5 inst_cell_31_61 (.BL(BL61),.BLN(BLN61),.WL(WL31));
sram_cell_6t_5 inst_cell_31_62 (.BL(BL62),.BLN(BLN62),.WL(WL31));
sram_cell_6t_5 inst_cell_31_63 (.BL(BL63),.BLN(BLN63),.WL(WL31));
sram_cell_6t_5 inst_cell_31_64 (.BL(BL64),.BLN(BLN64),.WL(WL31));
sram_cell_6t_5 inst_cell_31_65 (.BL(BL65),.BLN(BLN65),.WL(WL31));
sram_cell_6t_5 inst_cell_31_66 (.BL(BL66),.BLN(BLN66),.WL(WL31));
sram_cell_6t_5 inst_cell_31_67 (.BL(BL67),.BLN(BLN67),.WL(WL31));
sram_cell_6t_5 inst_cell_31_68 (.BL(BL68),.BLN(BLN68),.WL(WL31));
sram_cell_6t_5 inst_cell_31_69 (.BL(BL69),.BLN(BLN69),.WL(WL31));
sram_cell_6t_5 inst_cell_31_70 (.BL(BL70),.BLN(BLN70),.WL(WL31));
sram_cell_6t_5 inst_cell_31_71 (.BL(BL71),.BLN(BLN71),.WL(WL31));
sram_cell_6t_5 inst_cell_31_72 (.BL(BL72),.BLN(BLN72),.WL(WL31));
sram_cell_6t_5 inst_cell_31_73 (.BL(BL73),.BLN(BLN73),.WL(WL31));
sram_cell_6t_5 inst_cell_31_74 (.BL(BL74),.BLN(BLN74),.WL(WL31));
sram_cell_6t_5 inst_cell_31_75 (.BL(BL75),.BLN(BLN75),.WL(WL31));
sram_cell_6t_5 inst_cell_31_76 (.BL(BL76),.BLN(BLN76),.WL(WL31));
sram_cell_6t_5 inst_cell_31_77 (.BL(BL77),.BLN(BLN77),.WL(WL31));
sram_cell_6t_5 inst_cell_31_78 (.BL(BL78),.BLN(BLN78),.WL(WL31));
sram_cell_6t_5 inst_cell_31_79 (.BL(BL79),.BLN(BLN79),.WL(WL31));
sram_cell_6t_5 inst_cell_31_80 (.BL(BL80),.BLN(BLN80),.WL(WL31));
sram_cell_6t_5 inst_cell_31_81 (.BL(BL81),.BLN(BLN81),.WL(WL31));
sram_cell_6t_5 inst_cell_31_82 (.BL(BL82),.BLN(BLN82),.WL(WL31));
sram_cell_6t_5 inst_cell_31_83 (.BL(BL83),.BLN(BLN83),.WL(WL31));
sram_cell_6t_5 inst_cell_31_84 (.BL(BL84),.BLN(BLN84),.WL(WL31));
sram_cell_6t_5 inst_cell_31_85 (.BL(BL85),.BLN(BLN85),.WL(WL31));
sram_cell_6t_5 inst_cell_31_86 (.BL(BL86),.BLN(BLN86),.WL(WL31));
sram_cell_6t_5 inst_cell_31_87 (.BL(BL87),.BLN(BLN87),.WL(WL31));
sram_cell_6t_5 inst_cell_31_88 (.BL(BL88),.BLN(BLN88),.WL(WL31));
sram_cell_6t_5 inst_cell_31_89 (.BL(BL89),.BLN(BLN89),.WL(WL31));
sram_cell_6t_5 inst_cell_31_90 (.BL(BL90),.BLN(BLN90),.WL(WL31));
sram_cell_6t_5 inst_cell_31_91 (.BL(BL91),.BLN(BLN91),.WL(WL31));
sram_cell_6t_5 inst_cell_31_92 (.BL(BL92),.BLN(BLN92),.WL(WL31));
sram_cell_6t_5 inst_cell_31_93 (.BL(BL93),.BLN(BLN93),.WL(WL31));
sram_cell_6t_5 inst_cell_31_94 (.BL(BL94),.BLN(BLN94),.WL(WL31));
sram_cell_6t_5 inst_cell_31_95 (.BL(BL95),.BLN(BLN95),.WL(WL31));
sram_cell_6t_5 inst_cell_31_96 (.BL(BL96),.BLN(BLN96),.WL(WL31));
sram_cell_6t_5 inst_cell_31_97 (.BL(BL97),.BLN(BLN97),.WL(WL31));
sram_cell_6t_5 inst_cell_31_98 (.BL(BL98),.BLN(BLN98),.WL(WL31));
sram_cell_6t_5 inst_cell_31_99 (.BL(BL99),.BLN(BLN99),.WL(WL31));
sram_cell_6t_5 inst_cell_31_100 (.BL(BL100),.BLN(BLN100),.WL(WL31));
sram_cell_6t_5 inst_cell_31_101 (.BL(BL101),.BLN(BLN101),.WL(WL31));
sram_cell_6t_5 inst_cell_31_102 (.BL(BL102),.BLN(BLN102),.WL(WL31));
sram_cell_6t_5 inst_cell_31_103 (.BL(BL103),.BLN(BLN103),.WL(WL31));
sram_cell_6t_5 inst_cell_31_104 (.BL(BL104),.BLN(BLN104),.WL(WL31));
sram_cell_6t_5 inst_cell_31_105 (.BL(BL105),.BLN(BLN105),.WL(WL31));
sram_cell_6t_5 inst_cell_31_106 (.BL(BL106),.BLN(BLN106),.WL(WL31));
sram_cell_6t_5 inst_cell_31_107 (.BL(BL107),.BLN(BLN107),.WL(WL31));
sram_cell_6t_5 inst_cell_31_108 (.BL(BL108),.BLN(BLN108),.WL(WL31));
sram_cell_6t_5 inst_cell_31_109 (.BL(BL109),.BLN(BLN109),.WL(WL31));
sram_cell_6t_5 inst_cell_31_110 (.BL(BL110),.BLN(BLN110),.WL(WL31));
sram_cell_6t_5 inst_cell_31_111 (.BL(BL111),.BLN(BLN111),.WL(WL31));
sram_cell_6t_5 inst_cell_31_112 (.BL(BL112),.BLN(BLN112),.WL(WL31));
sram_cell_6t_5 inst_cell_31_113 (.BL(BL113),.BLN(BLN113),.WL(WL31));
sram_cell_6t_5 inst_cell_31_114 (.BL(BL114),.BLN(BLN114),.WL(WL31));
sram_cell_6t_5 inst_cell_31_115 (.BL(BL115),.BLN(BLN115),.WL(WL31));
sram_cell_6t_5 inst_cell_31_116 (.BL(BL116),.BLN(BLN116),.WL(WL31));
sram_cell_6t_5 inst_cell_31_117 (.BL(BL117),.BLN(BLN117),.WL(WL31));
sram_cell_6t_5 inst_cell_31_118 (.BL(BL118),.BLN(BLN118),.WL(WL31));
sram_cell_6t_5 inst_cell_31_119 (.BL(BL119),.BLN(BLN119),.WL(WL31));
sram_cell_6t_5 inst_cell_31_120 (.BL(BL120),.BLN(BLN120),.WL(WL31));
sram_cell_6t_5 inst_cell_31_121 (.BL(BL121),.BLN(BLN121),.WL(WL31));
sram_cell_6t_5 inst_cell_31_122 (.BL(BL122),.BLN(BLN122),.WL(WL31));
sram_cell_6t_5 inst_cell_31_123 (.BL(BL123),.BLN(BLN123),.WL(WL31));
sram_cell_6t_5 inst_cell_31_124 (.BL(BL124),.BLN(BLN124),.WL(WL31));
sram_cell_6t_5 inst_cell_31_125 (.BL(BL125),.BLN(BLN125),.WL(WL31));
sram_cell_6t_5 inst_cell_31_126 (.BL(BL126),.BLN(BLN126),.WL(WL31));
sram_cell_6t_5 inst_cell_31_127 (.BL(BL127),.BLN(BLN127),.WL(WL31));
sram_cell_6t_5 inst_cell_32_0 (.BL(BL0),.BLN(BLN0),.WL(WL32));
sram_cell_6t_5 inst_cell_32_1 (.BL(BL1),.BLN(BLN1),.WL(WL32));
sram_cell_6t_5 inst_cell_32_2 (.BL(BL2),.BLN(BLN2),.WL(WL32));
sram_cell_6t_5 inst_cell_32_3 (.BL(BL3),.BLN(BLN3),.WL(WL32));
sram_cell_6t_5 inst_cell_32_4 (.BL(BL4),.BLN(BLN4),.WL(WL32));
sram_cell_6t_5 inst_cell_32_5 (.BL(BL5),.BLN(BLN5),.WL(WL32));
sram_cell_6t_5 inst_cell_32_6 (.BL(BL6),.BLN(BLN6),.WL(WL32));
sram_cell_6t_5 inst_cell_32_7 (.BL(BL7),.BLN(BLN7),.WL(WL32));
sram_cell_6t_5 inst_cell_32_8 (.BL(BL8),.BLN(BLN8),.WL(WL32));
sram_cell_6t_5 inst_cell_32_9 (.BL(BL9),.BLN(BLN9),.WL(WL32));
sram_cell_6t_5 inst_cell_32_10 (.BL(BL10),.BLN(BLN10),.WL(WL32));
sram_cell_6t_5 inst_cell_32_11 (.BL(BL11),.BLN(BLN11),.WL(WL32));
sram_cell_6t_5 inst_cell_32_12 (.BL(BL12),.BLN(BLN12),.WL(WL32));
sram_cell_6t_5 inst_cell_32_13 (.BL(BL13),.BLN(BLN13),.WL(WL32));
sram_cell_6t_5 inst_cell_32_14 (.BL(BL14),.BLN(BLN14),.WL(WL32));
sram_cell_6t_5 inst_cell_32_15 (.BL(BL15),.BLN(BLN15),.WL(WL32));
sram_cell_6t_5 inst_cell_32_16 (.BL(BL16),.BLN(BLN16),.WL(WL32));
sram_cell_6t_5 inst_cell_32_17 (.BL(BL17),.BLN(BLN17),.WL(WL32));
sram_cell_6t_5 inst_cell_32_18 (.BL(BL18),.BLN(BLN18),.WL(WL32));
sram_cell_6t_5 inst_cell_32_19 (.BL(BL19),.BLN(BLN19),.WL(WL32));
sram_cell_6t_5 inst_cell_32_20 (.BL(BL20),.BLN(BLN20),.WL(WL32));
sram_cell_6t_5 inst_cell_32_21 (.BL(BL21),.BLN(BLN21),.WL(WL32));
sram_cell_6t_5 inst_cell_32_22 (.BL(BL22),.BLN(BLN22),.WL(WL32));
sram_cell_6t_5 inst_cell_32_23 (.BL(BL23),.BLN(BLN23),.WL(WL32));
sram_cell_6t_5 inst_cell_32_24 (.BL(BL24),.BLN(BLN24),.WL(WL32));
sram_cell_6t_5 inst_cell_32_25 (.BL(BL25),.BLN(BLN25),.WL(WL32));
sram_cell_6t_5 inst_cell_32_26 (.BL(BL26),.BLN(BLN26),.WL(WL32));
sram_cell_6t_5 inst_cell_32_27 (.BL(BL27),.BLN(BLN27),.WL(WL32));
sram_cell_6t_5 inst_cell_32_28 (.BL(BL28),.BLN(BLN28),.WL(WL32));
sram_cell_6t_5 inst_cell_32_29 (.BL(BL29),.BLN(BLN29),.WL(WL32));
sram_cell_6t_5 inst_cell_32_30 (.BL(BL30),.BLN(BLN30),.WL(WL32));
sram_cell_6t_5 inst_cell_32_31 (.BL(BL31),.BLN(BLN31),.WL(WL32));
sram_cell_6t_5 inst_cell_32_32 (.BL(BL32),.BLN(BLN32),.WL(WL32));
sram_cell_6t_5 inst_cell_32_33 (.BL(BL33),.BLN(BLN33),.WL(WL32));
sram_cell_6t_5 inst_cell_32_34 (.BL(BL34),.BLN(BLN34),.WL(WL32));
sram_cell_6t_5 inst_cell_32_35 (.BL(BL35),.BLN(BLN35),.WL(WL32));
sram_cell_6t_5 inst_cell_32_36 (.BL(BL36),.BLN(BLN36),.WL(WL32));
sram_cell_6t_5 inst_cell_32_37 (.BL(BL37),.BLN(BLN37),.WL(WL32));
sram_cell_6t_5 inst_cell_32_38 (.BL(BL38),.BLN(BLN38),.WL(WL32));
sram_cell_6t_5 inst_cell_32_39 (.BL(BL39),.BLN(BLN39),.WL(WL32));
sram_cell_6t_5 inst_cell_32_40 (.BL(BL40),.BLN(BLN40),.WL(WL32));
sram_cell_6t_5 inst_cell_32_41 (.BL(BL41),.BLN(BLN41),.WL(WL32));
sram_cell_6t_5 inst_cell_32_42 (.BL(BL42),.BLN(BLN42),.WL(WL32));
sram_cell_6t_5 inst_cell_32_43 (.BL(BL43),.BLN(BLN43),.WL(WL32));
sram_cell_6t_5 inst_cell_32_44 (.BL(BL44),.BLN(BLN44),.WL(WL32));
sram_cell_6t_5 inst_cell_32_45 (.BL(BL45),.BLN(BLN45),.WL(WL32));
sram_cell_6t_5 inst_cell_32_46 (.BL(BL46),.BLN(BLN46),.WL(WL32));
sram_cell_6t_5 inst_cell_32_47 (.BL(BL47),.BLN(BLN47),.WL(WL32));
sram_cell_6t_5 inst_cell_32_48 (.BL(BL48),.BLN(BLN48),.WL(WL32));
sram_cell_6t_5 inst_cell_32_49 (.BL(BL49),.BLN(BLN49),.WL(WL32));
sram_cell_6t_5 inst_cell_32_50 (.BL(BL50),.BLN(BLN50),.WL(WL32));
sram_cell_6t_5 inst_cell_32_51 (.BL(BL51),.BLN(BLN51),.WL(WL32));
sram_cell_6t_5 inst_cell_32_52 (.BL(BL52),.BLN(BLN52),.WL(WL32));
sram_cell_6t_5 inst_cell_32_53 (.BL(BL53),.BLN(BLN53),.WL(WL32));
sram_cell_6t_5 inst_cell_32_54 (.BL(BL54),.BLN(BLN54),.WL(WL32));
sram_cell_6t_5 inst_cell_32_55 (.BL(BL55),.BLN(BLN55),.WL(WL32));
sram_cell_6t_5 inst_cell_32_56 (.BL(BL56),.BLN(BLN56),.WL(WL32));
sram_cell_6t_5 inst_cell_32_57 (.BL(BL57),.BLN(BLN57),.WL(WL32));
sram_cell_6t_5 inst_cell_32_58 (.BL(BL58),.BLN(BLN58),.WL(WL32));
sram_cell_6t_5 inst_cell_32_59 (.BL(BL59),.BLN(BLN59),.WL(WL32));
sram_cell_6t_5 inst_cell_32_60 (.BL(BL60),.BLN(BLN60),.WL(WL32));
sram_cell_6t_5 inst_cell_32_61 (.BL(BL61),.BLN(BLN61),.WL(WL32));
sram_cell_6t_5 inst_cell_32_62 (.BL(BL62),.BLN(BLN62),.WL(WL32));
sram_cell_6t_5 inst_cell_32_63 (.BL(BL63),.BLN(BLN63),.WL(WL32));
sram_cell_6t_5 inst_cell_32_64 (.BL(BL64),.BLN(BLN64),.WL(WL32));
sram_cell_6t_5 inst_cell_32_65 (.BL(BL65),.BLN(BLN65),.WL(WL32));
sram_cell_6t_5 inst_cell_32_66 (.BL(BL66),.BLN(BLN66),.WL(WL32));
sram_cell_6t_5 inst_cell_32_67 (.BL(BL67),.BLN(BLN67),.WL(WL32));
sram_cell_6t_5 inst_cell_32_68 (.BL(BL68),.BLN(BLN68),.WL(WL32));
sram_cell_6t_5 inst_cell_32_69 (.BL(BL69),.BLN(BLN69),.WL(WL32));
sram_cell_6t_5 inst_cell_32_70 (.BL(BL70),.BLN(BLN70),.WL(WL32));
sram_cell_6t_5 inst_cell_32_71 (.BL(BL71),.BLN(BLN71),.WL(WL32));
sram_cell_6t_5 inst_cell_32_72 (.BL(BL72),.BLN(BLN72),.WL(WL32));
sram_cell_6t_5 inst_cell_32_73 (.BL(BL73),.BLN(BLN73),.WL(WL32));
sram_cell_6t_5 inst_cell_32_74 (.BL(BL74),.BLN(BLN74),.WL(WL32));
sram_cell_6t_5 inst_cell_32_75 (.BL(BL75),.BLN(BLN75),.WL(WL32));
sram_cell_6t_5 inst_cell_32_76 (.BL(BL76),.BLN(BLN76),.WL(WL32));
sram_cell_6t_5 inst_cell_32_77 (.BL(BL77),.BLN(BLN77),.WL(WL32));
sram_cell_6t_5 inst_cell_32_78 (.BL(BL78),.BLN(BLN78),.WL(WL32));
sram_cell_6t_5 inst_cell_32_79 (.BL(BL79),.BLN(BLN79),.WL(WL32));
sram_cell_6t_5 inst_cell_32_80 (.BL(BL80),.BLN(BLN80),.WL(WL32));
sram_cell_6t_5 inst_cell_32_81 (.BL(BL81),.BLN(BLN81),.WL(WL32));
sram_cell_6t_5 inst_cell_32_82 (.BL(BL82),.BLN(BLN82),.WL(WL32));
sram_cell_6t_5 inst_cell_32_83 (.BL(BL83),.BLN(BLN83),.WL(WL32));
sram_cell_6t_5 inst_cell_32_84 (.BL(BL84),.BLN(BLN84),.WL(WL32));
sram_cell_6t_5 inst_cell_32_85 (.BL(BL85),.BLN(BLN85),.WL(WL32));
sram_cell_6t_5 inst_cell_32_86 (.BL(BL86),.BLN(BLN86),.WL(WL32));
sram_cell_6t_5 inst_cell_32_87 (.BL(BL87),.BLN(BLN87),.WL(WL32));
sram_cell_6t_5 inst_cell_32_88 (.BL(BL88),.BLN(BLN88),.WL(WL32));
sram_cell_6t_5 inst_cell_32_89 (.BL(BL89),.BLN(BLN89),.WL(WL32));
sram_cell_6t_5 inst_cell_32_90 (.BL(BL90),.BLN(BLN90),.WL(WL32));
sram_cell_6t_5 inst_cell_32_91 (.BL(BL91),.BLN(BLN91),.WL(WL32));
sram_cell_6t_5 inst_cell_32_92 (.BL(BL92),.BLN(BLN92),.WL(WL32));
sram_cell_6t_5 inst_cell_32_93 (.BL(BL93),.BLN(BLN93),.WL(WL32));
sram_cell_6t_5 inst_cell_32_94 (.BL(BL94),.BLN(BLN94),.WL(WL32));
sram_cell_6t_5 inst_cell_32_95 (.BL(BL95),.BLN(BLN95),.WL(WL32));
sram_cell_6t_5 inst_cell_32_96 (.BL(BL96),.BLN(BLN96),.WL(WL32));
sram_cell_6t_5 inst_cell_32_97 (.BL(BL97),.BLN(BLN97),.WL(WL32));
sram_cell_6t_5 inst_cell_32_98 (.BL(BL98),.BLN(BLN98),.WL(WL32));
sram_cell_6t_5 inst_cell_32_99 (.BL(BL99),.BLN(BLN99),.WL(WL32));
sram_cell_6t_5 inst_cell_32_100 (.BL(BL100),.BLN(BLN100),.WL(WL32));
sram_cell_6t_5 inst_cell_32_101 (.BL(BL101),.BLN(BLN101),.WL(WL32));
sram_cell_6t_5 inst_cell_32_102 (.BL(BL102),.BLN(BLN102),.WL(WL32));
sram_cell_6t_5 inst_cell_32_103 (.BL(BL103),.BLN(BLN103),.WL(WL32));
sram_cell_6t_5 inst_cell_32_104 (.BL(BL104),.BLN(BLN104),.WL(WL32));
sram_cell_6t_5 inst_cell_32_105 (.BL(BL105),.BLN(BLN105),.WL(WL32));
sram_cell_6t_5 inst_cell_32_106 (.BL(BL106),.BLN(BLN106),.WL(WL32));
sram_cell_6t_5 inst_cell_32_107 (.BL(BL107),.BLN(BLN107),.WL(WL32));
sram_cell_6t_5 inst_cell_32_108 (.BL(BL108),.BLN(BLN108),.WL(WL32));
sram_cell_6t_5 inst_cell_32_109 (.BL(BL109),.BLN(BLN109),.WL(WL32));
sram_cell_6t_5 inst_cell_32_110 (.BL(BL110),.BLN(BLN110),.WL(WL32));
sram_cell_6t_5 inst_cell_32_111 (.BL(BL111),.BLN(BLN111),.WL(WL32));
sram_cell_6t_5 inst_cell_32_112 (.BL(BL112),.BLN(BLN112),.WL(WL32));
sram_cell_6t_5 inst_cell_32_113 (.BL(BL113),.BLN(BLN113),.WL(WL32));
sram_cell_6t_5 inst_cell_32_114 (.BL(BL114),.BLN(BLN114),.WL(WL32));
sram_cell_6t_5 inst_cell_32_115 (.BL(BL115),.BLN(BLN115),.WL(WL32));
sram_cell_6t_5 inst_cell_32_116 (.BL(BL116),.BLN(BLN116),.WL(WL32));
sram_cell_6t_5 inst_cell_32_117 (.BL(BL117),.BLN(BLN117),.WL(WL32));
sram_cell_6t_5 inst_cell_32_118 (.BL(BL118),.BLN(BLN118),.WL(WL32));
sram_cell_6t_5 inst_cell_32_119 (.BL(BL119),.BLN(BLN119),.WL(WL32));
sram_cell_6t_5 inst_cell_32_120 (.BL(BL120),.BLN(BLN120),.WL(WL32));
sram_cell_6t_5 inst_cell_32_121 (.BL(BL121),.BLN(BLN121),.WL(WL32));
sram_cell_6t_5 inst_cell_32_122 (.BL(BL122),.BLN(BLN122),.WL(WL32));
sram_cell_6t_5 inst_cell_32_123 (.BL(BL123),.BLN(BLN123),.WL(WL32));
sram_cell_6t_5 inst_cell_32_124 (.BL(BL124),.BLN(BLN124),.WL(WL32));
sram_cell_6t_5 inst_cell_32_125 (.BL(BL125),.BLN(BLN125),.WL(WL32));
sram_cell_6t_5 inst_cell_32_126 (.BL(BL126),.BLN(BLN126),.WL(WL32));
sram_cell_6t_5 inst_cell_32_127 (.BL(BL127),.BLN(BLN127),.WL(WL32));
sram_cell_6t_5 inst_cell_33_0 (.BL(BL0),.BLN(BLN0),.WL(WL33));
sram_cell_6t_5 inst_cell_33_1 (.BL(BL1),.BLN(BLN1),.WL(WL33));
sram_cell_6t_5 inst_cell_33_2 (.BL(BL2),.BLN(BLN2),.WL(WL33));
sram_cell_6t_5 inst_cell_33_3 (.BL(BL3),.BLN(BLN3),.WL(WL33));
sram_cell_6t_5 inst_cell_33_4 (.BL(BL4),.BLN(BLN4),.WL(WL33));
sram_cell_6t_5 inst_cell_33_5 (.BL(BL5),.BLN(BLN5),.WL(WL33));
sram_cell_6t_5 inst_cell_33_6 (.BL(BL6),.BLN(BLN6),.WL(WL33));
sram_cell_6t_5 inst_cell_33_7 (.BL(BL7),.BLN(BLN7),.WL(WL33));
sram_cell_6t_5 inst_cell_33_8 (.BL(BL8),.BLN(BLN8),.WL(WL33));
sram_cell_6t_5 inst_cell_33_9 (.BL(BL9),.BLN(BLN9),.WL(WL33));
sram_cell_6t_5 inst_cell_33_10 (.BL(BL10),.BLN(BLN10),.WL(WL33));
sram_cell_6t_5 inst_cell_33_11 (.BL(BL11),.BLN(BLN11),.WL(WL33));
sram_cell_6t_5 inst_cell_33_12 (.BL(BL12),.BLN(BLN12),.WL(WL33));
sram_cell_6t_5 inst_cell_33_13 (.BL(BL13),.BLN(BLN13),.WL(WL33));
sram_cell_6t_5 inst_cell_33_14 (.BL(BL14),.BLN(BLN14),.WL(WL33));
sram_cell_6t_5 inst_cell_33_15 (.BL(BL15),.BLN(BLN15),.WL(WL33));
sram_cell_6t_5 inst_cell_33_16 (.BL(BL16),.BLN(BLN16),.WL(WL33));
sram_cell_6t_5 inst_cell_33_17 (.BL(BL17),.BLN(BLN17),.WL(WL33));
sram_cell_6t_5 inst_cell_33_18 (.BL(BL18),.BLN(BLN18),.WL(WL33));
sram_cell_6t_5 inst_cell_33_19 (.BL(BL19),.BLN(BLN19),.WL(WL33));
sram_cell_6t_5 inst_cell_33_20 (.BL(BL20),.BLN(BLN20),.WL(WL33));
sram_cell_6t_5 inst_cell_33_21 (.BL(BL21),.BLN(BLN21),.WL(WL33));
sram_cell_6t_5 inst_cell_33_22 (.BL(BL22),.BLN(BLN22),.WL(WL33));
sram_cell_6t_5 inst_cell_33_23 (.BL(BL23),.BLN(BLN23),.WL(WL33));
sram_cell_6t_5 inst_cell_33_24 (.BL(BL24),.BLN(BLN24),.WL(WL33));
sram_cell_6t_5 inst_cell_33_25 (.BL(BL25),.BLN(BLN25),.WL(WL33));
sram_cell_6t_5 inst_cell_33_26 (.BL(BL26),.BLN(BLN26),.WL(WL33));
sram_cell_6t_5 inst_cell_33_27 (.BL(BL27),.BLN(BLN27),.WL(WL33));
sram_cell_6t_5 inst_cell_33_28 (.BL(BL28),.BLN(BLN28),.WL(WL33));
sram_cell_6t_5 inst_cell_33_29 (.BL(BL29),.BLN(BLN29),.WL(WL33));
sram_cell_6t_5 inst_cell_33_30 (.BL(BL30),.BLN(BLN30),.WL(WL33));
sram_cell_6t_5 inst_cell_33_31 (.BL(BL31),.BLN(BLN31),.WL(WL33));
sram_cell_6t_5 inst_cell_33_32 (.BL(BL32),.BLN(BLN32),.WL(WL33));
sram_cell_6t_5 inst_cell_33_33 (.BL(BL33),.BLN(BLN33),.WL(WL33));
sram_cell_6t_5 inst_cell_33_34 (.BL(BL34),.BLN(BLN34),.WL(WL33));
sram_cell_6t_5 inst_cell_33_35 (.BL(BL35),.BLN(BLN35),.WL(WL33));
sram_cell_6t_5 inst_cell_33_36 (.BL(BL36),.BLN(BLN36),.WL(WL33));
sram_cell_6t_5 inst_cell_33_37 (.BL(BL37),.BLN(BLN37),.WL(WL33));
sram_cell_6t_5 inst_cell_33_38 (.BL(BL38),.BLN(BLN38),.WL(WL33));
sram_cell_6t_5 inst_cell_33_39 (.BL(BL39),.BLN(BLN39),.WL(WL33));
sram_cell_6t_5 inst_cell_33_40 (.BL(BL40),.BLN(BLN40),.WL(WL33));
sram_cell_6t_5 inst_cell_33_41 (.BL(BL41),.BLN(BLN41),.WL(WL33));
sram_cell_6t_5 inst_cell_33_42 (.BL(BL42),.BLN(BLN42),.WL(WL33));
sram_cell_6t_5 inst_cell_33_43 (.BL(BL43),.BLN(BLN43),.WL(WL33));
sram_cell_6t_5 inst_cell_33_44 (.BL(BL44),.BLN(BLN44),.WL(WL33));
sram_cell_6t_5 inst_cell_33_45 (.BL(BL45),.BLN(BLN45),.WL(WL33));
sram_cell_6t_5 inst_cell_33_46 (.BL(BL46),.BLN(BLN46),.WL(WL33));
sram_cell_6t_5 inst_cell_33_47 (.BL(BL47),.BLN(BLN47),.WL(WL33));
sram_cell_6t_5 inst_cell_33_48 (.BL(BL48),.BLN(BLN48),.WL(WL33));
sram_cell_6t_5 inst_cell_33_49 (.BL(BL49),.BLN(BLN49),.WL(WL33));
sram_cell_6t_5 inst_cell_33_50 (.BL(BL50),.BLN(BLN50),.WL(WL33));
sram_cell_6t_5 inst_cell_33_51 (.BL(BL51),.BLN(BLN51),.WL(WL33));
sram_cell_6t_5 inst_cell_33_52 (.BL(BL52),.BLN(BLN52),.WL(WL33));
sram_cell_6t_5 inst_cell_33_53 (.BL(BL53),.BLN(BLN53),.WL(WL33));
sram_cell_6t_5 inst_cell_33_54 (.BL(BL54),.BLN(BLN54),.WL(WL33));
sram_cell_6t_5 inst_cell_33_55 (.BL(BL55),.BLN(BLN55),.WL(WL33));
sram_cell_6t_5 inst_cell_33_56 (.BL(BL56),.BLN(BLN56),.WL(WL33));
sram_cell_6t_5 inst_cell_33_57 (.BL(BL57),.BLN(BLN57),.WL(WL33));
sram_cell_6t_5 inst_cell_33_58 (.BL(BL58),.BLN(BLN58),.WL(WL33));
sram_cell_6t_5 inst_cell_33_59 (.BL(BL59),.BLN(BLN59),.WL(WL33));
sram_cell_6t_5 inst_cell_33_60 (.BL(BL60),.BLN(BLN60),.WL(WL33));
sram_cell_6t_5 inst_cell_33_61 (.BL(BL61),.BLN(BLN61),.WL(WL33));
sram_cell_6t_5 inst_cell_33_62 (.BL(BL62),.BLN(BLN62),.WL(WL33));
sram_cell_6t_5 inst_cell_33_63 (.BL(BL63),.BLN(BLN63),.WL(WL33));
sram_cell_6t_5 inst_cell_33_64 (.BL(BL64),.BLN(BLN64),.WL(WL33));
sram_cell_6t_5 inst_cell_33_65 (.BL(BL65),.BLN(BLN65),.WL(WL33));
sram_cell_6t_5 inst_cell_33_66 (.BL(BL66),.BLN(BLN66),.WL(WL33));
sram_cell_6t_5 inst_cell_33_67 (.BL(BL67),.BLN(BLN67),.WL(WL33));
sram_cell_6t_5 inst_cell_33_68 (.BL(BL68),.BLN(BLN68),.WL(WL33));
sram_cell_6t_5 inst_cell_33_69 (.BL(BL69),.BLN(BLN69),.WL(WL33));
sram_cell_6t_5 inst_cell_33_70 (.BL(BL70),.BLN(BLN70),.WL(WL33));
sram_cell_6t_5 inst_cell_33_71 (.BL(BL71),.BLN(BLN71),.WL(WL33));
sram_cell_6t_5 inst_cell_33_72 (.BL(BL72),.BLN(BLN72),.WL(WL33));
sram_cell_6t_5 inst_cell_33_73 (.BL(BL73),.BLN(BLN73),.WL(WL33));
sram_cell_6t_5 inst_cell_33_74 (.BL(BL74),.BLN(BLN74),.WL(WL33));
sram_cell_6t_5 inst_cell_33_75 (.BL(BL75),.BLN(BLN75),.WL(WL33));
sram_cell_6t_5 inst_cell_33_76 (.BL(BL76),.BLN(BLN76),.WL(WL33));
sram_cell_6t_5 inst_cell_33_77 (.BL(BL77),.BLN(BLN77),.WL(WL33));
sram_cell_6t_5 inst_cell_33_78 (.BL(BL78),.BLN(BLN78),.WL(WL33));
sram_cell_6t_5 inst_cell_33_79 (.BL(BL79),.BLN(BLN79),.WL(WL33));
sram_cell_6t_5 inst_cell_33_80 (.BL(BL80),.BLN(BLN80),.WL(WL33));
sram_cell_6t_5 inst_cell_33_81 (.BL(BL81),.BLN(BLN81),.WL(WL33));
sram_cell_6t_5 inst_cell_33_82 (.BL(BL82),.BLN(BLN82),.WL(WL33));
sram_cell_6t_5 inst_cell_33_83 (.BL(BL83),.BLN(BLN83),.WL(WL33));
sram_cell_6t_5 inst_cell_33_84 (.BL(BL84),.BLN(BLN84),.WL(WL33));
sram_cell_6t_5 inst_cell_33_85 (.BL(BL85),.BLN(BLN85),.WL(WL33));
sram_cell_6t_5 inst_cell_33_86 (.BL(BL86),.BLN(BLN86),.WL(WL33));
sram_cell_6t_5 inst_cell_33_87 (.BL(BL87),.BLN(BLN87),.WL(WL33));
sram_cell_6t_5 inst_cell_33_88 (.BL(BL88),.BLN(BLN88),.WL(WL33));
sram_cell_6t_5 inst_cell_33_89 (.BL(BL89),.BLN(BLN89),.WL(WL33));
sram_cell_6t_5 inst_cell_33_90 (.BL(BL90),.BLN(BLN90),.WL(WL33));
sram_cell_6t_5 inst_cell_33_91 (.BL(BL91),.BLN(BLN91),.WL(WL33));
sram_cell_6t_5 inst_cell_33_92 (.BL(BL92),.BLN(BLN92),.WL(WL33));
sram_cell_6t_5 inst_cell_33_93 (.BL(BL93),.BLN(BLN93),.WL(WL33));
sram_cell_6t_5 inst_cell_33_94 (.BL(BL94),.BLN(BLN94),.WL(WL33));
sram_cell_6t_5 inst_cell_33_95 (.BL(BL95),.BLN(BLN95),.WL(WL33));
sram_cell_6t_5 inst_cell_33_96 (.BL(BL96),.BLN(BLN96),.WL(WL33));
sram_cell_6t_5 inst_cell_33_97 (.BL(BL97),.BLN(BLN97),.WL(WL33));
sram_cell_6t_5 inst_cell_33_98 (.BL(BL98),.BLN(BLN98),.WL(WL33));
sram_cell_6t_5 inst_cell_33_99 (.BL(BL99),.BLN(BLN99),.WL(WL33));
sram_cell_6t_5 inst_cell_33_100 (.BL(BL100),.BLN(BLN100),.WL(WL33));
sram_cell_6t_5 inst_cell_33_101 (.BL(BL101),.BLN(BLN101),.WL(WL33));
sram_cell_6t_5 inst_cell_33_102 (.BL(BL102),.BLN(BLN102),.WL(WL33));
sram_cell_6t_5 inst_cell_33_103 (.BL(BL103),.BLN(BLN103),.WL(WL33));
sram_cell_6t_5 inst_cell_33_104 (.BL(BL104),.BLN(BLN104),.WL(WL33));
sram_cell_6t_5 inst_cell_33_105 (.BL(BL105),.BLN(BLN105),.WL(WL33));
sram_cell_6t_5 inst_cell_33_106 (.BL(BL106),.BLN(BLN106),.WL(WL33));
sram_cell_6t_5 inst_cell_33_107 (.BL(BL107),.BLN(BLN107),.WL(WL33));
sram_cell_6t_5 inst_cell_33_108 (.BL(BL108),.BLN(BLN108),.WL(WL33));
sram_cell_6t_5 inst_cell_33_109 (.BL(BL109),.BLN(BLN109),.WL(WL33));
sram_cell_6t_5 inst_cell_33_110 (.BL(BL110),.BLN(BLN110),.WL(WL33));
sram_cell_6t_5 inst_cell_33_111 (.BL(BL111),.BLN(BLN111),.WL(WL33));
sram_cell_6t_5 inst_cell_33_112 (.BL(BL112),.BLN(BLN112),.WL(WL33));
sram_cell_6t_5 inst_cell_33_113 (.BL(BL113),.BLN(BLN113),.WL(WL33));
sram_cell_6t_5 inst_cell_33_114 (.BL(BL114),.BLN(BLN114),.WL(WL33));
sram_cell_6t_5 inst_cell_33_115 (.BL(BL115),.BLN(BLN115),.WL(WL33));
sram_cell_6t_5 inst_cell_33_116 (.BL(BL116),.BLN(BLN116),.WL(WL33));
sram_cell_6t_5 inst_cell_33_117 (.BL(BL117),.BLN(BLN117),.WL(WL33));
sram_cell_6t_5 inst_cell_33_118 (.BL(BL118),.BLN(BLN118),.WL(WL33));
sram_cell_6t_5 inst_cell_33_119 (.BL(BL119),.BLN(BLN119),.WL(WL33));
sram_cell_6t_5 inst_cell_33_120 (.BL(BL120),.BLN(BLN120),.WL(WL33));
sram_cell_6t_5 inst_cell_33_121 (.BL(BL121),.BLN(BLN121),.WL(WL33));
sram_cell_6t_5 inst_cell_33_122 (.BL(BL122),.BLN(BLN122),.WL(WL33));
sram_cell_6t_5 inst_cell_33_123 (.BL(BL123),.BLN(BLN123),.WL(WL33));
sram_cell_6t_5 inst_cell_33_124 (.BL(BL124),.BLN(BLN124),.WL(WL33));
sram_cell_6t_5 inst_cell_33_125 (.BL(BL125),.BLN(BLN125),.WL(WL33));
sram_cell_6t_5 inst_cell_33_126 (.BL(BL126),.BLN(BLN126),.WL(WL33));
sram_cell_6t_5 inst_cell_33_127 (.BL(BL127),.BLN(BLN127),.WL(WL33));
sram_cell_6t_5 inst_cell_34_0 (.BL(BL0),.BLN(BLN0),.WL(WL34));
sram_cell_6t_5 inst_cell_34_1 (.BL(BL1),.BLN(BLN1),.WL(WL34));
sram_cell_6t_5 inst_cell_34_2 (.BL(BL2),.BLN(BLN2),.WL(WL34));
sram_cell_6t_5 inst_cell_34_3 (.BL(BL3),.BLN(BLN3),.WL(WL34));
sram_cell_6t_5 inst_cell_34_4 (.BL(BL4),.BLN(BLN4),.WL(WL34));
sram_cell_6t_5 inst_cell_34_5 (.BL(BL5),.BLN(BLN5),.WL(WL34));
sram_cell_6t_5 inst_cell_34_6 (.BL(BL6),.BLN(BLN6),.WL(WL34));
sram_cell_6t_5 inst_cell_34_7 (.BL(BL7),.BLN(BLN7),.WL(WL34));
sram_cell_6t_5 inst_cell_34_8 (.BL(BL8),.BLN(BLN8),.WL(WL34));
sram_cell_6t_5 inst_cell_34_9 (.BL(BL9),.BLN(BLN9),.WL(WL34));
sram_cell_6t_5 inst_cell_34_10 (.BL(BL10),.BLN(BLN10),.WL(WL34));
sram_cell_6t_5 inst_cell_34_11 (.BL(BL11),.BLN(BLN11),.WL(WL34));
sram_cell_6t_5 inst_cell_34_12 (.BL(BL12),.BLN(BLN12),.WL(WL34));
sram_cell_6t_5 inst_cell_34_13 (.BL(BL13),.BLN(BLN13),.WL(WL34));
sram_cell_6t_5 inst_cell_34_14 (.BL(BL14),.BLN(BLN14),.WL(WL34));
sram_cell_6t_5 inst_cell_34_15 (.BL(BL15),.BLN(BLN15),.WL(WL34));
sram_cell_6t_5 inst_cell_34_16 (.BL(BL16),.BLN(BLN16),.WL(WL34));
sram_cell_6t_5 inst_cell_34_17 (.BL(BL17),.BLN(BLN17),.WL(WL34));
sram_cell_6t_5 inst_cell_34_18 (.BL(BL18),.BLN(BLN18),.WL(WL34));
sram_cell_6t_5 inst_cell_34_19 (.BL(BL19),.BLN(BLN19),.WL(WL34));
sram_cell_6t_5 inst_cell_34_20 (.BL(BL20),.BLN(BLN20),.WL(WL34));
sram_cell_6t_5 inst_cell_34_21 (.BL(BL21),.BLN(BLN21),.WL(WL34));
sram_cell_6t_5 inst_cell_34_22 (.BL(BL22),.BLN(BLN22),.WL(WL34));
sram_cell_6t_5 inst_cell_34_23 (.BL(BL23),.BLN(BLN23),.WL(WL34));
sram_cell_6t_5 inst_cell_34_24 (.BL(BL24),.BLN(BLN24),.WL(WL34));
sram_cell_6t_5 inst_cell_34_25 (.BL(BL25),.BLN(BLN25),.WL(WL34));
sram_cell_6t_5 inst_cell_34_26 (.BL(BL26),.BLN(BLN26),.WL(WL34));
sram_cell_6t_5 inst_cell_34_27 (.BL(BL27),.BLN(BLN27),.WL(WL34));
sram_cell_6t_5 inst_cell_34_28 (.BL(BL28),.BLN(BLN28),.WL(WL34));
sram_cell_6t_5 inst_cell_34_29 (.BL(BL29),.BLN(BLN29),.WL(WL34));
sram_cell_6t_5 inst_cell_34_30 (.BL(BL30),.BLN(BLN30),.WL(WL34));
sram_cell_6t_5 inst_cell_34_31 (.BL(BL31),.BLN(BLN31),.WL(WL34));
sram_cell_6t_5 inst_cell_34_32 (.BL(BL32),.BLN(BLN32),.WL(WL34));
sram_cell_6t_5 inst_cell_34_33 (.BL(BL33),.BLN(BLN33),.WL(WL34));
sram_cell_6t_5 inst_cell_34_34 (.BL(BL34),.BLN(BLN34),.WL(WL34));
sram_cell_6t_5 inst_cell_34_35 (.BL(BL35),.BLN(BLN35),.WL(WL34));
sram_cell_6t_5 inst_cell_34_36 (.BL(BL36),.BLN(BLN36),.WL(WL34));
sram_cell_6t_5 inst_cell_34_37 (.BL(BL37),.BLN(BLN37),.WL(WL34));
sram_cell_6t_5 inst_cell_34_38 (.BL(BL38),.BLN(BLN38),.WL(WL34));
sram_cell_6t_5 inst_cell_34_39 (.BL(BL39),.BLN(BLN39),.WL(WL34));
sram_cell_6t_5 inst_cell_34_40 (.BL(BL40),.BLN(BLN40),.WL(WL34));
sram_cell_6t_5 inst_cell_34_41 (.BL(BL41),.BLN(BLN41),.WL(WL34));
sram_cell_6t_5 inst_cell_34_42 (.BL(BL42),.BLN(BLN42),.WL(WL34));
sram_cell_6t_5 inst_cell_34_43 (.BL(BL43),.BLN(BLN43),.WL(WL34));
sram_cell_6t_5 inst_cell_34_44 (.BL(BL44),.BLN(BLN44),.WL(WL34));
sram_cell_6t_5 inst_cell_34_45 (.BL(BL45),.BLN(BLN45),.WL(WL34));
sram_cell_6t_5 inst_cell_34_46 (.BL(BL46),.BLN(BLN46),.WL(WL34));
sram_cell_6t_5 inst_cell_34_47 (.BL(BL47),.BLN(BLN47),.WL(WL34));
sram_cell_6t_5 inst_cell_34_48 (.BL(BL48),.BLN(BLN48),.WL(WL34));
sram_cell_6t_5 inst_cell_34_49 (.BL(BL49),.BLN(BLN49),.WL(WL34));
sram_cell_6t_5 inst_cell_34_50 (.BL(BL50),.BLN(BLN50),.WL(WL34));
sram_cell_6t_5 inst_cell_34_51 (.BL(BL51),.BLN(BLN51),.WL(WL34));
sram_cell_6t_5 inst_cell_34_52 (.BL(BL52),.BLN(BLN52),.WL(WL34));
sram_cell_6t_5 inst_cell_34_53 (.BL(BL53),.BLN(BLN53),.WL(WL34));
sram_cell_6t_5 inst_cell_34_54 (.BL(BL54),.BLN(BLN54),.WL(WL34));
sram_cell_6t_5 inst_cell_34_55 (.BL(BL55),.BLN(BLN55),.WL(WL34));
sram_cell_6t_5 inst_cell_34_56 (.BL(BL56),.BLN(BLN56),.WL(WL34));
sram_cell_6t_5 inst_cell_34_57 (.BL(BL57),.BLN(BLN57),.WL(WL34));
sram_cell_6t_5 inst_cell_34_58 (.BL(BL58),.BLN(BLN58),.WL(WL34));
sram_cell_6t_5 inst_cell_34_59 (.BL(BL59),.BLN(BLN59),.WL(WL34));
sram_cell_6t_5 inst_cell_34_60 (.BL(BL60),.BLN(BLN60),.WL(WL34));
sram_cell_6t_5 inst_cell_34_61 (.BL(BL61),.BLN(BLN61),.WL(WL34));
sram_cell_6t_5 inst_cell_34_62 (.BL(BL62),.BLN(BLN62),.WL(WL34));
sram_cell_6t_5 inst_cell_34_63 (.BL(BL63),.BLN(BLN63),.WL(WL34));
sram_cell_6t_5 inst_cell_34_64 (.BL(BL64),.BLN(BLN64),.WL(WL34));
sram_cell_6t_5 inst_cell_34_65 (.BL(BL65),.BLN(BLN65),.WL(WL34));
sram_cell_6t_5 inst_cell_34_66 (.BL(BL66),.BLN(BLN66),.WL(WL34));
sram_cell_6t_5 inst_cell_34_67 (.BL(BL67),.BLN(BLN67),.WL(WL34));
sram_cell_6t_5 inst_cell_34_68 (.BL(BL68),.BLN(BLN68),.WL(WL34));
sram_cell_6t_5 inst_cell_34_69 (.BL(BL69),.BLN(BLN69),.WL(WL34));
sram_cell_6t_5 inst_cell_34_70 (.BL(BL70),.BLN(BLN70),.WL(WL34));
sram_cell_6t_5 inst_cell_34_71 (.BL(BL71),.BLN(BLN71),.WL(WL34));
sram_cell_6t_5 inst_cell_34_72 (.BL(BL72),.BLN(BLN72),.WL(WL34));
sram_cell_6t_5 inst_cell_34_73 (.BL(BL73),.BLN(BLN73),.WL(WL34));
sram_cell_6t_5 inst_cell_34_74 (.BL(BL74),.BLN(BLN74),.WL(WL34));
sram_cell_6t_5 inst_cell_34_75 (.BL(BL75),.BLN(BLN75),.WL(WL34));
sram_cell_6t_5 inst_cell_34_76 (.BL(BL76),.BLN(BLN76),.WL(WL34));
sram_cell_6t_5 inst_cell_34_77 (.BL(BL77),.BLN(BLN77),.WL(WL34));
sram_cell_6t_5 inst_cell_34_78 (.BL(BL78),.BLN(BLN78),.WL(WL34));
sram_cell_6t_5 inst_cell_34_79 (.BL(BL79),.BLN(BLN79),.WL(WL34));
sram_cell_6t_5 inst_cell_34_80 (.BL(BL80),.BLN(BLN80),.WL(WL34));
sram_cell_6t_5 inst_cell_34_81 (.BL(BL81),.BLN(BLN81),.WL(WL34));
sram_cell_6t_5 inst_cell_34_82 (.BL(BL82),.BLN(BLN82),.WL(WL34));
sram_cell_6t_5 inst_cell_34_83 (.BL(BL83),.BLN(BLN83),.WL(WL34));
sram_cell_6t_5 inst_cell_34_84 (.BL(BL84),.BLN(BLN84),.WL(WL34));
sram_cell_6t_5 inst_cell_34_85 (.BL(BL85),.BLN(BLN85),.WL(WL34));
sram_cell_6t_5 inst_cell_34_86 (.BL(BL86),.BLN(BLN86),.WL(WL34));
sram_cell_6t_5 inst_cell_34_87 (.BL(BL87),.BLN(BLN87),.WL(WL34));
sram_cell_6t_5 inst_cell_34_88 (.BL(BL88),.BLN(BLN88),.WL(WL34));
sram_cell_6t_5 inst_cell_34_89 (.BL(BL89),.BLN(BLN89),.WL(WL34));
sram_cell_6t_5 inst_cell_34_90 (.BL(BL90),.BLN(BLN90),.WL(WL34));
sram_cell_6t_5 inst_cell_34_91 (.BL(BL91),.BLN(BLN91),.WL(WL34));
sram_cell_6t_5 inst_cell_34_92 (.BL(BL92),.BLN(BLN92),.WL(WL34));
sram_cell_6t_5 inst_cell_34_93 (.BL(BL93),.BLN(BLN93),.WL(WL34));
sram_cell_6t_5 inst_cell_34_94 (.BL(BL94),.BLN(BLN94),.WL(WL34));
sram_cell_6t_5 inst_cell_34_95 (.BL(BL95),.BLN(BLN95),.WL(WL34));
sram_cell_6t_5 inst_cell_34_96 (.BL(BL96),.BLN(BLN96),.WL(WL34));
sram_cell_6t_5 inst_cell_34_97 (.BL(BL97),.BLN(BLN97),.WL(WL34));
sram_cell_6t_5 inst_cell_34_98 (.BL(BL98),.BLN(BLN98),.WL(WL34));
sram_cell_6t_5 inst_cell_34_99 (.BL(BL99),.BLN(BLN99),.WL(WL34));
sram_cell_6t_5 inst_cell_34_100 (.BL(BL100),.BLN(BLN100),.WL(WL34));
sram_cell_6t_5 inst_cell_34_101 (.BL(BL101),.BLN(BLN101),.WL(WL34));
sram_cell_6t_5 inst_cell_34_102 (.BL(BL102),.BLN(BLN102),.WL(WL34));
sram_cell_6t_5 inst_cell_34_103 (.BL(BL103),.BLN(BLN103),.WL(WL34));
sram_cell_6t_5 inst_cell_34_104 (.BL(BL104),.BLN(BLN104),.WL(WL34));
sram_cell_6t_5 inst_cell_34_105 (.BL(BL105),.BLN(BLN105),.WL(WL34));
sram_cell_6t_5 inst_cell_34_106 (.BL(BL106),.BLN(BLN106),.WL(WL34));
sram_cell_6t_5 inst_cell_34_107 (.BL(BL107),.BLN(BLN107),.WL(WL34));
sram_cell_6t_5 inst_cell_34_108 (.BL(BL108),.BLN(BLN108),.WL(WL34));
sram_cell_6t_5 inst_cell_34_109 (.BL(BL109),.BLN(BLN109),.WL(WL34));
sram_cell_6t_5 inst_cell_34_110 (.BL(BL110),.BLN(BLN110),.WL(WL34));
sram_cell_6t_5 inst_cell_34_111 (.BL(BL111),.BLN(BLN111),.WL(WL34));
sram_cell_6t_5 inst_cell_34_112 (.BL(BL112),.BLN(BLN112),.WL(WL34));
sram_cell_6t_5 inst_cell_34_113 (.BL(BL113),.BLN(BLN113),.WL(WL34));
sram_cell_6t_5 inst_cell_34_114 (.BL(BL114),.BLN(BLN114),.WL(WL34));
sram_cell_6t_5 inst_cell_34_115 (.BL(BL115),.BLN(BLN115),.WL(WL34));
sram_cell_6t_5 inst_cell_34_116 (.BL(BL116),.BLN(BLN116),.WL(WL34));
sram_cell_6t_5 inst_cell_34_117 (.BL(BL117),.BLN(BLN117),.WL(WL34));
sram_cell_6t_5 inst_cell_34_118 (.BL(BL118),.BLN(BLN118),.WL(WL34));
sram_cell_6t_5 inst_cell_34_119 (.BL(BL119),.BLN(BLN119),.WL(WL34));
sram_cell_6t_5 inst_cell_34_120 (.BL(BL120),.BLN(BLN120),.WL(WL34));
sram_cell_6t_5 inst_cell_34_121 (.BL(BL121),.BLN(BLN121),.WL(WL34));
sram_cell_6t_5 inst_cell_34_122 (.BL(BL122),.BLN(BLN122),.WL(WL34));
sram_cell_6t_5 inst_cell_34_123 (.BL(BL123),.BLN(BLN123),.WL(WL34));
sram_cell_6t_5 inst_cell_34_124 (.BL(BL124),.BLN(BLN124),.WL(WL34));
sram_cell_6t_5 inst_cell_34_125 (.BL(BL125),.BLN(BLN125),.WL(WL34));
sram_cell_6t_5 inst_cell_34_126 (.BL(BL126),.BLN(BLN126),.WL(WL34));
sram_cell_6t_5 inst_cell_34_127 (.BL(BL127),.BLN(BLN127),.WL(WL34));
sram_cell_6t_5 inst_cell_35_0 (.BL(BL0),.BLN(BLN0),.WL(WL35));
sram_cell_6t_5 inst_cell_35_1 (.BL(BL1),.BLN(BLN1),.WL(WL35));
sram_cell_6t_5 inst_cell_35_2 (.BL(BL2),.BLN(BLN2),.WL(WL35));
sram_cell_6t_5 inst_cell_35_3 (.BL(BL3),.BLN(BLN3),.WL(WL35));
sram_cell_6t_5 inst_cell_35_4 (.BL(BL4),.BLN(BLN4),.WL(WL35));
sram_cell_6t_5 inst_cell_35_5 (.BL(BL5),.BLN(BLN5),.WL(WL35));
sram_cell_6t_5 inst_cell_35_6 (.BL(BL6),.BLN(BLN6),.WL(WL35));
sram_cell_6t_5 inst_cell_35_7 (.BL(BL7),.BLN(BLN7),.WL(WL35));
sram_cell_6t_5 inst_cell_35_8 (.BL(BL8),.BLN(BLN8),.WL(WL35));
sram_cell_6t_5 inst_cell_35_9 (.BL(BL9),.BLN(BLN9),.WL(WL35));
sram_cell_6t_5 inst_cell_35_10 (.BL(BL10),.BLN(BLN10),.WL(WL35));
sram_cell_6t_5 inst_cell_35_11 (.BL(BL11),.BLN(BLN11),.WL(WL35));
sram_cell_6t_5 inst_cell_35_12 (.BL(BL12),.BLN(BLN12),.WL(WL35));
sram_cell_6t_5 inst_cell_35_13 (.BL(BL13),.BLN(BLN13),.WL(WL35));
sram_cell_6t_5 inst_cell_35_14 (.BL(BL14),.BLN(BLN14),.WL(WL35));
sram_cell_6t_5 inst_cell_35_15 (.BL(BL15),.BLN(BLN15),.WL(WL35));
sram_cell_6t_5 inst_cell_35_16 (.BL(BL16),.BLN(BLN16),.WL(WL35));
sram_cell_6t_5 inst_cell_35_17 (.BL(BL17),.BLN(BLN17),.WL(WL35));
sram_cell_6t_5 inst_cell_35_18 (.BL(BL18),.BLN(BLN18),.WL(WL35));
sram_cell_6t_5 inst_cell_35_19 (.BL(BL19),.BLN(BLN19),.WL(WL35));
sram_cell_6t_5 inst_cell_35_20 (.BL(BL20),.BLN(BLN20),.WL(WL35));
sram_cell_6t_5 inst_cell_35_21 (.BL(BL21),.BLN(BLN21),.WL(WL35));
sram_cell_6t_5 inst_cell_35_22 (.BL(BL22),.BLN(BLN22),.WL(WL35));
sram_cell_6t_5 inst_cell_35_23 (.BL(BL23),.BLN(BLN23),.WL(WL35));
sram_cell_6t_5 inst_cell_35_24 (.BL(BL24),.BLN(BLN24),.WL(WL35));
sram_cell_6t_5 inst_cell_35_25 (.BL(BL25),.BLN(BLN25),.WL(WL35));
sram_cell_6t_5 inst_cell_35_26 (.BL(BL26),.BLN(BLN26),.WL(WL35));
sram_cell_6t_5 inst_cell_35_27 (.BL(BL27),.BLN(BLN27),.WL(WL35));
sram_cell_6t_5 inst_cell_35_28 (.BL(BL28),.BLN(BLN28),.WL(WL35));
sram_cell_6t_5 inst_cell_35_29 (.BL(BL29),.BLN(BLN29),.WL(WL35));
sram_cell_6t_5 inst_cell_35_30 (.BL(BL30),.BLN(BLN30),.WL(WL35));
sram_cell_6t_5 inst_cell_35_31 (.BL(BL31),.BLN(BLN31),.WL(WL35));
sram_cell_6t_5 inst_cell_35_32 (.BL(BL32),.BLN(BLN32),.WL(WL35));
sram_cell_6t_5 inst_cell_35_33 (.BL(BL33),.BLN(BLN33),.WL(WL35));
sram_cell_6t_5 inst_cell_35_34 (.BL(BL34),.BLN(BLN34),.WL(WL35));
sram_cell_6t_5 inst_cell_35_35 (.BL(BL35),.BLN(BLN35),.WL(WL35));
sram_cell_6t_5 inst_cell_35_36 (.BL(BL36),.BLN(BLN36),.WL(WL35));
sram_cell_6t_5 inst_cell_35_37 (.BL(BL37),.BLN(BLN37),.WL(WL35));
sram_cell_6t_5 inst_cell_35_38 (.BL(BL38),.BLN(BLN38),.WL(WL35));
sram_cell_6t_5 inst_cell_35_39 (.BL(BL39),.BLN(BLN39),.WL(WL35));
sram_cell_6t_5 inst_cell_35_40 (.BL(BL40),.BLN(BLN40),.WL(WL35));
sram_cell_6t_5 inst_cell_35_41 (.BL(BL41),.BLN(BLN41),.WL(WL35));
sram_cell_6t_5 inst_cell_35_42 (.BL(BL42),.BLN(BLN42),.WL(WL35));
sram_cell_6t_5 inst_cell_35_43 (.BL(BL43),.BLN(BLN43),.WL(WL35));
sram_cell_6t_5 inst_cell_35_44 (.BL(BL44),.BLN(BLN44),.WL(WL35));
sram_cell_6t_5 inst_cell_35_45 (.BL(BL45),.BLN(BLN45),.WL(WL35));
sram_cell_6t_5 inst_cell_35_46 (.BL(BL46),.BLN(BLN46),.WL(WL35));
sram_cell_6t_5 inst_cell_35_47 (.BL(BL47),.BLN(BLN47),.WL(WL35));
sram_cell_6t_5 inst_cell_35_48 (.BL(BL48),.BLN(BLN48),.WL(WL35));
sram_cell_6t_5 inst_cell_35_49 (.BL(BL49),.BLN(BLN49),.WL(WL35));
sram_cell_6t_5 inst_cell_35_50 (.BL(BL50),.BLN(BLN50),.WL(WL35));
sram_cell_6t_5 inst_cell_35_51 (.BL(BL51),.BLN(BLN51),.WL(WL35));
sram_cell_6t_5 inst_cell_35_52 (.BL(BL52),.BLN(BLN52),.WL(WL35));
sram_cell_6t_5 inst_cell_35_53 (.BL(BL53),.BLN(BLN53),.WL(WL35));
sram_cell_6t_5 inst_cell_35_54 (.BL(BL54),.BLN(BLN54),.WL(WL35));
sram_cell_6t_5 inst_cell_35_55 (.BL(BL55),.BLN(BLN55),.WL(WL35));
sram_cell_6t_5 inst_cell_35_56 (.BL(BL56),.BLN(BLN56),.WL(WL35));
sram_cell_6t_5 inst_cell_35_57 (.BL(BL57),.BLN(BLN57),.WL(WL35));
sram_cell_6t_5 inst_cell_35_58 (.BL(BL58),.BLN(BLN58),.WL(WL35));
sram_cell_6t_5 inst_cell_35_59 (.BL(BL59),.BLN(BLN59),.WL(WL35));
sram_cell_6t_5 inst_cell_35_60 (.BL(BL60),.BLN(BLN60),.WL(WL35));
sram_cell_6t_5 inst_cell_35_61 (.BL(BL61),.BLN(BLN61),.WL(WL35));
sram_cell_6t_5 inst_cell_35_62 (.BL(BL62),.BLN(BLN62),.WL(WL35));
sram_cell_6t_5 inst_cell_35_63 (.BL(BL63),.BLN(BLN63),.WL(WL35));
sram_cell_6t_5 inst_cell_35_64 (.BL(BL64),.BLN(BLN64),.WL(WL35));
sram_cell_6t_5 inst_cell_35_65 (.BL(BL65),.BLN(BLN65),.WL(WL35));
sram_cell_6t_5 inst_cell_35_66 (.BL(BL66),.BLN(BLN66),.WL(WL35));
sram_cell_6t_5 inst_cell_35_67 (.BL(BL67),.BLN(BLN67),.WL(WL35));
sram_cell_6t_5 inst_cell_35_68 (.BL(BL68),.BLN(BLN68),.WL(WL35));
sram_cell_6t_5 inst_cell_35_69 (.BL(BL69),.BLN(BLN69),.WL(WL35));
sram_cell_6t_5 inst_cell_35_70 (.BL(BL70),.BLN(BLN70),.WL(WL35));
sram_cell_6t_5 inst_cell_35_71 (.BL(BL71),.BLN(BLN71),.WL(WL35));
sram_cell_6t_5 inst_cell_35_72 (.BL(BL72),.BLN(BLN72),.WL(WL35));
sram_cell_6t_5 inst_cell_35_73 (.BL(BL73),.BLN(BLN73),.WL(WL35));
sram_cell_6t_5 inst_cell_35_74 (.BL(BL74),.BLN(BLN74),.WL(WL35));
sram_cell_6t_5 inst_cell_35_75 (.BL(BL75),.BLN(BLN75),.WL(WL35));
sram_cell_6t_5 inst_cell_35_76 (.BL(BL76),.BLN(BLN76),.WL(WL35));
sram_cell_6t_5 inst_cell_35_77 (.BL(BL77),.BLN(BLN77),.WL(WL35));
sram_cell_6t_5 inst_cell_35_78 (.BL(BL78),.BLN(BLN78),.WL(WL35));
sram_cell_6t_5 inst_cell_35_79 (.BL(BL79),.BLN(BLN79),.WL(WL35));
sram_cell_6t_5 inst_cell_35_80 (.BL(BL80),.BLN(BLN80),.WL(WL35));
sram_cell_6t_5 inst_cell_35_81 (.BL(BL81),.BLN(BLN81),.WL(WL35));
sram_cell_6t_5 inst_cell_35_82 (.BL(BL82),.BLN(BLN82),.WL(WL35));
sram_cell_6t_5 inst_cell_35_83 (.BL(BL83),.BLN(BLN83),.WL(WL35));
sram_cell_6t_5 inst_cell_35_84 (.BL(BL84),.BLN(BLN84),.WL(WL35));
sram_cell_6t_5 inst_cell_35_85 (.BL(BL85),.BLN(BLN85),.WL(WL35));
sram_cell_6t_5 inst_cell_35_86 (.BL(BL86),.BLN(BLN86),.WL(WL35));
sram_cell_6t_5 inst_cell_35_87 (.BL(BL87),.BLN(BLN87),.WL(WL35));
sram_cell_6t_5 inst_cell_35_88 (.BL(BL88),.BLN(BLN88),.WL(WL35));
sram_cell_6t_5 inst_cell_35_89 (.BL(BL89),.BLN(BLN89),.WL(WL35));
sram_cell_6t_5 inst_cell_35_90 (.BL(BL90),.BLN(BLN90),.WL(WL35));
sram_cell_6t_5 inst_cell_35_91 (.BL(BL91),.BLN(BLN91),.WL(WL35));
sram_cell_6t_5 inst_cell_35_92 (.BL(BL92),.BLN(BLN92),.WL(WL35));
sram_cell_6t_5 inst_cell_35_93 (.BL(BL93),.BLN(BLN93),.WL(WL35));
sram_cell_6t_5 inst_cell_35_94 (.BL(BL94),.BLN(BLN94),.WL(WL35));
sram_cell_6t_5 inst_cell_35_95 (.BL(BL95),.BLN(BLN95),.WL(WL35));
sram_cell_6t_5 inst_cell_35_96 (.BL(BL96),.BLN(BLN96),.WL(WL35));
sram_cell_6t_5 inst_cell_35_97 (.BL(BL97),.BLN(BLN97),.WL(WL35));
sram_cell_6t_5 inst_cell_35_98 (.BL(BL98),.BLN(BLN98),.WL(WL35));
sram_cell_6t_5 inst_cell_35_99 (.BL(BL99),.BLN(BLN99),.WL(WL35));
sram_cell_6t_5 inst_cell_35_100 (.BL(BL100),.BLN(BLN100),.WL(WL35));
sram_cell_6t_5 inst_cell_35_101 (.BL(BL101),.BLN(BLN101),.WL(WL35));
sram_cell_6t_5 inst_cell_35_102 (.BL(BL102),.BLN(BLN102),.WL(WL35));
sram_cell_6t_5 inst_cell_35_103 (.BL(BL103),.BLN(BLN103),.WL(WL35));
sram_cell_6t_5 inst_cell_35_104 (.BL(BL104),.BLN(BLN104),.WL(WL35));
sram_cell_6t_5 inst_cell_35_105 (.BL(BL105),.BLN(BLN105),.WL(WL35));
sram_cell_6t_5 inst_cell_35_106 (.BL(BL106),.BLN(BLN106),.WL(WL35));
sram_cell_6t_5 inst_cell_35_107 (.BL(BL107),.BLN(BLN107),.WL(WL35));
sram_cell_6t_5 inst_cell_35_108 (.BL(BL108),.BLN(BLN108),.WL(WL35));
sram_cell_6t_5 inst_cell_35_109 (.BL(BL109),.BLN(BLN109),.WL(WL35));
sram_cell_6t_5 inst_cell_35_110 (.BL(BL110),.BLN(BLN110),.WL(WL35));
sram_cell_6t_5 inst_cell_35_111 (.BL(BL111),.BLN(BLN111),.WL(WL35));
sram_cell_6t_5 inst_cell_35_112 (.BL(BL112),.BLN(BLN112),.WL(WL35));
sram_cell_6t_5 inst_cell_35_113 (.BL(BL113),.BLN(BLN113),.WL(WL35));
sram_cell_6t_5 inst_cell_35_114 (.BL(BL114),.BLN(BLN114),.WL(WL35));
sram_cell_6t_5 inst_cell_35_115 (.BL(BL115),.BLN(BLN115),.WL(WL35));
sram_cell_6t_5 inst_cell_35_116 (.BL(BL116),.BLN(BLN116),.WL(WL35));
sram_cell_6t_5 inst_cell_35_117 (.BL(BL117),.BLN(BLN117),.WL(WL35));
sram_cell_6t_5 inst_cell_35_118 (.BL(BL118),.BLN(BLN118),.WL(WL35));
sram_cell_6t_5 inst_cell_35_119 (.BL(BL119),.BLN(BLN119),.WL(WL35));
sram_cell_6t_5 inst_cell_35_120 (.BL(BL120),.BLN(BLN120),.WL(WL35));
sram_cell_6t_5 inst_cell_35_121 (.BL(BL121),.BLN(BLN121),.WL(WL35));
sram_cell_6t_5 inst_cell_35_122 (.BL(BL122),.BLN(BLN122),.WL(WL35));
sram_cell_6t_5 inst_cell_35_123 (.BL(BL123),.BLN(BLN123),.WL(WL35));
sram_cell_6t_5 inst_cell_35_124 (.BL(BL124),.BLN(BLN124),.WL(WL35));
sram_cell_6t_5 inst_cell_35_125 (.BL(BL125),.BLN(BLN125),.WL(WL35));
sram_cell_6t_5 inst_cell_35_126 (.BL(BL126),.BLN(BLN126),.WL(WL35));
sram_cell_6t_5 inst_cell_35_127 (.BL(BL127),.BLN(BLN127),.WL(WL35));
sram_cell_6t_5 inst_cell_36_0 (.BL(BL0),.BLN(BLN0),.WL(WL36));
sram_cell_6t_5 inst_cell_36_1 (.BL(BL1),.BLN(BLN1),.WL(WL36));
sram_cell_6t_5 inst_cell_36_2 (.BL(BL2),.BLN(BLN2),.WL(WL36));
sram_cell_6t_5 inst_cell_36_3 (.BL(BL3),.BLN(BLN3),.WL(WL36));
sram_cell_6t_5 inst_cell_36_4 (.BL(BL4),.BLN(BLN4),.WL(WL36));
sram_cell_6t_5 inst_cell_36_5 (.BL(BL5),.BLN(BLN5),.WL(WL36));
sram_cell_6t_5 inst_cell_36_6 (.BL(BL6),.BLN(BLN6),.WL(WL36));
sram_cell_6t_5 inst_cell_36_7 (.BL(BL7),.BLN(BLN7),.WL(WL36));
sram_cell_6t_5 inst_cell_36_8 (.BL(BL8),.BLN(BLN8),.WL(WL36));
sram_cell_6t_5 inst_cell_36_9 (.BL(BL9),.BLN(BLN9),.WL(WL36));
sram_cell_6t_5 inst_cell_36_10 (.BL(BL10),.BLN(BLN10),.WL(WL36));
sram_cell_6t_5 inst_cell_36_11 (.BL(BL11),.BLN(BLN11),.WL(WL36));
sram_cell_6t_5 inst_cell_36_12 (.BL(BL12),.BLN(BLN12),.WL(WL36));
sram_cell_6t_5 inst_cell_36_13 (.BL(BL13),.BLN(BLN13),.WL(WL36));
sram_cell_6t_5 inst_cell_36_14 (.BL(BL14),.BLN(BLN14),.WL(WL36));
sram_cell_6t_5 inst_cell_36_15 (.BL(BL15),.BLN(BLN15),.WL(WL36));
sram_cell_6t_5 inst_cell_36_16 (.BL(BL16),.BLN(BLN16),.WL(WL36));
sram_cell_6t_5 inst_cell_36_17 (.BL(BL17),.BLN(BLN17),.WL(WL36));
sram_cell_6t_5 inst_cell_36_18 (.BL(BL18),.BLN(BLN18),.WL(WL36));
sram_cell_6t_5 inst_cell_36_19 (.BL(BL19),.BLN(BLN19),.WL(WL36));
sram_cell_6t_5 inst_cell_36_20 (.BL(BL20),.BLN(BLN20),.WL(WL36));
sram_cell_6t_5 inst_cell_36_21 (.BL(BL21),.BLN(BLN21),.WL(WL36));
sram_cell_6t_5 inst_cell_36_22 (.BL(BL22),.BLN(BLN22),.WL(WL36));
sram_cell_6t_5 inst_cell_36_23 (.BL(BL23),.BLN(BLN23),.WL(WL36));
sram_cell_6t_5 inst_cell_36_24 (.BL(BL24),.BLN(BLN24),.WL(WL36));
sram_cell_6t_5 inst_cell_36_25 (.BL(BL25),.BLN(BLN25),.WL(WL36));
sram_cell_6t_5 inst_cell_36_26 (.BL(BL26),.BLN(BLN26),.WL(WL36));
sram_cell_6t_5 inst_cell_36_27 (.BL(BL27),.BLN(BLN27),.WL(WL36));
sram_cell_6t_5 inst_cell_36_28 (.BL(BL28),.BLN(BLN28),.WL(WL36));
sram_cell_6t_5 inst_cell_36_29 (.BL(BL29),.BLN(BLN29),.WL(WL36));
sram_cell_6t_5 inst_cell_36_30 (.BL(BL30),.BLN(BLN30),.WL(WL36));
sram_cell_6t_5 inst_cell_36_31 (.BL(BL31),.BLN(BLN31),.WL(WL36));
sram_cell_6t_5 inst_cell_36_32 (.BL(BL32),.BLN(BLN32),.WL(WL36));
sram_cell_6t_5 inst_cell_36_33 (.BL(BL33),.BLN(BLN33),.WL(WL36));
sram_cell_6t_5 inst_cell_36_34 (.BL(BL34),.BLN(BLN34),.WL(WL36));
sram_cell_6t_5 inst_cell_36_35 (.BL(BL35),.BLN(BLN35),.WL(WL36));
sram_cell_6t_5 inst_cell_36_36 (.BL(BL36),.BLN(BLN36),.WL(WL36));
sram_cell_6t_5 inst_cell_36_37 (.BL(BL37),.BLN(BLN37),.WL(WL36));
sram_cell_6t_5 inst_cell_36_38 (.BL(BL38),.BLN(BLN38),.WL(WL36));
sram_cell_6t_5 inst_cell_36_39 (.BL(BL39),.BLN(BLN39),.WL(WL36));
sram_cell_6t_5 inst_cell_36_40 (.BL(BL40),.BLN(BLN40),.WL(WL36));
sram_cell_6t_5 inst_cell_36_41 (.BL(BL41),.BLN(BLN41),.WL(WL36));
sram_cell_6t_5 inst_cell_36_42 (.BL(BL42),.BLN(BLN42),.WL(WL36));
sram_cell_6t_5 inst_cell_36_43 (.BL(BL43),.BLN(BLN43),.WL(WL36));
sram_cell_6t_5 inst_cell_36_44 (.BL(BL44),.BLN(BLN44),.WL(WL36));
sram_cell_6t_5 inst_cell_36_45 (.BL(BL45),.BLN(BLN45),.WL(WL36));
sram_cell_6t_5 inst_cell_36_46 (.BL(BL46),.BLN(BLN46),.WL(WL36));
sram_cell_6t_5 inst_cell_36_47 (.BL(BL47),.BLN(BLN47),.WL(WL36));
sram_cell_6t_5 inst_cell_36_48 (.BL(BL48),.BLN(BLN48),.WL(WL36));
sram_cell_6t_5 inst_cell_36_49 (.BL(BL49),.BLN(BLN49),.WL(WL36));
sram_cell_6t_5 inst_cell_36_50 (.BL(BL50),.BLN(BLN50),.WL(WL36));
sram_cell_6t_5 inst_cell_36_51 (.BL(BL51),.BLN(BLN51),.WL(WL36));
sram_cell_6t_5 inst_cell_36_52 (.BL(BL52),.BLN(BLN52),.WL(WL36));
sram_cell_6t_5 inst_cell_36_53 (.BL(BL53),.BLN(BLN53),.WL(WL36));
sram_cell_6t_5 inst_cell_36_54 (.BL(BL54),.BLN(BLN54),.WL(WL36));
sram_cell_6t_5 inst_cell_36_55 (.BL(BL55),.BLN(BLN55),.WL(WL36));
sram_cell_6t_5 inst_cell_36_56 (.BL(BL56),.BLN(BLN56),.WL(WL36));
sram_cell_6t_5 inst_cell_36_57 (.BL(BL57),.BLN(BLN57),.WL(WL36));
sram_cell_6t_5 inst_cell_36_58 (.BL(BL58),.BLN(BLN58),.WL(WL36));
sram_cell_6t_5 inst_cell_36_59 (.BL(BL59),.BLN(BLN59),.WL(WL36));
sram_cell_6t_5 inst_cell_36_60 (.BL(BL60),.BLN(BLN60),.WL(WL36));
sram_cell_6t_5 inst_cell_36_61 (.BL(BL61),.BLN(BLN61),.WL(WL36));
sram_cell_6t_5 inst_cell_36_62 (.BL(BL62),.BLN(BLN62),.WL(WL36));
sram_cell_6t_5 inst_cell_36_63 (.BL(BL63),.BLN(BLN63),.WL(WL36));
sram_cell_6t_5 inst_cell_36_64 (.BL(BL64),.BLN(BLN64),.WL(WL36));
sram_cell_6t_5 inst_cell_36_65 (.BL(BL65),.BLN(BLN65),.WL(WL36));
sram_cell_6t_5 inst_cell_36_66 (.BL(BL66),.BLN(BLN66),.WL(WL36));
sram_cell_6t_5 inst_cell_36_67 (.BL(BL67),.BLN(BLN67),.WL(WL36));
sram_cell_6t_5 inst_cell_36_68 (.BL(BL68),.BLN(BLN68),.WL(WL36));
sram_cell_6t_5 inst_cell_36_69 (.BL(BL69),.BLN(BLN69),.WL(WL36));
sram_cell_6t_5 inst_cell_36_70 (.BL(BL70),.BLN(BLN70),.WL(WL36));
sram_cell_6t_5 inst_cell_36_71 (.BL(BL71),.BLN(BLN71),.WL(WL36));
sram_cell_6t_5 inst_cell_36_72 (.BL(BL72),.BLN(BLN72),.WL(WL36));
sram_cell_6t_5 inst_cell_36_73 (.BL(BL73),.BLN(BLN73),.WL(WL36));
sram_cell_6t_5 inst_cell_36_74 (.BL(BL74),.BLN(BLN74),.WL(WL36));
sram_cell_6t_5 inst_cell_36_75 (.BL(BL75),.BLN(BLN75),.WL(WL36));
sram_cell_6t_5 inst_cell_36_76 (.BL(BL76),.BLN(BLN76),.WL(WL36));
sram_cell_6t_5 inst_cell_36_77 (.BL(BL77),.BLN(BLN77),.WL(WL36));
sram_cell_6t_5 inst_cell_36_78 (.BL(BL78),.BLN(BLN78),.WL(WL36));
sram_cell_6t_5 inst_cell_36_79 (.BL(BL79),.BLN(BLN79),.WL(WL36));
sram_cell_6t_5 inst_cell_36_80 (.BL(BL80),.BLN(BLN80),.WL(WL36));
sram_cell_6t_5 inst_cell_36_81 (.BL(BL81),.BLN(BLN81),.WL(WL36));
sram_cell_6t_5 inst_cell_36_82 (.BL(BL82),.BLN(BLN82),.WL(WL36));
sram_cell_6t_5 inst_cell_36_83 (.BL(BL83),.BLN(BLN83),.WL(WL36));
sram_cell_6t_5 inst_cell_36_84 (.BL(BL84),.BLN(BLN84),.WL(WL36));
sram_cell_6t_5 inst_cell_36_85 (.BL(BL85),.BLN(BLN85),.WL(WL36));
sram_cell_6t_5 inst_cell_36_86 (.BL(BL86),.BLN(BLN86),.WL(WL36));
sram_cell_6t_5 inst_cell_36_87 (.BL(BL87),.BLN(BLN87),.WL(WL36));
sram_cell_6t_5 inst_cell_36_88 (.BL(BL88),.BLN(BLN88),.WL(WL36));
sram_cell_6t_5 inst_cell_36_89 (.BL(BL89),.BLN(BLN89),.WL(WL36));
sram_cell_6t_5 inst_cell_36_90 (.BL(BL90),.BLN(BLN90),.WL(WL36));
sram_cell_6t_5 inst_cell_36_91 (.BL(BL91),.BLN(BLN91),.WL(WL36));
sram_cell_6t_5 inst_cell_36_92 (.BL(BL92),.BLN(BLN92),.WL(WL36));
sram_cell_6t_5 inst_cell_36_93 (.BL(BL93),.BLN(BLN93),.WL(WL36));
sram_cell_6t_5 inst_cell_36_94 (.BL(BL94),.BLN(BLN94),.WL(WL36));
sram_cell_6t_5 inst_cell_36_95 (.BL(BL95),.BLN(BLN95),.WL(WL36));
sram_cell_6t_5 inst_cell_36_96 (.BL(BL96),.BLN(BLN96),.WL(WL36));
sram_cell_6t_5 inst_cell_36_97 (.BL(BL97),.BLN(BLN97),.WL(WL36));
sram_cell_6t_5 inst_cell_36_98 (.BL(BL98),.BLN(BLN98),.WL(WL36));
sram_cell_6t_5 inst_cell_36_99 (.BL(BL99),.BLN(BLN99),.WL(WL36));
sram_cell_6t_5 inst_cell_36_100 (.BL(BL100),.BLN(BLN100),.WL(WL36));
sram_cell_6t_5 inst_cell_36_101 (.BL(BL101),.BLN(BLN101),.WL(WL36));
sram_cell_6t_5 inst_cell_36_102 (.BL(BL102),.BLN(BLN102),.WL(WL36));
sram_cell_6t_5 inst_cell_36_103 (.BL(BL103),.BLN(BLN103),.WL(WL36));
sram_cell_6t_5 inst_cell_36_104 (.BL(BL104),.BLN(BLN104),.WL(WL36));
sram_cell_6t_5 inst_cell_36_105 (.BL(BL105),.BLN(BLN105),.WL(WL36));
sram_cell_6t_5 inst_cell_36_106 (.BL(BL106),.BLN(BLN106),.WL(WL36));
sram_cell_6t_5 inst_cell_36_107 (.BL(BL107),.BLN(BLN107),.WL(WL36));
sram_cell_6t_5 inst_cell_36_108 (.BL(BL108),.BLN(BLN108),.WL(WL36));
sram_cell_6t_5 inst_cell_36_109 (.BL(BL109),.BLN(BLN109),.WL(WL36));
sram_cell_6t_5 inst_cell_36_110 (.BL(BL110),.BLN(BLN110),.WL(WL36));
sram_cell_6t_5 inst_cell_36_111 (.BL(BL111),.BLN(BLN111),.WL(WL36));
sram_cell_6t_5 inst_cell_36_112 (.BL(BL112),.BLN(BLN112),.WL(WL36));
sram_cell_6t_5 inst_cell_36_113 (.BL(BL113),.BLN(BLN113),.WL(WL36));
sram_cell_6t_5 inst_cell_36_114 (.BL(BL114),.BLN(BLN114),.WL(WL36));
sram_cell_6t_5 inst_cell_36_115 (.BL(BL115),.BLN(BLN115),.WL(WL36));
sram_cell_6t_5 inst_cell_36_116 (.BL(BL116),.BLN(BLN116),.WL(WL36));
sram_cell_6t_5 inst_cell_36_117 (.BL(BL117),.BLN(BLN117),.WL(WL36));
sram_cell_6t_5 inst_cell_36_118 (.BL(BL118),.BLN(BLN118),.WL(WL36));
sram_cell_6t_5 inst_cell_36_119 (.BL(BL119),.BLN(BLN119),.WL(WL36));
sram_cell_6t_5 inst_cell_36_120 (.BL(BL120),.BLN(BLN120),.WL(WL36));
sram_cell_6t_5 inst_cell_36_121 (.BL(BL121),.BLN(BLN121),.WL(WL36));
sram_cell_6t_5 inst_cell_36_122 (.BL(BL122),.BLN(BLN122),.WL(WL36));
sram_cell_6t_5 inst_cell_36_123 (.BL(BL123),.BLN(BLN123),.WL(WL36));
sram_cell_6t_5 inst_cell_36_124 (.BL(BL124),.BLN(BLN124),.WL(WL36));
sram_cell_6t_5 inst_cell_36_125 (.BL(BL125),.BLN(BLN125),.WL(WL36));
sram_cell_6t_5 inst_cell_36_126 (.BL(BL126),.BLN(BLN126),.WL(WL36));
sram_cell_6t_5 inst_cell_36_127 (.BL(BL127),.BLN(BLN127),.WL(WL36));
sram_cell_6t_5 inst_cell_37_0 (.BL(BL0),.BLN(BLN0),.WL(WL37));
sram_cell_6t_5 inst_cell_37_1 (.BL(BL1),.BLN(BLN1),.WL(WL37));
sram_cell_6t_5 inst_cell_37_2 (.BL(BL2),.BLN(BLN2),.WL(WL37));
sram_cell_6t_5 inst_cell_37_3 (.BL(BL3),.BLN(BLN3),.WL(WL37));
sram_cell_6t_5 inst_cell_37_4 (.BL(BL4),.BLN(BLN4),.WL(WL37));
sram_cell_6t_5 inst_cell_37_5 (.BL(BL5),.BLN(BLN5),.WL(WL37));
sram_cell_6t_5 inst_cell_37_6 (.BL(BL6),.BLN(BLN6),.WL(WL37));
sram_cell_6t_5 inst_cell_37_7 (.BL(BL7),.BLN(BLN7),.WL(WL37));
sram_cell_6t_5 inst_cell_37_8 (.BL(BL8),.BLN(BLN8),.WL(WL37));
sram_cell_6t_5 inst_cell_37_9 (.BL(BL9),.BLN(BLN9),.WL(WL37));
sram_cell_6t_5 inst_cell_37_10 (.BL(BL10),.BLN(BLN10),.WL(WL37));
sram_cell_6t_5 inst_cell_37_11 (.BL(BL11),.BLN(BLN11),.WL(WL37));
sram_cell_6t_5 inst_cell_37_12 (.BL(BL12),.BLN(BLN12),.WL(WL37));
sram_cell_6t_5 inst_cell_37_13 (.BL(BL13),.BLN(BLN13),.WL(WL37));
sram_cell_6t_5 inst_cell_37_14 (.BL(BL14),.BLN(BLN14),.WL(WL37));
sram_cell_6t_5 inst_cell_37_15 (.BL(BL15),.BLN(BLN15),.WL(WL37));
sram_cell_6t_5 inst_cell_37_16 (.BL(BL16),.BLN(BLN16),.WL(WL37));
sram_cell_6t_5 inst_cell_37_17 (.BL(BL17),.BLN(BLN17),.WL(WL37));
sram_cell_6t_5 inst_cell_37_18 (.BL(BL18),.BLN(BLN18),.WL(WL37));
sram_cell_6t_5 inst_cell_37_19 (.BL(BL19),.BLN(BLN19),.WL(WL37));
sram_cell_6t_5 inst_cell_37_20 (.BL(BL20),.BLN(BLN20),.WL(WL37));
sram_cell_6t_5 inst_cell_37_21 (.BL(BL21),.BLN(BLN21),.WL(WL37));
sram_cell_6t_5 inst_cell_37_22 (.BL(BL22),.BLN(BLN22),.WL(WL37));
sram_cell_6t_5 inst_cell_37_23 (.BL(BL23),.BLN(BLN23),.WL(WL37));
sram_cell_6t_5 inst_cell_37_24 (.BL(BL24),.BLN(BLN24),.WL(WL37));
sram_cell_6t_5 inst_cell_37_25 (.BL(BL25),.BLN(BLN25),.WL(WL37));
sram_cell_6t_5 inst_cell_37_26 (.BL(BL26),.BLN(BLN26),.WL(WL37));
sram_cell_6t_5 inst_cell_37_27 (.BL(BL27),.BLN(BLN27),.WL(WL37));
sram_cell_6t_5 inst_cell_37_28 (.BL(BL28),.BLN(BLN28),.WL(WL37));
sram_cell_6t_5 inst_cell_37_29 (.BL(BL29),.BLN(BLN29),.WL(WL37));
sram_cell_6t_5 inst_cell_37_30 (.BL(BL30),.BLN(BLN30),.WL(WL37));
sram_cell_6t_5 inst_cell_37_31 (.BL(BL31),.BLN(BLN31),.WL(WL37));
sram_cell_6t_5 inst_cell_37_32 (.BL(BL32),.BLN(BLN32),.WL(WL37));
sram_cell_6t_5 inst_cell_37_33 (.BL(BL33),.BLN(BLN33),.WL(WL37));
sram_cell_6t_5 inst_cell_37_34 (.BL(BL34),.BLN(BLN34),.WL(WL37));
sram_cell_6t_5 inst_cell_37_35 (.BL(BL35),.BLN(BLN35),.WL(WL37));
sram_cell_6t_5 inst_cell_37_36 (.BL(BL36),.BLN(BLN36),.WL(WL37));
sram_cell_6t_5 inst_cell_37_37 (.BL(BL37),.BLN(BLN37),.WL(WL37));
sram_cell_6t_5 inst_cell_37_38 (.BL(BL38),.BLN(BLN38),.WL(WL37));
sram_cell_6t_5 inst_cell_37_39 (.BL(BL39),.BLN(BLN39),.WL(WL37));
sram_cell_6t_5 inst_cell_37_40 (.BL(BL40),.BLN(BLN40),.WL(WL37));
sram_cell_6t_5 inst_cell_37_41 (.BL(BL41),.BLN(BLN41),.WL(WL37));
sram_cell_6t_5 inst_cell_37_42 (.BL(BL42),.BLN(BLN42),.WL(WL37));
sram_cell_6t_5 inst_cell_37_43 (.BL(BL43),.BLN(BLN43),.WL(WL37));
sram_cell_6t_5 inst_cell_37_44 (.BL(BL44),.BLN(BLN44),.WL(WL37));
sram_cell_6t_5 inst_cell_37_45 (.BL(BL45),.BLN(BLN45),.WL(WL37));
sram_cell_6t_5 inst_cell_37_46 (.BL(BL46),.BLN(BLN46),.WL(WL37));
sram_cell_6t_5 inst_cell_37_47 (.BL(BL47),.BLN(BLN47),.WL(WL37));
sram_cell_6t_5 inst_cell_37_48 (.BL(BL48),.BLN(BLN48),.WL(WL37));
sram_cell_6t_5 inst_cell_37_49 (.BL(BL49),.BLN(BLN49),.WL(WL37));
sram_cell_6t_5 inst_cell_37_50 (.BL(BL50),.BLN(BLN50),.WL(WL37));
sram_cell_6t_5 inst_cell_37_51 (.BL(BL51),.BLN(BLN51),.WL(WL37));
sram_cell_6t_5 inst_cell_37_52 (.BL(BL52),.BLN(BLN52),.WL(WL37));
sram_cell_6t_5 inst_cell_37_53 (.BL(BL53),.BLN(BLN53),.WL(WL37));
sram_cell_6t_5 inst_cell_37_54 (.BL(BL54),.BLN(BLN54),.WL(WL37));
sram_cell_6t_5 inst_cell_37_55 (.BL(BL55),.BLN(BLN55),.WL(WL37));
sram_cell_6t_5 inst_cell_37_56 (.BL(BL56),.BLN(BLN56),.WL(WL37));
sram_cell_6t_5 inst_cell_37_57 (.BL(BL57),.BLN(BLN57),.WL(WL37));
sram_cell_6t_5 inst_cell_37_58 (.BL(BL58),.BLN(BLN58),.WL(WL37));
sram_cell_6t_5 inst_cell_37_59 (.BL(BL59),.BLN(BLN59),.WL(WL37));
sram_cell_6t_5 inst_cell_37_60 (.BL(BL60),.BLN(BLN60),.WL(WL37));
sram_cell_6t_5 inst_cell_37_61 (.BL(BL61),.BLN(BLN61),.WL(WL37));
sram_cell_6t_5 inst_cell_37_62 (.BL(BL62),.BLN(BLN62),.WL(WL37));
sram_cell_6t_5 inst_cell_37_63 (.BL(BL63),.BLN(BLN63),.WL(WL37));
sram_cell_6t_5 inst_cell_37_64 (.BL(BL64),.BLN(BLN64),.WL(WL37));
sram_cell_6t_5 inst_cell_37_65 (.BL(BL65),.BLN(BLN65),.WL(WL37));
sram_cell_6t_5 inst_cell_37_66 (.BL(BL66),.BLN(BLN66),.WL(WL37));
sram_cell_6t_5 inst_cell_37_67 (.BL(BL67),.BLN(BLN67),.WL(WL37));
sram_cell_6t_5 inst_cell_37_68 (.BL(BL68),.BLN(BLN68),.WL(WL37));
sram_cell_6t_5 inst_cell_37_69 (.BL(BL69),.BLN(BLN69),.WL(WL37));
sram_cell_6t_5 inst_cell_37_70 (.BL(BL70),.BLN(BLN70),.WL(WL37));
sram_cell_6t_5 inst_cell_37_71 (.BL(BL71),.BLN(BLN71),.WL(WL37));
sram_cell_6t_5 inst_cell_37_72 (.BL(BL72),.BLN(BLN72),.WL(WL37));
sram_cell_6t_5 inst_cell_37_73 (.BL(BL73),.BLN(BLN73),.WL(WL37));
sram_cell_6t_5 inst_cell_37_74 (.BL(BL74),.BLN(BLN74),.WL(WL37));
sram_cell_6t_5 inst_cell_37_75 (.BL(BL75),.BLN(BLN75),.WL(WL37));
sram_cell_6t_5 inst_cell_37_76 (.BL(BL76),.BLN(BLN76),.WL(WL37));
sram_cell_6t_5 inst_cell_37_77 (.BL(BL77),.BLN(BLN77),.WL(WL37));
sram_cell_6t_5 inst_cell_37_78 (.BL(BL78),.BLN(BLN78),.WL(WL37));
sram_cell_6t_5 inst_cell_37_79 (.BL(BL79),.BLN(BLN79),.WL(WL37));
sram_cell_6t_5 inst_cell_37_80 (.BL(BL80),.BLN(BLN80),.WL(WL37));
sram_cell_6t_5 inst_cell_37_81 (.BL(BL81),.BLN(BLN81),.WL(WL37));
sram_cell_6t_5 inst_cell_37_82 (.BL(BL82),.BLN(BLN82),.WL(WL37));
sram_cell_6t_5 inst_cell_37_83 (.BL(BL83),.BLN(BLN83),.WL(WL37));
sram_cell_6t_5 inst_cell_37_84 (.BL(BL84),.BLN(BLN84),.WL(WL37));
sram_cell_6t_5 inst_cell_37_85 (.BL(BL85),.BLN(BLN85),.WL(WL37));
sram_cell_6t_5 inst_cell_37_86 (.BL(BL86),.BLN(BLN86),.WL(WL37));
sram_cell_6t_5 inst_cell_37_87 (.BL(BL87),.BLN(BLN87),.WL(WL37));
sram_cell_6t_5 inst_cell_37_88 (.BL(BL88),.BLN(BLN88),.WL(WL37));
sram_cell_6t_5 inst_cell_37_89 (.BL(BL89),.BLN(BLN89),.WL(WL37));
sram_cell_6t_5 inst_cell_37_90 (.BL(BL90),.BLN(BLN90),.WL(WL37));
sram_cell_6t_5 inst_cell_37_91 (.BL(BL91),.BLN(BLN91),.WL(WL37));
sram_cell_6t_5 inst_cell_37_92 (.BL(BL92),.BLN(BLN92),.WL(WL37));
sram_cell_6t_5 inst_cell_37_93 (.BL(BL93),.BLN(BLN93),.WL(WL37));
sram_cell_6t_5 inst_cell_37_94 (.BL(BL94),.BLN(BLN94),.WL(WL37));
sram_cell_6t_5 inst_cell_37_95 (.BL(BL95),.BLN(BLN95),.WL(WL37));
sram_cell_6t_5 inst_cell_37_96 (.BL(BL96),.BLN(BLN96),.WL(WL37));
sram_cell_6t_5 inst_cell_37_97 (.BL(BL97),.BLN(BLN97),.WL(WL37));
sram_cell_6t_5 inst_cell_37_98 (.BL(BL98),.BLN(BLN98),.WL(WL37));
sram_cell_6t_5 inst_cell_37_99 (.BL(BL99),.BLN(BLN99),.WL(WL37));
sram_cell_6t_5 inst_cell_37_100 (.BL(BL100),.BLN(BLN100),.WL(WL37));
sram_cell_6t_5 inst_cell_37_101 (.BL(BL101),.BLN(BLN101),.WL(WL37));
sram_cell_6t_5 inst_cell_37_102 (.BL(BL102),.BLN(BLN102),.WL(WL37));
sram_cell_6t_5 inst_cell_37_103 (.BL(BL103),.BLN(BLN103),.WL(WL37));
sram_cell_6t_5 inst_cell_37_104 (.BL(BL104),.BLN(BLN104),.WL(WL37));
sram_cell_6t_5 inst_cell_37_105 (.BL(BL105),.BLN(BLN105),.WL(WL37));
sram_cell_6t_5 inst_cell_37_106 (.BL(BL106),.BLN(BLN106),.WL(WL37));
sram_cell_6t_5 inst_cell_37_107 (.BL(BL107),.BLN(BLN107),.WL(WL37));
sram_cell_6t_5 inst_cell_37_108 (.BL(BL108),.BLN(BLN108),.WL(WL37));
sram_cell_6t_5 inst_cell_37_109 (.BL(BL109),.BLN(BLN109),.WL(WL37));
sram_cell_6t_5 inst_cell_37_110 (.BL(BL110),.BLN(BLN110),.WL(WL37));
sram_cell_6t_5 inst_cell_37_111 (.BL(BL111),.BLN(BLN111),.WL(WL37));
sram_cell_6t_5 inst_cell_37_112 (.BL(BL112),.BLN(BLN112),.WL(WL37));
sram_cell_6t_5 inst_cell_37_113 (.BL(BL113),.BLN(BLN113),.WL(WL37));
sram_cell_6t_5 inst_cell_37_114 (.BL(BL114),.BLN(BLN114),.WL(WL37));
sram_cell_6t_5 inst_cell_37_115 (.BL(BL115),.BLN(BLN115),.WL(WL37));
sram_cell_6t_5 inst_cell_37_116 (.BL(BL116),.BLN(BLN116),.WL(WL37));
sram_cell_6t_5 inst_cell_37_117 (.BL(BL117),.BLN(BLN117),.WL(WL37));
sram_cell_6t_5 inst_cell_37_118 (.BL(BL118),.BLN(BLN118),.WL(WL37));
sram_cell_6t_5 inst_cell_37_119 (.BL(BL119),.BLN(BLN119),.WL(WL37));
sram_cell_6t_5 inst_cell_37_120 (.BL(BL120),.BLN(BLN120),.WL(WL37));
sram_cell_6t_5 inst_cell_37_121 (.BL(BL121),.BLN(BLN121),.WL(WL37));
sram_cell_6t_5 inst_cell_37_122 (.BL(BL122),.BLN(BLN122),.WL(WL37));
sram_cell_6t_5 inst_cell_37_123 (.BL(BL123),.BLN(BLN123),.WL(WL37));
sram_cell_6t_5 inst_cell_37_124 (.BL(BL124),.BLN(BLN124),.WL(WL37));
sram_cell_6t_5 inst_cell_37_125 (.BL(BL125),.BLN(BLN125),.WL(WL37));
sram_cell_6t_5 inst_cell_37_126 (.BL(BL126),.BLN(BLN126),.WL(WL37));
sram_cell_6t_5 inst_cell_37_127 (.BL(BL127),.BLN(BLN127),.WL(WL37));
sram_cell_6t_5 inst_cell_38_0 (.BL(BL0),.BLN(BLN0),.WL(WL38));
sram_cell_6t_5 inst_cell_38_1 (.BL(BL1),.BLN(BLN1),.WL(WL38));
sram_cell_6t_5 inst_cell_38_2 (.BL(BL2),.BLN(BLN2),.WL(WL38));
sram_cell_6t_5 inst_cell_38_3 (.BL(BL3),.BLN(BLN3),.WL(WL38));
sram_cell_6t_5 inst_cell_38_4 (.BL(BL4),.BLN(BLN4),.WL(WL38));
sram_cell_6t_5 inst_cell_38_5 (.BL(BL5),.BLN(BLN5),.WL(WL38));
sram_cell_6t_5 inst_cell_38_6 (.BL(BL6),.BLN(BLN6),.WL(WL38));
sram_cell_6t_5 inst_cell_38_7 (.BL(BL7),.BLN(BLN7),.WL(WL38));
sram_cell_6t_5 inst_cell_38_8 (.BL(BL8),.BLN(BLN8),.WL(WL38));
sram_cell_6t_5 inst_cell_38_9 (.BL(BL9),.BLN(BLN9),.WL(WL38));
sram_cell_6t_5 inst_cell_38_10 (.BL(BL10),.BLN(BLN10),.WL(WL38));
sram_cell_6t_5 inst_cell_38_11 (.BL(BL11),.BLN(BLN11),.WL(WL38));
sram_cell_6t_5 inst_cell_38_12 (.BL(BL12),.BLN(BLN12),.WL(WL38));
sram_cell_6t_5 inst_cell_38_13 (.BL(BL13),.BLN(BLN13),.WL(WL38));
sram_cell_6t_5 inst_cell_38_14 (.BL(BL14),.BLN(BLN14),.WL(WL38));
sram_cell_6t_5 inst_cell_38_15 (.BL(BL15),.BLN(BLN15),.WL(WL38));
sram_cell_6t_5 inst_cell_38_16 (.BL(BL16),.BLN(BLN16),.WL(WL38));
sram_cell_6t_5 inst_cell_38_17 (.BL(BL17),.BLN(BLN17),.WL(WL38));
sram_cell_6t_5 inst_cell_38_18 (.BL(BL18),.BLN(BLN18),.WL(WL38));
sram_cell_6t_5 inst_cell_38_19 (.BL(BL19),.BLN(BLN19),.WL(WL38));
sram_cell_6t_5 inst_cell_38_20 (.BL(BL20),.BLN(BLN20),.WL(WL38));
sram_cell_6t_5 inst_cell_38_21 (.BL(BL21),.BLN(BLN21),.WL(WL38));
sram_cell_6t_5 inst_cell_38_22 (.BL(BL22),.BLN(BLN22),.WL(WL38));
sram_cell_6t_5 inst_cell_38_23 (.BL(BL23),.BLN(BLN23),.WL(WL38));
sram_cell_6t_5 inst_cell_38_24 (.BL(BL24),.BLN(BLN24),.WL(WL38));
sram_cell_6t_5 inst_cell_38_25 (.BL(BL25),.BLN(BLN25),.WL(WL38));
sram_cell_6t_5 inst_cell_38_26 (.BL(BL26),.BLN(BLN26),.WL(WL38));
sram_cell_6t_5 inst_cell_38_27 (.BL(BL27),.BLN(BLN27),.WL(WL38));
sram_cell_6t_5 inst_cell_38_28 (.BL(BL28),.BLN(BLN28),.WL(WL38));
sram_cell_6t_5 inst_cell_38_29 (.BL(BL29),.BLN(BLN29),.WL(WL38));
sram_cell_6t_5 inst_cell_38_30 (.BL(BL30),.BLN(BLN30),.WL(WL38));
sram_cell_6t_5 inst_cell_38_31 (.BL(BL31),.BLN(BLN31),.WL(WL38));
sram_cell_6t_5 inst_cell_38_32 (.BL(BL32),.BLN(BLN32),.WL(WL38));
sram_cell_6t_5 inst_cell_38_33 (.BL(BL33),.BLN(BLN33),.WL(WL38));
sram_cell_6t_5 inst_cell_38_34 (.BL(BL34),.BLN(BLN34),.WL(WL38));
sram_cell_6t_5 inst_cell_38_35 (.BL(BL35),.BLN(BLN35),.WL(WL38));
sram_cell_6t_5 inst_cell_38_36 (.BL(BL36),.BLN(BLN36),.WL(WL38));
sram_cell_6t_5 inst_cell_38_37 (.BL(BL37),.BLN(BLN37),.WL(WL38));
sram_cell_6t_5 inst_cell_38_38 (.BL(BL38),.BLN(BLN38),.WL(WL38));
sram_cell_6t_5 inst_cell_38_39 (.BL(BL39),.BLN(BLN39),.WL(WL38));
sram_cell_6t_5 inst_cell_38_40 (.BL(BL40),.BLN(BLN40),.WL(WL38));
sram_cell_6t_5 inst_cell_38_41 (.BL(BL41),.BLN(BLN41),.WL(WL38));
sram_cell_6t_5 inst_cell_38_42 (.BL(BL42),.BLN(BLN42),.WL(WL38));
sram_cell_6t_5 inst_cell_38_43 (.BL(BL43),.BLN(BLN43),.WL(WL38));
sram_cell_6t_5 inst_cell_38_44 (.BL(BL44),.BLN(BLN44),.WL(WL38));
sram_cell_6t_5 inst_cell_38_45 (.BL(BL45),.BLN(BLN45),.WL(WL38));
sram_cell_6t_5 inst_cell_38_46 (.BL(BL46),.BLN(BLN46),.WL(WL38));
sram_cell_6t_5 inst_cell_38_47 (.BL(BL47),.BLN(BLN47),.WL(WL38));
sram_cell_6t_5 inst_cell_38_48 (.BL(BL48),.BLN(BLN48),.WL(WL38));
sram_cell_6t_5 inst_cell_38_49 (.BL(BL49),.BLN(BLN49),.WL(WL38));
sram_cell_6t_5 inst_cell_38_50 (.BL(BL50),.BLN(BLN50),.WL(WL38));
sram_cell_6t_5 inst_cell_38_51 (.BL(BL51),.BLN(BLN51),.WL(WL38));
sram_cell_6t_5 inst_cell_38_52 (.BL(BL52),.BLN(BLN52),.WL(WL38));
sram_cell_6t_5 inst_cell_38_53 (.BL(BL53),.BLN(BLN53),.WL(WL38));
sram_cell_6t_5 inst_cell_38_54 (.BL(BL54),.BLN(BLN54),.WL(WL38));
sram_cell_6t_5 inst_cell_38_55 (.BL(BL55),.BLN(BLN55),.WL(WL38));
sram_cell_6t_5 inst_cell_38_56 (.BL(BL56),.BLN(BLN56),.WL(WL38));
sram_cell_6t_5 inst_cell_38_57 (.BL(BL57),.BLN(BLN57),.WL(WL38));
sram_cell_6t_5 inst_cell_38_58 (.BL(BL58),.BLN(BLN58),.WL(WL38));
sram_cell_6t_5 inst_cell_38_59 (.BL(BL59),.BLN(BLN59),.WL(WL38));
sram_cell_6t_5 inst_cell_38_60 (.BL(BL60),.BLN(BLN60),.WL(WL38));
sram_cell_6t_5 inst_cell_38_61 (.BL(BL61),.BLN(BLN61),.WL(WL38));
sram_cell_6t_5 inst_cell_38_62 (.BL(BL62),.BLN(BLN62),.WL(WL38));
sram_cell_6t_5 inst_cell_38_63 (.BL(BL63),.BLN(BLN63),.WL(WL38));
sram_cell_6t_5 inst_cell_38_64 (.BL(BL64),.BLN(BLN64),.WL(WL38));
sram_cell_6t_5 inst_cell_38_65 (.BL(BL65),.BLN(BLN65),.WL(WL38));
sram_cell_6t_5 inst_cell_38_66 (.BL(BL66),.BLN(BLN66),.WL(WL38));
sram_cell_6t_5 inst_cell_38_67 (.BL(BL67),.BLN(BLN67),.WL(WL38));
sram_cell_6t_5 inst_cell_38_68 (.BL(BL68),.BLN(BLN68),.WL(WL38));
sram_cell_6t_5 inst_cell_38_69 (.BL(BL69),.BLN(BLN69),.WL(WL38));
sram_cell_6t_5 inst_cell_38_70 (.BL(BL70),.BLN(BLN70),.WL(WL38));
sram_cell_6t_5 inst_cell_38_71 (.BL(BL71),.BLN(BLN71),.WL(WL38));
sram_cell_6t_5 inst_cell_38_72 (.BL(BL72),.BLN(BLN72),.WL(WL38));
sram_cell_6t_5 inst_cell_38_73 (.BL(BL73),.BLN(BLN73),.WL(WL38));
sram_cell_6t_5 inst_cell_38_74 (.BL(BL74),.BLN(BLN74),.WL(WL38));
sram_cell_6t_5 inst_cell_38_75 (.BL(BL75),.BLN(BLN75),.WL(WL38));
sram_cell_6t_5 inst_cell_38_76 (.BL(BL76),.BLN(BLN76),.WL(WL38));
sram_cell_6t_5 inst_cell_38_77 (.BL(BL77),.BLN(BLN77),.WL(WL38));
sram_cell_6t_5 inst_cell_38_78 (.BL(BL78),.BLN(BLN78),.WL(WL38));
sram_cell_6t_5 inst_cell_38_79 (.BL(BL79),.BLN(BLN79),.WL(WL38));
sram_cell_6t_5 inst_cell_38_80 (.BL(BL80),.BLN(BLN80),.WL(WL38));
sram_cell_6t_5 inst_cell_38_81 (.BL(BL81),.BLN(BLN81),.WL(WL38));
sram_cell_6t_5 inst_cell_38_82 (.BL(BL82),.BLN(BLN82),.WL(WL38));
sram_cell_6t_5 inst_cell_38_83 (.BL(BL83),.BLN(BLN83),.WL(WL38));
sram_cell_6t_5 inst_cell_38_84 (.BL(BL84),.BLN(BLN84),.WL(WL38));
sram_cell_6t_5 inst_cell_38_85 (.BL(BL85),.BLN(BLN85),.WL(WL38));
sram_cell_6t_5 inst_cell_38_86 (.BL(BL86),.BLN(BLN86),.WL(WL38));
sram_cell_6t_5 inst_cell_38_87 (.BL(BL87),.BLN(BLN87),.WL(WL38));
sram_cell_6t_5 inst_cell_38_88 (.BL(BL88),.BLN(BLN88),.WL(WL38));
sram_cell_6t_5 inst_cell_38_89 (.BL(BL89),.BLN(BLN89),.WL(WL38));
sram_cell_6t_5 inst_cell_38_90 (.BL(BL90),.BLN(BLN90),.WL(WL38));
sram_cell_6t_5 inst_cell_38_91 (.BL(BL91),.BLN(BLN91),.WL(WL38));
sram_cell_6t_5 inst_cell_38_92 (.BL(BL92),.BLN(BLN92),.WL(WL38));
sram_cell_6t_5 inst_cell_38_93 (.BL(BL93),.BLN(BLN93),.WL(WL38));
sram_cell_6t_5 inst_cell_38_94 (.BL(BL94),.BLN(BLN94),.WL(WL38));
sram_cell_6t_5 inst_cell_38_95 (.BL(BL95),.BLN(BLN95),.WL(WL38));
sram_cell_6t_5 inst_cell_38_96 (.BL(BL96),.BLN(BLN96),.WL(WL38));
sram_cell_6t_5 inst_cell_38_97 (.BL(BL97),.BLN(BLN97),.WL(WL38));
sram_cell_6t_5 inst_cell_38_98 (.BL(BL98),.BLN(BLN98),.WL(WL38));
sram_cell_6t_5 inst_cell_38_99 (.BL(BL99),.BLN(BLN99),.WL(WL38));
sram_cell_6t_5 inst_cell_38_100 (.BL(BL100),.BLN(BLN100),.WL(WL38));
sram_cell_6t_5 inst_cell_38_101 (.BL(BL101),.BLN(BLN101),.WL(WL38));
sram_cell_6t_5 inst_cell_38_102 (.BL(BL102),.BLN(BLN102),.WL(WL38));
sram_cell_6t_5 inst_cell_38_103 (.BL(BL103),.BLN(BLN103),.WL(WL38));
sram_cell_6t_5 inst_cell_38_104 (.BL(BL104),.BLN(BLN104),.WL(WL38));
sram_cell_6t_5 inst_cell_38_105 (.BL(BL105),.BLN(BLN105),.WL(WL38));
sram_cell_6t_5 inst_cell_38_106 (.BL(BL106),.BLN(BLN106),.WL(WL38));
sram_cell_6t_5 inst_cell_38_107 (.BL(BL107),.BLN(BLN107),.WL(WL38));
sram_cell_6t_5 inst_cell_38_108 (.BL(BL108),.BLN(BLN108),.WL(WL38));
sram_cell_6t_5 inst_cell_38_109 (.BL(BL109),.BLN(BLN109),.WL(WL38));
sram_cell_6t_5 inst_cell_38_110 (.BL(BL110),.BLN(BLN110),.WL(WL38));
sram_cell_6t_5 inst_cell_38_111 (.BL(BL111),.BLN(BLN111),.WL(WL38));
sram_cell_6t_5 inst_cell_38_112 (.BL(BL112),.BLN(BLN112),.WL(WL38));
sram_cell_6t_5 inst_cell_38_113 (.BL(BL113),.BLN(BLN113),.WL(WL38));
sram_cell_6t_5 inst_cell_38_114 (.BL(BL114),.BLN(BLN114),.WL(WL38));
sram_cell_6t_5 inst_cell_38_115 (.BL(BL115),.BLN(BLN115),.WL(WL38));
sram_cell_6t_5 inst_cell_38_116 (.BL(BL116),.BLN(BLN116),.WL(WL38));
sram_cell_6t_5 inst_cell_38_117 (.BL(BL117),.BLN(BLN117),.WL(WL38));
sram_cell_6t_5 inst_cell_38_118 (.BL(BL118),.BLN(BLN118),.WL(WL38));
sram_cell_6t_5 inst_cell_38_119 (.BL(BL119),.BLN(BLN119),.WL(WL38));
sram_cell_6t_5 inst_cell_38_120 (.BL(BL120),.BLN(BLN120),.WL(WL38));
sram_cell_6t_5 inst_cell_38_121 (.BL(BL121),.BLN(BLN121),.WL(WL38));
sram_cell_6t_5 inst_cell_38_122 (.BL(BL122),.BLN(BLN122),.WL(WL38));
sram_cell_6t_5 inst_cell_38_123 (.BL(BL123),.BLN(BLN123),.WL(WL38));
sram_cell_6t_5 inst_cell_38_124 (.BL(BL124),.BLN(BLN124),.WL(WL38));
sram_cell_6t_5 inst_cell_38_125 (.BL(BL125),.BLN(BLN125),.WL(WL38));
sram_cell_6t_5 inst_cell_38_126 (.BL(BL126),.BLN(BLN126),.WL(WL38));
sram_cell_6t_5 inst_cell_38_127 (.BL(BL127),.BLN(BLN127),.WL(WL38));
sram_cell_6t_5 inst_cell_39_0 (.BL(BL0),.BLN(BLN0),.WL(WL39));
sram_cell_6t_5 inst_cell_39_1 (.BL(BL1),.BLN(BLN1),.WL(WL39));
sram_cell_6t_5 inst_cell_39_2 (.BL(BL2),.BLN(BLN2),.WL(WL39));
sram_cell_6t_5 inst_cell_39_3 (.BL(BL3),.BLN(BLN3),.WL(WL39));
sram_cell_6t_5 inst_cell_39_4 (.BL(BL4),.BLN(BLN4),.WL(WL39));
sram_cell_6t_5 inst_cell_39_5 (.BL(BL5),.BLN(BLN5),.WL(WL39));
sram_cell_6t_5 inst_cell_39_6 (.BL(BL6),.BLN(BLN6),.WL(WL39));
sram_cell_6t_5 inst_cell_39_7 (.BL(BL7),.BLN(BLN7),.WL(WL39));
sram_cell_6t_5 inst_cell_39_8 (.BL(BL8),.BLN(BLN8),.WL(WL39));
sram_cell_6t_5 inst_cell_39_9 (.BL(BL9),.BLN(BLN9),.WL(WL39));
sram_cell_6t_5 inst_cell_39_10 (.BL(BL10),.BLN(BLN10),.WL(WL39));
sram_cell_6t_5 inst_cell_39_11 (.BL(BL11),.BLN(BLN11),.WL(WL39));
sram_cell_6t_5 inst_cell_39_12 (.BL(BL12),.BLN(BLN12),.WL(WL39));
sram_cell_6t_5 inst_cell_39_13 (.BL(BL13),.BLN(BLN13),.WL(WL39));
sram_cell_6t_5 inst_cell_39_14 (.BL(BL14),.BLN(BLN14),.WL(WL39));
sram_cell_6t_5 inst_cell_39_15 (.BL(BL15),.BLN(BLN15),.WL(WL39));
sram_cell_6t_5 inst_cell_39_16 (.BL(BL16),.BLN(BLN16),.WL(WL39));
sram_cell_6t_5 inst_cell_39_17 (.BL(BL17),.BLN(BLN17),.WL(WL39));
sram_cell_6t_5 inst_cell_39_18 (.BL(BL18),.BLN(BLN18),.WL(WL39));
sram_cell_6t_5 inst_cell_39_19 (.BL(BL19),.BLN(BLN19),.WL(WL39));
sram_cell_6t_5 inst_cell_39_20 (.BL(BL20),.BLN(BLN20),.WL(WL39));
sram_cell_6t_5 inst_cell_39_21 (.BL(BL21),.BLN(BLN21),.WL(WL39));
sram_cell_6t_5 inst_cell_39_22 (.BL(BL22),.BLN(BLN22),.WL(WL39));
sram_cell_6t_5 inst_cell_39_23 (.BL(BL23),.BLN(BLN23),.WL(WL39));
sram_cell_6t_5 inst_cell_39_24 (.BL(BL24),.BLN(BLN24),.WL(WL39));
sram_cell_6t_5 inst_cell_39_25 (.BL(BL25),.BLN(BLN25),.WL(WL39));
sram_cell_6t_5 inst_cell_39_26 (.BL(BL26),.BLN(BLN26),.WL(WL39));
sram_cell_6t_5 inst_cell_39_27 (.BL(BL27),.BLN(BLN27),.WL(WL39));
sram_cell_6t_5 inst_cell_39_28 (.BL(BL28),.BLN(BLN28),.WL(WL39));
sram_cell_6t_5 inst_cell_39_29 (.BL(BL29),.BLN(BLN29),.WL(WL39));
sram_cell_6t_5 inst_cell_39_30 (.BL(BL30),.BLN(BLN30),.WL(WL39));
sram_cell_6t_5 inst_cell_39_31 (.BL(BL31),.BLN(BLN31),.WL(WL39));
sram_cell_6t_5 inst_cell_39_32 (.BL(BL32),.BLN(BLN32),.WL(WL39));
sram_cell_6t_5 inst_cell_39_33 (.BL(BL33),.BLN(BLN33),.WL(WL39));
sram_cell_6t_5 inst_cell_39_34 (.BL(BL34),.BLN(BLN34),.WL(WL39));
sram_cell_6t_5 inst_cell_39_35 (.BL(BL35),.BLN(BLN35),.WL(WL39));
sram_cell_6t_5 inst_cell_39_36 (.BL(BL36),.BLN(BLN36),.WL(WL39));
sram_cell_6t_5 inst_cell_39_37 (.BL(BL37),.BLN(BLN37),.WL(WL39));
sram_cell_6t_5 inst_cell_39_38 (.BL(BL38),.BLN(BLN38),.WL(WL39));
sram_cell_6t_5 inst_cell_39_39 (.BL(BL39),.BLN(BLN39),.WL(WL39));
sram_cell_6t_5 inst_cell_39_40 (.BL(BL40),.BLN(BLN40),.WL(WL39));
sram_cell_6t_5 inst_cell_39_41 (.BL(BL41),.BLN(BLN41),.WL(WL39));
sram_cell_6t_5 inst_cell_39_42 (.BL(BL42),.BLN(BLN42),.WL(WL39));
sram_cell_6t_5 inst_cell_39_43 (.BL(BL43),.BLN(BLN43),.WL(WL39));
sram_cell_6t_5 inst_cell_39_44 (.BL(BL44),.BLN(BLN44),.WL(WL39));
sram_cell_6t_5 inst_cell_39_45 (.BL(BL45),.BLN(BLN45),.WL(WL39));
sram_cell_6t_5 inst_cell_39_46 (.BL(BL46),.BLN(BLN46),.WL(WL39));
sram_cell_6t_5 inst_cell_39_47 (.BL(BL47),.BLN(BLN47),.WL(WL39));
sram_cell_6t_5 inst_cell_39_48 (.BL(BL48),.BLN(BLN48),.WL(WL39));
sram_cell_6t_5 inst_cell_39_49 (.BL(BL49),.BLN(BLN49),.WL(WL39));
sram_cell_6t_5 inst_cell_39_50 (.BL(BL50),.BLN(BLN50),.WL(WL39));
sram_cell_6t_5 inst_cell_39_51 (.BL(BL51),.BLN(BLN51),.WL(WL39));
sram_cell_6t_5 inst_cell_39_52 (.BL(BL52),.BLN(BLN52),.WL(WL39));
sram_cell_6t_5 inst_cell_39_53 (.BL(BL53),.BLN(BLN53),.WL(WL39));
sram_cell_6t_5 inst_cell_39_54 (.BL(BL54),.BLN(BLN54),.WL(WL39));
sram_cell_6t_5 inst_cell_39_55 (.BL(BL55),.BLN(BLN55),.WL(WL39));
sram_cell_6t_5 inst_cell_39_56 (.BL(BL56),.BLN(BLN56),.WL(WL39));
sram_cell_6t_5 inst_cell_39_57 (.BL(BL57),.BLN(BLN57),.WL(WL39));
sram_cell_6t_5 inst_cell_39_58 (.BL(BL58),.BLN(BLN58),.WL(WL39));
sram_cell_6t_5 inst_cell_39_59 (.BL(BL59),.BLN(BLN59),.WL(WL39));
sram_cell_6t_5 inst_cell_39_60 (.BL(BL60),.BLN(BLN60),.WL(WL39));
sram_cell_6t_5 inst_cell_39_61 (.BL(BL61),.BLN(BLN61),.WL(WL39));
sram_cell_6t_5 inst_cell_39_62 (.BL(BL62),.BLN(BLN62),.WL(WL39));
sram_cell_6t_5 inst_cell_39_63 (.BL(BL63),.BLN(BLN63),.WL(WL39));
sram_cell_6t_5 inst_cell_39_64 (.BL(BL64),.BLN(BLN64),.WL(WL39));
sram_cell_6t_5 inst_cell_39_65 (.BL(BL65),.BLN(BLN65),.WL(WL39));
sram_cell_6t_5 inst_cell_39_66 (.BL(BL66),.BLN(BLN66),.WL(WL39));
sram_cell_6t_5 inst_cell_39_67 (.BL(BL67),.BLN(BLN67),.WL(WL39));
sram_cell_6t_5 inst_cell_39_68 (.BL(BL68),.BLN(BLN68),.WL(WL39));
sram_cell_6t_5 inst_cell_39_69 (.BL(BL69),.BLN(BLN69),.WL(WL39));
sram_cell_6t_5 inst_cell_39_70 (.BL(BL70),.BLN(BLN70),.WL(WL39));
sram_cell_6t_5 inst_cell_39_71 (.BL(BL71),.BLN(BLN71),.WL(WL39));
sram_cell_6t_5 inst_cell_39_72 (.BL(BL72),.BLN(BLN72),.WL(WL39));
sram_cell_6t_5 inst_cell_39_73 (.BL(BL73),.BLN(BLN73),.WL(WL39));
sram_cell_6t_5 inst_cell_39_74 (.BL(BL74),.BLN(BLN74),.WL(WL39));
sram_cell_6t_5 inst_cell_39_75 (.BL(BL75),.BLN(BLN75),.WL(WL39));
sram_cell_6t_5 inst_cell_39_76 (.BL(BL76),.BLN(BLN76),.WL(WL39));
sram_cell_6t_5 inst_cell_39_77 (.BL(BL77),.BLN(BLN77),.WL(WL39));
sram_cell_6t_5 inst_cell_39_78 (.BL(BL78),.BLN(BLN78),.WL(WL39));
sram_cell_6t_5 inst_cell_39_79 (.BL(BL79),.BLN(BLN79),.WL(WL39));
sram_cell_6t_5 inst_cell_39_80 (.BL(BL80),.BLN(BLN80),.WL(WL39));
sram_cell_6t_5 inst_cell_39_81 (.BL(BL81),.BLN(BLN81),.WL(WL39));
sram_cell_6t_5 inst_cell_39_82 (.BL(BL82),.BLN(BLN82),.WL(WL39));
sram_cell_6t_5 inst_cell_39_83 (.BL(BL83),.BLN(BLN83),.WL(WL39));
sram_cell_6t_5 inst_cell_39_84 (.BL(BL84),.BLN(BLN84),.WL(WL39));
sram_cell_6t_5 inst_cell_39_85 (.BL(BL85),.BLN(BLN85),.WL(WL39));
sram_cell_6t_5 inst_cell_39_86 (.BL(BL86),.BLN(BLN86),.WL(WL39));
sram_cell_6t_5 inst_cell_39_87 (.BL(BL87),.BLN(BLN87),.WL(WL39));
sram_cell_6t_5 inst_cell_39_88 (.BL(BL88),.BLN(BLN88),.WL(WL39));
sram_cell_6t_5 inst_cell_39_89 (.BL(BL89),.BLN(BLN89),.WL(WL39));
sram_cell_6t_5 inst_cell_39_90 (.BL(BL90),.BLN(BLN90),.WL(WL39));
sram_cell_6t_5 inst_cell_39_91 (.BL(BL91),.BLN(BLN91),.WL(WL39));
sram_cell_6t_5 inst_cell_39_92 (.BL(BL92),.BLN(BLN92),.WL(WL39));
sram_cell_6t_5 inst_cell_39_93 (.BL(BL93),.BLN(BLN93),.WL(WL39));
sram_cell_6t_5 inst_cell_39_94 (.BL(BL94),.BLN(BLN94),.WL(WL39));
sram_cell_6t_5 inst_cell_39_95 (.BL(BL95),.BLN(BLN95),.WL(WL39));
sram_cell_6t_5 inst_cell_39_96 (.BL(BL96),.BLN(BLN96),.WL(WL39));
sram_cell_6t_5 inst_cell_39_97 (.BL(BL97),.BLN(BLN97),.WL(WL39));
sram_cell_6t_5 inst_cell_39_98 (.BL(BL98),.BLN(BLN98),.WL(WL39));
sram_cell_6t_5 inst_cell_39_99 (.BL(BL99),.BLN(BLN99),.WL(WL39));
sram_cell_6t_5 inst_cell_39_100 (.BL(BL100),.BLN(BLN100),.WL(WL39));
sram_cell_6t_5 inst_cell_39_101 (.BL(BL101),.BLN(BLN101),.WL(WL39));
sram_cell_6t_5 inst_cell_39_102 (.BL(BL102),.BLN(BLN102),.WL(WL39));
sram_cell_6t_5 inst_cell_39_103 (.BL(BL103),.BLN(BLN103),.WL(WL39));
sram_cell_6t_5 inst_cell_39_104 (.BL(BL104),.BLN(BLN104),.WL(WL39));
sram_cell_6t_5 inst_cell_39_105 (.BL(BL105),.BLN(BLN105),.WL(WL39));
sram_cell_6t_5 inst_cell_39_106 (.BL(BL106),.BLN(BLN106),.WL(WL39));
sram_cell_6t_5 inst_cell_39_107 (.BL(BL107),.BLN(BLN107),.WL(WL39));
sram_cell_6t_5 inst_cell_39_108 (.BL(BL108),.BLN(BLN108),.WL(WL39));
sram_cell_6t_5 inst_cell_39_109 (.BL(BL109),.BLN(BLN109),.WL(WL39));
sram_cell_6t_5 inst_cell_39_110 (.BL(BL110),.BLN(BLN110),.WL(WL39));
sram_cell_6t_5 inst_cell_39_111 (.BL(BL111),.BLN(BLN111),.WL(WL39));
sram_cell_6t_5 inst_cell_39_112 (.BL(BL112),.BLN(BLN112),.WL(WL39));
sram_cell_6t_5 inst_cell_39_113 (.BL(BL113),.BLN(BLN113),.WL(WL39));
sram_cell_6t_5 inst_cell_39_114 (.BL(BL114),.BLN(BLN114),.WL(WL39));
sram_cell_6t_5 inst_cell_39_115 (.BL(BL115),.BLN(BLN115),.WL(WL39));
sram_cell_6t_5 inst_cell_39_116 (.BL(BL116),.BLN(BLN116),.WL(WL39));
sram_cell_6t_5 inst_cell_39_117 (.BL(BL117),.BLN(BLN117),.WL(WL39));
sram_cell_6t_5 inst_cell_39_118 (.BL(BL118),.BLN(BLN118),.WL(WL39));
sram_cell_6t_5 inst_cell_39_119 (.BL(BL119),.BLN(BLN119),.WL(WL39));
sram_cell_6t_5 inst_cell_39_120 (.BL(BL120),.BLN(BLN120),.WL(WL39));
sram_cell_6t_5 inst_cell_39_121 (.BL(BL121),.BLN(BLN121),.WL(WL39));
sram_cell_6t_5 inst_cell_39_122 (.BL(BL122),.BLN(BLN122),.WL(WL39));
sram_cell_6t_5 inst_cell_39_123 (.BL(BL123),.BLN(BLN123),.WL(WL39));
sram_cell_6t_5 inst_cell_39_124 (.BL(BL124),.BLN(BLN124),.WL(WL39));
sram_cell_6t_5 inst_cell_39_125 (.BL(BL125),.BLN(BLN125),.WL(WL39));
sram_cell_6t_5 inst_cell_39_126 (.BL(BL126),.BLN(BLN126),.WL(WL39));
sram_cell_6t_5 inst_cell_39_127 (.BL(BL127),.BLN(BLN127),.WL(WL39));
sram_cell_6t_5 inst_cell_40_0 (.BL(BL0),.BLN(BLN0),.WL(WL40));
sram_cell_6t_5 inst_cell_40_1 (.BL(BL1),.BLN(BLN1),.WL(WL40));
sram_cell_6t_5 inst_cell_40_2 (.BL(BL2),.BLN(BLN2),.WL(WL40));
sram_cell_6t_5 inst_cell_40_3 (.BL(BL3),.BLN(BLN3),.WL(WL40));
sram_cell_6t_5 inst_cell_40_4 (.BL(BL4),.BLN(BLN4),.WL(WL40));
sram_cell_6t_5 inst_cell_40_5 (.BL(BL5),.BLN(BLN5),.WL(WL40));
sram_cell_6t_5 inst_cell_40_6 (.BL(BL6),.BLN(BLN6),.WL(WL40));
sram_cell_6t_5 inst_cell_40_7 (.BL(BL7),.BLN(BLN7),.WL(WL40));
sram_cell_6t_5 inst_cell_40_8 (.BL(BL8),.BLN(BLN8),.WL(WL40));
sram_cell_6t_5 inst_cell_40_9 (.BL(BL9),.BLN(BLN9),.WL(WL40));
sram_cell_6t_5 inst_cell_40_10 (.BL(BL10),.BLN(BLN10),.WL(WL40));
sram_cell_6t_5 inst_cell_40_11 (.BL(BL11),.BLN(BLN11),.WL(WL40));
sram_cell_6t_5 inst_cell_40_12 (.BL(BL12),.BLN(BLN12),.WL(WL40));
sram_cell_6t_5 inst_cell_40_13 (.BL(BL13),.BLN(BLN13),.WL(WL40));
sram_cell_6t_5 inst_cell_40_14 (.BL(BL14),.BLN(BLN14),.WL(WL40));
sram_cell_6t_5 inst_cell_40_15 (.BL(BL15),.BLN(BLN15),.WL(WL40));
sram_cell_6t_5 inst_cell_40_16 (.BL(BL16),.BLN(BLN16),.WL(WL40));
sram_cell_6t_5 inst_cell_40_17 (.BL(BL17),.BLN(BLN17),.WL(WL40));
sram_cell_6t_5 inst_cell_40_18 (.BL(BL18),.BLN(BLN18),.WL(WL40));
sram_cell_6t_5 inst_cell_40_19 (.BL(BL19),.BLN(BLN19),.WL(WL40));
sram_cell_6t_5 inst_cell_40_20 (.BL(BL20),.BLN(BLN20),.WL(WL40));
sram_cell_6t_5 inst_cell_40_21 (.BL(BL21),.BLN(BLN21),.WL(WL40));
sram_cell_6t_5 inst_cell_40_22 (.BL(BL22),.BLN(BLN22),.WL(WL40));
sram_cell_6t_5 inst_cell_40_23 (.BL(BL23),.BLN(BLN23),.WL(WL40));
sram_cell_6t_5 inst_cell_40_24 (.BL(BL24),.BLN(BLN24),.WL(WL40));
sram_cell_6t_5 inst_cell_40_25 (.BL(BL25),.BLN(BLN25),.WL(WL40));
sram_cell_6t_5 inst_cell_40_26 (.BL(BL26),.BLN(BLN26),.WL(WL40));
sram_cell_6t_5 inst_cell_40_27 (.BL(BL27),.BLN(BLN27),.WL(WL40));
sram_cell_6t_5 inst_cell_40_28 (.BL(BL28),.BLN(BLN28),.WL(WL40));
sram_cell_6t_5 inst_cell_40_29 (.BL(BL29),.BLN(BLN29),.WL(WL40));
sram_cell_6t_5 inst_cell_40_30 (.BL(BL30),.BLN(BLN30),.WL(WL40));
sram_cell_6t_5 inst_cell_40_31 (.BL(BL31),.BLN(BLN31),.WL(WL40));
sram_cell_6t_5 inst_cell_40_32 (.BL(BL32),.BLN(BLN32),.WL(WL40));
sram_cell_6t_5 inst_cell_40_33 (.BL(BL33),.BLN(BLN33),.WL(WL40));
sram_cell_6t_5 inst_cell_40_34 (.BL(BL34),.BLN(BLN34),.WL(WL40));
sram_cell_6t_5 inst_cell_40_35 (.BL(BL35),.BLN(BLN35),.WL(WL40));
sram_cell_6t_5 inst_cell_40_36 (.BL(BL36),.BLN(BLN36),.WL(WL40));
sram_cell_6t_5 inst_cell_40_37 (.BL(BL37),.BLN(BLN37),.WL(WL40));
sram_cell_6t_5 inst_cell_40_38 (.BL(BL38),.BLN(BLN38),.WL(WL40));
sram_cell_6t_5 inst_cell_40_39 (.BL(BL39),.BLN(BLN39),.WL(WL40));
sram_cell_6t_5 inst_cell_40_40 (.BL(BL40),.BLN(BLN40),.WL(WL40));
sram_cell_6t_5 inst_cell_40_41 (.BL(BL41),.BLN(BLN41),.WL(WL40));
sram_cell_6t_5 inst_cell_40_42 (.BL(BL42),.BLN(BLN42),.WL(WL40));
sram_cell_6t_5 inst_cell_40_43 (.BL(BL43),.BLN(BLN43),.WL(WL40));
sram_cell_6t_5 inst_cell_40_44 (.BL(BL44),.BLN(BLN44),.WL(WL40));
sram_cell_6t_5 inst_cell_40_45 (.BL(BL45),.BLN(BLN45),.WL(WL40));
sram_cell_6t_5 inst_cell_40_46 (.BL(BL46),.BLN(BLN46),.WL(WL40));
sram_cell_6t_5 inst_cell_40_47 (.BL(BL47),.BLN(BLN47),.WL(WL40));
sram_cell_6t_5 inst_cell_40_48 (.BL(BL48),.BLN(BLN48),.WL(WL40));
sram_cell_6t_5 inst_cell_40_49 (.BL(BL49),.BLN(BLN49),.WL(WL40));
sram_cell_6t_5 inst_cell_40_50 (.BL(BL50),.BLN(BLN50),.WL(WL40));
sram_cell_6t_5 inst_cell_40_51 (.BL(BL51),.BLN(BLN51),.WL(WL40));
sram_cell_6t_5 inst_cell_40_52 (.BL(BL52),.BLN(BLN52),.WL(WL40));
sram_cell_6t_5 inst_cell_40_53 (.BL(BL53),.BLN(BLN53),.WL(WL40));
sram_cell_6t_5 inst_cell_40_54 (.BL(BL54),.BLN(BLN54),.WL(WL40));
sram_cell_6t_5 inst_cell_40_55 (.BL(BL55),.BLN(BLN55),.WL(WL40));
sram_cell_6t_5 inst_cell_40_56 (.BL(BL56),.BLN(BLN56),.WL(WL40));
sram_cell_6t_5 inst_cell_40_57 (.BL(BL57),.BLN(BLN57),.WL(WL40));
sram_cell_6t_5 inst_cell_40_58 (.BL(BL58),.BLN(BLN58),.WL(WL40));
sram_cell_6t_5 inst_cell_40_59 (.BL(BL59),.BLN(BLN59),.WL(WL40));
sram_cell_6t_5 inst_cell_40_60 (.BL(BL60),.BLN(BLN60),.WL(WL40));
sram_cell_6t_5 inst_cell_40_61 (.BL(BL61),.BLN(BLN61),.WL(WL40));
sram_cell_6t_5 inst_cell_40_62 (.BL(BL62),.BLN(BLN62),.WL(WL40));
sram_cell_6t_5 inst_cell_40_63 (.BL(BL63),.BLN(BLN63),.WL(WL40));
sram_cell_6t_5 inst_cell_40_64 (.BL(BL64),.BLN(BLN64),.WL(WL40));
sram_cell_6t_5 inst_cell_40_65 (.BL(BL65),.BLN(BLN65),.WL(WL40));
sram_cell_6t_5 inst_cell_40_66 (.BL(BL66),.BLN(BLN66),.WL(WL40));
sram_cell_6t_5 inst_cell_40_67 (.BL(BL67),.BLN(BLN67),.WL(WL40));
sram_cell_6t_5 inst_cell_40_68 (.BL(BL68),.BLN(BLN68),.WL(WL40));
sram_cell_6t_5 inst_cell_40_69 (.BL(BL69),.BLN(BLN69),.WL(WL40));
sram_cell_6t_5 inst_cell_40_70 (.BL(BL70),.BLN(BLN70),.WL(WL40));
sram_cell_6t_5 inst_cell_40_71 (.BL(BL71),.BLN(BLN71),.WL(WL40));
sram_cell_6t_5 inst_cell_40_72 (.BL(BL72),.BLN(BLN72),.WL(WL40));
sram_cell_6t_5 inst_cell_40_73 (.BL(BL73),.BLN(BLN73),.WL(WL40));
sram_cell_6t_5 inst_cell_40_74 (.BL(BL74),.BLN(BLN74),.WL(WL40));
sram_cell_6t_5 inst_cell_40_75 (.BL(BL75),.BLN(BLN75),.WL(WL40));
sram_cell_6t_5 inst_cell_40_76 (.BL(BL76),.BLN(BLN76),.WL(WL40));
sram_cell_6t_5 inst_cell_40_77 (.BL(BL77),.BLN(BLN77),.WL(WL40));
sram_cell_6t_5 inst_cell_40_78 (.BL(BL78),.BLN(BLN78),.WL(WL40));
sram_cell_6t_5 inst_cell_40_79 (.BL(BL79),.BLN(BLN79),.WL(WL40));
sram_cell_6t_5 inst_cell_40_80 (.BL(BL80),.BLN(BLN80),.WL(WL40));
sram_cell_6t_5 inst_cell_40_81 (.BL(BL81),.BLN(BLN81),.WL(WL40));
sram_cell_6t_5 inst_cell_40_82 (.BL(BL82),.BLN(BLN82),.WL(WL40));
sram_cell_6t_5 inst_cell_40_83 (.BL(BL83),.BLN(BLN83),.WL(WL40));
sram_cell_6t_5 inst_cell_40_84 (.BL(BL84),.BLN(BLN84),.WL(WL40));
sram_cell_6t_5 inst_cell_40_85 (.BL(BL85),.BLN(BLN85),.WL(WL40));
sram_cell_6t_5 inst_cell_40_86 (.BL(BL86),.BLN(BLN86),.WL(WL40));
sram_cell_6t_5 inst_cell_40_87 (.BL(BL87),.BLN(BLN87),.WL(WL40));
sram_cell_6t_5 inst_cell_40_88 (.BL(BL88),.BLN(BLN88),.WL(WL40));
sram_cell_6t_5 inst_cell_40_89 (.BL(BL89),.BLN(BLN89),.WL(WL40));
sram_cell_6t_5 inst_cell_40_90 (.BL(BL90),.BLN(BLN90),.WL(WL40));
sram_cell_6t_5 inst_cell_40_91 (.BL(BL91),.BLN(BLN91),.WL(WL40));
sram_cell_6t_5 inst_cell_40_92 (.BL(BL92),.BLN(BLN92),.WL(WL40));
sram_cell_6t_5 inst_cell_40_93 (.BL(BL93),.BLN(BLN93),.WL(WL40));
sram_cell_6t_5 inst_cell_40_94 (.BL(BL94),.BLN(BLN94),.WL(WL40));
sram_cell_6t_5 inst_cell_40_95 (.BL(BL95),.BLN(BLN95),.WL(WL40));
sram_cell_6t_5 inst_cell_40_96 (.BL(BL96),.BLN(BLN96),.WL(WL40));
sram_cell_6t_5 inst_cell_40_97 (.BL(BL97),.BLN(BLN97),.WL(WL40));
sram_cell_6t_5 inst_cell_40_98 (.BL(BL98),.BLN(BLN98),.WL(WL40));
sram_cell_6t_5 inst_cell_40_99 (.BL(BL99),.BLN(BLN99),.WL(WL40));
sram_cell_6t_5 inst_cell_40_100 (.BL(BL100),.BLN(BLN100),.WL(WL40));
sram_cell_6t_5 inst_cell_40_101 (.BL(BL101),.BLN(BLN101),.WL(WL40));
sram_cell_6t_5 inst_cell_40_102 (.BL(BL102),.BLN(BLN102),.WL(WL40));
sram_cell_6t_5 inst_cell_40_103 (.BL(BL103),.BLN(BLN103),.WL(WL40));
sram_cell_6t_5 inst_cell_40_104 (.BL(BL104),.BLN(BLN104),.WL(WL40));
sram_cell_6t_5 inst_cell_40_105 (.BL(BL105),.BLN(BLN105),.WL(WL40));
sram_cell_6t_5 inst_cell_40_106 (.BL(BL106),.BLN(BLN106),.WL(WL40));
sram_cell_6t_5 inst_cell_40_107 (.BL(BL107),.BLN(BLN107),.WL(WL40));
sram_cell_6t_5 inst_cell_40_108 (.BL(BL108),.BLN(BLN108),.WL(WL40));
sram_cell_6t_5 inst_cell_40_109 (.BL(BL109),.BLN(BLN109),.WL(WL40));
sram_cell_6t_5 inst_cell_40_110 (.BL(BL110),.BLN(BLN110),.WL(WL40));
sram_cell_6t_5 inst_cell_40_111 (.BL(BL111),.BLN(BLN111),.WL(WL40));
sram_cell_6t_5 inst_cell_40_112 (.BL(BL112),.BLN(BLN112),.WL(WL40));
sram_cell_6t_5 inst_cell_40_113 (.BL(BL113),.BLN(BLN113),.WL(WL40));
sram_cell_6t_5 inst_cell_40_114 (.BL(BL114),.BLN(BLN114),.WL(WL40));
sram_cell_6t_5 inst_cell_40_115 (.BL(BL115),.BLN(BLN115),.WL(WL40));
sram_cell_6t_5 inst_cell_40_116 (.BL(BL116),.BLN(BLN116),.WL(WL40));
sram_cell_6t_5 inst_cell_40_117 (.BL(BL117),.BLN(BLN117),.WL(WL40));
sram_cell_6t_5 inst_cell_40_118 (.BL(BL118),.BLN(BLN118),.WL(WL40));
sram_cell_6t_5 inst_cell_40_119 (.BL(BL119),.BLN(BLN119),.WL(WL40));
sram_cell_6t_5 inst_cell_40_120 (.BL(BL120),.BLN(BLN120),.WL(WL40));
sram_cell_6t_5 inst_cell_40_121 (.BL(BL121),.BLN(BLN121),.WL(WL40));
sram_cell_6t_5 inst_cell_40_122 (.BL(BL122),.BLN(BLN122),.WL(WL40));
sram_cell_6t_5 inst_cell_40_123 (.BL(BL123),.BLN(BLN123),.WL(WL40));
sram_cell_6t_5 inst_cell_40_124 (.BL(BL124),.BLN(BLN124),.WL(WL40));
sram_cell_6t_5 inst_cell_40_125 (.BL(BL125),.BLN(BLN125),.WL(WL40));
sram_cell_6t_5 inst_cell_40_126 (.BL(BL126),.BLN(BLN126),.WL(WL40));
sram_cell_6t_5 inst_cell_40_127 (.BL(BL127),.BLN(BLN127),.WL(WL40));
sram_cell_6t_5 inst_cell_41_0 (.BL(BL0),.BLN(BLN0),.WL(WL41));
sram_cell_6t_5 inst_cell_41_1 (.BL(BL1),.BLN(BLN1),.WL(WL41));
sram_cell_6t_5 inst_cell_41_2 (.BL(BL2),.BLN(BLN2),.WL(WL41));
sram_cell_6t_5 inst_cell_41_3 (.BL(BL3),.BLN(BLN3),.WL(WL41));
sram_cell_6t_5 inst_cell_41_4 (.BL(BL4),.BLN(BLN4),.WL(WL41));
sram_cell_6t_5 inst_cell_41_5 (.BL(BL5),.BLN(BLN5),.WL(WL41));
sram_cell_6t_5 inst_cell_41_6 (.BL(BL6),.BLN(BLN6),.WL(WL41));
sram_cell_6t_5 inst_cell_41_7 (.BL(BL7),.BLN(BLN7),.WL(WL41));
sram_cell_6t_5 inst_cell_41_8 (.BL(BL8),.BLN(BLN8),.WL(WL41));
sram_cell_6t_5 inst_cell_41_9 (.BL(BL9),.BLN(BLN9),.WL(WL41));
sram_cell_6t_5 inst_cell_41_10 (.BL(BL10),.BLN(BLN10),.WL(WL41));
sram_cell_6t_5 inst_cell_41_11 (.BL(BL11),.BLN(BLN11),.WL(WL41));
sram_cell_6t_5 inst_cell_41_12 (.BL(BL12),.BLN(BLN12),.WL(WL41));
sram_cell_6t_5 inst_cell_41_13 (.BL(BL13),.BLN(BLN13),.WL(WL41));
sram_cell_6t_5 inst_cell_41_14 (.BL(BL14),.BLN(BLN14),.WL(WL41));
sram_cell_6t_5 inst_cell_41_15 (.BL(BL15),.BLN(BLN15),.WL(WL41));
sram_cell_6t_5 inst_cell_41_16 (.BL(BL16),.BLN(BLN16),.WL(WL41));
sram_cell_6t_5 inst_cell_41_17 (.BL(BL17),.BLN(BLN17),.WL(WL41));
sram_cell_6t_5 inst_cell_41_18 (.BL(BL18),.BLN(BLN18),.WL(WL41));
sram_cell_6t_5 inst_cell_41_19 (.BL(BL19),.BLN(BLN19),.WL(WL41));
sram_cell_6t_5 inst_cell_41_20 (.BL(BL20),.BLN(BLN20),.WL(WL41));
sram_cell_6t_5 inst_cell_41_21 (.BL(BL21),.BLN(BLN21),.WL(WL41));
sram_cell_6t_5 inst_cell_41_22 (.BL(BL22),.BLN(BLN22),.WL(WL41));
sram_cell_6t_5 inst_cell_41_23 (.BL(BL23),.BLN(BLN23),.WL(WL41));
sram_cell_6t_5 inst_cell_41_24 (.BL(BL24),.BLN(BLN24),.WL(WL41));
sram_cell_6t_5 inst_cell_41_25 (.BL(BL25),.BLN(BLN25),.WL(WL41));
sram_cell_6t_5 inst_cell_41_26 (.BL(BL26),.BLN(BLN26),.WL(WL41));
sram_cell_6t_5 inst_cell_41_27 (.BL(BL27),.BLN(BLN27),.WL(WL41));
sram_cell_6t_5 inst_cell_41_28 (.BL(BL28),.BLN(BLN28),.WL(WL41));
sram_cell_6t_5 inst_cell_41_29 (.BL(BL29),.BLN(BLN29),.WL(WL41));
sram_cell_6t_5 inst_cell_41_30 (.BL(BL30),.BLN(BLN30),.WL(WL41));
sram_cell_6t_5 inst_cell_41_31 (.BL(BL31),.BLN(BLN31),.WL(WL41));
sram_cell_6t_5 inst_cell_41_32 (.BL(BL32),.BLN(BLN32),.WL(WL41));
sram_cell_6t_5 inst_cell_41_33 (.BL(BL33),.BLN(BLN33),.WL(WL41));
sram_cell_6t_5 inst_cell_41_34 (.BL(BL34),.BLN(BLN34),.WL(WL41));
sram_cell_6t_5 inst_cell_41_35 (.BL(BL35),.BLN(BLN35),.WL(WL41));
sram_cell_6t_5 inst_cell_41_36 (.BL(BL36),.BLN(BLN36),.WL(WL41));
sram_cell_6t_5 inst_cell_41_37 (.BL(BL37),.BLN(BLN37),.WL(WL41));
sram_cell_6t_5 inst_cell_41_38 (.BL(BL38),.BLN(BLN38),.WL(WL41));
sram_cell_6t_5 inst_cell_41_39 (.BL(BL39),.BLN(BLN39),.WL(WL41));
sram_cell_6t_5 inst_cell_41_40 (.BL(BL40),.BLN(BLN40),.WL(WL41));
sram_cell_6t_5 inst_cell_41_41 (.BL(BL41),.BLN(BLN41),.WL(WL41));
sram_cell_6t_5 inst_cell_41_42 (.BL(BL42),.BLN(BLN42),.WL(WL41));
sram_cell_6t_5 inst_cell_41_43 (.BL(BL43),.BLN(BLN43),.WL(WL41));
sram_cell_6t_5 inst_cell_41_44 (.BL(BL44),.BLN(BLN44),.WL(WL41));
sram_cell_6t_5 inst_cell_41_45 (.BL(BL45),.BLN(BLN45),.WL(WL41));
sram_cell_6t_5 inst_cell_41_46 (.BL(BL46),.BLN(BLN46),.WL(WL41));
sram_cell_6t_5 inst_cell_41_47 (.BL(BL47),.BLN(BLN47),.WL(WL41));
sram_cell_6t_5 inst_cell_41_48 (.BL(BL48),.BLN(BLN48),.WL(WL41));
sram_cell_6t_5 inst_cell_41_49 (.BL(BL49),.BLN(BLN49),.WL(WL41));
sram_cell_6t_5 inst_cell_41_50 (.BL(BL50),.BLN(BLN50),.WL(WL41));
sram_cell_6t_5 inst_cell_41_51 (.BL(BL51),.BLN(BLN51),.WL(WL41));
sram_cell_6t_5 inst_cell_41_52 (.BL(BL52),.BLN(BLN52),.WL(WL41));
sram_cell_6t_5 inst_cell_41_53 (.BL(BL53),.BLN(BLN53),.WL(WL41));
sram_cell_6t_5 inst_cell_41_54 (.BL(BL54),.BLN(BLN54),.WL(WL41));
sram_cell_6t_5 inst_cell_41_55 (.BL(BL55),.BLN(BLN55),.WL(WL41));
sram_cell_6t_5 inst_cell_41_56 (.BL(BL56),.BLN(BLN56),.WL(WL41));
sram_cell_6t_5 inst_cell_41_57 (.BL(BL57),.BLN(BLN57),.WL(WL41));
sram_cell_6t_5 inst_cell_41_58 (.BL(BL58),.BLN(BLN58),.WL(WL41));
sram_cell_6t_5 inst_cell_41_59 (.BL(BL59),.BLN(BLN59),.WL(WL41));
sram_cell_6t_5 inst_cell_41_60 (.BL(BL60),.BLN(BLN60),.WL(WL41));
sram_cell_6t_5 inst_cell_41_61 (.BL(BL61),.BLN(BLN61),.WL(WL41));
sram_cell_6t_5 inst_cell_41_62 (.BL(BL62),.BLN(BLN62),.WL(WL41));
sram_cell_6t_5 inst_cell_41_63 (.BL(BL63),.BLN(BLN63),.WL(WL41));
sram_cell_6t_5 inst_cell_41_64 (.BL(BL64),.BLN(BLN64),.WL(WL41));
sram_cell_6t_5 inst_cell_41_65 (.BL(BL65),.BLN(BLN65),.WL(WL41));
sram_cell_6t_5 inst_cell_41_66 (.BL(BL66),.BLN(BLN66),.WL(WL41));
sram_cell_6t_5 inst_cell_41_67 (.BL(BL67),.BLN(BLN67),.WL(WL41));
sram_cell_6t_5 inst_cell_41_68 (.BL(BL68),.BLN(BLN68),.WL(WL41));
sram_cell_6t_5 inst_cell_41_69 (.BL(BL69),.BLN(BLN69),.WL(WL41));
sram_cell_6t_5 inst_cell_41_70 (.BL(BL70),.BLN(BLN70),.WL(WL41));
sram_cell_6t_5 inst_cell_41_71 (.BL(BL71),.BLN(BLN71),.WL(WL41));
sram_cell_6t_5 inst_cell_41_72 (.BL(BL72),.BLN(BLN72),.WL(WL41));
sram_cell_6t_5 inst_cell_41_73 (.BL(BL73),.BLN(BLN73),.WL(WL41));
sram_cell_6t_5 inst_cell_41_74 (.BL(BL74),.BLN(BLN74),.WL(WL41));
sram_cell_6t_5 inst_cell_41_75 (.BL(BL75),.BLN(BLN75),.WL(WL41));
sram_cell_6t_5 inst_cell_41_76 (.BL(BL76),.BLN(BLN76),.WL(WL41));
sram_cell_6t_5 inst_cell_41_77 (.BL(BL77),.BLN(BLN77),.WL(WL41));
sram_cell_6t_5 inst_cell_41_78 (.BL(BL78),.BLN(BLN78),.WL(WL41));
sram_cell_6t_5 inst_cell_41_79 (.BL(BL79),.BLN(BLN79),.WL(WL41));
sram_cell_6t_5 inst_cell_41_80 (.BL(BL80),.BLN(BLN80),.WL(WL41));
sram_cell_6t_5 inst_cell_41_81 (.BL(BL81),.BLN(BLN81),.WL(WL41));
sram_cell_6t_5 inst_cell_41_82 (.BL(BL82),.BLN(BLN82),.WL(WL41));
sram_cell_6t_5 inst_cell_41_83 (.BL(BL83),.BLN(BLN83),.WL(WL41));
sram_cell_6t_5 inst_cell_41_84 (.BL(BL84),.BLN(BLN84),.WL(WL41));
sram_cell_6t_5 inst_cell_41_85 (.BL(BL85),.BLN(BLN85),.WL(WL41));
sram_cell_6t_5 inst_cell_41_86 (.BL(BL86),.BLN(BLN86),.WL(WL41));
sram_cell_6t_5 inst_cell_41_87 (.BL(BL87),.BLN(BLN87),.WL(WL41));
sram_cell_6t_5 inst_cell_41_88 (.BL(BL88),.BLN(BLN88),.WL(WL41));
sram_cell_6t_5 inst_cell_41_89 (.BL(BL89),.BLN(BLN89),.WL(WL41));
sram_cell_6t_5 inst_cell_41_90 (.BL(BL90),.BLN(BLN90),.WL(WL41));
sram_cell_6t_5 inst_cell_41_91 (.BL(BL91),.BLN(BLN91),.WL(WL41));
sram_cell_6t_5 inst_cell_41_92 (.BL(BL92),.BLN(BLN92),.WL(WL41));
sram_cell_6t_5 inst_cell_41_93 (.BL(BL93),.BLN(BLN93),.WL(WL41));
sram_cell_6t_5 inst_cell_41_94 (.BL(BL94),.BLN(BLN94),.WL(WL41));
sram_cell_6t_5 inst_cell_41_95 (.BL(BL95),.BLN(BLN95),.WL(WL41));
sram_cell_6t_5 inst_cell_41_96 (.BL(BL96),.BLN(BLN96),.WL(WL41));
sram_cell_6t_5 inst_cell_41_97 (.BL(BL97),.BLN(BLN97),.WL(WL41));
sram_cell_6t_5 inst_cell_41_98 (.BL(BL98),.BLN(BLN98),.WL(WL41));
sram_cell_6t_5 inst_cell_41_99 (.BL(BL99),.BLN(BLN99),.WL(WL41));
sram_cell_6t_5 inst_cell_41_100 (.BL(BL100),.BLN(BLN100),.WL(WL41));
sram_cell_6t_5 inst_cell_41_101 (.BL(BL101),.BLN(BLN101),.WL(WL41));
sram_cell_6t_5 inst_cell_41_102 (.BL(BL102),.BLN(BLN102),.WL(WL41));
sram_cell_6t_5 inst_cell_41_103 (.BL(BL103),.BLN(BLN103),.WL(WL41));
sram_cell_6t_5 inst_cell_41_104 (.BL(BL104),.BLN(BLN104),.WL(WL41));
sram_cell_6t_5 inst_cell_41_105 (.BL(BL105),.BLN(BLN105),.WL(WL41));
sram_cell_6t_5 inst_cell_41_106 (.BL(BL106),.BLN(BLN106),.WL(WL41));
sram_cell_6t_5 inst_cell_41_107 (.BL(BL107),.BLN(BLN107),.WL(WL41));
sram_cell_6t_5 inst_cell_41_108 (.BL(BL108),.BLN(BLN108),.WL(WL41));
sram_cell_6t_5 inst_cell_41_109 (.BL(BL109),.BLN(BLN109),.WL(WL41));
sram_cell_6t_5 inst_cell_41_110 (.BL(BL110),.BLN(BLN110),.WL(WL41));
sram_cell_6t_5 inst_cell_41_111 (.BL(BL111),.BLN(BLN111),.WL(WL41));
sram_cell_6t_5 inst_cell_41_112 (.BL(BL112),.BLN(BLN112),.WL(WL41));
sram_cell_6t_5 inst_cell_41_113 (.BL(BL113),.BLN(BLN113),.WL(WL41));
sram_cell_6t_5 inst_cell_41_114 (.BL(BL114),.BLN(BLN114),.WL(WL41));
sram_cell_6t_5 inst_cell_41_115 (.BL(BL115),.BLN(BLN115),.WL(WL41));
sram_cell_6t_5 inst_cell_41_116 (.BL(BL116),.BLN(BLN116),.WL(WL41));
sram_cell_6t_5 inst_cell_41_117 (.BL(BL117),.BLN(BLN117),.WL(WL41));
sram_cell_6t_5 inst_cell_41_118 (.BL(BL118),.BLN(BLN118),.WL(WL41));
sram_cell_6t_5 inst_cell_41_119 (.BL(BL119),.BLN(BLN119),.WL(WL41));
sram_cell_6t_5 inst_cell_41_120 (.BL(BL120),.BLN(BLN120),.WL(WL41));
sram_cell_6t_5 inst_cell_41_121 (.BL(BL121),.BLN(BLN121),.WL(WL41));
sram_cell_6t_5 inst_cell_41_122 (.BL(BL122),.BLN(BLN122),.WL(WL41));
sram_cell_6t_5 inst_cell_41_123 (.BL(BL123),.BLN(BLN123),.WL(WL41));
sram_cell_6t_5 inst_cell_41_124 (.BL(BL124),.BLN(BLN124),.WL(WL41));
sram_cell_6t_5 inst_cell_41_125 (.BL(BL125),.BLN(BLN125),.WL(WL41));
sram_cell_6t_5 inst_cell_41_126 (.BL(BL126),.BLN(BLN126),.WL(WL41));
sram_cell_6t_5 inst_cell_41_127 (.BL(BL127),.BLN(BLN127),.WL(WL41));
sram_cell_6t_5 inst_cell_42_0 (.BL(BL0),.BLN(BLN0),.WL(WL42));
sram_cell_6t_5 inst_cell_42_1 (.BL(BL1),.BLN(BLN1),.WL(WL42));
sram_cell_6t_5 inst_cell_42_2 (.BL(BL2),.BLN(BLN2),.WL(WL42));
sram_cell_6t_5 inst_cell_42_3 (.BL(BL3),.BLN(BLN3),.WL(WL42));
sram_cell_6t_5 inst_cell_42_4 (.BL(BL4),.BLN(BLN4),.WL(WL42));
sram_cell_6t_5 inst_cell_42_5 (.BL(BL5),.BLN(BLN5),.WL(WL42));
sram_cell_6t_5 inst_cell_42_6 (.BL(BL6),.BLN(BLN6),.WL(WL42));
sram_cell_6t_5 inst_cell_42_7 (.BL(BL7),.BLN(BLN7),.WL(WL42));
sram_cell_6t_5 inst_cell_42_8 (.BL(BL8),.BLN(BLN8),.WL(WL42));
sram_cell_6t_5 inst_cell_42_9 (.BL(BL9),.BLN(BLN9),.WL(WL42));
sram_cell_6t_5 inst_cell_42_10 (.BL(BL10),.BLN(BLN10),.WL(WL42));
sram_cell_6t_5 inst_cell_42_11 (.BL(BL11),.BLN(BLN11),.WL(WL42));
sram_cell_6t_5 inst_cell_42_12 (.BL(BL12),.BLN(BLN12),.WL(WL42));
sram_cell_6t_5 inst_cell_42_13 (.BL(BL13),.BLN(BLN13),.WL(WL42));
sram_cell_6t_5 inst_cell_42_14 (.BL(BL14),.BLN(BLN14),.WL(WL42));
sram_cell_6t_5 inst_cell_42_15 (.BL(BL15),.BLN(BLN15),.WL(WL42));
sram_cell_6t_5 inst_cell_42_16 (.BL(BL16),.BLN(BLN16),.WL(WL42));
sram_cell_6t_5 inst_cell_42_17 (.BL(BL17),.BLN(BLN17),.WL(WL42));
sram_cell_6t_5 inst_cell_42_18 (.BL(BL18),.BLN(BLN18),.WL(WL42));
sram_cell_6t_5 inst_cell_42_19 (.BL(BL19),.BLN(BLN19),.WL(WL42));
sram_cell_6t_5 inst_cell_42_20 (.BL(BL20),.BLN(BLN20),.WL(WL42));
sram_cell_6t_5 inst_cell_42_21 (.BL(BL21),.BLN(BLN21),.WL(WL42));
sram_cell_6t_5 inst_cell_42_22 (.BL(BL22),.BLN(BLN22),.WL(WL42));
sram_cell_6t_5 inst_cell_42_23 (.BL(BL23),.BLN(BLN23),.WL(WL42));
sram_cell_6t_5 inst_cell_42_24 (.BL(BL24),.BLN(BLN24),.WL(WL42));
sram_cell_6t_5 inst_cell_42_25 (.BL(BL25),.BLN(BLN25),.WL(WL42));
sram_cell_6t_5 inst_cell_42_26 (.BL(BL26),.BLN(BLN26),.WL(WL42));
sram_cell_6t_5 inst_cell_42_27 (.BL(BL27),.BLN(BLN27),.WL(WL42));
sram_cell_6t_5 inst_cell_42_28 (.BL(BL28),.BLN(BLN28),.WL(WL42));
sram_cell_6t_5 inst_cell_42_29 (.BL(BL29),.BLN(BLN29),.WL(WL42));
sram_cell_6t_5 inst_cell_42_30 (.BL(BL30),.BLN(BLN30),.WL(WL42));
sram_cell_6t_5 inst_cell_42_31 (.BL(BL31),.BLN(BLN31),.WL(WL42));
sram_cell_6t_5 inst_cell_42_32 (.BL(BL32),.BLN(BLN32),.WL(WL42));
sram_cell_6t_5 inst_cell_42_33 (.BL(BL33),.BLN(BLN33),.WL(WL42));
sram_cell_6t_5 inst_cell_42_34 (.BL(BL34),.BLN(BLN34),.WL(WL42));
sram_cell_6t_5 inst_cell_42_35 (.BL(BL35),.BLN(BLN35),.WL(WL42));
sram_cell_6t_5 inst_cell_42_36 (.BL(BL36),.BLN(BLN36),.WL(WL42));
sram_cell_6t_5 inst_cell_42_37 (.BL(BL37),.BLN(BLN37),.WL(WL42));
sram_cell_6t_5 inst_cell_42_38 (.BL(BL38),.BLN(BLN38),.WL(WL42));
sram_cell_6t_5 inst_cell_42_39 (.BL(BL39),.BLN(BLN39),.WL(WL42));
sram_cell_6t_5 inst_cell_42_40 (.BL(BL40),.BLN(BLN40),.WL(WL42));
sram_cell_6t_5 inst_cell_42_41 (.BL(BL41),.BLN(BLN41),.WL(WL42));
sram_cell_6t_5 inst_cell_42_42 (.BL(BL42),.BLN(BLN42),.WL(WL42));
sram_cell_6t_5 inst_cell_42_43 (.BL(BL43),.BLN(BLN43),.WL(WL42));
sram_cell_6t_5 inst_cell_42_44 (.BL(BL44),.BLN(BLN44),.WL(WL42));
sram_cell_6t_5 inst_cell_42_45 (.BL(BL45),.BLN(BLN45),.WL(WL42));
sram_cell_6t_5 inst_cell_42_46 (.BL(BL46),.BLN(BLN46),.WL(WL42));
sram_cell_6t_5 inst_cell_42_47 (.BL(BL47),.BLN(BLN47),.WL(WL42));
sram_cell_6t_5 inst_cell_42_48 (.BL(BL48),.BLN(BLN48),.WL(WL42));
sram_cell_6t_5 inst_cell_42_49 (.BL(BL49),.BLN(BLN49),.WL(WL42));
sram_cell_6t_5 inst_cell_42_50 (.BL(BL50),.BLN(BLN50),.WL(WL42));
sram_cell_6t_5 inst_cell_42_51 (.BL(BL51),.BLN(BLN51),.WL(WL42));
sram_cell_6t_5 inst_cell_42_52 (.BL(BL52),.BLN(BLN52),.WL(WL42));
sram_cell_6t_5 inst_cell_42_53 (.BL(BL53),.BLN(BLN53),.WL(WL42));
sram_cell_6t_5 inst_cell_42_54 (.BL(BL54),.BLN(BLN54),.WL(WL42));
sram_cell_6t_5 inst_cell_42_55 (.BL(BL55),.BLN(BLN55),.WL(WL42));
sram_cell_6t_5 inst_cell_42_56 (.BL(BL56),.BLN(BLN56),.WL(WL42));
sram_cell_6t_5 inst_cell_42_57 (.BL(BL57),.BLN(BLN57),.WL(WL42));
sram_cell_6t_5 inst_cell_42_58 (.BL(BL58),.BLN(BLN58),.WL(WL42));
sram_cell_6t_5 inst_cell_42_59 (.BL(BL59),.BLN(BLN59),.WL(WL42));
sram_cell_6t_5 inst_cell_42_60 (.BL(BL60),.BLN(BLN60),.WL(WL42));
sram_cell_6t_5 inst_cell_42_61 (.BL(BL61),.BLN(BLN61),.WL(WL42));
sram_cell_6t_5 inst_cell_42_62 (.BL(BL62),.BLN(BLN62),.WL(WL42));
sram_cell_6t_5 inst_cell_42_63 (.BL(BL63),.BLN(BLN63),.WL(WL42));
sram_cell_6t_5 inst_cell_42_64 (.BL(BL64),.BLN(BLN64),.WL(WL42));
sram_cell_6t_5 inst_cell_42_65 (.BL(BL65),.BLN(BLN65),.WL(WL42));
sram_cell_6t_5 inst_cell_42_66 (.BL(BL66),.BLN(BLN66),.WL(WL42));
sram_cell_6t_5 inst_cell_42_67 (.BL(BL67),.BLN(BLN67),.WL(WL42));
sram_cell_6t_5 inst_cell_42_68 (.BL(BL68),.BLN(BLN68),.WL(WL42));
sram_cell_6t_5 inst_cell_42_69 (.BL(BL69),.BLN(BLN69),.WL(WL42));
sram_cell_6t_5 inst_cell_42_70 (.BL(BL70),.BLN(BLN70),.WL(WL42));
sram_cell_6t_5 inst_cell_42_71 (.BL(BL71),.BLN(BLN71),.WL(WL42));
sram_cell_6t_5 inst_cell_42_72 (.BL(BL72),.BLN(BLN72),.WL(WL42));
sram_cell_6t_5 inst_cell_42_73 (.BL(BL73),.BLN(BLN73),.WL(WL42));
sram_cell_6t_5 inst_cell_42_74 (.BL(BL74),.BLN(BLN74),.WL(WL42));
sram_cell_6t_5 inst_cell_42_75 (.BL(BL75),.BLN(BLN75),.WL(WL42));
sram_cell_6t_5 inst_cell_42_76 (.BL(BL76),.BLN(BLN76),.WL(WL42));
sram_cell_6t_5 inst_cell_42_77 (.BL(BL77),.BLN(BLN77),.WL(WL42));
sram_cell_6t_5 inst_cell_42_78 (.BL(BL78),.BLN(BLN78),.WL(WL42));
sram_cell_6t_5 inst_cell_42_79 (.BL(BL79),.BLN(BLN79),.WL(WL42));
sram_cell_6t_5 inst_cell_42_80 (.BL(BL80),.BLN(BLN80),.WL(WL42));
sram_cell_6t_5 inst_cell_42_81 (.BL(BL81),.BLN(BLN81),.WL(WL42));
sram_cell_6t_5 inst_cell_42_82 (.BL(BL82),.BLN(BLN82),.WL(WL42));
sram_cell_6t_5 inst_cell_42_83 (.BL(BL83),.BLN(BLN83),.WL(WL42));
sram_cell_6t_5 inst_cell_42_84 (.BL(BL84),.BLN(BLN84),.WL(WL42));
sram_cell_6t_5 inst_cell_42_85 (.BL(BL85),.BLN(BLN85),.WL(WL42));
sram_cell_6t_5 inst_cell_42_86 (.BL(BL86),.BLN(BLN86),.WL(WL42));
sram_cell_6t_5 inst_cell_42_87 (.BL(BL87),.BLN(BLN87),.WL(WL42));
sram_cell_6t_5 inst_cell_42_88 (.BL(BL88),.BLN(BLN88),.WL(WL42));
sram_cell_6t_5 inst_cell_42_89 (.BL(BL89),.BLN(BLN89),.WL(WL42));
sram_cell_6t_5 inst_cell_42_90 (.BL(BL90),.BLN(BLN90),.WL(WL42));
sram_cell_6t_5 inst_cell_42_91 (.BL(BL91),.BLN(BLN91),.WL(WL42));
sram_cell_6t_5 inst_cell_42_92 (.BL(BL92),.BLN(BLN92),.WL(WL42));
sram_cell_6t_5 inst_cell_42_93 (.BL(BL93),.BLN(BLN93),.WL(WL42));
sram_cell_6t_5 inst_cell_42_94 (.BL(BL94),.BLN(BLN94),.WL(WL42));
sram_cell_6t_5 inst_cell_42_95 (.BL(BL95),.BLN(BLN95),.WL(WL42));
sram_cell_6t_5 inst_cell_42_96 (.BL(BL96),.BLN(BLN96),.WL(WL42));
sram_cell_6t_5 inst_cell_42_97 (.BL(BL97),.BLN(BLN97),.WL(WL42));
sram_cell_6t_5 inst_cell_42_98 (.BL(BL98),.BLN(BLN98),.WL(WL42));
sram_cell_6t_5 inst_cell_42_99 (.BL(BL99),.BLN(BLN99),.WL(WL42));
sram_cell_6t_5 inst_cell_42_100 (.BL(BL100),.BLN(BLN100),.WL(WL42));
sram_cell_6t_5 inst_cell_42_101 (.BL(BL101),.BLN(BLN101),.WL(WL42));
sram_cell_6t_5 inst_cell_42_102 (.BL(BL102),.BLN(BLN102),.WL(WL42));
sram_cell_6t_5 inst_cell_42_103 (.BL(BL103),.BLN(BLN103),.WL(WL42));
sram_cell_6t_5 inst_cell_42_104 (.BL(BL104),.BLN(BLN104),.WL(WL42));
sram_cell_6t_5 inst_cell_42_105 (.BL(BL105),.BLN(BLN105),.WL(WL42));
sram_cell_6t_5 inst_cell_42_106 (.BL(BL106),.BLN(BLN106),.WL(WL42));
sram_cell_6t_5 inst_cell_42_107 (.BL(BL107),.BLN(BLN107),.WL(WL42));
sram_cell_6t_5 inst_cell_42_108 (.BL(BL108),.BLN(BLN108),.WL(WL42));
sram_cell_6t_5 inst_cell_42_109 (.BL(BL109),.BLN(BLN109),.WL(WL42));
sram_cell_6t_5 inst_cell_42_110 (.BL(BL110),.BLN(BLN110),.WL(WL42));
sram_cell_6t_5 inst_cell_42_111 (.BL(BL111),.BLN(BLN111),.WL(WL42));
sram_cell_6t_5 inst_cell_42_112 (.BL(BL112),.BLN(BLN112),.WL(WL42));
sram_cell_6t_5 inst_cell_42_113 (.BL(BL113),.BLN(BLN113),.WL(WL42));
sram_cell_6t_5 inst_cell_42_114 (.BL(BL114),.BLN(BLN114),.WL(WL42));
sram_cell_6t_5 inst_cell_42_115 (.BL(BL115),.BLN(BLN115),.WL(WL42));
sram_cell_6t_5 inst_cell_42_116 (.BL(BL116),.BLN(BLN116),.WL(WL42));
sram_cell_6t_5 inst_cell_42_117 (.BL(BL117),.BLN(BLN117),.WL(WL42));
sram_cell_6t_5 inst_cell_42_118 (.BL(BL118),.BLN(BLN118),.WL(WL42));
sram_cell_6t_5 inst_cell_42_119 (.BL(BL119),.BLN(BLN119),.WL(WL42));
sram_cell_6t_5 inst_cell_42_120 (.BL(BL120),.BLN(BLN120),.WL(WL42));
sram_cell_6t_5 inst_cell_42_121 (.BL(BL121),.BLN(BLN121),.WL(WL42));
sram_cell_6t_5 inst_cell_42_122 (.BL(BL122),.BLN(BLN122),.WL(WL42));
sram_cell_6t_5 inst_cell_42_123 (.BL(BL123),.BLN(BLN123),.WL(WL42));
sram_cell_6t_5 inst_cell_42_124 (.BL(BL124),.BLN(BLN124),.WL(WL42));
sram_cell_6t_5 inst_cell_42_125 (.BL(BL125),.BLN(BLN125),.WL(WL42));
sram_cell_6t_5 inst_cell_42_126 (.BL(BL126),.BLN(BLN126),.WL(WL42));
sram_cell_6t_5 inst_cell_42_127 (.BL(BL127),.BLN(BLN127),.WL(WL42));
sram_cell_6t_5 inst_cell_43_0 (.BL(BL0),.BLN(BLN0),.WL(WL43));
sram_cell_6t_5 inst_cell_43_1 (.BL(BL1),.BLN(BLN1),.WL(WL43));
sram_cell_6t_5 inst_cell_43_2 (.BL(BL2),.BLN(BLN2),.WL(WL43));
sram_cell_6t_5 inst_cell_43_3 (.BL(BL3),.BLN(BLN3),.WL(WL43));
sram_cell_6t_5 inst_cell_43_4 (.BL(BL4),.BLN(BLN4),.WL(WL43));
sram_cell_6t_5 inst_cell_43_5 (.BL(BL5),.BLN(BLN5),.WL(WL43));
sram_cell_6t_5 inst_cell_43_6 (.BL(BL6),.BLN(BLN6),.WL(WL43));
sram_cell_6t_5 inst_cell_43_7 (.BL(BL7),.BLN(BLN7),.WL(WL43));
sram_cell_6t_5 inst_cell_43_8 (.BL(BL8),.BLN(BLN8),.WL(WL43));
sram_cell_6t_5 inst_cell_43_9 (.BL(BL9),.BLN(BLN9),.WL(WL43));
sram_cell_6t_5 inst_cell_43_10 (.BL(BL10),.BLN(BLN10),.WL(WL43));
sram_cell_6t_5 inst_cell_43_11 (.BL(BL11),.BLN(BLN11),.WL(WL43));
sram_cell_6t_5 inst_cell_43_12 (.BL(BL12),.BLN(BLN12),.WL(WL43));
sram_cell_6t_5 inst_cell_43_13 (.BL(BL13),.BLN(BLN13),.WL(WL43));
sram_cell_6t_5 inst_cell_43_14 (.BL(BL14),.BLN(BLN14),.WL(WL43));
sram_cell_6t_5 inst_cell_43_15 (.BL(BL15),.BLN(BLN15),.WL(WL43));
sram_cell_6t_5 inst_cell_43_16 (.BL(BL16),.BLN(BLN16),.WL(WL43));
sram_cell_6t_5 inst_cell_43_17 (.BL(BL17),.BLN(BLN17),.WL(WL43));
sram_cell_6t_5 inst_cell_43_18 (.BL(BL18),.BLN(BLN18),.WL(WL43));
sram_cell_6t_5 inst_cell_43_19 (.BL(BL19),.BLN(BLN19),.WL(WL43));
sram_cell_6t_5 inst_cell_43_20 (.BL(BL20),.BLN(BLN20),.WL(WL43));
sram_cell_6t_5 inst_cell_43_21 (.BL(BL21),.BLN(BLN21),.WL(WL43));
sram_cell_6t_5 inst_cell_43_22 (.BL(BL22),.BLN(BLN22),.WL(WL43));
sram_cell_6t_5 inst_cell_43_23 (.BL(BL23),.BLN(BLN23),.WL(WL43));
sram_cell_6t_5 inst_cell_43_24 (.BL(BL24),.BLN(BLN24),.WL(WL43));
sram_cell_6t_5 inst_cell_43_25 (.BL(BL25),.BLN(BLN25),.WL(WL43));
sram_cell_6t_5 inst_cell_43_26 (.BL(BL26),.BLN(BLN26),.WL(WL43));
sram_cell_6t_5 inst_cell_43_27 (.BL(BL27),.BLN(BLN27),.WL(WL43));
sram_cell_6t_5 inst_cell_43_28 (.BL(BL28),.BLN(BLN28),.WL(WL43));
sram_cell_6t_5 inst_cell_43_29 (.BL(BL29),.BLN(BLN29),.WL(WL43));
sram_cell_6t_5 inst_cell_43_30 (.BL(BL30),.BLN(BLN30),.WL(WL43));
sram_cell_6t_5 inst_cell_43_31 (.BL(BL31),.BLN(BLN31),.WL(WL43));
sram_cell_6t_5 inst_cell_43_32 (.BL(BL32),.BLN(BLN32),.WL(WL43));
sram_cell_6t_5 inst_cell_43_33 (.BL(BL33),.BLN(BLN33),.WL(WL43));
sram_cell_6t_5 inst_cell_43_34 (.BL(BL34),.BLN(BLN34),.WL(WL43));
sram_cell_6t_5 inst_cell_43_35 (.BL(BL35),.BLN(BLN35),.WL(WL43));
sram_cell_6t_5 inst_cell_43_36 (.BL(BL36),.BLN(BLN36),.WL(WL43));
sram_cell_6t_5 inst_cell_43_37 (.BL(BL37),.BLN(BLN37),.WL(WL43));
sram_cell_6t_5 inst_cell_43_38 (.BL(BL38),.BLN(BLN38),.WL(WL43));
sram_cell_6t_5 inst_cell_43_39 (.BL(BL39),.BLN(BLN39),.WL(WL43));
sram_cell_6t_5 inst_cell_43_40 (.BL(BL40),.BLN(BLN40),.WL(WL43));
sram_cell_6t_5 inst_cell_43_41 (.BL(BL41),.BLN(BLN41),.WL(WL43));
sram_cell_6t_5 inst_cell_43_42 (.BL(BL42),.BLN(BLN42),.WL(WL43));
sram_cell_6t_5 inst_cell_43_43 (.BL(BL43),.BLN(BLN43),.WL(WL43));
sram_cell_6t_5 inst_cell_43_44 (.BL(BL44),.BLN(BLN44),.WL(WL43));
sram_cell_6t_5 inst_cell_43_45 (.BL(BL45),.BLN(BLN45),.WL(WL43));
sram_cell_6t_5 inst_cell_43_46 (.BL(BL46),.BLN(BLN46),.WL(WL43));
sram_cell_6t_5 inst_cell_43_47 (.BL(BL47),.BLN(BLN47),.WL(WL43));
sram_cell_6t_5 inst_cell_43_48 (.BL(BL48),.BLN(BLN48),.WL(WL43));
sram_cell_6t_5 inst_cell_43_49 (.BL(BL49),.BLN(BLN49),.WL(WL43));
sram_cell_6t_5 inst_cell_43_50 (.BL(BL50),.BLN(BLN50),.WL(WL43));
sram_cell_6t_5 inst_cell_43_51 (.BL(BL51),.BLN(BLN51),.WL(WL43));
sram_cell_6t_5 inst_cell_43_52 (.BL(BL52),.BLN(BLN52),.WL(WL43));
sram_cell_6t_5 inst_cell_43_53 (.BL(BL53),.BLN(BLN53),.WL(WL43));
sram_cell_6t_5 inst_cell_43_54 (.BL(BL54),.BLN(BLN54),.WL(WL43));
sram_cell_6t_5 inst_cell_43_55 (.BL(BL55),.BLN(BLN55),.WL(WL43));
sram_cell_6t_5 inst_cell_43_56 (.BL(BL56),.BLN(BLN56),.WL(WL43));
sram_cell_6t_5 inst_cell_43_57 (.BL(BL57),.BLN(BLN57),.WL(WL43));
sram_cell_6t_5 inst_cell_43_58 (.BL(BL58),.BLN(BLN58),.WL(WL43));
sram_cell_6t_5 inst_cell_43_59 (.BL(BL59),.BLN(BLN59),.WL(WL43));
sram_cell_6t_5 inst_cell_43_60 (.BL(BL60),.BLN(BLN60),.WL(WL43));
sram_cell_6t_5 inst_cell_43_61 (.BL(BL61),.BLN(BLN61),.WL(WL43));
sram_cell_6t_5 inst_cell_43_62 (.BL(BL62),.BLN(BLN62),.WL(WL43));
sram_cell_6t_5 inst_cell_43_63 (.BL(BL63),.BLN(BLN63),.WL(WL43));
sram_cell_6t_5 inst_cell_43_64 (.BL(BL64),.BLN(BLN64),.WL(WL43));
sram_cell_6t_5 inst_cell_43_65 (.BL(BL65),.BLN(BLN65),.WL(WL43));
sram_cell_6t_5 inst_cell_43_66 (.BL(BL66),.BLN(BLN66),.WL(WL43));
sram_cell_6t_5 inst_cell_43_67 (.BL(BL67),.BLN(BLN67),.WL(WL43));
sram_cell_6t_5 inst_cell_43_68 (.BL(BL68),.BLN(BLN68),.WL(WL43));
sram_cell_6t_5 inst_cell_43_69 (.BL(BL69),.BLN(BLN69),.WL(WL43));
sram_cell_6t_5 inst_cell_43_70 (.BL(BL70),.BLN(BLN70),.WL(WL43));
sram_cell_6t_5 inst_cell_43_71 (.BL(BL71),.BLN(BLN71),.WL(WL43));
sram_cell_6t_5 inst_cell_43_72 (.BL(BL72),.BLN(BLN72),.WL(WL43));
sram_cell_6t_5 inst_cell_43_73 (.BL(BL73),.BLN(BLN73),.WL(WL43));
sram_cell_6t_5 inst_cell_43_74 (.BL(BL74),.BLN(BLN74),.WL(WL43));
sram_cell_6t_5 inst_cell_43_75 (.BL(BL75),.BLN(BLN75),.WL(WL43));
sram_cell_6t_5 inst_cell_43_76 (.BL(BL76),.BLN(BLN76),.WL(WL43));
sram_cell_6t_5 inst_cell_43_77 (.BL(BL77),.BLN(BLN77),.WL(WL43));
sram_cell_6t_5 inst_cell_43_78 (.BL(BL78),.BLN(BLN78),.WL(WL43));
sram_cell_6t_5 inst_cell_43_79 (.BL(BL79),.BLN(BLN79),.WL(WL43));
sram_cell_6t_5 inst_cell_43_80 (.BL(BL80),.BLN(BLN80),.WL(WL43));
sram_cell_6t_5 inst_cell_43_81 (.BL(BL81),.BLN(BLN81),.WL(WL43));
sram_cell_6t_5 inst_cell_43_82 (.BL(BL82),.BLN(BLN82),.WL(WL43));
sram_cell_6t_5 inst_cell_43_83 (.BL(BL83),.BLN(BLN83),.WL(WL43));
sram_cell_6t_5 inst_cell_43_84 (.BL(BL84),.BLN(BLN84),.WL(WL43));
sram_cell_6t_5 inst_cell_43_85 (.BL(BL85),.BLN(BLN85),.WL(WL43));
sram_cell_6t_5 inst_cell_43_86 (.BL(BL86),.BLN(BLN86),.WL(WL43));
sram_cell_6t_5 inst_cell_43_87 (.BL(BL87),.BLN(BLN87),.WL(WL43));
sram_cell_6t_5 inst_cell_43_88 (.BL(BL88),.BLN(BLN88),.WL(WL43));
sram_cell_6t_5 inst_cell_43_89 (.BL(BL89),.BLN(BLN89),.WL(WL43));
sram_cell_6t_5 inst_cell_43_90 (.BL(BL90),.BLN(BLN90),.WL(WL43));
sram_cell_6t_5 inst_cell_43_91 (.BL(BL91),.BLN(BLN91),.WL(WL43));
sram_cell_6t_5 inst_cell_43_92 (.BL(BL92),.BLN(BLN92),.WL(WL43));
sram_cell_6t_5 inst_cell_43_93 (.BL(BL93),.BLN(BLN93),.WL(WL43));
sram_cell_6t_5 inst_cell_43_94 (.BL(BL94),.BLN(BLN94),.WL(WL43));
sram_cell_6t_5 inst_cell_43_95 (.BL(BL95),.BLN(BLN95),.WL(WL43));
sram_cell_6t_5 inst_cell_43_96 (.BL(BL96),.BLN(BLN96),.WL(WL43));
sram_cell_6t_5 inst_cell_43_97 (.BL(BL97),.BLN(BLN97),.WL(WL43));
sram_cell_6t_5 inst_cell_43_98 (.BL(BL98),.BLN(BLN98),.WL(WL43));
sram_cell_6t_5 inst_cell_43_99 (.BL(BL99),.BLN(BLN99),.WL(WL43));
sram_cell_6t_5 inst_cell_43_100 (.BL(BL100),.BLN(BLN100),.WL(WL43));
sram_cell_6t_5 inst_cell_43_101 (.BL(BL101),.BLN(BLN101),.WL(WL43));
sram_cell_6t_5 inst_cell_43_102 (.BL(BL102),.BLN(BLN102),.WL(WL43));
sram_cell_6t_5 inst_cell_43_103 (.BL(BL103),.BLN(BLN103),.WL(WL43));
sram_cell_6t_5 inst_cell_43_104 (.BL(BL104),.BLN(BLN104),.WL(WL43));
sram_cell_6t_5 inst_cell_43_105 (.BL(BL105),.BLN(BLN105),.WL(WL43));
sram_cell_6t_5 inst_cell_43_106 (.BL(BL106),.BLN(BLN106),.WL(WL43));
sram_cell_6t_5 inst_cell_43_107 (.BL(BL107),.BLN(BLN107),.WL(WL43));
sram_cell_6t_5 inst_cell_43_108 (.BL(BL108),.BLN(BLN108),.WL(WL43));
sram_cell_6t_5 inst_cell_43_109 (.BL(BL109),.BLN(BLN109),.WL(WL43));
sram_cell_6t_5 inst_cell_43_110 (.BL(BL110),.BLN(BLN110),.WL(WL43));
sram_cell_6t_5 inst_cell_43_111 (.BL(BL111),.BLN(BLN111),.WL(WL43));
sram_cell_6t_5 inst_cell_43_112 (.BL(BL112),.BLN(BLN112),.WL(WL43));
sram_cell_6t_5 inst_cell_43_113 (.BL(BL113),.BLN(BLN113),.WL(WL43));
sram_cell_6t_5 inst_cell_43_114 (.BL(BL114),.BLN(BLN114),.WL(WL43));
sram_cell_6t_5 inst_cell_43_115 (.BL(BL115),.BLN(BLN115),.WL(WL43));
sram_cell_6t_5 inst_cell_43_116 (.BL(BL116),.BLN(BLN116),.WL(WL43));
sram_cell_6t_5 inst_cell_43_117 (.BL(BL117),.BLN(BLN117),.WL(WL43));
sram_cell_6t_5 inst_cell_43_118 (.BL(BL118),.BLN(BLN118),.WL(WL43));
sram_cell_6t_5 inst_cell_43_119 (.BL(BL119),.BLN(BLN119),.WL(WL43));
sram_cell_6t_5 inst_cell_43_120 (.BL(BL120),.BLN(BLN120),.WL(WL43));
sram_cell_6t_5 inst_cell_43_121 (.BL(BL121),.BLN(BLN121),.WL(WL43));
sram_cell_6t_5 inst_cell_43_122 (.BL(BL122),.BLN(BLN122),.WL(WL43));
sram_cell_6t_5 inst_cell_43_123 (.BL(BL123),.BLN(BLN123),.WL(WL43));
sram_cell_6t_5 inst_cell_43_124 (.BL(BL124),.BLN(BLN124),.WL(WL43));
sram_cell_6t_5 inst_cell_43_125 (.BL(BL125),.BLN(BLN125),.WL(WL43));
sram_cell_6t_5 inst_cell_43_126 (.BL(BL126),.BLN(BLN126),.WL(WL43));
sram_cell_6t_5 inst_cell_43_127 (.BL(BL127),.BLN(BLN127),.WL(WL43));
sram_cell_6t_5 inst_cell_44_0 (.BL(BL0),.BLN(BLN0),.WL(WL44));
sram_cell_6t_5 inst_cell_44_1 (.BL(BL1),.BLN(BLN1),.WL(WL44));
sram_cell_6t_5 inst_cell_44_2 (.BL(BL2),.BLN(BLN2),.WL(WL44));
sram_cell_6t_5 inst_cell_44_3 (.BL(BL3),.BLN(BLN3),.WL(WL44));
sram_cell_6t_5 inst_cell_44_4 (.BL(BL4),.BLN(BLN4),.WL(WL44));
sram_cell_6t_5 inst_cell_44_5 (.BL(BL5),.BLN(BLN5),.WL(WL44));
sram_cell_6t_5 inst_cell_44_6 (.BL(BL6),.BLN(BLN6),.WL(WL44));
sram_cell_6t_5 inst_cell_44_7 (.BL(BL7),.BLN(BLN7),.WL(WL44));
sram_cell_6t_5 inst_cell_44_8 (.BL(BL8),.BLN(BLN8),.WL(WL44));
sram_cell_6t_5 inst_cell_44_9 (.BL(BL9),.BLN(BLN9),.WL(WL44));
sram_cell_6t_5 inst_cell_44_10 (.BL(BL10),.BLN(BLN10),.WL(WL44));
sram_cell_6t_5 inst_cell_44_11 (.BL(BL11),.BLN(BLN11),.WL(WL44));
sram_cell_6t_5 inst_cell_44_12 (.BL(BL12),.BLN(BLN12),.WL(WL44));
sram_cell_6t_5 inst_cell_44_13 (.BL(BL13),.BLN(BLN13),.WL(WL44));
sram_cell_6t_5 inst_cell_44_14 (.BL(BL14),.BLN(BLN14),.WL(WL44));
sram_cell_6t_5 inst_cell_44_15 (.BL(BL15),.BLN(BLN15),.WL(WL44));
sram_cell_6t_5 inst_cell_44_16 (.BL(BL16),.BLN(BLN16),.WL(WL44));
sram_cell_6t_5 inst_cell_44_17 (.BL(BL17),.BLN(BLN17),.WL(WL44));
sram_cell_6t_5 inst_cell_44_18 (.BL(BL18),.BLN(BLN18),.WL(WL44));
sram_cell_6t_5 inst_cell_44_19 (.BL(BL19),.BLN(BLN19),.WL(WL44));
sram_cell_6t_5 inst_cell_44_20 (.BL(BL20),.BLN(BLN20),.WL(WL44));
sram_cell_6t_5 inst_cell_44_21 (.BL(BL21),.BLN(BLN21),.WL(WL44));
sram_cell_6t_5 inst_cell_44_22 (.BL(BL22),.BLN(BLN22),.WL(WL44));
sram_cell_6t_5 inst_cell_44_23 (.BL(BL23),.BLN(BLN23),.WL(WL44));
sram_cell_6t_5 inst_cell_44_24 (.BL(BL24),.BLN(BLN24),.WL(WL44));
sram_cell_6t_5 inst_cell_44_25 (.BL(BL25),.BLN(BLN25),.WL(WL44));
sram_cell_6t_5 inst_cell_44_26 (.BL(BL26),.BLN(BLN26),.WL(WL44));
sram_cell_6t_5 inst_cell_44_27 (.BL(BL27),.BLN(BLN27),.WL(WL44));
sram_cell_6t_5 inst_cell_44_28 (.BL(BL28),.BLN(BLN28),.WL(WL44));
sram_cell_6t_5 inst_cell_44_29 (.BL(BL29),.BLN(BLN29),.WL(WL44));
sram_cell_6t_5 inst_cell_44_30 (.BL(BL30),.BLN(BLN30),.WL(WL44));
sram_cell_6t_5 inst_cell_44_31 (.BL(BL31),.BLN(BLN31),.WL(WL44));
sram_cell_6t_5 inst_cell_44_32 (.BL(BL32),.BLN(BLN32),.WL(WL44));
sram_cell_6t_5 inst_cell_44_33 (.BL(BL33),.BLN(BLN33),.WL(WL44));
sram_cell_6t_5 inst_cell_44_34 (.BL(BL34),.BLN(BLN34),.WL(WL44));
sram_cell_6t_5 inst_cell_44_35 (.BL(BL35),.BLN(BLN35),.WL(WL44));
sram_cell_6t_5 inst_cell_44_36 (.BL(BL36),.BLN(BLN36),.WL(WL44));
sram_cell_6t_5 inst_cell_44_37 (.BL(BL37),.BLN(BLN37),.WL(WL44));
sram_cell_6t_5 inst_cell_44_38 (.BL(BL38),.BLN(BLN38),.WL(WL44));
sram_cell_6t_5 inst_cell_44_39 (.BL(BL39),.BLN(BLN39),.WL(WL44));
sram_cell_6t_5 inst_cell_44_40 (.BL(BL40),.BLN(BLN40),.WL(WL44));
sram_cell_6t_5 inst_cell_44_41 (.BL(BL41),.BLN(BLN41),.WL(WL44));
sram_cell_6t_5 inst_cell_44_42 (.BL(BL42),.BLN(BLN42),.WL(WL44));
sram_cell_6t_5 inst_cell_44_43 (.BL(BL43),.BLN(BLN43),.WL(WL44));
sram_cell_6t_5 inst_cell_44_44 (.BL(BL44),.BLN(BLN44),.WL(WL44));
sram_cell_6t_5 inst_cell_44_45 (.BL(BL45),.BLN(BLN45),.WL(WL44));
sram_cell_6t_5 inst_cell_44_46 (.BL(BL46),.BLN(BLN46),.WL(WL44));
sram_cell_6t_5 inst_cell_44_47 (.BL(BL47),.BLN(BLN47),.WL(WL44));
sram_cell_6t_5 inst_cell_44_48 (.BL(BL48),.BLN(BLN48),.WL(WL44));
sram_cell_6t_5 inst_cell_44_49 (.BL(BL49),.BLN(BLN49),.WL(WL44));
sram_cell_6t_5 inst_cell_44_50 (.BL(BL50),.BLN(BLN50),.WL(WL44));
sram_cell_6t_5 inst_cell_44_51 (.BL(BL51),.BLN(BLN51),.WL(WL44));
sram_cell_6t_5 inst_cell_44_52 (.BL(BL52),.BLN(BLN52),.WL(WL44));
sram_cell_6t_5 inst_cell_44_53 (.BL(BL53),.BLN(BLN53),.WL(WL44));
sram_cell_6t_5 inst_cell_44_54 (.BL(BL54),.BLN(BLN54),.WL(WL44));
sram_cell_6t_5 inst_cell_44_55 (.BL(BL55),.BLN(BLN55),.WL(WL44));
sram_cell_6t_5 inst_cell_44_56 (.BL(BL56),.BLN(BLN56),.WL(WL44));
sram_cell_6t_5 inst_cell_44_57 (.BL(BL57),.BLN(BLN57),.WL(WL44));
sram_cell_6t_5 inst_cell_44_58 (.BL(BL58),.BLN(BLN58),.WL(WL44));
sram_cell_6t_5 inst_cell_44_59 (.BL(BL59),.BLN(BLN59),.WL(WL44));
sram_cell_6t_5 inst_cell_44_60 (.BL(BL60),.BLN(BLN60),.WL(WL44));
sram_cell_6t_5 inst_cell_44_61 (.BL(BL61),.BLN(BLN61),.WL(WL44));
sram_cell_6t_5 inst_cell_44_62 (.BL(BL62),.BLN(BLN62),.WL(WL44));
sram_cell_6t_5 inst_cell_44_63 (.BL(BL63),.BLN(BLN63),.WL(WL44));
sram_cell_6t_5 inst_cell_44_64 (.BL(BL64),.BLN(BLN64),.WL(WL44));
sram_cell_6t_5 inst_cell_44_65 (.BL(BL65),.BLN(BLN65),.WL(WL44));
sram_cell_6t_5 inst_cell_44_66 (.BL(BL66),.BLN(BLN66),.WL(WL44));
sram_cell_6t_5 inst_cell_44_67 (.BL(BL67),.BLN(BLN67),.WL(WL44));
sram_cell_6t_5 inst_cell_44_68 (.BL(BL68),.BLN(BLN68),.WL(WL44));
sram_cell_6t_5 inst_cell_44_69 (.BL(BL69),.BLN(BLN69),.WL(WL44));
sram_cell_6t_5 inst_cell_44_70 (.BL(BL70),.BLN(BLN70),.WL(WL44));
sram_cell_6t_5 inst_cell_44_71 (.BL(BL71),.BLN(BLN71),.WL(WL44));
sram_cell_6t_5 inst_cell_44_72 (.BL(BL72),.BLN(BLN72),.WL(WL44));
sram_cell_6t_5 inst_cell_44_73 (.BL(BL73),.BLN(BLN73),.WL(WL44));
sram_cell_6t_5 inst_cell_44_74 (.BL(BL74),.BLN(BLN74),.WL(WL44));
sram_cell_6t_5 inst_cell_44_75 (.BL(BL75),.BLN(BLN75),.WL(WL44));
sram_cell_6t_5 inst_cell_44_76 (.BL(BL76),.BLN(BLN76),.WL(WL44));
sram_cell_6t_5 inst_cell_44_77 (.BL(BL77),.BLN(BLN77),.WL(WL44));
sram_cell_6t_5 inst_cell_44_78 (.BL(BL78),.BLN(BLN78),.WL(WL44));
sram_cell_6t_5 inst_cell_44_79 (.BL(BL79),.BLN(BLN79),.WL(WL44));
sram_cell_6t_5 inst_cell_44_80 (.BL(BL80),.BLN(BLN80),.WL(WL44));
sram_cell_6t_5 inst_cell_44_81 (.BL(BL81),.BLN(BLN81),.WL(WL44));
sram_cell_6t_5 inst_cell_44_82 (.BL(BL82),.BLN(BLN82),.WL(WL44));
sram_cell_6t_5 inst_cell_44_83 (.BL(BL83),.BLN(BLN83),.WL(WL44));
sram_cell_6t_5 inst_cell_44_84 (.BL(BL84),.BLN(BLN84),.WL(WL44));
sram_cell_6t_5 inst_cell_44_85 (.BL(BL85),.BLN(BLN85),.WL(WL44));
sram_cell_6t_5 inst_cell_44_86 (.BL(BL86),.BLN(BLN86),.WL(WL44));
sram_cell_6t_5 inst_cell_44_87 (.BL(BL87),.BLN(BLN87),.WL(WL44));
sram_cell_6t_5 inst_cell_44_88 (.BL(BL88),.BLN(BLN88),.WL(WL44));
sram_cell_6t_5 inst_cell_44_89 (.BL(BL89),.BLN(BLN89),.WL(WL44));
sram_cell_6t_5 inst_cell_44_90 (.BL(BL90),.BLN(BLN90),.WL(WL44));
sram_cell_6t_5 inst_cell_44_91 (.BL(BL91),.BLN(BLN91),.WL(WL44));
sram_cell_6t_5 inst_cell_44_92 (.BL(BL92),.BLN(BLN92),.WL(WL44));
sram_cell_6t_5 inst_cell_44_93 (.BL(BL93),.BLN(BLN93),.WL(WL44));
sram_cell_6t_5 inst_cell_44_94 (.BL(BL94),.BLN(BLN94),.WL(WL44));
sram_cell_6t_5 inst_cell_44_95 (.BL(BL95),.BLN(BLN95),.WL(WL44));
sram_cell_6t_5 inst_cell_44_96 (.BL(BL96),.BLN(BLN96),.WL(WL44));
sram_cell_6t_5 inst_cell_44_97 (.BL(BL97),.BLN(BLN97),.WL(WL44));
sram_cell_6t_5 inst_cell_44_98 (.BL(BL98),.BLN(BLN98),.WL(WL44));
sram_cell_6t_5 inst_cell_44_99 (.BL(BL99),.BLN(BLN99),.WL(WL44));
sram_cell_6t_5 inst_cell_44_100 (.BL(BL100),.BLN(BLN100),.WL(WL44));
sram_cell_6t_5 inst_cell_44_101 (.BL(BL101),.BLN(BLN101),.WL(WL44));
sram_cell_6t_5 inst_cell_44_102 (.BL(BL102),.BLN(BLN102),.WL(WL44));
sram_cell_6t_5 inst_cell_44_103 (.BL(BL103),.BLN(BLN103),.WL(WL44));
sram_cell_6t_5 inst_cell_44_104 (.BL(BL104),.BLN(BLN104),.WL(WL44));
sram_cell_6t_5 inst_cell_44_105 (.BL(BL105),.BLN(BLN105),.WL(WL44));
sram_cell_6t_5 inst_cell_44_106 (.BL(BL106),.BLN(BLN106),.WL(WL44));
sram_cell_6t_5 inst_cell_44_107 (.BL(BL107),.BLN(BLN107),.WL(WL44));
sram_cell_6t_5 inst_cell_44_108 (.BL(BL108),.BLN(BLN108),.WL(WL44));
sram_cell_6t_5 inst_cell_44_109 (.BL(BL109),.BLN(BLN109),.WL(WL44));
sram_cell_6t_5 inst_cell_44_110 (.BL(BL110),.BLN(BLN110),.WL(WL44));
sram_cell_6t_5 inst_cell_44_111 (.BL(BL111),.BLN(BLN111),.WL(WL44));
sram_cell_6t_5 inst_cell_44_112 (.BL(BL112),.BLN(BLN112),.WL(WL44));
sram_cell_6t_5 inst_cell_44_113 (.BL(BL113),.BLN(BLN113),.WL(WL44));
sram_cell_6t_5 inst_cell_44_114 (.BL(BL114),.BLN(BLN114),.WL(WL44));
sram_cell_6t_5 inst_cell_44_115 (.BL(BL115),.BLN(BLN115),.WL(WL44));
sram_cell_6t_5 inst_cell_44_116 (.BL(BL116),.BLN(BLN116),.WL(WL44));
sram_cell_6t_5 inst_cell_44_117 (.BL(BL117),.BLN(BLN117),.WL(WL44));
sram_cell_6t_5 inst_cell_44_118 (.BL(BL118),.BLN(BLN118),.WL(WL44));
sram_cell_6t_5 inst_cell_44_119 (.BL(BL119),.BLN(BLN119),.WL(WL44));
sram_cell_6t_5 inst_cell_44_120 (.BL(BL120),.BLN(BLN120),.WL(WL44));
sram_cell_6t_5 inst_cell_44_121 (.BL(BL121),.BLN(BLN121),.WL(WL44));
sram_cell_6t_5 inst_cell_44_122 (.BL(BL122),.BLN(BLN122),.WL(WL44));
sram_cell_6t_5 inst_cell_44_123 (.BL(BL123),.BLN(BLN123),.WL(WL44));
sram_cell_6t_5 inst_cell_44_124 (.BL(BL124),.BLN(BLN124),.WL(WL44));
sram_cell_6t_5 inst_cell_44_125 (.BL(BL125),.BLN(BLN125),.WL(WL44));
sram_cell_6t_5 inst_cell_44_126 (.BL(BL126),.BLN(BLN126),.WL(WL44));
sram_cell_6t_5 inst_cell_44_127 (.BL(BL127),.BLN(BLN127),.WL(WL44));
sram_cell_6t_5 inst_cell_45_0 (.BL(BL0),.BLN(BLN0),.WL(WL45));
sram_cell_6t_5 inst_cell_45_1 (.BL(BL1),.BLN(BLN1),.WL(WL45));
sram_cell_6t_5 inst_cell_45_2 (.BL(BL2),.BLN(BLN2),.WL(WL45));
sram_cell_6t_5 inst_cell_45_3 (.BL(BL3),.BLN(BLN3),.WL(WL45));
sram_cell_6t_5 inst_cell_45_4 (.BL(BL4),.BLN(BLN4),.WL(WL45));
sram_cell_6t_5 inst_cell_45_5 (.BL(BL5),.BLN(BLN5),.WL(WL45));
sram_cell_6t_5 inst_cell_45_6 (.BL(BL6),.BLN(BLN6),.WL(WL45));
sram_cell_6t_5 inst_cell_45_7 (.BL(BL7),.BLN(BLN7),.WL(WL45));
sram_cell_6t_5 inst_cell_45_8 (.BL(BL8),.BLN(BLN8),.WL(WL45));
sram_cell_6t_5 inst_cell_45_9 (.BL(BL9),.BLN(BLN9),.WL(WL45));
sram_cell_6t_5 inst_cell_45_10 (.BL(BL10),.BLN(BLN10),.WL(WL45));
sram_cell_6t_5 inst_cell_45_11 (.BL(BL11),.BLN(BLN11),.WL(WL45));
sram_cell_6t_5 inst_cell_45_12 (.BL(BL12),.BLN(BLN12),.WL(WL45));
sram_cell_6t_5 inst_cell_45_13 (.BL(BL13),.BLN(BLN13),.WL(WL45));
sram_cell_6t_5 inst_cell_45_14 (.BL(BL14),.BLN(BLN14),.WL(WL45));
sram_cell_6t_5 inst_cell_45_15 (.BL(BL15),.BLN(BLN15),.WL(WL45));
sram_cell_6t_5 inst_cell_45_16 (.BL(BL16),.BLN(BLN16),.WL(WL45));
sram_cell_6t_5 inst_cell_45_17 (.BL(BL17),.BLN(BLN17),.WL(WL45));
sram_cell_6t_5 inst_cell_45_18 (.BL(BL18),.BLN(BLN18),.WL(WL45));
sram_cell_6t_5 inst_cell_45_19 (.BL(BL19),.BLN(BLN19),.WL(WL45));
sram_cell_6t_5 inst_cell_45_20 (.BL(BL20),.BLN(BLN20),.WL(WL45));
sram_cell_6t_5 inst_cell_45_21 (.BL(BL21),.BLN(BLN21),.WL(WL45));
sram_cell_6t_5 inst_cell_45_22 (.BL(BL22),.BLN(BLN22),.WL(WL45));
sram_cell_6t_5 inst_cell_45_23 (.BL(BL23),.BLN(BLN23),.WL(WL45));
sram_cell_6t_5 inst_cell_45_24 (.BL(BL24),.BLN(BLN24),.WL(WL45));
sram_cell_6t_5 inst_cell_45_25 (.BL(BL25),.BLN(BLN25),.WL(WL45));
sram_cell_6t_5 inst_cell_45_26 (.BL(BL26),.BLN(BLN26),.WL(WL45));
sram_cell_6t_5 inst_cell_45_27 (.BL(BL27),.BLN(BLN27),.WL(WL45));
sram_cell_6t_5 inst_cell_45_28 (.BL(BL28),.BLN(BLN28),.WL(WL45));
sram_cell_6t_5 inst_cell_45_29 (.BL(BL29),.BLN(BLN29),.WL(WL45));
sram_cell_6t_5 inst_cell_45_30 (.BL(BL30),.BLN(BLN30),.WL(WL45));
sram_cell_6t_5 inst_cell_45_31 (.BL(BL31),.BLN(BLN31),.WL(WL45));
sram_cell_6t_5 inst_cell_45_32 (.BL(BL32),.BLN(BLN32),.WL(WL45));
sram_cell_6t_5 inst_cell_45_33 (.BL(BL33),.BLN(BLN33),.WL(WL45));
sram_cell_6t_5 inst_cell_45_34 (.BL(BL34),.BLN(BLN34),.WL(WL45));
sram_cell_6t_5 inst_cell_45_35 (.BL(BL35),.BLN(BLN35),.WL(WL45));
sram_cell_6t_5 inst_cell_45_36 (.BL(BL36),.BLN(BLN36),.WL(WL45));
sram_cell_6t_5 inst_cell_45_37 (.BL(BL37),.BLN(BLN37),.WL(WL45));
sram_cell_6t_5 inst_cell_45_38 (.BL(BL38),.BLN(BLN38),.WL(WL45));
sram_cell_6t_5 inst_cell_45_39 (.BL(BL39),.BLN(BLN39),.WL(WL45));
sram_cell_6t_5 inst_cell_45_40 (.BL(BL40),.BLN(BLN40),.WL(WL45));
sram_cell_6t_5 inst_cell_45_41 (.BL(BL41),.BLN(BLN41),.WL(WL45));
sram_cell_6t_5 inst_cell_45_42 (.BL(BL42),.BLN(BLN42),.WL(WL45));
sram_cell_6t_5 inst_cell_45_43 (.BL(BL43),.BLN(BLN43),.WL(WL45));
sram_cell_6t_5 inst_cell_45_44 (.BL(BL44),.BLN(BLN44),.WL(WL45));
sram_cell_6t_5 inst_cell_45_45 (.BL(BL45),.BLN(BLN45),.WL(WL45));
sram_cell_6t_5 inst_cell_45_46 (.BL(BL46),.BLN(BLN46),.WL(WL45));
sram_cell_6t_5 inst_cell_45_47 (.BL(BL47),.BLN(BLN47),.WL(WL45));
sram_cell_6t_5 inst_cell_45_48 (.BL(BL48),.BLN(BLN48),.WL(WL45));
sram_cell_6t_5 inst_cell_45_49 (.BL(BL49),.BLN(BLN49),.WL(WL45));
sram_cell_6t_5 inst_cell_45_50 (.BL(BL50),.BLN(BLN50),.WL(WL45));
sram_cell_6t_5 inst_cell_45_51 (.BL(BL51),.BLN(BLN51),.WL(WL45));
sram_cell_6t_5 inst_cell_45_52 (.BL(BL52),.BLN(BLN52),.WL(WL45));
sram_cell_6t_5 inst_cell_45_53 (.BL(BL53),.BLN(BLN53),.WL(WL45));
sram_cell_6t_5 inst_cell_45_54 (.BL(BL54),.BLN(BLN54),.WL(WL45));
sram_cell_6t_5 inst_cell_45_55 (.BL(BL55),.BLN(BLN55),.WL(WL45));
sram_cell_6t_5 inst_cell_45_56 (.BL(BL56),.BLN(BLN56),.WL(WL45));
sram_cell_6t_5 inst_cell_45_57 (.BL(BL57),.BLN(BLN57),.WL(WL45));
sram_cell_6t_5 inst_cell_45_58 (.BL(BL58),.BLN(BLN58),.WL(WL45));
sram_cell_6t_5 inst_cell_45_59 (.BL(BL59),.BLN(BLN59),.WL(WL45));
sram_cell_6t_5 inst_cell_45_60 (.BL(BL60),.BLN(BLN60),.WL(WL45));
sram_cell_6t_5 inst_cell_45_61 (.BL(BL61),.BLN(BLN61),.WL(WL45));
sram_cell_6t_5 inst_cell_45_62 (.BL(BL62),.BLN(BLN62),.WL(WL45));
sram_cell_6t_5 inst_cell_45_63 (.BL(BL63),.BLN(BLN63),.WL(WL45));
sram_cell_6t_5 inst_cell_45_64 (.BL(BL64),.BLN(BLN64),.WL(WL45));
sram_cell_6t_5 inst_cell_45_65 (.BL(BL65),.BLN(BLN65),.WL(WL45));
sram_cell_6t_5 inst_cell_45_66 (.BL(BL66),.BLN(BLN66),.WL(WL45));
sram_cell_6t_5 inst_cell_45_67 (.BL(BL67),.BLN(BLN67),.WL(WL45));
sram_cell_6t_5 inst_cell_45_68 (.BL(BL68),.BLN(BLN68),.WL(WL45));
sram_cell_6t_5 inst_cell_45_69 (.BL(BL69),.BLN(BLN69),.WL(WL45));
sram_cell_6t_5 inst_cell_45_70 (.BL(BL70),.BLN(BLN70),.WL(WL45));
sram_cell_6t_5 inst_cell_45_71 (.BL(BL71),.BLN(BLN71),.WL(WL45));
sram_cell_6t_5 inst_cell_45_72 (.BL(BL72),.BLN(BLN72),.WL(WL45));
sram_cell_6t_5 inst_cell_45_73 (.BL(BL73),.BLN(BLN73),.WL(WL45));
sram_cell_6t_5 inst_cell_45_74 (.BL(BL74),.BLN(BLN74),.WL(WL45));
sram_cell_6t_5 inst_cell_45_75 (.BL(BL75),.BLN(BLN75),.WL(WL45));
sram_cell_6t_5 inst_cell_45_76 (.BL(BL76),.BLN(BLN76),.WL(WL45));
sram_cell_6t_5 inst_cell_45_77 (.BL(BL77),.BLN(BLN77),.WL(WL45));
sram_cell_6t_5 inst_cell_45_78 (.BL(BL78),.BLN(BLN78),.WL(WL45));
sram_cell_6t_5 inst_cell_45_79 (.BL(BL79),.BLN(BLN79),.WL(WL45));
sram_cell_6t_5 inst_cell_45_80 (.BL(BL80),.BLN(BLN80),.WL(WL45));
sram_cell_6t_5 inst_cell_45_81 (.BL(BL81),.BLN(BLN81),.WL(WL45));
sram_cell_6t_5 inst_cell_45_82 (.BL(BL82),.BLN(BLN82),.WL(WL45));
sram_cell_6t_5 inst_cell_45_83 (.BL(BL83),.BLN(BLN83),.WL(WL45));
sram_cell_6t_5 inst_cell_45_84 (.BL(BL84),.BLN(BLN84),.WL(WL45));
sram_cell_6t_5 inst_cell_45_85 (.BL(BL85),.BLN(BLN85),.WL(WL45));
sram_cell_6t_5 inst_cell_45_86 (.BL(BL86),.BLN(BLN86),.WL(WL45));
sram_cell_6t_5 inst_cell_45_87 (.BL(BL87),.BLN(BLN87),.WL(WL45));
sram_cell_6t_5 inst_cell_45_88 (.BL(BL88),.BLN(BLN88),.WL(WL45));
sram_cell_6t_5 inst_cell_45_89 (.BL(BL89),.BLN(BLN89),.WL(WL45));
sram_cell_6t_5 inst_cell_45_90 (.BL(BL90),.BLN(BLN90),.WL(WL45));
sram_cell_6t_5 inst_cell_45_91 (.BL(BL91),.BLN(BLN91),.WL(WL45));
sram_cell_6t_5 inst_cell_45_92 (.BL(BL92),.BLN(BLN92),.WL(WL45));
sram_cell_6t_5 inst_cell_45_93 (.BL(BL93),.BLN(BLN93),.WL(WL45));
sram_cell_6t_5 inst_cell_45_94 (.BL(BL94),.BLN(BLN94),.WL(WL45));
sram_cell_6t_5 inst_cell_45_95 (.BL(BL95),.BLN(BLN95),.WL(WL45));
sram_cell_6t_5 inst_cell_45_96 (.BL(BL96),.BLN(BLN96),.WL(WL45));
sram_cell_6t_5 inst_cell_45_97 (.BL(BL97),.BLN(BLN97),.WL(WL45));
sram_cell_6t_5 inst_cell_45_98 (.BL(BL98),.BLN(BLN98),.WL(WL45));
sram_cell_6t_5 inst_cell_45_99 (.BL(BL99),.BLN(BLN99),.WL(WL45));
sram_cell_6t_5 inst_cell_45_100 (.BL(BL100),.BLN(BLN100),.WL(WL45));
sram_cell_6t_5 inst_cell_45_101 (.BL(BL101),.BLN(BLN101),.WL(WL45));
sram_cell_6t_5 inst_cell_45_102 (.BL(BL102),.BLN(BLN102),.WL(WL45));
sram_cell_6t_5 inst_cell_45_103 (.BL(BL103),.BLN(BLN103),.WL(WL45));
sram_cell_6t_5 inst_cell_45_104 (.BL(BL104),.BLN(BLN104),.WL(WL45));
sram_cell_6t_5 inst_cell_45_105 (.BL(BL105),.BLN(BLN105),.WL(WL45));
sram_cell_6t_5 inst_cell_45_106 (.BL(BL106),.BLN(BLN106),.WL(WL45));
sram_cell_6t_5 inst_cell_45_107 (.BL(BL107),.BLN(BLN107),.WL(WL45));
sram_cell_6t_5 inst_cell_45_108 (.BL(BL108),.BLN(BLN108),.WL(WL45));
sram_cell_6t_5 inst_cell_45_109 (.BL(BL109),.BLN(BLN109),.WL(WL45));
sram_cell_6t_5 inst_cell_45_110 (.BL(BL110),.BLN(BLN110),.WL(WL45));
sram_cell_6t_5 inst_cell_45_111 (.BL(BL111),.BLN(BLN111),.WL(WL45));
sram_cell_6t_5 inst_cell_45_112 (.BL(BL112),.BLN(BLN112),.WL(WL45));
sram_cell_6t_5 inst_cell_45_113 (.BL(BL113),.BLN(BLN113),.WL(WL45));
sram_cell_6t_5 inst_cell_45_114 (.BL(BL114),.BLN(BLN114),.WL(WL45));
sram_cell_6t_5 inst_cell_45_115 (.BL(BL115),.BLN(BLN115),.WL(WL45));
sram_cell_6t_5 inst_cell_45_116 (.BL(BL116),.BLN(BLN116),.WL(WL45));
sram_cell_6t_5 inst_cell_45_117 (.BL(BL117),.BLN(BLN117),.WL(WL45));
sram_cell_6t_5 inst_cell_45_118 (.BL(BL118),.BLN(BLN118),.WL(WL45));
sram_cell_6t_5 inst_cell_45_119 (.BL(BL119),.BLN(BLN119),.WL(WL45));
sram_cell_6t_5 inst_cell_45_120 (.BL(BL120),.BLN(BLN120),.WL(WL45));
sram_cell_6t_5 inst_cell_45_121 (.BL(BL121),.BLN(BLN121),.WL(WL45));
sram_cell_6t_5 inst_cell_45_122 (.BL(BL122),.BLN(BLN122),.WL(WL45));
sram_cell_6t_5 inst_cell_45_123 (.BL(BL123),.BLN(BLN123),.WL(WL45));
sram_cell_6t_5 inst_cell_45_124 (.BL(BL124),.BLN(BLN124),.WL(WL45));
sram_cell_6t_5 inst_cell_45_125 (.BL(BL125),.BLN(BLN125),.WL(WL45));
sram_cell_6t_5 inst_cell_45_126 (.BL(BL126),.BLN(BLN126),.WL(WL45));
sram_cell_6t_5 inst_cell_45_127 (.BL(BL127),.BLN(BLN127),.WL(WL45));
sram_cell_6t_5 inst_cell_46_0 (.BL(BL0),.BLN(BLN0),.WL(WL46));
sram_cell_6t_5 inst_cell_46_1 (.BL(BL1),.BLN(BLN1),.WL(WL46));
sram_cell_6t_5 inst_cell_46_2 (.BL(BL2),.BLN(BLN2),.WL(WL46));
sram_cell_6t_5 inst_cell_46_3 (.BL(BL3),.BLN(BLN3),.WL(WL46));
sram_cell_6t_5 inst_cell_46_4 (.BL(BL4),.BLN(BLN4),.WL(WL46));
sram_cell_6t_5 inst_cell_46_5 (.BL(BL5),.BLN(BLN5),.WL(WL46));
sram_cell_6t_5 inst_cell_46_6 (.BL(BL6),.BLN(BLN6),.WL(WL46));
sram_cell_6t_5 inst_cell_46_7 (.BL(BL7),.BLN(BLN7),.WL(WL46));
sram_cell_6t_5 inst_cell_46_8 (.BL(BL8),.BLN(BLN8),.WL(WL46));
sram_cell_6t_5 inst_cell_46_9 (.BL(BL9),.BLN(BLN9),.WL(WL46));
sram_cell_6t_5 inst_cell_46_10 (.BL(BL10),.BLN(BLN10),.WL(WL46));
sram_cell_6t_5 inst_cell_46_11 (.BL(BL11),.BLN(BLN11),.WL(WL46));
sram_cell_6t_5 inst_cell_46_12 (.BL(BL12),.BLN(BLN12),.WL(WL46));
sram_cell_6t_5 inst_cell_46_13 (.BL(BL13),.BLN(BLN13),.WL(WL46));
sram_cell_6t_5 inst_cell_46_14 (.BL(BL14),.BLN(BLN14),.WL(WL46));
sram_cell_6t_5 inst_cell_46_15 (.BL(BL15),.BLN(BLN15),.WL(WL46));
sram_cell_6t_5 inst_cell_46_16 (.BL(BL16),.BLN(BLN16),.WL(WL46));
sram_cell_6t_5 inst_cell_46_17 (.BL(BL17),.BLN(BLN17),.WL(WL46));
sram_cell_6t_5 inst_cell_46_18 (.BL(BL18),.BLN(BLN18),.WL(WL46));
sram_cell_6t_5 inst_cell_46_19 (.BL(BL19),.BLN(BLN19),.WL(WL46));
sram_cell_6t_5 inst_cell_46_20 (.BL(BL20),.BLN(BLN20),.WL(WL46));
sram_cell_6t_5 inst_cell_46_21 (.BL(BL21),.BLN(BLN21),.WL(WL46));
sram_cell_6t_5 inst_cell_46_22 (.BL(BL22),.BLN(BLN22),.WL(WL46));
sram_cell_6t_5 inst_cell_46_23 (.BL(BL23),.BLN(BLN23),.WL(WL46));
sram_cell_6t_5 inst_cell_46_24 (.BL(BL24),.BLN(BLN24),.WL(WL46));
sram_cell_6t_5 inst_cell_46_25 (.BL(BL25),.BLN(BLN25),.WL(WL46));
sram_cell_6t_5 inst_cell_46_26 (.BL(BL26),.BLN(BLN26),.WL(WL46));
sram_cell_6t_5 inst_cell_46_27 (.BL(BL27),.BLN(BLN27),.WL(WL46));
sram_cell_6t_5 inst_cell_46_28 (.BL(BL28),.BLN(BLN28),.WL(WL46));
sram_cell_6t_5 inst_cell_46_29 (.BL(BL29),.BLN(BLN29),.WL(WL46));
sram_cell_6t_5 inst_cell_46_30 (.BL(BL30),.BLN(BLN30),.WL(WL46));
sram_cell_6t_5 inst_cell_46_31 (.BL(BL31),.BLN(BLN31),.WL(WL46));
sram_cell_6t_5 inst_cell_46_32 (.BL(BL32),.BLN(BLN32),.WL(WL46));
sram_cell_6t_5 inst_cell_46_33 (.BL(BL33),.BLN(BLN33),.WL(WL46));
sram_cell_6t_5 inst_cell_46_34 (.BL(BL34),.BLN(BLN34),.WL(WL46));
sram_cell_6t_5 inst_cell_46_35 (.BL(BL35),.BLN(BLN35),.WL(WL46));
sram_cell_6t_5 inst_cell_46_36 (.BL(BL36),.BLN(BLN36),.WL(WL46));
sram_cell_6t_5 inst_cell_46_37 (.BL(BL37),.BLN(BLN37),.WL(WL46));
sram_cell_6t_5 inst_cell_46_38 (.BL(BL38),.BLN(BLN38),.WL(WL46));
sram_cell_6t_5 inst_cell_46_39 (.BL(BL39),.BLN(BLN39),.WL(WL46));
sram_cell_6t_5 inst_cell_46_40 (.BL(BL40),.BLN(BLN40),.WL(WL46));
sram_cell_6t_5 inst_cell_46_41 (.BL(BL41),.BLN(BLN41),.WL(WL46));
sram_cell_6t_5 inst_cell_46_42 (.BL(BL42),.BLN(BLN42),.WL(WL46));
sram_cell_6t_5 inst_cell_46_43 (.BL(BL43),.BLN(BLN43),.WL(WL46));
sram_cell_6t_5 inst_cell_46_44 (.BL(BL44),.BLN(BLN44),.WL(WL46));
sram_cell_6t_5 inst_cell_46_45 (.BL(BL45),.BLN(BLN45),.WL(WL46));
sram_cell_6t_5 inst_cell_46_46 (.BL(BL46),.BLN(BLN46),.WL(WL46));
sram_cell_6t_5 inst_cell_46_47 (.BL(BL47),.BLN(BLN47),.WL(WL46));
sram_cell_6t_5 inst_cell_46_48 (.BL(BL48),.BLN(BLN48),.WL(WL46));
sram_cell_6t_5 inst_cell_46_49 (.BL(BL49),.BLN(BLN49),.WL(WL46));
sram_cell_6t_5 inst_cell_46_50 (.BL(BL50),.BLN(BLN50),.WL(WL46));
sram_cell_6t_5 inst_cell_46_51 (.BL(BL51),.BLN(BLN51),.WL(WL46));
sram_cell_6t_5 inst_cell_46_52 (.BL(BL52),.BLN(BLN52),.WL(WL46));
sram_cell_6t_5 inst_cell_46_53 (.BL(BL53),.BLN(BLN53),.WL(WL46));
sram_cell_6t_5 inst_cell_46_54 (.BL(BL54),.BLN(BLN54),.WL(WL46));
sram_cell_6t_5 inst_cell_46_55 (.BL(BL55),.BLN(BLN55),.WL(WL46));
sram_cell_6t_5 inst_cell_46_56 (.BL(BL56),.BLN(BLN56),.WL(WL46));
sram_cell_6t_5 inst_cell_46_57 (.BL(BL57),.BLN(BLN57),.WL(WL46));
sram_cell_6t_5 inst_cell_46_58 (.BL(BL58),.BLN(BLN58),.WL(WL46));
sram_cell_6t_5 inst_cell_46_59 (.BL(BL59),.BLN(BLN59),.WL(WL46));
sram_cell_6t_5 inst_cell_46_60 (.BL(BL60),.BLN(BLN60),.WL(WL46));
sram_cell_6t_5 inst_cell_46_61 (.BL(BL61),.BLN(BLN61),.WL(WL46));
sram_cell_6t_5 inst_cell_46_62 (.BL(BL62),.BLN(BLN62),.WL(WL46));
sram_cell_6t_5 inst_cell_46_63 (.BL(BL63),.BLN(BLN63),.WL(WL46));
sram_cell_6t_5 inst_cell_46_64 (.BL(BL64),.BLN(BLN64),.WL(WL46));
sram_cell_6t_5 inst_cell_46_65 (.BL(BL65),.BLN(BLN65),.WL(WL46));
sram_cell_6t_5 inst_cell_46_66 (.BL(BL66),.BLN(BLN66),.WL(WL46));
sram_cell_6t_5 inst_cell_46_67 (.BL(BL67),.BLN(BLN67),.WL(WL46));
sram_cell_6t_5 inst_cell_46_68 (.BL(BL68),.BLN(BLN68),.WL(WL46));
sram_cell_6t_5 inst_cell_46_69 (.BL(BL69),.BLN(BLN69),.WL(WL46));
sram_cell_6t_5 inst_cell_46_70 (.BL(BL70),.BLN(BLN70),.WL(WL46));
sram_cell_6t_5 inst_cell_46_71 (.BL(BL71),.BLN(BLN71),.WL(WL46));
sram_cell_6t_5 inst_cell_46_72 (.BL(BL72),.BLN(BLN72),.WL(WL46));
sram_cell_6t_5 inst_cell_46_73 (.BL(BL73),.BLN(BLN73),.WL(WL46));
sram_cell_6t_5 inst_cell_46_74 (.BL(BL74),.BLN(BLN74),.WL(WL46));
sram_cell_6t_5 inst_cell_46_75 (.BL(BL75),.BLN(BLN75),.WL(WL46));
sram_cell_6t_5 inst_cell_46_76 (.BL(BL76),.BLN(BLN76),.WL(WL46));
sram_cell_6t_5 inst_cell_46_77 (.BL(BL77),.BLN(BLN77),.WL(WL46));
sram_cell_6t_5 inst_cell_46_78 (.BL(BL78),.BLN(BLN78),.WL(WL46));
sram_cell_6t_5 inst_cell_46_79 (.BL(BL79),.BLN(BLN79),.WL(WL46));
sram_cell_6t_5 inst_cell_46_80 (.BL(BL80),.BLN(BLN80),.WL(WL46));
sram_cell_6t_5 inst_cell_46_81 (.BL(BL81),.BLN(BLN81),.WL(WL46));
sram_cell_6t_5 inst_cell_46_82 (.BL(BL82),.BLN(BLN82),.WL(WL46));
sram_cell_6t_5 inst_cell_46_83 (.BL(BL83),.BLN(BLN83),.WL(WL46));
sram_cell_6t_5 inst_cell_46_84 (.BL(BL84),.BLN(BLN84),.WL(WL46));
sram_cell_6t_5 inst_cell_46_85 (.BL(BL85),.BLN(BLN85),.WL(WL46));
sram_cell_6t_5 inst_cell_46_86 (.BL(BL86),.BLN(BLN86),.WL(WL46));
sram_cell_6t_5 inst_cell_46_87 (.BL(BL87),.BLN(BLN87),.WL(WL46));
sram_cell_6t_5 inst_cell_46_88 (.BL(BL88),.BLN(BLN88),.WL(WL46));
sram_cell_6t_5 inst_cell_46_89 (.BL(BL89),.BLN(BLN89),.WL(WL46));
sram_cell_6t_5 inst_cell_46_90 (.BL(BL90),.BLN(BLN90),.WL(WL46));
sram_cell_6t_5 inst_cell_46_91 (.BL(BL91),.BLN(BLN91),.WL(WL46));
sram_cell_6t_5 inst_cell_46_92 (.BL(BL92),.BLN(BLN92),.WL(WL46));
sram_cell_6t_5 inst_cell_46_93 (.BL(BL93),.BLN(BLN93),.WL(WL46));
sram_cell_6t_5 inst_cell_46_94 (.BL(BL94),.BLN(BLN94),.WL(WL46));
sram_cell_6t_5 inst_cell_46_95 (.BL(BL95),.BLN(BLN95),.WL(WL46));
sram_cell_6t_5 inst_cell_46_96 (.BL(BL96),.BLN(BLN96),.WL(WL46));
sram_cell_6t_5 inst_cell_46_97 (.BL(BL97),.BLN(BLN97),.WL(WL46));
sram_cell_6t_5 inst_cell_46_98 (.BL(BL98),.BLN(BLN98),.WL(WL46));
sram_cell_6t_5 inst_cell_46_99 (.BL(BL99),.BLN(BLN99),.WL(WL46));
sram_cell_6t_5 inst_cell_46_100 (.BL(BL100),.BLN(BLN100),.WL(WL46));
sram_cell_6t_5 inst_cell_46_101 (.BL(BL101),.BLN(BLN101),.WL(WL46));
sram_cell_6t_5 inst_cell_46_102 (.BL(BL102),.BLN(BLN102),.WL(WL46));
sram_cell_6t_5 inst_cell_46_103 (.BL(BL103),.BLN(BLN103),.WL(WL46));
sram_cell_6t_5 inst_cell_46_104 (.BL(BL104),.BLN(BLN104),.WL(WL46));
sram_cell_6t_5 inst_cell_46_105 (.BL(BL105),.BLN(BLN105),.WL(WL46));
sram_cell_6t_5 inst_cell_46_106 (.BL(BL106),.BLN(BLN106),.WL(WL46));
sram_cell_6t_5 inst_cell_46_107 (.BL(BL107),.BLN(BLN107),.WL(WL46));
sram_cell_6t_5 inst_cell_46_108 (.BL(BL108),.BLN(BLN108),.WL(WL46));
sram_cell_6t_5 inst_cell_46_109 (.BL(BL109),.BLN(BLN109),.WL(WL46));
sram_cell_6t_5 inst_cell_46_110 (.BL(BL110),.BLN(BLN110),.WL(WL46));
sram_cell_6t_5 inst_cell_46_111 (.BL(BL111),.BLN(BLN111),.WL(WL46));
sram_cell_6t_5 inst_cell_46_112 (.BL(BL112),.BLN(BLN112),.WL(WL46));
sram_cell_6t_5 inst_cell_46_113 (.BL(BL113),.BLN(BLN113),.WL(WL46));
sram_cell_6t_5 inst_cell_46_114 (.BL(BL114),.BLN(BLN114),.WL(WL46));
sram_cell_6t_5 inst_cell_46_115 (.BL(BL115),.BLN(BLN115),.WL(WL46));
sram_cell_6t_5 inst_cell_46_116 (.BL(BL116),.BLN(BLN116),.WL(WL46));
sram_cell_6t_5 inst_cell_46_117 (.BL(BL117),.BLN(BLN117),.WL(WL46));
sram_cell_6t_5 inst_cell_46_118 (.BL(BL118),.BLN(BLN118),.WL(WL46));
sram_cell_6t_5 inst_cell_46_119 (.BL(BL119),.BLN(BLN119),.WL(WL46));
sram_cell_6t_5 inst_cell_46_120 (.BL(BL120),.BLN(BLN120),.WL(WL46));
sram_cell_6t_5 inst_cell_46_121 (.BL(BL121),.BLN(BLN121),.WL(WL46));
sram_cell_6t_5 inst_cell_46_122 (.BL(BL122),.BLN(BLN122),.WL(WL46));
sram_cell_6t_5 inst_cell_46_123 (.BL(BL123),.BLN(BLN123),.WL(WL46));
sram_cell_6t_5 inst_cell_46_124 (.BL(BL124),.BLN(BLN124),.WL(WL46));
sram_cell_6t_5 inst_cell_46_125 (.BL(BL125),.BLN(BLN125),.WL(WL46));
sram_cell_6t_5 inst_cell_46_126 (.BL(BL126),.BLN(BLN126),.WL(WL46));
sram_cell_6t_5 inst_cell_46_127 (.BL(BL127),.BLN(BLN127),.WL(WL46));
sram_cell_6t_5 inst_cell_47_0 (.BL(BL0),.BLN(BLN0),.WL(WL47));
sram_cell_6t_5 inst_cell_47_1 (.BL(BL1),.BLN(BLN1),.WL(WL47));
sram_cell_6t_5 inst_cell_47_2 (.BL(BL2),.BLN(BLN2),.WL(WL47));
sram_cell_6t_5 inst_cell_47_3 (.BL(BL3),.BLN(BLN3),.WL(WL47));
sram_cell_6t_5 inst_cell_47_4 (.BL(BL4),.BLN(BLN4),.WL(WL47));
sram_cell_6t_5 inst_cell_47_5 (.BL(BL5),.BLN(BLN5),.WL(WL47));
sram_cell_6t_5 inst_cell_47_6 (.BL(BL6),.BLN(BLN6),.WL(WL47));
sram_cell_6t_5 inst_cell_47_7 (.BL(BL7),.BLN(BLN7),.WL(WL47));
sram_cell_6t_5 inst_cell_47_8 (.BL(BL8),.BLN(BLN8),.WL(WL47));
sram_cell_6t_5 inst_cell_47_9 (.BL(BL9),.BLN(BLN9),.WL(WL47));
sram_cell_6t_5 inst_cell_47_10 (.BL(BL10),.BLN(BLN10),.WL(WL47));
sram_cell_6t_5 inst_cell_47_11 (.BL(BL11),.BLN(BLN11),.WL(WL47));
sram_cell_6t_5 inst_cell_47_12 (.BL(BL12),.BLN(BLN12),.WL(WL47));
sram_cell_6t_5 inst_cell_47_13 (.BL(BL13),.BLN(BLN13),.WL(WL47));
sram_cell_6t_5 inst_cell_47_14 (.BL(BL14),.BLN(BLN14),.WL(WL47));
sram_cell_6t_5 inst_cell_47_15 (.BL(BL15),.BLN(BLN15),.WL(WL47));
sram_cell_6t_5 inst_cell_47_16 (.BL(BL16),.BLN(BLN16),.WL(WL47));
sram_cell_6t_5 inst_cell_47_17 (.BL(BL17),.BLN(BLN17),.WL(WL47));
sram_cell_6t_5 inst_cell_47_18 (.BL(BL18),.BLN(BLN18),.WL(WL47));
sram_cell_6t_5 inst_cell_47_19 (.BL(BL19),.BLN(BLN19),.WL(WL47));
sram_cell_6t_5 inst_cell_47_20 (.BL(BL20),.BLN(BLN20),.WL(WL47));
sram_cell_6t_5 inst_cell_47_21 (.BL(BL21),.BLN(BLN21),.WL(WL47));
sram_cell_6t_5 inst_cell_47_22 (.BL(BL22),.BLN(BLN22),.WL(WL47));
sram_cell_6t_5 inst_cell_47_23 (.BL(BL23),.BLN(BLN23),.WL(WL47));
sram_cell_6t_5 inst_cell_47_24 (.BL(BL24),.BLN(BLN24),.WL(WL47));
sram_cell_6t_5 inst_cell_47_25 (.BL(BL25),.BLN(BLN25),.WL(WL47));
sram_cell_6t_5 inst_cell_47_26 (.BL(BL26),.BLN(BLN26),.WL(WL47));
sram_cell_6t_5 inst_cell_47_27 (.BL(BL27),.BLN(BLN27),.WL(WL47));
sram_cell_6t_5 inst_cell_47_28 (.BL(BL28),.BLN(BLN28),.WL(WL47));
sram_cell_6t_5 inst_cell_47_29 (.BL(BL29),.BLN(BLN29),.WL(WL47));
sram_cell_6t_5 inst_cell_47_30 (.BL(BL30),.BLN(BLN30),.WL(WL47));
sram_cell_6t_5 inst_cell_47_31 (.BL(BL31),.BLN(BLN31),.WL(WL47));
sram_cell_6t_5 inst_cell_47_32 (.BL(BL32),.BLN(BLN32),.WL(WL47));
sram_cell_6t_5 inst_cell_47_33 (.BL(BL33),.BLN(BLN33),.WL(WL47));
sram_cell_6t_5 inst_cell_47_34 (.BL(BL34),.BLN(BLN34),.WL(WL47));
sram_cell_6t_5 inst_cell_47_35 (.BL(BL35),.BLN(BLN35),.WL(WL47));
sram_cell_6t_5 inst_cell_47_36 (.BL(BL36),.BLN(BLN36),.WL(WL47));
sram_cell_6t_5 inst_cell_47_37 (.BL(BL37),.BLN(BLN37),.WL(WL47));
sram_cell_6t_5 inst_cell_47_38 (.BL(BL38),.BLN(BLN38),.WL(WL47));
sram_cell_6t_5 inst_cell_47_39 (.BL(BL39),.BLN(BLN39),.WL(WL47));
sram_cell_6t_5 inst_cell_47_40 (.BL(BL40),.BLN(BLN40),.WL(WL47));
sram_cell_6t_5 inst_cell_47_41 (.BL(BL41),.BLN(BLN41),.WL(WL47));
sram_cell_6t_5 inst_cell_47_42 (.BL(BL42),.BLN(BLN42),.WL(WL47));
sram_cell_6t_5 inst_cell_47_43 (.BL(BL43),.BLN(BLN43),.WL(WL47));
sram_cell_6t_5 inst_cell_47_44 (.BL(BL44),.BLN(BLN44),.WL(WL47));
sram_cell_6t_5 inst_cell_47_45 (.BL(BL45),.BLN(BLN45),.WL(WL47));
sram_cell_6t_5 inst_cell_47_46 (.BL(BL46),.BLN(BLN46),.WL(WL47));
sram_cell_6t_5 inst_cell_47_47 (.BL(BL47),.BLN(BLN47),.WL(WL47));
sram_cell_6t_5 inst_cell_47_48 (.BL(BL48),.BLN(BLN48),.WL(WL47));
sram_cell_6t_5 inst_cell_47_49 (.BL(BL49),.BLN(BLN49),.WL(WL47));
sram_cell_6t_5 inst_cell_47_50 (.BL(BL50),.BLN(BLN50),.WL(WL47));
sram_cell_6t_5 inst_cell_47_51 (.BL(BL51),.BLN(BLN51),.WL(WL47));
sram_cell_6t_5 inst_cell_47_52 (.BL(BL52),.BLN(BLN52),.WL(WL47));
sram_cell_6t_5 inst_cell_47_53 (.BL(BL53),.BLN(BLN53),.WL(WL47));
sram_cell_6t_5 inst_cell_47_54 (.BL(BL54),.BLN(BLN54),.WL(WL47));
sram_cell_6t_5 inst_cell_47_55 (.BL(BL55),.BLN(BLN55),.WL(WL47));
sram_cell_6t_5 inst_cell_47_56 (.BL(BL56),.BLN(BLN56),.WL(WL47));
sram_cell_6t_5 inst_cell_47_57 (.BL(BL57),.BLN(BLN57),.WL(WL47));
sram_cell_6t_5 inst_cell_47_58 (.BL(BL58),.BLN(BLN58),.WL(WL47));
sram_cell_6t_5 inst_cell_47_59 (.BL(BL59),.BLN(BLN59),.WL(WL47));
sram_cell_6t_5 inst_cell_47_60 (.BL(BL60),.BLN(BLN60),.WL(WL47));
sram_cell_6t_5 inst_cell_47_61 (.BL(BL61),.BLN(BLN61),.WL(WL47));
sram_cell_6t_5 inst_cell_47_62 (.BL(BL62),.BLN(BLN62),.WL(WL47));
sram_cell_6t_5 inst_cell_47_63 (.BL(BL63),.BLN(BLN63),.WL(WL47));
sram_cell_6t_5 inst_cell_47_64 (.BL(BL64),.BLN(BLN64),.WL(WL47));
sram_cell_6t_5 inst_cell_47_65 (.BL(BL65),.BLN(BLN65),.WL(WL47));
sram_cell_6t_5 inst_cell_47_66 (.BL(BL66),.BLN(BLN66),.WL(WL47));
sram_cell_6t_5 inst_cell_47_67 (.BL(BL67),.BLN(BLN67),.WL(WL47));
sram_cell_6t_5 inst_cell_47_68 (.BL(BL68),.BLN(BLN68),.WL(WL47));
sram_cell_6t_5 inst_cell_47_69 (.BL(BL69),.BLN(BLN69),.WL(WL47));
sram_cell_6t_5 inst_cell_47_70 (.BL(BL70),.BLN(BLN70),.WL(WL47));
sram_cell_6t_5 inst_cell_47_71 (.BL(BL71),.BLN(BLN71),.WL(WL47));
sram_cell_6t_5 inst_cell_47_72 (.BL(BL72),.BLN(BLN72),.WL(WL47));
sram_cell_6t_5 inst_cell_47_73 (.BL(BL73),.BLN(BLN73),.WL(WL47));
sram_cell_6t_5 inst_cell_47_74 (.BL(BL74),.BLN(BLN74),.WL(WL47));
sram_cell_6t_5 inst_cell_47_75 (.BL(BL75),.BLN(BLN75),.WL(WL47));
sram_cell_6t_5 inst_cell_47_76 (.BL(BL76),.BLN(BLN76),.WL(WL47));
sram_cell_6t_5 inst_cell_47_77 (.BL(BL77),.BLN(BLN77),.WL(WL47));
sram_cell_6t_5 inst_cell_47_78 (.BL(BL78),.BLN(BLN78),.WL(WL47));
sram_cell_6t_5 inst_cell_47_79 (.BL(BL79),.BLN(BLN79),.WL(WL47));
sram_cell_6t_5 inst_cell_47_80 (.BL(BL80),.BLN(BLN80),.WL(WL47));
sram_cell_6t_5 inst_cell_47_81 (.BL(BL81),.BLN(BLN81),.WL(WL47));
sram_cell_6t_5 inst_cell_47_82 (.BL(BL82),.BLN(BLN82),.WL(WL47));
sram_cell_6t_5 inst_cell_47_83 (.BL(BL83),.BLN(BLN83),.WL(WL47));
sram_cell_6t_5 inst_cell_47_84 (.BL(BL84),.BLN(BLN84),.WL(WL47));
sram_cell_6t_5 inst_cell_47_85 (.BL(BL85),.BLN(BLN85),.WL(WL47));
sram_cell_6t_5 inst_cell_47_86 (.BL(BL86),.BLN(BLN86),.WL(WL47));
sram_cell_6t_5 inst_cell_47_87 (.BL(BL87),.BLN(BLN87),.WL(WL47));
sram_cell_6t_5 inst_cell_47_88 (.BL(BL88),.BLN(BLN88),.WL(WL47));
sram_cell_6t_5 inst_cell_47_89 (.BL(BL89),.BLN(BLN89),.WL(WL47));
sram_cell_6t_5 inst_cell_47_90 (.BL(BL90),.BLN(BLN90),.WL(WL47));
sram_cell_6t_5 inst_cell_47_91 (.BL(BL91),.BLN(BLN91),.WL(WL47));
sram_cell_6t_5 inst_cell_47_92 (.BL(BL92),.BLN(BLN92),.WL(WL47));
sram_cell_6t_5 inst_cell_47_93 (.BL(BL93),.BLN(BLN93),.WL(WL47));
sram_cell_6t_5 inst_cell_47_94 (.BL(BL94),.BLN(BLN94),.WL(WL47));
sram_cell_6t_5 inst_cell_47_95 (.BL(BL95),.BLN(BLN95),.WL(WL47));
sram_cell_6t_5 inst_cell_47_96 (.BL(BL96),.BLN(BLN96),.WL(WL47));
sram_cell_6t_5 inst_cell_47_97 (.BL(BL97),.BLN(BLN97),.WL(WL47));
sram_cell_6t_5 inst_cell_47_98 (.BL(BL98),.BLN(BLN98),.WL(WL47));
sram_cell_6t_5 inst_cell_47_99 (.BL(BL99),.BLN(BLN99),.WL(WL47));
sram_cell_6t_5 inst_cell_47_100 (.BL(BL100),.BLN(BLN100),.WL(WL47));
sram_cell_6t_5 inst_cell_47_101 (.BL(BL101),.BLN(BLN101),.WL(WL47));
sram_cell_6t_5 inst_cell_47_102 (.BL(BL102),.BLN(BLN102),.WL(WL47));
sram_cell_6t_5 inst_cell_47_103 (.BL(BL103),.BLN(BLN103),.WL(WL47));
sram_cell_6t_5 inst_cell_47_104 (.BL(BL104),.BLN(BLN104),.WL(WL47));
sram_cell_6t_5 inst_cell_47_105 (.BL(BL105),.BLN(BLN105),.WL(WL47));
sram_cell_6t_5 inst_cell_47_106 (.BL(BL106),.BLN(BLN106),.WL(WL47));
sram_cell_6t_5 inst_cell_47_107 (.BL(BL107),.BLN(BLN107),.WL(WL47));
sram_cell_6t_5 inst_cell_47_108 (.BL(BL108),.BLN(BLN108),.WL(WL47));
sram_cell_6t_5 inst_cell_47_109 (.BL(BL109),.BLN(BLN109),.WL(WL47));
sram_cell_6t_5 inst_cell_47_110 (.BL(BL110),.BLN(BLN110),.WL(WL47));
sram_cell_6t_5 inst_cell_47_111 (.BL(BL111),.BLN(BLN111),.WL(WL47));
sram_cell_6t_5 inst_cell_47_112 (.BL(BL112),.BLN(BLN112),.WL(WL47));
sram_cell_6t_5 inst_cell_47_113 (.BL(BL113),.BLN(BLN113),.WL(WL47));
sram_cell_6t_5 inst_cell_47_114 (.BL(BL114),.BLN(BLN114),.WL(WL47));
sram_cell_6t_5 inst_cell_47_115 (.BL(BL115),.BLN(BLN115),.WL(WL47));
sram_cell_6t_5 inst_cell_47_116 (.BL(BL116),.BLN(BLN116),.WL(WL47));
sram_cell_6t_5 inst_cell_47_117 (.BL(BL117),.BLN(BLN117),.WL(WL47));
sram_cell_6t_5 inst_cell_47_118 (.BL(BL118),.BLN(BLN118),.WL(WL47));
sram_cell_6t_5 inst_cell_47_119 (.BL(BL119),.BLN(BLN119),.WL(WL47));
sram_cell_6t_5 inst_cell_47_120 (.BL(BL120),.BLN(BLN120),.WL(WL47));
sram_cell_6t_5 inst_cell_47_121 (.BL(BL121),.BLN(BLN121),.WL(WL47));
sram_cell_6t_5 inst_cell_47_122 (.BL(BL122),.BLN(BLN122),.WL(WL47));
sram_cell_6t_5 inst_cell_47_123 (.BL(BL123),.BLN(BLN123),.WL(WL47));
sram_cell_6t_5 inst_cell_47_124 (.BL(BL124),.BLN(BLN124),.WL(WL47));
sram_cell_6t_5 inst_cell_47_125 (.BL(BL125),.BLN(BLN125),.WL(WL47));
sram_cell_6t_5 inst_cell_47_126 (.BL(BL126),.BLN(BLN126),.WL(WL47));
sram_cell_6t_5 inst_cell_47_127 (.BL(BL127),.BLN(BLN127),.WL(WL47));
sram_cell_6t_5 inst_cell_48_0 (.BL(BL0),.BLN(BLN0),.WL(WL48));
sram_cell_6t_5 inst_cell_48_1 (.BL(BL1),.BLN(BLN1),.WL(WL48));
sram_cell_6t_5 inst_cell_48_2 (.BL(BL2),.BLN(BLN2),.WL(WL48));
sram_cell_6t_5 inst_cell_48_3 (.BL(BL3),.BLN(BLN3),.WL(WL48));
sram_cell_6t_5 inst_cell_48_4 (.BL(BL4),.BLN(BLN4),.WL(WL48));
sram_cell_6t_5 inst_cell_48_5 (.BL(BL5),.BLN(BLN5),.WL(WL48));
sram_cell_6t_5 inst_cell_48_6 (.BL(BL6),.BLN(BLN6),.WL(WL48));
sram_cell_6t_5 inst_cell_48_7 (.BL(BL7),.BLN(BLN7),.WL(WL48));
sram_cell_6t_5 inst_cell_48_8 (.BL(BL8),.BLN(BLN8),.WL(WL48));
sram_cell_6t_5 inst_cell_48_9 (.BL(BL9),.BLN(BLN9),.WL(WL48));
sram_cell_6t_5 inst_cell_48_10 (.BL(BL10),.BLN(BLN10),.WL(WL48));
sram_cell_6t_5 inst_cell_48_11 (.BL(BL11),.BLN(BLN11),.WL(WL48));
sram_cell_6t_5 inst_cell_48_12 (.BL(BL12),.BLN(BLN12),.WL(WL48));
sram_cell_6t_5 inst_cell_48_13 (.BL(BL13),.BLN(BLN13),.WL(WL48));
sram_cell_6t_5 inst_cell_48_14 (.BL(BL14),.BLN(BLN14),.WL(WL48));
sram_cell_6t_5 inst_cell_48_15 (.BL(BL15),.BLN(BLN15),.WL(WL48));
sram_cell_6t_5 inst_cell_48_16 (.BL(BL16),.BLN(BLN16),.WL(WL48));
sram_cell_6t_5 inst_cell_48_17 (.BL(BL17),.BLN(BLN17),.WL(WL48));
sram_cell_6t_5 inst_cell_48_18 (.BL(BL18),.BLN(BLN18),.WL(WL48));
sram_cell_6t_5 inst_cell_48_19 (.BL(BL19),.BLN(BLN19),.WL(WL48));
sram_cell_6t_5 inst_cell_48_20 (.BL(BL20),.BLN(BLN20),.WL(WL48));
sram_cell_6t_5 inst_cell_48_21 (.BL(BL21),.BLN(BLN21),.WL(WL48));
sram_cell_6t_5 inst_cell_48_22 (.BL(BL22),.BLN(BLN22),.WL(WL48));
sram_cell_6t_5 inst_cell_48_23 (.BL(BL23),.BLN(BLN23),.WL(WL48));
sram_cell_6t_5 inst_cell_48_24 (.BL(BL24),.BLN(BLN24),.WL(WL48));
sram_cell_6t_5 inst_cell_48_25 (.BL(BL25),.BLN(BLN25),.WL(WL48));
sram_cell_6t_5 inst_cell_48_26 (.BL(BL26),.BLN(BLN26),.WL(WL48));
sram_cell_6t_5 inst_cell_48_27 (.BL(BL27),.BLN(BLN27),.WL(WL48));
sram_cell_6t_5 inst_cell_48_28 (.BL(BL28),.BLN(BLN28),.WL(WL48));
sram_cell_6t_5 inst_cell_48_29 (.BL(BL29),.BLN(BLN29),.WL(WL48));
sram_cell_6t_5 inst_cell_48_30 (.BL(BL30),.BLN(BLN30),.WL(WL48));
sram_cell_6t_5 inst_cell_48_31 (.BL(BL31),.BLN(BLN31),.WL(WL48));
sram_cell_6t_5 inst_cell_48_32 (.BL(BL32),.BLN(BLN32),.WL(WL48));
sram_cell_6t_5 inst_cell_48_33 (.BL(BL33),.BLN(BLN33),.WL(WL48));
sram_cell_6t_5 inst_cell_48_34 (.BL(BL34),.BLN(BLN34),.WL(WL48));
sram_cell_6t_5 inst_cell_48_35 (.BL(BL35),.BLN(BLN35),.WL(WL48));
sram_cell_6t_5 inst_cell_48_36 (.BL(BL36),.BLN(BLN36),.WL(WL48));
sram_cell_6t_5 inst_cell_48_37 (.BL(BL37),.BLN(BLN37),.WL(WL48));
sram_cell_6t_5 inst_cell_48_38 (.BL(BL38),.BLN(BLN38),.WL(WL48));
sram_cell_6t_5 inst_cell_48_39 (.BL(BL39),.BLN(BLN39),.WL(WL48));
sram_cell_6t_5 inst_cell_48_40 (.BL(BL40),.BLN(BLN40),.WL(WL48));
sram_cell_6t_5 inst_cell_48_41 (.BL(BL41),.BLN(BLN41),.WL(WL48));
sram_cell_6t_5 inst_cell_48_42 (.BL(BL42),.BLN(BLN42),.WL(WL48));
sram_cell_6t_5 inst_cell_48_43 (.BL(BL43),.BLN(BLN43),.WL(WL48));
sram_cell_6t_5 inst_cell_48_44 (.BL(BL44),.BLN(BLN44),.WL(WL48));
sram_cell_6t_5 inst_cell_48_45 (.BL(BL45),.BLN(BLN45),.WL(WL48));
sram_cell_6t_5 inst_cell_48_46 (.BL(BL46),.BLN(BLN46),.WL(WL48));
sram_cell_6t_5 inst_cell_48_47 (.BL(BL47),.BLN(BLN47),.WL(WL48));
sram_cell_6t_5 inst_cell_48_48 (.BL(BL48),.BLN(BLN48),.WL(WL48));
sram_cell_6t_5 inst_cell_48_49 (.BL(BL49),.BLN(BLN49),.WL(WL48));
sram_cell_6t_5 inst_cell_48_50 (.BL(BL50),.BLN(BLN50),.WL(WL48));
sram_cell_6t_5 inst_cell_48_51 (.BL(BL51),.BLN(BLN51),.WL(WL48));
sram_cell_6t_5 inst_cell_48_52 (.BL(BL52),.BLN(BLN52),.WL(WL48));
sram_cell_6t_5 inst_cell_48_53 (.BL(BL53),.BLN(BLN53),.WL(WL48));
sram_cell_6t_5 inst_cell_48_54 (.BL(BL54),.BLN(BLN54),.WL(WL48));
sram_cell_6t_5 inst_cell_48_55 (.BL(BL55),.BLN(BLN55),.WL(WL48));
sram_cell_6t_5 inst_cell_48_56 (.BL(BL56),.BLN(BLN56),.WL(WL48));
sram_cell_6t_5 inst_cell_48_57 (.BL(BL57),.BLN(BLN57),.WL(WL48));
sram_cell_6t_5 inst_cell_48_58 (.BL(BL58),.BLN(BLN58),.WL(WL48));
sram_cell_6t_5 inst_cell_48_59 (.BL(BL59),.BLN(BLN59),.WL(WL48));
sram_cell_6t_5 inst_cell_48_60 (.BL(BL60),.BLN(BLN60),.WL(WL48));
sram_cell_6t_5 inst_cell_48_61 (.BL(BL61),.BLN(BLN61),.WL(WL48));
sram_cell_6t_5 inst_cell_48_62 (.BL(BL62),.BLN(BLN62),.WL(WL48));
sram_cell_6t_5 inst_cell_48_63 (.BL(BL63),.BLN(BLN63),.WL(WL48));
sram_cell_6t_5 inst_cell_48_64 (.BL(BL64),.BLN(BLN64),.WL(WL48));
sram_cell_6t_5 inst_cell_48_65 (.BL(BL65),.BLN(BLN65),.WL(WL48));
sram_cell_6t_5 inst_cell_48_66 (.BL(BL66),.BLN(BLN66),.WL(WL48));
sram_cell_6t_5 inst_cell_48_67 (.BL(BL67),.BLN(BLN67),.WL(WL48));
sram_cell_6t_5 inst_cell_48_68 (.BL(BL68),.BLN(BLN68),.WL(WL48));
sram_cell_6t_5 inst_cell_48_69 (.BL(BL69),.BLN(BLN69),.WL(WL48));
sram_cell_6t_5 inst_cell_48_70 (.BL(BL70),.BLN(BLN70),.WL(WL48));
sram_cell_6t_5 inst_cell_48_71 (.BL(BL71),.BLN(BLN71),.WL(WL48));
sram_cell_6t_5 inst_cell_48_72 (.BL(BL72),.BLN(BLN72),.WL(WL48));
sram_cell_6t_5 inst_cell_48_73 (.BL(BL73),.BLN(BLN73),.WL(WL48));
sram_cell_6t_5 inst_cell_48_74 (.BL(BL74),.BLN(BLN74),.WL(WL48));
sram_cell_6t_5 inst_cell_48_75 (.BL(BL75),.BLN(BLN75),.WL(WL48));
sram_cell_6t_5 inst_cell_48_76 (.BL(BL76),.BLN(BLN76),.WL(WL48));
sram_cell_6t_5 inst_cell_48_77 (.BL(BL77),.BLN(BLN77),.WL(WL48));
sram_cell_6t_5 inst_cell_48_78 (.BL(BL78),.BLN(BLN78),.WL(WL48));
sram_cell_6t_5 inst_cell_48_79 (.BL(BL79),.BLN(BLN79),.WL(WL48));
sram_cell_6t_5 inst_cell_48_80 (.BL(BL80),.BLN(BLN80),.WL(WL48));
sram_cell_6t_5 inst_cell_48_81 (.BL(BL81),.BLN(BLN81),.WL(WL48));
sram_cell_6t_5 inst_cell_48_82 (.BL(BL82),.BLN(BLN82),.WL(WL48));
sram_cell_6t_5 inst_cell_48_83 (.BL(BL83),.BLN(BLN83),.WL(WL48));
sram_cell_6t_5 inst_cell_48_84 (.BL(BL84),.BLN(BLN84),.WL(WL48));
sram_cell_6t_5 inst_cell_48_85 (.BL(BL85),.BLN(BLN85),.WL(WL48));
sram_cell_6t_5 inst_cell_48_86 (.BL(BL86),.BLN(BLN86),.WL(WL48));
sram_cell_6t_5 inst_cell_48_87 (.BL(BL87),.BLN(BLN87),.WL(WL48));
sram_cell_6t_5 inst_cell_48_88 (.BL(BL88),.BLN(BLN88),.WL(WL48));
sram_cell_6t_5 inst_cell_48_89 (.BL(BL89),.BLN(BLN89),.WL(WL48));
sram_cell_6t_5 inst_cell_48_90 (.BL(BL90),.BLN(BLN90),.WL(WL48));
sram_cell_6t_5 inst_cell_48_91 (.BL(BL91),.BLN(BLN91),.WL(WL48));
sram_cell_6t_5 inst_cell_48_92 (.BL(BL92),.BLN(BLN92),.WL(WL48));
sram_cell_6t_5 inst_cell_48_93 (.BL(BL93),.BLN(BLN93),.WL(WL48));
sram_cell_6t_5 inst_cell_48_94 (.BL(BL94),.BLN(BLN94),.WL(WL48));
sram_cell_6t_5 inst_cell_48_95 (.BL(BL95),.BLN(BLN95),.WL(WL48));
sram_cell_6t_5 inst_cell_48_96 (.BL(BL96),.BLN(BLN96),.WL(WL48));
sram_cell_6t_5 inst_cell_48_97 (.BL(BL97),.BLN(BLN97),.WL(WL48));
sram_cell_6t_5 inst_cell_48_98 (.BL(BL98),.BLN(BLN98),.WL(WL48));
sram_cell_6t_5 inst_cell_48_99 (.BL(BL99),.BLN(BLN99),.WL(WL48));
sram_cell_6t_5 inst_cell_48_100 (.BL(BL100),.BLN(BLN100),.WL(WL48));
sram_cell_6t_5 inst_cell_48_101 (.BL(BL101),.BLN(BLN101),.WL(WL48));
sram_cell_6t_5 inst_cell_48_102 (.BL(BL102),.BLN(BLN102),.WL(WL48));
sram_cell_6t_5 inst_cell_48_103 (.BL(BL103),.BLN(BLN103),.WL(WL48));
sram_cell_6t_5 inst_cell_48_104 (.BL(BL104),.BLN(BLN104),.WL(WL48));
sram_cell_6t_5 inst_cell_48_105 (.BL(BL105),.BLN(BLN105),.WL(WL48));
sram_cell_6t_5 inst_cell_48_106 (.BL(BL106),.BLN(BLN106),.WL(WL48));
sram_cell_6t_5 inst_cell_48_107 (.BL(BL107),.BLN(BLN107),.WL(WL48));
sram_cell_6t_5 inst_cell_48_108 (.BL(BL108),.BLN(BLN108),.WL(WL48));
sram_cell_6t_5 inst_cell_48_109 (.BL(BL109),.BLN(BLN109),.WL(WL48));
sram_cell_6t_5 inst_cell_48_110 (.BL(BL110),.BLN(BLN110),.WL(WL48));
sram_cell_6t_5 inst_cell_48_111 (.BL(BL111),.BLN(BLN111),.WL(WL48));
sram_cell_6t_5 inst_cell_48_112 (.BL(BL112),.BLN(BLN112),.WL(WL48));
sram_cell_6t_5 inst_cell_48_113 (.BL(BL113),.BLN(BLN113),.WL(WL48));
sram_cell_6t_5 inst_cell_48_114 (.BL(BL114),.BLN(BLN114),.WL(WL48));
sram_cell_6t_5 inst_cell_48_115 (.BL(BL115),.BLN(BLN115),.WL(WL48));
sram_cell_6t_5 inst_cell_48_116 (.BL(BL116),.BLN(BLN116),.WL(WL48));
sram_cell_6t_5 inst_cell_48_117 (.BL(BL117),.BLN(BLN117),.WL(WL48));
sram_cell_6t_5 inst_cell_48_118 (.BL(BL118),.BLN(BLN118),.WL(WL48));
sram_cell_6t_5 inst_cell_48_119 (.BL(BL119),.BLN(BLN119),.WL(WL48));
sram_cell_6t_5 inst_cell_48_120 (.BL(BL120),.BLN(BLN120),.WL(WL48));
sram_cell_6t_5 inst_cell_48_121 (.BL(BL121),.BLN(BLN121),.WL(WL48));
sram_cell_6t_5 inst_cell_48_122 (.BL(BL122),.BLN(BLN122),.WL(WL48));
sram_cell_6t_5 inst_cell_48_123 (.BL(BL123),.BLN(BLN123),.WL(WL48));
sram_cell_6t_5 inst_cell_48_124 (.BL(BL124),.BLN(BLN124),.WL(WL48));
sram_cell_6t_5 inst_cell_48_125 (.BL(BL125),.BLN(BLN125),.WL(WL48));
sram_cell_6t_5 inst_cell_48_126 (.BL(BL126),.BLN(BLN126),.WL(WL48));
sram_cell_6t_5 inst_cell_48_127 (.BL(BL127),.BLN(BLN127),.WL(WL48));
sram_cell_6t_5 inst_cell_49_0 (.BL(BL0),.BLN(BLN0),.WL(WL49));
sram_cell_6t_5 inst_cell_49_1 (.BL(BL1),.BLN(BLN1),.WL(WL49));
sram_cell_6t_5 inst_cell_49_2 (.BL(BL2),.BLN(BLN2),.WL(WL49));
sram_cell_6t_5 inst_cell_49_3 (.BL(BL3),.BLN(BLN3),.WL(WL49));
sram_cell_6t_5 inst_cell_49_4 (.BL(BL4),.BLN(BLN4),.WL(WL49));
sram_cell_6t_5 inst_cell_49_5 (.BL(BL5),.BLN(BLN5),.WL(WL49));
sram_cell_6t_5 inst_cell_49_6 (.BL(BL6),.BLN(BLN6),.WL(WL49));
sram_cell_6t_5 inst_cell_49_7 (.BL(BL7),.BLN(BLN7),.WL(WL49));
sram_cell_6t_5 inst_cell_49_8 (.BL(BL8),.BLN(BLN8),.WL(WL49));
sram_cell_6t_5 inst_cell_49_9 (.BL(BL9),.BLN(BLN9),.WL(WL49));
sram_cell_6t_5 inst_cell_49_10 (.BL(BL10),.BLN(BLN10),.WL(WL49));
sram_cell_6t_5 inst_cell_49_11 (.BL(BL11),.BLN(BLN11),.WL(WL49));
sram_cell_6t_5 inst_cell_49_12 (.BL(BL12),.BLN(BLN12),.WL(WL49));
sram_cell_6t_5 inst_cell_49_13 (.BL(BL13),.BLN(BLN13),.WL(WL49));
sram_cell_6t_5 inst_cell_49_14 (.BL(BL14),.BLN(BLN14),.WL(WL49));
sram_cell_6t_5 inst_cell_49_15 (.BL(BL15),.BLN(BLN15),.WL(WL49));
sram_cell_6t_5 inst_cell_49_16 (.BL(BL16),.BLN(BLN16),.WL(WL49));
sram_cell_6t_5 inst_cell_49_17 (.BL(BL17),.BLN(BLN17),.WL(WL49));
sram_cell_6t_5 inst_cell_49_18 (.BL(BL18),.BLN(BLN18),.WL(WL49));
sram_cell_6t_5 inst_cell_49_19 (.BL(BL19),.BLN(BLN19),.WL(WL49));
sram_cell_6t_5 inst_cell_49_20 (.BL(BL20),.BLN(BLN20),.WL(WL49));
sram_cell_6t_5 inst_cell_49_21 (.BL(BL21),.BLN(BLN21),.WL(WL49));
sram_cell_6t_5 inst_cell_49_22 (.BL(BL22),.BLN(BLN22),.WL(WL49));
sram_cell_6t_5 inst_cell_49_23 (.BL(BL23),.BLN(BLN23),.WL(WL49));
sram_cell_6t_5 inst_cell_49_24 (.BL(BL24),.BLN(BLN24),.WL(WL49));
sram_cell_6t_5 inst_cell_49_25 (.BL(BL25),.BLN(BLN25),.WL(WL49));
sram_cell_6t_5 inst_cell_49_26 (.BL(BL26),.BLN(BLN26),.WL(WL49));
sram_cell_6t_5 inst_cell_49_27 (.BL(BL27),.BLN(BLN27),.WL(WL49));
sram_cell_6t_5 inst_cell_49_28 (.BL(BL28),.BLN(BLN28),.WL(WL49));
sram_cell_6t_5 inst_cell_49_29 (.BL(BL29),.BLN(BLN29),.WL(WL49));
sram_cell_6t_5 inst_cell_49_30 (.BL(BL30),.BLN(BLN30),.WL(WL49));
sram_cell_6t_5 inst_cell_49_31 (.BL(BL31),.BLN(BLN31),.WL(WL49));
sram_cell_6t_5 inst_cell_49_32 (.BL(BL32),.BLN(BLN32),.WL(WL49));
sram_cell_6t_5 inst_cell_49_33 (.BL(BL33),.BLN(BLN33),.WL(WL49));
sram_cell_6t_5 inst_cell_49_34 (.BL(BL34),.BLN(BLN34),.WL(WL49));
sram_cell_6t_5 inst_cell_49_35 (.BL(BL35),.BLN(BLN35),.WL(WL49));
sram_cell_6t_5 inst_cell_49_36 (.BL(BL36),.BLN(BLN36),.WL(WL49));
sram_cell_6t_5 inst_cell_49_37 (.BL(BL37),.BLN(BLN37),.WL(WL49));
sram_cell_6t_5 inst_cell_49_38 (.BL(BL38),.BLN(BLN38),.WL(WL49));
sram_cell_6t_5 inst_cell_49_39 (.BL(BL39),.BLN(BLN39),.WL(WL49));
sram_cell_6t_5 inst_cell_49_40 (.BL(BL40),.BLN(BLN40),.WL(WL49));
sram_cell_6t_5 inst_cell_49_41 (.BL(BL41),.BLN(BLN41),.WL(WL49));
sram_cell_6t_5 inst_cell_49_42 (.BL(BL42),.BLN(BLN42),.WL(WL49));
sram_cell_6t_5 inst_cell_49_43 (.BL(BL43),.BLN(BLN43),.WL(WL49));
sram_cell_6t_5 inst_cell_49_44 (.BL(BL44),.BLN(BLN44),.WL(WL49));
sram_cell_6t_5 inst_cell_49_45 (.BL(BL45),.BLN(BLN45),.WL(WL49));
sram_cell_6t_5 inst_cell_49_46 (.BL(BL46),.BLN(BLN46),.WL(WL49));
sram_cell_6t_5 inst_cell_49_47 (.BL(BL47),.BLN(BLN47),.WL(WL49));
sram_cell_6t_5 inst_cell_49_48 (.BL(BL48),.BLN(BLN48),.WL(WL49));
sram_cell_6t_5 inst_cell_49_49 (.BL(BL49),.BLN(BLN49),.WL(WL49));
sram_cell_6t_5 inst_cell_49_50 (.BL(BL50),.BLN(BLN50),.WL(WL49));
sram_cell_6t_5 inst_cell_49_51 (.BL(BL51),.BLN(BLN51),.WL(WL49));
sram_cell_6t_5 inst_cell_49_52 (.BL(BL52),.BLN(BLN52),.WL(WL49));
sram_cell_6t_5 inst_cell_49_53 (.BL(BL53),.BLN(BLN53),.WL(WL49));
sram_cell_6t_5 inst_cell_49_54 (.BL(BL54),.BLN(BLN54),.WL(WL49));
sram_cell_6t_5 inst_cell_49_55 (.BL(BL55),.BLN(BLN55),.WL(WL49));
sram_cell_6t_5 inst_cell_49_56 (.BL(BL56),.BLN(BLN56),.WL(WL49));
sram_cell_6t_5 inst_cell_49_57 (.BL(BL57),.BLN(BLN57),.WL(WL49));
sram_cell_6t_5 inst_cell_49_58 (.BL(BL58),.BLN(BLN58),.WL(WL49));
sram_cell_6t_5 inst_cell_49_59 (.BL(BL59),.BLN(BLN59),.WL(WL49));
sram_cell_6t_5 inst_cell_49_60 (.BL(BL60),.BLN(BLN60),.WL(WL49));
sram_cell_6t_5 inst_cell_49_61 (.BL(BL61),.BLN(BLN61),.WL(WL49));
sram_cell_6t_5 inst_cell_49_62 (.BL(BL62),.BLN(BLN62),.WL(WL49));
sram_cell_6t_5 inst_cell_49_63 (.BL(BL63),.BLN(BLN63),.WL(WL49));
sram_cell_6t_5 inst_cell_49_64 (.BL(BL64),.BLN(BLN64),.WL(WL49));
sram_cell_6t_5 inst_cell_49_65 (.BL(BL65),.BLN(BLN65),.WL(WL49));
sram_cell_6t_5 inst_cell_49_66 (.BL(BL66),.BLN(BLN66),.WL(WL49));
sram_cell_6t_5 inst_cell_49_67 (.BL(BL67),.BLN(BLN67),.WL(WL49));
sram_cell_6t_5 inst_cell_49_68 (.BL(BL68),.BLN(BLN68),.WL(WL49));
sram_cell_6t_5 inst_cell_49_69 (.BL(BL69),.BLN(BLN69),.WL(WL49));
sram_cell_6t_5 inst_cell_49_70 (.BL(BL70),.BLN(BLN70),.WL(WL49));
sram_cell_6t_5 inst_cell_49_71 (.BL(BL71),.BLN(BLN71),.WL(WL49));
sram_cell_6t_5 inst_cell_49_72 (.BL(BL72),.BLN(BLN72),.WL(WL49));
sram_cell_6t_5 inst_cell_49_73 (.BL(BL73),.BLN(BLN73),.WL(WL49));
sram_cell_6t_5 inst_cell_49_74 (.BL(BL74),.BLN(BLN74),.WL(WL49));
sram_cell_6t_5 inst_cell_49_75 (.BL(BL75),.BLN(BLN75),.WL(WL49));
sram_cell_6t_5 inst_cell_49_76 (.BL(BL76),.BLN(BLN76),.WL(WL49));
sram_cell_6t_5 inst_cell_49_77 (.BL(BL77),.BLN(BLN77),.WL(WL49));
sram_cell_6t_5 inst_cell_49_78 (.BL(BL78),.BLN(BLN78),.WL(WL49));
sram_cell_6t_5 inst_cell_49_79 (.BL(BL79),.BLN(BLN79),.WL(WL49));
sram_cell_6t_5 inst_cell_49_80 (.BL(BL80),.BLN(BLN80),.WL(WL49));
sram_cell_6t_5 inst_cell_49_81 (.BL(BL81),.BLN(BLN81),.WL(WL49));
sram_cell_6t_5 inst_cell_49_82 (.BL(BL82),.BLN(BLN82),.WL(WL49));
sram_cell_6t_5 inst_cell_49_83 (.BL(BL83),.BLN(BLN83),.WL(WL49));
sram_cell_6t_5 inst_cell_49_84 (.BL(BL84),.BLN(BLN84),.WL(WL49));
sram_cell_6t_5 inst_cell_49_85 (.BL(BL85),.BLN(BLN85),.WL(WL49));
sram_cell_6t_5 inst_cell_49_86 (.BL(BL86),.BLN(BLN86),.WL(WL49));
sram_cell_6t_5 inst_cell_49_87 (.BL(BL87),.BLN(BLN87),.WL(WL49));
sram_cell_6t_5 inst_cell_49_88 (.BL(BL88),.BLN(BLN88),.WL(WL49));
sram_cell_6t_5 inst_cell_49_89 (.BL(BL89),.BLN(BLN89),.WL(WL49));
sram_cell_6t_5 inst_cell_49_90 (.BL(BL90),.BLN(BLN90),.WL(WL49));
sram_cell_6t_5 inst_cell_49_91 (.BL(BL91),.BLN(BLN91),.WL(WL49));
sram_cell_6t_5 inst_cell_49_92 (.BL(BL92),.BLN(BLN92),.WL(WL49));
sram_cell_6t_5 inst_cell_49_93 (.BL(BL93),.BLN(BLN93),.WL(WL49));
sram_cell_6t_5 inst_cell_49_94 (.BL(BL94),.BLN(BLN94),.WL(WL49));
sram_cell_6t_5 inst_cell_49_95 (.BL(BL95),.BLN(BLN95),.WL(WL49));
sram_cell_6t_5 inst_cell_49_96 (.BL(BL96),.BLN(BLN96),.WL(WL49));
sram_cell_6t_5 inst_cell_49_97 (.BL(BL97),.BLN(BLN97),.WL(WL49));
sram_cell_6t_5 inst_cell_49_98 (.BL(BL98),.BLN(BLN98),.WL(WL49));
sram_cell_6t_5 inst_cell_49_99 (.BL(BL99),.BLN(BLN99),.WL(WL49));
sram_cell_6t_5 inst_cell_49_100 (.BL(BL100),.BLN(BLN100),.WL(WL49));
sram_cell_6t_5 inst_cell_49_101 (.BL(BL101),.BLN(BLN101),.WL(WL49));
sram_cell_6t_5 inst_cell_49_102 (.BL(BL102),.BLN(BLN102),.WL(WL49));
sram_cell_6t_5 inst_cell_49_103 (.BL(BL103),.BLN(BLN103),.WL(WL49));
sram_cell_6t_5 inst_cell_49_104 (.BL(BL104),.BLN(BLN104),.WL(WL49));
sram_cell_6t_5 inst_cell_49_105 (.BL(BL105),.BLN(BLN105),.WL(WL49));
sram_cell_6t_5 inst_cell_49_106 (.BL(BL106),.BLN(BLN106),.WL(WL49));
sram_cell_6t_5 inst_cell_49_107 (.BL(BL107),.BLN(BLN107),.WL(WL49));
sram_cell_6t_5 inst_cell_49_108 (.BL(BL108),.BLN(BLN108),.WL(WL49));
sram_cell_6t_5 inst_cell_49_109 (.BL(BL109),.BLN(BLN109),.WL(WL49));
sram_cell_6t_5 inst_cell_49_110 (.BL(BL110),.BLN(BLN110),.WL(WL49));
sram_cell_6t_5 inst_cell_49_111 (.BL(BL111),.BLN(BLN111),.WL(WL49));
sram_cell_6t_5 inst_cell_49_112 (.BL(BL112),.BLN(BLN112),.WL(WL49));
sram_cell_6t_5 inst_cell_49_113 (.BL(BL113),.BLN(BLN113),.WL(WL49));
sram_cell_6t_5 inst_cell_49_114 (.BL(BL114),.BLN(BLN114),.WL(WL49));
sram_cell_6t_5 inst_cell_49_115 (.BL(BL115),.BLN(BLN115),.WL(WL49));
sram_cell_6t_5 inst_cell_49_116 (.BL(BL116),.BLN(BLN116),.WL(WL49));
sram_cell_6t_5 inst_cell_49_117 (.BL(BL117),.BLN(BLN117),.WL(WL49));
sram_cell_6t_5 inst_cell_49_118 (.BL(BL118),.BLN(BLN118),.WL(WL49));
sram_cell_6t_5 inst_cell_49_119 (.BL(BL119),.BLN(BLN119),.WL(WL49));
sram_cell_6t_5 inst_cell_49_120 (.BL(BL120),.BLN(BLN120),.WL(WL49));
sram_cell_6t_5 inst_cell_49_121 (.BL(BL121),.BLN(BLN121),.WL(WL49));
sram_cell_6t_5 inst_cell_49_122 (.BL(BL122),.BLN(BLN122),.WL(WL49));
sram_cell_6t_5 inst_cell_49_123 (.BL(BL123),.BLN(BLN123),.WL(WL49));
sram_cell_6t_5 inst_cell_49_124 (.BL(BL124),.BLN(BLN124),.WL(WL49));
sram_cell_6t_5 inst_cell_49_125 (.BL(BL125),.BLN(BLN125),.WL(WL49));
sram_cell_6t_5 inst_cell_49_126 (.BL(BL126),.BLN(BLN126),.WL(WL49));
sram_cell_6t_5 inst_cell_49_127 (.BL(BL127),.BLN(BLN127),.WL(WL49));
sram_cell_6t_5 inst_cell_50_0 (.BL(BL0),.BLN(BLN0),.WL(WL50));
sram_cell_6t_5 inst_cell_50_1 (.BL(BL1),.BLN(BLN1),.WL(WL50));
sram_cell_6t_5 inst_cell_50_2 (.BL(BL2),.BLN(BLN2),.WL(WL50));
sram_cell_6t_5 inst_cell_50_3 (.BL(BL3),.BLN(BLN3),.WL(WL50));
sram_cell_6t_5 inst_cell_50_4 (.BL(BL4),.BLN(BLN4),.WL(WL50));
sram_cell_6t_5 inst_cell_50_5 (.BL(BL5),.BLN(BLN5),.WL(WL50));
sram_cell_6t_5 inst_cell_50_6 (.BL(BL6),.BLN(BLN6),.WL(WL50));
sram_cell_6t_5 inst_cell_50_7 (.BL(BL7),.BLN(BLN7),.WL(WL50));
sram_cell_6t_5 inst_cell_50_8 (.BL(BL8),.BLN(BLN8),.WL(WL50));
sram_cell_6t_5 inst_cell_50_9 (.BL(BL9),.BLN(BLN9),.WL(WL50));
sram_cell_6t_5 inst_cell_50_10 (.BL(BL10),.BLN(BLN10),.WL(WL50));
sram_cell_6t_5 inst_cell_50_11 (.BL(BL11),.BLN(BLN11),.WL(WL50));
sram_cell_6t_5 inst_cell_50_12 (.BL(BL12),.BLN(BLN12),.WL(WL50));
sram_cell_6t_5 inst_cell_50_13 (.BL(BL13),.BLN(BLN13),.WL(WL50));
sram_cell_6t_5 inst_cell_50_14 (.BL(BL14),.BLN(BLN14),.WL(WL50));
sram_cell_6t_5 inst_cell_50_15 (.BL(BL15),.BLN(BLN15),.WL(WL50));
sram_cell_6t_5 inst_cell_50_16 (.BL(BL16),.BLN(BLN16),.WL(WL50));
sram_cell_6t_5 inst_cell_50_17 (.BL(BL17),.BLN(BLN17),.WL(WL50));
sram_cell_6t_5 inst_cell_50_18 (.BL(BL18),.BLN(BLN18),.WL(WL50));
sram_cell_6t_5 inst_cell_50_19 (.BL(BL19),.BLN(BLN19),.WL(WL50));
sram_cell_6t_5 inst_cell_50_20 (.BL(BL20),.BLN(BLN20),.WL(WL50));
sram_cell_6t_5 inst_cell_50_21 (.BL(BL21),.BLN(BLN21),.WL(WL50));
sram_cell_6t_5 inst_cell_50_22 (.BL(BL22),.BLN(BLN22),.WL(WL50));
sram_cell_6t_5 inst_cell_50_23 (.BL(BL23),.BLN(BLN23),.WL(WL50));
sram_cell_6t_5 inst_cell_50_24 (.BL(BL24),.BLN(BLN24),.WL(WL50));
sram_cell_6t_5 inst_cell_50_25 (.BL(BL25),.BLN(BLN25),.WL(WL50));
sram_cell_6t_5 inst_cell_50_26 (.BL(BL26),.BLN(BLN26),.WL(WL50));
sram_cell_6t_5 inst_cell_50_27 (.BL(BL27),.BLN(BLN27),.WL(WL50));
sram_cell_6t_5 inst_cell_50_28 (.BL(BL28),.BLN(BLN28),.WL(WL50));
sram_cell_6t_5 inst_cell_50_29 (.BL(BL29),.BLN(BLN29),.WL(WL50));
sram_cell_6t_5 inst_cell_50_30 (.BL(BL30),.BLN(BLN30),.WL(WL50));
sram_cell_6t_5 inst_cell_50_31 (.BL(BL31),.BLN(BLN31),.WL(WL50));
sram_cell_6t_5 inst_cell_50_32 (.BL(BL32),.BLN(BLN32),.WL(WL50));
sram_cell_6t_5 inst_cell_50_33 (.BL(BL33),.BLN(BLN33),.WL(WL50));
sram_cell_6t_5 inst_cell_50_34 (.BL(BL34),.BLN(BLN34),.WL(WL50));
sram_cell_6t_5 inst_cell_50_35 (.BL(BL35),.BLN(BLN35),.WL(WL50));
sram_cell_6t_5 inst_cell_50_36 (.BL(BL36),.BLN(BLN36),.WL(WL50));
sram_cell_6t_5 inst_cell_50_37 (.BL(BL37),.BLN(BLN37),.WL(WL50));
sram_cell_6t_5 inst_cell_50_38 (.BL(BL38),.BLN(BLN38),.WL(WL50));
sram_cell_6t_5 inst_cell_50_39 (.BL(BL39),.BLN(BLN39),.WL(WL50));
sram_cell_6t_5 inst_cell_50_40 (.BL(BL40),.BLN(BLN40),.WL(WL50));
sram_cell_6t_5 inst_cell_50_41 (.BL(BL41),.BLN(BLN41),.WL(WL50));
sram_cell_6t_5 inst_cell_50_42 (.BL(BL42),.BLN(BLN42),.WL(WL50));
sram_cell_6t_5 inst_cell_50_43 (.BL(BL43),.BLN(BLN43),.WL(WL50));
sram_cell_6t_5 inst_cell_50_44 (.BL(BL44),.BLN(BLN44),.WL(WL50));
sram_cell_6t_5 inst_cell_50_45 (.BL(BL45),.BLN(BLN45),.WL(WL50));
sram_cell_6t_5 inst_cell_50_46 (.BL(BL46),.BLN(BLN46),.WL(WL50));
sram_cell_6t_5 inst_cell_50_47 (.BL(BL47),.BLN(BLN47),.WL(WL50));
sram_cell_6t_5 inst_cell_50_48 (.BL(BL48),.BLN(BLN48),.WL(WL50));
sram_cell_6t_5 inst_cell_50_49 (.BL(BL49),.BLN(BLN49),.WL(WL50));
sram_cell_6t_5 inst_cell_50_50 (.BL(BL50),.BLN(BLN50),.WL(WL50));
sram_cell_6t_5 inst_cell_50_51 (.BL(BL51),.BLN(BLN51),.WL(WL50));
sram_cell_6t_5 inst_cell_50_52 (.BL(BL52),.BLN(BLN52),.WL(WL50));
sram_cell_6t_5 inst_cell_50_53 (.BL(BL53),.BLN(BLN53),.WL(WL50));
sram_cell_6t_5 inst_cell_50_54 (.BL(BL54),.BLN(BLN54),.WL(WL50));
sram_cell_6t_5 inst_cell_50_55 (.BL(BL55),.BLN(BLN55),.WL(WL50));
sram_cell_6t_5 inst_cell_50_56 (.BL(BL56),.BLN(BLN56),.WL(WL50));
sram_cell_6t_5 inst_cell_50_57 (.BL(BL57),.BLN(BLN57),.WL(WL50));
sram_cell_6t_5 inst_cell_50_58 (.BL(BL58),.BLN(BLN58),.WL(WL50));
sram_cell_6t_5 inst_cell_50_59 (.BL(BL59),.BLN(BLN59),.WL(WL50));
sram_cell_6t_5 inst_cell_50_60 (.BL(BL60),.BLN(BLN60),.WL(WL50));
sram_cell_6t_5 inst_cell_50_61 (.BL(BL61),.BLN(BLN61),.WL(WL50));
sram_cell_6t_5 inst_cell_50_62 (.BL(BL62),.BLN(BLN62),.WL(WL50));
sram_cell_6t_5 inst_cell_50_63 (.BL(BL63),.BLN(BLN63),.WL(WL50));
sram_cell_6t_5 inst_cell_50_64 (.BL(BL64),.BLN(BLN64),.WL(WL50));
sram_cell_6t_5 inst_cell_50_65 (.BL(BL65),.BLN(BLN65),.WL(WL50));
sram_cell_6t_5 inst_cell_50_66 (.BL(BL66),.BLN(BLN66),.WL(WL50));
sram_cell_6t_5 inst_cell_50_67 (.BL(BL67),.BLN(BLN67),.WL(WL50));
sram_cell_6t_5 inst_cell_50_68 (.BL(BL68),.BLN(BLN68),.WL(WL50));
sram_cell_6t_5 inst_cell_50_69 (.BL(BL69),.BLN(BLN69),.WL(WL50));
sram_cell_6t_5 inst_cell_50_70 (.BL(BL70),.BLN(BLN70),.WL(WL50));
sram_cell_6t_5 inst_cell_50_71 (.BL(BL71),.BLN(BLN71),.WL(WL50));
sram_cell_6t_5 inst_cell_50_72 (.BL(BL72),.BLN(BLN72),.WL(WL50));
sram_cell_6t_5 inst_cell_50_73 (.BL(BL73),.BLN(BLN73),.WL(WL50));
sram_cell_6t_5 inst_cell_50_74 (.BL(BL74),.BLN(BLN74),.WL(WL50));
sram_cell_6t_5 inst_cell_50_75 (.BL(BL75),.BLN(BLN75),.WL(WL50));
sram_cell_6t_5 inst_cell_50_76 (.BL(BL76),.BLN(BLN76),.WL(WL50));
sram_cell_6t_5 inst_cell_50_77 (.BL(BL77),.BLN(BLN77),.WL(WL50));
sram_cell_6t_5 inst_cell_50_78 (.BL(BL78),.BLN(BLN78),.WL(WL50));
sram_cell_6t_5 inst_cell_50_79 (.BL(BL79),.BLN(BLN79),.WL(WL50));
sram_cell_6t_5 inst_cell_50_80 (.BL(BL80),.BLN(BLN80),.WL(WL50));
sram_cell_6t_5 inst_cell_50_81 (.BL(BL81),.BLN(BLN81),.WL(WL50));
sram_cell_6t_5 inst_cell_50_82 (.BL(BL82),.BLN(BLN82),.WL(WL50));
sram_cell_6t_5 inst_cell_50_83 (.BL(BL83),.BLN(BLN83),.WL(WL50));
sram_cell_6t_5 inst_cell_50_84 (.BL(BL84),.BLN(BLN84),.WL(WL50));
sram_cell_6t_5 inst_cell_50_85 (.BL(BL85),.BLN(BLN85),.WL(WL50));
sram_cell_6t_5 inst_cell_50_86 (.BL(BL86),.BLN(BLN86),.WL(WL50));
sram_cell_6t_5 inst_cell_50_87 (.BL(BL87),.BLN(BLN87),.WL(WL50));
sram_cell_6t_5 inst_cell_50_88 (.BL(BL88),.BLN(BLN88),.WL(WL50));
sram_cell_6t_5 inst_cell_50_89 (.BL(BL89),.BLN(BLN89),.WL(WL50));
sram_cell_6t_5 inst_cell_50_90 (.BL(BL90),.BLN(BLN90),.WL(WL50));
sram_cell_6t_5 inst_cell_50_91 (.BL(BL91),.BLN(BLN91),.WL(WL50));
sram_cell_6t_5 inst_cell_50_92 (.BL(BL92),.BLN(BLN92),.WL(WL50));
sram_cell_6t_5 inst_cell_50_93 (.BL(BL93),.BLN(BLN93),.WL(WL50));
sram_cell_6t_5 inst_cell_50_94 (.BL(BL94),.BLN(BLN94),.WL(WL50));
sram_cell_6t_5 inst_cell_50_95 (.BL(BL95),.BLN(BLN95),.WL(WL50));
sram_cell_6t_5 inst_cell_50_96 (.BL(BL96),.BLN(BLN96),.WL(WL50));
sram_cell_6t_5 inst_cell_50_97 (.BL(BL97),.BLN(BLN97),.WL(WL50));
sram_cell_6t_5 inst_cell_50_98 (.BL(BL98),.BLN(BLN98),.WL(WL50));
sram_cell_6t_5 inst_cell_50_99 (.BL(BL99),.BLN(BLN99),.WL(WL50));
sram_cell_6t_5 inst_cell_50_100 (.BL(BL100),.BLN(BLN100),.WL(WL50));
sram_cell_6t_5 inst_cell_50_101 (.BL(BL101),.BLN(BLN101),.WL(WL50));
sram_cell_6t_5 inst_cell_50_102 (.BL(BL102),.BLN(BLN102),.WL(WL50));
sram_cell_6t_5 inst_cell_50_103 (.BL(BL103),.BLN(BLN103),.WL(WL50));
sram_cell_6t_5 inst_cell_50_104 (.BL(BL104),.BLN(BLN104),.WL(WL50));
sram_cell_6t_5 inst_cell_50_105 (.BL(BL105),.BLN(BLN105),.WL(WL50));
sram_cell_6t_5 inst_cell_50_106 (.BL(BL106),.BLN(BLN106),.WL(WL50));
sram_cell_6t_5 inst_cell_50_107 (.BL(BL107),.BLN(BLN107),.WL(WL50));
sram_cell_6t_5 inst_cell_50_108 (.BL(BL108),.BLN(BLN108),.WL(WL50));
sram_cell_6t_5 inst_cell_50_109 (.BL(BL109),.BLN(BLN109),.WL(WL50));
sram_cell_6t_5 inst_cell_50_110 (.BL(BL110),.BLN(BLN110),.WL(WL50));
sram_cell_6t_5 inst_cell_50_111 (.BL(BL111),.BLN(BLN111),.WL(WL50));
sram_cell_6t_5 inst_cell_50_112 (.BL(BL112),.BLN(BLN112),.WL(WL50));
sram_cell_6t_5 inst_cell_50_113 (.BL(BL113),.BLN(BLN113),.WL(WL50));
sram_cell_6t_5 inst_cell_50_114 (.BL(BL114),.BLN(BLN114),.WL(WL50));
sram_cell_6t_5 inst_cell_50_115 (.BL(BL115),.BLN(BLN115),.WL(WL50));
sram_cell_6t_5 inst_cell_50_116 (.BL(BL116),.BLN(BLN116),.WL(WL50));
sram_cell_6t_5 inst_cell_50_117 (.BL(BL117),.BLN(BLN117),.WL(WL50));
sram_cell_6t_5 inst_cell_50_118 (.BL(BL118),.BLN(BLN118),.WL(WL50));
sram_cell_6t_5 inst_cell_50_119 (.BL(BL119),.BLN(BLN119),.WL(WL50));
sram_cell_6t_5 inst_cell_50_120 (.BL(BL120),.BLN(BLN120),.WL(WL50));
sram_cell_6t_5 inst_cell_50_121 (.BL(BL121),.BLN(BLN121),.WL(WL50));
sram_cell_6t_5 inst_cell_50_122 (.BL(BL122),.BLN(BLN122),.WL(WL50));
sram_cell_6t_5 inst_cell_50_123 (.BL(BL123),.BLN(BLN123),.WL(WL50));
sram_cell_6t_5 inst_cell_50_124 (.BL(BL124),.BLN(BLN124),.WL(WL50));
sram_cell_6t_5 inst_cell_50_125 (.BL(BL125),.BLN(BLN125),.WL(WL50));
sram_cell_6t_5 inst_cell_50_126 (.BL(BL126),.BLN(BLN126),.WL(WL50));
sram_cell_6t_5 inst_cell_50_127 (.BL(BL127),.BLN(BLN127),.WL(WL50));
sram_cell_6t_5 inst_cell_51_0 (.BL(BL0),.BLN(BLN0),.WL(WL51));
sram_cell_6t_5 inst_cell_51_1 (.BL(BL1),.BLN(BLN1),.WL(WL51));
sram_cell_6t_5 inst_cell_51_2 (.BL(BL2),.BLN(BLN2),.WL(WL51));
sram_cell_6t_5 inst_cell_51_3 (.BL(BL3),.BLN(BLN3),.WL(WL51));
sram_cell_6t_5 inst_cell_51_4 (.BL(BL4),.BLN(BLN4),.WL(WL51));
sram_cell_6t_5 inst_cell_51_5 (.BL(BL5),.BLN(BLN5),.WL(WL51));
sram_cell_6t_5 inst_cell_51_6 (.BL(BL6),.BLN(BLN6),.WL(WL51));
sram_cell_6t_5 inst_cell_51_7 (.BL(BL7),.BLN(BLN7),.WL(WL51));
sram_cell_6t_5 inst_cell_51_8 (.BL(BL8),.BLN(BLN8),.WL(WL51));
sram_cell_6t_5 inst_cell_51_9 (.BL(BL9),.BLN(BLN9),.WL(WL51));
sram_cell_6t_5 inst_cell_51_10 (.BL(BL10),.BLN(BLN10),.WL(WL51));
sram_cell_6t_5 inst_cell_51_11 (.BL(BL11),.BLN(BLN11),.WL(WL51));
sram_cell_6t_5 inst_cell_51_12 (.BL(BL12),.BLN(BLN12),.WL(WL51));
sram_cell_6t_5 inst_cell_51_13 (.BL(BL13),.BLN(BLN13),.WL(WL51));
sram_cell_6t_5 inst_cell_51_14 (.BL(BL14),.BLN(BLN14),.WL(WL51));
sram_cell_6t_5 inst_cell_51_15 (.BL(BL15),.BLN(BLN15),.WL(WL51));
sram_cell_6t_5 inst_cell_51_16 (.BL(BL16),.BLN(BLN16),.WL(WL51));
sram_cell_6t_5 inst_cell_51_17 (.BL(BL17),.BLN(BLN17),.WL(WL51));
sram_cell_6t_5 inst_cell_51_18 (.BL(BL18),.BLN(BLN18),.WL(WL51));
sram_cell_6t_5 inst_cell_51_19 (.BL(BL19),.BLN(BLN19),.WL(WL51));
sram_cell_6t_5 inst_cell_51_20 (.BL(BL20),.BLN(BLN20),.WL(WL51));
sram_cell_6t_5 inst_cell_51_21 (.BL(BL21),.BLN(BLN21),.WL(WL51));
sram_cell_6t_5 inst_cell_51_22 (.BL(BL22),.BLN(BLN22),.WL(WL51));
sram_cell_6t_5 inst_cell_51_23 (.BL(BL23),.BLN(BLN23),.WL(WL51));
sram_cell_6t_5 inst_cell_51_24 (.BL(BL24),.BLN(BLN24),.WL(WL51));
sram_cell_6t_5 inst_cell_51_25 (.BL(BL25),.BLN(BLN25),.WL(WL51));
sram_cell_6t_5 inst_cell_51_26 (.BL(BL26),.BLN(BLN26),.WL(WL51));
sram_cell_6t_5 inst_cell_51_27 (.BL(BL27),.BLN(BLN27),.WL(WL51));
sram_cell_6t_5 inst_cell_51_28 (.BL(BL28),.BLN(BLN28),.WL(WL51));
sram_cell_6t_5 inst_cell_51_29 (.BL(BL29),.BLN(BLN29),.WL(WL51));
sram_cell_6t_5 inst_cell_51_30 (.BL(BL30),.BLN(BLN30),.WL(WL51));
sram_cell_6t_5 inst_cell_51_31 (.BL(BL31),.BLN(BLN31),.WL(WL51));
sram_cell_6t_5 inst_cell_51_32 (.BL(BL32),.BLN(BLN32),.WL(WL51));
sram_cell_6t_5 inst_cell_51_33 (.BL(BL33),.BLN(BLN33),.WL(WL51));
sram_cell_6t_5 inst_cell_51_34 (.BL(BL34),.BLN(BLN34),.WL(WL51));
sram_cell_6t_5 inst_cell_51_35 (.BL(BL35),.BLN(BLN35),.WL(WL51));
sram_cell_6t_5 inst_cell_51_36 (.BL(BL36),.BLN(BLN36),.WL(WL51));
sram_cell_6t_5 inst_cell_51_37 (.BL(BL37),.BLN(BLN37),.WL(WL51));
sram_cell_6t_5 inst_cell_51_38 (.BL(BL38),.BLN(BLN38),.WL(WL51));
sram_cell_6t_5 inst_cell_51_39 (.BL(BL39),.BLN(BLN39),.WL(WL51));
sram_cell_6t_5 inst_cell_51_40 (.BL(BL40),.BLN(BLN40),.WL(WL51));
sram_cell_6t_5 inst_cell_51_41 (.BL(BL41),.BLN(BLN41),.WL(WL51));
sram_cell_6t_5 inst_cell_51_42 (.BL(BL42),.BLN(BLN42),.WL(WL51));
sram_cell_6t_5 inst_cell_51_43 (.BL(BL43),.BLN(BLN43),.WL(WL51));
sram_cell_6t_5 inst_cell_51_44 (.BL(BL44),.BLN(BLN44),.WL(WL51));
sram_cell_6t_5 inst_cell_51_45 (.BL(BL45),.BLN(BLN45),.WL(WL51));
sram_cell_6t_5 inst_cell_51_46 (.BL(BL46),.BLN(BLN46),.WL(WL51));
sram_cell_6t_5 inst_cell_51_47 (.BL(BL47),.BLN(BLN47),.WL(WL51));
sram_cell_6t_5 inst_cell_51_48 (.BL(BL48),.BLN(BLN48),.WL(WL51));
sram_cell_6t_5 inst_cell_51_49 (.BL(BL49),.BLN(BLN49),.WL(WL51));
sram_cell_6t_5 inst_cell_51_50 (.BL(BL50),.BLN(BLN50),.WL(WL51));
sram_cell_6t_5 inst_cell_51_51 (.BL(BL51),.BLN(BLN51),.WL(WL51));
sram_cell_6t_5 inst_cell_51_52 (.BL(BL52),.BLN(BLN52),.WL(WL51));
sram_cell_6t_5 inst_cell_51_53 (.BL(BL53),.BLN(BLN53),.WL(WL51));
sram_cell_6t_5 inst_cell_51_54 (.BL(BL54),.BLN(BLN54),.WL(WL51));
sram_cell_6t_5 inst_cell_51_55 (.BL(BL55),.BLN(BLN55),.WL(WL51));
sram_cell_6t_5 inst_cell_51_56 (.BL(BL56),.BLN(BLN56),.WL(WL51));
sram_cell_6t_5 inst_cell_51_57 (.BL(BL57),.BLN(BLN57),.WL(WL51));
sram_cell_6t_5 inst_cell_51_58 (.BL(BL58),.BLN(BLN58),.WL(WL51));
sram_cell_6t_5 inst_cell_51_59 (.BL(BL59),.BLN(BLN59),.WL(WL51));
sram_cell_6t_5 inst_cell_51_60 (.BL(BL60),.BLN(BLN60),.WL(WL51));
sram_cell_6t_5 inst_cell_51_61 (.BL(BL61),.BLN(BLN61),.WL(WL51));
sram_cell_6t_5 inst_cell_51_62 (.BL(BL62),.BLN(BLN62),.WL(WL51));
sram_cell_6t_5 inst_cell_51_63 (.BL(BL63),.BLN(BLN63),.WL(WL51));
sram_cell_6t_5 inst_cell_51_64 (.BL(BL64),.BLN(BLN64),.WL(WL51));
sram_cell_6t_5 inst_cell_51_65 (.BL(BL65),.BLN(BLN65),.WL(WL51));
sram_cell_6t_5 inst_cell_51_66 (.BL(BL66),.BLN(BLN66),.WL(WL51));
sram_cell_6t_5 inst_cell_51_67 (.BL(BL67),.BLN(BLN67),.WL(WL51));
sram_cell_6t_5 inst_cell_51_68 (.BL(BL68),.BLN(BLN68),.WL(WL51));
sram_cell_6t_5 inst_cell_51_69 (.BL(BL69),.BLN(BLN69),.WL(WL51));
sram_cell_6t_5 inst_cell_51_70 (.BL(BL70),.BLN(BLN70),.WL(WL51));
sram_cell_6t_5 inst_cell_51_71 (.BL(BL71),.BLN(BLN71),.WL(WL51));
sram_cell_6t_5 inst_cell_51_72 (.BL(BL72),.BLN(BLN72),.WL(WL51));
sram_cell_6t_5 inst_cell_51_73 (.BL(BL73),.BLN(BLN73),.WL(WL51));
sram_cell_6t_5 inst_cell_51_74 (.BL(BL74),.BLN(BLN74),.WL(WL51));
sram_cell_6t_5 inst_cell_51_75 (.BL(BL75),.BLN(BLN75),.WL(WL51));
sram_cell_6t_5 inst_cell_51_76 (.BL(BL76),.BLN(BLN76),.WL(WL51));
sram_cell_6t_5 inst_cell_51_77 (.BL(BL77),.BLN(BLN77),.WL(WL51));
sram_cell_6t_5 inst_cell_51_78 (.BL(BL78),.BLN(BLN78),.WL(WL51));
sram_cell_6t_5 inst_cell_51_79 (.BL(BL79),.BLN(BLN79),.WL(WL51));
sram_cell_6t_5 inst_cell_51_80 (.BL(BL80),.BLN(BLN80),.WL(WL51));
sram_cell_6t_5 inst_cell_51_81 (.BL(BL81),.BLN(BLN81),.WL(WL51));
sram_cell_6t_5 inst_cell_51_82 (.BL(BL82),.BLN(BLN82),.WL(WL51));
sram_cell_6t_5 inst_cell_51_83 (.BL(BL83),.BLN(BLN83),.WL(WL51));
sram_cell_6t_5 inst_cell_51_84 (.BL(BL84),.BLN(BLN84),.WL(WL51));
sram_cell_6t_5 inst_cell_51_85 (.BL(BL85),.BLN(BLN85),.WL(WL51));
sram_cell_6t_5 inst_cell_51_86 (.BL(BL86),.BLN(BLN86),.WL(WL51));
sram_cell_6t_5 inst_cell_51_87 (.BL(BL87),.BLN(BLN87),.WL(WL51));
sram_cell_6t_5 inst_cell_51_88 (.BL(BL88),.BLN(BLN88),.WL(WL51));
sram_cell_6t_5 inst_cell_51_89 (.BL(BL89),.BLN(BLN89),.WL(WL51));
sram_cell_6t_5 inst_cell_51_90 (.BL(BL90),.BLN(BLN90),.WL(WL51));
sram_cell_6t_5 inst_cell_51_91 (.BL(BL91),.BLN(BLN91),.WL(WL51));
sram_cell_6t_5 inst_cell_51_92 (.BL(BL92),.BLN(BLN92),.WL(WL51));
sram_cell_6t_5 inst_cell_51_93 (.BL(BL93),.BLN(BLN93),.WL(WL51));
sram_cell_6t_5 inst_cell_51_94 (.BL(BL94),.BLN(BLN94),.WL(WL51));
sram_cell_6t_5 inst_cell_51_95 (.BL(BL95),.BLN(BLN95),.WL(WL51));
sram_cell_6t_5 inst_cell_51_96 (.BL(BL96),.BLN(BLN96),.WL(WL51));
sram_cell_6t_5 inst_cell_51_97 (.BL(BL97),.BLN(BLN97),.WL(WL51));
sram_cell_6t_5 inst_cell_51_98 (.BL(BL98),.BLN(BLN98),.WL(WL51));
sram_cell_6t_5 inst_cell_51_99 (.BL(BL99),.BLN(BLN99),.WL(WL51));
sram_cell_6t_5 inst_cell_51_100 (.BL(BL100),.BLN(BLN100),.WL(WL51));
sram_cell_6t_5 inst_cell_51_101 (.BL(BL101),.BLN(BLN101),.WL(WL51));
sram_cell_6t_5 inst_cell_51_102 (.BL(BL102),.BLN(BLN102),.WL(WL51));
sram_cell_6t_5 inst_cell_51_103 (.BL(BL103),.BLN(BLN103),.WL(WL51));
sram_cell_6t_5 inst_cell_51_104 (.BL(BL104),.BLN(BLN104),.WL(WL51));
sram_cell_6t_5 inst_cell_51_105 (.BL(BL105),.BLN(BLN105),.WL(WL51));
sram_cell_6t_5 inst_cell_51_106 (.BL(BL106),.BLN(BLN106),.WL(WL51));
sram_cell_6t_5 inst_cell_51_107 (.BL(BL107),.BLN(BLN107),.WL(WL51));
sram_cell_6t_5 inst_cell_51_108 (.BL(BL108),.BLN(BLN108),.WL(WL51));
sram_cell_6t_5 inst_cell_51_109 (.BL(BL109),.BLN(BLN109),.WL(WL51));
sram_cell_6t_5 inst_cell_51_110 (.BL(BL110),.BLN(BLN110),.WL(WL51));
sram_cell_6t_5 inst_cell_51_111 (.BL(BL111),.BLN(BLN111),.WL(WL51));
sram_cell_6t_5 inst_cell_51_112 (.BL(BL112),.BLN(BLN112),.WL(WL51));
sram_cell_6t_5 inst_cell_51_113 (.BL(BL113),.BLN(BLN113),.WL(WL51));
sram_cell_6t_5 inst_cell_51_114 (.BL(BL114),.BLN(BLN114),.WL(WL51));
sram_cell_6t_5 inst_cell_51_115 (.BL(BL115),.BLN(BLN115),.WL(WL51));
sram_cell_6t_5 inst_cell_51_116 (.BL(BL116),.BLN(BLN116),.WL(WL51));
sram_cell_6t_5 inst_cell_51_117 (.BL(BL117),.BLN(BLN117),.WL(WL51));
sram_cell_6t_5 inst_cell_51_118 (.BL(BL118),.BLN(BLN118),.WL(WL51));
sram_cell_6t_5 inst_cell_51_119 (.BL(BL119),.BLN(BLN119),.WL(WL51));
sram_cell_6t_5 inst_cell_51_120 (.BL(BL120),.BLN(BLN120),.WL(WL51));
sram_cell_6t_5 inst_cell_51_121 (.BL(BL121),.BLN(BLN121),.WL(WL51));
sram_cell_6t_5 inst_cell_51_122 (.BL(BL122),.BLN(BLN122),.WL(WL51));
sram_cell_6t_5 inst_cell_51_123 (.BL(BL123),.BLN(BLN123),.WL(WL51));
sram_cell_6t_5 inst_cell_51_124 (.BL(BL124),.BLN(BLN124),.WL(WL51));
sram_cell_6t_5 inst_cell_51_125 (.BL(BL125),.BLN(BLN125),.WL(WL51));
sram_cell_6t_5 inst_cell_51_126 (.BL(BL126),.BLN(BLN126),.WL(WL51));
sram_cell_6t_5 inst_cell_51_127 (.BL(BL127),.BLN(BLN127),.WL(WL51));
sram_cell_6t_5 inst_cell_52_0 (.BL(BL0),.BLN(BLN0),.WL(WL52));
sram_cell_6t_5 inst_cell_52_1 (.BL(BL1),.BLN(BLN1),.WL(WL52));
sram_cell_6t_5 inst_cell_52_2 (.BL(BL2),.BLN(BLN2),.WL(WL52));
sram_cell_6t_5 inst_cell_52_3 (.BL(BL3),.BLN(BLN3),.WL(WL52));
sram_cell_6t_5 inst_cell_52_4 (.BL(BL4),.BLN(BLN4),.WL(WL52));
sram_cell_6t_5 inst_cell_52_5 (.BL(BL5),.BLN(BLN5),.WL(WL52));
sram_cell_6t_5 inst_cell_52_6 (.BL(BL6),.BLN(BLN6),.WL(WL52));
sram_cell_6t_5 inst_cell_52_7 (.BL(BL7),.BLN(BLN7),.WL(WL52));
sram_cell_6t_5 inst_cell_52_8 (.BL(BL8),.BLN(BLN8),.WL(WL52));
sram_cell_6t_5 inst_cell_52_9 (.BL(BL9),.BLN(BLN9),.WL(WL52));
sram_cell_6t_5 inst_cell_52_10 (.BL(BL10),.BLN(BLN10),.WL(WL52));
sram_cell_6t_5 inst_cell_52_11 (.BL(BL11),.BLN(BLN11),.WL(WL52));
sram_cell_6t_5 inst_cell_52_12 (.BL(BL12),.BLN(BLN12),.WL(WL52));
sram_cell_6t_5 inst_cell_52_13 (.BL(BL13),.BLN(BLN13),.WL(WL52));
sram_cell_6t_5 inst_cell_52_14 (.BL(BL14),.BLN(BLN14),.WL(WL52));
sram_cell_6t_5 inst_cell_52_15 (.BL(BL15),.BLN(BLN15),.WL(WL52));
sram_cell_6t_5 inst_cell_52_16 (.BL(BL16),.BLN(BLN16),.WL(WL52));
sram_cell_6t_5 inst_cell_52_17 (.BL(BL17),.BLN(BLN17),.WL(WL52));
sram_cell_6t_5 inst_cell_52_18 (.BL(BL18),.BLN(BLN18),.WL(WL52));
sram_cell_6t_5 inst_cell_52_19 (.BL(BL19),.BLN(BLN19),.WL(WL52));
sram_cell_6t_5 inst_cell_52_20 (.BL(BL20),.BLN(BLN20),.WL(WL52));
sram_cell_6t_5 inst_cell_52_21 (.BL(BL21),.BLN(BLN21),.WL(WL52));
sram_cell_6t_5 inst_cell_52_22 (.BL(BL22),.BLN(BLN22),.WL(WL52));
sram_cell_6t_5 inst_cell_52_23 (.BL(BL23),.BLN(BLN23),.WL(WL52));
sram_cell_6t_5 inst_cell_52_24 (.BL(BL24),.BLN(BLN24),.WL(WL52));
sram_cell_6t_5 inst_cell_52_25 (.BL(BL25),.BLN(BLN25),.WL(WL52));
sram_cell_6t_5 inst_cell_52_26 (.BL(BL26),.BLN(BLN26),.WL(WL52));
sram_cell_6t_5 inst_cell_52_27 (.BL(BL27),.BLN(BLN27),.WL(WL52));
sram_cell_6t_5 inst_cell_52_28 (.BL(BL28),.BLN(BLN28),.WL(WL52));
sram_cell_6t_5 inst_cell_52_29 (.BL(BL29),.BLN(BLN29),.WL(WL52));
sram_cell_6t_5 inst_cell_52_30 (.BL(BL30),.BLN(BLN30),.WL(WL52));
sram_cell_6t_5 inst_cell_52_31 (.BL(BL31),.BLN(BLN31),.WL(WL52));
sram_cell_6t_5 inst_cell_52_32 (.BL(BL32),.BLN(BLN32),.WL(WL52));
sram_cell_6t_5 inst_cell_52_33 (.BL(BL33),.BLN(BLN33),.WL(WL52));
sram_cell_6t_5 inst_cell_52_34 (.BL(BL34),.BLN(BLN34),.WL(WL52));
sram_cell_6t_5 inst_cell_52_35 (.BL(BL35),.BLN(BLN35),.WL(WL52));
sram_cell_6t_5 inst_cell_52_36 (.BL(BL36),.BLN(BLN36),.WL(WL52));
sram_cell_6t_5 inst_cell_52_37 (.BL(BL37),.BLN(BLN37),.WL(WL52));
sram_cell_6t_5 inst_cell_52_38 (.BL(BL38),.BLN(BLN38),.WL(WL52));
sram_cell_6t_5 inst_cell_52_39 (.BL(BL39),.BLN(BLN39),.WL(WL52));
sram_cell_6t_5 inst_cell_52_40 (.BL(BL40),.BLN(BLN40),.WL(WL52));
sram_cell_6t_5 inst_cell_52_41 (.BL(BL41),.BLN(BLN41),.WL(WL52));
sram_cell_6t_5 inst_cell_52_42 (.BL(BL42),.BLN(BLN42),.WL(WL52));
sram_cell_6t_5 inst_cell_52_43 (.BL(BL43),.BLN(BLN43),.WL(WL52));
sram_cell_6t_5 inst_cell_52_44 (.BL(BL44),.BLN(BLN44),.WL(WL52));
sram_cell_6t_5 inst_cell_52_45 (.BL(BL45),.BLN(BLN45),.WL(WL52));
sram_cell_6t_5 inst_cell_52_46 (.BL(BL46),.BLN(BLN46),.WL(WL52));
sram_cell_6t_5 inst_cell_52_47 (.BL(BL47),.BLN(BLN47),.WL(WL52));
sram_cell_6t_5 inst_cell_52_48 (.BL(BL48),.BLN(BLN48),.WL(WL52));
sram_cell_6t_5 inst_cell_52_49 (.BL(BL49),.BLN(BLN49),.WL(WL52));
sram_cell_6t_5 inst_cell_52_50 (.BL(BL50),.BLN(BLN50),.WL(WL52));
sram_cell_6t_5 inst_cell_52_51 (.BL(BL51),.BLN(BLN51),.WL(WL52));
sram_cell_6t_5 inst_cell_52_52 (.BL(BL52),.BLN(BLN52),.WL(WL52));
sram_cell_6t_5 inst_cell_52_53 (.BL(BL53),.BLN(BLN53),.WL(WL52));
sram_cell_6t_5 inst_cell_52_54 (.BL(BL54),.BLN(BLN54),.WL(WL52));
sram_cell_6t_5 inst_cell_52_55 (.BL(BL55),.BLN(BLN55),.WL(WL52));
sram_cell_6t_5 inst_cell_52_56 (.BL(BL56),.BLN(BLN56),.WL(WL52));
sram_cell_6t_5 inst_cell_52_57 (.BL(BL57),.BLN(BLN57),.WL(WL52));
sram_cell_6t_5 inst_cell_52_58 (.BL(BL58),.BLN(BLN58),.WL(WL52));
sram_cell_6t_5 inst_cell_52_59 (.BL(BL59),.BLN(BLN59),.WL(WL52));
sram_cell_6t_5 inst_cell_52_60 (.BL(BL60),.BLN(BLN60),.WL(WL52));
sram_cell_6t_5 inst_cell_52_61 (.BL(BL61),.BLN(BLN61),.WL(WL52));
sram_cell_6t_5 inst_cell_52_62 (.BL(BL62),.BLN(BLN62),.WL(WL52));
sram_cell_6t_5 inst_cell_52_63 (.BL(BL63),.BLN(BLN63),.WL(WL52));
sram_cell_6t_5 inst_cell_52_64 (.BL(BL64),.BLN(BLN64),.WL(WL52));
sram_cell_6t_5 inst_cell_52_65 (.BL(BL65),.BLN(BLN65),.WL(WL52));
sram_cell_6t_5 inst_cell_52_66 (.BL(BL66),.BLN(BLN66),.WL(WL52));
sram_cell_6t_5 inst_cell_52_67 (.BL(BL67),.BLN(BLN67),.WL(WL52));
sram_cell_6t_5 inst_cell_52_68 (.BL(BL68),.BLN(BLN68),.WL(WL52));
sram_cell_6t_5 inst_cell_52_69 (.BL(BL69),.BLN(BLN69),.WL(WL52));
sram_cell_6t_5 inst_cell_52_70 (.BL(BL70),.BLN(BLN70),.WL(WL52));
sram_cell_6t_5 inst_cell_52_71 (.BL(BL71),.BLN(BLN71),.WL(WL52));
sram_cell_6t_5 inst_cell_52_72 (.BL(BL72),.BLN(BLN72),.WL(WL52));
sram_cell_6t_5 inst_cell_52_73 (.BL(BL73),.BLN(BLN73),.WL(WL52));
sram_cell_6t_5 inst_cell_52_74 (.BL(BL74),.BLN(BLN74),.WL(WL52));
sram_cell_6t_5 inst_cell_52_75 (.BL(BL75),.BLN(BLN75),.WL(WL52));
sram_cell_6t_5 inst_cell_52_76 (.BL(BL76),.BLN(BLN76),.WL(WL52));
sram_cell_6t_5 inst_cell_52_77 (.BL(BL77),.BLN(BLN77),.WL(WL52));
sram_cell_6t_5 inst_cell_52_78 (.BL(BL78),.BLN(BLN78),.WL(WL52));
sram_cell_6t_5 inst_cell_52_79 (.BL(BL79),.BLN(BLN79),.WL(WL52));
sram_cell_6t_5 inst_cell_52_80 (.BL(BL80),.BLN(BLN80),.WL(WL52));
sram_cell_6t_5 inst_cell_52_81 (.BL(BL81),.BLN(BLN81),.WL(WL52));
sram_cell_6t_5 inst_cell_52_82 (.BL(BL82),.BLN(BLN82),.WL(WL52));
sram_cell_6t_5 inst_cell_52_83 (.BL(BL83),.BLN(BLN83),.WL(WL52));
sram_cell_6t_5 inst_cell_52_84 (.BL(BL84),.BLN(BLN84),.WL(WL52));
sram_cell_6t_5 inst_cell_52_85 (.BL(BL85),.BLN(BLN85),.WL(WL52));
sram_cell_6t_5 inst_cell_52_86 (.BL(BL86),.BLN(BLN86),.WL(WL52));
sram_cell_6t_5 inst_cell_52_87 (.BL(BL87),.BLN(BLN87),.WL(WL52));
sram_cell_6t_5 inst_cell_52_88 (.BL(BL88),.BLN(BLN88),.WL(WL52));
sram_cell_6t_5 inst_cell_52_89 (.BL(BL89),.BLN(BLN89),.WL(WL52));
sram_cell_6t_5 inst_cell_52_90 (.BL(BL90),.BLN(BLN90),.WL(WL52));
sram_cell_6t_5 inst_cell_52_91 (.BL(BL91),.BLN(BLN91),.WL(WL52));
sram_cell_6t_5 inst_cell_52_92 (.BL(BL92),.BLN(BLN92),.WL(WL52));
sram_cell_6t_5 inst_cell_52_93 (.BL(BL93),.BLN(BLN93),.WL(WL52));
sram_cell_6t_5 inst_cell_52_94 (.BL(BL94),.BLN(BLN94),.WL(WL52));
sram_cell_6t_5 inst_cell_52_95 (.BL(BL95),.BLN(BLN95),.WL(WL52));
sram_cell_6t_5 inst_cell_52_96 (.BL(BL96),.BLN(BLN96),.WL(WL52));
sram_cell_6t_5 inst_cell_52_97 (.BL(BL97),.BLN(BLN97),.WL(WL52));
sram_cell_6t_5 inst_cell_52_98 (.BL(BL98),.BLN(BLN98),.WL(WL52));
sram_cell_6t_5 inst_cell_52_99 (.BL(BL99),.BLN(BLN99),.WL(WL52));
sram_cell_6t_5 inst_cell_52_100 (.BL(BL100),.BLN(BLN100),.WL(WL52));
sram_cell_6t_5 inst_cell_52_101 (.BL(BL101),.BLN(BLN101),.WL(WL52));
sram_cell_6t_5 inst_cell_52_102 (.BL(BL102),.BLN(BLN102),.WL(WL52));
sram_cell_6t_5 inst_cell_52_103 (.BL(BL103),.BLN(BLN103),.WL(WL52));
sram_cell_6t_5 inst_cell_52_104 (.BL(BL104),.BLN(BLN104),.WL(WL52));
sram_cell_6t_5 inst_cell_52_105 (.BL(BL105),.BLN(BLN105),.WL(WL52));
sram_cell_6t_5 inst_cell_52_106 (.BL(BL106),.BLN(BLN106),.WL(WL52));
sram_cell_6t_5 inst_cell_52_107 (.BL(BL107),.BLN(BLN107),.WL(WL52));
sram_cell_6t_5 inst_cell_52_108 (.BL(BL108),.BLN(BLN108),.WL(WL52));
sram_cell_6t_5 inst_cell_52_109 (.BL(BL109),.BLN(BLN109),.WL(WL52));
sram_cell_6t_5 inst_cell_52_110 (.BL(BL110),.BLN(BLN110),.WL(WL52));
sram_cell_6t_5 inst_cell_52_111 (.BL(BL111),.BLN(BLN111),.WL(WL52));
sram_cell_6t_5 inst_cell_52_112 (.BL(BL112),.BLN(BLN112),.WL(WL52));
sram_cell_6t_5 inst_cell_52_113 (.BL(BL113),.BLN(BLN113),.WL(WL52));
sram_cell_6t_5 inst_cell_52_114 (.BL(BL114),.BLN(BLN114),.WL(WL52));
sram_cell_6t_5 inst_cell_52_115 (.BL(BL115),.BLN(BLN115),.WL(WL52));
sram_cell_6t_5 inst_cell_52_116 (.BL(BL116),.BLN(BLN116),.WL(WL52));
sram_cell_6t_5 inst_cell_52_117 (.BL(BL117),.BLN(BLN117),.WL(WL52));
sram_cell_6t_5 inst_cell_52_118 (.BL(BL118),.BLN(BLN118),.WL(WL52));
sram_cell_6t_5 inst_cell_52_119 (.BL(BL119),.BLN(BLN119),.WL(WL52));
sram_cell_6t_5 inst_cell_52_120 (.BL(BL120),.BLN(BLN120),.WL(WL52));
sram_cell_6t_5 inst_cell_52_121 (.BL(BL121),.BLN(BLN121),.WL(WL52));
sram_cell_6t_5 inst_cell_52_122 (.BL(BL122),.BLN(BLN122),.WL(WL52));
sram_cell_6t_5 inst_cell_52_123 (.BL(BL123),.BLN(BLN123),.WL(WL52));
sram_cell_6t_5 inst_cell_52_124 (.BL(BL124),.BLN(BLN124),.WL(WL52));
sram_cell_6t_5 inst_cell_52_125 (.BL(BL125),.BLN(BLN125),.WL(WL52));
sram_cell_6t_5 inst_cell_52_126 (.BL(BL126),.BLN(BLN126),.WL(WL52));
sram_cell_6t_5 inst_cell_52_127 (.BL(BL127),.BLN(BLN127),.WL(WL52));
sram_cell_6t_5 inst_cell_53_0 (.BL(BL0),.BLN(BLN0),.WL(WL53));
sram_cell_6t_5 inst_cell_53_1 (.BL(BL1),.BLN(BLN1),.WL(WL53));
sram_cell_6t_5 inst_cell_53_2 (.BL(BL2),.BLN(BLN2),.WL(WL53));
sram_cell_6t_5 inst_cell_53_3 (.BL(BL3),.BLN(BLN3),.WL(WL53));
sram_cell_6t_5 inst_cell_53_4 (.BL(BL4),.BLN(BLN4),.WL(WL53));
sram_cell_6t_5 inst_cell_53_5 (.BL(BL5),.BLN(BLN5),.WL(WL53));
sram_cell_6t_5 inst_cell_53_6 (.BL(BL6),.BLN(BLN6),.WL(WL53));
sram_cell_6t_5 inst_cell_53_7 (.BL(BL7),.BLN(BLN7),.WL(WL53));
sram_cell_6t_5 inst_cell_53_8 (.BL(BL8),.BLN(BLN8),.WL(WL53));
sram_cell_6t_5 inst_cell_53_9 (.BL(BL9),.BLN(BLN9),.WL(WL53));
sram_cell_6t_5 inst_cell_53_10 (.BL(BL10),.BLN(BLN10),.WL(WL53));
sram_cell_6t_5 inst_cell_53_11 (.BL(BL11),.BLN(BLN11),.WL(WL53));
sram_cell_6t_5 inst_cell_53_12 (.BL(BL12),.BLN(BLN12),.WL(WL53));
sram_cell_6t_5 inst_cell_53_13 (.BL(BL13),.BLN(BLN13),.WL(WL53));
sram_cell_6t_5 inst_cell_53_14 (.BL(BL14),.BLN(BLN14),.WL(WL53));
sram_cell_6t_5 inst_cell_53_15 (.BL(BL15),.BLN(BLN15),.WL(WL53));
sram_cell_6t_5 inst_cell_53_16 (.BL(BL16),.BLN(BLN16),.WL(WL53));
sram_cell_6t_5 inst_cell_53_17 (.BL(BL17),.BLN(BLN17),.WL(WL53));
sram_cell_6t_5 inst_cell_53_18 (.BL(BL18),.BLN(BLN18),.WL(WL53));
sram_cell_6t_5 inst_cell_53_19 (.BL(BL19),.BLN(BLN19),.WL(WL53));
sram_cell_6t_5 inst_cell_53_20 (.BL(BL20),.BLN(BLN20),.WL(WL53));
sram_cell_6t_5 inst_cell_53_21 (.BL(BL21),.BLN(BLN21),.WL(WL53));
sram_cell_6t_5 inst_cell_53_22 (.BL(BL22),.BLN(BLN22),.WL(WL53));
sram_cell_6t_5 inst_cell_53_23 (.BL(BL23),.BLN(BLN23),.WL(WL53));
sram_cell_6t_5 inst_cell_53_24 (.BL(BL24),.BLN(BLN24),.WL(WL53));
sram_cell_6t_5 inst_cell_53_25 (.BL(BL25),.BLN(BLN25),.WL(WL53));
sram_cell_6t_5 inst_cell_53_26 (.BL(BL26),.BLN(BLN26),.WL(WL53));
sram_cell_6t_5 inst_cell_53_27 (.BL(BL27),.BLN(BLN27),.WL(WL53));
sram_cell_6t_5 inst_cell_53_28 (.BL(BL28),.BLN(BLN28),.WL(WL53));
sram_cell_6t_5 inst_cell_53_29 (.BL(BL29),.BLN(BLN29),.WL(WL53));
sram_cell_6t_5 inst_cell_53_30 (.BL(BL30),.BLN(BLN30),.WL(WL53));
sram_cell_6t_5 inst_cell_53_31 (.BL(BL31),.BLN(BLN31),.WL(WL53));
sram_cell_6t_5 inst_cell_53_32 (.BL(BL32),.BLN(BLN32),.WL(WL53));
sram_cell_6t_5 inst_cell_53_33 (.BL(BL33),.BLN(BLN33),.WL(WL53));
sram_cell_6t_5 inst_cell_53_34 (.BL(BL34),.BLN(BLN34),.WL(WL53));
sram_cell_6t_5 inst_cell_53_35 (.BL(BL35),.BLN(BLN35),.WL(WL53));
sram_cell_6t_5 inst_cell_53_36 (.BL(BL36),.BLN(BLN36),.WL(WL53));
sram_cell_6t_5 inst_cell_53_37 (.BL(BL37),.BLN(BLN37),.WL(WL53));
sram_cell_6t_5 inst_cell_53_38 (.BL(BL38),.BLN(BLN38),.WL(WL53));
sram_cell_6t_5 inst_cell_53_39 (.BL(BL39),.BLN(BLN39),.WL(WL53));
sram_cell_6t_5 inst_cell_53_40 (.BL(BL40),.BLN(BLN40),.WL(WL53));
sram_cell_6t_5 inst_cell_53_41 (.BL(BL41),.BLN(BLN41),.WL(WL53));
sram_cell_6t_5 inst_cell_53_42 (.BL(BL42),.BLN(BLN42),.WL(WL53));
sram_cell_6t_5 inst_cell_53_43 (.BL(BL43),.BLN(BLN43),.WL(WL53));
sram_cell_6t_5 inst_cell_53_44 (.BL(BL44),.BLN(BLN44),.WL(WL53));
sram_cell_6t_5 inst_cell_53_45 (.BL(BL45),.BLN(BLN45),.WL(WL53));
sram_cell_6t_5 inst_cell_53_46 (.BL(BL46),.BLN(BLN46),.WL(WL53));
sram_cell_6t_5 inst_cell_53_47 (.BL(BL47),.BLN(BLN47),.WL(WL53));
sram_cell_6t_5 inst_cell_53_48 (.BL(BL48),.BLN(BLN48),.WL(WL53));
sram_cell_6t_5 inst_cell_53_49 (.BL(BL49),.BLN(BLN49),.WL(WL53));
sram_cell_6t_5 inst_cell_53_50 (.BL(BL50),.BLN(BLN50),.WL(WL53));
sram_cell_6t_5 inst_cell_53_51 (.BL(BL51),.BLN(BLN51),.WL(WL53));
sram_cell_6t_5 inst_cell_53_52 (.BL(BL52),.BLN(BLN52),.WL(WL53));
sram_cell_6t_5 inst_cell_53_53 (.BL(BL53),.BLN(BLN53),.WL(WL53));
sram_cell_6t_5 inst_cell_53_54 (.BL(BL54),.BLN(BLN54),.WL(WL53));
sram_cell_6t_5 inst_cell_53_55 (.BL(BL55),.BLN(BLN55),.WL(WL53));
sram_cell_6t_5 inst_cell_53_56 (.BL(BL56),.BLN(BLN56),.WL(WL53));
sram_cell_6t_5 inst_cell_53_57 (.BL(BL57),.BLN(BLN57),.WL(WL53));
sram_cell_6t_5 inst_cell_53_58 (.BL(BL58),.BLN(BLN58),.WL(WL53));
sram_cell_6t_5 inst_cell_53_59 (.BL(BL59),.BLN(BLN59),.WL(WL53));
sram_cell_6t_5 inst_cell_53_60 (.BL(BL60),.BLN(BLN60),.WL(WL53));
sram_cell_6t_5 inst_cell_53_61 (.BL(BL61),.BLN(BLN61),.WL(WL53));
sram_cell_6t_5 inst_cell_53_62 (.BL(BL62),.BLN(BLN62),.WL(WL53));
sram_cell_6t_5 inst_cell_53_63 (.BL(BL63),.BLN(BLN63),.WL(WL53));
sram_cell_6t_5 inst_cell_53_64 (.BL(BL64),.BLN(BLN64),.WL(WL53));
sram_cell_6t_5 inst_cell_53_65 (.BL(BL65),.BLN(BLN65),.WL(WL53));
sram_cell_6t_5 inst_cell_53_66 (.BL(BL66),.BLN(BLN66),.WL(WL53));
sram_cell_6t_5 inst_cell_53_67 (.BL(BL67),.BLN(BLN67),.WL(WL53));
sram_cell_6t_5 inst_cell_53_68 (.BL(BL68),.BLN(BLN68),.WL(WL53));
sram_cell_6t_5 inst_cell_53_69 (.BL(BL69),.BLN(BLN69),.WL(WL53));
sram_cell_6t_5 inst_cell_53_70 (.BL(BL70),.BLN(BLN70),.WL(WL53));
sram_cell_6t_5 inst_cell_53_71 (.BL(BL71),.BLN(BLN71),.WL(WL53));
sram_cell_6t_5 inst_cell_53_72 (.BL(BL72),.BLN(BLN72),.WL(WL53));
sram_cell_6t_5 inst_cell_53_73 (.BL(BL73),.BLN(BLN73),.WL(WL53));
sram_cell_6t_5 inst_cell_53_74 (.BL(BL74),.BLN(BLN74),.WL(WL53));
sram_cell_6t_5 inst_cell_53_75 (.BL(BL75),.BLN(BLN75),.WL(WL53));
sram_cell_6t_5 inst_cell_53_76 (.BL(BL76),.BLN(BLN76),.WL(WL53));
sram_cell_6t_5 inst_cell_53_77 (.BL(BL77),.BLN(BLN77),.WL(WL53));
sram_cell_6t_5 inst_cell_53_78 (.BL(BL78),.BLN(BLN78),.WL(WL53));
sram_cell_6t_5 inst_cell_53_79 (.BL(BL79),.BLN(BLN79),.WL(WL53));
sram_cell_6t_5 inst_cell_53_80 (.BL(BL80),.BLN(BLN80),.WL(WL53));
sram_cell_6t_5 inst_cell_53_81 (.BL(BL81),.BLN(BLN81),.WL(WL53));
sram_cell_6t_5 inst_cell_53_82 (.BL(BL82),.BLN(BLN82),.WL(WL53));
sram_cell_6t_5 inst_cell_53_83 (.BL(BL83),.BLN(BLN83),.WL(WL53));
sram_cell_6t_5 inst_cell_53_84 (.BL(BL84),.BLN(BLN84),.WL(WL53));
sram_cell_6t_5 inst_cell_53_85 (.BL(BL85),.BLN(BLN85),.WL(WL53));
sram_cell_6t_5 inst_cell_53_86 (.BL(BL86),.BLN(BLN86),.WL(WL53));
sram_cell_6t_5 inst_cell_53_87 (.BL(BL87),.BLN(BLN87),.WL(WL53));
sram_cell_6t_5 inst_cell_53_88 (.BL(BL88),.BLN(BLN88),.WL(WL53));
sram_cell_6t_5 inst_cell_53_89 (.BL(BL89),.BLN(BLN89),.WL(WL53));
sram_cell_6t_5 inst_cell_53_90 (.BL(BL90),.BLN(BLN90),.WL(WL53));
sram_cell_6t_5 inst_cell_53_91 (.BL(BL91),.BLN(BLN91),.WL(WL53));
sram_cell_6t_5 inst_cell_53_92 (.BL(BL92),.BLN(BLN92),.WL(WL53));
sram_cell_6t_5 inst_cell_53_93 (.BL(BL93),.BLN(BLN93),.WL(WL53));
sram_cell_6t_5 inst_cell_53_94 (.BL(BL94),.BLN(BLN94),.WL(WL53));
sram_cell_6t_5 inst_cell_53_95 (.BL(BL95),.BLN(BLN95),.WL(WL53));
sram_cell_6t_5 inst_cell_53_96 (.BL(BL96),.BLN(BLN96),.WL(WL53));
sram_cell_6t_5 inst_cell_53_97 (.BL(BL97),.BLN(BLN97),.WL(WL53));
sram_cell_6t_5 inst_cell_53_98 (.BL(BL98),.BLN(BLN98),.WL(WL53));
sram_cell_6t_5 inst_cell_53_99 (.BL(BL99),.BLN(BLN99),.WL(WL53));
sram_cell_6t_5 inst_cell_53_100 (.BL(BL100),.BLN(BLN100),.WL(WL53));
sram_cell_6t_5 inst_cell_53_101 (.BL(BL101),.BLN(BLN101),.WL(WL53));
sram_cell_6t_5 inst_cell_53_102 (.BL(BL102),.BLN(BLN102),.WL(WL53));
sram_cell_6t_5 inst_cell_53_103 (.BL(BL103),.BLN(BLN103),.WL(WL53));
sram_cell_6t_5 inst_cell_53_104 (.BL(BL104),.BLN(BLN104),.WL(WL53));
sram_cell_6t_5 inst_cell_53_105 (.BL(BL105),.BLN(BLN105),.WL(WL53));
sram_cell_6t_5 inst_cell_53_106 (.BL(BL106),.BLN(BLN106),.WL(WL53));
sram_cell_6t_5 inst_cell_53_107 (.BL(BL107),.BLN(BLN107),.WL(WL53));
sram_cell_6t_5 inst_cell_53_108 (.BL(BL108),.BLN(BLN108),.WL(WL53));
sram_cell_6t_5 inst_cell_53_109 (.BL(BL109),.BLN(BLN109),.WL(WL53));
sram_cell_6t_5 inst_cell_53_110 (.BL(BL110),.BLN(BLN110),.WL(WL53));
sram_cell_6t_5 inst_cell_53_111 (.BL(BL111),.BLN(BLN111),.WL(WL53));
sram_cell_6t_5 inst_cell_53_112 (.BL(BL112),.BLN(BLN112),.WL(WL53));
sram_cell_6t_5 inst_cell_53_113 (.BL(BL113),.BLN(BLN113),.WL(WL53));
sram_cell_6t_5 inst_cell_53_114 (.BL(BL114),.BLN(BLN114),.WL(WL53));
sram_cell_6t_5 inst_cell_53_115 (.BL(BL115),.BLN(BLN115),.WL(WL53));
sram_cell_6t_5 inst_cell_53_116 (.BL(BL116),.BLN(BLN116),.WL(WL53));
sram_cell_6t_5 inst_cell_53_117 (.BL(BL117),.BLN(BLN117),.WL(WL53));
sram_cell_6t_5 inst_cell_53_118 (.BL(BL118),.BLN(BLN118),.WL(WL53));
sram_cell_6t_5 inst_cell_53_119 (.BL(BL119),.BLN(BLN119),.WL(WL53));
sram_cell_6t_5 inst_cell_53_120 (.BL(BL120),.BLN(BLN120),.WL(WL53));
sram_cell_6t_5 inst_cell_53_121 (.BL(BL121),.BLN(BLN121),.WL(WL53));
sram_cell_6t_5 inst_cell_53_122 (.BL(BL122),.BLN(BLN122),.WL(WL53));
sram_cell_6t_5 inst_cell_53_123 (.BL(BL123),.BLN(BLN123),.WL(WL53));
sram_cell_6t_5 inst_cell_53_124 (.BL(BL124),.BLN(BLN124),.WL(WL53));
sram_cell_6t_5 inst_cell_53_125 (.BL(BL125),.BLN(BLN125),.WL(WL53));
sram_cell_6t_5 inst_cell_53_126 (.BL(BL126),.BLN(BLN126),.WL(WL53));
sram_cell_6t_5 inst_cell_53_127 (.BL(BL127),.BLN(BLN127),.WL(WL53));
sram_cell_6t_5 inst_cell_54_0 (.BL(BL0),.BLN(BLN0),.WL(WL54));
sram_cell_6t_5 inst_cell_54_1 (.BL(BL1),.BLN(BLN1),.WL(WL54));
sram_cell_6t_5 inst_cell_54_2 (.BL(BL2),.BLN(BLN2),.WL(WL54));
sram_cell_6t_5 inst_cell_54_3 (.BL(BL3),.BLN(BLN3),.WL(WL54));
sram_cell_6t_5 inst_cell_54_4 (.BL(BL4),.BLN(BLN4),.WL(WL54));
sram_cell_6t_5 inst_cell_54_5 (.BL(BL5),.BLN(BLN5),.WL(WL54));
sram_cell_6t_5 inst_cell_54_6 (.BL(BL6),.BLN(BLN6),.WL(WL54));
sram_cell_6t_5 inst_cell_54_7 (.BL(BL7),.BLN(BLN7),.WL(WL54));
sram_cell_6t_5 inst_cell_54_8 (.BL(BL8),.BLN(BLN8),.WL(WL54));
sram_cell_6t_5 inst_cell_54_9 (.BL(BL9),.BLN(BLN9),.WL(WL54));
sram_cell_6t_5 inst_cell_54_10 (.BL(BL10),.BLN(BLN10),.WL(WL54));
sram_cell_6t_5 inst_cell_54_11 (.BL(BL11),.BLN(BLN11),.WL(WL54));
sram_cell_6t_5 inst_cell_54_12 (.BL(BL12),.BLN(BLN12),.WL(WL54));
sram_cell_6t_5 inst_cell_54_13 (.BL(BL13),.BLN(BLN13),.WL(WL54));
sram_cell_6t_5 inst_cell_54_14 (.BL(BL14),.BLN(BLN14),.WL(WL54));
sram_cell_6t_5 inst_cell_54_15 (.BL(BL15),.BLN(BLN15),.WL(WL54));
sram_cell_6t_5 inst_cell_54_16 (.BL(BL16),.BLN(BLN16),.WL(WL54));
sram_cell_6t_5 inst_cell_54_17 (.BL(BL17),.BLN(BLN17),.WL(WL54));
sram_cell_6t_5 inst_cell_54_18 (.BL(BL18),.BLN(BLN18),.WL(WL54));
sram_cell_6t_5 inst_cell_54_19 (.BL(BL19),.BLN(BLN19),.WL(WL54));
sram_cell_6t_5 inst_cell_54_20 (.BL(BL20),.BLN(BLN20),.WL(WL54));
sram_cell_6t_5 inst_cell_54_21 (.BL(BL21),.BLN(BLN21),.WL(WL54));
sram_cell_6t_5 inst_cell_54_22 (.BL(BL22),.BLN(BLN22),.WL(WL54));
sram_cell_6t_5 inst_cell_54_23 (.BL(BL23),.BLN(BLN23),.WL(WL54));
sram_cell_6t_5 inst_cell_54_24 (.BL(BL24),.BLN(BLN24),.WL(WL54));
sram_cell_6t_5 inst_cell_54_25 (.BL(BL25),.BLN(BLN25),.WL(WL54));
sram_cell_6t_5 inst_cell_54_26 (.BL(BL26),.BLN(BLN26),.WL(WL54));
sram_cell_6t_5 inst_cell_54_27 (.BL(BL27),.BLN(BLN27),.WL(WL54));
sram_cell_6t_5 inst_cell_54_28 (.BL(BL28),.BLN(BLN28),.WL(WL54));
sram_cell_6t_5 inst_cell_54_29 (.BL(BL29),.BLN(BLN29),.WL(WL54));
sram_cell_6t_5 inst_cell_54_30 (.BL(BL30),.BLN(BLN30),.WL(WL54));
sram_cell_6t_5 inst_cell_54_31 (.BL(BL31),.BLN(BLN31),.WL(WL54));
sram_cell_6t_5 inst_cell_54_32 (.BL(BL32),.BLN(BLN32),.WL(WL54));
sram_cell_6t_5 inst_cell_54_33 (.BL(BL33),.BLN(BLN33),.WL(WL54));
sram_cell_6t_5 inst_cell_54_34 (.BL(BL34),.BLN(BLN34),.WL(WL54));
sram_cell_6t_5 inst_cell_54_35 (.BL(BL35),.BLN(BLN35),.WL(WL54));
sram_cell_6t_5 inst_cell_54_36 (.BL(BL36),.BLN(BLN36),.WL(WL54));
sram_cell_6t_5 inst_cell_54_37 (.BL(BL37),.BLN(BLN37),.WL(WL54));
sram_cell_6t_5 inst_cell_54_38 (.BL(BL38),.BLN(BLN38),.WL(WL54));
sram_cell_6t_5 inst_cell_54_39 (.BL(BL39),.BLN(BLN39),.WL(WL54));
sram_cell_6t_5 inst_cell_54_40 (.BL(BL40),.BLN(BLN40),.WL(WL54));
sram_cell_6t_5 inst_cell_54_41 (.BL(BL41),.BLN(BLN41),.WL(WL54));
sram_cell_6t_5 inst_cell_54_42 (.BL(BL42),.BLN(BLN42),.WL(WL54));
sram_cell_6t_5 inst_cell_54_43 (.BL(BL43),.BLN(BLN43),.WL(WL54));
sram_cell_6t_5 inst_cell_54_44 (.BL(BL44),.BLN(BLN44),.WL(WL54));
sram_cell_6t_5 inst_cell_54_45 (.BL(BL45),.BLN(BLN45),.WL(WL54));
sram_cell_6t_5 inst_cell_54_46 (.BL(BL46),.BLN(BLN46),.WL(WL54));
sram_cell_6t_5 inst_cell_54_47 (.BL(BL47),.BLN(BLN47),.WL(WL54));
sram_cell_6t_5 inst_cell_54_48 (.BL(BL48),.BLN(BLN48),.WL(WL54));
sram_cell_6t_5 inst_cell_54_49 (.BL(BL49),.BLN(BLN49),.WL(WL54));
sram_cell_6t_5 inst_cell_54_50 (.BL(BL50),.BLN(BLN50),.WL(WL54));
sram_cell_6t_5 inst_cell_54_51 (.BL(BL51),.BLN(BLN51),.WL(WL54));
sram_cell_6t_5 inst_cell_54_52 (.BL(BL52),.BLN(BLN52),.WL(WL54));
sram_cell_6t_5 inst_cell_54_53 (.BL(BL53),.BLN(BLN53),.WL(WL54));
sram_cell_6t_5 inst_cell_54_54 (.BL(BL54),.BLN(BLN54),.WL(WL54));
sram_cell_6t_5 inst_cell_54_55 (.BL(BL55),.BLN(BLN55),.WL(WL54));
sram_cell_6t_5 inst_cell_54_56 (.BL(BL56),.BLN(BLN56),.WL(WL54));
sram_cell_6t_5 inst_cell_54_57 (.BL(BL57),.BLN(BLN57),.WL(WL54));
sram_cell_6t_5 inst_cell_54_58 (.BL(BL58),.BLN(BLN58),.WL(WL54));
sram_cell_6t_5 inst_cell_54_59 (.BL(BL59),.BLN(BLN59),.WL(WL54));
sram_cell_6t_5 inst_cell_54_60 (.BL(BL60),.BLN(BLN60),.WL(WL54));
sram_cell_6t_5 inst_cell_54_61 (.BL(BL61),.BLN(BLN61),.WL(WL54));
sram_cell_6t_5 inst_cell_54_62 (.BL(BL62),.BLN(BLN62),.WL(WL54));
sram_cell_6t_5 inst_cell_54_63 (.BL(BL63),.BLN(BLN63),.WL(WL54));
sram_cell_6t_5 inst_cell_54_64 (.BL(BL64),.BLN(BLN64),.WL(WL54));
sram_cell_6t_5 inst_cell_54_65 (.BL(BL65),.BLN(BLN65),.WL(WL54));
sram_cell_6t_5 inst_cell_54_66 (.BL(BL66),.BLN(BLN66),.WL(WL54));
sram_cell_6t_5 inst_cell_54_67 (.BL(BL67),.BLN(BLN67),.WL(WL54));
sram_cell_6t_5 inst_cell_54_68 (.BL(BL68),.BLN(BLN68),.WL(WL54));
sram_cell_6t_5 inst_cell_54_69 (.BL(BL69),.BLN(BLN69),.WL(WL54));
sram_cell_6t_5 inst_cell_54_70 (.BL(BL70),.BLN(BLN70),.WL(WL54));
sram_cell_6t_5 inst_cell_54_71 (.BL(BL71),.BLN(BLN71),.WL(WL54));
sram_cell_6t_5 inst_cell_54_72 (.BL(BL72),.BLN(BLN72),.WL(WL54));
sram_cell_6t_5 inst_cell_54_73 (.BL(BL73),.BLN(BLN73),.WL(WL54));
sram_cell_6t_5 inst_cell_54_74 (.BL(BL74),.BLN(BLN74),.WL(WL54));
sram_cell_6t_5 inst_cell_54_75 (.BL(BL75),.BLN(BLN75),.WL(WL54));
sram_cell_6t_5 inst_cell_54_76 (.BL(BL76),.BLN(BLN76),.WL(WL54));
sram_cell_6t_5 inst_cell_54_77 (.BL(BL77),.BLN(BLN77),.WL(WL54));
sram_cell_6t_5 inst_cell_54_78 (.BL(BL78),.BLN(BLN78),.WL(WL54));
sram_cell_6t_5 inst_cell_54_79 (.BL(BL79),.BLN(BLN79),.WL(WL54));
sram_cell_6t_5 inst_cell_54_80 (.BL(BL80),.BLN(BLN80),.WL(WL54));
sram_cell_6t_5 inst_cell_54_81 (.BL(BL81),.BLN(BLN81),.WL(WL54));
sram_cell_6t_5 inst_cell_54_82 (.BL(BL82),.BLN(BLN82),.WL(WL54));
sram_cell_6t_5 inst_cell_54_83 (.BL(BL83),.BLN(BLN83),.WL(WL54));
sram_cell_6t_5 inst_cell_54_84 (.BL(BL84),.BLN(BLN84),.WL(WL54));
sram_cell_6t_5 inst_cell_54_85 (.BL(BL85),.BLN(BLN85),.WL(WL54));
sram_cell_6t_5 inst_cell_54_86 (.BL(BL86),.BLN(BLN86),.WL(WL54));
sram_cell_6t_5 inst_cell_54_87 (.BL(BL87),.BLN(BLN87),.WL(WL54));
sram_cell_6t_5 inst_cell_54_88 (.BL(BL88),.BLN(BLN88),.WL(WL54));
sram_cell_6t_5 inst_cell_54_89 (.BL(BL89),.BLN(BLN89),.WL(WL54));
sram_cell_6t_5 inst_cell_54_90 (.BL(BL90),.BLN(BLN90),.WL(WL54));
sram_cell_6t_5 inst_cell_54_91 (.BL(BL91),.BLN(BLN91),.WL(WL54));
sram_cell_6t_5 inst_cell_54_92 (.BL(BL92),.BLN(BLN92),.WL(WL54));
sram_cell_6t_5 inst_cell_54_93 (.BL(BL93),.BLN(BLN93),.WL(WL54));
sram_cell_6t_5 inst_cell_54_94 (.BL(BL94),.BLN(BLN94),.WL(WL54));
sram_cell_6t_5 inst_cell_54_95 (.BL(BL95),.BLN(BLN95),.WL(WL54));
sram_cell_6t_5 inst_cell_54_96 (.BL(BL96),.BLN(BLN96),.WL(WL54));
sram_cell_6t_5 inst_cell_54_97 (.BL(BL97),.BLN(BLN97),.WL(WL54));
sram_cell_6t_5 inst_cell_54_98 (.BL(BL98),.BLN(BLN98),.WL(WL54));
sram_cell_6t_5 inst_cell_54_99 (.BL(BL99),.BLN(BLN99),.WL(WL54));
sram_cell_6t_5 inst_cell_54_100 (.BL(BL100),.BLN(BLN100),.WL(WL54));
sram_cell_6t_5 inst_cell_54_101 (.BL(BL101),.BLN(BLN101),.WL(WL54));
sram_cell_6t_5 inst_cell_54_102 (.BL(BL102),.BLN(BLN102),.WL(WL54));
sram_cell_6t_5 inst_cell_54_103 (.BL(BL103),.BLN(BLN103),.WL(WL54));
sram_cell_6t_5 inst_cell_54_104 (.BL(BL104),.BLN(BLN104),.WL(WL54));
sram_cell_6t_5 inst_cell_54_105 (.BL(BL105),.BLN(BLN105),.WL(WL54));
sram_cell_6t_5 inst_cell_54_106 (.BL(BL106),.BLN(BLN106),.WL(WL54));
sram_cell_6t_5 inst_cell_54_107 (.BL(BL107),.BLN(BLN107),.WL(WL54));
sram_cell_6t_5 inst_cell_54_108 (.BL(BL108),.BLN(BLN108),.WL(WL54));
sram_cell_6t_5 inst_cell_54_109 (.BL(BL109),.BLN(BLN109),.WL(WL54));
sram_cell_6t_5 inst_cell_54_110 (.BL(BL110),.BLN(BLN110),.WL(WL54));
sram_cell_6t_5 inst_cell_54_111 (.BL(BL111),.BLN(BLN111),.WL(WL54));
sram_cell_6t_5 inst_cell_54_112 (.BL(BL112),.BLN(BLN112),.WL(WL54));
sram_cell_6t_5 inst_cell_54_113 (.BL(BL113),.BLN(BLN113),.WL(WL54));
sram_cell_6t_5 inst_cell_54_114 (.BL(BL114),.BLN(BLN114),.WL(WL54));
sram_cell_6t_5 inst_cell_54_115 (.BL(BL115),.BLN(BLN115),.WL(WL54));
sram_cell_6t_5 inst_cell_54_116 (.BL(BL116),.BLN(BLN116),.WL(WL54));
sram_cell_6t_5 inst_cell_54_117 (.BL(BL117),.BLN(BLN117),.WL(WL54));
sram_cell_6t_5 inst_cell_54_118 (.BL(BL118),.BLN(BLN118),.WL(WL54));
sram_cell_6t_5 inst_cell_54_119 (.BL(BL119),.BLN(BLN119),.WL(WL54));
sram_cell_6t_5 inst_cell_54_120 (.BL(BL120),.BLN(BLN120),.WL(WL54));
sram_cell_6t_5 inst_cell_54_121 (.BL(BL121),.BLN(BLN121),.WL(WL54));
sram_cell_6t_5 inst_cell_54_122 (.BL(BL122),.BLN(BLN122),.WL(WL54));
sram_cell_6t_5 inst_cell_54_123 (.BL(BL123),.BLN(BLN123),.WL(WL54));
sram_cell_6t_5 inst_cell_54_124 (.BL(BL124),.BLN(BLN124),.WL(WL54));
sram_cell_6t_5 inst_cell_54_125 (.BL(BL125),.BLN(BLN125),.WL(WL54));
sram_cell_6t_5 inst_cell_54_126 (.BL(BL126),.BLN(BLN126),.WL(WL54));
sram_cell_6t_5 inst_cell_54_127 (.BL(BL127),.BLN(BLN127),.WL(WL54));
sram_cell_6t_5 inst_cell_55_0 (.BL(BL0),.BLN(BLN0),.WL(WL55));
sram_cell_6t_5 inst_cell_55_1 (.BL(BL1),.BLN(BLN1),.WL(WL55));
sram_cell_6t_5 inst_cell_55_2 (.BL(BL2),.BLN(BLN2),.WL(WL55));
sram_cell_6t_5 inst_cell_55_3 (.BL(BL3),.BLN(BLN3),.WL(WL55));
sram_cell_6t_5 inst_cell_55_4 (.BL(BL4),.BLN(BLN4),.WL(WL55));
sram_cell_6t_5 inst_cell_55_5 (.BL(BL5),.BLN(BLN5),.WL(WL55));
sram_cell_6t_5 inst_cell_55_6 (.BL(BL6),.BLN(BLN6),.WL(WL55));
sram_cell_6t_5 inst_cell_55_7 (.BL(BL7),.BLN(BLN7),.WL(WL55));
sram_cell_6t_5 inst_cell_55_8 (.BL(BL8),.BLN(BLN8),.WL(WL55));
sram_cell_6t_5 inst_cell_55_9 (.BL(BL9),.BLN(BLN9),.WL(WL55));
sram_cell_6t_5 inst_cell_55_10 (.BL(BL10),.BLN(BLN10),.WL(WL55));
sram_cell_6t_5 inst_cell_55_11 (.BL(BL11),.BLN(BLN11),.WL(WL55));
sram_cell_6t_5 inst_cell_55_12 (.BL(BL12),.BLN(BLN12),.WL(WL55));
sram_cell_6t_5 inst_cell_55_13 (.BL(BL13),.BLN(BLN13),.WL(WL55));
sram_cell_6t_5 inst_cell_55_14 (.BL(BL14),.BLN(BLN14),.WL(WL55));
sram_cell_6t_5 inst_cell_55_15 (.BL(BL15),.BLN(BLN15),.WL(WL55));
sram_cell_6t_5 inst_cell_55_16 (.BL(BL16),.BLN(BLN16),.WL(WL55));
sram_cell_6t_5 inst_cell_55_17 (.BL(BL17),.BLN(BLN17),.WL(WL55));
sram_cell_6t_5 inst_cell_55_18 (.BL(BL18),.BLN(BLN18),.WL(WL55));
sram_cell_6t_5 inst_cell_55_19 (.BL(BL19),.BLN(BLN19),.WL(WL55));
sram_cell_6t_5 inst_cell_55_20 (.BL(BL20),.BLN(BLN20),.WL(WL55));
sram_cell_6t_5 inst_cell_55_21 (.BL(BL21),.BLN(BLN21),.WL(WL55));
sram_cell_6t_5 inst_cell_55_22 (.BL(BL22),.BLN(BLN22),.WL(WL55));
sram_cell_6t_5 inst_cell_55_23 (.BL(BL23),.BLN(BLN23),.WL(WL55));
sram_cell_6t_5 inst_cell_55_24 (.BL(BL24),.BLN(BLN24),.WL(WL55));
sram_cell_6t_5 inst_cell_55_25 (.BL(BL25),.BLN(BLN25),.WL(WL55));
sram_cell_6t_5 inst_cell_55_26 (.BL(BL26),.BLN(BLN26),.WL(WL55));
sram_cell_6t_5 inst_cell_55_27 (.BL(BL27),.BLN(BLN27),.WL(WL55));
sram_cell_6t_5 inst_cell_55_28 (.BL(BL28),.BLN(BLN28),.WL(WL55));
sram_cell_6t_5 inst_cell_55_29 (.BL(BL29),.BLN(BLN29),.WL(WL55));
sram_cell_6t_5 inst_cell_55_30 (.BL(BL30),.BLN(BLN30),.WL(WL55));
sram_cell_6t_5 inst_cell_55_31 (.BL(BL31),.BLN(BLN31),.WL(WL55));
sram_cell_6t_5 inst_cell_55_32 (.BL(BL32),.BLN(BLN32),.WL(WL55));
sram_cell_6t_5 inst_cell_55_33 (.BL(BL33),.BLN(BLN33),.WL(WL55));
sram_cell_6t_5 inst_cell_55_34 (.BL(BL34),.BLN(BLN34),.WL(WL55));
sram_cell_6t_5 inst_cell_55_35 (.BL(BL35),.BLN(BLN35),.WL(WL55));
sram_cell_6t_5 inst_cell_55_36 (.BL(BL36),.BLN(BLN36),.WL(WL55));
sram_cell_6t_5 inst_cell_55_37 (.BL(BL37),.BLN(BLN37),.WL(WL55));
sram_cell_6t_5 inst_cell_55_38 (.BL(BL38),.BLN(BLN38),.WL(WL55));
sram_cell_6t_5 inst_cell_55_39 (.BL(BL39),.BLN(BLN39),.WL(WL55));
sram_cell_6t_5 inst_cell_55_40 (.BL(BL40),.BLN(BLN40),.WL(WL55));
sram_cell_6t_5 inst_cell_55_41 (.BL(BL41),.BLN(BLN41),.WL(WL55));
sram_cell_6t_5 inst_cell_55_42 (.BL(BL42),.BLN(BLN42),.WL(WL55));
sram_cell_6t_5 inst_cell_55_43 (.BL(BL43),.BLN(BLN43),.WL(WL55));
sram_cell_6t_5 inst_cell_55_44 (.BL(BL44),.BLN(BLN44),.WL(WL55));
sram_cell_6t_5 inst_cell_55_45 (.BL(BL45),.BLN(BLN45),.WL(WL55));
sram_cell_6t_5 inst_cell_55_46 (.BL(BL46),.BLN(BLN46),.WL(WL55));
sram_cell_6t_5 inst_cell_55_47 (.BL(BL47),.BLN(BLN47),.WL(WL55));
sram_cell_6t_5 inst_cell_55_48 (.BL(BL48),.BLN(BLN48),.WL(WL55));
sram_cell_6t_5 inst_cell_55_49 (.BL(BL49),.BLN(BLN49),.WL(WL55));
sram_cell_6t_5 inst_cell_55_50 (.BL(BL50),.BLN(BLN50),.WL(WL55));
sram_cell_6t_5 inst_cell_55_51 (.BL(BL51),.BLN(BLN51),.WL(WL55));
sram_cell_6t_5 inst_cell_55_52 (.BL(BL52),.BLN(BLN52),.WL(WL55));
sram_cell_6t_5 inst_cell_55_53 (.BL(BL53),.BLN(BLN53),.WL(WL55));
sram_cell_6t_5 inst_cell_55_54 (.BL(BL54),.BLN(BLN54),.WL(WL55));
sram_cell_6t_5 inst_cell_55_55 (.BL(BL55),.BLN(BLN55),.WL(WL55));
sram_cell_6t_5 inst_cell_55_56 (.BL(BL56),.BLN(BLN56),.WL(WL55));
sram_cell_6t_5 inst_cell_55_57 (.BL(BL57),.BLN(BLN57),.WL(WL55));
sram_cell_6t_5 inst_cell_55_58 (.BL(BL58),.BLN(BLN58),.WL(WL55));
sram_cell_6t_5 inst_cell_55_59 (.BL(BL59),.BLN(BLN59),.WL(WL55));
sram_cell_6t_5 inst_cell_55_60 (.BL(BL60),.BLN(BLN60),.WL(WL55));
sram_cell_6t_5 inst_cell_55_61 (.BL(BL61),.BLN(BLN61),.WL(WL55));
sram_cell_6t_5 inst_cell_55_62 (.BL(BL62),.BLN(BLN62),.WL(WL55));
sram_cell_6t_5 inst_cell_55_63 (.BL(BL63),.BLN(BLN63),.WL(WL55));
sram_cell_6t_5 inst_cell_55_64 (.BL(BL64),.BLN(BLN64),.WL(WL55));
sram_cell_6t_5 inst_cell_55_65 (.BL(BL65),.BLN(BLN65),.WL(WL55));
sram_cell_6t_5 inst_cell_55_66 (.BL(BL66),.BLN(BLN66),.WL(WL55));
sram_cell_6t_5 inst_cell_55_67 (.BL(BL67),.BLN(BLN67),.WL(WL55));
sram_cell_6t_5 inst_cell_55_68 (.BL(BL68),.BLN(BLN68),.WL(WL55));
sram_cell_6t_5 inst_cell_55_69 (.BL(BL69),.BLN(BLN69),.WL(WL55));
sram_cell_6t_5 inst_cell_55_70 (.BL(BL70),.BLN(BLN70),.WL(WL55));
sram_cell_6t_5 inst_cell_55_71 (.BL(BL71),.BLN(BLN71),.WL(WL55));
sram_cell_6t_5 inst_cell_55_72 (.BL(BL72),.BLN(BLN72),.WL(WL55));
sram_cell_6t_5 inst_cell_55_73 (.BL(BL73),.BLN(BLN73),.WL(WL55));
sram_cell_6t_5 inst_cell_55_74 (.BL(BL74),.BLN(BLN74),.WL(WL55));
sram_cell_6t_5 inst_cell_55_75 (.BL(BL75),.BLN(BLN75),.WL(WL55));
sram_cell_6t_5 inst_cell_55_76 (.BL(BL76),.BLN(BLN76),.WL(WL55));
sram_cell_6t_5 inst_cell_55_77 (.BL(BL77),.BLN(BLN77),.WL(WL55));
sram_cell_6t_5 inst_cell_55_78 (.BL(BL78),.BLN(BLN78),.WL(WL55));
sram_cell_6t_5 inst_cell_55_79 (.BL(BL79),.BLN(BLN79),.WL(WL55));
sram_cell_6t_5 inst_cell_55_80 (.BL(BL80),.BLN(BLN80),.WL(WL55));
sram_cell_6t_5 inst_cell_55_81 (.BL(BL81),.BLN(BLN81),.WL(WL55));
sram_cell_6t_5 inst_cell_55_82 (.BL(BL82),.BLN(BLN82),.WL(WL55));
sram_cell_6t_5 inst_cell_55_83 (.BL(BL83),.BLN(BLN83),.WL(WL55));
sram_cell_6t_5 inst_cell_55_84 (.BL(BL84),.BLN(BLN84),.WL(WL55));
sram_cell_6t_5 inst_cell_55_85 (.BL(BL85),.BLN(BLN85),.WL(WL55));
sram_cell_6t_5 inst_cell_55_86 (.BL(BL86),.BLN(BLN86),.WL(WL55));
sram_cell_6t_5 inst_cell_55_87 (.BL(BL87),.BLN(BLN87),.WL(WL55));
sram_cell_6t_5 inst_cell_55_88 (.BL(BL88),.BLN(BLN88),.WL(WL55));
sram_cell_6t_5 inst_cell_55_89 (.BL(BL89),.BLN(BLN89),.WL(WL55));
sram_cell_6t_5 inst_cell_55_90 (.BL(BL90),.BLN(BLN90),.WL(WL55));
sram_cell_6t_5 inst_cell_55_91 (.BL(BL91),.BLN(BLN91),.WL(WL55));
sram_cell_6t_5 inst_cell_55_92 (.BL(BL92),.BLN(BLN92),.WL(WL55));
sram_cell_6t_5 inst_cell_55_93 (.BL(BL93),.BLN(BLN93),.WL(WL55));
sram_cell_6t_5 inst_cell_55_94 (.BL(BL94),.BLN(BLN94),.WL(WL55));
sram_cell_6t_5 inst_cell_55_95 (.BL(BL95),.BLN(BLN95),.WL(WL55));
sram_cell_6t_5 inst_cell_55_96 (.BL(BL96),.BLN(BLN96),.WL(WL55));
sram_cell_6t_5 inst_cell_55_97 (.BL(BL97),.BLN(BLN97),.WL(WL55));
sram_cell_6t_5 inst_cell_55_98 (.BL(BL98),.BLN(BLN98),.WL(WL55));
sram_cell_6t_5 inst_cell_55_99 (.BL(BL99),.BLN(BLN99),.WL(WL55));
sram_cell_6t_5 inst_cell_55_100 (.BL(BL100),.BLN(BLN100),.WL(WL55));
sram_cell_6t_5 inst_cell_55_101 (.BL(BL101),.BLN(BLN101),.WL(WL55));
sram_cell_6t_5 inst_cell_55_102 (.BL(BL102),.BLN(BLN102),.WL(WL55));
sram_cell_6t_5 inst_cell_55_103 (.BL(BL103),.BLN(BLN103),.WL(WL55));
sram_cell_6t_5 inst_cell_55_104 (.BL(BL104),.BLN(BLN104),.WL(WL55));
sram_cell_6t_5 inst_cell_55_105 (.BL(BL105),.BLN(BLN105),.WL(WL55));
sram_cell_6t_5 inst_cell_55_106 (.BL(BL106),.BLN(BLN106),.WL(WL55));
sram_cell_6t_5 inst_cell_55_107 (.BL(BL107),.BLN(BLN107),.WL(WL55));
sram_cell_6t_5 inst_cell_55_108 (.BL(BL108),.BLN(BLN108),.WL(WL55));
sram_cell_6t_5 inst_cell_55_109 (.BL(BL109),.BLN(BLN109),.WL(WL55));
sram_cell_6t_5 inst_cell_55_110 (.BL(BL110),.BLN(BLN110),.WL(WL55));
sram_cell_6t_5 inst_cell_55_111 (.BL(BL111),.BLN(BLN111),.WL(WL55));
sram_cell_6t_5 inst_cell_55_112 (.BL(BL112),.BLN(BLN112),.WL(WL55));
sram_cell_6t_5 inst_cell_55_113 (.BL(BL113),.BLN(BLN113),.WL(WL55));
sram_cell_6t_5 inst_cell_55_114 (.BL(BL114),.BLN(BLN114),.WL(WL55));
sram_cell_6t_5 inst_cell_55_115 (.BL(BL115),.BLN(BLN115),.WL(WL55));
sram_cell_6t_5 inst_cell_55_116 (.BL(BL116),.BLN(BLN116),.WL(WL55));
sram_cell_6t_5 inst_cell_55_117 (.BL(BL117),.BLN(BLN117),.WL(WL55));
sram_cell_6t_5 inst_cell_55_118 (.BL(BL118),.BLN(BLN118),.WL(WL55));
sram_cell_6t_5 inst_cell_55_119 (.BL(BL119),.BLN(BLN119),.WL(WL55));
sram_cell_6t_5 inst_cell_55_120 (.BL(BL120),.BLN(BLN120),.WL(WL55));
sram_cell_6t_5 inst_cell_55_121 (.BL(BL121),.BLN(BLN121),.WL(WL55));
sram_cell_6t_5 inst_cell_55_122 (.BL(BL122),.BLN(BLN122),.WL(WL55));
sram_cell_6t_5 inst_cell_55_123 (.BL(BL123),.BLN(BLN123),.WL(WL55));
sram_cell_6t_5 inst_cell_55_124 (.BL(BL124),.BLN(BLN124),.WL(WL55));
sram_cell_6t_5 inst_cell_55_125 (.BL(BL125),.BLN(BLN125),.WL(WL55));
sram_cell_6t_5 inst_cell_55_126 (.BL(BL126),.BLN(BLN126),.WL(WL55));
sram_cell_6t_5 inst_cell_55_127 (.BL(BL127),.BLN(BLN127),.WL(WL55));
sram_cell_6t_5 inst_cell_56_0 (.BL(BL0),.BLN(BLN0),.WL(WL56));
sram_cell_6t_5 inst_cell_56_1 (.BL(BL1),.BLN(BLN1),.WL(WL56));
sram_cell_6t_5 inst_cell_56_2 (.BL(BL2),.BLN(BLN2),.WL(WL56));
sram_cell_6t_5 inst_cell_56_3 (.BL(BL3),.BLN(BLN3),.WL(WL56));
sram_cell_6t_5 inst_cell_56_4 (.BL(BL4),.BLN(BLN4),.WL(WL56));
sram_cell_6t_5 inst_cell_56_5 (.BL(BL5),.BLN(BLN5),.WL(WL56));
sram_cell_6t_5 inst_cell_56_6 (.BL(BL6),.BLN(BLN6),.WL(WL56));
sram_cell_6t_5 inst_cell_56_7 (.BL(BL7),.BLN(BLN7),.WL(WL56));
sram_cell_6t_5 inst_cell_56_8 (.BL(BL8),.BLN(BLN8),.WL(WL56));
sram_cell_6t_5 inst_cell_56_9 (.BL(BL9),.BLN(BLN9),.WL(WL56));
sram_cell_6t_5 inst_cell_56_10 (.BL(BL10),.BLN(BLN10),.WL(WL56));
sram_cell_6t_5 inst_cell_56_11 (.BL(BL11),.BLN(BLN11),.WL(WL56));
sram_cell_6t_5 inst_cell_56_12 (.BL(BL12),.BLN(BLN12),.WL(WL56));
sram_cell_6t_5 inst_cell_56_13 (.BL(BL13),.BLN(BLN13),.WL(WL56));
sram_cell_6t_5 inst_cell_56_14 (.BL(BL14),.BLN(BLN14),.WL(WL56));
sram_cell_6t_5 inst_cell_56_15 (.BL(BL15),.BLN(BLN15),.WL(WL56));
sram_cell_6t_5 inst_cell_56_16 (.BL(BL16),.BLN(BLN16),.WL(WL56));
sram_cell_6t_5 inst_cell_56_17 (.BL(BL17),.BLN(BLN17),.WL(WL56));
sram_cell_6t_5 inst_cell_56_18 (.BL(BL18),.BLN(BLN18),.WL(WL56));
sram_cell_6t_5 inst_cell_56_19 (.BL(BL19),.BLN(BLN19),.WL(WL56));
sram_cell_6t_5 inst_cell_56_20 (.BL(BL20),.BLN(BLN20),.WL(WL56));
sram_cell_6t_5 inst_cell_56_21 (.BL(BL21),.BLN(BLN21),.WL(WL56));
sram_cell_6t_5 inst_cell_56_22 (.BL(BL22),.BLN(BLN22),.WL(WL56));
sram_cell_6t_5 inst_cell_56_23 (.BL(BL23),.BLN(BLN23),.WL(WL56));
sram_cell_6t_5 inst_cell_56_24 (.BL(BL24),.BLN(BLN24),.WL(WL56));
sram_cell_6t_5 inst_cell_56_25 (.BL(BL25),.BLN(BLN25),.WL(WL56));
sram_cell_6t_5 inst_cell_56_26 (.BL(BL26),.BLN(BLN26),.WL(WL56));
sram_cell_6t_5 inst_cell_56_27 (.BL(BL27),.BLN(BLN27),.WL(WL56));
sram_cell_6t_5 inst_cell_56_28 (.BL(BL28),.BLN(BLN28),.WL(WL56));
sram_cell_6t_5 inst_cell_56_29 (.BL(BL29),.BLN(BLN29),.WL(WL56));
sram_cell_6t_5 inst_cell_56_30 (.BL(BL30),.BLN(BLN30),.WL(WL56));
sram_cell_6t_5 inst_cell_56_31 (.BL(BL31),.BLN(BLN31),.WL(WL56));
sram_cell_6t_5 inst_cell_56_32 (.BL(BL32),.BLN(BLN32),.WL(WL56));
sram_cell_6t_5 inst_cell_56_33 (.BL(BL33),.BLN(BLN33),.WL(WL56));
sram_cell_6t_5 inst_cell_56_34 (.BL(BL34),.BLN(BLN34),.WL(WL56));
sram_cell_6t_5 inst_cell_56_35 (.BL(BL35),.BLN(BLN35),.WL(WL56));
sram_cell_6t_5 inst_cell_56_36 (.BL(BL36),.BLN(BLN36),.WL(WL56));
sram_cell_6t_5 inst_cell_56_37 (.BL(BL37),.BLN(BLN37),.WL(WL56));
sram_cell_6t_5 inst_cell_56_38 (.BL(BL38),.BLN(BLN38),.WL(WL56));
sram_cell_6t_5 inst_cell_56_39 (.BL(BL39),.BLN(BLN39),.WL(WL56));
sram_cell_6t_5 inst_cell_56_40 (.BL(BL40),.BLN(BLN40),.WL(WL56));
sram_cell_6t_5 inst_cell_56_41 (.BL(BL41),.BLN(BLN41),.WL(WL56));
sram_cell_6t_5 inst_cell_56_42 (.BL(BL42),.BLN(BLN42),.WL(WL56));
sram_cell_6t_5 inst_cell_56_43 (.BL(BL43),.BLN(BLN43),.WL(WL56));
sram_cell_6t_5 inst_cell_56_44 (.BL(BL44),.BLN(BLN44),.WL(WL56));
sram_cell_6t_5 inst_cell_56_45 (.BL(BL45),.BLN(BLN45),.WL(WL56));
sram_cell_6t_5 inst_cell_56_46 (.BL(BL46),.BLN(BLN46),.WL(WL56));
sram_cell_6t_5 inst_cell_56_47 (.BL(BL47),.BLN(BLN47),.WL(WL56));
sram_cell_6t_5 inst_cell_56_48 (.BL(BL48),.BLN(BLN48),.WL(WL56));
sram_cell_6t_5 inst_cell_56_49 (.BL(BL49),.BLN(BLN49),.WL(WL56));
sram_cell_6t_5 inst_cell_56_50 (.BL(BL50),.BLN(BLN50),.WL(WL56));
sram_cell_6t_5 inst_cell_56_51 (.BL(BL51),.BLN(BLN51),.WL(WL56));
sram_cell_6t_5 inst_cell_56_52 (.BL(BL52),.BLN(BLN52),.WL(WL56));
sram_cell_6t_5 inst_cell_56_53 (.BL(BL53),.BLN(BLN53),.WL(WL56));
sram_cell_6t_5 inst_cell_56_54 (.BL(BL54),.BLN(BLN54),.WL(WL56));
sram_cell_6t_5 inst_cell_56_55 (.BL(BL55),.BLN(BLN55),.WL(WL56));
sram_cell_6t_5 inst_cell_56_56 (.BL(BL56),.BLN(BLN56),.WL(WL56));
sram_cell_6t_5 inst_cell_56_57 (.BL(BL57),.BLN(BLN57),.WL(WL56));
sram_cell_6t_5 inst_cell_56_58 (.BL(BL58),.BLN(BLN58),.WL(WL56));
sram_cell_6t_5 inst_cell_56_59 (.BL(BL59),.BLN(BLN59),.WL(WL56));
sram_cell_6t_5 inst_cell_56_60 (.BL(BL60),.BLN(BLN60),.WL(WL56));
sram_cell_6t_5 inst_cell_56_61 (.BL(BL61),.BLN(BLN61),.WL(WL56));
sram_cell_6t_5 inst_cell_56_62 (.BL(BL62),.BLN(BLN62),.WL(WL56));
sram_cell_6t_5 inst_cell_56_63 (.BL(BL63),.BLN(BLN63),.WL(WL56));
sram_cell_6t_5 inst_cell_56_64 (.BL(BL64),.BLN(BLN64),.WL(WL56));
sram_cell_6t_5 inst_cell_56_65 (.BL(BL65),.BLN(BLN65),.WL(WL56));
sram_cell_6t_5 inst_cell_56_66 (.BL(BL66),.BLN(BLN66),.WL(WL56));
sram_cell_6t_5 inst_cell_56_67 (.BL(BL67),.BLN(BLN67),.WL(WL56));
sram_cell_6t_5 inst_cell_56_68 (.BL(BL68),.BLN(BLN68),.WL(WL56));
sram_cell_6t_5 inst_cell_56_69 (.BL(BL69),.BLN(BLN69),.WL(WL56));
sram_cell_6t_5 inst_cell_56_70 (.BL(BL70),.BLN(BLN70),.WL(WL56));
sram_cell_6t_5 inst_cell_56_71 (.BL(BL71),.BLN(BLN71),.WL(WL56));
sram_cell_6t_5 inst_cell_56_72 (.BL(BL72),.BLN(BLN72),.WL(WL56));
sram_cell_6t_5 inst_cell_56_73 (.BL(BL73),.BLN(BLN73),.WL(WL56));
sram_cell_6t_5 inst_cell_56_74 (.BL(BL74),.BLN(BLN74),.WL(WL56));
sram_cell_6t_5 inst_cell_56_75 (.BL(BL75),.BLN(BLN75),.WL(WL56));
sram_cell_6t_5 inst_cell_56_76 (.BL(BL76),.BLN(BLN76),.WL(WL56));
sram_cell_6t_5 inst_cell_56_77 (.BL(BL77),.BLN(BLN77),.WL(WL56));
sram_cell_6t_5 inst_cell_56_78 (.BL(BL78),.BLN(BLN78),.WL(WL56));
sram_cell_6t_5 inst_cell_56_79 (.BL(BL79),.BLN(BLN79),.WL(WL56));
sram_cell_6t_5 inst_cell_56_80 (.BL(BL80),.BLN(BLN80),.WL(WL56));
sram_cell_6t_5 inst_cell_56_81 (.BL(BL81),.BLN(BLN81),.WL(WL56));
sram_cell_6t_5 inst_cell_56_82 (.BL(BL82),.BLN(BLN82),.WL(WL56));
sram_cell_6t_5 inst_cell_56_83 (.BL(BL83),.BLN(BLN83),.WL(WL56));
sram_cell_6t_5 inst_cell_56_84 (.BL(BL84),.BLN(BLN84),.WL(WL56));
sram_cell_6t_5 inst_cell_56_85 (.BL(BL85),.BLN(BLN85),.WL(WL56));
sram_cell_6t_5 inst_cell_56_86 (.BL(BL86),.BLN(BLN86),.WL(WL56));
sram_cell_6t_5 inst_cell_56_87 (.BL(BL87),.BLN(BLN87),.WL(WL56));
sram_cell_6t_5 inst_cell_56_88 (.BL(BL88),.BLN(BLN88),.WL(WL56));
sram_cell_6t_5 inst_cell_56_89 (.BL(BL89),.BLN(BLN89),.WL(WL56));
sram_cell_6t_5 inst_cell_56_90 (.BL(BL90),.BLN(BLN90),.WL(WL56));
sram_cell_6t_5 inst_cell_56_91 (.BL(BL91),.BLN(BLN91),.WL(WL56));
sram_cell_6t_5 inst_cell_56_92 (.BL(BL92),.BLN(BLN92),.WL(WL56));
sram_cell_6t_5 inst_cell_56_93 (.BL(BL93),.BLN(BLN93),.WL(WL56));
sram_cell_6t_5 inst_cell_56_94 (.BL(BL94),.BLN(BLN94),.WL(WL56));
sram_cell_6t_5 inst_cell_56_95 (.BL(BL95),.BLN(BLN95),.WL(WL56));
sram_cell_6t_5 inst_cell_56_96 (.BL(BL96),.BLN(BLN96),.WL(WL56));
sram_cell_6t_5 inst_cell_56_97 (.BL(BL97),.BLN(BLN97),.WL(WL56));
sram_cell_6t_5 inst_cell_56_98 (.BL(BL98),.BLN(BLN98),.WL(WL56));
sram_cell_6t_5 inst_cell_56_99 (.BL(BL99),.BLN(BLN99),.WL(WL56));
sram_cell_6t_5 inst_cell_56_100 (.BL(BL100),.BLN(BLN100),.WL(WL56));
sram_cell_6t_5 inst_cell_56_101 (.BL(BL101),.BLN(BLN101),.WL(WL56));
sram_cell_6t_5 inst_cell_56_102 (.BL(BL102),.BLN(BLN102),.WL(WL56));
sram_cell_6t_5 inst_cell_56_103 (.BL(BL103),.BLN(BLN103),.WL(WL56));
sram_cell_6t_5 inst_cell_56_104 (.BL(BL104),.BLN(BLN104),.WL(WL56));
sram_cell_6t_5 inst_cell_56_105 (.BL(BL105),.BLN(BLN105),.WL(WL56));
sram_cell_6t_5 inst_cell_56_106 (.BL(BL106),.BLN(BLN106),.WL(WL56));
sram_cell_6t_5 inst_cell_56_107 (.BL(BL107),.BLN(BLN107),.WL(WL56));
sram_cell_6t_5 inst_cell_56_108 (.BL(BL108),.BLN(BLN108),.WL(WL56));
sram_cell_6t_5 inst_cell_56_109 (.BL(BL109),.BLN(BLN109),.WL(WL56));
sram_cell_6t_5 inst_cell_56_110 (.BL(BL110),.BLN(BLN110),.WL(WL56));
sram_cell_6t_5 inst_cell_56_111 (.BL(BL111),.BLN(BLN111),.WL(WL56));
sram_cell_6t_5 inst_cell_56_112 (.BL(BL112),.BLN(BLN112),.WL(WL56));
sram_cell_6t_5 inst_cell_56_113 (.BL(BL113),.BLN(BLN113),.WL(WL56));
sram_cell_6t_5 inst_cell_56_114 (.BL(BL114),.BLN(BLN114),.WL(WL56));
sram_cell_6t_5 inst_cell_56_115 (.BL(BL115),.BLN(BLN115),.WL(WL56));
sram_cell_6t_5 inst_cell_56_116 (.BL(BL116),.BLN(BLN116),.WL(WL56));
sram_cell_6t_5 inst_cell_56_117 (.BL(BL117),.BLN(BLN117),.WL(WL56));
sram_cell_6t_5 inst_cell_56_118 (.BL(BL118),.BLN(BLN118),.WL(WL56));
sram_cell_6t_5 inst_cell_56_119 (.BL(BL119),.BLN(BLN119),.WL(WL56));
sram_cell_6t_5 inst_cell_56_120 (.BL(BL120),.BLN(BLN120),.WL(WL56));
sram_cell_6t_5 inst_cell_56_121 (.BL(BL121),.BLN(BLN121),.WL(WL56));
sram_cell_6t_5 inst_cell_56_122 (.BL(BL122),.BLN(BLN122),.WL(WL56));
sram_cell_6t_5 inst_cell_56_123 (.BL(BL123),.BLN(BLN123),.WL(WL56));
sram_cell_6t_5 inst_cell_56_124 (.BL(BL124),.BLN(BLN124),.WL(WL56));
sram_cell_6t_5 inst_cell_56_125 (.BL(BL125),.BLN(BLN125),.WL(WL56));
sram_cell_6t_5 inst_cell_56_126 (.BL(BL126),.BLN(BLN126),.WL(WL56));
sram_cell_6t_5 inst_cell_56_127 (.BL(BL127),.BLN(BLN127),.WL(WL56));
sram_cell_6t_5 inst_cell_57_0 (.BL(BL0),.BLN(BLN0),.WL(WL57));
sram_cell_6t_5 inst_cell_57_1 (.BL(BL1),.BLN(BLN1),.WL(WL57));
sram_cell_6t_5 inst_cell_57_2 (.BL(BL2),.BLN(BLN2),.WL(WL57));
sram_cell_6t_5 inst_cell_57_3 (.BL(BL3),.BLN(BLN3),.WL(WL57));
sram_cell_6t_5 inst_cell_57_4 (.BL(BL4),.BLN(BLN4),.WL(WL57));
sram_cell_6t_5 inst_cell_57_5 (.BL(BL5),.BLN(BLN5),.WL(WL57));
sram_cell_6t_5 inst_cell_57_6 (.BL(BL6),.BLN(BLN6),.WL(WL57));
sram_cell_6t_5 inst_cell_57_7 (.BL(BL7),.BLN(BLN7),.WL(WL57));
sram_cell_6t_5 inst_cell_57_8 (.BL(BL8),.BLN(BLN8),.WL(WL57));
sram_cell_6t_5 inst_cell_57_9 (.BL(BL9),.BLN(BLN9),.WL(WL57));
sram_cell_6t_5 inst_cell_57_10 (.BL(BL10),.BLN(BLN10),.WL(WL57));
sram_cell_6t_5 inst_cell_57_11 (.BL(BL11),.BLN(BLN11),.WL(WL57));
sram_cell_6t_5 inst_cell_57_12 (.BL(BL12),.BLN(BLN12),.WL(WL57));
sram_cell_6t_5 inst_cell_57_13 (.BL(BL13),.BLN(BLN13),.WL(WL57));
sram_cell_6t_5 inst_cell_57_14 (.BL(BL14),.BLN(BLN14),.WL(WL57));
sram_cell_6t_5 inst_cell_57_15 (.BL(BL15),.BLN(BLN15),.WL(WL57));
sram_cell_6t_5 inst_cell_57_16 (.BL(BL16),.BLN(BLN16),.WL(WL57));
sram_cell_6t_5 inst_cell_57_17 (.BL(BL17),.BLN(BLN17),.WL(WL57));
sram_cell_6t_5 inst_cell_57_18 (.BL(BL18),.BLN(BLN18),.WL(WL57));
sram_cell_6t_5 inst_cell_57_19 (.BL(BL19),.BLN(BLN19),.WL(WL57));
sram_cell_6t_5 inst_cell_57_20 (.BL(BL20),.BLN(BLN20),.WL(WL57));
sram_cell_6t_5 inst_cell_57_21 (.BL(BL21),.BLN(BLN21),.WL(WL57));
sram_cell_6t_5 inst_cell_57_22 (.BL(BL22),.BLN(BLN22),.WL(WL57));
sram_cell_6t_5 inst_cell_57_23 (.BL(BL23),.BLN(BLN23),.WL(WL57));
sram_cell_6t_5 inst_cell_57_24 (.BL(BL24),.BLN(BLN24),.WL(WL57));
sram_cell_6t_5 inst_cell_57_25 (.BL(BL25),.BLN(BLN25),.WL(WL57));
sram_cell_6t_5 inst_cell_57_26 (.BL(BL26),.BLN(BLN26),.WL(WL57));
sram_cell_6t_5 inst_cell_57_27 (.BL(BL27),.BLN(BLN27),.WL(WL57));
sram_cell_6t_5 inst_cell_57_28 (.BL(BL28),.BLN(BLN28),.WL(WL57));
sram_cell_6t_5 inst_cell_57_29 (.BL(BL29),.BLN(BLN29),.WL(WL57));
sram_cell_6t_5 inst_cell_57_30 (.BL(BL30),.BLN(BLN30),.WL(WL57));
sram_cell_6t_5 inst_cell_57_31 (.BL(BL31),.BLN(BLN31),.WL(WL57));
sram_cell_6t_5 inst_cell_57_32 (.BL(BL32),.BLN(BLN32),.WL(WL57));
sram_cell_6t_5 inst_cell_57_33 (.BL(BL33),.BLN(BLN33),.WL(WL57));
sram_cell_6t_5 inst_cell_57_34 (.BL(BL34),.BLN(BLN34),.WL(WL57));
sram_cell_6t_5 inst_cell_57_35 (.BL(BL35),.BLN(BLN35),.WL(WL57));
sram_cell_6t_5 inst_cell_57_36 (.BL(BL36),.BLN(BLN36),.WL(WL57));
sram_cell_6t_5 inst_cell_57_37 (.BL(BL37),.BLN(BLN37),.WL(WL57));
sram_cell_6t_5 inst_cell_57_38 (.BL(BL38),.BLN(BLN38),.WL(WL57));
sram_cell_6t_5 inst_cell_57_39 (.BL(BL39),.BLN(BLN39),.WL(WL57));
sram_cell_6t_5 inst_cell_57_40 (.BL(BL40),.BLN(BLN40),.WL(WL57));
sram_cell_6t_5 inst_cell_57_41 (.BL(BL41),.BLN(BLN41),.WL(WL57));
sram_cell_6t_5 inst_cell_57_42 (.BL(BL42),.BLN(BLN42),.WL(WL57));
sram_cell_6t_5 inst_cell_57_43 (.BL(BL43),.BLN(BLN43),.WL(WL57));
sram_cell_6t_5 inst_cell_57_44 (.BL(BL44),.BLN(BLN44),.WL(WL57));
sram_cell_6t_5 inst_cell_57_45 (.BL(BL45),.BLN(BLN45),.WL(WL57));
sram_cell_6t_5 inst_cell_57_46 (.BL(BL46),.BLN(BLN46),.WL(WL57));
sram_cell_6t_5 inst_cell_57_47 (.BL(BL47),.BLN(BLN47),.WL(WL57));
sram_cell_6t_5 inst_cell_57_48 (.BL(BL48),.BLN(BLN48),.WL(WL57));
sram_cell_6t_5 inst_cell_57_49 (.BL(BL49),.BLN(BLN49),.WL(WL57));
sram_cell_6t_5 inst_cell_57_50 (.BL(BL50),.BLN(BLN50),.WL(WL57));
sram_cell_6t_5 inst_cell_57_51 (.BL(BL51),.BLN(BLN51),.WL(WL57));
sram_cell_6t_5 inst_cell_57_52 (.BL(BL52),.BLN(BLN52),.WL(WL57));
sram_cell_6t_5 inst_cell_57_53 (.BL(BL53),.BLN(BLN53),.WL(WL57));
sram_cell_6t_5 inst_cell_57_54 (.BL(BL54),.BLN(BLN54),.WL(WL57));
sram_cell_6t_5 inst_cell_57_55 (.BL(BL55),.BLN(BLN55),.WL(WL57));
sram_cell_6t_5 inst_cell_57_56 (.BL(BL56),.BLN(BLN56),.WL(WL57));
sram_cell_6t_5 inst_cell_57_57 (.BL(BL57),.BLN(BLN57),.WL(WL57));
sram_cell_6t_5 inst_cell_57_58 (.BL(BL58),.BLN(BLN58),.WL(WL57));
sram_cell_6t_5 inst_cell_57_59 (.BL(BL59),.BLN(BLN59),.WL(WL57));
sram_cell_6t_5 inst_cell_57_60 (.BL(BL60),.BLN(BLN60),.WL(WL57));
sram_cell_6t_5 inst_cell_57_61 (.BL(BL61),.BLN(BLN61),.WL(WL57));
sram_cell_6t_5 inst_cell_57_62 (.BL(BL62),.BLN(BLN62),.WL(WL57));
sram_cell_6t_5 inst_cell_57_63 (.BL(BL63),.BLN(BLN63),.WL(WL57));
sram_cell_6t_5 inst_cell_57_64 (.BL(BL64),.BLN(BLN64),.WL(WL57));
sram_cell_6t_5 inst_cell_57_65 (.BL(BL65),.BLN(BLN65),.WL(WL57));
sram_cell_6t_5 inst_cell_57_66 (.BL(BL66),.BLN(BLN66),.WL(WL57));
sram_cell_6t_5 inst_cell_57_67 (.BL(BL67),.BLN(BLN67),.WL(WL57));
sram_cell_6t_5 inst_cell_57_68 (.BL(BL68),.BLN(BLN68),.WL(WL57));
sram_cell_6t_5 inst_cell_57_69 (.BL(BL69),.BLN(BLN69),.WL(WL57));
sram_cell_6t_5 inst_cell_57_70 (.BL(BL70),.BLN(BLN70),.WL(WL57));
sram_cell_6t_5 inst_cell_57_71 (.BL(BL71),.BLN(BLN71),.WL(WL57));
sram_cell_6t_5 inst_cell_57_72 (.BL(BL72),.BLN(BLN72),.WL(WL57));
sram_cell_6t_5 inst_cell_57_73 (.BL(BL73),.BLN(BLN73),.WL(WL57));
sram_cell_6t_5 inst_cell_57_74 (.BL(BL74),.BLN(BLN74),.WL(WL57));
sram_cell_6t_5 inst_cell_57_75 (.BL(BL75),.BLN(BLN75),.WL(WL57));
sram_cell_6t_5 inst_cell_57_76 (.BL(BL76),.BLN(BLN76),.WL(WL57));
sram_cell_6t_5 inst_cell_57_77 (.BL(BL77),.BLN(BLN77),.WL(WL57));
sram_cell_6t_5 inst_cell_57_78 (.BL(BL78),.BLN(BLN78),.WL(WL57));
sram_cell_6t_5 inst_cell_57_79 (.BL(BL79),.BLN(BLN79),.WL(WL57));
sram_cell_6t_5 inst_cell_57_80 (.BL(BL80),.BLN(BLN80),.WL(WL57));
sram_cell_6t_5 inst_cell_57_81 (.BL(BL81),.BLN(BLN81),.WL(WL57));
sram_cell_6t_5 inst_cell_57_82 (.BL(BL82),.BLN(BLN82),.WL(WL57));
sram_cell_6t_5 inst_cell_57_83 (.BL(BL83),.BLN(BLN83),.WL(WL57));
sram_cell_6t_5 inst_cell_57_84 (.BL(BL84),.BLN(BLN84),.WL(WL57));
sram_cell_6t_5 inst_cell_57_85 (.BL(BL85),.BLN(BLN85),.WL(WL57));
sram_cell_6t_5 inst_cell_57_86 (.BL(BL86),.BLN(BLN86),.WL(WL57));
sram_cell_6t_5 inst_cell_57_87 (.BL(BL87),.BLN(BLN87),.WL(WL57));
sram_cell_6t_5 inst_cell_57_88 (.BL(BL88),.BLN(BLN88),.WL(WL57));
sram_cell_6t_5 inst_cell_57_89 (.BL(BL89),.BLN(BLN89),.WL(WL57));
sram_cell_6t_5 inst_cell_57_90 (.BL(BL90),.BLN(BLN90),.WL(WL57));
sram_cell_6t_5 inst_cell_57_91 (.BL(BL91),.BLN(BLN91),.WL(WL57));
sram_cell_6t_5 inst_cell_57_92 (.BL(BL92),.BLN(BLN92),.WL(WL57));
sram_cell_6t_5 inst_cell_57_93 (.BL(BL93),.BLN(BLN93),.WL(WL57));
sram_cell_6t_5 inst_cell_57_94 (.BL(BL94),.BLN(BLN94),.WL(WL57));
sram_cell_6t_5 inst_cell_57_95 (.BL(BL95),.BLN(BLN95),.WL(WL57));
sram_cell_6t_5 inst_cell_57_96 (.BL(BL96),.BLN(BLN96),.WL(WL57));
sram_cell_6t_5 inst_cell_57_97 (.BL(BL97),.BLN(BLN97),.WL(WL57));
sram_cell_6t_5 inst_cell_57_98 (.BL(BL98),.BLN(BLN98),.WL(WL57));
sram_cell_6t_5 inst_cell_57_99 (.BL(BL99),.BLN(BLN99),.WL(WL57));
sram_cell_6t_5 inst_cell_57_100 (.BL(BL100),.BLN(BLN100),.WL(WL57));
sram_cell_6t_5 inst_cell_57_101 (.BL(BL101),.BLN(BLN101),.WL(WL57));
sram_cell_6t_5 inst_cell_57_102 (.BL(BL102),.BLN(BLN102),.WL(WL57));
sram_cell_6t_5 inst_cell_57_103 (.BL(BL103),.BLN(BLN103),.WL(WL57));
sram_cell_6t_5 inst_cell_57_104 (.BL(BL104),.BLN(BLN104),.WL(WL57));
sram_cell_6t_5 inst_cell_57_105 (.BL(BL105),.BLN(BLN105),.WL(WL57));
sram_cell_6t_5 inst_cell_57_106 (.BL(BL106),.BLN(BLN106),.WL(WL57));
sram_cell_6t_5 inst_cell_57_107 (.BL(BL107),.BLN(BLN107),.WL(WL57));
sram_cell_6t_5 inst_cell_57_108 (.BL(BL108),.BLN(BLN108),.WL(WL57));
sram_cell_6t_5 inst_cell_57_109 (.BL(BL109),.BLN(BLN109),.WL(WL57));
sram_cell_6t_5 inst_cell_57_110 (.BL(BL110),.BLN(BLN110),.WL(WL57));
sram_cell_6t_5 inst_cell_57_111 (.BL(BL111),.BLN(BLN111),.WL(WL57));
sram_cell_6t_5 inst_cell_57_112 (.BL(BL112),.BLN(BLN112),.WL(WL57));
sram_cell_6t_5 inst_cell_57_113 (.BL(BL113),.BLN(BLN113),.WL(WL57));
sram_cell_6t_5 inst_cell_57_114 (.BL(BL114),.BLN(BLN114),.WL(WL57));
sram_cell_6t_5 inst_cell_57_115 (.BL(BL115),.BLN(BLN115),.WL(WL57));
sram_cell_6t_5 inst_cell_57_116 (.BL(BL116),.BLN(BLN116),.WL(WL57));
sram_cell_6t_5 inst_cell_57_117 (.BL(BL117),.BLN(BLN117),.WL(WL57));
sram_cell_6t_5 inst_cell_57_118 (.BL(BL118),.BLN(BLN118),.WL(WL57));
sram_cell_6t_5 inst_cell_57_119 (.BL(BL119),.BLN(BLN119),.WL(WL57));
sram_cell_6t_5 inst_cell_57_120 (.BL(BL120),.BLN(BLN120),.WL(WL57));
sram_cell_6t_5 inst_cell_57_121 (.BL(BL121),.BLN(BLN121),.WL(WL57));
sram_cell_6t_5 inst_cell_57_122 (.BL(BL122),.BLN(BLN122),.WL(WL57));
sram_cell_6t_5 inst_cell_57_123 (.BL(BL123),.BLN(BLN123),.WL(WL57));
sram_cell_6t_5 inst_cell_57_124 (.BL(BL124),.BLN(BLN124),.WL(WL57));
sram_cell_6t_5 inst_cell_57_125 (.BL(BL125),.BLN(BLN125),.WL(WL57));
sram_cell_6t_5 inst_cell_57_126 (.BL(BL126),.BLN(BLN126),.WL(WL57));
sram_cell_6t_5 inst_cell_57_127 (.BL(BL127),.BLN(BLN127),.WL(WL57));
sram_cell_6t_5 inst_cell_58_0 (.BL(BL0),.BLN(BLN0),.WL(WL58));
sram_cell_6t_5 inst_cell_58_1 (.BL(BL1),.BLN(BLN1),.WL(WL58));
sram_cell_6t_5 inst_cell_58_2 (.BL(BL2),.BLN(BLN2),.WL(WL58));
sram_cell_6t_5 inst_cell_58_3 (.BL(BL3),.BLN(BLN3),.WL(WL58));
sram_cell_6t_5 inst_cell_58_4 (.BL(BL4),.BLN(BLN4),.WL(WL58));
sram_cell_6t_5 inst_cell_58_5 (.BL(BL5),.BLN(BLN5),.WL(WL58));
sram_cell_6t_5 inst_cell_58_6 (.BL(BL6),.BLN(BLN6),.WL(WL58));
sram_cell_6t_5 inst_cell_58_7 (.BL(BL7),.BLN(BLN7),.WL(WL58));
sram_cell_6t_5 inst_cell_58_8 (.BL(BL8),.BLN(BLN8),.WL(WL58));
sram_cell_6t_5 inst_cell_58_9 (.BL(BL9),.BLN(BLN9),.WL(WL58));
sram_cell_6t_5 inst_cell_58_10 (.BL(BL10),.BLN(BLN10),.WL(WL58));
sram_cell_6t_5 inst_cell_58_11 (.BL(BL11),.BLN(BLN11),.WL(WL58));
sram_cell_6t_5 inst_cell_58_12 (.BL(BL12),.BLN(BLN12),.WL(WL58));
sram_cell_6t_5 inst_cell_58_13 (.BL(BL13),.BLN(BLN13),.WL(WL58));
sram_cell_6t_5 inst_cell_58_14 (.BL(BL14),.BLN(BLN14),.WL(WL58));
sram_cell_6t_5 inst_cell_58_15 (.BL(BL15),.BLN(BLN15),.WL(WL58));
sram_cell_6t_5 inst_cell_58_16 (.BL(BL16),.BLN(BLN16),.WL(WL58));
sram_cell_6t_5 inst_cell_58_17 (.BL(BL17),.BLN(BLN17),.WL(WL58));
sram_cell_6t_5 inst_cell_58_18 (.BL(BL18),.BLN(BLN18),.WL(WL58));
sram_cell_6t_5 inst_cell_58_19 (.BL(BL19),.BLN(BLN19),.WL(WL58));
sram_cell_6t_5 inst_cell_58_20 (.BL(BL20),.BLN(BLN20),.WL(WL58));
sram_cell_6t_5 inst_cell_58_21 (.BL(BL21),.BLN(BLN21),.WL(WL58));
sram_cell_6t_5 inst_cell_58_22 (.BL(BL22),.BLN(BLN22),.WL(WL58));
sram_cell_6t_5 inst_cell_58_23 (.BL(BL23),.BLN(BLN23),.WL(WL58));
sram_cell_6t_5 inst_cell_58_24 (.BL(BL24),.BLN(BLN24),.WL(WL58));
sram_cell_6t_5 inst_cell_58_25 (.BL(BL25),.BLN(BLN25),.WL(WL58));
sram_cell_6t_5 inst_cell_58_26 (.BL(BL26),.BLN(BLN26),.WL(WL58));
sram_cell_6t_5 inst_cell_58_27 (.BL(BL27),.BLN(BLN27),.WL(WL58));
sram_cell_6t_5 inst_cell_58_28 (.BL(BL28),.BLN(BLN28),.WL(WL58));
sram_cell_6t_5 inst_cell_58_29 (.BL(BL29),.BLN(BLN29),.WL(WL58));
sram_cell_6t_5 inst_cell_58_30 (.BL(BL30),.BLN(BLN30),.WL(WL58));
sram_cell_6t_5 inst_cell_58_31 (.BL(BL31),.BLN(BLN31),.WL(WL58));
sram_cell_6t_5 inst_cell_58_32 (.BL(BL32),.BLN(BLN32),.WL(WL58));
sram_cell_6t_5 inst_cell_58_33 (.BL(BL33),.BLN(BLN33),.WL(WL58));
sram_cell_6t_5 inst_cell_58_34 (.BL(BL34),.BLN(BLN34),.WL(WL58));
sram_cell_6t_5 inst_cell_58_35 (.BL(BL35),.BLN(BLN35),.WL(WL58));
sram_cell_6t_5 inst_cell_58_36 (.BL(BL36),.BLN(BLN36),.WL(WL58));
sram_cell_6t_5 inst_cell_58_37 (.BL(BL37),.BLN(BLN37),.WL(WL58));
sram_cell_6t_5 inst_cell_58_38 (.BL(BL38),.BLN(BLN38),.WL(WL58));
sram_cell_6t_5 inst_cell_58_39 (.BL(BL39),.BLN(BLN39),.WL(WL58));
sram_cell_6t_5 inst_cell_58_40 (.BL(BL40),.BLN(BLN40),.WL(WL58));
sram_cell_6t_5 inst_cell_58_41 (.BL(BL41),.BLN(BLN41),.WL(WL58));
sram_cell_6t_5 inst_cell_58_42 (.BL(BL42),.BLN(BLN42),.WL(WL58));
sram_cell_6t_5 inst_cell_58_43 (.BL(BL43),.BLN(BLN43),.WL(WL58));
sram_cell_6t_5 inst_cell_58_44 (.BL(BL44),.BLN(BLN44),.WL(WL58));
sram_cell_6t_5 inst_cell_58_45 (.BL(BL45),.BLN(BLN45),.WL(WL58));
sram_cell_6t_5 inst_cell_58_46 (.BL(BL46),.BLN(BLN46),.WL(WL58));
sram_cell_6t_5 inst_cell_58_47 (.BL(BL47),.BLN(BLN47),.WL(WL58));
sram_cell_6t_5 inst_cell_58_48 (.BL(BL48),.BLN(BLN48),.WL(WL58));
sram_cell_6t_5 inst_cell_58_49 (.BL(BL49),.BLN(BLN49),.WL(WL58));
sram_cell_6t_5 inst_cell_58_50 (.BL(BL50),.BLN(BLN50),.WL(WL58));
sram_cell_6t_5 inst_cell_58_51 (.BL(BL51),.BLN(BLN51),.WL(WL58));
sram_cell_6t_5 inst_cell_58_52 (.BL(BL52),.BLN(BLN52),.WL(WL58));
sram_cell_6t_5 inst_cell_58_53 (.BL(BL53),.BLN(BLN53),.WL(WL58));
sram_cell_6t_5 inst_cell_58_54 (.BL(BL54),.BLN(BLN54),.WL(WL58));
sram_cell_6t_5 inst_cell_58_55 (.BL(BL55),.BLN(BLN55),.WL(WL58));
sram_cell_6t_5 inst_cell_58_56 (.BL(BL56),.BLN(BLN56),.WL(WL58));
sram_cell_6t_5 inst_cell_58_57 (.BL(BL57),.BLN(BLN57),.WL(WL58));
sram_cell_6t_5 inst_cell_58_58 (.BL(BL58),.BLN(BLN58),.WL(WL58));
sram_cell_6t_5 inst_cell_58_59 (.BL(BL59),.BLN(BLN59),.WL(WL58));
sram_cell_6t_5 inst_cell_58_60 (.BL(BL60),.BLN(BLN60),.WL(WL58));
sram_cell_6t_5 inst_cell_58_61 (.BL(BL61),.BLN(BLN61),.WL(WL58));
sram_cell_6t_5 inst_cell_58_62 (.BL(BL62),.BLN(BLN62),.WL(WL58));
sram_cell_6t_5 inst_cell_58_63 (.BL(BL63),.BLN(BLN63),.WL(WL58));
sram_cell_6t_5 inst_cell_58_64 (.BL(BL64),.BLN(BLN64),.WL(WL58));
sram_cell_6t_5 inst_cell_58_65 (.BL(BL65),.BLN(BLN65),.WL(WL58));
sram_cell_6t_5 inst_cell_58_66 (.BL(BL66),.BLN(BLN66),.WL(WL58));
sram_cell_6t_5 inst_cell_58_67 (.BL(BL67),.BLN(BLN67),.WL(WL58));
sram_cell_6t_5 inst_cell_58_68 (.BL(BL68),.BLN(BLN68),.WL(WL58));
sram_cell_6t_5 inst_cell_58_69 (.BL(BL69),.BLN(BLN69),.WL(WL58));
sram_cell_6t_5 inst_cell_58_70 (.BL(BL70),.BLN(BLN70),.WL(WL58));
sram_cell_6t_5 inst_cell_58_71 (.BL(BL71),.BLN(BLN71),.WL(WL58));
sram_cell_6t_5 inst_cell_58_72 (.BL(BL72),.BLN(BLN72),.WL(WL58));
sram_cell_6t_5 inst_cell_58_73 (.BL(BL73),.BLN(BLN73),.WL(WL58));
sram_cell_6t_5 inst_cell_58_74 (.BL(BL74),.BLN(BLN74),.WL(WL58));
sram_cell_6t_5 inst_cell_58_75 (.BL(BL75),.BLN(BLN75),.WL(WL58));
sram_cell_6t_5 inst_cell_58_76 (.BL(BL76),.BLN(BLN76),.WL(WL58));
sram_cell_6t_5 inst_cell_58_77 (.BL(BL77),.BLN(BLN77),.WL(WL58));
sram_cell_6t_5 inst_cell_58_78 (.BL(BL78),.BLN(BLN78),.WL(WL58));
sram_cell_6t_5 inst_cell_58_79 (.BL(BL79),.BLN(BLN79),.WL(WL58));
sram_cell_6t_5 inst_cell_58_80 (.BL(BL80),.BLN(BLN80),.WL(WL58));
sram_cell_6t_5 inst_cell_58_81 (.BL(BL81),.BLN(BLN81),.WL(WL58));
sram_cell_6t_5 inst_cell_58_82 (.BL(BL82),.BLN(BLN82),.WL(WL58));
sram_cell_6t_5 inst_cell_58_83 (.BL(BL83),.BLN(BLN83),.WL(WL58));
sram_cell_6t_5 inst_cell_58_84 (.BL(BL84),.BLN(BLN84),.WL(WL58));
sram_cell_6t_5 inst_cell_58_85 (.BL(BL85),.BLN(BLN85),.WL(WL58));
sram_cell_6t_5 inst_cell_58_86 (.BL(BL86),.BLN(BLN86),.WL(WL58));
sram_cell_6t_5 inst_cell_58_87 (.BL(BL87),.BLN(BLN87),.WL(WL58));
sram_cell_6t_5 inst_cell_58_88 (.BL(BL88),.BLN(BLN88),.WL(WL58));
sram_cell_6t_5 inst_cell_58_89 (.BL(BL89),.BLN(BLN89),.WL(WL58));
sram_cell_6t_5 inst_cell_58_90 (.BL(BL90),.BLN(BLN90),.WL(WL58));
sram_cell_6t_5 inst_cell_58_91 (.BL(BL91),.BLN(BLN91),.WL(WL58));
sram_cell_6t_5 inst_cell_58_92 (.BL(BL92),.BLN(BLN92),.WL(WL58));
sram_cell_6t_5 inst_cell_58_93 (.BL(BL93),.BLN(BLN93),.WL(WL58));
sram_cell_6t_5 inst_cell_58_94 (.BL(BL94),.BLN(BLN94),.WL(WL58));
sram_cell_6t_5 inst_cell_58_95 (.BL(BL95),.BLN(BLN95),.WL(WL58));
sram_cell_6t_5 inst_cell_58_96 (.BL(BL96),.BLN(BLN96),.WL(WL58));
sram_cell_6t_5 inst_cell_58_97 (.BL(BL97),.BLN(BLN97),.WL(WL58));
sram_cell_6t_5 inst_cell_58_98 (.BL(BL98),.BLN(BLN98),.WL(WL58));
sram_cell_6t_5 inst_cell_58_99 (.BL(BL99),.BLN(BLN99),.WL(WL58));
sram_cell_6t_5 inst_cell_58_100 (.BL(BL100),.BLN(BLN100),.WL(WL58));
sram_cell_6t_5 inst_cell_58_101 (.BL(BL101),.BLN(BLN101),.WL(WL58));
sram_cell_6t_5 inst_cell_58_102 (.BL(BL102),.BLN(BLN102),.WL(WL58));
sram_cell_6t_5 inst_cell_58_103 (.BL(BL103),.BLN(BLN103),.WL(WL58));
sram_cell_6t_5 inst_cell_58_104 (.BL(BL104),.BLN(BLN104),.WL(WL58));
sram_cell_6t_5 inst_cell_58_105 (.BL(BL105),.BLN(BLN105),.WL(WL58));
sram_cell_6t_5 inst_cell_58_106 (.BL(BL106),.BLN(BLN106),.WL(WL58));
sram_cell_6t_5 inst_cell_58_107 (.BL(BL107),.BLN(BLN107),.WL(WL58));
sram_cell_6t_5 inst_cell_58_108 (.BL(BL108),.BLN(BLN108),.WL(WL58));
sram_cell_6t_5 inst_cell_58_109 (.BL(BL109),.BLN(BLN109),.WL(WL58));
sram_cell_6t_5 inst_cell_58_110 (.BL(BL110),.BLN(BLN110),.WL(WL58));
sram_cell_6t_5 inst_cell_58_111 (.BL(BL111),.BLN(BLN111),.WL(WL58));
sram_cell_6t_5 inst_cell_58_112 (.BL(BL112),.BLN(BLN112),.WL(WL58));
sram_cell_6t_5 inst_cell_58_113 (.BL(BL113),.BLN(BLN113),.WL(WL58));
sram_cell_6t_5 inst_cell_58_114 (.BL(BL114),.BLN(BLN114),.WL(WL58));
sram_cell_6t_5 inst_cell_58_115 (.BL(BL115),.BLN(BLN115),.WL(WL58));
sram_cell_6t_5 inst_cell_58_116 (.BL(BL116),.BLN(BLN116),.WL(WL58));
sram_cell_6t_5 inst_cell_58_117 (.BL(BL117),.BLN(BLN117),.WL(WL58));
sram_cell_6t_5 inst_cell_58_118 (.BL(BL118),.BLN(BLN118),.WL(WL58));
sram_cell_6t_5 inst_cell_58_119 (.BL(BL119),.BLN(BLN119),.WL(WL58));
sram_cell_6t_5 inst_cell_58_120 (.BL(BL120),.BLN(BLN120),.WL(WL58));
sram_cell_6t_5 inst_cell_58_121 (.BL(BL121),.BLN(BLN121),.WL(WL58));
sram_cell_6t_5 inst_cell_58_122 (.BL(BL122),.BLN(BLN122),.WL(WL58));
sram_cell_6t_5 inst_cell_58_123 (.BL(BL123),.BLN(BLN123),.WL(WL58));
sram_cell_6t_5 inst_cell_58_124 (.BL(BL124),.BLN(BLN124),.WL(WL58));
sram_cell_6t_5 inst_cell_58_125 (.BL(BL125),.BLN(BLN125),.WL(WL58));
sram_cell_6t_5 inst_cell_58_126 (.BL(BL126),.BLN(BLN126),.WL(WL58));
sram_cell_6t_5 inst_cell_58_127 (.BL(BL127),.BLN(BLN127),.WL(WL58));
sram_cell_6t_5 inst_cell_59_0 (.BL(BL0),.BLN(BLN0),.WL(WL59));
sram_cell_6t_5 inst_cell_59_1 (.BL(BL1),.BLN(BLN1),.WL(WL59));
sram_cell_6t_5 inst_cell_59_2 (.BL(BL2),.BLN(BLN2),.WL(WL59));
sram_cell_6t_5 inst_cell_59_3 (.BL(BL3),.BLN(BLN3),.WL(WL59));
sram_cell_6t_5 inst_cell_59_4 (.BL(BL4),.BLN(BLN4),.WL(WL59));
sram_cell_6t_5 inst_cell_59_5 (.BL(BL5),.BLN(BLN5),.WL(WL59));
sram_cell_6t_5 inst_cell_59_6 (.BL(BL6),.BLN(BLN6),.WL(WL59));
sram_cell_6t_5 inst_cell_59_7 (.BL(BL7),.BLN(BLN7),.WL(WL59));
sram_cell_6t_5 inst_cell_59_8 (.BL(BL8),.BLN(BLN8),.WL(WL59));
sram_cell_6t_5 inst_cell_59_9 (.BL(BL9),.BLN(BLN9),.WL(WL59));
sram_cell_6t_5 inst_cell_59_10 (.BL(BL10),.BLN(BLN10),.WL(WL59));
sram_cell_6t_5 inst_cell_59_11 (.BL(BL11),.BLN(BLN11),.WL(WL59));
sram_cell_6t_5 inst_cell_59_12 (.BL(BL12),.BLN(BLN12),.WL(WL59));
sram_cell_6t_5 inst_cell_59_13 (.BL(BL13),.BLN(BLN13),.WL(WL59));
sram_cell_6t_5 inst_cell_59_14 (.BL(BL14),.BLN(BLN14),.WL(WL59));
sram_cell_6t_5 inst_cell_59_15 (.BL(BL15),.BLN(BLN15),.WL(WL59));
sram_cell_6t_5 inst_cell_59_16 (.BL(BL16),.BLN(BLN16),.WL(WL59));
sram_cell_6t_5 inst_cell_59_17 (.BL(BL17),.BLN(BLN17),.WL(WL59));
sram_cell_6t_5 inst_cell_59_18 (.BL(BL18),.BLN(BLN18),.WL(WL59));
sram_cell_6t_5 inst_cell_59_19 (.BL(BL19),.BLN(BLN19),.WL(WL59));
sram_cell_6t_5 inst_cell_59_20 (.BL(BL20),.BLN(BLN20),.WL(WL59));
sram_cell_6t_5 inst_cell_59_21 (.BL(BL21),.BLN(BLN21),.WL(WL59));
sram_cell_6t_5 inst_cell_59_22 (.BL(BL22),.BLN(BLN22),.WL(WL59));
sram_cell_6t_5 inst_cell_59_23 (.BL(BL23),.BLN(BLN23),.WL(WL59));
sram_cell_6t_5 inst_cell_59_24 (.BL(BL24),.BLN(BLN24),.WL(WL59));
sram_cell_6t_5 inst_cell_59_25 (.BL(BL25),.BLN(BLN25),.WL(WL59));
sram_cell_6t_5 inst_cell_59_26 (.BL(BL26),.BLN(BLN26),.WL(WL59));
sram_cell_6t_5 inst_cell_59_27 (.BL(BL27),.BLN(BLN27),.WL(WL59));
sram_cell_6t_5 inst_cell_59_28 (.BL(BL28),.BLN(BLN28),.WL(WL59));
sram_cell_6t_5 inst_cell_59_29 (.BL(BL29),.BLN(BLN29),.WL(WL59));
sram_cell_6t_5 inst_cell_59_30 (.BL(BL30),.BLN(BLN30),.WL(WL59));
sram_cell_6t_5 inst_cell_59_31 (.BL(BL31),.BLN(BLN31),.WL(WL59));
sram_cell_6t_5 inst_cell_59_32 (.BL(BL32),.BLN(BLN32),.WL(WL59));
sram_cell_6t_5 inst_cell_59_33 (.BL(BL33),.BLN(BLN33),.WL(WL59));
sram_cell_6t_5 inst_cell_59_34 (.BL(BL34),.BLN(BLN34),.WL(WL59));
sram_cell_6t_5 inst_cell_59_35 (.BL(BL35),.BLN(BLN35),.WL(WL59));
sram_cell_6t_5 inst_cell_59_36 (.BL(BL36),.BLN(BLN36),.WL(WL59));
sram_cell_6t_5 inst_cell_59_37 (.BL(BL37),.BLN(BLN37),.WL(WL59));
sram_cell_6t_5 inst_cell_59_38 (.BL(BL38),.BLN(BLN38),.WL(WL59));
sram_cell_6t_5 inst_cell_59_39 (.BL(BL39),.BLN(BLN39),.WL(WL59));
sram_cell_6t_5 inst_cell_59_40 (.BL(BL40),.BLN(BLN40),.WL(WL59));
sram_cell_6t_5 inst_cell_59_41 (.BL(BL41),.BLN(BLN41),.WL(WL59));
sram_cell_6t_5 inst_cell_59_42 (.BL(BL42),.BLN(BLN42),.WL(WL59));
sram_cell_6t_5 inst_cell_59_43 (.BL(BL43),.BLN(BLN43),.WL(WL59));
sram_cell_6t_5 inst_cell_59_44 (.BL(BL44),.BLN(BLN44),.WL(WL59));
sram_cell_6t_5 inst_cell_59_45 (.BL(BL45),.BLN(BLN45),.WL(WL59));
sram_cell_6t_5 inst_cell_59_46 (.BL(BL46),.BLN(BLN46),.WL(WL59));
sram_cell_6t_5 inst_cell_59_47 (.BL(BL47),.BLN(BLN47),.WL(WL59));
sram_cell_6t_5 inst_cell_59_48 (.BL(BL48),.BLN(BLN48),.WL(WL59));
sram_cell_6t_5 inst_cell_59_49 (.BL(BL49),.BLN(BLN49),.WL(WL59));
sram_cell_6t_5 inst_cell_59_50 (.BL(BL50),.BLN(BLN50),.WL(WL59));
sram_cell_6t_5 inst_cell_59_51 (.BL(BL51),.BLN(BLN51),.WL(WL59));
sram_cell_6t_5 inst_cell_59_52 (.BL(BL52),.BLN(BLN52),.WL(WL59));
sram_cell_6t_5 inst_cell_59_53 (.BL(BL53),.BLN(BLN53),.WL(WL59));
sram_cell_6t_5 inst_cell_59_54 (.BL(BL54),.BLN(BLN54),.WL(WL59));
sram_cell_6t_5 inst_cell_59_55 (.BL(BL55),.BLN(BLN55),.WL(WL59));
sram_cell_6t_5 inst_cell_59_56 (.BL(BL56),.BLN(BLN56),.WL(WL59));
sram_cell_6t_5 inst_cell_59_57 (.BL(BL57),.BLN(BLN57),.WL(WL59));
sram_cell_6t_5 inst_cell_59_58 (.BL(BL58),.BLN(BLN58),.WL(WL59));
sram_cell_6t_5 inst_cell_59_59 (.BL(BL59),.BLN(BLN59),.WL(WL59));
sram_cell_6t_5 inst_cell_59_60 (.BL(BL60),.BLN(BLN60),.WL(WL59));
sram_cell_6t_5 inst_cell_59_61 (.BL(BL61),.BLN(BLN61),.WL(WL59));
sram_cell_6t_5 inst_cell_59_62 (.BL(BL62),.BLN(BLN62),.WL(WL59));
sram_cell_6t_5 inst_cell_59_63 (.BL(BL63),.BLN(BLN63),.WL(WL59));
sram_cell_6t_5 inst_cell_59_64 (.BL(BL64),.BLN(BLN64),.WL(WL59));
sram_cell_6t_5 inst_cell_59_65 (.BL(BL65),.BLN(BLN65),.WL(WL59));
sram_cell_6t_5 inst_cell_59_66 (.BL(BL66),.BLN(BLN66),.WL(WL59));
sram_cell_6t_5 inst_cell_59_67 (.BL(BL67),.BLN(BLN67),.WL(WL59));
sram_cell_6t_5 inst_cell_59_68 (.BL(BL68),.BLN(BLN68),.WL(WL59));
sram_cell_6t_5 inst_cell_59_69 (.BL(BL69),.BLN(BLN69),.WL(WL59));
sram_cell_6t_5 inst_cell_59_70 (.BL(BL70),.BLN(BLN70),.WL(WL59));
sram_cell_6t_5 inst_cell_59_71 (.BL(BL71),.BLN(BLN71),.WL(WL59));
sram_cell_6t_5 inst_cell_59_72 (.BL(BL72),.BLN(BLN72),.WL(WL59));
sram_cell_6t_5 inst_cell_59_73 (.BL(BL73),.BLN(BLN73),.WL(WL59));
sram_cell_6t_5 inst_cell_59_74 (.BL(BL74),.BLN(BLN74),.WL(WL59));
sram_cell_6t_5 inst_cell_59_75 (.BL(BL75),.BLN(BLN75),.WL(WL59));
sram_cell_6t_5 inst_cell_59_76 (.BL(BL76),.BLN(BLN76),.WL(WL59));
sram_cell_6t_5 inst_cell_59_77 (.BL(BL77),.BLN(BLN77),.WL(WL59));
sram_cell_6t_5 inst_cell_59_78 (.BL(BL78),.BLN(BLN78),.WL(WL59));
sram_cell_6t_5 inst_cell_59_79 (.BL(BL79),.BLN(BLN79),.WL(WL59));
sram_cell_6t_5 inst_cell_59_80 (.BL(BL80),.BLN(BLN80),.WL(WL59));
sram_cell_6t_5 inst_cell_59_81 (.BL(BL81),.BLN(BLN81),.WL(WL59));
sram_cell_6t_5 inst_cell_59_82 (.BL(BL82),.BLN(BLN82),.WL(WL59));
sram_cell_6t_5 inst_cell_59_83 (.BL(BL83),.BLN(BLN83),.WL(WL59));
sram_cell_6t_5 inst_cell_59_84 (.BL(BL84),.BLN(BLN84),.WL(WL59));
sram_cell_6t_5 inst_cell_59_85 (.BL(BL85),.BLN(BLN85),.WL(WL59));
sram_cell_6t_5 inst_cell_59_86 (.BL(BL86),.BLN(BLN86),.WL(WL59));
sram_cell_6t_5 inst_cell_59_87 (.BL(BL87),.BLN(BLN87),.WL(WL59));
sram_cell_6t_5 inst_cell_59_88 (.BL(BL88),.BLN(BLN88),.WL(WL59));
sram_cell_6t_5 inst_cell_59_89 (.BL(BL89),.BLN(BLN89),.WL(WL59));
sram_cell_6t_5 inst_cell_59_90 (.BL(BL90),.BLN(BLN90),.WL(WL59));
sram_cell_6t_5 inst_cell_59_91 (.BL(BL91),.BLN(BLN91),.WL(WL59));
sram_cell_6t_5 inst_cell_59_92 (.BL(BL92),.BLN(BLN92),.WL(WL59));
sram_cell_6t_5 inst_cell_59_93 (.BL(BL93),.BLN(BLN93),.WL(WL59));
sram_cell_6t_5 inst_cell_59_94 (.BL(BL94),.BLN(BLN94),.WL(WL59));
sram_cell_6t_5 inst_cell_59_95 (.BL(BL95),.BLN(BLN95),.WL(WL59));
sram_cell_6t_5 inst_cell_59_96 (.BL(BL96),.BLN(BLN96),.WL(WL59));
sram_cell_6t_5 inst_cell_59_97 (.BL(BL97),.BLN(BLN97),.WL(WL59));
sram_cell_6t_5 inst_cell_59_98 (.BL(BL98),.BLN(BLN98),.WL(WL59));
sram_cell_6t_5 inst_cell_59_99 (.BL(BL99),.BLN(BLN99),.WL(WL59));
sram_cell_6t_5 inst_cell_59_100 (.BL(BL100),.BLN(BLN100),.WL(WL59));
sram_cell_6t_5 inst_cell_59_101 (.BL(BL101),.BLN(BLN101),.WL(WL59));
sram_cell_6t_5 inst_cell_59_102 (.BL(BL102),.BLN(BLN102),.WL(WL59));
sram_cell_6t_5 inst_cell_59_103 (.BL(BL103),.BLN(BLN103),.WL(WL59));
sram_cell_6t_5 inst_cell_59_104 (.BL(BL104),.BLN(BLN104),.WL(WL59));
sram_cell_6t_5 inst_cell_59_105 (.BL(BL105),.BLN(BLN105),.WL(WL59));
sram_cell_6t_5 inst_cell_59_106 (.BL(BL106),.BLN(BLN106),.WL(WL59));
sram_cell_6t_5 inst_cell_59_107 (.BL(BL107),.BLN(BLN107),.WL(WL59));
sram_cell_6t_5 inst_cell_59_108 (.BL(BL108),.BLN(BLN108),.WL(WL59));
sram_cell_6t_5 inst_cell_59_109 (.BL(BL109),.BLN(BLN109),.WL(WL59));
sram_cell_6t_5 inst_cell_59_110 (.BL(BL110),.BLN(BLN110),.WL(WL59));
sram_cell_6t_5 inst_cell_59_111 (.BL(BL111),.BLN(BLN111),.WL(WL59));
sram_cell_6t_5 inst_cell_59_112 (.BL(BL112),.BLN(BLN112),.WL(WL59));
sram_cell_6t_5 inst_cell_59_113 (.BL(BL113),.BLN(BLN113),.WL(WL59));
sram_cell_6t_5 inst_cell_59_114 (.BL(BL114),.BLN(BLN114),.WL(WL59));
sram_cell_6t_5 inst_cell_59_115 (.BL(BL115),.BLN(BLN115),.WL(WL59));
sram_cell_6t_5 inst_cell_59_116 (.BL(BL116),.BLN(BLN116),.WL(WL59));
sram_cell_6t_5 inst_cell_59_117 (.BL(BL117),.BLN(BLN117),.WL(WL59));
sram_cell_6t_5 inst_cell_59_118 (.BL(BL118),.BLN(BLN118),.WL(WL59));
sram_cell_6t_5 inst_cell_59_119 (.BL(BL119),.BLN(BLN119),.WL(WL59));
sram_cell_6t_5 inst_cell_59_120 (.BL(BL120),.BLN(BLN120),.WL(WL59));
sram_cell_6t_5 inst_cell_59_121 (.BL(BL121),.BLN(BLN121),.WL(WL59));
sram_cell_6t_5 inst_cell_59_122 (.BL(BL122),.BLN(BLN122),.WL(WL59));
sram_cell_6t_5 inst_cell_59_123 (.BL(BL123),.BLN(BLN123),.WL(WL59));
sram_cell_6t_5 inst_cell_59_124 (.BL(BL124),.BLN(BLN124),.WL(WL59));
sram_cell_6t_5 inst_cell_59_125 (.BL(BL125),.BLN(BLN125),.WL(WL59));
sram_cell_6t_5 inst_cell_59_126 (.BL(BL126),.BLN(BLN126),.WL(WL59));
sram_cell_6t_5 inst_cell_59_127 (.BL(BL127),.BLN(BLN127),.WL(WL59));
sram_cell_6t_5 inst_cell_60_0 (.BL(BL0),.BLN(BLN0),.WL(WL60));
sram_cell_6t_5 inst_cell_60_1 (.BL(BL1),.BLN(BLN1),.WL(WL60));
sram_cell_6t_5 inst_cell_60_2 (.BL(BL2),.BLN(BLN2),.WL(WL60));
sram_cell_6t_5 inst_cell_60_3 (.BL(BL3),.BLN(BLN3),.WL(WL60));
sram_cell_6t_5 inst_cell_60_4 (.BL(BL4),.BLN(BLN4),.WL(WL60));
sram_cell_6t_5 inst_cell_60_5 (.BL(BL5),.BLN(BLN5),.WL(WL60));
sram_cell_6t_5 inst_cell_60_6 (.BL(BL6),.BLN(BLN6),.WL(WL60));
sram_cell_6t_5 inst_cell_60_7 (.BL(BL7),.BLN(BLN7),.WL(WL60));
sram_cell_6t_5 inst_cell_60_8 (.BL(BL8),.BLN(BLN8),.WL(WL60));
sram_cell_6t_5 inst_cell_60_9 (.BL(BL9),.BLN(BLN9),.WL(WL60));
sram_cell_6t_5 inst_cell_60_10 (.BL(BL10),.BLN(BLN10),.WL(WL60));
sram_cell_6t_5 inst_cell_60_11 (.BL(BL11),.BLN(BLN11),.WL(WL60));
sram_cell_6t_5 inst_cell_60_12 (.BL(BL12),.BLN(BLN12),.WL(WL60));
sram_cell_6t_5 inst_cell_60_13 (.BL(BL13),.BLN(BLN13),.WL(WL60));
sram_cell_6t_5 inst_cell_60_14 (.BL(BL14),.BLN(BLN14),.WL(WL60));
sram_cell_6t_5 inst_cell_60_15 (.BL(BL15),.BLN(BLN15),.WL(WL60));
sram_cell_6t_5 inst_cell_60_16 (.BL(BL16),.BLN(BLN16),.WL(WL60));
sram_cell_6t_5 inst_cell_60_17 (.BL(BL17),.BLN(BLN17),.WL(WL60));
sram_cell_6t_5 inst_cell_60_18 (.BL(BL18),.BLN(BLN18),.WL(WL60));
sram_cell_6t_5 inst_cell_60_19 (.BL(BL19),.BLN(BLN19),.WL(WL60));
sram_cell_6t_5 inst_cell_60_20 (.BL(BL20),.BLN(BLN20),.WL(WL60));
sram_cell_6t_5 inst_cell_60_21 (.BL(BL21),.BLN(BLN21),.WL(WL60));
sram_cell_6t_5 inst_cell_60_22 (.BL(BL22),.BLN(BLN22),.WL(WL60));
sram_cell_6t_5 inst_cell_60_23 (.BL(BL23),.BLN(BLN23),.WL(WL60));
sram_cell_6t_5 inst_cell_60_24 (.BL(BL24),.BLN(BLN24),.WL(WL60));
sram_cell_6t_5 inst_cell_60_25 (.BL(BL25),.BLN(BLN25),.WL(WL60));
sram_cell_6t_5 inst_cell_60_26 (.BL(BL26),.BLN(BLN26),.WL(WL60));
sram_cell_6t_5 inst_cell_60_27 (.BL(BL27),.BLN(BLN27),.WL(WL60));
sram_cell_6t_5 inst_cell_60_28 (.BL(BL28),.BLN(BLN28),.WL(WL60));
sram_cell_6t_5 inst_cell_60_29 (.BL(BL29),.BLN(BLN29),.WL(WL60));
sram_cell_6t_5 inst_cell_60_30 (.BL(BL30),.BLN(BLN30),.WL(WL60));
sram_cell_6t_5 inst_cell_60_31 (.BL(BL31),.BLN(BLN31),.WL(WL60));
sram_cell_6t_5 inst_cell_60_32 (.BL(BL32),.BLN(BLN32),.WL(WL60));
sram_cell_6t_5 inst_cell_60_33 (.BL(BL33),.BLN(BLN33),.WL(WL60));
sram_cell_6t_5 inst_cell_60_34 (.BL(BL34),.BLN(BLN34),.WL(WL60));
sram_cell_6t_5 inst_cell_60_35 (.BL(BL35),.BLN(BLN35),.WL(WL60));
sram_cell_6t_5 inst_cell_60_36 (.BL(BL36),.BLN(BLN36),.WL(WL60));
sram_cell_6t_5 inst_cell_60_37 (.BL(BL37),.BLN(BLN37),.WL(WL60));
sram_cell_6t_5 inst_cell_60_38 (.BL(BL38),.BLN(BLN38),.WL(WL60));
sram_cell_6t_5 inst_cell_60_39 (.BL(BL39),.BLN(BLN39),.WL(WL60));
sram_cell_6t_5 inst_cell_60_40 (.BL(BL40),.BLN(BLN40),.WL(WL60));
sram_cell_6t_5 inst_cell_60_41 (.BL(BL41),.BLN(BLN41),.WL(WL60));
sram_cell_6t_5 inst_cell_60_42 (.BL(BL42),.BLN(BLN42),.WL(WL60));
sram_cell_6t_5 inst_cell_60_43 (.BL(BL43),.BLN(BLN43),.WL(WL60));
sram_cell_6t_5 inst_cell_60_44 (.BL(BL44),.BLN(BLN44),.WL(WL60));
sram_cell_6t_5 inst_cell_60_45 (.BL(BL45),.BLN(BLN45),.WL(WL60));
sram_cell_6t_5 inst_cell_60_46 (.BL(BL46),.BLN(BLN46),.WL(WL60));
sram_cell_6t_5 inst_cell_60_47 (.BL(BL47),.BLN(BLN47),.WL(WL60));
sram_cell_6t_5 inst_cell_60_48 (.BL(BL48),.BLN(BLN48),.WL(WL60));
sram_cell_6t_5 inst_cell_60_49 (.BL(BL49),.BLN(BLN49),.WL(WL60));
sram_cell_6t_5 inst_cell_60_50 (.BL(BL50),.BLN(BLN50),.WL(WL60));
sram_cell_6t_5 inst_cell_60_51 (.BL(BL51),.BLN(BLN51),.WL(WL60));
sram_cell_6t_5 inst_cell_60_52 (.BL(BL52),.BLN(BLN52),.WL(WL60));
sram_cell_6t_5 inst_cell_60_53 (.BL(BL53),.BLN(BLN53),.WL(WL60));
sram_cell_6t_5 inst_cell_60_54 (.BL(BL54),.BLN(BLN54),.WL(WL60));
sram_cell_6t_5 inst_cell_60_55 (.BL(BL55),.BLN(BLN55),.WL(WL60));
sram_cell_6t_5 inst_cell_60_56 (.BL(BL56),.BLN(BLN56),.WL(WL60));
sram_cell_6t_5 inst_cell_60_57 (.BL(BL57),.BLN(BLN57),.WL(WL60));
sram_cell_6t_5 inst_cell_60_58 (.BL(BL58),.BLN(BLN58),.WL(WL60));
sram_cell_6t_5 inst_cell_60_59 (.BL(BL59),.BLN(BLN59),.WL(WL60));
sram_cell_6t_5 inst_cell_60_60 (.BL(BL60),.BLN(BLN60),.WL(WL60));
sram_cell_6t_5 inst_cell_60_61 (.BL(BL61),.BLN(BLN61),.WL(WL60));
sram_cell_6t_5 inst_cell_60_62 (.BL(BL62),.BLN(BLN62),.WL(WL60));
sram_cell_6t_5 inst_cell_60_63 (.BL(BL63),.BLN(BLN63),.WL(WL60));
sram_cell_6t_5 inst_cell_60_64 (.BL(BL64),.BLN(BLN64),.WL(WL60));
sram_cell_6t_5 inst_cell_60_65 (.BL(BL65),.BLN(BLN65),.WL(WL60));
sram_cell_6t_5 inst_cell_60_66 (.BL(BL66),.BLN(BLN66),.WL(WL60));
sram_cell_6t_5 inst_cell_60_67 (.BL(BL67),.BLN(BLN67),.WL(WL60));
sram_cell_6t_5 inst_cell_60_68 (.BL(BL68),.BLN(BLN68),.WL(WL60));
sram_cell_6t_5 inst_cell_60_69 (.BL(BL69),.BLN(BLN69),.WL(WL60));
sram_cell_6t_5 inst_cell_60_70 (.BL(BL70),.BLN(BLN70),.WL(WL60));
sram_cell_6t_5 inst_cell_60_71 (.BL(BL71),.BLN(BLN71),.WL(WL60));
sram_cell_6t_5 inst_cell_60_72 (.BL(BL72),.BLN(BLN72),.WL(WL60));
sram_cell_6t_5 inst_cell_60_73 (.BL(BL73),.BLN(BLN73),.WL(WL60));
sram_cell_6t_5 inst_cell_60_74 (.BL(BL74),.BLN(BLN74),.WL(WL60));
sram_cell_6t_5 inst_cell_60_75 (.BL(BL75),.BLN(BLN75),.WL(WL60));
sram_cell_6t_5 inst_cell_60_76 (.BL(BL76),.BLN(BLN76),.WL(WL60));
sram_cell_6t_5 inst_cell_60_77 (.BL(BL77),.BLN(BLN77),.WL(WL60));
sram_cell_6t_5 inst_cell_60_78 (.BL(BL78),.BLN(BLN78),.WL(WL60));
sram_cell_6t_5 inst_cell_60_79 (.BL(BL79),.BLN(BLN79),.WL(WL60));
sram_cell_6t_5 inst_cell_60_80 (.BL(BL80),.BLN(BLN80),.WL(WL60));
sram_cell_6t_5 inst_cell_60_81 (.BL(BL81),.BLN(BLN81),.WL(WL60));
sram_cell_6t_5 inst_cell_60_82 (.BL(BL82),.BLN(BLN82),.WL(WL60));
sram_cell_6t_5 inst_cell_60_83 (.BL(BL83),.BLN(BLN83),.WL(WL60));
sram_cell_6t_5 inst_cell_60_84 (.BL(BL84),.BLN(BLN84),.WL(WL60));
sram_cell_6t_5 inst_cell_60_85 (.BL(BL85),.BLN(BLN85),.WL(WL60));
sram_cell_6t_5 inst_cell_60_86 (.BL(BL86),.BLN(BLN86),.WL(WL60));
sram_cell_6t_5 inst_cell_60_87 (.BL(BL87),.BLN(BLN87),.WL(WL60));
sram_cell_6t_5 inst_cell_60_88 (.BL(BL88),.BLN(BLN88),.WL(WL60));
sram_cell_6t_5 inst_cell_60_89 (.BL(BL89),.BLN(BLN89),.WL(WL60));
sram_cell_6t_5 inst_cell_60_90 (.BL(BL90),.BLN(BLN90),.WL(WL60));
sram_cell_6t_5 inst_cell_60_91 (.BL(BL91),.BLN(BLN91),.WL(WL60));
sram_cell_6t_5 inst_cell_60_92 (.BL(BL92),.BLN(BLN92),.WL(WL60));
sram_cell_6t_5 inst_cell_60_93 (.BL(BL93),.BLN(BLN93),.WL(WL60));
sram_cell_6t_5 inst_cell_60_94 (.BL(BL94),.BLN(BLN94),.WL(WL60));
sram_cell_6t_5 inst_cell_60_95 (.BL(BL95),.BLN(BLN95),.WL(WL60));
sram_cell_6t_5 inst_cell_60_96 (.BL(BL96),.BLN(BLN96),.WL(WL60));
sram_cell_6t_5 inst_cell_60_97 (.BL(BL97),.BLN(BLN97),.WL(WL60));
sram_cell_6t_5 inst_cell_60_98 (.BL(BL98),.BLN(BLN98),.WL(WL60));
sram_cell_6t_5 inst_cell_60_99 (.BL(BL99),.BLN(BLN99),.WL(WL60));
sram_cell_6t_5 inst_cell_60_100 (.BL(BL100),.BLN(BLN100),.WL(WL60));
sram_cell_6t_5 inst_cell_60_101 (.BL(BL101),.BLN(BLN101),.WL(WL60));
sram_cell_6t_5 inst_cell_60_102 (.BL(BL102),.BLN(BLN102),.WL(WL60));
sram_cell_6t_5 inst_cell_60_103 (.BL(BL103),.BLN(BLN103),.WL(WL60));
sram_cell_6t_5 inst_cell_60_104 (.BL(BL104),.BLN(BLN104),.WL(WL60));
sram_cell_6t_5 inst_cell_60_105 (.BL(BL105),.BLN(BLN105),.WL(WL60));
sram_cell_6t_5 inst_cell_60_106 (.BL(BL106),.BLN(BLN106),.WL(WL60));
sram_cell_6t_5 inst_cell_60_107 (.BL(BL107),.BLN(BLN107),.WL(WL60));
sram_cell_6t_5 inst_cell_60_108 (.BL(BL108),.BLN(BLN108),.WL(WL60));
sram_cell_6t_5 inst_cell_60_109 (.BL(BL109),.BLN(BLN109),.WL(WL60));
sram_cell_6t_5 inst_cell_60_110 (.BL(BL110),.BLN(BLN110),.WL(WL60));
sram_cell_6t_5 inst_cell_60_111 (.BL(BL111),.BLN(BLN111),.WL(WL60));
sram_cell_6t_5 inst_cell_60_112 (.BL(BL112),.BLN(BLN112),.WL(WL60));
sram_cell_6t_5 inst_cell_60_113 (.BL(BL113),.BLN(BLN113),.WL(WL60));
sram_cell_6t_5 inst_cell_60_114 (.BL(BL114),.BLN(BLN114),.WL(WL60));
sram_cell_6t_5 inst_cell_60_115 (.BL(BL115),.BLN(BLN115),.WL(WL60));
sram_cell_6t_5 inst_cell_60_116 (.BL(BL116),.BLN(BLN116),.WL(WL60));
sram_cell_6t_5 inst_cell_60_117 (.BL(BL117),.BLN(BLN117),.WL(WL60));
sram_cell_6t_5 inst_cell_60_118 (.BL(BL118),.BLN(BLN118),.WL(WL60));
sram_cell_6t_5 inst_cell_60_119 (.BL(BL119),.BLN(BLN119),.WL(WL60));
sram_cell_6t_5 inst_cell_60_120 (.BL(BL120),.BLN(BLN120),.WL(WL60));
sram_cell_6t_5 inst_cell_60_121 (.BL(BL121),.BLN(BLN121),.WL(WL60));
sram_cell_6t_5 inst_cell_60_122 (.BL(BL122),.BLN(BLN122),.WL(WL60));
sram_cell_6t_5 inst_cell_60_123 (.BL(BL123),.BLN(BLN123),.WL(WL60));
sram_cell_6t_5 inst_cell_60_124 (.BL(BL124),.BLN(BLN124),.WL(WL60));
sram_cell_6t_5 inst_cell_60_125 (.BL(BL125),.BLN(BLN125),.WL(WL60));
sram_cell_6t_5 inst_cell_60_126 (.BL(BL126),.BLN(BLN126),.WL(WL60));
sram_cell_6t_5 inst_cell_60_127 (.BL(BL127),.BLN(BLN127),.WL(WL60));
sram_cell_6t_5 inst_cell_61_0 (.BL(BL0),.BLN(BLN0),.WL(WL61));
sram_cell_6t_5 inst_cell_61_1 (.BL(BL1),.BLN(BLN1),.WL(WL61));
sram_cell_6t_5 inst_cell_61_2 (.BL(BL2),.BLN(BLN2),.WL(WL61));
sram_cell_6t_5 inst_cell_61_3 (.BL(BL3),.BLN(BLN3),.WL(WL61));
sram_cell_6t_5 inst_cell_61_4 (.BL(BL4),.BLN(BLN4),.WL(WL61));
sram_cell_6t_5 inst_cell_61_5 (.BL(BL5),.BLN(BLN5),.WL(WL61));
sram_cell_6t_5 inst_cell_61_6 (.BL(BL6),.BLN(BLN6),.WL(WL61));
sram_cell_6t_5 inst_cell_61_7 (.BL(BL7),.BLN(BLN7),.WL(WL61));
sram_cell_6t_5 inst_cell_61_8 (.BL(BL8),.BLN(BLN8),.WL(WL61));
sram_cell_6t_5 inst_cell_61_9 (.BL(BL9),.BLN(BLN9),.WL(WL61));
sram_cell_6t_5 inst_cell_61_10 (.BL(BL10),.BLN(BLN10),.WL(WL61));
sram_cell_6t_5 inst_cell_61_11 (.BL(BL11),.BLN(BLN11),.WL(WL61));
sram_cell_6t_5 inst_cell_61_12 (.BL(BL12),.BLN(BLN12),.WL(WL61));
sram_cell_6t_5 inst_cell_61_13 (.BL(BL13),.BLN(BLN13),.WL(WL61));
sram_cell_6t_5 inst_cell_61_14 (.BL(BL14),.BLN(BLN14),.WL(WL61));
sram_cell_6t_5 inst_cell_61_15 (.BL(BL15),.BLN(BLN15),.WL(WL61));
sram_cell_6t_5 inst_cell_61_16 (.BL(BL16),.BLN(BLN16),.WL(WL61));
sram_cell_6t_5 inst_cell_61_17 (.BL(BL17),.BLN(BLN17),.WL(WL61));
sram_cell_6t_5 inst_cell_61_18 (.BL(BL18),.BLN(BLN18),.WL(WL61));
sram_cell_6t_5 inst_cell_61_19 (.BL(BL19),.BLN(BLN19),.WL(WL61));
sram_cell_6t_5 inst_cell_61_20 (.BL(BL20),.BLN(BLN20),.WL(WL61));
sram_cell_6t_5 inst_cell_61_21 (.BL(BL21),.BLN(BLN21),.WL(WL61));
sram_cell_6t_5 inst_cell_61_22 (.BL(BL22),.BLN(BLN22),.WL(WL61));
sram_cell_6t_5 inst_cell_61_23 (.BL(BL23),.BLN(BLN23),.WL(WL61));
sram_cell_6t_5 inst_cell_61_24 (.BL(BL24),.BLN(BLN24),.WL(WL61));
sram_cell_6t_5 inst_cell_61_25 (.BL(BL25),.BLN(BLN25),.WL(WL61));
sram_cell_6t_5 inst_cell_61_26 (.BL(BL26),.BLN(BLN26),.WL(WL61));
sram_cell_6t_5 inst_cell_61_27 (.BL(BL27),.BLN(BLN27),.WL(WL61));
sram_cell_6t_5 inst_cell_61_28 (.BL(BL28),.BLN(BLN28),.WL(WL61));
sram_cell_6t_5 inst_cell_61_29 (.BL(BL29),.BLN(BLN29),.WL(WL61));
sram_cell_6t_5 inst_cell_61_30 (.BL(BL30),.BLN(BLN30),.WL(WL61));
sram_cell_6t_5 inst_cell_61_31 (.BL(BL31),.BLN(BLN31),.WL(WL61));
sram_cell_6t_5 inst_cell_61_32 (.BL(BL32),.BLN(BLN32),.WL(WL61));
sram_cell_6t_5 inst_cell_61_33 (.BL(BL33),.BLN(BLN33),.WL(WL61));
sram_cell_6t_5 inst_cell_61_34 (.BL(BL34),.BLN(BLN34),.WL(WL61));
sram_cell_6t_5 inst_cell_61_35 (.BL(BL35),.BLN(BLN35),.WL(WL61));
sram_cell_6t_5 inst_cell_61_36 (.BL(BL36),.BLN(BLN36),.WL(WL61));
sram_cell_6t_5 inst_cell_61_37 (.BL(BL37),.BLN(BLN37),.WL(WL61));
sram_cell_6t_5 inst_cell_61_38 (.BL(BL38),.BLN(BLN38),.WL(WL61));
sram_cell_6t_5 inst_cell_61_39 (.BL(BL39),.BLN(BLN39),.WL(WL61));
sram_cell_6t_5 inst_cell_61_40 (.BL(BL40),.BLN(BLN40),.WL(WL61));
sram_cell_6t_5 inst_cell_61_41 (.BL(BL41),.BLN(BLN41),.WL(WL61));
sram_cell_6t_5 inst_cell_61_42 (.BL(BL42),.BLN(BLN42),.WL(WL61));
sram_cell_6t_5 inst_cell_61_43 (.BL(BL43),.BLN(BLN43),.WL(WL61));
sram_cell_6t_5 inst_cell_61_44 (.BL(BL44),.BLN(BLN44),.WL(WL61));
sram_cell_6t_5 inst_cell_61_45 (.BL(BL45),.BLN(BLN45),.WL(WL61));
sram_cell_6t_5 inst_cell_61_46 (.BL(BL46),.BLN(BLN46),.WL(WL61));
sram_cell_6t_5 inst_cell_61_47 (.BL(BL47),.BLN(BLN47),.WL(WL61));
sram_cell_6t_5 inst_cell_61_48 (.BL(BL48),.BLN(BLN48),.WL(WL61));
sram_cell_6t_5 inst_cell_61_49 (.BL(BL49),.BLN(BLN49),.WL(WL61));
sram_cell_6t_5 inst_cell_61_50 (.BL(BL50),.BLN(BLN50),.WL(WL61));
sram_cell_6t_5 inst_cell_61_51 (.BL(BL51),.BLN(BLN51),.WL(WL61));
sram_cell_6t_5 inst_cell_61_52 (.BL(BL52),.BLN(BLN52),.WL(WL61));
sram_cell_6t_5 inst_cell_61_53 (.BL(BL53),.BLN(BLN53),.WL(WL61));
sram_cell_6t_5 inst_cell_61_54 (.BL(BL54),.BLN(BLN54),.WL(WL61));
sram_cell_6t_5 inst_cell_61_55 (.BL(BL55),.BLN(BLN55),.WL(WL61));
sram_cell_6t_5 inst_cell_61_56 (.BL(BL56),.BLN(BLN56),.WL(WL61));
sram_cell_6t_5 inst_cell_61_57 (.BL(BL57),.BLN(BLN57),.WL(WL61));
sram_cell_6t_5 inst_cell_61_58 (.BL(BL58),.BLN(BLN58),.WL(WL61));
sram_cell_6t_5 inst_cell_61_59 (.BL(BL59),.BLN(BLN59),.WL(WL61));
sram_cell_6t_5 inst_cell_61_60 (.BL(BL60),.BLN(BLN60),.WL(WL61));
sram_cell_6t_5 inst_cell_61_61 (.BL(BL61),.BLN(BLN61),.WL(WL61));
sram_cell_6t_5 inst_cell_61_62 (.BL(BL62),.BLN(BLN62),.WL(WL61));
sram_cell_6t_5 inst_cell_61_63 (.BL(BL63),.BLN(BLN63),.WL(WL61));
sram_cell_6t_5 inst_cell_61_64 (.BL(BL64),.BLN(BLN64),.WL(WL61));
sram_cell_6t_5 inst_cell_61_65 (.BL(BL65),.BLN(BLN65),.WL(WL61));
sram_cell_6t_5 inst_cell_61_66 (.BL(BL66),.BLN(BLN66),.WL(WL61));
sram_cell_6t_5 inst_cell_61_67 (.BL(BL67),.BLN(BLN67),.WL(WL61));
sram_cell_6t_5 inst_cell_61_68 (.BL(BL68),.BLN(BLN68),.WL(WL61));
sram_cell_6t_5 inst_cell_61_69 (.BL(BL69),.BLN(BLN69),.WL(WL61));
sram_cell_6t_5 inst_cell_61_70 (.BL(BL70),.BLN(BLN70),.WL(WL61));
sram_cell_6t_5 inst_cell_61_71 (.BL(BL71),.BLN(BLN71),.WL(WL61));
sram_cell_6t_5 inst_cell_61_72 (.BL(BL72),.BLN(BLN72),.WL(WL61));
sram_cell_6t_5 inst_cell_61_73 (.BL(BL73),.BLN(BLN73),.WL(WL61));
sram_cell_6t_5 inst_cell_61_74 (.BL(BL74),.BLN(BLN74),.WL(WL61));
sram_cell_6t_5 inst_cell_61_75 (.BL(BL75),.BLN(BLN75),.WL(WL61));
sram_cell_6t_5 inst_cell_61_76 (.BL(BL76),.BLN(BLN76),.WL(WL61));
sram_cell_6t_5 inst_cell_61_77 (.BL(BL77),.BLN(BLN77),.WL(WL61));
sram_cell_6t_5 inst_cell_61_78 (.BL(BL78),.BLN(BLN78),.WL(WL61));
sram_cell_6t_5 inst_cell_61_79 (.BL(BL79),.BLN(BLN79),.WL(WL61));
sram_cell_6t_5 inst_cell_61_80 (.BL(BL80),.BLN(BLN80),.WL(WL61));
sram_cell_6t_5 inst_cell_61_81 (.BL(BL81),.BLN(BLN81),.WL(WL61));
sram_cell_6t_5 inst_cell_61_82 (.BL(BL82),.BLN(BLN82),.WL(WL61));
sram_cell_6t_5 inst_cell_61_83 (.BL(BL83),.BLN(BLN83),.WL(WL61));
sram_cell_6t_5 inst_cell_61_84 (.BL(BL84),.BLN(BLN84),.WL(WL61));
sram_cell_6t_5 inst_cell_61_85 (.BL(BL85),.BLN(BLN85),.WL(WL61));
sram_cell_6t_5 inst_cell_61_86 (.BL(BL86),.BLN(BLN86),.WL(WL61));
sram_cell_6t_5 inst_cell_61_87 (.BL(BL87),.BLN(BLN87),.WL(WL61));
sram_cell_6t_5 inst_cell_61_88 (.BL(BL88),.BLN(BLN88),.WL(WL61));
sram_cell_6t_5 inst_cell_61_89 (.BL(BL89),.BLN(BLN89),.WL(WL61));
sram_cell_6t_5 inst_cell_61_90 (.BL(BL90),.BLN(BLN90),.WL(WL61));
sram_cell_6t_5 inst_cell_61_91 (.BL(BL91),.BLN(BLN91),.WL(WL61));
sram_cell_6t_5 inst_cell_61_92 (.BL(BL92),.BLN(BLN92),.WL(WL61));
sram_cell_6t_5 inst_cell_61_93 (.BL(BL93),.BLN(BLN93),.WL(WL61));
sram_cell_6t_5 inst_cell_61_94 (.BL(BL94),.BLN(BLN94),.WL(WL61));
sram_cell_6t_5 inst_cell_61_95 (.BL(BL95),.BLN(BLN95),.WL(WL61));
sram_cell_6t_5 inst_cell_61_96 (.BL(BL96),.BLN(BLN96),.WL(WL61));
sram_cell_6t_5 inst_cell_61_97 (.BL(BL97),.BLN(BLN97),.WL(WL61));
sram_cell_6t_5 inst_cell_61_98 (.BL(BL98),.BLN(BLN98),.WL(WL61));
sram_cell_6t_5 inst_cell_61_99 (.BL(BL99),.BLN(BLN99),.WL(WL61));
sram_cell_6t_5 inst_cell_61_100 (.BL(BL100),.BLN(BLN100),.WL(WL61));
sram_cell_6t_5 inst_cell_61_101 (.BL(BL101),.BLN(BLN101),.WL(WL61));
sram_cell_6t_5 inst_cell_61_102 (.BL(BL102),.BLN(BLN102),.WL(WL61));
sram_cell_6t_5 inst_cell_61_103 (.BL(BL103),.BLN(BLN103),.WL(WL61));
sram_cell_6t_5 inst_cell_61_104 (.BL(BL104),.BLN(BLN104),.WL(WL61));
sram_cell_6t_5 inst_cell_61_105 (.BL(BL105),.BLN(BLN105),.WL(WL61));
sram_cell_6t_5 inst_cell_61_106 (.BL(BL106),.BLN(BLN106),.WL(WL61));
sram_cell_6t_5 inst_cell_61_107 (.BL(BL107),.BLN(BLN107),.WL(WL61));
sram_cell_6t_5 inst_cell_61_108 (.BL(BL108),.BLN(BLN108),.WL(WL61));
sram_cell_6t_5 inst_cell_61_109 (.BL(BL109),.BLN(BLN109),.WL(WL61));
sram_cell_6t_5 inst_cell_61_110 (.BL(BL110),.BLN(BLN110),.WL(WL61));
sram_cell_6t_5 inst_cell_61_111 (.BL(BL111),.BLN(BLN111),.WL(WL61));
sram_cell_6t_5 inst_cell_61_112 (.BL(BL112),.BLN(BLN112),.WL(WL61));
sram_cell_6t_5 inst_cell_61_113 (.BL(BL113),.BLN(BLN113),.WL(WL61));
sram_cell_6t_5 inst_cell_61_114 (.BL(BL114),.BLN(BLN114),.WL(WL61));
sram_cell_6t_5 inst_cell_61_115 (.BL(BL115),.BLN(BLN115),.WL(WL61));
sram_cell_6t_5 inst_cell_61_116 (.BL(BL116),.BLN(BLN116),.WL(WL61));
sram_cell_6t_5 inst_cell_61_117 (.BL(BL117),.BLN(BLN117),.WL(WL61));
sram_cell_6t_5 inst_cell_61_118 (.BL(BL118),.BLN(BLN118),.WL(WL61));
sram_cell_6t_5 inst_cell_61_119 (.BL(BL119),.BLN(BLN119),.WL(WL61));
sram_cell_6t_5 inst_cell_61_120 (.BL(BL120),.BLN(BLN120),.WL(WL61));
sram_cell_6t_5 inst_cell_61_121 (.BL(BL121),.BLN(BLN121),.WL(WL61));
sram_cell_6t_5 inst_cell_61_122 (.BL(BL122),.BLN(BLN122),.WL(WL61));
sram_cell_6t_5 inst_cell_61_123 (.BL(BL123),.BLN(BLN123),.WL(WL61));
sram_cell_6t_5 inst_cell_61_124 (.BL(BL124),.BLN(BLN124),.WL(WL61));
sram_cell_6t_5 inst_cell_61_125 (.BL(BL125),.BLN(BLN125),.WL(WL61));
sram_cell_6t_5 inst_cell_61_126 (.BL(BL126),.BLN(BLN126),.WL(WL61));
sram_cell_6t_5 inst_cell_61_127 (.BL(BL127),.BLN(BLN127),.WL(WL61));
sram_cell_6t_5 inst_cell_62_0 (.BL(BL0),.BLN(BLN0),.WL(WL62));
sram_cell_6t_5 inst_cell_62_1 (.BL(BL1),.BLN(BLN1),.WL(WL62));
sram_cell_6t_5 inst_cell_62_2 (.BL(BL2),.BLN(BLN2),.WL(WL62));
sram_cell_6t_5 inst_cell_62_3 (.BL(BL3),.BLN(BLN3),.WL(WL62));
sram_cell_6t_5 inst_cell_62_4 (.BL(BL4),.BLN(BLN4),.WL(WL62));
sram_cell_6t_5 inst_cell_62_5 (.BL(BL5),.BLN(BLN5),.WL(WL62));
sram_cell_6t_5 inst_cell_62_6 (.BL(BL6),.BLN(BLN6),.WL(WL62));
sram_cell_6t_5 inst_cell_62_7 (.BL(BL7),.BLN(BLN7),.WL(WL62));
sram_cell_6t_5 inst_cell_62_8 (.BL(BL8),.BLN(BLN8),.WL(WL62));
sram_cell_6t_5 inst_cell_62_9 (.BL(BL9),.BLN(BLN9),.WL(WL62));
sram_cell_6t_5 inst_cell_62_10 (.BL(BL10),.BLN(BLN10),.WL(WL62));
sram_cell_6t_5 inst_cell_62_11 (.BL(BL11),.BLN(BLN11),.WL(WL62));
sram_cell_6t_5 inst_cell_62_12 (.BL(BL12),.BLN(BLN12),.WL(WL62));
sram_cell_6t_5 inst_cell_62_13 (.BL(BL13),.BLN(BLN13),.WL(WL62));
sram_cell_6t_5 inst_cell_62_14 (.BL(BL14),.BLN(BLN14),.WL(WL62));
sram_cell_6t_5 inst_cell_62_15 (.BL(BL15),.BLN(BLN15),.WL(WL62));
sram_cell_6t_5 inst_cell_62_16 (.BL(BL16),.BLN(BLN16),.WL(WL62));
sram_cell_6t_5 inst_cell_62_17 (.BL(BL17),.BLN(BLN17),.WL(WL62));
sram_cell_6t_5 inst_cell_62_18 (.BL(BL18),.BLN(BLN18),.WL(WL62));
sram_cell_6t_5 inst_cell_62_19 (.BL(BL19),.BLN(BLN19),.WL(WL62));
sram_cell_6t_5 inst_cell_62_20 (.BL(BL20),.BLN(BLN20),.WL(WL62));
sram_cell_6t_5 inst_cell_62_21 (.BL(BL21),.BLN(BLN21),.WL(WL62));
sram_cell_6t_5 inst_cell_62_22 (.BL(BL22),.BLN(BLN22),.WL(WL62));
sram_cell_6t_5 inst_cell_62_23 (.BL(BL23),.BLN(BLN23),.WL(WL62));
sram_cell_6t_5 inst_cell_62_24 (.BL(BL24),.BLN(BLN24),.WL(WL62));
sram_cell_6t_5 inst_cell_62_25 (.BL(BL25),.BLN(BLN25),.WL(WL62));
sram_cell_6t_5 inst_cell_62_26 (.BL(BL26),.BLN(BLN26),.WL(WL62));
sram_cell_6t_5 inst_cell_62_27 (.BL(BL27),.BLN(BLN27),.WL(WL62));
sram_cell_6t_5 inst_cell_62_28 (.BL(BL28),.BLN(BLN28),.WL(WL62));
sram_cell_6t_5 inst_cell_62_29 (.BL(BL29),.BLN(BLN29),.WL(WL62));
sram_cell_6t_5 inst_cell_62_30 (.BL(BL30),.BLN(BLN30),.WL(WL62));
sram_cell_6t_5 inst_cell_62_31 (.BL(BL31),.BLN(BLN31),.WL(WL62));
sram_cell_6t_5 inst_cell_62_32 (.BL(BL32),.BLN(BLN32),.WL(WL62));
sram_cell_6t_5 inst_cell_62_33 (.BL(BL33),.BLN(BLN33),.WL(WL62));
sram_cell_6t_5 inst_cell_62_34 (.BL(BL34),.BLN(BLN34),.WL(WL62));
sram_cell_6t_5 inst_cell_62_35 (.BL(BL35),.BLN(BLN35),.WL(WL62));
sram_cell_6t_5 inst_cell_62_36 (.BL(BL36),.BLN(BLN36),.WL(WL62));
sram_cell_6t_5 inst_cell_62_37 (.BL(BL37),.BLN(BLN37),.WL(WL62));
sram_cell_6t_5 inst_cell_62_38 (.BL(BL38),.BLN(BLN38),.WL(WL62));
sram_cell_6t_5 inst_cell_62_39 (.BL(BL39),.BLN(BLN39),.WL(WL62));
sram_cell_6t_5 inst_cell_62_40 (.BL(BL40),.BLN(BLN40),.WL(WL62));
sram_cell_6t_5 inst_cell_62_41 (.BL(BL41),.BLN(BLN41),.WL(WL62));
sram_cell_6t_5 inst_cell_62_42 (.BL(BL42),.BLN(BLN42),.WL(WL62));
sram_cell_6t_5 inst_cell_62_43 (.BL(BL43),.BLN(BLN43),.WL(WL62));
sram_cell_6t_5 inst_cell_62_44 (.BL(BL44),.BLN(BLN44),.WL(WL62));
sram_cell_6t_5 inst_cell_62_45 (.BL(BL45),.BLN(BLN45),.WL(WL62));
sram_cell_6t_5 inst_cell_62_46 (.BL(BL46),.BLN(BLN46),.WL(WL62));
sram_cell_6t_5 inst_cell_62_47 (.BL(BL47),.BLN(BLN47),.WL(WL62));
sram_cell_6t_5 inst_cell_62_48 (.BL(BL48),.BLN(BLN48),.WL(WL62));
sram_cell_6t_5 inst_cell_62_49 (.BL(BL49),.BLN(BLN49),.WL(WL62));
sram_cell_6t_5 inst_cell_62_50 (.BL(BL50),.BLN(BLN50),.WL(WL62));
sram_cell_6t_5 inst_cell_62_51 (.BL(BL51),.BLN(BLN51),.WL(WL62));
sram_cell_6t_5 inst_cell_62_52 (.BL(BL52),.BLN(BLN52),.WL(WL62));
sram_cell_6t_5 inst_cell_62_53 (.BL(BL53),.BLN(BLN53),.WL(WL62));
sram_cell_6t_5 inst_cell_62_54 (.BL(BL54),.BLN(BLN54),.WL(WL62));
sram_cell_6t_5 inst_cell_62_55 (.BL(BL55),.BLN(BLN55),.WL(WL62));
sram_cell_6t_5 inst_cell_62_56 (.BL(BL56),.BLN(BLN56),.WL(WL62));
sram_cell_6t_5 inst_cell_62_57 (.BL(BL57),.BLN(BLN57),.WL(WL62));
sram_cell_6t_5 inst_cell_62_58 (.BL(BL58),.BLN(BLN58),.WL(WL62));
sram_cell_6t_5 inst_cell_62_59 (.BL(BL59),.BLN(BLN59),.WL(WL62));
sram_cell_6t_5 inst_cell_62_60 (.BL(BL60),.BLN(BLN60),.WL(WL62));
sram_cell_6t_5 inst_cell_62_61 (.BL(BL61),.BLN(BLN61),.WL(WL62));
sram_cell_6t_5 inst_cell_62_62 (.BL(BL62),.BLN(BLN62),.WL(WL62));
sram_cell_6t_5 inst_cell_62_63 (.BL(BL63),.BLN(BLN63),.WL(WL62));
sram_cell_6t_5 inst_cell_62_64 (.BL(BL64),.BLN(BLN64),.WL(WL62));
sram_cell_6t_5 inst_cell_62_65 (.BL(BL65),.BLN(BLN65),.WL(WL62));
sram_cell_6t_5 inst_cell_62_66 (.BL(BL66),.BLN(BLN66),.WL(WL62));
sram_cell_6t_5 inst_cell_62_67 (.BL(BL67),.BLN(BLN67),.WL(WL62));
sram_cell_6t_5 inst_cell_62_68 (.BL(BL68),.BLN(BLN68),.WL(WL62));
sram_cell_6t_5 inst_cell_62_69 (.BL(BL69),.BLN(BLN69),.WL(WL62));
sram_cell_6t_5 inst_cell_62_70 (.BL(BL70),.BLN(BLN70),.WL(WL62));
sram_cell_6t_5 inst_cell_62_71 (.BL(BL71),.BLN(BLN71),.WL(WL62));
sram_cell_6t_5 inst_cell_62_72 (.BL(BL72),.BLN(BLN72),.WL(WL62));
sram_cell_6t_5 inst_cell_62_73 (.BL(BL73),.BLN(BLN73),.WL(WL62));
sram_cell_6t_5 inst_cell_62_74 (.BL(BL74),.BLN(BLN74),.WL(WL62));
sram_cell_6t_5 inst_cell_62_75 (.BL(BL75),.BLN(BLN75),.WL(WL62));
sram_cell_6t_5 inst_cell_62_76 (.BL(BL76),.BLN(BLN76),.WL(WL62));
sram_cell_6t_5 inst_cell_62_77 (.BL(BL77),.BLN(BLN77),.WL(WL62));
sram_cell_6t_5 inst_cell_62_78 (.BL(BL78),.BLN(BLN78),.WL(WL62));
sram_cell_6t_5 inst_cell_62_79 (.BL(BL79),.BLN(BLN79),.WL(WL62));
sram_cell_6t_5 inst_cell_62_80 (.BL(BL80),.BLN(BLN80),.WL(WL62));
sram_cell_6t_5 inst_cell_62_81 (.BL(BL81),.BLN(BLN81),.WL(WL62));
sram_cell_6t_5 inst_cell_62_82 (.BL(BL82),.BLN(BLN82),.WL(WL62));
sram_cell_6t_5 inst_cell_62_83 (.BL(BL83),.BLN(BLN83),.WL(WL62));
sram_cell_6t_5 inst_cell_62_84 (.BL(BL84),.BLN(BLN84),.WL(WL62));
sram_cell_6t_5 inst_cell_62_85 (.BL(BL85),.BLN(BLN85),.WL(WL62));
sram_cell_6t_5 inst_cell_62_86 (.BL(BL86),.BLN(BLN86),.WL(WL62));
sram_cell_6t_5 inst_cell_62_87 (.BL(BL87),.BLN(BLN87),.WL(WL62));
sram_cell_6t_5 inst_cell_62_88 (.BL(BL88),.BLN(BLN88),.WL(WL62));
sram_cell_6t_5 inst_cell_62_89 (.BL(BL89),.BLN(BLN89),.WL(WL62));
sram_cell_6t_5 inst_cell_62_90 (.BL(BL90),.BLN(BLN90),.WL(WL62));
sram_cell_6t_5 inst_cell_62_91 (.BL(BL91),.BLN(BLN91),.WL(WL62));
sram_cell_6t_5 inst_cell_62_92 (.BL(BL92),.BLN(BLN92),.WL(WL62));
sram_cell_6t_5 inst_cell_62_93 (.BL(BL93),.BLN(BLN93),.WL(WL62));
sram_cell_6t_5 inst_cell_62_94 (.BL(BL94),.BLN(BLN94),.WL(WL62));
sram_cell_6t_5 inst_cell_62_95 (.BL(BL95),.BLN(BLN95),.WL(WL62));
sram_cell_6t_5 inst_cell_62_96 (.BL(BL96),.BLN(BLN96),.WL(WL62));
sram_cell_6t_5 inst_cell_62_97 (.BL(BL97),.BLN(BLN97),.WL(WL62));
sram_cell_6t_5 inst_cell_62_98 (.BL(BL98),.BLN(BLN98),.WL(WL62));
sram_cell_6t_5 inst_cell_62_99 (.BL(BL99),.BLN(BLN99),.WL(WL62));
sram_cell_6t_5 inst_cell_62_100 (.BL(BL100),.BLN(BLN100),.WL(WL62));
sram_cell_6t_5 inst_cell_62_101 (.BL(BL101),.BLN(BLN101),.WL(WL62));
sram_cell_6t_5 inst_cell_62_102 (.BL(BL102),.BLN(BLN102),.WL(WL62));
sram_cell_6t_5 inst_cell_62_103 (.BL(BL103),.BLN(BLN103),.WL(WL62));
sram_cell_6t_5 inst_cell_62_104 (.BL(BL104),.BLN(BLN104),.WL(WL62));
sram_cell_6t_5 inst_cell_62_105 (.BL(BL105),.BLN(BLN105),.WL(WL62));
sram_cell_6t_5 inst_cell_62_106 (.BL(BL106),.BLN(BLN106),.WL(WL62));
sram_cell_6t_5 inst_cell_62_107 (.BL(BL107),.BLN(BLN107),.WL(WL62));
sram_cell_6t_5 inst_cell_62_108 (.BL(BL108),.BLN(BLN108),.WL(WL62));
sram_cell_6t_5 inst_cell_62_109 (.BL(BL109),.BLN(BLN109),.WL(WL62));
sram_cell_6t_5 inst_cell_62_110 (.BL(BL110),.BLN(BLN110),.WL(WL62));
sram_cell_6t_5 inst_cell_62_111 (.BL(BL111),.BLN(BLN111),.WL(WL62));
sram_cell_6t_5 inst_cell_62_112 (.BL(BL112),.BLN(BLN112),.WL(WL62));
sram_cell_6t_5 inst_cell_62_113 (.BL(BL113),.BLN(BLN113),.WL(WL62));
sram_cell_6t_5 inst_cell_62_114 (.BL(BL114),.BLN(BLN114),.WL(WL62));
sram_cell_6t_5 inst_cell_62_115 (.BL(BL115),.BLN(BLN115),.WL(WL62));
sram_cell_6t_5 inst_cell_62_116 (.BL(BL116),.BLN(BLN116),.WL(WL62));
sram_cell_6t_5 inst_cell_62_117 (.BL(BL117),.BLN(BLN117),.WL(WL62));
sram_cell_6t_5 inst_cell_62_118 (.BL(BL118),.BLN(BLN118),.WL(WL62));
sram_cell_6t_5 inst_cell_62_119 (.BL(BL119),.BLN(BLN119),.WL(WL62));
sram_cell_6t_5 inst_cell_62_120 (.BL(BL120),.BLN(BLN120),.WL(WL62));
sram_cell_6t_5 inst_cell_62_121 (.BL(BL121),.BLN(BLN121),.WL(WL62));
sram_cell_6t_5 inst_cell_62_122 (.BL(BL122),.BLN(BLN122),.WL(WL62));
sram_cell_6t_5 inst_cell_62_123 (.BL(BL123),.BLN(BLN123),.WL(WL62));
sram_cell_6t_5 inst_cell_62_124 (.BL(BL124),.BLN(BLN124),.WL(WL62));
sram_cell_6t_5 inst_cell_62_125 (.BL(BL125),.BLN(BLN125),.WL(WL62));
sram_cell_6t_5 inst_cell_62_126 (.BL(BL126),.BLN(BLN126),.WL(WL62));
sram_cell_6t_5 inst_cell_62_127 (.BL(BL127),.BLN(BLN127),.WL(WL62));
sram_cell_6t_5 inst_cell_63_0 (.BL(BL0),.BLN(BLN0),.WL(WL63));
sram_cell_6t_5 inst_cell_63_1 (.BL(BL1),.BLN(BLN1),.WL(WL63));
sram_cell_6t_5 inst_cell_63_2 (.BL(BL2),.BLN(BLN2),.WL(WL63));
sram_cell_6t_5 inst_cell_63_3 (.BL(BL3),.BLN(BLN3),.WL(WL63));
sram_cell_6t_5 inst_cell_63_4 (.BL(BL4),.BLN(BLN4),.WL(WL63));
sram_cell_6t_5 inst_cell_63_5 (.BL(BL5),.BLN(BLN5),.WL(WL63));
sram_cell_6t_5 inst_cell_63_6 (.BL(BL6),.BLN(BLN6),.WL(WL63));
sram_cell_6t_5 inst_cell_63_7 (.BL(BL7),.BLN(BLN7),.WL(WL63));
sram_cell_6t_5 inst_cell_63_8 (.BL(BL8),.BLN(BLN8),.WL(WL63));
sram_cell_6t_5 inst_cell_63_9 (.BL(BL9),.BLN(BLN9),.WL(WL63));
sram_cell_6t_5 inst_cell_63_10 (.BL(BL10),.BLN(BLN10),.WL(WL63));
sram_cell_6t_5 inst_cell_63_11 (.BL(BL11),.BLN(BLN11),.WL(WL63));
sram_cell_6t_5 inst_cell_63_12 (.BL(BL12),.BLN(BLN12),.WL(WL63));
sram_cell_6t_5 inst_cell_63_13 (.BL(BL13),.BLN(BLN13),.WL(WL63));
sram_cell_6t_5 inst_cell_63_14 (.BL(BL14),.BLN(BLN14),.WL(WL63));
sram_cell_6t_5 inst_cell_63_15 (.BL(BL15),.BLN(BLN15),.WL(WL63));
sram_cell_6t_5 inst_cell_63_16 (.BL(BL16),.BLN(BLN16),.WL(WL63));
sram_cell_6t_5 inst_cell_63_17 (.BL(BL17),.BLN(BLN17),.WL(WL63));
sram_cell_6t_5 inst_cell_63_18 (.BL(BL18),.BLN(BLN18),.WL(WL63));
sram_cell_6t_5 inst_cell_63_19 (.BL(BL19),.BLN(BLN19),.WL(WL63));
sram_cell_6t_5 inst_cell_63_20 (.BL(BL20),.BLN(BLN20),.WL(WL63));
sram_cell_6t_5 inst_cell_63_21 (.BL(BL21),.BLN(BLN21),.WL(WL63));
sram_cell_6t_5 inst_cell_63_22 (.BL(BL22),.BLN(BLN22),.WL(WL63));
sram_cell_6t_5 inst_cell_63_23 (.BL(BL23),.BLN(BLN23),.WL(WL63));
sram_cell_6t_5 inst_cell_63_24 (.BL(BL24),.BLN(BLN24),.WL(WL63));
sram_cell_6t_5 inst_cell_63_25 (.BL(BL25),.BLN(BLN25),.WL(WL63));
sram_cell_6t_5 inst_cell_63_26 (.BL(BL26),.BLN(BLN26),.WL(WL63));
sram_cell_6t_5 inst_cell_63_27 (.BL(BL27),.BLN(BLN27),.WL(WL63));
sram_cell_6t_5 inst_cell_63_28 (.BL(BL28),.BLN(BLN28),.WL(WL63));
sram_cell_6t_5 inst_cell_63_29 (.BL(BL29),.BLN(BLN29),.WL(WL63));
sram_cell_6t_5 inst_cell_63_30 (.BL(BL30),.BLN(BLN30),.WL(WL63));
sram_cell_6t_5 inst_cell_63_31 (.BL(BL31),.BLN(BLN31),.WL(WL63));
sram_cell_6t_5 inst_cell_63_32 (.BL(BL32),.BLN(BLN32),.WL(WL63));
sram_cell_6t_5 inst_cell_63_33 (.BL(BL33),.BLN(BLN33),.WL(WL63));
sram_cell_6t_5 inst_cell_63_34 (.BL(BL34),.BLN(BLN34),.WL(WL63));
sram_cell_6t_5 inst_cell_63_35 (.BL(BL35),.BLN(BLN35),.WL(WL63));
sram_cell_6t_5 inst_cell_63_36 (.BL(BL36),.BLN(BLN36),.WL(WL63));
sram_cell_6t_5 inst_cell_63_37 (.BL(BL37),.BLN(BLN37),.WL(WL63));
sram_cell_6t_5 inst_cell_63_38 (.BL(BL38),.BLN(BLN38),.WL(WL63));
sram_cell_6t_5 inst_cell_63_39 (.BL(BL39),.BLN(BLN39),.WL(WL63));
sram_cell_6t_5 inst_cell_63_40 (.BL(BL40),.BLN(BLN40),.WL(WL63));
sram_cell_6t_5 inst_cell_63_41 (.BL(BL41),.BLN(BLN41),.WL(WL63));
sram_cell_6t_5 inst_cell_63_42 (.BL(BL42),.BLN(BLN42),.WL(WL63));
sram_cell_6t_5 inst_cell_63_43 (.BL(BL43),.BLN(BLN43),.WL(WL63));
sram_cell_6t_5 inst_cell_63_44 (.BL(BL44),.BLN(BLN44),.WL(WL63));
sram_cell_6t_5 inst_cell_63_45 (.BL(BL45),.BLN(BLN45),.WL(WL63));
sram_cell_6t_5 inst_cell_63_46 (.BL(BL46),.BLN(BLN46),.WL(WL63));
sram_cell_6t_5 inst_cell_63_47 (.BL(BL47),.BLN(BLN47),.WL(WL63));
sram_cell_6t_5 inst_cell_63_48 (.BL(BL48),.BLN(BLN48),.WL(WL63));
sram_cell_6t_5 inst_cell_63_49 (.BL(BL49),.BLN(BLN49),.WL(WL63));
sram_cell_6t_5 inst_cell_63_50 (.BL(BL50),.BLN(BLN50),.WL(WL63));
sram_cell_6t_5 inst_cell_63_51 (.BL(BL51),.BLN(BLN51),.WL(WL63));
sram_cell_6t_5 inst_cell_63_52 (.BL(BL52),.BLN(BLN52),.WL(WL63));
sram_cell_6t_5 inst_cell_63_53 (.BL(BL53),.BLN(BLN53),.WL(WL63));
sram_cell_6t_5 inst_cell_63_54 (.BL(BL54),.BLN(BLN54),.WL(WL63));
sram_cell_6t_5 inst_cell_63_55 (.BL(BL55),.BLN(BLN55),.WL(WL63));
sram_cell_6t_5 inst_cell_63_56 (.BL(BL56),.BLN(BLN56),.WL(WL63));
sram_cell_6t_5 inst_cell_63_57 (.BL(BL57),.BLN(BLN57),.WL(WL63));
sram_cell_6t_5 inst_cell_63_58 (.BL(BL58),.BLN(BLN58),.WL(WL63));
sram_cell_6t_5 inst_cell_63_59 (.BL(BL59),.BLN(BLN59),.WL(WL63));
sram_cell_6t_5 inst_cell_63_60 (.BL(BL60),.BLN(BLN60),.WL(WL63));
sram_cell_6t_5 inst_cell_63_61 (.BL(BL61),.BLN(BLN61),.WL(WL63));
sram_cell_6t_5 inst_cell_63_62 (.BL(BL62),.BLN(BLN62),.WL(WL63));
sram_cell_6t_5 inst_cell_63_63 (.BL(BL63),.BLN(BLN63),.WL(WL63));
sram_cell_6t_5 inst_cell_63_64 (.BL(BL64),.BLN(BLN64),.WL(WL63));
sram_cell_6t_5 inst_cell_63_65 (.BL(BL65),.BLN(BLN65),.WL(WL63));
sram_cell_6t_5 inst_cell_63_66 (.BL(BL66),.BLN(BLN66),.WL(WL63));
sram_cell_6t_5 inst_cell_63_67 (.BL(BL67),.BLN(BLN67),.WL(WL63));
sram_cell_6t_5 inst_cell_63_68 (.BL(BL68),.BLN(BLN68),.WL(WL63));
sram_cell_6t_5 inst_cell_63_69 (.BL(BL69),.BLN(BLN69),.WL(WL63));
sram_cell_6t_5 inst_cell_63_70 (.BL(BL70),.BLN(BLN70),.WL(WL63));
sram_cell_6t_5 inst_cell_63_71 (.BL(BL71),.BLN(BLN71),.WL(WL63));
sram_cell_6t_5 inst_cell_63_72 (.BL(BL72),.BLN(BLN72),.WL(WL63));
sram_cell_6t_5 inst_cell_63_73 (.BL(BL73),.BLN(BLN73),.WL(WL63));
sram_cell_6t_5 inst_cell_63_74 (.BL(BL74),.BLN(BLN74),.WL(WL63));
sram_cell_6t_5 inst_cell_63_75 (.BL(BL75),.BLN(BLN75),.WL(WL63));
sram_cell_6t_5 inst_cell_63_76 (.BL(BL76),.BLN(BLN76),.WL(WL63));
sram_cell_6t_5 inst_cell_63_77 (.BL(BL77),.BLN(BLN77),.WL(WL63));
sram_cell_6t_5 inst_cell_63_78 (.BL(BL78),.BLN(BLN78),.WL(WL63));
sram_cell_6t_5 inst_cell_63_79 (.BL(BL79),.BLN(BLN79),.WL(WL63));
sram_cell_6t_5 inst_cell_63_80 (.BL(BL80),.BLN(BLN80),.WL(WL63));
sram_cell_6t_5 inst_cell_63_81 (.BL(BL81),.BLN(BLN81),.WL(WL63));
sram_cell_6t_5 inst_cell_63_82 (.BL(BL82),.BLN(BLN82),.WL(WL63));
sram_cell_6t_5 inst_cell_63_83 (.BL(BL83),.BLN(BLN83),.WL(WL63));
sram_cell_6t_5 inst_cell_63_84 (.BL(BL84),.BLN(BLN84),.WL(WL63));
sram_cell_6t_5 inst_cell_63_85 (.BL(BL85),.BLN(BLN85),.WL(WL63));
sram_cell_6t_5 inst_cell_63_86 (.BL(BL86),.BLN(BLN86),.WL(WL63));
sram_cell_6t_5 inst_cell_63_87 (.BL(BL87),.BLN(BLN87),.WL(WL63));
sram_cell_6t_5 inst_cell_63_88 (.BL(BL88),.BLN(BLN88),.WL(WL63));
sram_cell_6t_5 inst_cell_63_89 (.BL(BL89),.BLN(BLN89),.WL(WL63));
sram_cell_6t_5 inst_cell_63_90 (.BL(BL90),.BLN(BLN90),.WL(WL63));
sram_cell_6t_5 inst_cell_63_91 (.BL(BL91),.BLN(BLN91),.WL(WL63));
sram_cell_6t_5 inst_cell_63_92 (.BL(BL92),.BLN(BLN92),.WL(WL63));
sram_cell_6t_5 inst_cell_63_93 (.BL(BL93),.BLN(BLN93),.WL(WL63));
sram_cell_6t_5 inst_cell_63_94 (.BL(BL94),.BLN(BLN94),.WL(WL63));
sram_cell_6t_5 inst_cell_63_95 (.BL(BL95),.BLN(BLN95),.WL(WL63));
sram_cell_6t_5 inst_cell_63_96 (.BL(BL96),.BLN(BLN96),.WL(WL63));
sram_cell_6t_5 inst_cell_63_97 (.BL(BL97),.BLN(BLN97),.WL(WL63));
sram_cell_6t_5 inst_cell_63_98 (.BL(BL98),.BLN(BLN98),.WL(WL63));
sram_cell_6t_5 inst_cell_63_99 (.BL(BL99),.BLN(BLN99),.WL(WL63));
sram_cell_6t_5 inst_cell_63_100 (.BL(BL100),.BLN(BLN100),.WL(WL63));
sram_cell_6t_5 inst_cell_63_101 (.BL(BL101),.BLN(BLN101),.WL(WL63));
sram_cell_6t_5 inst_cell_63_102 (.BL(BL102),.BLN(BLN102),.WL(WL63));
sram_cell_6t_5 inst_cell_63_103 (.BL(BL103),.BLN(BLN103),.WL(WL63));
sram_cell_6t_5 inst_cell_63_104 (.BL(BL104),.BLN(BLN104),.WL(WL63));
sram_cell_6t_5 inst_cell_63_105 (.BL(BL105),.BLN(BLN105),.WL(WL63));
sram_cell_6t_5 inst_cell_63_106 (.BL(BL106),.BLN(BLN106),.WL(WL63));
sram_cell_6t_5 inst_cell_63_107 (.BL(BL107),.BLN(BLN107),.WL(WL63));
sram_cell_6t_5 inst_cell_63_108 (.BL(BL108),.BLN(BLN108),.WL(WL63));
sram_cell_6t_5 inst_cell_63_109 (.BL(BL109),.BLN(BLN109),.WL(WL63));
sram_cell_6t_5 inst_cell_63_110 (.BL(BL110),.BLN(BLN110),.WL(WL63));
sram_cell_6t_5 inst_cell_63_111 (.BL(BL111),.BLN(BLN111),.WL(WL63));
sram_cell_6t_5 inst_cell_63_112 (.BL(BL112),.BLN(BLN112),.WL(WL63));
sram_cell_6t_5 inst_cell_63_113 (.BL(BL113),.BLN(BLN113),.WL(WL63));
sram_cell_6t_5 inst_cell_63_114 (.BL(BL114),.BLN(BLN114),.WL(WL63));
sram_cell_6t_5 inst_cell_63_115 (.BL(BL115),.BLN(BLN115),.WL(WL63));
sram_cell_6t_5 inst_cell_63_116 (.BL(BL116),.BLN(BLN116),.WL(WL63));
sram_cell_6t_5 inst_cell_63_117 (.BL(BL117),.BLN(BLN117),.WL(WL63));
sram_cell_6t_5 inst_cell_63_118 (.BL(BL118),.BLN(BLN118),.WL(WL63));
sram_cell_6t_5 inst_cell_63_119 (.BL(BL119),.BLN(BLN119),.WL(WL63));
sram_cell_6t_5 inst_cell_63_120 (.BL(BL120),.BLN(BLN120),.WL(WL63));
sram_cell_6t_5 inst_cell_63_121 (.BL(BL121),.BLN(BLN121),.WL(WL63));
sram_cell_6t_5 inst_cell_63_122 (.BL(BL122),.BLN(BLN122),.WL(WL63));
sram_cell_6t_5 inst_cell_63_123 (.BL(BL123),.BLN(BLN123),.WL(WL63));
sram_cell_6t_5 inst_cell_63_124 (.BL(BL124),.BLN(BLN124),.WL(WL63));
sram_cell_6t_5 inst_cell_63_125 (.BL(BL125),.BLN(BLN125),.WL(WL63));
sram_cell_6t_5 inst_cell_63_126 (.BL(BL126),.BLN(BLN126),.WL(WL63));
sram_cell_6t_5 inst_cell_63_127 (.BL(BL127),.BLN(BLN127),.WL(WL63));
sram_cell_6t_5 inst_cell_64_0 (.BL(BL0),.BLN(BLN0),.WL(WL64));
sram_cell_6t_5 inst_cell_64_1 (.BL(BL1),.BLN(BLN1),.WL(WL64));
sram_cell_6t_5 inst_cell_64_2 (.BL(BL2),.BLN(BLN2),.WL(WL64));
sram_cell_6t_5 inst_cell_64_3 (.BL(BL3),.BLN(BLN3),.WL(WL64));
sram_cell_6t_5 inst_cell_64_4 (.BL(BL4),.BLN(BLN4),.WL(WL64));
sram_cell_6t_5 inst_cell_64_5 (.BL(BL5),.BLN(BLN5),.WL(WL64));
sram_cell_6t_5 inst_cell_64_6 (.BL(BL6),.BLN(BLN6),.WL(WL64));
sram_cell_6t_5 inst_cell_64_7 (.BL(BL7),.BLN(BLN7),.WL(WL64));
sram_cell_6t_5 inst_cell_64_8 (.BL(BL8),.BLN(BLN8),.WL(WL64));
sram_cell_6t_5 inst_cell_64_9 (.BL(BL9),.BLN(BLN9),.WL(WL64));
sram_cell_6t_5 inst_cell_64_10 (.BL(BL10),.BLN(BLN10),.WL(WL64));
sram_cell_6t_5 inst_cell_64_11 (.BL(BL11),.BLN(BLN11),.WL(WL64));
sram_cell_6t_5 inst_cell_64_12 (.BL(BL12),.BLN(BLN12),.WL(WL64));
sram_cell_6t_5 inst_cell_64_13 (.BL(BL13),.BLN(BLN13),.WL(WL64));
sram_cell_6t_5 inst_cell_64_14 (.BL(BL14),.BLN(BLN14),.WL(WL64));
sram_cell_6t_5 inst_cell_64_15 (.BL(BL15),.BLN(BLN15),.WL(WL64));
sram_cell_6t_5 inst_cell_64_16 (.BL(BL16),.BLN(BLN16),.WL(WL64));
sram_cell_6t_5 inst_cell_64_17 (.BL(BL17),.BLN(BLN17),.WL(WL64));
sram_cell_6t_5 inst_cell_64_18 (.BL(BL18),.BLN(BLN18),.WL(WL64));
sram_cell_6t_5 inst_cell_64_19 (.BL(BL19),.BLN(BLN19),.WL(WL64));
sram_cell_6t_5 inst_cell_64_20 (.BL(BL20),.BLN(BLN20),.WL(WL64));
sram_cell_6t_5 inst_cell_64_21 (.BL(BL21),.BLN(BLN21),.WL(WL64));
sram_cell_6t_5 inst_cell_64_22 (.BL(BL22),.BLN(BLN22),.WL(WL64));
sram_cell_6t_5 inst_cell_64_23 (.BL(BL23),.BLN(BLN23),.WL(WL64));
sram_cell_6t_5 inst_cell_64_24 (.BL(BL24),.BLN(BLN24),.WL(WL64));
sram_cell_6t_5 inst_cell_64_25 (.BL(BL25),.BLN(BLN25),.WL(WL64));
sram_cell_6t_5 inst_cell_64_26 (.BL(BL26),.BLN(BLN26),.WL(WL64));
sram_cell_6t_5 inst_cell_64_27 (.BL(BL27),.BLN(BLN27),.WL(WL64));
sram_cell_6t_5 inst_cell_64_28 (.BL(BL28),.BLN(BLN28),.WL(WL64));
sram_cell_6t_5 inst_cell_64_29 (.BL(BL29),.BLN(BLN29),.WL(WL64));
sram_cell_6t_5 inst_cell_64_30 (.BL(BL30),.BLN(BLN30),.WL(WL64));
sram_cell_6t_5 inst_cell_64_31 (.BL(BL31),.BLN(BLN31),.WL(WL64));
sram_cell_6t_5 inst_cell_64_32 (.BL(BL32),.BLN(BLN32),.WL(WL64));
sram_cell_6t_5 inst_cell_64_33 (.BL(BL33),.BLN(BLN33),.WL(WL64));
sram_cell_6t_5 inst_cell_64_34 (.BL(BL34),.BLN(BLN34),.WL(WL64));
sram_cell_6t_5 inst_cell_64_35 (.BL(BL35),.BLN(BLN35),.WL(WL64));
sram_cell_6t_5 inst_cell_64_36 (.BL(BL36),.BLN(BLN36),.WL(WL64));
sram_cell_6t_5 inst_cell_64_37 (.BL(BL37),.BLN(BLN37),.WL(WL64));
sram_cell_6t_5 inst_cell_64_38 (.BL(BL38),.BLN(BLN38),.WL(WL64));
sram_cell_6t_5 inst_cell_64_39 (.BL(BL39),.BLN(BLN39),.WL(WL64));
sram_cell_6t_5 inst_cell_64_40 (.BL(BL40),.BLN(BLN40),.WL(WL64));
sram_cell_6t_5 inst_cell_64_41 (.BL(BL41),.BLN(BLN41),.WL(WL64));
sram_cell_6t_5 inst_cell_64_42 (.BL(BL42),.BLN(BLN42),.WL(WL64));
sram_cell_6t_5 inst_cell_64_43 (.BL(BL43),.BLN(BLN43),.WL(WL64));
sram_cell_6t_5 inst_cell_64_44 (.BL(BL44),.BLN(BLN44),.WL(WL64));
sram_cell_6t_5 inst_cell_64_45 (.BL(BL45),.BLN(BLN45),.WL(WL64));
sram_cell_6t_5 inst_cell_64_46 (.BL(BL46),.BLN(BLN46),.WL(WL64));
sram_cell_6t_5 inst_cell_64_47 (.BL(BL47),.BLN(BLN47),.WL(WL64));
sram_cell_6t_5 inst_cell_64_48 (.BL(BL48),.BLN(BLN48),.WL(WL64));
sram_cell_6t_5 inst_cell_64_49 (.BL(BL49),.BLN(BLN49),.WL(WL64));
sram_cell_6t_5 inst_cell_64_50 (.BL(BL50),.BLN(BLN50),.WL(WL64));
sram_cell_6t_5 inst_cell_64_51 (.BL(BL51),.BLN(BLN51),.WL(WL64));
sram_cell_6t_5 inst_cell_64_52 (.BL(BL52),.BLN(BLN52),.WL(WL64));
sram_cell_6t_5 inst_cell_64_53 (.BL(BL53),.BLN(BLN53),.WL(WL64));
sram_cell_6t_5 inst_cell_64_54 (.BL(BL54),.BLN(BLN54),.WL(WL64));
sram_cell_6t_5 inst_cell_64_55 (.BL(BL55),.BLN(BLN55),.WL(WL64));
sram_cell_6t_5 inst_cell_64_56 (.BL(BL56),.BLN(BLN56),.WL(WL64));
sram_cell_6t_5 inst_cell_64_57 (.BL(BL57),.BLN(BLN57),.WL(WL64));
sram_cell_6t_5 inst_cell_64_58 (.BL(BL58),.BLN(BLN58),.WL(WL64));
sram_cell_6t_5 inst_cell_64_59 (.BL(BL59),.BLN(BLN59),.WL(WL64));
sram_cell_6t_5 inst_cell_64_60 (.BL(BL60),.BLN(BLN60),.WL(WL64));
sram_cell_6t_5 inst_cell_64_61 (.BL(BL61),.BLN(BLN61),.WL(WL64));
sram_cell_6t_5 inst_cell_64_62 (.BL(BL62),.BLN(BLN62),.WL(WL64));
sram_cell_6t_5 inst_cell_64_63 (.BL(BL63),.BLN(BLN63),.WL(WL64));
sram_cell_6t_5 inst_cell_64_64 (.BL(BL64),.BLN(BLN64),.WL(WL64));
sram_cell_6t_5 inst_cell_64_65 (.BL(BL65),.BLN(BLN65),.WL(WL64));
sram_cell_6t_5 inst_cell_64_66 (.BL(BL66),.BLN(BLN66),.WL(WL64));
sram_cell_6t_5 inst_cell_64_67 (.BL(BL67),.BLN(BLN67),.WL(WL64));
sram_cell_6t_5 inst_cell_64_68 (.BL(BL68),.BLN(BLN68),.WL(WL64));
sram_cell_6t_5 inst_cell_64_69 (.BL(BL69),.BLN(BLN69),.WL(WL64));
sram_cell_6t_5 inst_cell_64_70 (.BL(BL70),.BLN(BLN70),.WL(WL64));
sram_cell_6t_5 inst_cell_64_71 (.BL(BL71),.BLN(BLN71),.WL(WL64));
sram_cell_6t_5 inst_cell_64_72 (.BL(BL72),.BLN(BLN72),.WL(WL64));
sram_cell_6t_5 inst_cell_64_73 (.BL(BL73),.BLN(BLN73),.WL(WL64));
sram_cell_6t_5 inst_cell_64_74 (.BL(BL74),.BLN(BLN74),.WL(WL64));
sram_cell_6t_5 inst_cell_64_75 (.BL(BL75),.BLN(BLN75),.WL(WL64));
sram_cell_6t_5 inst_cell_64_76 (.BL(BL76),.BLN(BLN76),.WL(WL64));
sram_cell_6t_5 inst_cell_64_77 (.BL(BL77),.BLN(BLN77),.WL(WL64));
sram_cell_6t_5 inst_cell_64_78 (.BL(BL78),.BLN(BLN78),.WL(WL64));
sram_cell_6t_5 inst_cell_64_79 (.BL(BL79),.BLN(BLN79),.WL(WL64));
sram_cell_6t_5 inst_cell_64_80 (.BL(BL80),.BLN(BLN80),.WL(WL64));
sram_cell_6t_5 inst_cell_64_81 (.BL(BL81),.BLN(BLN81),.WL(WL64));
sram_cell_6t_5 inst_cell_64_82 (.BL(BL82),.BLN(BLN82),.WL(WL64));
sram_cell_6t_5 inst_cell_64_83 (.BL(BL83),.BLN(BLN83),.WL(WL64));
sram_cell_6t_5 inst_cell_64_84 (.BL(BL84),.BLN(BLN84),.WL(WL64));
sram_cell_6t_5 inst_cell_64_85 (.BL(BL85),.BLN(BLN85),.WL(WL64));
sram_cell_6t_5 inst_cell_64_86 (.BL(BL86),.BLN(BLN86),.WL(WL64));
sram_cell_6t_5 inst_cell_64_87 (.BL(BL87),.BLN(BLN87),.WL(WL64));
sram_cell_6t_5 inst_cell_64_88 (.BL(BL88),.BLN(BLN88),.WL(WL64));
sram_cell_6t_5 inst_cell_64_89 (.BL(BL89),.BLN(BLN89),.WL(WL64));
sram_cell_6t_5 inst_cell_64_90 (.BL(BL90),.BLN(BLN90),.WL(WL64));
sram_cell_6t_5 inst_cell_64_91 (.BL(BL91),.BLN(BLN91),.WL(WL64));
sram_cell_6t_5 inst_cell_64_92 (.BL(BL92),.BLN(BLN92),.WL(WL64));
sram_cell_6t_5 inst_cell_64_93 (.BL(BL93),.BLN(BLN93),.WL(WL64));
sram_cell_6t_5 inst_cell_64_94 (.BL(BL94),.BLN(BLN94),.WL(WL64));
sram_cell_6t_5 inst_cell_64_95 (.BL(BL95),.BLN(BLN95),.WL(WL64));
sram_cell_6t_5 inst_cell_64_96 (.BL(BL96),.BLN(BLN96),.WL(WL64));
sram_cell_6t_5 inst_cell_64_97 (.BL(BL97),.BLN(BLN97),.WL(WL64));
sram_cell_6t_5 inst_cell_64_98 (.BL(BL98),.BLN(BLN98),.WL(WL64));
sram_cell_6t_5 inst_cell_64_99 (.BL(BL99),.BLN(BLN99),.WL(WL64));
sram_cell_6t_5 inst_cell_64_100 (.BL(BL100),.BLN(BLN100),.WL(WL64));
sram_cell_6t_5 inst_cell_64_101 (.BL(BL101),.BLN(BLN101),.WL(WL64));
sram_cell_6t_5 inst_cell_64_102 (.BL(BL102),.BLN(BLN102),.WL(WL64));
sram_cell_6t_5 inst_cell_64_103 (.BL(BL103),.BLN(BLN103),.WL(WL64));
sram_cell_6t_5 inst_cell_64_104 (.BL(BL104),.BLN(BLN104),.WL(WL64));
sram_cell_6t_5 inst_cell_64_105 (.BL(BL105),.BLN(BLN105),.WL(WL64));
sram_cell_6t_5 inst_cell_64_106 (.BL(BL106),.BLN(BLN106),.WL(WL64));
sram_cell_6t_5 inst_cell_64_107 (.BL(BL107),.BLN(BLN107),.WL(WL64));
sram_cell_6t_5 inst_cell_64_108 (.BL(BL108),.BLN(BLN108),.WL(WL64));
sram_cell_6t_5 inst_cell_64_109 (.BL(BL109),.BLN(BLN109),.WL(WL64));
sram_cell_6t_5 inst_cell_64_110 (.BL(BL110),.BLN(BLN110),.WL(WL64));
sram_cell_6t_5 inst_cell_64_111 (.BL(BL111),.BLN(BLN111),.WL(WL64));
sram_cell_6t_5 inst_cell_64_112 (.BL(BL112),.BLN(BLN112),.WL(WL64));
sram_cell_6t_5 inst_cell_64_113 (.BL(BL113),.BLN(BLN113),.WL(WL64));
sram_cell_6t_5 inst_cell_64_114 (.BL(BL114),.BLN(BLN114),.WL(WL64));
sram_cell_6t_5 inst_cell_64_115 (.BL(BL115),.BLN(BLN115),.WL(WL64));
sram_cell_6t_5 inst_cell_64_116 (.BL(BL116),.BLN(BLN116),.WL(WL64));
sram_cell_6t_5 inst_cell_64_117 (.BL(BL117),.BLN(BLN117),.WL(WL64));
sram_cell_6t_5 inst_cell_64_118 (.BL(BL118),.BLN(BLN118),.WL(WL64));
sram_cell_6t_5 inst_cell_64_119 (.BL(BL119),.BLN(BLN119),.WL(WL64));
sram_cell_6t_5 inst_cell_64_120 (.BL(BL120),.BLN(BLN120),.WL(WL64));
sram_cell_6t_5 inst_cell_64_121 (.BL(BL121),.BLN(BLN121),.WL(WL64));
sram_cell_6t_5 inst_cell_64_122 (.BL(BL122),.BLN(BLN122),.WL(WL64));
sram_cell_6t_5 inst_cell_64_123 (.BL(BL123),.BLN(BLN123),.WL(WL64));
sram_cell_6t_5 inst_cell_64_124 (.BL(BL124),.BLN(BLN124),.WL(WL64));
sram_cell_6t_5 inst_cell_64_125 (.BL(BL125),.BLN(BLN125),.WL(WL64));
sram_cell_6t_5 inst_cell_64_126 (.BL(BL126),.BLN(BLN126),.WL(WL64));
sram_cell_6t_5 inst_cell_64_127 (.BL(BL127),.BLN(BLN127),.WL(WL64));
sram_cell_6t_5 inst_cell_65_0 (.BL(BL0),.BLN(BLN0),.WL(WL65));
sram_cell_6t_5 inst_cell_65_1 (.BL(BL1),.BLN(BLN1),.WL(WL65));
sram_cell_6t_5 inst_cell_65_2 (.BL(BL2),.BLN(BLN2),.WL(WL65));
sram_cell_6t_5 inst_cell_65_3 (.BL(BL3),.BLN(BLN3),.WL(WL65));
sram_cell_6t_5 inst_cell_65_4 (.BL(BL4),.BLN(BLN4),.WL(WL65));
sram_cell_6t_5 inst_cell_65_5 (.BL(BL5),.BLN(BLN5),.WL(WL65));
sram_cell_6t_5 inst_cell_65_6 (.BL(BL6),.BLN(BLN6),.WL(WL65));
sram_cell_6t_5 inst_cell_65_7 (.BL(BL7),.BLN(BLN7),.WL(WL65));
sram_cell_6t_5 inst_cell_65_8 (.BL(BL8),.BLN(BLN8),.WL(WL65));
sram_cell_6t_5 inst_cell_65_9 (.BL(BL9),.BLN(BLN9),.WL(WL65));
sram_cell_6t_5 inst_cell_65_10 (.BL(BL10),.BLN(BLN10),.WL(WL65));
sram_cell_6t_5 inst_cell_65_11 (.BL(BL11),.BLN(BLN11),.WL(WL65));
sram_cell_6t_5 inst_cell_65_12 (.BL(BL12),.BLN(BLN12),.WL(WL65));
sram_cell_6t_5 inst_cell_65_13 (.BL(BL13),.BLN(BLN13),.WL(WL65));
sram_cell_6t_5 inst_cell_65_14 (.BL(BL14),.BLN(BLN14),.WL(WL65));
sram_cell_6t_5 inst_cell_65_15 (.BL(BL15),.BLN(BLN15),.WL(WL65));
sram_cell_6t_5 inst_cell_65_16 (.BL(BL16),.BLN(BLN16),.WL(WL65));
sram_cell_6t_5 inst_cell_65_17 (.BL(BL17),.BLN(BLN17),.WL(WL65));
sram_cell_6t_5 inst_cell_65_18 (.BL(BL18),.BLN(BLN18),.WL(WL65));
sram_cell_6t_5 inst_cell_65_19 (.BL(BL19),.BLN(BLN19),.WL(WL65));
sram_cell_6t_5 inst_cell_65_20 (.BL(BL20),.BLN(BLN20),.WL(WL65));
sram_cell_6t_5 inst_cell_65_21 (.BL(BL21),.BLN(BLN21),.WL(WL65));
sram_cell_6t_5 inst_cell_65_22 (.BL(BL22),.BLN(BLN22),.WL(WL65));
sram_cell_6t_5 inst_cell_65_23 (.BL(BL23),.BLN(BLN23),.WL(WL65));
sram_cell_6t_5 inst_cell_65_24 (.BL(BL24),.BLN(BLN24),.WL(WL65));
sram_cell_6t_5 inst_cell_65_25 (.BL(BL25),.BLN(BLN25),.WL(WL65));
sram_cell_6t_5 inst_cell_65_26 (.BL(BL26),.BLN(BLN26),.WL(WL65));
sram_cell_6t_5 inst_cell_65_27 (.BL(BL27),.BLN(BLN27),.WL(WL65));
sram_cell_6t_5 inst_cell_65_28 (.BL(BL28),.BLN(BLN28),.WL(WL65));
sram_cell_6t_5 inst_cell_65_29 (.BL(BL29),.BLN(BLN29),.WL(WL65));
sram_cell_6t_5 inst_cell_65_30 (.BL(BL30),.BLN(BLN30),.WL(WL65));
sram_cell_6t_5 inst_cell_65_31 (.BL(BL31),.BLN(BLN31),.WL(WL65));
sram_cell_6t_5 inst_cell_65_32 (.BL(BL32),.BLN(BLN32),.WL(WL65));
sram_cell_6t_5 inst_cell_65_33 (.BL(BL33),.BLN(BLN33),.WL(WL65));
sram_cell_6t_5 inst_cell_65_34 (.BL(BL34),.BLN(BLN34),.WL(WL65));
sram_cell_6t_5 inst_cell_65_35 (.BL(BL35),.BLN(BLN35),.WL(WL65));
sram_cell_6t_5 inst_cell_65_36 (.BL(BL36),.BLN(BLN36),.WL(WL65));
sram_cell_6t_5 inst_cell_65_37 (.BL(BL37),.BLN(BLN37),.WL(WL65));
sram_cell_6t_5 inst_cell_65_38 (.BL(BL38),.BLN(BLN38),.WL(WL65));
sram_cell_6t_5 inst_cell_65_39 (.BL(BL39),.BLN(BLN39),.WL(WL65));
sram_cell_6t_5 inst_cell_65_40 (.BL(BL40),.BLN(BLN40),.WL(WL65));
sram_cell_6t_5 inst_cell_65_41 (.BL(BL41),.BLN(BLN41),.WL(WL65));
sram_cell_6t_5 inst_cell_65_42 (.BL(BL42),.BLN(BLN42),.WL(WL65));
sram_cell_6t_5 inst_cell_65_43 (.BL(BL43),.BLN(BLN43),.WL(WL65));
sram_cell_6t_5 inst_cell_65_44 (.BL(BL44),.BLN(BLN44),.WL(WL65));
sram_cell_6t_5 inst_cell_65_45 (.BL(BL45),.BLN(BLN45),.WL(WL65));
sram_cell_6t_5 inst_cell_65_46 (.BL(BL46),.BLN(BLN46),.WL(WL65));
sram_cell_6t_5 inst_cell_65_47 (.BL(BL47),.BLN(BLN47),.WL(WL65));
sram_cell_6t_5 inst_cell_65_48 (.BL(BL48),.BLN(BLN48),.WL(WL65));
sram_cell_6t_5 inst_cell_65_49 (.BL(BL49),.BLN(BLN49),.WL(WL65));
sram_cell_6t_5 inst_cell_65_50 (.BL(BL50),.BLN(BLN50),.WL(WL65));
sram_cell_6t_5 inst_cell_65_51 (.BL(BL51),.BLN(BLN51),.WL(WL65));
sram_cell_6t_5 inst_cell_65_52 (.BL(BL52),.BLN(BLN52),.WL(WL65));
sram_cell_6t_5 inst_cell_65_53 (.BL(BL53),.BLN(BLN53),.WL(WL65));
sram_cell_6t_5 inst_cell_65_54 (.BL(BL54),.BLN(BLN54),.WL(WL65));
sram_cell_6t_5 inst_cell_65_55 (.BL(BL55),.BLN(BLN55),.WL(WL65));
sram_cell_6t_5 inst_cell_65_56 (.BL(BL56),.BLN(BLN56),.WL(WL65));
sram_cell_6t_5 inst_cell_65_57 (.BL(BL57),.BLN(BLN57),.WL(WL65));
sram_cell_6t_5 inst_cell_65_58 (.BL(BL58),.BLN(BLN58),.WL(WL65));
sram_cell_6t_5 inst_cell_65_59 (.BL(BL59),.BLN(BLN59),.WL(WL65));
sram_cell_6t_5 inst_cell_65_60 (.BL(BL60),.BLN(BLN60),.WL(WL65));
sram_cell_6t_5 inst_cell_65_61 (.BL(BL61),.BLN(BLN61),.WL(WL65));
sram_cell_6t_5 inst_cell_65_62 (.BL(BL62),.BLN(BLN62),.WL(WL65));
sram_cell_6t_5 inst_cell_65_63 (.BL(BL63),.BLN(BLN63),.WL(WL65));
sram_cell_6t_5 inst_cell_65_64 (.BL(BL64),.BLN(BLN64),.WL(WL65));
sram_cell_6t_5 inst_cell_65_65 (.BL(BL65),.BLN(BLN65),.WL(WL65));
sram_cell_6t_5 inst_cell_65_66 (.BL(BL66),.BLN(BLN66),.WL(WL65));
sram_cell_6t_5 inst_cell_65_67 (.BL(BL67),.BLN(BLN67),.WL(WL65));
sram_cell_6t_5 inst_cell_65_68 (.BL(BL68),.BLN(BLN68),.WL(WL65));
sram_cell_6t_5 inst_cell_65_69 (.BL(BL69),.BLN(BLN69),.WL(WL65));
sram_cell_6t_5 inst_cell_65_70 (.BL(BL70),.BLN(BLN70),.WL(WL65));
sram_cell_6t_5 inst_cell_65_71 (.BL(BL71),.BLN(BLN71),.WL(WL65));
sram_cell_6t_5 inst_cell_65_72 (.BL(BL72),.BLN(BLN72),.WL(WL65));
sram_cell_6t_5 inst_cell_65_73 (.BL(BL73),.BLN(BLN73),.WL(WL65));
sram_cell_6t_5 inst_cell_65_74 (.BL(BL74),.BLN(BLN74),.WL(WL65));
sram_cell_6t_5 inst_cell_65_75 (.BL(BL75),.BLN(BLN75),.WL(WL65));
sram_cell_6t_5 inst_cell_65_76 (.BL(BL76),.BLN(BLN76),.WL(WL65));
sram_cell_6t_5 inst_cell_65_77 (.BL(BL77),.BLN(BLN77),.WL(WL65));
sram_cell_6t_5 inst_cell_65_78 (.BL(BL78),.BLN(BLN78),.WL(WL65));
sram_cell_6t_5 inst_cell_65_79 (.BL(BL79),.BLN(BLN79),.WL(WL65));
sram_cell_6t_5 inst_cell_65_80 (.BL(BL80),.BLN(BLN80),.WL(WL65));
sram_cell_6t_5 inst_cell_65_81 (.BL(BL81),.BLN(BLN81),.WL(WL65));
sram_cell_6t_5 inst_cell_65_82 (.BL(BL82),.BLN(BLN82),.WL(WL65));
sram_cell_6t_5 inst_cell_65_83 (.BL(BL83),.BLN(BLN83),.WL(WL65));
sram_cell_6t_5 inst_cell_65_84 (.BL(BL84),.BLN(BLN84),.WL(WL65));
sram_cell_6t_5 inst_cell_65_85 (.BL(BL85),.BLN(BLN85),.WL(WL65));
sram_cell_6t_5 inst_cell_65_86 (.BL(BL86),.BLN(BLN86),.WL(WL65));
sram_cell_6t_5 inst_cell_65_87 (.BL(BL87),.BLN(BLN87),.WL(WL65));
sram_cell_6t_5 inst_cell_65_88 (.BL(BL88),.BLN(BLN88),.WL(WL65));
sram_cell_6t_5 inst_cell_65_89 (.BL(BL89),.BLN(BLN89),.WL(WL65));
sram_cell_6t_5 inst_cell_65_90 (.BL(BL90),.BLN(BLN90),.WL(WL65));
sram_cell_6t_5 inst_cell_65_91 (.BL(BL91),.BLN(BLN91),.WL(WL65));
sram_cell_6t_5 inst_cell_65_92 (.BL(BL92),.BLN(BLN92),.WL(WL65));
sram_cell_6t_5 inst_cell_65_93 (.BL(BL93),.BLN(BLN93),.WL(WL65));
sram_cell_6t_5 inst_cell_65_94 (.BL(BL94),.BLN(BLN94),.WL(WL65));
sram_cell_6t_5 inst_cell_65_95 (.BL(BL95),.BLN(BLN95),.WL(WL65));
sram_cell_6t_5 inst_cell_65_96 (.BL(BL96),.BLN(BLN96),.WL(WL65));
sram_cell_6t_5 inst_cell_65_97 (.BL(BL97),.BLN(BLN97),.WL(WL65));
sram_cell_6t_5 inst_cell_65_98 (.BL(BL98),.BLN(BLN98),.WL(WL65));
sram_cell_6t_5 inst_cell_65_99 (.BL(BL99),.BLN(BLN99),.WL(WL65));
sram_cell_6t_5 inst_cell_65_100 (.BL(BL100),.BLN(BLN100),.WL(WL65));
sram_cell_6t_5 inst_cell_65_101 (.BL(BL101),.BLN(BLN101),.WL(WL65));
sram_cell_6t_5 inst_cell_65_102 (.BL(BL102),.BLN(BLN102),.WL(WL65));
sram_cell_6t_5 inst_cell_65_103 (.BL(BL103),.BLN(BLN103),.WL(WL65));
sram_cell_6t_5 inst_cell_65_104 (.BL(BL104),.BLN(BLN104),.WL(WL65));
sram_cell_6t_5 inst_cell_65_105 (.BL(BL105),.BLN(BLN105),.WL(WL65));
sram_cell_6t_5 inst_cell_65_106 (.BL(BL106),.BLN(BLN106),.WL(WL65));
sram_cell_6t_5 inst_cell_65_107 (.BL(BL107),.BLN(BLN107),.WL(WL65));
sram_cell_6t_5 inst_cell_65_108 (.BL(BL108),.BLN(BLN108),.WL(WL65));
sram_cell_6t_5 inst_cell_65_109 (.BL(BL109),.BLN(BLN109),.WL(WL65));
sram_cell_6t_5 inst_cell_65_110 (.BL(BL110),.BLN(BLN110),.WL(WL65));
sram_cell_6t_5 inst_cell_65_111 (.BL(BL111),.BLN(BLN111),.WL(WL65));
sram_cell_6t_5 inst_cell_65_112 (.BL(BL112),.BLN(BLN112),.WL(WL65));
sram_cell_6t_5 inst_cell_65_113 (.BL(BL113),.BLN(BLN113),.WL(WL65));
sram_cell_6t_5 inst_cell_65_114 (.BL(BL114),.BLN(BLN114),.WL(WL65));
sram_cell_6t_5 inst_cell_65_115 (.BL(BL115),.BLN(BLN115),.WL(WL65));
sram_cell_6t_5 inst_cell_65_116 (.BL(BL116),.BLN(BLN116),.WL(WL65));
sram_cell_6t_5 inst_cell_65_117 (.BL(BL117),.BLN(BLN117),.WL(WL65));
sram_cell_6t_5 inst_cell_65_118 (.BL(BL118),.BLN(BLN118),.WL(WL65));
sram_cell_6t_5 inst_cell_65_119 (.BL(BL119),.BLN(BLN119),.WL(WL65));
sram_cell_6t_5 inst_cell_65_120 (.BL(BL120),.BLN(BLN120),.WL(WL65));
sram_cell_6t_5 inst_cell_65_121 (.BL(BL121),.BLN(BLN121),.WL(WL65));
sram_cell_6t_5 inst_cell_65_122 (.BL(BL122),.BLN(BLN122),.WL(WL65));
sram_cell_6t_5 inst_cell_65_123 (.BL(BL123),.BLN(BLN123),.WL(WL65));
sram_cell_6t_5 inst_cell_65_124 (.BL(BL124),.BLN(BLN124),.WL(WL65));
sram_cell_6t_5 inst_cell_65_125 (.BL(BL125),.BLN(BLN125),.WL(WL65));
sram_cell_6t_5 inst_cell_65_126 (.BL(BL126),.BLN(BLN126),.WL(WL65));
sram_cell_6t_5 inst_cell_65_127 (.BL(BL127),.BLN(BLN127),.WL(WL65));
sram_cell_6t_5 inst_cell_66_0 (.BL(BL0),.BLN(BLN0),.WL(WL66));
sram_cell_6t_5 inst_cell_66_1 (.BL(BL1),.BLN(BLN1),.WL(WL66));
sram_cell_6t_5 inst_cell_66_2 (.BL(BL2),.BLN(BLN2),.WL(WL66));
sram_cell_6t_5 inst_cell_66_3 (.BL(BL3),.BLN(BLN3),.WL(WL66));
sram_cell_6t_5 inst_cell_66_4 (.BL(BL4),.BLN(BLN4),.WL(WL66));
sram_cell_6t_5 inst_cell_66_5 (.BL(BL5),.BLN(BLN5),.WL(WL66));
sram_cell_6t_5 inst_cell_66_6 (.BL(BL6),.BLN(BLN6),.WL(WL66));
sram_cell_6t_5 inst_cell_66_7 (.BL(BL7),.BLN(BLN7),.WL(WL66));
sram_cell_6t_5 inst_cell_66_8 (.BL(BL8),.BLN(BLN8),.WL(WL66));
sram_cell_6t_5 inst_cell_66_9 (.BL(BL9),.BLN(BLN9),.WL(WL66));
sram_cell_6t_5 inst_cell_66_10 (.BL(BL10),.BLN(BLN10),.WL(WL66));
sram_cell_6t_5 inst_cell_66_11 (.BL(BL11),.BLN(BLN11),.WL(WL66));
sram_cell_6t_5 inst_cell_66_12 (.BL(BL12),.BLN(BLN12),.WL(WL66));
sram_cell_6t_5 inst_cell_66_13 (.BL(BL13),.BLN(BLN13),.WL(WL66));
sram_cell_6t_5 inst_cell_66_14 (.BL(BL14),.BLN(BLN14),.WL(WL66));
sram_cell_6t_5 inst_cell_66_15 (.BL(BL15),.BLN(BLN15),.WL(WL66));
sram_cell_6t_5 inst_cell_66_16 (.BL(BL16),.BLN(BLN16),.WL(WL66));
sram_cell_6t_5 inst_cell_66_17 (.BL(BL17),.BLN(BLN17),.WL(WL66));
sram_cell_6t_5 inst_cell_66_18 (.BL(BL18),.BLN(BLN18),.WL(WL66));
sram_cell_6t_5 inst_cell_66_19 (.BL(BL19),.BLN(BLN19),.WL(WL66));
sram_cell_6t_5 inst_cell_66_20 (.BL(BL20),.BLN(BLN20),.WL(WL66));
sram_cell_6t_5 inst_cell_66_21 (.BL(BL21),.BLN(BLN21),.WL(WL66));
sram_cell_6t_5 inst_cell_66_22 (.BL(BL22),.BLN(BLN22),.WL(WL66));
sram_cell_6t_5 inst_cell_66_23 (.BL(BL23),.BLN(BLN23),.WL(WL66));
sram_cell_6t_5 inst_cell_66_24 (.BL(BL24),.BLN(BLN24),.WL(WL66));
sram_cell_6t_5 inst_cell_66_25 (.BL(BL25),.BLN(BLN25),.WL(WL66));
sram_cell_6t_5 inst_cell_66_26 (.BL(BL26),.BLN(BLN26),.WL(WL66));
sram_cell_6t_5 inst_cell_66_27 (.BL(BL27),.BLN(BLN27),.WL(WL66));
sram_cell_6t_5 inst_cell_66_28 (.BL(BL28),.BLN(BLN28),.WL(WL66));
sram_cell_6t_5 inst_cell_66_29 (.BL(BL29),.BLN(BLN29),.WL(WL66));
sram_cell_6t_5 inst_cell_66_30 (.BL(BL30),.BLN(BLN30),.WL(WL66));
sram_cell_6t_5 inst_cell_66_31 (.BL(BL31),.BLN(BLN31),.WL(WL66));
sram_cell_6t_5 inst_cell_66_32 (.BL(BL32),.BLN(BLN32),.WL(WL66));
sram_cell_6t_5 inst_cell_66_33 (.BL(BL33),.BLN(BLN33),.WL(WL66));
sram_cell_6t_5 inst_cell_66_34 (.BL(BL34),.BLN(BLN34),.WL(WL66));
sram_cell_6t_5 inst_cell_66_35 (.BL(BL35),.BLN(BLN35),.WL(WL66));
sram_cell_6t_5 inst_cell_66_36 (.BL(BL36),.BLN(BLN36),.WL(WL66));
sram_cell_6t_5 inst_cell_66_37 (.BL(BL37),.BLN(BLN37),.WL(WL66));
sram_cell_6t_5 inst_cell_66_38 (.BL(BL38),.BLN(BLN38),.WL(WL66));
sram_cell_6t_5 inst_cell_66_39 (.BL(BL39),.BLN(BLN39),.WL(WL66));
sram_cell_6t_5 inst_cell_66_40 (.BL(BL40),.BLN(BLN40),.WL(WL66));
sram_cell_6t_5 inst_cell_66_41 (.BL(BL41),.BLN(BLN41),.WL(WL66));
sram_cell_6t_5 inst_cell_66_42 (.BL(BL42),.BLN(BLN42),.WL(WL66));
sram_cell_6t_5 inst_cell_66_43 (.BL(BL43),.BLN(BLN43),.WL(WL66));
sram_cell_6t_5 inst_cell_66_44 (.BL(BL44),.BLN(BLN44),.WL(WL66));
sram_cell_6t_5 inst_cell_66_45 (.BL(BL45),.BLN(BLN45),.WL(WL66));
sram_cell_6t_5 inst_cell_66_46 (.BL(BL46),.BLN(BLN46),.WL(WL66));
sram_cell_6t_5 inst_cell_66_47 (.BL(BL47),.BLN(BLN47),.WL(WL66));
sram_cell_6t_5 inst_cell_66_48 (.BL(BL48),.BLN(BLN48),.WL(WL66));
sram_cell_6t_5 inst_cell_66_49 (.BL(BL49),.BLN(BLN49),.WL(WL66));
sram_cell_6t_5 inst_cell_66_50 (.BL(BL50),.BLN(BLN50),.WL(WL66));
sram_cell_6t_5 inst_cell_66_51 (.BL(BL51),.BLN(BLN51),.WL(WL66));
sram_cell_6t_5 inst_cell_66_52 (.BL(BL52),.BLN(BLN52),.WL(WL66));
sram_cell_6t_5 inst_cell_66_53 (.BL(BL53),.BLN(BLN53),.WL(WL66));
sram_cell_6t_5 inst_cell_66_54 (.BL(BL54),.BLN(BLN54),.WL(WL66));
sram_cell_6t_5 inst_cell_66_55 (.BL(BL55),.BLN(BLN55),.WL(WL66));
sram_cell_6t_5 inst_cell_66_56 (.BL(BL56),.BLN(BLN56),.WL(WL66));
sram_cell_6t_5 inst_cell_66_57 (.BL(BL57),.BLN(BLN57),.WL(WL66));
sram_cell_6t_5 inst_cell_66_58 (.BL(BL58),.BLN(BLN58),.WL(WL66));
sram_cell_6t_5 inst_cell_66_59 (.BL(BL59),.BLN(BLN59),.WL(WL66));
sram_cell_6t_5 inst_cell_66_60 (.BL(BL60),.BLN(BLN60),.WL(WL66));
sram_cell_6t_5 inst_cell_66_61 (.BL(BL61),.BLN(BLN61),.WL(WL66));
sram_cell_6t_5 inst_cell_66_62 (.BL(BL62),.BLN(BLN62),.WL(WL66));
sram_cell_6t_5 inst_cell_66_63 (.BL(BL63),.BLN(BLN63),.WL(WL66));
sram_cell_6t_5 inst_cell_66_64 (.BL(BL64),.BLN(BLN64),.WL(WL66));
sram_cell_6t_5 inst_cell_66_65 (.BL(BL65),.BLN(BLN65),.WL(WL66));
sram_cell_6t_5 inst_cell_66_66 (.BL(BL66),.BLN(BLN66),.WL(WL66));
sram_cell_6t_5 inst_cell_66_67 (.BL(BL67),.BLN(BLN67),.WL(WL66));
sram_cell_6t_5 inst_cell_66_68 (.BL(BL68),.BLN(BLN68),.WL(WL66));
sram_cell_6t_5 inst_cell_66_69 (.BL(BL69),.BLN(BLN69),.WL(WL66));
sram_cell_6t_5 inst_cell_66_70 (.BL(BL70),.BLN(BLN70),.WL(WL66));
sram_cell_6t_5 inst_cell_66_71 (.BL(BL71),.BLN(BLN71),.WL(WL66));
sram_cell_6t_5 inst_cell_66_72 (.BL(BL72),.BLN(BLN72),.WL(WL66));
sram_cell_6t_5 inst_cell_66_73 (.BL(BL73),.BLN(BLN73),.WL(WL66));
sram_cell_6t_5 inst_cell_66_74 (.BL(BL74),.BLN(BLN74),.WL(WL66));
sram_cell_6t_5 inst_cell_66_75 (.BL(BL75),.BLN(BLN75),.WL(WL66));
sram_cell_6t_5 inst_cell_66_76 (.BL(BL76),.BLN(BLN76),.WL(WL66));
sram_cell_6t_5 inst_cell_66_77 (.BL(BL77),.BLN(BLN77),.WL(WL66));
sram_cell_6t_5 inst_cell_66_78 (.BL(BL78),.BLN(BLN78),.WL(WL66));
sram_cell_6t_5 inst_cell_66_79 (.BL(BL79),.BLN(BLN79),.WL(WL66));
sram_cell_6t_5 inst_cell_66_80 (.BL(BL80),.BLN(BLN80),.WL(WL66));
sram_cell_6t_5 inst_cell_66_81 (.BL(BL81),.BLN(BLN81),.WL(WL66));
sram_cell_6t_5 inst_cell_66_82 (.BL(BL82),.BLN(BLN82),.WL(WL66));
sram_cell_6t_5 inst_cell_66_83 (.BL(BL83),.BLN(BLN83),.WL(WL66));
sram_cell_6t_5 inst_cell_66_84 (.BL(BL84),.BLN(BLN84),.WL(WL66));
sram_cell_6t_5 inst_cell_66_85 (.BL(BL85),.BLN(BLN85),.WL(WL66));
sram_cell_6t_5 inst_cell_66_86 (.BL(BL86),.BLN(BLN86),.WL(WL66));
sram_cell_6t_5 inst_cell_66_87 (.BL(BL87),.BLN(BLN87),.WL(WL66));
sram_cell_6t_5 inst_cell_66_88 (.BL(BL88),.BLN(BLN88),.WL(WL66));
sram_cell_6t_5 inst_cell_66_89 (.BL(BL89),.BLN(BLN89),.WL(WL66));
sram_cell_6t_5 inst_cell_66_90 (.BL(BL90),.BLN(BLN90),.WL(WL66));
sram_cell_6t_5 inst_cell_66_91 (.BL(BL91),.BLN(BLN91),.WL(WL66));
sram_cell_6t_5 inst_cell_66_92 (.BL(BL92),.BLN(BLN92),.WL(WL66));
sram_cell_6t_5 inst_cell_66_93 (.BL(BL93),.BLN(BLN93),.WL(WL66));
sram_cell_6t_5 inst_cell_66_94 (.BL(BL94),.BLN(BLN94),.WL(WL66));
sram_cell_6t_5 inst_cell_66_95 (.BL(BL95),.BLN(BLN95),.WL(WL66));
sram_cell_6t_5 inst_cell_66_96 (.BL(BL96),.BLN(BLN96),.WL(WL66));
sram_cell_6t_5 inst_cell_66_97 (.BL(BL97),.BLN(BLN97),.WL(WL66));
sram_cell_6t_5 inst_cell_66_98 (.BL(BL98),.BLN(BLN98),.WL(WL66));
sram_cell_6t_5 inst_cell_66_99 (.BL(BL99),.BLN(BLN99),.WL(WL66));
sram_cell_6t_5 inst_cell_66_100 (.BL(BL100),.BLN(BLN100),.WL(WL66));
sram_cell_6t_5 inst_cell_66_101 (.BL(BL101),.BLN(BLN101),.WL(WL66));
sram_cell_6t_5 inst_cell_66_102 (.BL(BL102),.BLN(BLN102),.WL(WL66));
sram_cell_6t_5 inst_cell_66_103 (.BL(BL103),.BLN(BLN103),.WL(WL66));
sram_cell_6t_5 inst_cell_66_104 (.BL(BL104),.BLN(BLN104),.WL(WL66));
sram_cell_6t_5 inst_cell_66_105 (.BL(BL105),.BLN(BLN105),.WL(WL66));
sram_cell_6t_5 inst_cell_66_106 (.BL(BL106),.BLN(BLN106),.WL(WL66));
sram_cell_6t_5 inst_cell_66_107 (.BL(BL107),.BLN(BLN107),.WL(WL66));
sram_cell_6t_5 inst_cell_66_108 (.BL(BL108),.BLN(BLN108),.WL(WL66));
sram_cell_6t_5 inst_cell_66_109 (.BL(BL109),.BLN(BLN109),.WL(WL66));
sram_cell_6t_5 inst_cell_66_110 (.BL(BL110),.BLN(BLN110),.WL(WL66));
sram_cell_6t_5 inst_cell_66_111 (.BL(BL111),.BLN(BLN111),.WL(WL66));
sram_cell_6t_5 inst_cell_66_112 (.BL(BL112),.BLN(BLN112),.WL(WL66));
sram_cell_6t_5 inst_cell_66_113 (.BL(BL113),.BLN(BLN113),.WL(WL66));
sram_cell_6t_5 inst_cell_66_114 (.BL(BL114),.BLN(BLN114),.WL(WL66));
sram_cell_6t_5 inst_cell_66_115 (.BL(BL115),.BLN(BLN115),.WL(WL66));
sram_cell_6t_5 inst_cell_66_116 (.BL(BL116),.BLN(BLN116),.WL(WL66));
sram_cell_6t_5 inst_cell_66_117 (.BL(BL117),.BLN(BLN117),.WL(WL66));
sram_cell_6t_5 inst_cell_66_118 (.BL(BL118),.BLN(BLN118),.WL(WL66));
sram_cell_6t_5 inst_cell_66_119 (.BL(BL119),.BLN(BLN119),.WL(WL66));
sram_cell_6t_5 inst_cell_66_120 (.BL(BL120),.BLN(BLN120),.WL(WL66));
sram_cell_6t_5 inst_cell_66_121 (.BL(BL121),.BLN(BLN121),.WL(WL66));
sram_cell_6t_5 inst_cell_66_122 (.BL(BL122),.BLN(BLN122),.WL(WL66));
sram_cell_6t_5 inst_cell_66_123 (.BL(BL123),.BLN(BLN123),.WL(WL66));
sram_cell_6t_5 inst_cell_66_124 (.BL(BL124),.BLN(BLN124),.WL(WL66));
sram_cell_6t_5 inst_cell_66_125 (.BL(BL125),.BLN(BLN125),.WL(WL66));
sram_cell_6t_5 inst_cell_66_126 (.BL(BL126),.BLN(BLN126),.WL(WL66));
sram_cell_6t_5 inst_cell_66_127 (.BL(BL127),.BLN(BLN127),.WL(WL66));
sram_cell_6t_5 inst_cell_67_0 (.BL(BL0),.BLN(BLN0),.WL(WL67));
sram_cell_6t_5 inst_cell_67_1 (.BL(BL1),.BLN(BLN1),.WL(WL67));
sram_cell_6t_5 inst_cell_67_2 (.BL(BL2),.BLN(BLN2),.WL(WL67));
sram_cell_6t_5 inst_cell_67_3 (.BL(BL3),.BLN(BLN3),.WL(WL67));
sram_cell_6t_5 inst_cell_67_4 (.BL(BL4),.BLN(BLN4),.WL(WL67));
sram_cell_6t_5 inst_cell_67_5 (.BL(BL5),.BLN(BLN5),.WL(WL67));
sram_cell_6t_5 inst_cell_67_6 (.BL(BL6),.BLN(BLN6),.WL(WL67));
sram_cell_6t_5 inst_cell_67_7 (.BL(BL7),.BLN(BLN7),.WL(WL67));
sram_cell_6t_5 inst_cell_67_8 (.BL(BL8),.BLN(BLN8),.WL(WL67));
sram_cell_6t_5 inst_cell_67_9 (.BL(BL9),.BLN(BLN9),.WL(WL67));
sram_cell_6t_5 inst_cell_67_10 (.BL(BL10),.BLN(BLN10),.WL(WL67));
sram_cell_6t_5 inst_cell_67_11 (.BL(BL11),.BLN(BLN11),.WL(WL67));
sram_cell_6t_5 inst_cell_67_12 (.BL(BL12),.BLN(BLN12),.WL(WL67));
sram_cell_6t_5 inst_cell_67_13 (.BL(BL13),.BLN(BLN13),.WL(WL67));
sram_cell_6t_5 inst_cell_67_14 (.BL(BL14),.BLN(BLN14),.WL(WL67));
sram_cell_6t_5 inst_cell_67_15 (.BL(BL15),.BLN(BLN15),.WL(WL67));
sram_cell_6t_5 inst_cell_67_16 (.BL(BL16),.BLN(BLN16),.WL(WL67));
sram_cell_6t_5 inst_cell_67_17 (.BL(BL17),.BLN(BLN17),.WL(WL67));
sram_cell_6t_5 inst_cell_67_18 (.BL(BL18),.BLN(BLN18),.WL(WL67));
sram_cell_6t_5 inst_cell_67_19 (.BL(BL19),.BLN(BLN19),.WL(WL67));
sram_cell_6t_5 inst_cell_67_20 (.BL(BL20),.BLN(BLN20),.WL(WL67));
sram_cell_6t_5 inst_cell_67_21 (.BL(BL21),.BLN(BLN21),.WL(WL67));
sram_cell_6t_5 inst_cell_67_22 (.BL(BL22),.BLN(BLN22),.WL(WL67));
sram_cell_6t_5 inst_cell_67_23 (.BL(BL23),.BLN(BLN23),.WL(WL67));
sram_cell_6t_5 inst_cell_67_24 (.BL(BL24),.BLN(BLN24),.WL(WL67));
sram_cell_6t_5 inst_cell_67_25 (.BL(BL25),.BLN(BLN25),.WL(WL67));
sram_cell_6t_5 inst_cell_67_26 (.BL(BL26),.BLN(BLN26),.WL(WL67));
sram_cell_6t_5 inst_cell_67_27 (.BL(BL27),.BLN(BLN27),.WL(WL67));
sram_cell_6t_5 inst_cell_67_28 (.BL(BL28),.BLN(BLN28),.WL(WL67));
sram_cell_6t_5 inst_cell_67_29 (.BL(BL29),.BLN(BLN29),.WL(WL67));
sram_cell_6t_5 inst_cell_67_30 (.BL(BL30),.BLN(BLN30),.WL(WL67));
sram_cell_6t_5 inst_cell_67_31 (.BL(BL31),.BLN(BLN31),.WL(WL67));
sram_cell_6t_5 inst_cell_67_32 (.BL(BL32),.BLN(BLN32),.WL(WL67));
sram_cell_6t_5 inst_cell_67_33 (.BL(BL33),.BLN(BLN33),.WL(WL67));
sram_cell_6t_5 inst_cell_67_34 (.BL(BL34),.BLN(BLN34),.WL(WL67));
sram_cell_6t_5 inst_cell_67_35 (.BL(BL35),.BLN(BLN35),.WL(WL67));
sram_cell_6t_5 inst_cell_67_36 (.BL(BL36),.BLN(BLN36),.WL(WL67));
sram_cell_6t_5 inst_cell_67_37 (.BL(BL37),.BLN(BLN37),.WL(WL67));
sram_cell_6t_5 inst_cell_67_38 (.BL(BL38),.BLN(BLN38),.WL(WL67));
sram_cell_6t_5 inst_cell_67_39 (.BL(BL39),.BLN(BLN39),.WL(WL67));
sram_cell_6t_5 inst_cell_67_40 (.BL(BL40),.BLN(BLN40),.WL(WL67));
sram_cell_6t_5 inst_cell_67_41 (.BL(BL41),.BLN(BLN41),.WL(WL67));
sram_cell_6t_5 inst_cell_67_42 (.BL(BL42),.BLN(BLN42),.WL(WL67));
sram_cell_6t_5 inst_cell_67_43 (.BL(BL43),.BLN(BLN43),.WL(WL67));
sram_cell_6t_5 inst_cell_67_44 (.BL(BL44),.BLN(BLN44),.WL(WL67));
sram_cell_6t_5 inst_cell_67_45 (.BL(BL45),.BLN(BLN45),.WL(WL67));
sram_cell_6t_5 inst_cell_67_46 (.BL(BL46),.BLN(BLN46),.WL(WL67));
sram_cell_6t_5 inst_cell_67_47 (.BL(BL47),.BLN(BLN47),.WL(WL67));
sram_cell_6t_5 inst_cell_67_48 (.BL(BL48),.BLN(BLN48),.WL(WL67));
sram_cell_6t_5 inst_cell_67_49 (.BL(BL49),.BLN(BLN49),.WL(WL67));
sram_cell_6t_5 inst_cell_67_50 (.BL(BL50),.BLN(BLN50),.WL(WL67));
sram_cell_6t_5 inst_cell_67_51 (.BL(BL51),.BLN(BLN51),.WL(WL67));
sram_cell_6t_5 inst_cell_67_52 (.BL(BL52),.BLN(BLN52),.WL(WL67));
sram_cell_6t_5 inst_cell_67_53 (.BL(BL53),.BLN(BLN53),.WL(WL67));
sram_cell_6t_5 inst_cell_67_54 (.BL(BL54),.BLN(BLN54),.WL(WL67));
sram_cell_6t_5 inst_cell_67_55 (.BL(BL55),.BLN(BLN55),.WL(WL67));
sram_cell_6t_5 inst_cell_67_56 (.BL(BL56),.BLN(BLN56),.WL(WL67));
sram_cell_6t_5 inst_cell_67_57 (.BL(BL57),.BLN(BLN57),.WL(WL67));
sram_cell_6t_5 inst_cell_67_58 (.BL(BL58),.BLN(BLN58),.WL(WL67));
sram_cell_6t_5 inst_cell_67_59 (.BL(BL59),.BLN(BLN59),.WL(WL67));
sram_cell_6t_5 inst_cell_67_60 (.BL(BL60),.BLN(BLN60),.WL(WL67));
sram_cell_6t_5 inst_cell_67_61 (.BL(BL61),.BLN(BLN61),.WL(WL67));
sram_cell_6t_5 inst_cell_67_62 (.BL(BL62),.BLN(BLN62),.WL(WL67));
sram_cell_6t_5 inst_cell_67_63 (.BL(BL63),.BLN(BLN63),.WL(WL67));
sram_cell_6t_5 inst_cell_67_64 (.BL(BL64),.BLN(BLN64),.WL(WL67));
sram_cell_6t_5 inst_cell_67_65 (.BL(BL65),.BLN(BLN65),.WL(WL67));
sram_cell_6t_5 inst_cell_67_66 (.BL(BL66),.BLN(BLN66),.WL(WL67));
sram_cell_6t_5 inst_cell_67_67 (.BL(BL67),.BLN(BLN67),.WL(WL67));
sram_cell_6t_5 inst_cell_67_68 (.BL(BL68),.BLN(BLN68),.WL(WL67));
sram_cell_6t_5 inst_cell_67_69 (.BL(BL69),.BLN(BLN69),.WL(WL67));
sram_cell_6t_5 inst_cell_67_70 (.BL(BL70),.BLN(BLN70),.WL(WL67));
sram_cell_6t_5 inst_cell_67_71 (.BL(BL71),.BLN(BLN71),.WL(WL67));
sram_cell_6t_5 inst_cell_67_72 (.BL(BL72),.BLN(BLN72),.WL(WL67));
sram_cell_6t_5 inst_cell_67_73 (.BL(BL73),.BLN(BLN73),.WL(WL67));
sram_cell_6t_5 inst_cell_67_74 (.BL(BL74),.BLN(BLN74),.WL(WL67));
sram_cell_6t_5 inst_cell_67_75 (.BL(BL75),.BLN(BLN75),.WL(WL67));
sram_cell_6t_5 inst_cell_67_76 (.BL(BL76),.BLN(BLN76),.WL(WL67));
sram_cell_6t_5 inst_cell_67_77 (.BL(BL77),.BLN(BLN77),.WL(WL67));
sram_cell_6t_5 inst_cell_67_78 (.BL(BL78),.BLN(BLN78),.WL(WL67));
sram_cell_6t_5 inst_cell_67_79 (.BL(BL79),.BLN(BLN79),.WL(WL67));
sram_cell_6t_5 inst_cell_67_80 (.BL(BL80),.BLN(BLN80),.WL(WL67));
sram_cell_6t_5 inst_cell_67_81 (.BL(BL81),.BLN(BLN81),.WL(WL67));
sram_cell_6t_5 inst_cell_67_82 (.BL(BL82),.BLN(BLN82),.WL(WL67));
sram_cell_6t_5 inst_cell_67_83 (.BL(BL83),.BLN(BLN83),.WL(WL67));
sram_cell_6t_5 inst_cell_67_84 (.BL(BL84),.BLN(BLN84),.WL(WL67));
sram_cell_6t_5 inst_cell_67_85 (.BL(BL85),.BLN(BLN85),.WL(WL67));
sram_cell_6t_5 inst_cell_67_86 (.BL(BL86),.BLN(BLN86),.WL(WL67));
sram_cell_6t_5 inst_cell_67_87 (.BL(BL87),.BLN(BLN87),.WL(WL67));
sram_cell_6t_5 inst_cell_67_88 (.BL(BL88),.BLN(BLN88),.WL(WL67));
sram_cell_6t_5 inst_cell_67_89 (.BL(BL89),.BLN(BLN89),.WL(WL67));
sram_cell_6t_5 inst_cell_67_90 (.BL(BL90),.BLN(BLN90),.WL(WL67));
sram_cell_6t_5 inst_cell_67_91 (.BL(BL91),.BLN(BLN91),.WL(WL67));
sram_cell_6t_5 inst_cell_67_92 (.BL(BL92),.BLN(BLN92),.WL(WL67));
sram_cell_6t_5 inst_cell_67_93 (.BL(BL93),.BLN(BLN93),.WL(WL67));
sram_cell_6t_5 inst_cell_67_94 (.BL(BL94),.BLN(BLN94),.WL(WL67));
sram_cell_6t_5 inst_cell_67_95 (.BL(BL95),.BLN(BLN95),.WL(WL67));
sram_cell_6t_5 inst_cell_67_96 (.BL(BL96),.BLN(BLN96),.WL(WL67));
sram_cell_6t_5 inst_cell_67_97 (.BL(BL97),.BLN(BLN97),.WL(WL67));
sram_cell_6t_5 inst_cell_67_98 (.BL(BL98),.BLN(BLN98),.WL(WL67));
sram_cell_6t_5 inst_cell_67_99 (.BL(BL99),.BLN(BLN99),.WL(WL67));
sram_cell_6t_5 inst_cell_67_100 (.BL(BL100),.BLN(BLN100),.WL(WL67));
sram_cell_6t_5 inst_cell_67_101 (.BL(BL101),.BLN(BLN101),.WL(WL67));
sram_cell_6t_5 inst_cell_67_102 (.BL(BL102),.BLN(BLN102),.WL(WL67));
sram_cell_6t_5 inst_cell_67_103 (.BL(BL103),.BLN(BLN103),.WL(WL67));
sram_cell_6t_5 inst_cell_67_104 (.BL(BL104),.BLN(BLN104),.WL(WL67));
sram_cell_6t_5 inst_cell_67_105 (.BL(BL105),.BLN(BLN105),.WL(WL67));
sram_cell_6t_5 inst_cell_67_106 (.BL(BL106),.BLN(BLN106),.WL(WL67));
sram_cell_6t_5 inst_cell_67_107 (.BL(BL107),.BLN(BLN107),.WL(WL67));
sram_cell_6t_5 inst_cell_67_108 (.BL(BL108),.BLN(BLN108),.WL(WL67));
sram_cell_6t_5 inst_cell_67_109 (.BL(BL109),.BLN(BLN109),.WL(WL67));
sram_cell_6t_5 inst_cell_67_110 (.BL(BL110),.BLN(BLN110),.WL(WL67));
sram_cell_6t_5 inst_cell_67_111 (.BL(BL111),.BLN(BLN111),.WL(WL67));
sram_cell_6t_5 inst_cell_67_112 (.BL(BL112),.BLN(BLN112),.WL(WL67));
sram_cell_6t_5 inst_cell_67_113 (.BL(BL113),.BLN(BLN113),.WL(WL67));
sram_cell_6t_5 inst_cell_67_114 (.BL(BL114),.BLN(BLN114),.WL(WL67));
sram_cell_6t_5 inst_cell_67_115 (.BL(BL115),.BLN(BLN115),.WL(WL67));
sram_cell_6t_5 inst_cell_67_116 (.BL(BL116),.BLN(BLN116),.WL(WL67));
sram_cell_6t_5 inst_cell_67_117 (.BL(BL117),.BLN(BLN117),.WL(WL67));
sram_cell_6t_5 inst_cell_67_118 (.BL(BL118),.BLN(BLN118),.WL(WL67));
sram_cell_6t_5 inst_cell_67_119 (.BL(BL119),.BLN(BLN119),.WL(WL67));
sram_cell_6t_5 inst_cell_67_120 (.BL(BL120),.BLN(BLN120),.WL(WL67));
sram_cell_6t_5 inst_cell_67_121 (.BL(BL121),.BLN(BLN121),.WL(WL67));
sram_cell_6t_5 inst_cell_67_122 (.BL(BL122),.BLN(BLN122),.WL(WL67));
sram_cell_6t_5 inst_cell_67_123 (.BL(BL123),.BLN(BLN123),.WL(WL67));
sram_cell_6t_5 inst_cell_67_124 (.BL(BL124),.BLN(BLN124),.WL(WL67));
sram_cell_6t_5 inst_cell_67_125 (.BL(BL125),.BLN(BLN125),.WL(WL67));
sram_cell_6t_5 inst_cell_67_126 (.BL(BL126),.BLN(BLN126),.WL(WL67));
sram_cell_6t_5 inst_cell_67_127 (.BL(BL127),.BLN(BLN127),.WL(WL67));
sram_cell_6t_5 inst_cell_68_0 (.BL(BL0),.BLN(BLN0),.WL(WL68));
sram_cell_6t_5 inst_cell_68_1 (.BL(BL1),.BLN(BLN1),.WL(WL68));
sram_cell_6t_5 inst_cell_68_2 (.BL(BL2),.BLN(BLN2),.WL(WL68));
sram_cell_6t_5 inst_cell_68_3 (.BL(BL3),.BLN(BLN3),.WL(WL68));
sram_cell_6t_5 inst_cell_68_4 (.BL(BL4),.BLN(BLN4),.WL(WL68));
sram_cell_6t_5 inst_cell_68_5 (.BL(BL5),.BLN(BLN5),.WL(WL68));
sram_cell_6t_5 inst_cell_68_6 (.BL(BL6),.BLN(BLN6),.WL(WL68));
sram_cell_6t_5 inst_cell_68_7 (.BL(BL7),.BLN(BLN7),.WL(WL68));
sram_cell_6t_5 inst_cell_68_8 (.BL(BL8),.BLN(BLN8),.WL(WL68));
sram_cell_6t_5 inst_cell_68_9 (.BL(BL9),.BLN(BLN9),.WL(WL68));
sram_cell_6t_5 inst_cell_68_10 (.BL(BL10),.BLN(BLN10),.WL(WL68));
sram_cell_6t_5 inst_cell_68_11 (.BL(BL11),.BLN(BLN11),.WL(WL68));
sram_cell_6t_5 inst_cell_68_12 (.BL(BL12),.BLN(BLN12),.WL(WL68));
sram_cell_6t_5 inst_cell_68_13 (.BL(BL13),.BLN(BLN13),.WL(WL68));
sram_cell_6t_5 inst_cell_68_14 (.BL(BL14),.BLN(BLN14),.WL(WL68));
sram_cell_6t_5 inst_cell_68_15 (.BL(BL15),.BLN(BLN15),.WL(WL68));
sram_cell_6t_5 inst_cell_68_16 (.BL(BL16),.BLN(BLN16),.WL(WL68));
sram_cell_6t_5 inst_cell_68_17 (.BL(BL17),.BLN(BLN17),.WL(WL68));
sram_cell_6t_5 inst_cell_68_18 (.BL(BL18),.BLN(BLN18),.WL(WL68));
sram_cell_6t_5 inst_cell_68_19 (.BL(BL19),.BLN(BLN19),.WL(WL68));
sram_cell_6t_5 inst_cell_68_20 (.BL(BL20),.BLN(BLN20),.WL(WL68));
sram_cell_6t_5 inst_cell_68_21 (.BL(BL21),.BLN(BLN21),.WL(WL68));
sram_cell_6t_5 inst_cell_68_22 (.BL(BL22),.BLN(BLN22),.WL(WL68));
sram_cell_6t_5 inst_cell_68_23 (.BL(BL23),.BLN(BLN23),.WL(WL68));
sram_cell_6t_5 inst_cell_68_24 (.BL(BL24),.BLN(BLN24),.WL(WL68));
sram_cell_6t_5 inst_cell_68_25 (.BL(BL25),.BLN(BLN25),.WL(WL68));
sram_cell_6t_5 inst_cell_68_26 (.BL(BL26),.BLN(BLN26),.WL(WL68));
sram_cell_6t_5 inst_cell_68_27 (.BL(BL27),.BLN(BLN27),.WL(WL68));
sram_cell_6t_5 inst_cell_68_28 (.BL(BL28),.BLN(BLN28),.WL(WL68));
sram_cell_6t_5 inst_cell_68_29 (.BL(BL29),.BLN(BLN29),.WL(WL68));
sram_cell_6t_5 inst_cell_68_30 (.BL(BL30),.BLN(BLN30),.WL(WL68));
sram_cell_6t_5 inst_cell_68_31 (.BL(BL31),.BLN(BLN31),.WL(WL68));
sram_cell_6t_5 inst_cell_68_32 (.BL(BL32),.BLN(BLN32),.WL(WL68));
sram_cell_6t_5 inst_cell_68_33 (.BL(BL33),.BLN(BLN33),.WL(WL68));
sram_cell_6t_5 inst_cell_68_34 (.BL(BL34),.BLN(BLN34),.WL(WL68));
sram_cell_6t_5 inst_cell_68_35 (.BL(BL35),.BLN(BLN35),.WL(WL68));
sram_cell_6t_5 inst_cell_68_36 (.BL(BL36),.BLN(BLN36),.WL(WL68));
sram_cell_6t_5 inst_cell_68_37 (.BL(BL37),.BLN(BLN37),.WL(WL68));
sram_cell_6t_5 inst_cell_68_38 (.BL(BL38),.BLN(BLN38),.WL(WL68));
sram_cell_6t_5 inst_cell_68_39 (.BL(BL39),.BLN(BLN39),.WL(WL68));
sram_cell_6t_5 inst_cell_68_40 (.BL(BL40),.BLN(BLN40),.WL(WL68));
sram_cell_6t_5 inst_cell_68_41 (.BL(BL41),.BLN(BLN41),.WL(WL68));
sram_cell_6t_5 inst_cell_68_42 (.BL(BL42),.BLN(BLN42),.WL(WL68));
sram_cell_6t_5 inst_cell_68_43 (.BL(BL43),.BLN(BLN43),.WL(WL68));
sram_cell_6t_5 inst_cell_68_44 (.BL(BL44),.BLN(BLN44),.WL(WL68));
sram_cell_6t_5 inst_cell_68_45 (.BL(BL45),.BLN(BLN45),.WL(WL68));
sram_cell_6t_5 inst_cell_68_46 (.BL(BL46),.BLN(BLN46),.WL(WL68));
sram_cell_6t_5 inst_cell_68_47 (.BL(BL47),.BLN(BLN47),.WL(WL68));
sram_cell_6t_5 inst_cell_68_48 (.BL(BL48),.BLN(BLN48),.WL(WL68));
sram_cell_6t_5 inst_cell_68_49 (.BL(BL49),.BLN(BLN49),.WL(WL68));
sram_cell_6t_5 inst_cell_68_50 (.BL(BL50),.BLN(BLN50),.WL(WL68));
sram_cell_6t_5 inst_cell_68_51 (.BL(BL51),.BLN(BLN51),.WL(WL68));
sram_cell_6t_5 inst_cell_68_52 (.BL(BL52),.BLN(BLN52),.WL(WL68));
sram_cell_6t_5 inst_cell_68_53 (.BL(BL53),.BLN(BLN53),.WL(WL68));
sram_cell_6t_5 inst_cell_68_54 (.BL(BL54),.BLN(BLN54),.WL(WL68));
sram_cell_6t_5 inst_cell_68_55 (.BL(BL55),.BLN(BLN55),.WL(WL68));
sram_cell_6t_5 inst_cell_68_56 (.BL(BL56),.BLN(BLN56),.WL(WL68));
sram_cell_6t_5 inst_cell_68_57 (.BL(BL57),.BLN(BLN57),.WL(WL68));
sram_cell_6t_5 inst_cell_68_58 (.BL(BL58),.BLN(BLN58),.WL(WL68));
sram_cell_6t_5 inst_cell_68_59 (.BL(BL59),.BLN(BLN59),.WL(WL68));
sram_cell_6t_5 inst_cell_68_60 (.BL(BL60),.BLN(BLN60),.WL(WL68));
sram_cell_6t_5 inst_cell_68_61 (.BL(BL61),.BLN(BLN61),.WL(WL68));
sram_cell_6t_5 inst_cell_68_62 (.BL(BL62),.BLN(BLN62),.WL(WL68));
sram_cell_6t_5 inst_cell_68_63 (.BL(BL63),.BLN(BLN63),.WL(WL68));
sram_cell_6t_5 inst_cell_68_64 (.BL(BL64),.BLN(BLN64),.WL(WL68));
sram_cell_6t_5 inst_cell_68_65 (.BL(BL65),.BLN(BLN65),.WL(WL68));
sram_cell_6t_5 inst_cell_68_66 (.BL(BL66),.BLN(BLN66),.WL(WL68));
sram_cell_6t_5 inst_cell_68_67 (.BL(BL67),.BLN(BLN67),.WL(WL68));
sram_cell_6t_5 inst_cell_68_68 (.BL(BL68),.BLN(BLN68),.WL(WL68));
sram_cell_6t_5 inst_cell_68_69 (.BL(BL69),.BLN(BLN69),.WL(WL68));
sram_cell_6t_5 inst_cell_68_70 (.BL(BL70),.BLN(BLN70),.WL(WL68));
sram_cell_6t_5 inst_cell_68_71 (.BL(BL71),.BLN(BLN71),.WL(WL68));
sram_cell_6t_5 inst_cell_68_72 (.BL(BL72),.BLN(BLN72),.WL(WL68));
sram_cell_6t_5 inst_cell_68_73 (.BL(BL73),.BLN(BLN73),.WL(WL68));
sram_cell_6t_5 inst_cell_68_74 (.BL(BL74),.BLN(BLN74),.WL(WL68));
sram_cell_6t_5 inst_cell_68_75 (.BL(BL75),.BLN(BLN75),.WL(WL68));
sram_cell_6t_5 inst_cell_68_76 (.BL(BL76),.BLN(BLN76),.WL(WL68));
sram_cell_6t_5 inst_cell_68_77 (.BL(BL77),.BLN(BLN77),.WL(WL68));
sram_cell_6t_5 inst_cell_68_78 (.BL(BL78),.BLN(BLN78),.WL(WL68));
sram_cell_6t_5 inst_cell_68_79 (.BL(BL79),.BLN(BLN79),.WL(WL68));
sram_cell_6t_5 inst_cell_68_80 (.BL(BL80),.BLN(BLN80),.WL(WL68));
sram_cell_6t_5 inst_cell_68_81 (.BL(BL81),.BLN(BLN81),.WL(WL68));
sram_cell_6t_5 inst_cell_68_82 (.BL(BL82),.BLN(BLN82),.WL(WL68));
sram_cell_6t_5 inst_cell_68_83 (.BL(BL83),.BLN(BLN83),.WL(WL68));
sram_cell_6t_5 inst_cell_68_84 (.BL(BL84),.BLN(BLN84),.WL(WL68));
sram_cell_6t_5 inst_cell_68_85 (.BL(BL85),.BLN(BLN85),.WL(WL68));
sram_cell_6t_5 inst_cell_68_86 (.BL(BL86),.BLN(BLN86),.WL(WL68));
sram_cell_6t_5 inst_cell_68_87 (.BL(BL87),.BLN(BLN87),.WL(WL68));
sram_cell_6t_5 inst_cell_68_88 (.BL(BL88),.BLN(BLN88),.WL(WL68));
sram_cell_6t_5 inst_cell_68_89 (.BL(BL89),.BLN(BLN89),.WL(WL68));
sram_cell_6t_5 inst_cell_68_90 (.BL(BL90),.BLN(BLN90),.WL(WL68));
sram_cell_6t_5 inst_cell_68_91 (.BL(BL91),.BLN(BLN91),.WL(WL68));
sram_cell_6t_5 inst_cell_68_92 (.BL(BL92),.BLN(BLN92),.WL(WL68));
sram_cell_6t_5 inst_cell_68_93 (.BL(BL93),.BLN(BLN93),.WL(WL68));
sram_cell_6t_5 inst_cell_68_94 (.BL(BL94),.BLN(BLN94),.WL(WL68));
sram_cell_6t_5 inst_cell_68_95 (.BL(BL95),.BLN(BLN95),.WL(WL68));
sram_cell_6t_5 inst_cell_68_96 (.BL(BL96),.BLN(BLN96),.WL(WL68));
sram_cell_6t_5 inst_cell_68_97 (.BL(BL97),.BLN(BLN97),.WL(WL68));
sram_cell_6t_5 inst_cell_68_98 (.BL(BL98),.BLN(BLN98),.WL(WL68));
sram_cell_6t_5 inst_cell_68_99 (.BL(BL99),.BLN(BLN99),.WL(WL68));
sram_cell_6t_5 inst_cell_68_100 (.BL(BL100),.BLN(BLN100),.WL(WL68));
sram_cell_6t_5 inst_cell_68_101 (.BL(BL101),.BLN(BLN101),.WL(WL68));
sram_cell_6t_5 inst_cell_68_102 (.BL(BL102),.BLN(BLN102),.WL(WL68));
sram_cell_6t_5 inst_cell_68_103 (.BL(BL103),.BLN(BLN103),.WL(WL68));
sram_cell_6t_5 inst_cell_68_104 (.BL(BL104),.BLN(BLN104),.WL(WL68));
sram_cell_6t_5 inst_cell_68_105 (.BL(BL105),.BLN(BLN105),.WL(WL68));
sram_cell_6t_5 inst_cell_68_106 (.BL(BL106),.BLN(BLN106),.WL(WL68));
sram_cell_6t_5 inst_cell_68_107 (.BL(BL107),.BLN(BLN107),.WL(WL68));
sram_cell_6t_5 inst_cell_68_108 (.BL(BL108),.BLN(BLN108),.WL(WL68));
sram_cell_6t_5 inst_cell_68_109 (.BL(BL109),.BLN(BLN109),.WL(WL68));
sram_cell_6t_5 inst_cell_68_110 (.BL(BL110),.BLN(BLN110),.WL(WL68));
sram_cell_6t_5 inst_cell_68_111 (.BL(BL111),.BLN(BLN111),.WL(WL68));
sram_cell_6t_5 inst_cell_68_112 (.BL(BL112),.BLN(BLN112),.WL(WL68));
sram_cell_6t_5 inst_cell_68_113 (.BL(BL113),.BLN(BLN113),.WL(WL68));
sram_cell_6t_5 inst_cell_68_114 (.BL(BL114),.BLN(BLN114),.WL(WL68));
sram_cell_6t_5 inst_cell_68_115 (.BL(BL115),.BLN(BLN115),.WL(WL68));
sram_cell_6t_5 inst_cell_68_116 (.BL(BL116),.BLN(BLN116),.WL(WL68));
sram_cell_6t_5 inst_cell_68_117 (.BL(BL117),.BLN(BLN117),.WL(WL68));
sram_cell_6t_5 inst_cell_68_118 (.BL(BL118),.BLN(BLN118),.WL(WL68));
sram_cell_6t_5 inst_cell_68_119 (.BL(BL119),.BLN(BLN119),.WL(WL68));
sram_cell_6t_5 inst_cell_68_120 (.BL(BL120),.BLN(BLN120),.WL(WL68));
sram_cell_6t_5 inst_cell_68_121 (.BL(BL121),.BLN(BLN121),.WL(WL68));
sram_cell_6t_5 inst_cell_68_122 (.BL(BL122),.BLN(BLN122),.WL(WL68));
sram_cell_6t_5 inst_cell_68_123 (.BL(BL123),.BLN(BLN123),.WL(WL68));
sram_cell_6t_5 inst_cell_68_124 (.BL(BL124),.BLN(BLN124),.WL(WL68));
sram_cell_6t_5 inst_cell_68_125 (.BL(BL125),.BLN(BLN125),.WL(WL68));
sram_cell_6t_5 inst_cell_68_126 (.BL(BL126),.BLN(BLN126),.WL(WL68));
sram_cell_6t_5 inst_cell_68_127 (.BL(BL127),.BLN(BLN127),.WL(WL68));
sram_cell_6t_5 inst_cell_69_0 (.BL(BL0),.BLN(BLN0),.WL(WL69));
sram_cell_6t_5 inst_cell_69_1 (.BL(BL1),.BLN(BLN1),.WL(WL69));
sram_cell_6t_5 inst_cell_69_2 (.BL(BL2),.BLN(BLN2),.WL(WL69));
sram_cell_6t_5 inst_cell_69_3 (.BL(BL3),.BLN(BLN3),.WL(WL69));
sram_cell_6t_5 inst_cell_69_4 (.BL(BL4),.BLN(BLN4),.WL(WL69));
sram_cell_6t_5 inst_cell_69_5 (.BL(BL5),.BLN(BLN5),.WL(WL69));
sram_cell_6t_5 inst_cell_69_6 (.BL(BL6),.BLN(BLN6),.WL(WL69));
sram_cell_6t_5 inst_cell_69_7 (.BL(BL7),.BLN(BLN7),.WL(WL69));
sram_cell_6t_5 inst_cell_69_8 (.BL(BL8),.BLN(BLN8),.WL(WL69));
sram_cell_6t_5 inst_cell_69_9 (.BL(BL9),.BLN(BLN9),.WL(WL69));
sram_cell_6t_5 inst_cell_69_10 (.BL(BL10),.BLN(BLN10),.WL(WL69));
sram_cell_6t_5 inst_cell_69_11 (.BL(BL11),.BLN(BLN11),.WL(WL69));
sram_cell_6t_5 inst_cell_69_12 (.BL(BL12),.BLN(BLN12),.WL(WL69));
sram_cell_6t_5 inst_cell_69_13 (.BL(BL13),.BLN(BLN13),.WL(WL69));
sram_cell_6t_5 inst_cell_69_14 (.BL(BL14),.BLN(BLN14),.WL(WL69));
sram_cell_6t_5 inst_cell_69_15 (.BL(BL15),.BLN(BLN15),.WL(WL69));
sram_cell_6t_5 inst_cell_69_16 (.BL(BL16),.BLN(BLN16),.WL(WL69));
sram_cell_6t_5 inst_cell_69_17 (.BL(BL17),.BLN(BLN17),.WL(WL69));
sram_cell_6t_5 inst_cell_69_18 (.BL(BL18),.BLN(BLN18),.WL(WL69));
sram_cell_6t_5 inst_cell_69_19 (.BL(BL19),.BLN(BLN19),.WL(WL69));
sram_cell_6t_5 inst_cell_69_20 (.BL(BL20),.BLN(BLN20),.WL(WL69));
sram_cell_6t_5 inst_cell_69_21 (.BL(BL21),.BLN(BLN21),.WL(WL69));
sram_cell_6t_5 inst_cell_69_22 (.BL(BL22),.BLN(BLN22),.WL(WL69));
sram_cell_6t_5 inst_cell_69_23 (.BL(BL23),.BLN(BLN23),.WL(WL69));
sram_cell_6t_5 inst_cell_69_24 (.BL(BL24),.BLN(BLN24),.WL(WL69));
sram_cell_6t_5 inst_cell_69_25 (.BL(BL25),.BLN(BLN25),.WL(WL69));
sram_cell_6t_5 inst_cell_69_26 (.BL(BL26),.BLN(BLN26),.WL(WL69));
sram_cell_6t_5 inst_cell_69_27 (.BL(BL27),.BLN(BLN27),.WL(WL69));
sram_cell_6t_5 inst_cell_69_28 (.BL(BL28),.BLN(BLN28),.WL(WL69));
sram_cell_6t_5 inst_cell_69_29 (.BL(BL29),.BLN(BLN29),.WL(WL69));
sram_cell_6t_5 inst_cell_69_30 (.BL(BL30),.BLN(BLN30),.WL(WL69));
sram_cell_6t_5 inst_cell_69_31 (.BL(BL31),.BLN(BLN31),.WL(WL69));
sram_cell_6t_5 inst_cell_69_32 (.BL(BL32),.BLN(BLN32),.WL(WL69));
sram_cell_6t_5 inst_cell_69_33 (.BL(BL33),.BLN(BLN33),.WL(WL69));
sram_cell_6t_5 inst_cell_69_34 (.BL(BL34),.BLN(BLN34),.WL(WL69));
sram_cell_6t_5 inst_cell_69_35 (.BL(BL35),.BLN(BLN35),.WL(WL69));
sram_cell_6t_5 inst_cell_69_36 (.BL(BL36),.BLN(BLN36),.WL(WL69));
sram_cell_6t_5 inst_cell_69_37 (.BL(BL37),.BLN(BLN37),.WL(WL69));
sram_cell_6t_5 inst_cell_69_38 (.BL(BL38),.BLN(BLN38),.WL(WL69));
sram_cell_6t_5 inst_cell_69_39 (.BL(BL39),.BLN(BLN39),.WL(WL69));
sram_cell_6t_5 inst_cell_69_40 (.BL(BL40),.BLN(BLN40),.WL(WL69));
sram_cell_6t_5 inst_cell_69_41 (.BL(BL41),.BLN(BLN41),.WL(WL69));
sram_cell_6t_5 inst_cell_69_42 (.BL(BL42),.BLN(BLN42),.WL(WL69));
sram_cell_6t_5 inst_cell_69_43 (.BL(BL43),.BLN(BLN43),.WL(WL69));
sram_cell_6t_5 inst_cell_69_44 (.BL(BL44),.BLN(BLN44),.WL(WL69));
sram_cell_6t_5 inst_cell_69_45 (.BL(BL45),.BLN(BLN45),.WL(WL69));
sram_cell_6t_5 inst_cell_69_46 (.BL(BL46),.BLN(BLN46),.WL(WL69));
sram_cell_6t_5 inst_cell_69_47 (.BL(BL47),.BLN(BLN47),.WL(WL69));
sram_cell_6t_5 inst_cell_69_48 (.BL(BL48),.BLN(BLN48),.WL(WL69));
sram_cell_6t_5 inst_cell_69_49 (.BL(BL49),.BLN(BLN49),.WL(WL69));
sram_cell_6t_5 inst_cell_69_50 (.BL(BL50),.BLN(BLN50),.WL(WL69));
sram_cell_6t_5 inst_cell_69_51 (.BL(BL51),.BLN(BLN51),.WL(WL69));
sram_cell_6t_5 inst_cell_69_52 (.BL(BL52),.BLN(BLN52),.WL(WL69));
sram_cell_6t_5 inst_cell_69_53 (.BL(BL53),.BLN(BLN53),.WL(WL69));
sram_cell_6t_5 inst_cell_69_54 (.BL(BL54),.BLN(BLN54),.WL(WL69));
sram_cell_6t_5 inst_cell_69_55 (.BL(BL55),.BLN(BLN55),.WL(WL69));
sram_cell_6t_5 inst_cell_69_56 (.BL(BL56),.BLN(BLN56),.WL(WL69));
sram_cell_6t_5 inst_cell_69_57 (.BL(BL57),.BLN(BLN57),.WL(WL69));
sram_cell_6t_5 inst_cell_69_58 (.BL(BL58),.BLN(BLN58),.WL(WL69));
sram_cell_6t_5 inst_cell_69_59 (.BL(BL59),.BLN(BLN59),.WL(WL69));
sram_cell_6t_5 inst_cell_69_60 (.BL(BL60),.BLN(BLN60),.WL(WL69));
sram_cell_6t_5 inst_cell_69_61 (.BL(BL61),.BLN(BLN61),.WL(WL69));
sram_cell_6t_5 inst_cell_69_62 (.BL(BL62),.BLN(BLN62),.WL(WL69));
sram_cell_6t_5 inst_cell_69_63 (.BL(BL63),.BLN(BLN63),.WL(WL69));
sram_cell_6t_5 inst_cell_69_64 (.BL(BL64),.BLN(BLN64),.WL(WL69));
sram_cell_6t_5 inst_cell_69_65 (.BL(BL65),.BLN(BLN65),.WL(WL69));
sram_cell_6t_5 inst_cell_69_66 (.BL(BL66),.BLN(BLN66),.WL(WL69));
sram_cell_6t_5 inst_cell_69_67 (.BL(BL67),.BLN(BLN67),.WL(WL69));
sram_cell_6t_5 inst_cell_69_68 (.BL(BL68),.BLN(BLN68),.WL(WL69));
sram_cell_6t_5 inst_cell_69_69 (.BL(BL69),.BLN(BLN69),.WL(WL69));
sram_cell_6t_5 inst_cell_69_70 (.BL(BL70),.BLN(BLN70),.WL(WL69));
sram_cell_6t_5 inst_cell_69_71 (.BL(BL71),.BLN(BLN71),.WL(WL69));
sram_cell_6t_5 inst_cell_69_72 (.BL(BL72),.BLN(BLN72),.WL(WL69));
sram_cell_6t_5 inst_cell_69_73 (.BL(BL73),.BLN(BLN73),.WL(WL69));
sram_cell_6t_5 inst_cell_69_74 (.BL(BL74),.BLN(BLN74),.WL(WL69));
sram_cell_6t_5 inst_cell_69_75 (.BL(BL75),.BLN(BLN75),.WL(WL69));
sram_cell_6t_5 inst_cell_69_76 (.BL(BL76),.BLN(BLN76),.WL(WL69));
sram_cell_6t_5 inst_cell_69_77 (.BL(BL77),.BLN(BLN77),.WL(WL69));
sram_cell_6t_5 inst_cell_69_78 (.BL(BL78),.BLN(BLN78),.WL(WL69));
sram_cell_6t_5 inst_cell_69_79 (.BL(BL79),.BLN(BLN79),.WL(WL69));
sram_cell_6t_5 inst_cell_69_80 (.BL(BL80),.BLN(BLN80),.WL(WL69));
sram_cell_6t_5 inst_cell_69_81 (.BL(BL81),.BLN(BLN81),.WL(WL69));
sram_cell_6t_5 inst_cell_69_82 (.BL(BL82),.BLN(BLN82),.WL(WL69));
sram_cell_6t_5 inst_cell_69_83 (.BL(BL83),.BLN(BLN83),.WL(WL69));
sram_cell_6t_5 inst_cell_69_84 (.BL(BL84),.BLN(BLN84),.WL(WL69));
sram_cell_6t_5 inst_cell_69_85 (.BL(BL85),.BLN(BLN85),.WL(WL69));
sram_cell_6t_5 inst_cell_69_86 (.BL(BL86),.BLN(BLN86),.WL(WL69));
sram_cell_6t_5 inst_cell_69_87 (.BL(BL87),.BLN(BLN87),.WL(WL69));
sram_cell_6t_5 inst_cell_69_88 (.BL(BL88),.BLN(BLN88),.WL(WL69));
sram_cell_6t_5 inst_cell_69_89 (.BL(BL89),.BLN(BLN89),.WL(WL69));
sram_cell_6t_5 inst_cell_69_90 (.BL(BL90),.BLN(BLN90),.WL(WL69));
sram_cell_6t_5 inst_cell_69_91 (.BL(BL91),.BLN(BLN91),.WL(WL69));
sram_cell_6t_5 inst_cell_69_92 (.BL(BL92),.BLN(BLN92),.WL(WL69));
sram_cell_6t_5 inst_cell_69_93 (.BL(BL93),.BLN(BLN93),.WL(WL69));
sram_cell_6t_5 inst_cell_69_94 (.BL(BL94),.BLN(BLN94),.WL(WL69));
sram_cell_6t_5 inst_cell_69_95 (.BL(BL95),.BLN(BLN95),.WL(WL69));
sram_cell_6t_5 inst_cell_69_96 (.BL(BL96),.BLN(BLN96),.WL(WL69));
sram_cell_6t_5 inst_cell_69_97 (.BL(BL97),.BLN(BLN97),.WL(WL69));
sram_cell_6t_5 inst_cell_69_98 (.BL(BL98),.BLN(BLN98),.WL(WL69));
sram_cell_6t_5 inst_cell_69_99 (.BL(BL99),.BLN(BLN99),.WL(WL69));
sram_cell_6t_5 inst_cell_69_100 (.BL(BL100),.BLN(BLN100),.WL(WL69));
sram_cell_6t_5 inst_cell_69_101 (.BL(BL101),.BLN(BLN101),.WL(WL69));
sram_cell_6t_5 inst_cell_69_102 (.BL(BL102),.BLN(BLN102),.WL(WL69));
sram_cell_6t_5 inst_cell_69_103 (.BL(BL103),.BLN(BLN103),.WL(WL69));
sram_cell_6t_5 inst_cell_69_104 (.BL(BL104),.BLN(BLN104),.WL(WL69));
sram_cell_6t_5 inst_cell_69_105 (.BL(BL105),.BLN(BLN105),.WL(WL69));
sram_cell_6t_5 inst_cell_69_106 (.BL(BL106),.BLN(BLN106),.WL(WL69));
sram_cell_6t_5 inst_cell_69_107 (.BL(BL107),.BLN(BLN107),.WL(WL69));
sram_cell_6t_5 inst_cell_69_108 (.BL(BL108),.BLN(BLN108),.WL(WL69));
sram_cell_6t_5 inst_cell_69_109 (.BL(BL109),.BLN(BLN109),.WL(WL69));
sram_cell_6t_5 inst_cell_69_110 (.BL(BL110),.BLN(BLN110),.WL(WL69));
sram_cell_6t_5 inst_cell_69_111 (.BL(BL111),.BLN(BLN111),.WL(WL69));
sram_cell_6t_5 inst_cell_69_112 (.BL(BL112),.BLN(BLN112),.WL(WL69));
sram_cell_6t_5 inst_cell_69_113 (.BL(BL113),.BLN(BLN113),.WL(WL69));
sram_cell_6t_5 inst_cell_69_114 (.BL(BL114),.BLN(BLN114),.WL(WL69));
sram_cell_6t_5 inst_cell_69_115 (.BL(BL115),.BLN(BLN115),.WL(WL69));
sram_cell_6t_5 inst_cell_69_116 (.BL(BL116),.BLN(BLN116),.WL(WL69));
sram_cell_6t_5 inst_cell_69_117 (.BL(BL117),.BLN(BLN117),.WL(WL69));
sram_cell_6t_5 inst_cell_69_118 (.BL(BL118),.BLN(BLN118),.WL(WL69));
sram_cell_6t_5 inst_cell_69_119 (.BL(BL119),.BLN(BLN119),.WL(WL69));
sram_cell_6t_5 inst_cell_69_120 (.BL(BL120),.BLN(BLN120),.WL(WL69));
sram_cell_6t_5 inst_cell_69_121 (.BL(BL121),.BLN(BLN121),.WL(WL69));
sram_cell_6t_5 inst_cell_69_122 (.BL(BL122),.BLN(BLN122),.WL(WL69));
sram_cell_6t_5 inst_cell_69_123 (.BL(BL123),.BLN(BLN123),.WL(WL69));
sram_cell_6t_5 inst_cell_69_124 (.BL(BL124),.BLN(BLN124),.WL(WL69));
sram_cell_6t_5 inst_cell_69_125 (.BL(BL125),.BLN(BLN125),.WL(WL69));
sram_cell_6t_5 inst_cell_69_126 (.BL(BL126),.BLN(BLN126),.WL(WL69));
sram_cell_6t_5 inst_cell_69_127 (.BL(BL127),.BLN(BLN127),.WL(WL69));
sram_cell_6t_5 inst_cell_70_0 (.BL(BL0),.BLN(BLN0),.WL(WL70));
sram_cell_6t_5 inst_cell_70_1 (.BL(BL1),.BLN(BLN1),.WL(WL70));
sram_cell_6t_5 inst_cell_70_2 (.BL(BL2),.BLN(BLN2),.WL(WL70));
sram_cell_6t_5 inst_cell_70_3 (.BL(BL3),.BLN(BLN3),.WL(WL70));
sram_cell_6t_5 inst_cell_70_4 (.BL(BL4),.BLN(BLN4),.WL(WL70));
sram_cell_6t_5 inst_cell_70_5 (.BL(BL5),.BLN(BLN5),.WL(WL70));
sram_cell_6t_5 inst_cell_70_6 (.BL(BL6),.BLN(BLN6),.WL(WL70));
sram_cell_6t_5 inst_cell_70_7 (.BL(BL7),.BLN(BLN7),.WL(WL70));
sram_cell_6t_5 inst_cell_70_8 (.BL(BL8),.BLN(BLN8),.WL(WL70));
sram_cell_6t_5 inst_cell_70_9 (.BL(BL9),.BLN(BLN9),.WL(WL70));
sram_cell_6t_5 inst_cell_70_10 (.BL(BL10),.BLN(BLN10),.WL(WL70));
sram_cell_6t_5 inst_cell_70_11 (.BL(BL11),.BLN(BLN11),.WL(WL70));
sram_cell_6t_5 inst_cell_70_12 (.BL(BL12),.BLN(BLN12),.WL(WL70));
sram_cell_6t_5 inst_cell_70_13 (.BL(BL13),.BLN(BLN13),.WL(WL70));
sram_cell_6t_5 inst_cell_70_14 (.BL(BL14),.BLN(BLN14),.WL(WL70));
sram_cell_6t_5 inst_cell_70_15 (.BL(BL15),.BLN(BLN15),.WL(WL70));
sram_cell_6t_5 inst_cell_70_16 (.BL(BL16),.BLN(BLN16),.WL(WL70));
sram_cell_6t_5 inst_cell_70_17 (.BL(BL17),.BLN(BLN17),.WL(WL70));
sram_cell_6t_5 inst_cell_70_18 (.BL(BL18),.BLN(BLN18),.WL(WL70));
sram_cell_6t_5 inst_cell_70_19 (.BL(BL19),.BLN(BLN19),.WL(WL70));
sram_cell_6t_5 inst_cell_70_20 (.BL(BL20),.BLN(BLN20),.WL(WL70));
sram_cell_6t_5 inst_cell_70_21 (.BL(BL21),.BLN(BLN21),.WL(WL70));
sram_cell_6t_5 inst_cell_70_22 (.BL(BL22),.BLN(BLN22),.WL(WL70));
sram_cell_6t_5 inst_cell_70_23 (.BL(BL23),.BLN(BLN23),.WL(WL70));
sram_cell_6t_5 inst_cell_70_24 (.BL(BL24),.BLN(BLN24),.WL(WL70));
sram_cell_6t_5 inst_cell_70_25 (.BL(BL25),.BLN(BLN25),.WL(WL70));
sram_cell_6t_5 inst_cell_70_26 (.BL(BL26),.BLN(BLN26),.WL(WL70));
sram_cell_6t_5 inst_cell_70_27 (.BL(BL27),.BLN(BLN27),.WL(WL70));
sram_cell_6t_5 inst_cell_70_28 (.BL(BL28),.BLN(BLN28),.WL(WL70));
sram_cell_6t_5 inst_cell_70_29 (.BL(BL29),.BLN(BLN29),.WL(WL70));
sram_cell_6t_5 inst_cell_70_30 (.BL(BL30),.BLN(BLN30),.WL(WL70));
sram_cell_6t_5 inst_cell_70_31 (.BL(BL31),.BLN(BLN31),.WL(WL70));
sram_cell_6t_5 inst_cell_70_32 (.BL(BL32),.BLN(BLN32),.WL(WL70));
sram_cell_6t_5 inst_cell_70_33 (.BL(BL33),.BLN(BLN33),.WL(WL70));
sram_cell_6t_5 inst_cell_70_34 (.BL(BL34),.BLN(BLN34),.WL(WL70));
sram_cell_6t_5 inst_cell_70_35 (.BL(BL35),.BLN(BLN35),.WL(WL70));
sram_cell_6t_5 inst_cell_70_36 (.BL(BL36),.BLN(BLN36),.WL(WL70));
sram_cell_6t_5 inst_cell_70_37 (.BL(BL37),.BLN(BLN37),.WL(WL70));
sram_cell_6t_5 inst_cell_70_38 (.BL(BL38),.BLN(BLN38),.WL(WL70));
sram_cell_6t_5 inst_cell_70_39 (.BL(BL39),.BLN(BLN39),.WL(WL70));
sram_cell_6t_5 inst_cell_70_40 (.BL(BL40),.BLN(BLN40),.WL(WL70));
sram_cell_6t_5 inst_cell_70_41 (.BL(BL41),.BLN(BLN41),.WL(WL70));
sram_cell_6t_5 inst_cell_70_42 (.BL(BL42),.BLN(BLN42),.WL(WL70));
sram_cell_6t_5 inst_cell_70_43 (.BL(BL43),.BLN(BLN43),.WL(WL70));
sram_cell_6t_5 inst_cell_70_44 (.BL(BL44),.BLN(BLN44),.WL(WL70));
sram_cell_6t_5 inst_cell_70_45 (.BL(BL45),.BLN(BLN45),.WL(WL70));
sram_cell_6t_5 inst_cell_70_46 (.BL(BL46),.BLN(BLN46),.WL(WL70));
sram_cell_6t_5 inst_cell_70_47 (.BL(BL47),.BLN(BLN47),.WL(WL70));
sram_cell_6t_5 inst_cell_70_48 (.BL(BL48),.BLN(BLN48),.WL(WL70));
sram_cell_6t_5 inst_cell_70_49 (.BL(BL49),.BLN(BLN49),.WL(WL70));
sram_cell_6t_5 inst_cell_70_50 (.BL(BL50),.BLN(BLN50),.WL(WL70));
sram_cell_6t_5 inst_cell_70_51 (.BL(BL51),.BLN(BLN51),.WL(WL70));
sram_cell_6t_5 inst_cell_70_52 (.BL(BL52),.BLN(BLN52),.WL(WL70));
sram_cell_6t_5 inst_cell_70_53 (.BL(BL53),.BLN(BLN53),.WL(WL70));
sram_cell_6t_5 inst_cell_70_54 (.BL(BL54),.BLN(BLN54),.WL(WL70));
sram_cell_6t_5 inst_cell_70_55 (.BL(BL55),.BLN(BLN55),.WL(WL70));
sram_cell_6t_5 inst_cell_70_56 (.BL(BL56),.BLN(BLN56),.WL(WL70));
sram_cell_6t_5 inst_cell_70_57 (.BL(BL57),.BLN(BLN57),.WL(WL70));
sram_cell_6t_5 inst_cell_70_58 (.BL(BL58),.BLN(BLN58),.WL(WL70));
sram_cell_6t_5 inst_cell_70_59 (.BL(BL59),.BLN(BLN59),.WL(WL70));
sram_cell_6t_5 inst_cell_70_60 (.BL(BL60),.BLN(BLN60),.WL(WL70));
sram_cell_6t_5 inst_cell_70_61 (.BL(BL61),.BLN(BLN61),.WL(WL70));
sram_cell_6t_5 inst_cell_70_62 (.BL(BL62),.BLN(BLN62),.WL(WL70));
sram_cell_6t_5 inst_cell_70_63 (.BL(BL63),.BLN(BLN63),.WL(WL70));
sram_cell_6t_5 inst_cell_70_64 (.BL(BL64),.BLN(BLN64),.WL(WL70));
sram_cell_6t_5 inst_cell_70_65 (.BL(BL65),.BLN(BLN65),.WL(WL70));
sram_cell_6t_5 inst_cell_70_66 (.BL(BL66),.BLN(BLN66),.WL(WL70));
sram_cell_6t_5 inst_cell_70_67 (.BL(BL67),.BLN(BLN67),.WL(WL70));
sram_cell_6t_5 inst_cell_70_68 (.BL(BL68),.BLN(BLN68),.WL(WL70));
sram_cell_6t_5 inst_cell_70_69 (.BL(BL69),.BLN(BLN69),.WL(WL70));
sram_cell_6t_5 inst_cell_70_70 (.BL(BL70),.BLN(BLN70),.WL(WL70));
sram_cell_6t_5 inst_cell_70_71 (.BL(BL71),.BLN(BLN71),.WL(WL70));
sram_cell_6t_5 inst_cell_70_72 (.BL(BL72),.BLN(BLN72),.WL(WL70));
sram_cell_6t_5 inst_cell_70_73 (.BL(BL73),.BLN(BLN73),.WL(WL70));
sram_cell_6t_5 inst_cell_70_74 (.BL(BL74),.BLN(BLN74),.WL(WL70));
sram_cell_6t_5 inst_cell_70_75 (.BL(BL75),.BLN(BLN75),.WL(WL70));
sram_cell_6t_5 inst_cell_70_76 (.BL(BL76),.BLN(BLN76),.WL(WL70));
sram_cell_6t_5 inst_cell_70_77 (.BL(BL77),.BLN(BLN77),.WL(WL70));
sram_cell_6t_5 inst_cell_70_78 (.BL(BL78),.BLN(BLN78),.WL(WL70));
sram_cell_6t_5 inst_cell_70_79 (.BL(BL79),.BLN(BLN79),.WL(WL70));
sram_cell_6t_5 inst_cell_70_80 (.BL(BL80),.BLN(BLN80),.WL(WL70));
sram_cell_6t_5 inst_cell_70_81 (.BL(BL81),.BLN(BLN81),.WL(WL70));
sram_cell_6t_5 inst_cell_70_82 (.BL(BL82),.BLN(BLN82),.WL(WL70));
sram_cell_6t_5 inst_cell_70_83 (.BL(BL83),.BLN(BLN83),.WL(WL70));
sram_cell_6t_5 inst_cell_70_84 (.BL(BL84),.BLN(BLN84),.WL(WL70));
sram_cell_6t_5 inst_cell_70_85 (.BL(BL85),.BLN(BLN85),.WL(WL70));
sram_cell_6t_5 inst_cell_70_86 (.BL(BL86),.BLN(BLN86),.WL(WL70));
sram_cell_6t_5 inst_cell_70_87 (.BL(BL87),.BLN(BLN87),.WL(WL70));
sram_cell_6t_5 inst_cell_70_88 (.BL(BL88),.BLN(BLN88),.WL(WL70));
sram_cell_6t_5 inst_cell_70_89 (.BL(BL89),.BLN(BLN89),.WL(WL70));
sram_cell_6t_5 inst_cell_70_90 (.BL(BL90),.BLN(BLN90),.WL(WL70));
sram_cell_6t_5 inst_cell_70_91 (.BL(BL91),.BLN(BLN91),.WL(WL70));
sram_cell_6t_5 inst_cell_70_92 (.BL(BL92),.BLN(BLN92),.WL(WL70));
sram_cell_6t_5 inst_cell_70_93 (.BL(BL93),.BLN(BLN93),.WL(WL70));
sram_cell_6t_5 inst_cell_70_94 (.BL(BL94),.BLN(BLN94),.WL(WL70));
sram_cell_6t_5 inst_cell_70_95 (.BL(BL95),.BLN(BLN95),.WL(WL70));
sram_cell_6t_5 inst_cell_70_96 (.BL(BL96),.BLN(BLN96),.WL(WL70));
sram_cell_6t_5 inst_cell_70_97 (.BL(BL97),.BLN(BLN97),.WL(WL70));
sram_cell_6t_5 inst_cell_70_98 (.BL(BL98),.BLN(BLN98),.WL(WL70));
sram_cell_6t_5 inst_cell_70_99 (.BL(BL99),.BLN(BLN99),.WL(WL70));
sram_cell_6t_5 inst_cell_70_100 (.BL(BL100),.BLN(BLN100),.WL(WL70));
sram_cell_6t_5 inst_cell_70_101 (.BL(BL101),.BLN(BLN101),.WL(WL70));
sram_cell_6t_5 inst_cell_70_102 (.BL(BL102),.BLN(BLN102),.WL(WL70));
sram_cell_6t_5 inst_cell_70_103 (.BL(BL103),.BLN(BLN103),.WL(WL70));
sram_cell_6t_5 inst_cell_70_104 (.BL(BL104),.BLN(BLN104),.WL(WL70));
sram_cell_6t_5 inst_cell_70_105 (.BL(BL105),.BLN(BLN105),.WL(WL70));
sram_cell_6t_5 inst_cell_70_106 (.BL(BL106),.BLN(BLN106),.WL(WL70));
sram_cell_6t_5 inst_cell_70_107 (.BL(BL107),.BLN(BLN107),.WL(WL70));
sram_cell_6t_5 inst_cell_70_108 (.BL(BL108),.BLN(BLN108),.WL(WL70));
sram_cell_6t_5 inst_cell_70_109 (.BL(BL109),.BLN(BLN109),.WL(WL70));
sram_cell_6t_5 inst_cell_70_110 (.BL(BL110),.BLN(BLN110),.WL(WL70));
sram_cell_6t_5 inst_cell_70_111 (.BL(BL111),.BLN(BLN111),.WL(WL70));
sram_cell_6t_5 inst_cell_70_112 (.BL(BL112),.BLN(BLN112),.WL(WL70));
sram_cell_6t_5 inst_cell_70_113 (.BL(BL113),.BLN(BLN113),.WL(WL70));
sram_cell_6t_5 inst_cell_70_114 (.BL(BL114),.BLN(BLN114),.WL(WL70));
sram_cell_6t_5 inst_cell_70_115 (.BL(BL115),.BLN(BLN115),.WL(WL70));
sram_cell_6t_5 inst_cell_70_116 (.BL(BL116),.BLN(BLN116),.WL(WL70));
sram_cell_6t_5 inst_cell_70_117 (.BL(BL117),.BLN(BLN117),.WL(WL70));
sram_cell_6t_5 inst_cell_70_118 (.BL(BL118),.BLN(BLN118),.WL(WL70));
sram_cell_6t_5 inst_cell_70_119 (.BL(BL119),.BLN(BLN119),.WL(WL70));
sram_cell_6t_5 inst_cell_70_120 (.BL(BL120),.BLN(BLN120),.WL(WL70));
sram_cell_6t_5 inst_cell_70_121 (.BL(BL121),.BLN(BLN121),.WL(WL70));
sram_cell_6t_5 inst_cell_70_122 (.BL(BL122),.BLN(BLN122),.WL(WL70));
sram_cell_6t_5 inst_cell_70_123 (.BL(BL123),.BLN(BLN123),.WL(WL70));
sram_cell_6t_5 inst_cell_70_124 (.BL(BL124),.BLN(BLN124),.WL(WL70));
sram_cell_6t_5 inst_cell_70_125 (.BL(BL125),.BLN(BLN125),.WL(WL70));
sram_cell_6t_5 inst_cell_70_126 (.BL(BL126),.BLN(BLN126),.WL(WL70));
sram_cell_6t_5 inst_cell_70_127 (.BL(BL127),.BLN(BLN127),.WL(WL70));
sram_cell_6t_5 inst_cell_71_0 (.BL(BL0),.BLN(BLN0),.WL(WL71));
sram_cell_6t_5 inst_cell_71_1 (.BL(BL1),.BLN(BLN1),.WL(WL71));
sram_cell_6t_5 inst_cell_71_2 (.BL(BL2),.BLN(BLN2),.WL(WL71));
sram_cell_6t_5 inst_cell_71_3 (.BL(BL3),.BLN(BLN3),.WL(WL71));
sram_cell_6t_5 inst_cell_71_4 (.BL(BL4),.BLN(BLN4),.WL(WL71));
sram_cell_6t_5 inst_cell_71_5 (.BL(BL5),.BLN(BLN5),.WL(WL71));
sram_cell_6t_5 inst_cell_71_6 (.BL(BL6),.BLN(BLN6),.WL(WL71));
sram_cell_6t_5 inst_cell_71_7 (.BL(BL7),.BLN(BLN7),.WL(WL71));
sram_cell_6t_5 inst_cell_71_8 (.BL(BL8),.BLN(BLN8),.WL(WL71));
sram_cell_6t_5 inst_cell_71_9 (.BL(BL9),.BLN(BLN9),.WL(WL71));
sram_cell_6t_5 inst_cell_71_10 (.BL(BL10),.BLN(BLN10),.WL(WL71));
sram_cell_6t_5 inst_cell_71_11 (.BL(BL11),.BLN(BLN11),.WL(WL71));
sram_cell_6t_5 inst_cell_71_12 (.BL(BL12),.BLN(BLN12),.WL(WL71));
sram_cell_6t_5 inst_cell_71_13 (.BL(BL13),.BLN(BLN13),.WL(WL71));
sram_cell_6t_5 inst_cell_71_14 (.BL(BL14),.BLN(BLN14),.WL(WL71));
sram_cell_6t_5 inst_cell_71_15 (.BL(BL15),.BLN(BLN15),.WL(WL71));
sram_cell_6t_5 inst_cell_71_16 (.BL(BL16),.BLN(BLN16),.WL(WL71));
sram_cell_6t_5 inst_cell_71_17 (.BL(BL17),.BLN(BLN17),.WL(WL71));
sram_cell_6t_5 inst_cell_71_18 (.BL(BL18),.BLN(BLN18),.WL(WL71));
sram_cell_6t_5 inst_cell_71_19 (.BL(BL19),.BLN(BLN19),.WL(WL71));
sram_cell_6t_5 inst_cell_71_20 (.BL(BL20),.BLN(BLN20),.WL(WL71));
sram_cell_6t_5 inst_cell_71_21 (.BL(BL21),.BLN(BLN21),.WL(WL71));
sram_cell_6t_5 inst_cell_71_22 (.BL(BL22),.BLN(BLN22),.WL(WL71));
sram_cell_6t_5 inst_cell_71_23 (.BL(BL23),.BLN(BLN23),.WL(WL71));
sram_cell_6t_5 inst_cell_71_24 (.BL(BL24),.BLN(BLN24),.WL(WL71));
sram_cell_6t_5 inst_cell_71_25 (.BL(BL25),.BLN(BLN25),.WL(WL71));
sram_cell_6t_5 inst_cell_71_26 (.BL(BL26),.BLN(BLN26),.WL(WL71));
sram_cell_6t_5 inst_cell_71_27 (.BL(BL27),.BLN(BLN27),.WL(WL71));
sram_cell_6t_5 inst_cell_71_28 (.BL(BL28),.BLN(BLN28),.WL(WL71));
sram_cell_6t_5 inst_cell_71_29 (.BL(BL29),.BLN(BLN29),.WL(WL71));
sram_cell_6t_5 inst_cell_71_30 (.BL(BL30),.BLN(BLN30),.WL(WL71));
sram_cell_6t_5 inst_cell_71_31 (.BL(BL31),.BLN(BLN31),.WL(WL71));
sram_cell_6t_5 inst_cell_71_32 (.BL(BL32),.BLN(BLN32),.WL(WL71));
sram_cell_6t_5 inst_cell_71_33 (.BL(BL33),.BLN(BLN33),.WL(WL71));
sram_cell_6t_5 inst_cell_71_34 (.BL(BL34),.BLN(BLN34),.WL(WL71));
sram_cell_6t_5 inst_cell_71_35 (.BL(BL35),.BLN(BLN35),.WL(WL71));
sram_cell_6t_5 inst_cell_71_36 (.BL(BL36),.BLN(BLN36),.WL(WL71));
sram_cell_6t_5 inst_cell_71_37 (.BL(BL37),.BLN(BLN37),.WL(WL71));
sram_cell_6t_5 inst_cell_71_38 (.BL(BL38),.BLN(BLN38),.WL(WL71));
sram_cell_6t_5 inst_cell_71_39 (.BL(BL39),.BLN(BLN39),.WL(WL71));
sram_cell_6t_5 inst_cell_71_40 (.BL(BL40),.BLN(BLN40),.WL(WL71));
sram_cell_6t_5 inst_cell_71_41 (.BL(BL41),.BLN(BLN41),.WL(WL71));
sram_cell_6t_5 inst_cell_71_42 (.BL(BL42),.BLN(BLN42),.WL(WL71));
sram_cell_6t_5 inst_cell_71_43 (.BL(BL43),.BLN(BLN43),.WL(WL71));
sram_cell_6t_5 inst_cell_71_44 (.BL(BL44),.BLN(BLN44),.WL(WL71));
sram_cell_6t_5 inst_cell_71_45 (.BL(BL45),.BLN(BLN45),.WL(WL71));
sram_cell_6t_5 inst_cell_71_46 (.BL(BL46),.BLN(BLN46),.WL(WL71));
sram_cell_6t_5 inst_cell_71_47 (.BL(BL47),.BLN(BLN47),.WL(WL71));
sram_cell_6t_5 inst_cell_71_48 (.BL(BL48),.BLN(BLN48),.WL(WL71));
sram_cell_6t_5 inst_cell_71_49 (.BL(BL49),.BLN(BLN49),.WL(WL71));
sram_cell_6t_5 inst_cell_71_50 (.BL(BL50),.BLN(BLN50),.WL(WL71));
sram_cell_6t_5 inst_cell_71_51 (.BL(BL51),.BLN(BLN51),.WL(WL71));
sram_cell_6t_5 inst_cell_71_52 (.BL(BL52),.BLN(BLN52),.WL(WL71));
sram_cell_6t_5 inst_cell_71_53 (.BL(BL53),.BLN(BLN53),.WL(WL71));
sram_cell_6t_5 inst_cell_71_54 (.BL(BL54),.BLN(BLN54),.WL(WL71));
sram_cell_6t_5 inst_cell_71_55 (.BL(BL55),.BLN(BLN55),.WL(WL71));
sram_cell_6t_5 inst_cell_71_56 (.BL(BL56),.BLN(BLN56),.WL(WL71));
sram_cell_6t_5 inst_cell_71_57 (.BL(BL57),.BLN(BLN57),.WL(WL71));
sram_cell_6t_5 inst_cell_71_58 (.BL(BL58),.BLN(BLN58),.WL(WL71));
sram_cell_6t_5 inst_cell_71_59 (.BL(BL59),.BLN(BLN59),.WL(WL71));
sram_cell_6t_5 inst_cell_71_60 (.BL(BL60),.BLN(BLN60),.WL(WL71));
sram_cell_6t_5 inst_cell_71_61 (.BL(BL61),.BLN(BLN61),.WL(WL71));
sram_cell_6t_5 inst_cell_71_62 (.BL(BL62),.BLN(BLN62),.WL(WL71));
sram_cell_6t_5 inst_cell_71_63 (.BL(BL63),.BLN(BLN63),.WL(WL71));
sram_cell_6t_5 inst_cell_71_64 (.BL(BL64),.BLN(BLN64),.WL(WL71));
sram_cell_6t_5 inst_cell_71_65 (.BL(BL65),.BLN(BLN65),.WL(WL71));
sram_cell_6t_5 inst_cell_71_66 (.BL(BL66),.BLN(BLN66),.WL(WL71));
sram_cell_6t_5 inst_cell_71_67 (.BL(BL67),.BLN(BLN67),.WL(WL71));
sram_cell_6t_5 inst_cell_71_68 (.BL(BL68),.BLN(BLN68),.WL(WL71));
sram_cell_6t_5 inst_cell_71_69 (.BL(BL69),.BLN(BLN69),.WL(WL71));
sram_cell_6t_5 inst_cell_71_70 (.BL(BL70),.BLN(BLN70),.WL(WL71));
sram_cell_6t_5 inst_cell_71_71 (.BL(BL71),.BLN(BLN71),.WL(WL71));
sram_cell_6t_5 inst_cell_71_72 (.BL(BL72),.BLN(BLN72),.WL(WL71));
sram_cell_6t_5 inst_cell_71_73 (.BL(BL73),.BLN(BLN73),.WL(WL71));
sram_cell_6t_5 inst_cell_71_74 (.BL(BL74),.BLN(BLN74),.WL(WL71));
sram_cell_6t_5 inst_cell_71_75 (.BL(BL75),.BLN(BLN75),.WL(WL71));
sram_cell_6t_5 inst_cell_71_76 (.BL(BL76),.BLN(BLN76),.WL(WL71));
sram_cell_6t_5 inst_cell_71_77 (.BL(BL77),.BLN(BLN77),.WL(WL71));
sram_cell_6t_5 inst_cell_71_78 (.BL(BL78),.BLN(BLN78),.WL(WL71));
sram_cell_6t_5 inst_cell_71_79 (.BL(BL79),.BLN(BLN79),.WL(WL71));
sram_cell_6t_5 inst_cell_71_80 (.BL(BL80),.BLN(BLN80),.WL(WL71));
sram_cell_6t_5 inst_cell_71_81 (.BL(BL81),.BLN(BLN81),.WL(WL71));
sram_cell_6t_5 inst_cell_71_82 (.BL(BL82),.BLN(BLN82),.WL(WL71));
sram_cell_6t_5 inst_cell_71_83 (.BL(BL83),.BLN(BLN83),.WL(WL71));
sram_cell_6t_5 inst_cell_71_84 (.BL(BL84),.BLN(BLN84),.WL(WL71));
sram_cell_6t_5 inst_cell_71_85 (.BL(BL85),.BLN(BLN85),.WL(WL71));
sram_cell_6t_5 inst_cell_71_86 (.BL(BL86),.BLN(BLN86),.WL(WL71));
sram_cell_6t_5 inst_cell_71_87 (.BL(BL87),.BLN(BLN87),.WL(WL71));
sram_cell_6t_5 inst_cell_71_88 (.BL(BL88),.BLN(BLN88),.WL(WL71));
sram_cell_6t_5 inst_cell_71_89 (.BL(BL89),.BLN(BLN89),.WL(WL71));
sram_cell_6t_5 inst_cell_71_90 (.BL(BL90),.BLN(BLN90),.WL(WL71));
sram_cell_6t_5 inst_cell_71_91 (.BL(BL91),.BLN(BLN91),.WL(WL71));
sram_cell_6t_5 inst_cell_71_92 (.BL(BL92),.BLN(BLN92),.WL(WL71));
sram_cell_6t_5 inst_cell_71_93 (.BL(BL93),.BLN(BLN93),.WL(WL71));
sram_cell_6t_5 inst_cell_71_94 (.BL(BL94),.BLN(BLN94),.WL(WL71));
sram_cell_6t_5 inst_cell_71_95 (.BL(BL95),.BLN(BLN95),.WL(WL71));
sram_cell_6t_5 inst_cell_71_96 (.BL(BL96),.BLN(BLN96),.WL(WL71));
sram_cell_6t_5 inst_cell_71_97 (.BL(BL97),.BLN(BLN97),.WL(WL71));
sram_cell_6t_5 inst_cell_71_98 (.BL(BL98),.BLN(BLN98),.WL(WL71));
sram_cell_6t_5 inst_cell_71_99 (.BL(BL99),.BLN(BLN99),.WL(WL71));
sram_cell_6t_5 inst_cell_71_100 (.BL(BL100),.BLN(BLN100),.WL(WL71));
sram_cell_6t_5 inst_cell_71_101 (.BL(BL101),.BLN(BLN101),.WL(WL71));
sram_cell_6t_5 inst_cell_71_102 (.BL(BL102),.BLN(BLN102),.WL(WL71));
sram_cell_6t_5 inst_cell_71_103 (.BL(BL103),.BLN(BLN103),.WL(WL71));
sram_cell_6t_5 inst_cell_71_104 (.BL(BL104),.BLN(BLN104),.WL(WL71));
sram_cell_6t_5 inst_cell_71_105 (.BL(BL105),.BLN(BLN105),.WL(WL71));
sram_cell_6t_5 inst_cell_71_106 (.BL(BL106),.BLN(BLN106),.WL(WL71));
sram_cell_6t_5 inst_cell_71_107 (.BL(BL107),.BLN(BLN107),.WL(WL71));
sram_cell_6t_5 inst_cell_71_108 (.BL(BL108),.BLN(BLN108),.WL(WL71));
sram_cell_6t_5 inst_cell_71_109 (.BL(BL109),.BLN(BLN109),.WL(WL71));
sram_cell_6t_5 inst_cell_71_110 (.BL(BL110),.BLN(BLN110),.WL(WL71));
sram_cell_6t_5 inst_cell_71_111 (.BL(BL111),.BLN(BLN111),.WL(WL71));
sram_cell_6t_5 inst_cell_71_112 (.BL(BL112),.BLN(BLN112),.WL(WL71));
sram_cell_6t_5 inst_cell_71_113 (.BL(BL113),.BLN(BLN113),.WL(WL71));
sram_cell_6t_5 inst_cell_71_114 (.BL(BL114),.BLN(BLN114),.WL(WL71));
sram_cell_6t_5 inst_cell_71_115 (.BL(BL115),.BLN(BLN115),.WL(WL71));
sram_cell_6t_5 inst_cell_71_116 (.BL(BL116),.BLN(BLN116),.WL(WL71));
sram_cell_6t_5 inst_cell_71_117 (.BL(BL117),.BLN(BLN117),.WL(WL71));
sram_cell_6t_5 inst_cell_71_118 (.BL(BL118),.BLN(BLN118),.WL(WL71));
sram_cell_6t_5 inst_cell_71_119 (.BL(BL119),.BLN(BLN119),.WL(WL71));
sram_cell_6t_5 inst_cell_71_120 (.BL(BL120),.BLN(BLN120),.WL(WL71));
sram_cell_6t_5 inst_cell_71_121 (.BL(BL121),.BLN(BLN121),.WL(WL71));
sram_cell_6t_5 inst_cell_71_122 (.BL(BL122),.BLN(BLN122),.WL(WL71));
sram_cell_6t_5 inst_cell_71_123 (.BL(BL123),.BLN(BLN123),.WL(WL71));
sram_cell_6t_5 inst_cell_71_124 (.BL(BL124),.BLN(BLN124),.WL(WL71));
sram_cell_6t_5 inst_cell_71_125 (.BL(BL125),.BLN(BLN125),.WL(WL71));
sram_cell_6t_5 inst_cell_71_126 (.BL(BL126),.BLN(BLN126),.WL(WL71));
sram_cell_6t_5 inst_cell_71_127 (.BL(BL127),.BLN(BLN127),.WL(WL71));
sram_cell_6t_5 inst_cell_72_0 (.BL(BL0),.BLN(BLN0),.WL(WL72));
sram_cell_6t_5 inst_cell_72_1 (.BL(BL1),.BLN(BLN1),.WL(WL72));
sram_cell_6t_5 inst_cell_72_2 (.BL(BL2),.BLN(BLN2),.WL(WL72));
sram_cell_6t_5 inst_cell_72_3 (.BL(BL3),.BLN(BLN3),.WL(WL72));
sram_cell_6t_5 inst_cell_72_4 (.BL(BL4),.BLN(BLN4),.WL(WL72));
sram_cell_6t_5 inst_cell_72_5 (.BL(BL5),.BLN(BLN5),.WL(WL72));
sram_cell_6t_5 inst_cell_72_6 (.BL(BL6),.BLN(BLN6),.WL(WL72));
sram_cell_6t_5 inst_cell_72_7 (.BL(BL7),.BLN(BLN7),.WL(WL72));
sram_cell_6t_5 inst_cell_72_8 (.BL(BL8),.BLN(BLN8),.WL(WL72));
sram_cell_6t_5 inst_cell_72_9 (.BL(BL9),.BLN(BLN9),.WL(WL72));
sram_cell_6t_5 inst_cell_72_10 (.BL(BL10),.BLN(BLN10),.WL(WL72));
sram_cell_6t_5 inst_cell_72_11 (.BL(BL11),.BLN(BLN11),.WL(WL72));
sram_cell_6t_5 inst_cell_72_12 (.BL(BL12),.BLN(BLN12),.WL(WL72));
sram_cell_6t_5 inst_cell_72_13 (.BL(BL13),.BLN(BLN13),.WL(WL72));
sram_cell_6t_5 inst_cell_72_14 (.BL(BL14),.BLN(BLN14),.WL(WL72));
sram_cell_6t_5 inst_cell_72_15 (.BL(BL15),.BLN(BLN15),.WL(WL72));
sram_cell_6t_5 inst_cell_72_16 (.BL(BL16),.BLN(BLN16),.WL(WL72));
sram_cell_6t_5 inst_cell_72_17 (.BL(BL17),.BLN(BLN17),.WL(WL72));
sram_cell_6t_5 inst_cell_72_18 (.BL(BL18),.BLN(BLN18),.WL(WL72));
sram_cell_6t_5 inst_cell_72_19 (.BL(BL19),.BLN(BLN19),.WL(WL72));
sram_cell_6t_5 inst_cell_72_20 (.BL(BL20),.BLN(BLN20),.WL(WL72));
sram_cell_6t_5 inst_cell_72_21 (.BL(BL21),.BLN(BLN21),.WL(WL72));
sram_cell_6t_5 inst_cell_72_22 (.BL(BL22),.BLN(BLN22),.WL(WL72));
sram_cell_6t_5 inst_cell_72_23 (.BL(BL23),.BLN(BLN23),.WL(WL72));
sram_cell_6t_5 inst_cell_72_24 (.BL(BL24),.BLN(BLN24),.WL(WL72));
sram_cell_6t_5 inst_cell_72_25 (.BL(BL25),.BLN(BLN25),.WL(WL72));
sram_cell_6t_5 inst_cell_72_26 (.BL(BL26),.BLN(BLN26),.WL(WL72));
sram_cell_6t_5 inst_cell_72_27 (.BL(BL27),.BLN(BLN27),.WL(WL72));
sram_cell_6t_5 inst_cell_72_28 (.BL(BL28),.BLN(BLN28),.WL(WL72));
sram_cell_6t_5 inst_cell_72_29 (.BL(BL29),.BLN(BLN29),.WL(WL72));
sram_cell_6t_5 inst_cell_72_30 (.BL(BL30),.BLN(BLN30),.WL(WL72));
sram_cell_6t_5 inst_cell_72_31 (.BL(BL31),.BLN(BLN31),.WL(WL72));
sram_cell_6t_5 inst_cell_72_32 (.BL(BL32),.BLN(BLN32),.WL(WL72));
sram_cell_6t_5 inst_cell_72_33 (.BL(BL33),.BLN(BLN33),.WL(WL72));
sram_cell_6t_5 inst_cell_72_34 (.BL(BL34),.BLN(BLN34),.WL(WL72));
sram_cell_6t_5 inst_cell_72_35 (.BL(BL35),.BLN(BLN35),.WL(WL72));
sram_cell_6t_5 inst_cell_72_36 (.BL(BL36),.BLN(BLN36),.WL(WL72));
sram_cell_6t_5 inst_cell_72_37 (.BL(BL37),.BLN(BLN37),.WL(WL72));
sram_cell_6t_5 inst_cell_72_38 (.BL(BL38),.BLN(BLN38),.WL(WL72));
sram_cell_6t_5 inst_cell_72_39 (.BL(BL39),.BLN(BLN39),.WL(WL72));
sram_cell_6t_5 inst_cell_72_40 (.BL(BL40),.BLN(BLN40),.WL(WL72));
sram_cell_6t_5 inst_cell_72_41 (.BL(BL41),.BLN(BLN41),.WL(WL72));
sram_cell_6t_5 inst_cell_72_42 (.BL(BL42),.BLN(BLN42),.WL(WL72));
sram_cell_6t_5 inst_cell_72_43 (.BL(BL43),.BLN(BLN43),.WL(WL72));
sram_cell_6t_5 inst_cell_72_44 (.BL(BL44),.BLN(BLN44),.WL(WL72));
sram_cell_6t_5 inst_cell_72_45 (.BL(BL45),.BLN(BLN45),.WL(WL72));
sram_cell_6t_5 inst_cell_72_46 (.BL(BL46),.BLN(BLN46),.WL(WL72));
sram_cell_6t_5 inst_cell_72_47 (.BL(BL47),.BLN(BLN47),.WL(WL72));
sram_cell_6t_5 inst_cell_72_48 (.BL(BL48),.BLN(BLN48),.WL(WL72));
sram_cell_6t_5 inst_cell_72_49 (.BL(BL49),.BLN(BLN49),.WL(WL72));
sram_cell_6t_5 inst_cell_72_50 (.BL(BL50),.BLN(BLN50),.WL(WL72));
sram_cell_6t_5 inst_cell_72_51 (.BL(BL51),.BLN(BLN51),.WL(WL72));
sram_cell_6t_5 inst_cell_72_52 (.BL(BL52),.BLN(BLN52),.WL(WL72));
sram_cell_6t_5 inst_cell_72_53 (.BL(BL53),.BLN(BLN53),.WL(WL72));
sram_cell_6t_5 inst_cell_72_54 (.BL(BL54),.BLN(BLN54),.WL(WL72));
sram_cell_6t_5 inst_cell_72_55 (.BL(BL55),.BLN(BLN55),.WL(WL72));
sram_cell_6t_5 inst_cell_72_56 (.BL(BL56),.BLN(BLN56),.WL(WL72));
sram_cell_6t_5 inst_cell_72_57 (.BL(BL57),.BLN(BLN57),.WL(WL72));
sram_cell_6t_5 inst_cell_72_58 (.BL(BL58),.BLN(BLN58),.WL(WL72));
sram_cell_6t_5 inst_cell_72_59 (.BL(BL59),.BLN(BLN59),.WL(WL72));
sram_cell_6t_5 inst_cell_72_60 (.BL(BL60),.BLN(BLN60),.WL(WL72));
sram_cell_6t_5 inst_cell_72_61 (.BL(BL61),.BLN(BLN61),.WL(WL72));
sram_cell_6t_5 inst_cell_72_62 (.BL(BL62),.BLN(BLN62),.WL(WL72));
sram_cell_6t_5 inst_cell_72_63 (.BL(BL63),.BLN(BLN63),.WL(WL72));
sram_cell_6t_5 inst_cell_72_64 (.BL(BL64),.BLN(BLN64),.WL(WL72));
sram_cell_6t_5 inst_cell_72_65 (.BL(BL65),.BLN(BLN65),.WL(WL72));
sram_cell_6t_5 inst_cell_72_66 (.BL(BL66),.BLN(BLN66),.WL(WL72));
sram_cell_6t_5 inst_cell_72_67 (.BL(BL67),.BLN(BLN67),.WL(WL72));
sram_cell_6t_5 inst_cell_72_68 (.BL(BL68),.BLN(BLN68),.WL(WL72));
sram_cell_6t_5 inst_cell_72_69 (.BL(BL69),.BLN(BLN69),.WL(WL72));
sram_cell_6t_5 inst_cell_72_70 (.BL(BL70),.BLN(BLN70),.WL(WL72));
sram_cell_6t_5 inst_cell_72_71 (.BL(BL71),.BLN(BLN71),.WL(WL72));
sram_cell_6t_5 inst_cell_72_72 (.BL(BL72),.BLN(BLN72),.WL(WL72));
sram_cell_6t_5 inst_cell_72_73 (.BL(BL73),.BLN(BLN73),.WL(WL72));
sram_cell_6t_5 inst_cell_72_74 (.BL(BL74),.BLN(BLN74),.WL(WL72));
sram_cell_6t_5 inst_cell_72_75 (.BL(BL75),.BLN(BLN75),.WL(WL72));
sram_cell_6t_5 inst_cell_72_76 (.BL(BL76),.BLN(BLN76),.WL(WL72));
sram_cell_6t_5 inst_cell_72_77 (.BL(BL77),.BLN(BLN77),.WL(WL72));
sram_cell_6t_5 inst_cell_72_78 (.BL(BL78),.BLN(BLN78),.WL(WL72));
sram_cell_6t_5 inst_cell_72_79 (.BL(BL79),.BLN(BLN79),.WL(WL72));
sram_cell_6t_5 inst_cell_72_80 (.BL(BL80),.BLN(BLN80),.WL(WL72));
sram_cell_6t_5 inst_cell_72_81 (.BL(BL81),.BLN(BLN81),.WL(WL72));
sram_cell_6t_5 inst_cell_72_82 (.BL(BL82),.BLN(BLN82),.WL(WL72));
sram_cell_6t_5 inst_cell_72_83 (.BL(BL83),.BLN(BLN83),.WL(WL72));
sram_cell_6t_5 inst_cell_72_84 (.BL(BL84),.BLN(BLN84),.WL(WL72));
sram_cell_6t_5 inst_cell_72_85 (.BL(BL85),.BLN(BLN85),.WL(WL72));
sram_cell_6t_5 inst_cell_72_86 (.BL(BL86),.BLN(BLN86),.WL(WL72));
sram_cell_6t_5 inst_cell_72_87 (.BL(BL87),.BLN(BLN87),.WL(WL72));
sram_cell_6t_5 inst_cell_72_88 (.BL(BL88),.BLN(BLN88),.WL(WL72));
sram_cell_6t_5 inst_cell_72_89 (.BL(BL89),.BLN(BLN89),.WL(WL72));
sram_cell_6t_5 inst_cell_72_90 (.BL(BL90),.BLN(BLN90),.WL(WL72));
sram_cell_6t_5 inst_cell_72_91 (.BL(BL91),.BLN(BLN91),.WL(WL72));
sram_cell_6t_5 inst_cell_72_92 (.BL(BL92),.BLN(BLN92),.WL(WL72));
sram_cell_6t_5 inst_cell_72_93 (.BL(BL93),.BLN(BLN93),.WL(WL72));
sram_cell_6t_5 inst_cell_72_94 (.BL(BL94),.BLN(BLN94),.WL(WL72));
sram_cell_6t_5 inst_cell_72_95 (.BL(BL95),.BLN(BLN95),.WL(WL72));
sram_cell_6t_5 inst_cell_72_96 (.BL(BL96),.BLN(BLN96),.WL(WL72));
sram_cell_6t_5 inst_cell_72_97 (.BL(BL97),.BLN(BLN97),.WL(WL72));
sram_cell_6t_5 inst_cell_72_98 (.BL(BL98),.BLN(BLN98),.WL(WL72));
sram_cell_6t_5 inst_cell_72_99 (.BL(BL99),.BLN(BLN99),.WL(WL72));
sram_cell_6t_5 inst_cell_72_100 (.BL(BL100),.BLN(BLN100),.WL(WL72));
sram_cell_6t_5 inst_cell_72_101 (.BL(BL101),.BLN(BLN101),.WL(WL72));
sram_cell_6t_5 inst_cell_72_102 (.BL(BL102),.BLN(BLN102),.WL(WL72));
sram_cell_6t_5 inst_cell_72_103 (.BL(BL103),.BLN(BLN103),.WL(WL72));
sram_cell_6t_5 inst_cell_72_104 (.BL(BL104),.BLN(BLN104),.WL(WL72));
sram_cell_6t_5 inst_cell_72_105 (.BL(BL105),.BLN(BLN105),.WL(WL72));
sram_cell_6t_5 inst_cell_72_106 (.BL(BL106),.BLN(BLN106),.WL(WL72));
sram_cell_6t_5 inst_cell_72_107 (.BL(BL107),.BLN(BLN107),.WL(WL72));
sram_cell_6t_5 inst_cell_72_108 (.BL(BL108),.BLN(BLN108),.WL(WL72));
sram_cell_6t_5 inst_cell_72_109 (.BL(BL109),.BLN(BLN109),.WL(WL72));
sram_cell_6t_5 inst_cell_72_110 (.BL(BL110),.BLN(BLN110),.WL(WL72));
sram_cell_6t_5 inst_cell_72_111 (.BL(BL111),.BLN(BLN111),.WL(WL72));
sram_cell_6t_5 inst_cell_72_112 (.BL(BL112),.BLN(BLN112),.WL(WL72));
sram_cell_6t_5 inst_cell_72_113 (.BL(BL113),.BLN(BLN113),.WL(WL72));
sram_cell_6t_5 inst_cell_72_114 (.BL(BL114),.BLN(BLN114),.WL(WL72));
sram_cell_6t_5 inst_cell_72_115 (.BL(BL115),.BLN(BLN115),.WL(WL72));
sram_cell_6t_5 inst_cell_72_116 (.BL(BL116),.BLN(BLN116),.WL(WL72));
sram_cell_6t_5 inst_cell_72_117 (.BL(BL117),.BLN(BLN117),.WL(WL72));
sram_cell_6t_5 inst_cell_72_118 (.BL(BL118),.BLN(BLN118),.WL(WL72));
sram_cell_6t_5 inst_cell_72_119 (.BL(BL119),.BLN(BLN119),.WL(WL72));
sram_cell_6t_5 inst_cell_72_120 (.BL(BL120),.BLN(BLN120),.WL(WL72));
sram_cell_6t_5 inst_cell_72_121 (.BL(BL121),.BLN(BLN121),.WL(WL72));
sram_cell_6t_5 inst_cell_72_122 (.BL(BL122),.BLN(BLN122),.WL(WL72));
sram_cell_6t_5 inst_cell_72_123 (.BL(BL123),.BLN(BLN123),.WL(WL72));
sram_cell_6t_5 inst_cell_72_124 (.BL(BL124),.BLN(BLN124),.WL(WL72));
sram_cell_6t_5 inst_cell_72_125 (.BL(BL125),.BLN(BLN125),.WL(WL72));
sram_cell_6t_5 inst_cell_72_126 (.BL(BL126),.BLN(BLN126),.WL(WL72));
sram_cell_6t_5 inst_cell_72_127 (.BL(BL127),.BLN(BLN127),.WL(WL72));
sram_cell_6t_5 inst_cell_73_0 (.BL(BL0),.BLN(BLN0),.WL(WL73));
sram_cell_6t_5 inst_cell_73_1 (.BL(BL1),.BLN(BLN1),.WL(WL73));
sram_cell_6t_5 inst_cell_73_2 (.BL(BL2),.BLN(BLN2),.WL(WL73));
sram_cell_6t_5 inst_cell_73_3 (.BL(BL3),.BLN(BLN3),.WL(WL73));
sram_cell_6t_5 inst_cell_73_4 (.BL(BL4),.BLN(BLN4),.WL(WL73));
sram_cell_6t_5 inst_cell_73_5 (.BL(BL5),.BLN(BLN5),.WL(WL73));
sram_cell_6t_5 inst_cell_73_6 (.BL(BL6),.BLN(BLN6),.WL(WL73));
sram_cell_6t_5 inst_cell_73_7 (.BL(BL7),.BLN(BLN7),.WL(WL73));
sram_cell_6t_5 inst_cell_73_8 (.BL(BL8),.BLN(BLN8),.WL(WL73));
sram_cell_6t_5 inst_cell_73_9 (.BL(BL9),.BLN(BLN9),.WL(WL73));
sram_cell_6t_5 inst_cell_73_10 (.BL(BL10),.BLN(BLN10),.WL(WL73));
sram_cell_6t_5 inst_cell_73_11 (.BL(BL11),.BLN(BLN11),.WL(WL73));
sram_cell_6t_5 inst_cell_73_12 (.BL(BL12),.BLN(BLN12),.WL(WL73));
sram_cell_6t_5 inst_cell_73_13 (.BL(BL13),.BLN(BLN13),.WL(WL73));
sram_cell_6t_5 inst_cell_73_14 (.BL(BL14),.BLN(BLN14),.WL(WL73));
sram_cell_6t_5 inst_cell_73_15 (.BL(BL15),.BLN(BLN15),.WL(WL73));
sram_cell_6t_5 inst_cell_73_16 (.BL(BL16),.BLN(BLN16),.WL(WL73));
sram_cell_6t_5 inst_cell_73_17 (.BL(BL17),.BLN(BLN17),.WL(WL73));
sram_cell_6t_5 inst_cell_73_18 (.BL(BL18),.BLN(BLN18),.WL(WL73));
sram_cell_6t_5 inst_cell_73_19 (.BL(BL19),.BLN(BLN19),.WL(WL73));
sram_cell_6t_5 inst_cell_73_20 (.BL(BL20),.BLN(BLN20),.WL(WL73));
sram_cell_6t_5 inst_cell_73_21 (.BL(BL21),.BLN(BLN21),.WL(WL73));
sram_cell_6t_5 inst_cell_73_22 (.BL(BL22),.BLN(BLN22),.WL(WL73));
sram_cell_6t_5 inst_cell_73_23 (.BL(BL23),.BLN(BLN23),.WL(WL73));
sram_cell_6t_5 inst_cell_73_24 (.BL(BL24),.BLN(BLN24),.WL(WL73));
sram_cell_6t_5 inst_cell_73_25 (.BL(BL25),.BLN(BLN25),.WL(WL73));
sram_cell_6t_5 inst_cell_73_26 (.BL(BL26),.BLN(BLN26),.WL(WL73));
sram_cell_6t_5 inst_cell_73_27 (.BL(BL27),.BLN(BLN27),.WL(WL73));
sram_cell_6t_5 inst_cell_73_28 (.BL(BL28),.BLN(BLN28),.WL(WL73));
sram_cell_6t_5 inst_cell_73_29 (.BL(BL29),.BLN(BLN29),.WL(WL73));
sram_cell_6t_5 inst_cell_73_30 (.BL(BL30),.BLN(BLN30),.WL(WL73));
sram_cell_6t_5 inst_cell_73_31 (.BL(BL31),.BLN(BLN31),.WL(WL73));
sram_cell_6t_5 inst_cell_73_32 (.BL(BL32),.BLN(BLN32),.WL(WL73));
sram_cell_6t_5 inst_cell_73_33 (.BL(BL33),.BLN(BLN33),.WL(WL73));
sram_cell_6t_5 inst_cell_73_34 (.BL(BL34),.BLN(BLN34),.WL(WL73));
sram_cell_6t_5 inst_cell_73_35 (.BL(BL35),.BLN(BLN35),.WL(WL73));
sram_cell_6t_5 inst_cell_73_36 (.BL(BL36),.BLN(BLN36),.WL(WL73));
sram_cell_6t_5 inst_cell_73_37 (.BL(BL37),.BLN(BLN37),.WL(WL73));
sram_cell_6t_5 inst_cell_73_38 (.BL(BL38),.BLN(BLN38),.WL(WL73));
sram_cell_6t_5 inst_cell_73_39 (.BL(BL39),.BLN(BLN39),.WL(WL73));
sram_cell_6t_5 inst_cell_73_40 (.BL(BL40),.BLN(BLN40),.WL(WL73));
sram_cell_6t_5 inst_cell_73_41 (.BL(BL41),.BLN(BLN41),.WL(WL73));
sram_cell_6t_5 inst_cell_73_42 (.BL(BL42),.BLN(BLN42),.WL(WL73));
sram_cell_6t_5 inst_cell_73_43 (.BL(BL43),.BLN(BLN43),.WL(WL73));
sram_cell_6t_5 inst_cell_73_44 (.BL(BL44),.BLN(BLN44),.WL(WL73));
sram_cell_6t_5 inst_cell_73_45 (.BL(BL45),.BLN(BLN45),.WL(WL73));
sram_cell_6t_5 inst_cell_73_46 (.BL(BL46),.BLN(BLN46),.WL(WL73));
sram_cell_6t_5 inst_cell_73_47 (.BL(BL47),.BLN(BLN47),.WL(WL73));
sram_cell_6t_5 inst_cell_73_48 (.BL(BL48),.BLN(BLN48),.WL(WL73));
sram_cell_6t_5 inst_cell_73_49 (.BL(BL49),.BLN(BLN49),.WL(WL73));
sram_cell_6t_5 inst_cell_73_50 (.BL(BL50),.BLN(BLN50),.WL(WL73));
sram_cell_6t_5 inst_cell_73_51 (.BL(BL51),.BLN(BLN51),.WL(WL73));
sram_cell_6t_5 inst_cell_73_52 (.BL(BL52),.BLN(BLN52),.WL(WL73));
sram_cell_6t_5 inst_cell_73_53 (.BL(BL53),.BLN(BLN53),.WL(WL73));
sram_cell_6t_5 inst_cell_73_54 (.BL(BL54),.BLN(BLN54),.WL(WL73));
sram_cell_6t_5 inst_cell_73_55 (.BL(BL55),.BLN(BLN55),.WL(WL73));
sram_cell_6t_5 inst_cell_73_56 (.BL(BL56),.BLN(BLN56),.WL(WL73));
sram_cell_6t_5 inst_cell_73_57 (.BL(BL57),.BLN(BLN57),.WL(WL73));
sram_cell_6t_5 inst_cell_73_58 (.BL(BL58),.BLN(BLN58),.WL(WL73));
sram_cell_6t_5 inst_cell_73_59 (.BL(BL59),.BLN(BLN59),.WL(WL73));
sram_cell_6t_5 inst_cell_73_60 (.BL(BL60),.BLN(BLN60),.WL(WL73));
sram_cell_6t_5 inst_cell_73_61 (.BL(BL61),.BLN(BLN61),.WL(WL73));
sram_cell_6t_5 inst_cell_73_62 (.BL(BL62),.BLN(BLN62),.WL(WL73));
sram_cell_6t_5 inst_cell_73_63 (.BL(BL63),.BLN(BLN63),.WL(WL73));
sram_cell_6t_5 inst_cell_73_64 (.BL(BL64),.BLN(BLN64),.WL(WL73));
sram_cell_6t_5 inst_cell_73_65 (.BL(BL65),.BLN(BLN65),.WL(WL73));
sram_cell_6t_5 inst_cell_73_66 (.BL(BL66),.BLN(BLN66),.WL(WL73));
sram_cell_6t_5 inst_cell_73_67 (.BL(BL67),.BLN(BLN67),.WL(WL73));
sram_cell_6t_5 inst_cell_73_68 (.BL(BL68),.BLN(BLN68),.WL(WL73));
sram_cell_6t_5 inst_cell_73_69 (.BL(BL69),.BLN(BLN69),.WL(WL73));
sram_cell_6t_5 inst_cell_73_70 (.BL(BL70),.BLN(BLN70),.WL(WL73));
sram_cell_6t_5 inst_cell_73_71 (.BL(BL71),.BLN(BLN71),.WL(WL73));
sram_cell_6t_5 inst_cell_73_72 (.BL(BL72),.BLN(BLN72),.WL(WL73));
sram_cell_6t_5 inst_cell_73_73 (.BL(BL73),.BLN(BLN73),.WL(WL73));
sram_cell_6t_5 inst_cell_73_74 (.BL(BL74),.BLN(BLN74),.WL(WL73));
sram_cell_6t_5 inst_cell_73_75 (.BL(BL75),.BLN(BLN75),.WL(WL73));
sram_cell_6t_5 inst_cell_73_76 (.BL(BL76),.BLN(BLN76),.WL(WL73));
sram_cell_6t_5 inst_cell_73_77 (.BL(BL77),.BLN(BLN77),.WL(WL73));
sram_cell_6t_5 inst_cell_73_78 (.BL(BL78),.BLN(BLN78),.WL(WL73));
sram_cell_6t_5 inst_cell_73_79 (.BL(BL79),.BLN(BLN79),.WL(WL73));
sram_cell_6t_5 inst_cell_73_80 (.BL(BL80),.BLN(BLN80),.WL(WL73));
sram_cell_6t_5 inst_cell_73_81 (.BL(BL81),.BLN(BLN81),.WL(WL73));
sram_cell_6t_5 inst_cell_73_82 (.BL(BL82),.BLN(BLN82),.WL(WL73));
sram_cell_6t_5 inst_cell_73_83 (.BL(BL83),.BLN(BLN83),.WL(WL73));
sram_cell_6t_5 inst_cell_73_84 (.BL(BL84),.BLN(BLN84),.WL(WL73));
sram_cell_6t_5 inst_cell_73_85 (.BL(BL85),.BLN(BLN85),.WL(WL73));
sram_cell_6t_5 inst_cell_73_86 (.BL(BL86),.BLN(BLN86),.WL(WL73));
sram_cell_6t_5 inst_cell_73_87 (.BL(BL87),.BLN(BLN87),.WL(WL73));
sram_cell_6t_5 inst_cell_73_88 (.BL(BL88),.BLN(BLN88),.WL(WL73));
sram_cell_6t_5 inst_cell_73_89 (.BL(BL89),.BLN(BLN89),.WL(WL73));
sram_cell_6t_5 inst_cell_73_90 (.BL(BL90),.BLN(BLN90),.WL(WL73));
sram_cell_6t_5 inst_cell_73_91 (.BL(BL91),.BLN(BLN91),.WL(WL73));
sram_cell_6t_5 inst_cell_73_92 (.BL(BL92),.BLN(BLN92),.WL(WL73));
sram_cell_6t_5 inst_cell_73_93 (.BL(BL93),.BLN(BLN93),.WL(WL73));
sram_cell_6t_5 inst_cell_73_94 (.BL(BL94),.BLN(BLN94),.WL(WL73));
sram_cell_6t_5 inst_cell_73_95 (.BL(BL95),.BLN(BLN95),.WL(WL73));
sram_cell_6t_5 inst_cell_73_96 (.BL(BL96),.BLN(BLN96),.WL(WL73));
sram_cell_6t_5 inst_cell_73_97 (.BL(BL97),.BLN(BLN97),.WL(WL73));
sram_cell_6t_5 inst_cell_73_98 (.BL(BL98),.BLN(BLN98),.WL(WL73));
sram_cell_6t_5 inst_cell_73_99 (.BL(BL99),.BLN(BLN99),.WL(WL73));
sram_cell_6t_5 inst_cell_73_100 (.BL(BL100),.BLN(BLN100),.WL(WL73));
sram_cell_6t_5 inst_cell_73_101 (.BL(BL101),.BLN(BLN101),.WL(WL73));
sram_cell_6t_5 inst_cell_73_102 (.BL(BL102),.BLN(BLN102),.WL(WL73));
sram_cell_6t_5 inst_cell_73_103 (.BL(BL103),.BLN(BLN103),.WL(WL73));
sram_cell_6t_5 inst_cell_73_104 (.BL(BL104),.BLN(BLN104),.WL(WL73));
sram_cell_6t_5 inst_cell_73_105 (.BL(BL105),.BLN(BLN105),.WL(WL73));
sram_cell_6t_5 inst_cell_73_106 (.BL(BL106),.BLN(BLN106),.WL(WL73));
sram_cell_6t_5 inst_cell_73_107 (.BL(BL107),.BLN(BLN107),.WL(WL73));
sram_cell_6t_5 inst_cell_73_108 (.BL(BL108),.BLN(BLN108),.WL(WL73));
sram_cell_6t_5 inst_cell_73_109 (.BL(BL109),.BLN(BLN109),.WL(WL73));
sram_cell_6t_5 inst_cell_73_110 (.BL(BL110),.BLN(BLN110),.WL(WL73));
sram_cell_6t_5 inst_cell_73_111 (.BL(BL111),.BLN(BLN111),.WL(WL73));
sram_cell_6t_5 inst_cell_73_112 (.BL(BL112),.BLN(BLN112),.WL(WL73));
sram_cell_6t_5 inst_cell_73_113 (.BL(BL113),.BLN(BLN113),.WL(WL73));
sram_cell_6t_5 inst_cell_73_114 (.BL(BL114),.BLN(BLN114),.WL(WL73));
sram_cell_6t_5 inst_cell_73_115 (.BL(BL115),.BLN(BLN115),.WL(WL73));
sram_cell_6t_5 inst_cell_73_116 (.BL(BL116),.BLN(BLN116),.WL(WL73));
sram_cell_6t_5 inst_cell_73_117 (.BL(BL117),.BLN(BLN117),.WL(WL73));
sram_cell_6t_5 inst_cell_73_118 (.BL(BL118),.BLN(BLN118),.WL(WL73));
sram_cell_6t_5 inst_cell_73_119 (.BL(BL119),.BLN(BLN119),.WL(WL73));
sram_cell_6t_5 inst_cell_73_120 (.BL(BL120),.BLN(BLN120),.WL(WL73));
sram_cell_6t_5 inst_cell_73_121 (.BL(BL121),.BLN(BLN121),.WL(WL73));
sram_cell_6t_5 inst_cell_73_122 (.BL(BL122),.BLN(BLN122),.WL(WL73));
sram_cell_6t_5 inst_cell_73_123 (.BL(BL123),.BLN(BLN123),.WL(WL73));
sram_cell_6t_5 inst_cell_73_124 (.BL(BL124),.BLN(BLN124),.WL(WL73));
sram_cell_6t_5 inst_cell_73_125 (.BL(BL125),.BLN(BLN125),.WL(WL73));
sram_cell_6t_5 inst_cell_73_126 (.BL(BL126),.BLN(BLN126),.WL(WL73));
sram_cell_6t_5 inst_cell_73_127 (.BL(BL127),.BLN(BLN127),.WL(WL73));
sram_cell_6t_5 inst_cell_74_0 (.BL(BL0),.BLN(BLN0),.WL(WL74));
sram_cell_6t_5 inst_cell_74_1 (.BL(BL1),.BLN(BLN1),.WL(WL74));
sram_cell_6t_5 inst_cell_74_2 (.BL(BL2),.BLN(BLN2),.WL(WL74));
sram_cell_6t_5 inst_cell_74_3 (.BL(BL3),.BLN(BLN3),.WL(WL74));
sram_cell_6t_5 inst_cell_74_4 (.BL(BL4),.BLN(BLN4),.WL(WL74));
sram_cell_6t_5 inst_cell_74_5 (.BL(BL5),.BLN(BLN5),.WL(WL74));
sram_cell_6t_5 inst_cell_74_6 (.BL(BL6),.BLN(BLN6),.WL(WL74));
sram_cell_6t_5 inst_cell_74_7 (.BL(BL7),.BLN(BLN7),.WL(WL74));
sram_cell_6t_5 inst_cell_74_8 (.BL(BL8),.BLN(BLN8),.WL(WL74));
sram_cell_6t_5 inst_cell_74_9 (.BL(BL9),.BLN(BLN9),.WL(WL74));
sram_cell_6t_5 inst_cell_74_10 (.BL(BL10),.BLN(BLN10),.WL(WL74));
sram_cell_6t_5 inst_cell_74_11 (.BL(BL11),.BLN(BLN11),.WL(WL74));
sram_cell_6t_5 inst_cell_74_12 (.BL(BL12),.BLN(BLN12),.WL(WL74));
sram_cell_6t_5 inst_cell_74_13 (.BL(BL13),.BLN(BLN13),.WL(WL74));
sram_cell_6t_5 inst_cell_74_14 (.BL(BL14),.BLN(BLN14),.WL(WL74));
sram_cell_6t_5 inst_cell_74_15 (.BL(BL15),.BLN(BLN15),.WL(WL74));
sram_cell_6t_5 inst_cell_74_16 (.BL(BL16),.BLN(BLN16),.WL(WL74));
sram_cell_6t_5 inst_cell_74_17 (.BL(BL17),.BLN(BLN17),.WL(WL74));
sram_cell_6t_5 inst_cell_74_18 (.BL(BL18),.BLN(BLN18),.WL(WL74));
sram_cell_6t_5 inst_cell_74_19 (.BL(BL19),.BLN(BLN19),.WL(WL74));
sram_cell_6t_5 inst_cell_74_20 (.BL(BL20),.BLN(BLN20),.WL(WL74));
sram_cell_6t_5 inst_cell_74_21 (.BL(BL21),.BLN(BLN21),.WL(WL74));
sram_cell_6t_5 inst_cell_74_22 (.BL(BL22),.BLN(BLN22),.WL(WL74));
sram_cell_6t_5 inst_cell_74_23 (.BL(BL23),.BLN(BLN23),.WL(WL74));
sram_cell_6t_5 inst_cell_74_24 (.BL(BL24),.BLN(BLN24),.WL(WL74));
sram_cell_6t_5 inst_cell_74_25 (.BL(BL25),.BLN(BLN25),.WL(WL74));
sram_cell_6t_5 inst_cell_74_26 (.BL(BL26),.BLN(BLN26),.WL(WL74));
sram_cell_6t_5 inst_cell_74_27 (.BL(BL27),.BLN(BLN27),.WL(WL74));
sram_cell_6t_5 inst_cell_74_28 (.BL(BL28),.BLN(BLN28),.WL(WL74));
sram_cell_6t_5 inst_cell_74_29 (.BL(BL29),.BLN(BLN29),.WL(WL74));
sram_cell_6t_5 inst_cell_74_30 (.BL(BL30),.BLN(BLN30),.WL(WL74));
sram_cell_6t_5 inst_cell_74_31 (.BL(BL31),.BLN(BLN31),.WL(WL74));
sram_cell_6t_5 inst_cell_74_32 (.BL(BL32),.BLN(BLN32),.WL(WL74));
sram_cell_6t_5 inst_cell_74_33 (.BL(BL33),.BLN(BLN33),.WL(WL74));
sram_cell_6t_5 inst_cell_74_34 (.BL(BL34),.BLN(BLN34),.WL(WL74));
sram_cell_6t_5 inst_cell_74_35 (.BL(BL35),.BLN(BLN35),.WL(WL74));
sram_cell_6t_5 inst_cell_74_36 (.BL(BL36),.BLN(BLN36),.WL(WL74));
sram_cell_6t_5 inst_cell_74_37 (.BL(BL37),.BLN(BLN37),.WL(WL74));
sram_cell_6t_5 inst_cell_74_38 (.BL(BL38),.BLN(BLN38),.WL(WL74));
sram_cell_6t_5 inst_cell_74_39 (.BL(BL39),.BLN(BLN39),.WL(WL74));
sram_cell_6t_5 inst_cell_74_40 (.BL(BL40),.BLN(BLN40),.WL(WL74));
sram_cell_6t_5 inst_cell_74_41 (.BL(BL41),.BLN(BLN41),.WL(WL74));
sram_cell_6t_5 inst_cell_74_42 (.BL(BL42),.BLN(BLN42),.WL(WL74));
sram_cell_6t_5 inst_cell_74_43 (.BL(BL43),.BLN(BLN43),.WL(WL74));
sram_cell_6t_5 inst_cell_74_44 (.BL(BL44),.BLN(BLN44),.WL(WL74));
sram_cell_6t_5 inst_cell_74_45 (.BL(BL45),.BLN(BLN45),.WL(WL74));
sram_cell_6t_5 inst_cell_74_46 (.BL(BL46),.BLN(BLN46),.WL(WL74));
sram_cell_6t_5 inst_cell_74_47 (.BL(BL47),.BLN(BLN47),.WL(WL74));
sram_cell_6t_5 inst_cell_74_48 (.BL(BL48),.BLN(BLN48),.WL(WL74));
sram_cell_6t_5 inst_cell_74_49 (.BL(BL49),.BLN(BLN49),.WL(WL74));
sram_cell_6t_5 inst_cell_74_50 (.BL(BL50),.BLN(BLN50),.WL(WL74));
sram_cell_6t_5 inst_cell_74_51 (.BL(BL51),.BLN(BLN51),.WL(WL74));
sram_cell_6t_5 inst_cell_74_52 (.BL(BL52),.BLN(BLN52),.WL(WL74));
sram_cell_6t_5 inst_cell_74_53 (.BL(BL53),.BLN(BLN53),.WL(WL74));
sram_cell_6t_5 inst_cell_74_54 (.BL(BL54),.BLN(BLN54),.WL(WL74));
sram_cell_6t_5 inst_cell_74_55 (.BL(BL55),.BLN(BLN55),.WL(WL74));
sram_cell_6t_5 inst_cell_74_56 (.BL(BL56),.BLN(BLN56),.WL(WL74));
sram_cell_6t_5 inst_cell_74_57 (.BL(BL57),.BLN(BLN57),.WL(WL74));
sram_cell_6t_5 inst_cell_74_58 (.BL(BL58),.BLN(BLN58),.WL(WL74));
sram_cell_6t_5 inst_cell_74_59 (.BL(BL59),.BLN(BLN59),.WL(WL74));
sram_cell_6t_5 inst_cell_74_60 (.BL(BL60),.BLN(BLN60),.WL(WL74));
sram_cell_6t_5 inst_cell_74_61 (.BL(BL61),.BLN(BLN61),.WL(WL74));
sram_cell_6t_5 inst_cell_74_62 (.BL(BL62),.BLN(BLN62),.WL(WL74));
sram_cell_6t_5 inst_cell_74_63 (.BL(BL63),.BLN(BLN63),.WL(WL74));
sram_cell_6t_5 inst_cell_74_64 (.BL(BL64),.BLN(BLN64),.WL(WL74));
sram_cell_6t_5 inst_cell_74_65 (.BL(BL65),.BLN(BLN65),.WL(WL74));
sram_cell_6t_5 inst_cell_74_66 (.BL(BL66),.BLN(BLN66),.WL(WL74));
sram_cell_6t_5 inst_cell_74_67 (.BL(BL67),.BLN(BLN67),.WL(WL74));
sram_cell_6t_5 inst_cell_74_68 (.BL(BL68),.BLN(BLN68),.WL(WL74));
sram_cell_6t_5 inst_cell_74_69 (.BL(BL69),.BLN(BLN69),.WL(WL74));
sram_cell_6t_5 inst_cell_74_70 (.BL(BL70),.BLN(BLN70),.WL(WL74));
sram_cell_6t_5 inst_cell_74_71 (.BL(BL71),.BLN(BLN71),.WL(WL74));
sram_cell_6t_5 inst_cell_74_72 (.BL(BL72),.BLN(BLN72),.WL(WL74));
sram_cell_6t_5 inst_cell_74_73 (.BL(BL73),.BLN(BLN73),.WL(WL74));
sram_cell_6t_5 inst_cell_74_74 (.BL(BL74),.BLN(BLN74),.WL(WL74));
sram_cell_6t_5 inst_cell_74_75 (.BL(BL75),.BLN(BLN75),.WL(WL74));
sram_cell_6t_5 inst_cell_74_76 (.BL(BL76),.BLN(BLN76),.WL(WL74));
sram_cell_6t_5 inst_cell_74_77 (.BL(BL77),.BLN(BLN77),.WL(WL74));
sram_cell_6t_5 inst_cell_74_78 (.BL(BL78),.BLN(BLN78),.WL(WL74));
sram_cell_6t_5 inst_cell_74_79 (.BL(BL79),.BLN(BLN79),.WL(WL74));
sram_cell_6t_5 inst_cell_74_80 (.BL(BL80),.BLN(BLN80),.WL(WL74));
sram_cell_6t_5 inst_cell_74_81 (.BL(BL81),.BLN(BLN81),.WL(WL74));
sram_cell_6t_5 inst_cell_74_82 (.BL(BL82),.BLN(BLN82),.WL(WL74));
sram_cell_6t_5 inst_cell_74_83 (.BL(BL83),.BLN(BLN83),.WL(WL74));
sram_cell_6t_5 inst_cell_74_84 (.BL(BL84),.BLN(BLN84),.WL(WL74));
sram_cell_6t_5 inst_cell_74_85 (.BL(BL85),.BLN(BLN85),.WL(WL74));
sram_cell_6t_5 inst_cell_74_86 (.BL(BL86),.BLN(BLN86),.WL(WL74));
sram_cell_6t_5 inst_cell_74_87 (.BL(BL87),.BLN(BLN87),.WL(WL74));
sram_cell_6t_5 inst_cell_74_88 (.BL(BL88),.BLN(BLN88),.WL(WL74));
sram_cell_6t_5 inst_cell_74_89 (.BL(BL89),.BLN(BLN89),.WL(WL74));
sram_cell_6t_5 inst_cell_74_90 (.BL(BL90),.BLN(BLN90),.WL(WL74));
sram_cell_6t_5 inst_cell_74_91 (.BL(BL91),.BLN(BLN91),.WL(WL74));
sram_cell_6t_5 inst_cell_74_92 (.BL(BL92),.BLN(BLN92),.WL(WL74));
sram_cell_6t_5 inst_cell_74_93 (.BL(BL93),.BLN(BLN93),.WL(WL74));
sram_cell_6t_5 inst_cell_74_94 (.BL(BL94),.BLN(BLN94),.WL(WL74));
sram_cell_6t_5 inst_cell_74_95 (.BL(BL95),.BLN(BLN95),.WL(WL74));
sram_cell_6t_5 inst_cell_74_96 (.BL(BL96),.BLN(BLN96),.WL(WL74));
sram_cell_6t_5 inst_cell_74_97 (.BL(BL97),.BLN(BLN97),.WL(WL74));
sram_cell_6t_5 inst_cell_74_98 (.BL(BL98),.BLN(BLN98),.WL(WL74));
sram_cell_6t_5 inst_cell_74_99 (.BL(BL99),.BLN(BLN99),.WL(WL74));
sram_cell_6t_5 inst_cell_74_100 (.BL(BL100),.BLN(BLN100),.WL(WL74));
sram_cell_6t_5 inst_cell_74_101 (.BL(BL101),.BLN(BLN101),.WL(WL74));
sram_cell_6t_5 inst_cell_74_102 (.BL(BL102),.BLN(BLN102),.WL(WL74));
sram_cell_6t_5 inst_cell_74_103 (.BL(BL103),.BLN(BLN103),.WL(WL74));
sram_cell_6t_5 inst_cell_74_104 (.BL(BL104),.BLN(BLN104),.WL(WL74));
sram_cell_6t_5 inst_cell_74_105 (.BL(BL105),.BLN(BLN105),.WL(WL74));
sram_cell_6t_5 inst_cell_74_106 (.BL(BL106),.BLN(BLN106),.WL(WL74));
sram_cell_6t_5 inst_cell_74_107 (.BL(BL107),.BLN(BLN107),.WL(WL74));
sram_cell_6t_5 inst_cell_74_108 (.BL(BL108),.BLN(BLN108),.WL(WL74));
sram_cell_6t_5 inst_cell_74_109 (.BL(BL109),.BLN(BLN109),.WL(WL74));
sram_cell_6t_5 inst_cell_74_110 (.BL(BL110),.BLN(BLN110),.WL(WL74));
sram_cell_6t_5 inst_cell_74_111 (.BL(BL111),.BLN(BLN111),.WL(WL74));
sram_cell_6t_5 inst_cell_74_112 (.BL(BL112),.BLN(BLN112),.WL(WL74));
sram_cell_6t_5 inst_cell_74_113 (.BL(BL113),.BLN(BLN113),.WL(WL74));
sram_cell_6t_5 inst_cell_74_114 (.BL(BL114),.BLN(BLN114),.WL(WL74));
sram_cell_6t_5 inst_cell_74_115 (.BL(BL115),.BLN(BLN115),.WL(WL74));
sram_cell_6t_5 inst_cell_74_116 (.BL(BL116),.BLN(BLN116),.WL(WL74));
sram_cell_6t_5 inst_cell_74_117 (.BL(BL117),.BLN(BLN117),.WL(WL74));
sram_cell_6t_5 inst_cell_74_118 (.BL(BL118),.BLN(BLN118),.WL(WL74));
sram_cell_6t_5 inst_cell_74_119 (.BL(BL119),.BLN(BLN119),.WL(WL74));
sram_cell_6t_5 inst_cell_74_120 (.BL(BL120),.BLN(BLN120),.WL(WL74));
sram_cell_6t_5 inst_cell_74_121 (.BL(BL121),.BLN(BLN121),.WL(WL74));
sram_cell_6t_5 inst_cell_74_122 (.BL(BL122),.BLN(BLN122),.WL(WL74));
sram_cell_6t_5 inst_cell_74_123 (.BL(BL123),.BLN(BLN123),.WL(WL74));
sram_cell_6t_5 inst_cell_74_124 (.BL(BL124),.BLN(BLN124),.WL(WL74));
sram_cell_6t_5 inst_cell_74_125 (.BL(BL125),.BLN(BLN125),.WL(WL74));
sram_cell_6t_5 inst_cell_74_126 (.BL(BL126),.BLN(BLN126),.WL(WL74));
sram_cell_6t_5 inst_cell_74_127 (.BL(BL127),.BLN(BLN127),.WL(WL74));
sram_cell_6t_5 inst_cell_75_0 (.BL(BL0),.BLN(BLN0),.WL(WL75));
sram_cell_6t_5 inst_cell_75_1 (.BL(BL1),.BLN(BLN1),.WL(WL75));
sram_cell_6t_5 inst_cell_75_2 (.BL(BL2),.BLN(BLN2),.WL(WL75));
sram_cell_6t_5 inst_cell_75_3 (.BL(BL3),.BLN(BLN3),.WL(WL75));
sram_cell_6t_5 inst_cell_75_4 (.BL(BL4),.BLN(BLN4),.WL(WL75));
sram_cell_6t_5 inst_cell_75_5 (.BL(BL5),.BLN(BLN5),.WL(WL75));
sram_cell_6t_5 inst_cell_75_6 (.BL(BL6),.BLN(BLN6),.WL(WL75));
sram_cell_6t_5 inst_cell_75_7 (.BL(BL7),.BLN(BLN7),.WL(WL75));
sram_cell_6t_5 inst_cell_75_8 (.BL(BL8),.BLN(BLN8),.WL(WL75));
sram_cell_6t_5 inst_cell_75_9 (.BL(BL9),.BLN(BLN9),.WL(WL75));
sram_cell_6t_5 inst_cell_75_10 (.BL(BL10),.BLN(BLN10),.WL(WL75));
sram_cell_6t_5 inst_cell_75_11 (.BL(BL11),.BLN(BLN11),.WL(WL75));
sram_cell_6t_5 inst_cell_75_12 (.BL(BL12),.BLN(BLN12),.WL(WL75));
sram_cell_6t_5 inst_cell_75_13 (.BL(BL13),.BLN(BLN13),.WL(WL75));
sram_cell_6t_5 inst_cell_75_14 (.BL(BL14),.BLN(BLN14),.WL(WL75));
sram_cell_6t_5 inst_cell_75_15 (.BL(BL15),.BLN(BLN15),.WL(WL75));
sram_cell_6t_5 inst_cell_75_16 (.BL(BL16),.BLN(BLN16),.WL(WL75));
sram_cell_6t_5 inst_cell_75_17 (.BL(BL17),.BLN(BLN17),.WL(WL75));
sram_cell_6t_5 inst_cell_75_18 (.BL(BL18),.BLN(BLN18),.WL(WL75));
sram_cell_6t_5 inst_cell_75_19 (.BL(BL19),.BLN(BLN19),.WL(WL75));
sram_cell_6t_5 inst_cell_75_20 (.BL(BL20),.BLN(BLN20),.WL(WL75));
sram_cell_6t_5 inst_cell_75_21 (.BL(BL21),.BLN(BLN21),.WL(WL75));
sram_cell_6t_5 inst_cell_75_22 (.BL(BL22),.BLN(BLN22),.WL(WL75));
sram_cell_6t_5 inst_cell_75_23 (.BL(BL23),.BLN(BLN23),.WL(WL75));
sram_cell_6t_5 inst_cell_75_24 (.BL(BL24),.BLN(BLN24),.WL(WL75));
sram_cell_6t_5 inst_cell_75_25 (.BL(BL25),.BLN(BLN25),.WL(WL75));
sram_cell_6t_5 inst_cell_75_26 (.BL(BL26),.BLN(BLN26),.WL(WL75));
sram_cell_6t_5 inst_cell_75_27 (.BL(BL27),.BLN(BLN27),.WL(WL75));
sram_cell_6t_5 inst_cell_75_28 (.BL(BL28),.BLN(BLN28),.WL(WL75));
sram_cell_6t_5 inst_cell_75_29 (.BL(BL29),.BLN(BLN29),.WL(WL75));
sram_cell_6t_5 inst_cell_75_30 (.BL(BL30),.BLN(BLN30),.WL(WL75));
sram_cell_6t_5 inst_cell_75_31 (.BL(BL31),.BLN(BLN31),.WL(WL75));
sram_cell_6t_5 inst_cell_75_32 (.BL(BL32),.BLN(BLN32),.WL(WL75));
sram_cell_6t_5 inst_cell_75_33 (.BL(BL33),.BLN(BLN33),.WL(WL75));
sram_cell_6t_5 inst_cell_75_34 (.BL(BL34),.BLN(BLN34),.WL(WL75));
sram_cell_6t_5 inst_cell_75_35 (.BL(BL35),.BLN(BLN35),.WL(WL75));
sram_cell_6t_5 inst_cell_75_36 (.BL(BL36),.BLN(BLN36),.WL(WL75));
sram_cell_6t_5 inst_cell_75_37 (.BL(BL37),.BLN(BLN37),.WL(WL75));
sram_cell_6t_5 inst_cell_75_38 (.BL(BL38),.BLN(BLN38),.WL(WL75));
sram_cell_6t_5 inst_cell_75_39 (.BL(BL39),.BLN(BLN39),.WL(WL75));
sram_cell_6t_5 inst_cell_75_40 (.BL(BL40),.BLN(BLN40),.WL(WL75));
sram_cell_6t_5 inst_cell_75_41 (.BL(BL41),.BLN(BLN41),.WL(WL75));
sram_cell_6t_5 inst_cell_75_42 (.BL(BL42),.BLN(BLN42),.WL(WL75));
sram_cell_6t_5 inst_cell_75_43 (.BL(BL43),.BLN(BLN43),.WL(WL75));
sram_cell_6t_5 inst_cell_75_44 (.BL(BL44),.BLN(BLN44),.WL(WL75));
sram_cell_6t_5 inst_cell_75_45 (.BL(BL45),.BLN(BLN45),.WL(WL75));
sram_cell_6t_5 inst_cell_75_46 (.BL(BL46),.BLN(BLN46),.WL(WL75));
sram_cell_6t_5 inst_cell_75_47 (.BL(BL47),.BLN(BLN47),.WL(WL75));
sram_cell_6t_5 inst_cell_75_48 (.BL(BL48),.BLN(BLN48),.WL(WL75));
sram_cell_6t_5 inst_cell_75_49 (.BL(BL49),.BLN(BLN49),.WL(WL75));
sram_cell_6t_5 inst_cell_75_50 (.BL(BL50),.BLN(BLN50),.WL(WL75));
sram_cell_6t_5 inst_cell_75_51 (.BL(BL51),.BLN(BLN51),.WL(WL75));
sram_cell_6t_5 inst_cell_75_52 (.BL(BL52),.BLN(BLN52),.WL(WL75));
sram_cell_6t_5 inst_cell_75_53 (.BL(BL53),.BLN(BLN53),.WL(WL75));
sram_cell_6t_5 inst_cell_75_54 (.BL(BL54),.BLN(BLN54),.WL(WL75));
sram_cell_6t_5 inst_cell_75_55 (.BL(BL55),.BLN(BLN55),.WL(WL75));
sram_cell_6t_5 inst_cell_75_56 (.BL(BL56),.BLN(BLN56),.WL(WL75));
sram_cell_6t_5 inst_cell_75_57 (.BL(BL57),.BLN(BLN57),.WL(WL75));
sram_cell_6t_5 inst_cell_75_58 (.BL(BL58),.BLN(BLN58),.WL(WL75));
sram_cell_6t_5 inst_cell_75_59 (.BL(BL59),.BLN(BLN59),.WL(WL75));
sram_cell_6t_5 inst_cell_75_60 (.BL(BL60),.BLN(BLN60),.WL(WL75));
sram_cell_6t_5 inst_cell_75_61 (.BL(BL61),.BLN(BLN61),.WL(WL75));
sram_cell_6t_5 inst_cell_75_62 (.BL(BL62),.BLN(BLN62),.WL(WL75));
sram_cell_6t_5 inst_cell_75_63 (.BL(BL63),.BLN(BLN63),.WL(WL75));
sram_cell_6t_5 inst_cell_75_64 (.BL(BL64),.BLN(BLN64),.WL(WL75));
sram_cell_6t_5 inst_cell_75_65 (.BL(BL65),.BLN(BLN65),.WL(WL75));
sram_cell_6t_5 inst_cell_75_66 (.BL(BL66),.BLN(BLN66),.WL(WL75));
sram_cell_6t_5 inst_cell_75_67 (.BL(BL67),.BLN(BLN67),.WL(WL75));
sram_cell_6t_5 inst_cell_75_68 (.BL(BL68),.BLN(BLN68),.WL(WL75));
sram_cell_6t_5 inst_cell_75_69 (.BL(BL69),.BLN(BLN69),.WL(WL75));
sram_cell_6t_5 inst_cell_75_70 (.BL(BL70),.BLN(BLN70),.WL(WL75));
sram_cell_6t_5 inst_cell_75_71 (.BL(BL71),.BLN(BLN71),.WL(WL75));
sram_cell_6t_5 inst_cell_75_72 (.BL(BL72),.BLN(BLN72),.WL(WL75));
sram_cell_6t_5 inst_cell_75_73 (.BL(BL73),.BLN(BLN73),.WL(WL75));
sram_cell_6t_5 inst_cell_75_74 (.BL(BL74),.BLN(BLN74),.WL(WL75));
sram_cell_6t_5 inst_cell_75_75 (.BL(BL75),.BLN(BLN75),.WL(WL75));
sram_cell_6t_5 inst_cell_75_76 (.BL(BL76),.BLN(BLN76),.WL(WL75));
sram_cell_6t_5 inst_cell_75_77 (.BL(BL77),.BLN(BLN77),.WL(WL75));
sram_cell_6t_5 inst_cell_75_78 (.BL(BL78),.BLN(BLN78),.WL(WL75));
sram_cell_6t_5 inst_cell_75_79 (.BL(BL79),.BLN(BLN79),.WL(WL75));
sram_cell_6t_5 inst_cell_75_80 (.BL(BL80),.BLN(BLN80),.WL(WL75));
sram_cell_6t_5 inst_cell_75_81 (.BL(BL81),.BLN(BLN81),.WL(WL75));
sram_cell_6t_5 inst_cell_75_82 (.BL(BL82),.BLN(BLN82),.WL(WL75));
sram_cell_6t_5 inst_cell_75_83 (.BL(BL83),.BLN(BLN83),.WL(WL75));
sram_cell_6t_5 inst_cell_75_84 (.BL(BL84),.BLN(BLN84),.WL(WL75));
sram_cell_6t_5 inst_cell_75_85 (.BL(BL85),.BLN(BLN85),.WL(WL75));
sram_cell_6t_5 inst_cell_75_86 (.BL(BL86),.BLN(BLN86),.WL(WL75));
sram_cell_6t_5 inst_cell_75_87 (.BL(BL87),.BLN(BLN87),.WL(WL75));
sram_cell_6t_5 inst_cell_75_88 (.BL(BL88),.BLN(BLN88),.WL(WL75));
sram_cell_6t_5 inst_cell_75_89 (.BL(BL89),.BLN(BLN89),.WL(WL75));
sram_cell_6t_5 inst_cell_75_90 (.BL(BL90),.BLN(BLN90),.WL(WL75));
sram_cell_6t_5 inst_cell_75_91 (.BL(BL91),.BLN(BLN91),.WL(WL75));
sram_cell_6t_5 inst_cell_75_92 (.BL(BL92),.BLN(BLN92),.WL(WL75));
sram_cell_6t_5 inst_cell_75_93 (.BL(BL93),.BLN(BLN93),.WL(WL75));
sram_cell_6t_5 inst_cell_75_94 (.BL(BL94),.BLN(BLN94),.WL(WL75));
sram_cell_6t_5 inst_cell_75_95 (.BL(BL95),.BLN(BLN95),.WL(WL75));
sram_cell_6t_5 inst_cell_75_96 (.BL(BL96),.BLN(BLN96),.WL(WL75));
sram_cell_6t_5 inst_cell_75_97 (.BL(BL97),.BLN(BLN97),.WL(WL75));
sram_cell_6t_5 inst_cell_75_98 (.BL(BL98),.BLN(BLN98),.WL(WL75));
sram_cell_6t_5 inst_cell_75_99 (.BL(BL99),.BLN(BLN99),.WL(WL75));
sram_cell_6t_5 inst_cell_75_100 (.BL(BL100),.BLN(BLN100),.WL(WL75));
sram_cell_6t_5 inst_cell_75_101 (.BL(BL101),.BLN(BLN101),.WL(WL75));
sram_cell_6t_5 inst_cell_75_102 (.BL(BL102),.BLN(BLN102),.WL(WL75));
sram_cell_6t_5 inst_cell_75_103 (.BL(BL103),.BLN(BLN103),.WL(WL75));
sram_cell_6t_5 inst_cell_75_104 (.BL(BL104),.BLN(BLN104),.WL(WL75));
sram_cell_6t_5 inst_cell_75_105 (.BL(BL105),.BLN(BLN105),.WL(WL75));
sram_cell_6t_5 inst_cell_75_106 (.BL(BL106),.BLN(BLN106),.WL(WL75));
sram_cell_6t_5 inst_cell_75_107 (.BL(BL107),.BLN(BLN107),.WL(WL75));
sram_cell_6t_5 inst_cell_75_108 (.BL(BL108),.BLN(BLN108),.WL(WL75));
sram_cell_6t_5 inst_cell_75_109 (.BL(BL109),.BLN(BLN109),.WL(WL75));
sram_cell_6t_5 inst_cell_75_110 (.BL(BL110),.BLN(BLN110),.WL(WL75));
sram_cell_6t_5 inst_cell_75_111 (.BL(BL111),.BLN(BLN111),.WL(WL75));
sram_cell_6t_5 inst_cell_75_112 (.BL(BL112),.BLN(BLN112),.WL(WL75));
sram_cell_6t_5 inst_cell_75_113 (.BL(BL113),.BLN(BLN113),.WL(WL75));
sram_cell_6t_5 inst_cell_75_114 (.BL(BL114),.BLN(BLN114),.WL(WL75));
sram_cell_6t_5 inst_cell_75_115 (.BL(BL115),.BLN(BLN115),.WL(WL75));
sram_cell_6t_5 inst_cell_75_116 (.BL(BL116),.BLN(BLN116),.WL(WL75));
sram_cell_6t_5 inst_cell_75_117 (.BL(BL117),.BLN(BLN117),.WL(WL75));
sram_cell_6t_5 inst_cell_75_118 (.BL(BL118),.BLN(BLN118),.WL(WL75));
sram_cell_6t_5 inst_cell_75_119 (.BL(BL119),.BLN(BLN119),.WL(WL75));
sram_cell_6t_5 inst_cell_75_120 (.BL(BL120),.BLN(BLN120),.WL(WL75));
sram_cell_6t_5 inst_cell_75_121 (.BL(BL121),.BLN(BLN121),.WL(WL75));
sram_cell_6t_5 inst_cell_75_122 (.BL(BL122),.BLN(BLN122),.WL(WL75));
sram_cell_6t_5 inst_cell_75_123 (.BL(BL123),.BLN(BLN123),.WL(WL75));
sram_cell_6t_5 inst_cell_75_124 (.BL(BL124),.BLN(BLN124),.WL(WL75));
sram_cell_6t_5 inst_cell_75_125 (.BL(BL125),.BLN(BLN125),.WL(WL75));
sram_cell_6t_5 inst_cell_75_126 (.BL(BL126),.BLN(BLN126),.WL(WL75));
sram_cell_6t_5 inst_cell_75_127 (.BL(BL127),.BLN(BLN127),.WL(WL75));
sram_cell_6t_5 inst_cell_76_0 (.BL(BL0),.BLN(BLN0),.WL(WL76));
sram_cell_6t_5 inst_cell_76_1 (.BL(BL1),.BLN(BLN1),.WL(WL76));
sram_cell_6t_5 inst_cell_76_2 (.BL(BL2),.BLN(BLN2),.WL(WL76));
sram_cell_6t_5 inst_cell_76_3 (.BL(BL3),.BLN(BLN3),.WL(WL76));
sram_cell_6t_5 inst_cell_76_4 (.BL(BL4),.BLN(BLN4),.WL(WL76));
sram_cell_6t_5 inst_cell_76_5 (.BL(BL5),.BLN(BLN5),.WL(WL76));
sram_cell_6t_5 inst_cell_76_6 (.BL(BL6),.BLN(BLN6),.WL(WL76));
sram_cell_6t_5 inst_cell_76_7 (.BL(BL7),.BLN(BLN7),.WL(WL76));
sram_cell_6t_5 inst_cell_76_8 (.BL(BL8),.BLN(BLN8),.WL(WL76));
sram_cell_6t_5 inst_cell_76_9 (.BL(BL9),.BLN(BLN9),.WL(WL76));
sram_cell_6t_5 inst_cell_76_10 (.BL(BL10),.BLN(BLN10),.WL(WL76));
sram_cell_6t_5 inst_cell_76_11 (.BL(BL11),.BLN(BLN11),.WL(WL76));
sram_cell_6t_5 inst_cell_76_12 (.BL(BL12),.BLN(BLN12),.WL(WL76));
sram_cell_6t_5 inst_cell_76_13 (.BL(BL13),.BLN(BLN13),.WL(WL76));
sram_cell_6t_5 inst_cell_76_14 (.BL(BL14),.BLN(BLN14),.WL(WL76));
sram_cell_6t_5 inst_cell_76_15 (.BL(BL15),.BLN(BLN15),.WL(WL76));
sram_cell_6t_5 inst_cell_76_16 (.BL(BL16),.BLN(BLN16),.WL(WL76));
sram_cell_6t_5 inst_cell_76_17 (.BL(BL17),.BLN(BLN17),.WL(WL76));
sram_cell_6t_5 inst_cell_76_18 (.BL(BL18),.BLN(BLN18),.WL(WL76));
sram_cell_6t_5 inst_cell_76_19 (.BL(BL19),.BLN(BLN19),.WL(WL76));
sram_cell_6t_5 inst_cell_76_20 (.BL(BL20),.BLN(BLN20),.WL(WL76));
sram_cell_6t_5 inst_cell_76_21 (.BL(BL21),.BLN(BLN21),.WL(WL76));
sram_cell_6t_5 inst_cell_76_22 (.BL(BL22),.BLN(BLN22),.WL(WL76));
sram_cell_6t_5 inst_cell_76_23 (.BL(BL23),.BLN(BLN23),.WL(WL76));
sram_cell_6t_5 inst_cell_76_24 (.BL(BL24),.BLN(BLN24),.WL(WL76));
sram_cell_6t_5 inst_cell_76_25 (.BL(BL25),.BLN(BLN25),.WL(WL76));
sram_cell_6t_5 inst_cell_76_26 (.BL(BL26),.BLN(BLN26),.WL(WL76));
sram_cell_6t_5 inst_cell_76_27 (.BL(BL27),.BLN(BLN27),.WL(WL76));
sram_cell_6t_5 inst_cell_76_28 (.BL(BL28),.BLN(BLN28),.WL(WL76));
sram_cell_6t_5 inst_cell_76_29 (.BL(BL29),.BLN(BLN29),.WL(WL76));
sram_cell_6t_5 inst_cell_76_30 (.BL(BL30),.BLN(BLN30),.WL(WL76));
sram_cell_6t_5 inst_cell_76_31 (.BL(BL31),.BLN(BLN31),.WL(WL76));
sram_cell_6t_5 inst_cell_76_32 (.BL(BL32),.BLN(BLN32),.WL(WL76));
sram_cell_6t_5 inst_cell_76_33 (.BL(BL33),.BLN(BLN33),.WL(WL76));
sram_cell_6t_5 inst_cell_76_34 (.BL(BL34),.BLN(BLN34),.WL(WL76));
sram_cell_6t_5 inst_cell_76_35 (.BL(BL35),.BLN(BLN35),.WL(WL76));
sram_cell_6t_5 inst_cell_76_36 (.BL(BL36),.BLN(BLN36),.WL(WL76));
sram_cell_6t_5 inst_cell_76_37 (.BL(BL37),.BLN(BLN37),.WL(WL76));
sram_cell_6t_5 inst_cell_76_38 (.BL(BL38),.BLN(BLN38),.WL(WL76));
sram_cell_6t_5 inst_cell_76_39 (.BL(BL39),.BLN(BLN39),.WL(WL76));
sram_cell_6t_5 inst_cell_76_40 (.BL(BL40),.BLN(BLN40),.WL(WL76));
sram_cell_6t_5 inst_cell_76_41 (.BL(BL41),.BLN(BLN41),.WL(WL76));
sram_cell_6t_5 inst_cell_76_42 (.BL(BL42),.BLN(BLN42),.WL(WL76));
sram_cell_6t_5 inst_cell_76_43 (.BL(BL43),.BLN(BLN43),.WL(WL76));
sram_cell_6t_5 inst_cell_76_44 (.BL(BL44),.BLN(BLN44),.WL(WL76));
sram_cell_6t_5 inst_cell_76_45 (.BL(BL45),.BLN(BLN45),.WL(WL76));
sram_cell_6t_5 inst_cell_76_46 (.BL(BL46),.BLN(BLN46),.WL(WL76));
sram_cell_6t_5 inst_cell_76_47 (.BL(BL47),.BLN(BLN47),.WL(WL76));
sram_cell_6t_5 inst_cell_76_48 (.BL(BL48),.BLN(BLN48),.WL(WL76));
sram_cell_6t_5 inst_cell_76_49 (.BL(BL49),.BLN(BLN49),.WL(WL76));
sram_cell_6t_5 inst_cell_76_50 (.BL(BL50),.BLN(BLN50),.WL(WL76));
sram_cell_6t_5 inst_cell_76_51 (.BL(BL51),.BLN(BLN51),.WL(WL76));
sram_cell_6t_5 inst_cell_76_52 (.BL(BL52),.BLN(BLN52),.WL(WL76));
sram_cell_6t_5 inst_cell_76_53 (.BL(BL53),.BLN(BLN53),.WL(WL76));
sram_cell_6t_5 inst_cell_76_54 (.BL(BL54),.BLN(BLN54),.WL(WL76));
sram_cell_6t_5 inst_cell_76_55 (.BL(BL55),.BLN(BLN55),.WL(WL76));
sram_cell_6t_5 inst_cell_76_56 (.BL(BL56),.BLN(BLN56),.WL(WL76));
sram_cell_6t_5 inst_cell_76_57 (.BL(BL57),.BLN(BLN57),.WL(WL76));
sram_cell_6t_5 inst_cell_76_58 (.BL(BL58),.BLN(BLN58),.WL(WL76));
sram_cell_6t_5 inst_cell_76_59 (.BL(BL59),.BLN(BLN59),.WL(WL76));
sram_cell_6t_5 inst_cell_76_60 (.BL(BL60),.BLN(BLN60),.WL(WL76));
sram_cell_6t_5 inst_cell_76_61 (.BL(BL61),.BLN(BLN61),.WL(WL76));
sram_cell_6t_5 inst_cell_76_62 (.BL(BL62),.BLN(BLN62),.WL(WL76));
sram_cell_6t_5 inst_cell_76_63 (.BL(BL63),.BLN(BLN63),.WL(WL76));
sram_cell_6t_5 inst_cell_76_64 (.BL(BL64),.BLN(BLN64),.WL(WL76));
sram_cell_6t_5 inst_cell_76_65 (.BL(BL65),.BLN(BLN65),.WL(WL76));
sram_cell_6t_5 inst_cell_76_66 (.BL(BL66),.BLN(BLN66),.WL(WL76));
sram_cell_6t_5 inst_cell_76_67 (.BL(BL67),.BLN(BLN67),.WL(WL76));
sram_cell_6t_5 inst_cell_76_68 (.BL(BL68),.BLN(BLN68),.WL(WL76));
sram_cell_6t_5 inst_cell_76_69 (.BL(BL69),.BLN(BLN69),.WL(WL76));
sram_cell_6t_5 inst_cell_76_70 (.BL(BL70),.BLN(BLN70),.WL(WL76));
sram_cell_6t_5 inst_cell_76_71 (.BL(BL71),.BLN(BLN71),.WL(WL76));
sram_cell_6t_5 inst_cell_76_72 (.BL(BL72),.BLN(BLN72),.WL(WL76));
sram_cell_6t_5 inst_cell_76_73 (.BL(BL73),.BLN(BLN73),.WL(WL76));
sram_cell_6t_5 inst_cell_76_74 (.BL(BL74),.BLN(BLN74),.WL(WL76));
sram_cell_6t_5 inst_cell_76_75 (.BL(BL75),.BLN(BLN75),.WL(WL76));
sram_cell_6t_5 inst_cell_76_76 (.BL(BL76),.BLN(BLN76),.WL(WL76));
sram_cell_6t_5 inst_cell_76_77 (.BL(BL77),.BLN(BLN77),.WL(WL76));
sram_cell_6t_5 inst_cell_76_78 (.BL(BL78),.BLN(BLN78),.WL(WL76));
sram_cell_6t_5 inst_cell_76_79 (.BL(BL79),.BLN(BLN79),.WL(WL76));
sram_cell_6t_5 inst_cell_76_80 (.BL(BL80),.BLN(BLN80),.WL(WL76));
sram_cell_6t_5 inst_cell_76_81 (.BL(BL81),.BLN(BLN81),.WL(WL76));
sram_cell_6t_5 inst_cell_76_82 (.BL(BL82),.BLN(BLN82),.WL(WL76));
sram_cell_6t_5 inst_cell_76_83 (.BL(BL83),.BLN(BLN83),.WL(WL76));
sram_cell_6t_5 inst_cell_76_84 (.BL(BL84),.BLN(BLN84),.WL(WL76));
sram_cell_6t_5 inst_cell_76_85 (.BL(BL85),.BLN(BLN85),.WL(WL76));
sram_cell_6t_5 inst_cell_76_86 (.BL(BL86),.BLN(BLN86),.WL(WL76));
sram_cell_6t_5 inst_cell_76_87 (.BL(BL87),.BLN(BLN87),.WL(WL76));
sram_cell_6t_5 inst_cell_76_88 (.BL(BL88),.BLN(BLN88),.WL(WL76));
sram_cell_6t_5 inst_cell_76_89 (.BL(BL89),.BLN(BLN89),.WL(WL76));
sram_cell_6t_5 inst_cell_76_90 (.BL(BL90),.BLN(BLN90),.WL(WL76));
sram_cell_6t_5 inst_cell_76_91 (.BL(BL91),.BLN(BLN91),.WL(WL76));
sram_cell_6t_5 inst_cell_76_92 (.BL(BL92),.BLN(BLN92),.WL(WL76));
sram_cell_6t_5 inst_cell_76_93 (.BL(BL93),.BLN(BLN93),.WL(WL76));
sram_cell_6t_5 inst_cell_76_94 (.BL(BL94),.BLN(BLN94),.WL(WL76));
sram_cell_6t_5 inst_cell_76_95 (.BL(BL95),.BLN(BLN95),.WL(WL76));
sram_cell_6t_5 inst_cell_76_96 (.BL(BL96),.BLN(BLN96),.WL(WL76));
sram_cell_6t_5 inst_cell_76_97 (.BL(BL97),.BLN(BLN97),.WL(WL76));
sram_cell_6t_5 inst_cell_76_98 (.BL(BL98),.BLN(BLN98),.WL(WL76));
sram_cell_6t_5 inst_cell_76_99 (.BL(BL99),.BLN(BLN99),.WL(WL76));
sram_cell_6t_5 inst_cell_76_100 (.BL(BL100),.BLN(BLN100),.WL(WL76));
sram_cell_6t_5 inst_cell_76_101 (.BL(BL101),.BLN(BLN101),.WL(WL76));
sram_cell_6t_5 inst_cell_76_102 (.BL(BL102),.BLN(BLN102),.WL(WL76));
sram_cell_6t_5 inst_cell_76_103 (.BL(BL103),.BLN(BLN103),.WL(WL76));
sram_cell_6t_5 inst_cell_76_104 (.BL(BL104),.BLN(BLN104),.WL(WL76));
sram_cell_6t_5 inst_cell_76_105 (.BL(BL105),.BLN(BLN105),.WL(WL76));
sram_cell_6t_5 inst_cell_76_106 (.BL(BL106),.BLN(BLN106),.WL(WL76));
sram_cell_6t_5 inst_cell_76_107 (.BL(BL107),.BLN(BLN107),.WL(WL76));
sram_cell_6t_5 inst_cell_76_108 (.BL(BL108),.BLN(BLN108),.WL(WL76));
sram_cell_6t_5 inst_cell_76_109 (.BL(BL109),.BLN(BLN109),.WL(WL76));
sram_cell_6t_5 inst_cell_76_110 (.BL(BL110),.BLN(BLN110),.WL(WL76));
sram_cell_6t_5 inst_cell_76_111 (.BL(BL111),.BLN(BLN111),.WL(WL76));
sram_cell_6t_5 inst_cell_76_112 (.BL(BL112),.BLN(BLN112),.WL(WL76));
sram_cell_6t_5 inst_cell_76_113 (.BL(BL113),.BLN(BLN113),.WL(WL76));
sram_cell_6t_5 inst_cell_76_114 (.BL(BL114),.BLN(BLN114),.WL(WL76));
sram_cell_6t_5 inst_cell_76_115 (.BL(BL115),.BLN(BLN115),.WL(WL76));
sram_cell_6t_5 inst_cell_76_116 (.BL(BL116),.BLN(BLN116),.WL(WL76));
sram_cell_6t_5 inst_cell_76_117 (.BL(BL117),.BLN(BLN117),.WL(WL76));
sram_cell_6t_5 inst_cell_76_118 (.BL(BL118),.BLN(BLN118),.WL(WL76));
sram_cell_6t_5 inst_cell_76_119 (.BL(BL119),.BLN(BLN119),.WL(WL76));
sram_cell_6t_5 inst_cell_76_120 (.BL(BL120),.BLN(BLN120),.WL(WL76));
sram_cell_6t_5 inst_cell_76_121 (.BL(BL121),.BLN(BLN121),.WL(WL76));
sram_cell_6t_5 inst_cell_76_122 (.BL(BL122),.BLN(BLN122),.WL(WL76));
sram_cell_6t_5 inst_cell_76_123 (.BL(BL123),.BLN(BLN123),.WL(WL76));
sram_cell_6t_5 inst_cell_76_124 (.BL(BL124),.BLN(BLN124),.WL(WL76));
sram_cell_6t_5 inst_cell_76_125 (.BL(BL125),.BLN(BLN125),.WL(WL76));
sram_cell_6t_5 inst_cell_76_126 (.BL(BL126),.BLN(BLN126),.WL(WL76));
sram_cell_6t_5 inst_cell_76_127 (.BL(BL127),.BLN(BLN127),.WL(WL76));
sram_cell_6t_5 inst_cell_77_0 (.BL(BL0),.BLN(BLN0),.WL(WL77));
sram_cell_6t_5 inst_cell_77_1 (.BL(BL1),.BLN(BLN1),.WL(WL77));
sram_cell_6t_5 inst_cell_77_2 (.BL(BL2),.BLN(BLN2),.WL(WL77));
sram_cell_6t_5 inst_cell_77_3 (.BL(BL3),.BLN(BLN3),.WL(WL77));
sram_cell_6t_5 inst_cell_77_4 (.BL(BL4),.BLN(BLN4),.WL(WL77));
sram_cell_6t_5 inst_cell_77_5 (.BL(BL5),.BLN(BLN5),.WL(WL77));
sram_cell_6t_5 inst_cell_77_6 (.BL(BL6),.BLN(BLN6),.WL(WL77));
sram_cell_6t_5 inst_cell_77_7 (.BL(BL7),.BLN(BLN7),.WL(WL77));
sram_cell_6t_5 inst_cell_77_8 (.BL(BL8),.BLN(BLN8),.WL(WL77));
sram_cell_6t_5 inst_cell_77_9 (.BL(BL9),.BLN(BLN9),.WL(WL77));
sram_cell_6t_5 inst_cell_77_10 (.BL(BL10),.BLN(BLN10),.WL(WL77));
sram_cell_6t_5 inst_cell_77_11 (.BL(BL11),.BLN(BLN11),.WL(WL77));
sram_cell_6t_5 inst_cell_77_12 (.BL(BL12),.BLN(BLN12),.WL(WL77));
sram_cell_6t_5 inst_cell_77_13 (.BL(BL13),.BLN(BLN13),.WL(WL77));
sram_cell_6t_5 inst_cell_77_14 (.BL(BL14),.BLN(BLN14),.WL(WL77));
sram_cell_6t_5 inst_cell_77_15 (.BL(BL15),.BLN(BLN15),.WL(WL77));
sram_cell_6t_5 inst_cell_77_16 (.BL(BL16),.BLN(BLN16),.WL(WL77));
sram_cell_6t_5 inst_cell_77_17 (.BL(BL17),.BLN(BLN17),.WL(WL77));
sram_cell_6t_5 inst_cell_77_18 (.BL(BL18),.BLN(BLN18),.WL(WL77));
sram_cell_6t_5 inst_cell_77_19 (.BL(BL19),.BLN(BLN19),.WL(WL77));
sram_cell_6t_5 inst_cell_77_20 (.BL(BL20),.BLN(BLN20),.WL(WL77));
sram_cell_6t_5 inst_cell_77_21 (.BL(BL21),.BLN(BLN21),.WL(WL77));
sram_cell_6t_5 inst_cell_77_22 (.BL(BL22),.BLN(BLN22),.WL(WL77));
sram_cell_6t_5 inst_cell_77_23 (.BL(BL23),.BLN(BLN23),.WL(WL77));
sram_cell_6t_5 inst_cell_77_24 (.BL(BL24),.BLN(BLN24),.WL(WL77));
sram_cell_6t_5 inst_cell_77_25 (.BL(BL25),.BLN(BLN25),.WL(WL77));
sram_cell_6t_5 inst_cell_77_26 (.BL(BL26),.BLN(BLN26),.WL(WL77));
sram_cell_6t_5 inst_cell_77_27 (.BL(BL27),.BLN(BLN27),.WL(WL77));
sram_cell_6t_5 inst_cell_77_28 (.BL(BL28),.BLN(BLN28),.WL(WL77));
sram_cell_6t_5 inst_cell_77_29 (.BL(BL29),.BLN(BLN29),.WL(WL77));
sram_cell_6t_5 inst_cell_77_30 (.BL(BL30),.BLN(BLN30),.WL(WL77));
sram_cell_6t_5 inst_cell_77_31 (.BL(BL31),.BLN(BLN31),.WL(WL77));
sram_cell_6t_5 inst_cell_77_32 (.BL(BL32),.BLN(BLN32),.WL(WL77));
sram_cell_6t_5 inst_cell_77_33 (.BL(BL33),.BLN(BLN33),.WL(WL77));
sram_cell_6t_5 inst_cell_77_34 (.BL(BL34),.BLN(BLN34),.WL(WL77));
sram_cell_6t_5 inst_cell_77_35 (.BL(BL35),.BLN(BLN35),.WL(WL77));
sram_cell_6t_5 inst_cell_77_36 (.BL(BL36),.BLN(BLN36),.WL(WL77));
sram_cell_6t_5 inst_cell_77_37 (.BL(BL37),.BLN(BLN37),.WL(WL77));
sram_cell_6t_5 inst_cell_77_38 (.BL(BL38),.BLN(BLN38),.WL(WL77));
sram_cell_6t_5 inst_cell_77_39 (.BL(BL39),.BLN(BLN39),.WL(WL77));
sram_cell_6t_5 inst_cell_77_40 (.BL(BL40),.BLN(BLN40),.WL(WL77));
sram_cell_6t_5 inst_cell_77_41 (.BL(BL41),.BLN(BLN41),.WL(WL77));
sram_cell_6t_5 inst_cell_77_42 (.BL(BL42),.BLN(BLN42),.WL(WL77));
sram_cell_6t_5 inst_cell_77_43 (.BL(BL43),.BLN(BLN43),.WL(WL77));
sram_cell_6t_5 inst_cell_77_44 (.BL(BL44),.BLN(BLN44),.WL(WL77));
sram_cell_6t_5 inst_cell_77_45 (.BL(BL45),.BLN(BLN45),.WL(WL77));
sram_cell_6t_5 inst_cell_77_46 (.BL(BL46),.BLN(BLN46),.WL(WL77));
sram_cell_6t_5 inst_cell_77_47 (.BL(BL47),.BLN(BLN47),.WL(WL77));
sram_cell_6t_5 inst_cell_77_48 (.BL(BL48),.BLN(BLN48),.WL(WL77));
sram_cell_6t_5 inst_cell_77_49 (.BL(BL49),.BLN(BLN49),.WL(WL77));
sram_cell_6t_5 inst_cell_77_50 (.BL(BL50),.BLN(BLN50),.WL(WL77));
sram_cell_6t_5 inst_cell_77_51 (.BL(BL51),.BLN(BLN51),.WL(WL77));
sram_cell_6t_5 inst_cell_77_52 (.BL(BL52),.BLN(BLN52),.WL(WL77));
sram_cell_6t_5 inst_cell_77_53 (.BL(BL53),.BLN(BLN53),.WL(WL77));
sram_cell_6t_5 inst_cell_77_54 (.BL(BL54),.BLN(BLN54),.WL(WL77));
sram_cell_6t_5 inst_cell_77_55 (.BL(BL55),.BLN(BLN55),.WL(WL77));
sram_cell_6t_5 inst_cell_77_56 (.BL(BL56),.BLN(BLN56),.WL(WL77));
sram_cell_6t_5 inst_cell_77_57 (.BL(BL57),.BLN(BLN57),.WL(WL77));
sram_cell_6t_5 inst_cell_77_58 (.BL(BL58),.BLN(BLN58),.WL(WL77));
sram_cell_6t_5 inst_cell_77_59 (.BL(BL59),.BLN(BLN59),.WL(WL77));
sram_cell_6t_5 inst_cell_77_60 (.BL(BL60),.BLN(BLN60),.WL(WL77));
sram_cell_6t_5 inst_cell_77_61 (.BL(BL61),.BLN(BLN61),.WL(WL77));
sram_cell_6t_5 inst_cell_77_62 (.BL(BL62),.BLN(BLN62),.WL(WL77));
sram_cell_6t_5 inst_cell_77_63 (.BL(BL63),.BLN(BLN63),.WL(WL77));
sram_cell_6t_5 inst_cell_77_64 (.BL(BL64),.BLN(BLN64),.WL(WL77));
sram_cell_6t_5 inst_cell_77_65 (.BL(BL65),.BLN(BLN65),.WL(WL77));
sram_cell_6t_5 inst_cell_77_66 (.BL(BL66),.BLN(BLN66),.WL(WL77));
sram_cell_6t_5 inst_cell_77_67 (.BL(BL67),.BLN(BLN67),.WL(WL77));
sram_cell_6t_5 inst_cell_77_68 (.BL(BL68),.BLN(BLN68),.WL(WL77));
sram_cell_6t_5 inst_cell_77_69 (.BL(BL69),.BLN(BLN69),.WL(WL77));
sram_cell_6t_5 inst_cell_77_70 (.BL(BL70),.BLN(BLN70),.WL(WL77));
sram_cell_6t_5 inst_cell_77_71 (.BL(BL71),.BLN(BLN71),.WL(WL77));
sram_cell_6t_5 inst_cell_77_72 (.BL(BL72),.BLN(BLN72),.WL(WL77));
sram_cell_6t_5 inst_cell_77_73 (.BL(BL73),.BLN(BLN73),.WL(WL77));
sram_cell_6t_5 inst_cell_77_74 (.BL(BL74),.BLN(BLN74),.WL(WL77));
sram_cell_6t_5 inst_cell_77_75 (.BL(BL75),.BLN(BLN75),.WL(WL77));
sram_cell_6t_5 inst_cell_77_76 (.BL(BL76),.BLN(BLN76),.WL(WL77));
sram_cell_6t_5 inst_cell_77_77 (.BL(BL77),.BLN(BLN77),.WL(WL77));
sram_cell_6t_5 inst_cell_77_78 (.BL(BL78),.BLN(BLN78),.WL(WL77));
sram_cell_6t_5 inst_cell_77_79 (.BL(BL79),.BLN(BLN79),.WL(WL77));
sram_cell_6t_5 inst_cell_77_80 (.BL(BL80),.BLN(BLN80),.WL(WL77));
sram_cell_6t_5 inst_cell_77_81 (.BL(BL81),.BLN(BLN81),.WL(WL77));
sram_cell_6t_5 inst_cell_77_82 (.BL(BL82),.BLN(BLN82),.WL(WL77));
sram_cell_6t_5 inst_cell_77_83 (.BL(BL83),.BLN(BLN83),.WL(WL77));
sram_cell_6t_5 inst_cell_77_84 (.BL(BL84),.BLN(BLN84),.WL(WL77));
sram_cell_6t_5 inst_cell_77_85 (.BL(BL85),.BLN(BLN85),.WL(WL77));
sram_cell_6t_5 inst_cell_77_86 (.BL(BL86),.BLN(BLN86),.WL(WL77));
sram_cell_6t_5 inst_cell_77_87 (.BL(BL87),.BLN(BLN87),.WL(WL77));
sram_cell_6t_5 inst_cell_77_88 (.BL(BL88),.BLN(BLN88),.WL(WL77));
sram_cell_6t_5 inst_cell_77_89 (.BL(BL89),.BLN(BLN89),.WL(WL77));
sram_cell_6t_5 inst_cell_77_90 (.BL(BL90),.BLN(BLN90),.WL(WL77));
sram_cell_6t_5 inst_cell_77_91 (.BL(BL91),.BLN(BLN91),.WL(WL77));
sram_cell_6t_5 inst_cell_77_92 (.BL(BL92),.BLN(BLN92),.WL(WL77));
sram_cell_6t_5 inst_cell_77_93 (.BL(BL93),.BLN(BLN93),.WL(WL77));
sram_cell_6t_5 inst_cell_77_94 (.BL(BL94),.BLN(BLN94),.WL(WL77));
sram_cell_6t_5 inst_cell_77_95 (.BL(BL95),.BLN(BLN95),.WL(WL77));
sram_cell_6t_5 inst_cell_77_96 (.BL(BL96),.BLN(BLN96),.WL(WL77));
sram_cell_6t_5 inst_cell_77_97 (.BL(BL97),.BLN(BLN97),.WL(WL77));
sram_cell_6t_5 inst_cell_77_98 (.BL(BL98),.BLN(BLN98),.WL(WL77));
sram_cell_6t_5 inst_cell_77_99 (.BL(BL99),.BLN(BLN99),.WL(WL77));
sram_cell_6t_5 inst_cell_77_100 (.BL(BL100),.BLN(BLN100),.WL(WL77));
sram_cell_6t_5 inst_cell_77_101 (.BL(BL101),.BLN(BLN101),.WL(WL77));
sram_cell_6t_5 inst_cell_77_102 (.BL(BL102),.BLN(BLN102),.WL(WL77));
sram_cell_6t_5 inst_cell_77_103 (.BL(BL103),.BLN(BLN103),.WL(WL77));
sram_cell_6t_5 inst_cell_77_104 (.BL(BL104),.BLN(BLN104),.WL(WL77));
sram_cell_6t_5 inst_cell_77_105 (.BL(BL105),.BLN(BLN105),.WL(WL77));
sram_cell_6t_5 inst_cell_77_106 (.BL(BL106),.BLN(BLN106),.WL(WL77));
sram_cell_6t_5 inst_cell_77_107 (.BL(BL107),.BLN(BLN107),.WL(WL77));
sram_cell_6t_5 inst_cell_77_108 (.BL(BL108),.BLN(BLN108),.WL(WL77));
sram_cell_6t_5 inst_cell_77_109 (.BL(BL109),.BLN(BLN109),.WL(WL77));
sram_cell_6t_5 inst_cell_77_110 (.BL(BL110),.BLN(BLN110),.WL(WL77));
sram_cell_6t_5 inst_cell_77_111 (.BL(BL111),.BLN(BLN111),.WL(WL77));
sram_cell_6t_5 inst_cell_77_112 (.BL(BL112),.BLN(BLN112),.WL(WL77));
sram_cell_6t_5 inst_cell_77_113 (.BL(BL113),.BLN(BLN113),.WL(WL77));
sram_cell_6t_5 inst_cell_77_114 (.BL(BL114),.BLN(BLN114),.WL(WL77));
sram_cell_6t_5 inst_cell_77_115 (.BL(BL115),.BLN(BLN115),.WL(WL77));
sram_cell_6t_5 inst_cell_77_116 (.BL(BL116),.BLN(BLN116),.WL(WL77));
sram_cell_6t_5 inst_cell_77_117 (.BL(BL117),.BLN(BLN117),.WL(WL77));
sram_cell_6t_5 inst_cell_77_118 (.BL(BL118),.BLN(BLN118),.WL(WL77));
sram_cell_6t_5 inst_cell_77_119 (.BL(BL119),.BLN(BLN119),.WL(WL77));
sram_cell_6t_5 inst_cell_77_120 (.BL(BL120),.BLN(BLN120),.WL(WL77));
sram_cell_6t_5 inst_cell_77_121 (.BL(BL121),.BLN(BLN121),.WL(WL77));
sram_cell_6t_5 inst_cell_77_122 (.BL(BL122),.BLN(BLN122),.WL(WL77));
sram_cell_6t_5 inst_cell_77_123 (.BL(BL123),.BLN(BLN123),.WL(WL77));
sram_cell_6t_5 inst_cell_77_124 (.BL(BL124),.BLN(BLN124),.WL(WL77));
sram_cell_6t_5 inst_cell_77_125 (.BL(BL125),.BLN(BLN125),.WL(WL77));
sram_cell_6t_5 inst_cell_77_126 (.BL(BL126),.BLN(BLN126),.WL(WL77));
sram_cell_6t_5 inst_cell_77_127 (.BL(BL127),.BLN(BLN127),.WL(WL77));
sram_cell_6t_5 inst_cell_78_0 (.BL(BL0),.BLN(BLN0),.WL(WL78));
sram_cell_6t_5 inst_cell_78_1 (.BL(BL1),.BLN(BLN1),.WL(WL78));
sram_cell_6t_5 inst_cell_78_2 (.BL(BL2),.BLN(BLN2),.WL(WL78));
sram_cell_6t_5 inst_cell_78_3 (.BL(BL3),.BLN(BLN3),.WL(WL78));
sram_cell_6t_5 inst_cell_78_4 (.BL(BL4),.BLN(BLN4),.WL(WL78));
sram_cell_6t_5 inst_cell_78_5 (.BL(BL5),.BLN(BLN5),.WL(WL78));
sram_cell_6t_5 inst_cell_78_6 (.BL(BL6),.BLN(BLN6),.WL(WL78));
sram_cell_6t_5 inst_cell_78_7 (.BL(BL7),.BLN(BLN7),.WL(WL78));
sram_cell_6t_5 inst_cell_78_8 (.BL(BL8),.BLN(BLN8),.WL(WL78));
sram_cell_6t_5 inst_cell_78_9 (.BL(BL9),.BLN(BLN9),.WL(WL78));
sram_cell_6t_5 inst_cell_78_10 (.BL(BL10),.BLN(BLN10),.WL(WL78));
sram_cell_6t_5 inst_cell_78_11 (.BL(BL11),.BLN(BLN11),.WL(WL78));
sram_cell_6t_5 inst_cell_78_12 (.BL(BL12),.BLN(BLN12),.WL(WL78));
sram_cell_6t_5 inst_cell_78_13 (.BL(BL13),.BLN(BLN13),.WL(WL78));
sram_cell_6t_5 inst_cell_78_14 (.BL(BL14),.BLN(BLN14),.WL(WL78));
sram_cell_6t_5 inst_cell_78_15 (.BL(BL15),.BLN(BLN15),.WL(WL78));
sram_cell_6t_5 inst_cell_78_16 (.BL(BL16),.BLN(BLN16),.WL(WL78));
sram_cell_6t_5 inst_cell_78_17 (.BL(BL17),.BLN(BLN17),.WL(WL78));
sram_cell_6t_5 inst_cell_78_18 (.BL(BL18),.BLN(BLN18),.WL(WL78));
sram_cell_6t_5 inst_cell_78_19 (.BL(BL19),.BLN(BLN19),.WL(WL78));
sram_cell_6t_5 inst_cell_78_20 (.BL(BL20),.BLN(BLN20),.WL(WL78));
sram_cell_6t_5 inst_cell_78_21 (.BL(BL21),.BLN(BLN21),.WL(WL78));
sram_cell_6t_5 inst_cell_78_22 (.BL(BL22),.BLN(BLN22),.WL(WL78));
sram_cell_6t_5 inst_cell_78_23 (.BL(BL23),.BLN(BLN23),.WL(WL78));
sram_cell_6t_5 inst_cell_78_24 (.BL(BL24),.BLN(BLN24),.WL(WL78));
sram_cell_6t_5 inst_cell_78_25 (.BL(BL25),.BLN(BLN25),.WL(WL78));
sram_cell_6t_5 inst_cell_78_26 (.BL(BL26),.BLN(BLN26),.WL(WL78));
sram_cell_6t_5 inst_cell_78_27 (.BL(BL27),.BLN(BLN27),.WL(WL78));
sram_cell_6t_5 inst_cell_78_28 (.BL(BL28),.BLN(BLN28),.WL(WL78));
sram_cell_6t_5 inst_cell_78_29 (.BL(BL29),.BLN(BLN29),.WL(WL78));
sram_cell_6t_5 inst_cell_78_30 (.BL(BL30),.BLN(BLN30),.WL(WL78));
sram_cell_6t_5 inst_cell_78_31 (.BL(BL31),.BLN(BLN31),.WL(WL78));
sram_cell_6t_5 inst_cell_78_32 (.BL(BL32),.BLN(BLN32),.WL(WL78));
sram_cell_6t_5 inst_cell_78_33 (.BL(BL33),.BLN(BLN33),.WL(WL78));
sram_cell_6t_5 inst_cell_78_34 (.BL(BL34),.BLN(BLN34),.WL(WL78));
sram_cell_6t_5 inst_cell_78_35 (.BL(BL35),.BLN(BLN35),.WL(WL78));
sram_cell_6t_5 inst_cell_78_36 (.BL(BL36),.BLN(BLN36),.WL(WL78));
sram_cell_6t_5 inst_cell_78_37 (.BL(BL37),.BLN(BLN37),.WL(WL78));
sram_cell_6t_5 inst_cell_78_38 (.BL(BL38),.BLN(BLN38),.WL(WL78));
sram_cell_6t_5 inst_cell_78_39 (.BL(BL39),.BLN(BLN39),.WL(WL78));
sram_cell_6t_5 inst_cell_78_40 (.BL(BL40),.BLN(BLN40),.WL(WL78));
sram_cell_6t_5 inst_cell_78_41 (.BL(BL41),.BLN(BLN41),.WL(WL78));
sram_cell_6t_5 inst_cell_78_42 (.BL(BL42),.BLN(BLN42),.WL(WL78));
sram_cell_6t_5 inst_cell_78_43 (.BL(BL43),.BLN(BLN43),.WL(WL78));
sram_cell_6t_5 inst_cell_78_44 (.BL(BL44),.BLN(BLN44),.WL(WL78));
sram_cell_6t_5 inst_cell_78_45 (.BL(BL45),.BLN(BLN45),.WL(WL78));
sram_cell_6t_5 inst_cell_78_46 (.BL(BL46),.BLN(BLN46),.WL(WL78));
sram_cell_6t_5 inst_cell_78_47 (.BL(BL47),.BLN(BLN47),.WL(WL78));
sram_cell_6t_5 inst_cell_78_48 (.BL(BL48),.BLN(BLN48),.WL(WL78));
sram_cell_6t_5 inst_cell_78_49 (.BL(BL49),.BLN(BLN49),.WL(WL78));
sram_cell_6t_5 inst_cell_78_50 (.BL(BL50),.BLN(BLN50),.WL(WL78));
sram_cell_6t_5 inst_cell_78_51 (.BL(BL51),.BLN(BLN51),.WL(WL78));
sram_cell_6t_5 inst_cell_78_52 (.BL(BL52),.BLN(BLN52),.WL(WL78));
sram_cell_6t_5 inst_cell_78_53 (.BL(BL53),.BLN(BLN53),.WL(WL78));
sram_cell_6t_5 inst_cell_78_54 (.BL(BL54),.BLN(BLN54),.WL(WL78));
sram_cell_6t_5 inst_cell_78_55 (.BL(BL55),.BLN(BLN55),.WL(WL78));
sram_cell_6t_5 inst_cell_78_56 (.BL(BL56),.BLN(BLN56),.WL(WL78));
sram_cell_6t_5 inst_cell_78_57 (.BL(BL57),.BLN(BLN57),.WL(WL78));
sram_cell_6t_5 inst_cell_78_58 (.BL(BL58),.BLN(BLN58),.WL(WL78));
sram_cell_6t_5 inst_cell_78_59 (.BL(BL59),.BLN(BLN59),.WL(WL78));
sram_cell_6t_5 inst_cell_78_60 (.BL(BL60),.BLN(BLN60),.WL(WL78));
sram_cell_6t_5 inst_cell_78_61 (.BL(BL61),.BLN(BLN61),.WL(WL78));
sram_cell_6t_5 inst_cell_78_62 (.BL(BL62),.BLN(BLN62),.WL(WL78));
sram_cell_6t_5 inst_cell_78_63 (.BL(BL63),.BLN(BLN63),.WL(WL78));
sram_cell_6t_5 inst_cell_78_64 (.BL(BL64),.BLN(BLN64),.WL(WL78));
sram_cell_6t_5 inst_cell_78_65 (.BL(BL65),.BLN(BLN65),.WL(WL78));
sram_cell_6t_5 inst_cell_78_66 (.BL(BL66),.BLN(BLN66),.WL(WL78));
sram_cell_6t_5 inst_cell_78_67 (.BL(BL67),.BLN(BLN67),.WL(WL78));
sram_cell_6t_5 inst_cell_78_68 (.BL(BL68),.BLN(BLN68),.WL(WL78));
sram_cell_6t_5 inst_cell_78_69 (.BL(BL69),.BLN(BLN69),.WL(WL78));
sram_cell_6t_5 inst_cell_78_70 (.BL(BL70),.BLN(BLN70),.WL(WL78));
sram_cell_6t_5 inst_cell_78_71 (.BL(BL71),.BLN(BLN71),.WL(WL78));
sram_cell_6t_5 inst_cell_78_72 (.BL(BL72),.BLN(BLN72),.WL(WL78));
sram_cell_6t_5 inst_cell_78_73 (.BL(BL73),.BLN(BLN73),.WL(WL78));
sram_cell_6t_5 inst_cell_78_74 (.BL(BL74),.BLN(BLN74),.WL(WL78));
sram_cell_6t_5 inst_cell_78_75 (.BL(BL75),.BLN(BLN75),.WL(WL78));
sram_cell_6t_5 inst_cell_78_76 (.BL(BL76),.BLN(BLN76),.WL(WL78));
sram_cell_6t_5 inst_cell_78_77 (.BL(BL77),.BLN(BLN77),.WL(WL78));
sram_cell_6t_5 inst_cell_78_78 (.BL(BL78),.BLN(BLN78),.WL(WL78));
sram_cell_6t_5 inst_cell_78_79 (.BL(BL79),.BLN(BLN79),.WL(WL78));
sram_cell_6t_5 inst_cell_78_80 (.BL(BL80),.BLN(BLN80),.WL(WL78));
sram_cell_6t_5 inst_cell_78_81 (.BL(BL81),.BLN(BLN81),.WL(WL78));
sram_cell_6t_5 inst_cell_78_82 (.BL(BL82),.BLN(BLN82),.WL(WL78));
sram_cell_6t_5 inst_cell_78_83 (.BL(BL83),.BLN(BLN83),.WL(WL78));
sram_cell_6t_5 inst_cell_78_84 (.BL(BL84),.BLN(BLN84),.WL(WL78));
sram_cell_6t_5 inst_cell_78_85 (.BL(BL85),.BLN(BLN85),.WL(WL78));
sram_cell_6t_5 inst_cell_78_86 (.BL(BL86),.BLN(BLN86),.WL(WL78));
sram_cell_6t_5 inst_cell_78_87 (.BL(BL87),.BLN(BLN87),.WL(WL78));
sram_cell_6t_5 inst_cell_78_88 (.BL(BL88),.BLN(BLN88),.WL(WL78));
sram_cell_6t_5 inst_cell_78_89 (.BL(BL89),.BLN(BLN89),.WL(WL78));
sram_cell_6t_5 inst_cell_78_90 (.BL(BL90),.BLN(BLN90),.WL(WL78));
sram_cell_6t_5 inst_cell_78_91 (.BL(BL91),.BLN(BLN91),.WL(WL78));
sram_cell_6t_5 inst_cell_78_92 (.BL(BL92),.BLN(BLN92),.WL(WL78));
sram_cell_6t_5 inst_cell_78_93 (.BL(BL93),.BLN(BLN93),.WL(WL78));
sram_cell_6t_5 inst_cell_78_94 (.BL(BL94),.BLN(BLN94),.WL(WL78));
sram_cell_6t_5 inst_cell_78_95 (.BL(BL95),.BLN(BLN95),.WL(WL78));
sram_cell_6t_5 inst_cell_78_96 (.BL(BL96),.BLN(BLN96),.WL(WL78));
sram_cell_6t_5 inst_cell_78_97 (.BL(BL97),.BLN(BLN97),.WL(WL78));
sram_cell_6t_5 inst_cell_78_98 (.BL(BL98),.BLN(BLN98),.WL(WL78));
sram_cell_6t_5 inst_cell_78_99 (.BL(BL99),.BLN(BLN99),.WL(WL78));
sram_cell_6t_5 inst_cell_78_100 (.BL(BL100),.BLN(BLN100),.WL(WL78));
sram_cell_6t_5 inst_cell_78_101 (.BL(BL101),.BLN(BLN101),.WL(WL78));
sram_cell_6t_5 inst_cell_78_102 (.BL(BL102),.BLN(BLN102),.WL(WL78));
sram_cell_6t_5 inst_cell_78_103 (.BL(BL103),.BLN(BLN103),.WL(WL78));
sram_cell_6t_5 inst_cell_78_104 (.BL(BL104),.BLN(BLN104),.WL(WL78));
sram_cell_6t_5 inst_cell_78_105 (.BL(BL105),.BLN(BLN105),.WL(WL78));
sram_cell_6t_5 inst_cell_78_106 (.BL(BL106),.BLN(BLN106),.WL(WL78));
sram_cell_6t_5 inst_cell_78_107 (.BL(BL107),.BLN(BLN107),.WL(WL78));
sram_cell_6t_5 inst_cell_78_108 (.BL(BL108),.BLN(BLN108),.WL(WL78));
sram_cell_6t_5 inst_cell_78_109 (.BL(BL109),.BLN(BLN109),.WL(WL78));
sram_cell_6t_5 inst_cell_78_110 (.BL(BL110),.BLN(BLN110),.WL(WL78));
sram_cell_6t_5 inst_cell_78_111 (.BL(BL111),.BLN(BLN111),.WL(WL78));
sram_cell_6t_5 inst_cell_78_112 (.BL(BL112),.BLN(BLN112),.WL(WL78));
sram_cell_6t_5 inst_cell_78_113 (.BL(BL113),.BLN(BLN113),.WL(WL78));
sram_cell_6t_5 inst_cell_78_114 (.BL(BL114),.BLN(BLN114),.WL(WL78));
sram_cell_6t_5 inst_cell_78_115 (.BL(BL115),.BLN(BLN115),.WL(WL78));
sram_cell_6t_5 inst_cell_78_116 (.BL(BL116),.BLN(BLN116),.WL(WL78));
sram_cell_6t_5 inst_cell_78_117 (.BL(BL117),.BLN(BLN117),.WL(WL78));
sram_cell_6t_5 inst_cell_78_118 (.BL(BL118),.BLN(BLN118),.WL(WL78));
sram_cell_6t_5 inst_cell_78_119 (.BL(BL119),.BLN(BLN119),.WL(WL78));
sram_cell_6t_5 inst_cell_78_120 (.BL(BL120),.BLN(BLN120),.WL(WL78));
sram_cell_6t_5 inst_cell_78_121 (.BL(BL121),.BLN(BLN121),.WL(WL78));
sram_cell_6t_5 inst_cell_78_122 (.BL(BL122),.BLN(BLN122),.WL(WL78));
sram_cell_6t_5 inst_cell_78_123 (.BL(BL123),.BLN(BLN123),.WL(WL78));
sram_cell_6t_5 inst_cell_78_124 (.BL(BL124),.BLN(BLN124),.WL(WL78));
sram_cell_6t_5 inst_cell_78_125 (.BL(BL125),.BLN(BLN125),.WL(WL78));
sram_cell_6t_5 inst_cell_78_126 (.BL(BL126),.BLN(BLN126),.WL(WL78));
sram_cell_6t_5 inst_cell_78_127 (.BL(BL127),.BLN(BLN127),.WL(WL78));
sram_cell_6t_5 inst_cell_79_0 (.BL(BL0),.BLN(BLN0),.WL(WL79));
sram_cell_6t_5 inst_cell_79_1 (.BL(BL1),.BLN(BLN1),.WL(WL79));
sram_cell_6t_5 inst_cell_79_2 (.BL(BL2),.BLN(BLN2),.WL(WL79));
sram_cell_6t_5 inst_cell_79_3 (.BL(BL3),.BLN(BLN3),.WL(WL79));
sram_cell_6t_5 inst_cell_79_4 (.BL(BL4),.BLN(BLN4),.WL(WL79));
sram_cell_6t_5 inst_cell_79_5 (.BL(BL5),.BLN(BLN5),.WL(WL79));
sram_cell_6t_5 inst_cell_79_6 (.BL(BL6),.BLN(BLN6),.WL(WL79));
sram_cell_6t_5 inst_cell_79_7 (.BL(BL7),.BLN(BLN7),.WL(WL79));
sram_cell_6t_5 inst_cell_79_8 (.BL(BL8),.BLN(BLN8),.WL(WL79));
sram_cell_6t_5 inst_cell_79_9 (.BL(BL9),.BLN(BLN9),.WL(WL79));
sram_cell_6t_5 inst_cell_79_10 (.BL(BL10),.BLN(BLN10),.WL(WL79));
sram_cell_6t_5 inst_cell_79_11 (.BL(BL11),.BLN(BLN11),.WL(WL79));
sram_cell_6t_5 inst_cell_79_12 (.BL(BL12),.BLN(BLN12),.WL(WL79));
sram_cell_6t_5 inst_cell_79_13 (.BL(BL13),.BLN(BLN13),.WL(WL79));
sram_cell_6t_5 inst_cell_79_14 (.BL(BL14),.BLN(BLN14),.WL(WL79));
sram_cell_6t_5 inst_cell_79_15 (.BL(BL15),.BLN(BLN15),.WL(WL79));
sram_cell_6t_5 inst_cell_79_16 (.BL(BL16),.BLN(BLN16),.WL(WL79));
sram_cell_6t_5 inst_cell_79_17 (.BL(BL17),.BLN(BLN17),.WL(WL79));
sram_cell_6t_5 inst_cell_79_18 (.BL(BL18),.BLN(BLN18),.WL(WL79));
sram_cell_6t_5 inst_cell_79_19 (.BL(BL19),.BLN(BLN19),.WL(WL79));
sram_cell_6t_5 inst_cell_79_20 (.BL(BL20),.BLN(BLN20),.WL(WL79));
sram_cell_6t_5 inst_cell_79_21 (.BL(BL21),.BLN(BLN21),.WL(WL79));
sram_cell_6t_5 inst_cell_79_22 (.BL(BL22),.BLN(BLN22),.WL(WL79));
sram_cell_6t_5 inst_cell_79_23 (.BL(BL23),.BLN(BLN23),.WL(WL79));
sram_cell_6t_5 inst_cell_79_24 (.BL(BL24),.BLN(BLN24),.WL(WL79));
sram_cell_6t_5 inst_cell_79_25 (.BL(BL25),.BLN(BLN25),.WL(WL79));
sram_cell_6t_5 inst_cell_79_26 (.BL(BL26),.BLN(BLN26),.WL(WL79));
sram_cell_6t_5 inst_cell_79_27 (.BL(BL27),.BLN(BLN27),.WL(WL79));
sram_cell_6t_5 inst_cell_79_28 (.BL(BL28),.BLN(BLN28),.WL(WL79));
sram_cell_6t_5 inst_cell_79_29 (.BL(BL29),.BLN(BLN29),.WL(WL79));
sram_cell_6t_5 inst_cell_79_30 (.BL(BL30),.BLN(BLN30),.WL(WL79));
sram_cell_6t_5 inst_cell_79_31 (.BL(BL31),.BLN(BLN31),.WL(WL79));
sram_cell_6t_5 inst_cell_79_32 (.BL(BL32),.BLN(BLN32),.WL(WL79));
sram_cell_6t_5 inst_cell_79_33 (.BL(BL33),.BLN(BLN33),.WL(WL79));
sram_cell_6t_5 inst_cell_79_34 (.BL(BL34),.BLN(BLN34),.WL(WL79));
sram_cell_6t_5 inst_cell_79_35 (.BL(BL35),.BLN(BLN35),.WL(WL79));
sram_cell_6t_5 inst_cell_79_36 (.BL(BL36),.BLN(BLN36),.WL(WL79));
sram_cell_6t_5 inst_cell_79_37 (.BL(BL37),.BLN(BLN37),.WL(WL79));
sram_cell_6t_5 inst_cell_79_38 (.BL(BL38),.BLN(BLN38),.WL(WL79));
sram_cell_6t_5 inst_cell_79_39 (.BL(BL39),.BLN(BLN39),.WL(WL79));
sram_cell_6t_5 inst_cell_79_40 (.BL(BL40),.BLN(BLN40),.WL(WL79));
sram_cell_6t_5 inst_cell_79_41 (.BL(BL41),.BLN(BLN41),.WL(WL79));
sram_cell_6t_5 inst_cell_79_42 (.BL(BL42),.BLN(BLN42),.WL(WL79));
sram_cell_6t_5 inst_cell_79_43 (.BL(BL43),.BLN(BLN43),.WL(WL79));
sram_cell_6t_5 inst_cell_79_44 (.BL(BL44),.BLN(BLN44),.WL(WL79));
sram_cell_6t_5 inst_cell_79_45 (.BL(BL45),.BLN(BLN45),.WL(WL79));
sram_cell_6t_5 inst_cell_79_46 (.BL(BL46),.BLN(BLN46),.WL(WL79));
sram_cell_6t_5 inst_cell_79_47 (.BL(BL47),.BLN(BLN47),.WL(WL79));
sram_cell_6t_5 inst_cell_79_48 (.BL(BL48),.BLN(BLN48),.WL(WL79));
sram_cell_6t_5 inst_cell_79_49 (.BL(BL49),.BLN(BLN49),.WL(WL79));
sram_cell_6t_5 inst_cell_79_50 (.BL(BL50),.BLN(BLN50),.WL(WL79));
sram_cell_6t_5 inst_cell_79_51 (.BL(BL51),.BLN(BLN51),.WL(WL79));
sram_cell_6t_5 inst_cell_79_52 (.BL(BL52),.BLN(BLN52),.WL(WL79));
sram_cell_6t_5 inst_cell_79_53 (.BL(BL53),.BLN(BLN53),.WL(WL79));
sram_cell_6t_5 inst_cell_79_54 (.BL(BL54),.BLN(BLN54),.WL(WL79));
sram_cell_6t_5 inst_cell_79_55 (.BL(BL55),.BLN(BLN55),.WL(WL79));
sram_cell_6t_5 inst_cell_79_56 (.BL(BL56),.BLN(BLN56),.WL(WL79));
sram_cell_6t_5 inst_cell_79_57 (.BL(BL57),.BLN(BLN57),.WL(WL79));
sram_cell_6t_5 inst_cell_79_58 (.BL(BL58),.BLN(BLN58),.WL(WL79));
sram_cell_6t_5 inst_cell_79_59 (.BL(BL59),.BLN(BLN59),.WL(WL79));
sram_cell_6t_5 inst_cell_79_60 (.BL(BL60),.BLN(BLN60),.WL(WL79));
sram_cell_6t_5 inst_cell_79_61 (.BL(BL61),.BLN(BLN61),.WL(WL79));
sram_cell_6t_5 inst_cell_79_62 (.BL(BL62),.BLN(BLN62),.WL(WL79));
sram_cell_6t_5 inst_cell_79_63 (.BL(BL63),.BLN(BLN63),.WL(WL79));
sram_cell_6t_5 inst_cell_79_64 (.BL(BL64),.BLN(BLN64),.WL(WL79));
sram_cell_6t_5 inst_cell_79_65 (.BL(BL65),.BLN(BLN65),.WL(WL79));
sram_cell_6t_5 inst_cell_79_66 (.BL(BL66),.BLN(BLN66),.WL(WL79));
sram_cell_6t_5 inst_cell_79_67 (.BL(BL67),.BLN(BLN67),.WL(WL79));
sram_cell_6t_5 inst_cell_79_68 (.BL(BL68),.BLN(BLN68),.WL(WL79));
sram_cell_6t_5 inst_cell_79_69 (.BL(BL69),.BLN(BLN69),.WL(WL79));
sram_cell_6t_5 inst_cell_79_70 (.BL(BL70),.BLN(BLN70),.WL(WL79));
sram_cell_6t_5 inst_cell_79_71 (.BL(BL71),.BLN(BLN71),.WL(WL79));
sram_cell_6t_5 inst_cell_79_72 (.BL(BL72),.BLN(BLN72),.WL(WL79));
sram_cell_6t_5 inst_cell_79_73 (.BL(BL73),.BLN(BLN73),.WL(WL79));
sram_cell_6t_5 inst_cell_79_74 (.BL(BL74),.BLN(BLN74),.WL(WL79));
sram_cell_6t_5 inst_cell_79_75 (.BL(BL75),.BLN(BLN75),.WL(WL79));
sram_cell_6t_5 inst_cell_79_76 (.BL(BL76),.BLN(BLN76),.WL(WL79));
sram_cell_6t_5 inst_cell_79_77 (.BL(BL77),.BLN(BLN77),.WL(WL79));
sram_cell_6t_5 inst_cell_79_78 (.BL(BL78),.BLN(BLN78),.WL(WL79));
sram_cell_6t_5 inst_cell_79_79 (.BL(BL79),.BLN(BLN79),.WL(WL79));
sram_cell_6t_5 inst_cell_79_80 (.BL(BL80),.BLN(BLN80),.WL(WL79));
sram_cell_6t_5 inst_cell_79_81 (.BL(BL81),.BLN(BLN81),.WL(WL79));
sram_cell_6t_5 inst_cell_79_82 (.BL(BL82),.BLN(BLN82),.WL(WL79));
sram_cell_6t_5 inst_cell_79_83 (.BL(BL83),.BLN(BLN83),.WL(WL79));
sram_cell_6t_5 inst_cell_79_84 (.BL(BL84),.BLN(BLN84),.WL(WL79));
sram_cell_6t_5 inst_cell_79_85 (.BL(BL85),.BLN(BLN85),.WL(WL79));
sram_cell_6t_5 inst_cell_79_86 (.BL(BL86),.BLN(BLN86),.WL(WL79));
sram_cell_6t_5 inst_cell_79_87 (.BL(BL87),.BLN(BLN87),.WL(WL79));
sram_cell_6t_5 inst_cell_79_88 (.BL(BL88),.BLN(BLN88),.WL(WL79));
sram_cell_6t_5 inst_cell_79_89 (.BL(BL89),.BLN(BLN89),.WL(WL79));
sram_cell_6t_5 inst_cell_79_90 (.BL(BL90),.BLN(BLN90),.WL(WL79));
sram_cell_6t_5 inst_cell_79_91 (.BL(BL91),.BLN(BLN91),.WL(WL79));
sram_cell_6t_5 inst_cell_79_92 (.BL(BL92),.BLN(BLN92),.WL(WL79));
sram_cell_6t_5 inst_cell_79_93 (.BL(BL93),.BLN(BLN93),.WL(WL79));
sram_cell_6t_5 inst_cell_79_94 (.BL(BL94),.BLN(BLN94),.WL(WL79));
sram_cell_6t_5 inst_cell_79_95 (.BL(BL95),.BLN(BLN95),.WL(WL79));
sram_cell_6t_5 inst_cell_79_96 (.BL(BL96),.BLN(BLN96),.WL(WL79));
sram_cell_6t_5 inst_cell_79_97 (.BL(BL97),.BLN(BLN97),.WL(WL79));
sram_cell_6t_5 inst_cell_79_98 (.BL(BL98),.BLN(BLN98),.WL(WL79));
sram_cell_6t_5 inst_cell_79_99 (.BL(BL99),.BLN(BLN99),.WL(WL79));
sram_cell_6t_5 inst_cell_79_100 (.BL(BL100),.BLN(BLN100),.WL(WL79));
sram_cell_6t_5 inst_cell_79_101 (.BL(BL101),.BLN(BLN101),.WL(WL79));
sram_cell_6t_5 inst_cell_79_102 (.BL(BL102),.BLN(BLN102),.WL(WL79));
sram_cell_6t_5 inst_cell_79_103 (.BL(BL103),.BLN(BLN103),.WL(WL79));
sram_cell_6t_5 inst_cell_79_104 (.BL(BL104),.BLN(BLN104),.WL(WL79));
sram_cell_6t_5 inst_cell_79_105 (.BL(BL105),.BLN(BLN105),.WL(WL79));
sram_cell_6t_5 inst_cell_79_106 (.BL(BL106),.BLN(BLN106),.WL(WL79));
sram_cell_6t_5 inst_cell_79_107 (.BL(BL107),.BLN(BLN107),.WL(WL79));
sram_cell_6t_5 inst_cell_79_108 (.BL(BL108),.BLN(BLN108),.WL(WL79));
sram_cell_6t_5 inst_cell_79_109 (.BL(BL109),.BLN(BLN109),.WL(WL79));
sram_cell_6t_5 inst_cell_79_110 (.BL(BL110),.BLN(BLN110),.WL(WL79));
sram_cell_6t_5 inst_cell_79_111 (.BL(BL111),.BLN(BLN111),.WL(WL79));
sram_cell_6t_5 inst_cell_79_112 (.BL(BL112),.BLN(BLN112),.WL(WL79));
sram_cell_6t_5 inst_cell_79_113 (.BL(BL113),.BLN(BLN113),.WL(WL79));
sram_cell_6t_5 inst_cell_79_114 (.BL(BL114),.BLN(BLN114),.WL(WL79));
sram_cell_6t_5 inst_cell_79_115 (.BL(BL115),.BLN(BLN115),.WL(WL79));
sram_cell_6t_5 inst_cell_79_116 (.BL(BL116),.BLN(BLN116),.WL(WL79));
sram_cell_6t_5 inst_cell_79_117 (.BL(BL117),.BLN(BLN117),.WL(WL79));
sram_cell_6t_5 inst_cell_79_118 (.BL(BL118),.BLN(BLN118),.WL(WL79));
sram_cell_6t_5 inst_cell_79_119 (.BL(BL119),.BLN(BLN119),.WL(WL79));
sram_cell_6t_5 inst_cell_79_120 (.BL(BL120),.BLN(BLN120),.WL(WL79));
sram_cell_6t_5 inst_cell_79_121 (.BL(BL121),.BLN(BLN121),.WL(WL79));
sram_cell_6t_5 inst_cell_79_122 (.BL(BL122),.BLN(BLN122),.WL(WL79));
sram_cell_6t_5 inst_cell_79_123 (.BL(BL123),.BLN(BLN123),.WL(WL79));
sram_cell_6t_5 inst_cell_79_124 (.BL(BL124),.BLN(BLN124),.WL(WL79));
sram_cell_6t_5 inst_cell_79_125 (.BL(BL125),.BLN(BLN125),.WL(WL79));
sram_cell_6t_5 inst_cell_79_126 (.BL(BL126),.BLN(BLN126),.WL(WL79));
sram_cell_6t_5 inst_cell_79_127 (.BL(BL127),.BLN(BLN127),.WL(WL79));
sram_cell_6t_5 inst_cell_80_0 (.BL(BL0),.BLN(BLN0),.WL(WL80));
sram_cell_6t_5 inst_cell_80_1 (.BL(BL1),.BLN(BLN1),.WL(WL80));
sram_cell_6t_5 inst_cell_80_2 (.BL(BL2),.BLN(BLN2),.WL(WL80));
sram_cell_6t_5 inst_cell_80_3 (.BL(BL3),.BLN(BLN3),.WL(WL80));
sram_cell_6t_5 inst_cell_80_4 (.BL(BL4),.BLN(BLN4),.WL(WL80));
sram_cell_6t_5 inst_cell_80_5 (.BL(BL5),.BLN(BLN5),.WL(WL80));
sram_cell_6t_5 inst_cell_80_6 (.BL(BL6),.BLN(BLN6),.WL(WL80));
sram_cell_6t_5 inst_cell_80_7 (.BL(BL7),.BLN(BLN7),.WL(WL80));
sram_cell_6t_5 inst_cell_80_8 (.BL(BL8),.BLN(BLN8),.WL(WL80));
sram_cell_6t_5 inst_cell_80_9 (.BL(BL9),.BLN(BLN9),.WL(WL80));
sram_cell_6t_5 inst_cell_80_10 (.BL(BL10),.BLN(BLN10),.WL(WL80));
sram_cell_6t_5 inst_cell_80_11 (.BL(BL11),.BLN(BLN11),.WL(WL80));
sram_cell_6t_5 inst_cell_80_12 (.BL(BL12),.BLN(BLN12),.WL(WL80));
sram_cell_6t_5 inst_cell_80_13 (.BL(BL13),.BLN(BLN13),.WL(WL80));
sram_cell_6t_5 inst_cell_80_14 (.BL(BL14),.BLN(BLN14),.WL(WL80));
sram_cell_6t_5 inst_cell_80_15 (.BL(BL15),.BLN(BLN15),.WL(WL80));
sram_cell_6t_5 inst_cell_80_16 (.BL(BL16),.BLN(BLN16),.WL(WL80));
sram_cell_6t_5 inst_cell_80_17 (.BL(BL17),.BLN(BLN17),.WL(WL80));
sram_cell_6t_5 inst_cell_80_18 (.BL(BL18),.BLN(BLN18),.WL(WL80));
sram_cell_6t_5 inst_cell_80_19 (.BL(BL19),.BLN(BLN19),.WL(WL80));
sram_cell_6t_5 inst_cell_80_20 (.BL(BL20),.BLN(BLN20),.WL(WL80));
sram_cell_6t_5 inst_cell_80_21 (.BL(BL21),.BLN(BLN21),.WL(WL80));
sram_cell_6t_5 inst_cell_80_22 (.BL(BL22),.BLN(BLN22),.WL(WL80));
sram_cell_6t_5 inst_cell_80_23 (.BL(BL23),.BLN(BLN23),.WL(WL80));
sram_cell_6t_5 inst_cell_80_24 (.BL(BL24),.BLN(BLN24),.WL(WL80));
sram_cell_6t_5 inst_cell_80_25 (.BL(BL25),.BLN(BLN25),.WL(WL80));
sram_cell_6t_5 inst_cell_80_26 (.BL(BL26),.BLN(BLN26),.WL(WL80));
sram_cell_6t_5 inst_cell_80_27 (.BL(BL27),.BLN(BLN27),.WL(WL80));
sram_cell_6t_5 inst_cell_80_28 (.BL(BL28),.BLN(BLN28),.WL(WL80));
sram_cell_6t_5 inst_cell_80_29 (.BL(BL29),.BLN(BLN29),.WL(WL80));
sram_cell_6t_5 inst_cell_80_30 (.BL(BL30),.BLN(BLN30),.WL(WL80));
sram_cell_6t_5 inst_cell_80_31 (.BL(BL31),.BLN(BLN31),.WL(WL80));
sram_cell_6t_5 inst_cell_80_32 (.BL(BL32),.BLN(BLN32),.WL(WL80));
sram_cell_6t_5 inst_cell_80_33 (.BL(BL33),.BLN(BLN33),.WL(WL80));
sram_cell_6t_5 inst_cell_80_34 (.BL(BL34),.BLN(BLN34),.WL(WL80));
sram_cell_6t_5 inst_cell_80_35 (.BL(BL35),.BLN(BLN35),.WL(WL80));
sram_cell_6t_5 inst_cell_80_36 (.BL(BL36),.BLN(BLN36),.WL(WL80));
sram_cell_6t_5 inst_cell_80_37 (.BL(BL37),.BLN(BLN37),.WL(WL80));
sram_cell_6t_5 inst_cell_80_38 (.BL(BL38),.BLN(BLN38),.WL(WL80));
sram_cell_6t_5 inst_cell_80_39 (.BL(BL39),.BLN(BLN39),.WL(WL80));
sram_cell_6t_5 inst_cell_80_40 (.BL(BL40),.BLN(BLN40),.WL(WL80));
sram_cell_6t_5 inst_cell_80_41 (.BL(BL41),.BLN(BLN41),.WL(WL80));
sram_cell_6t_5 inst_cell_80_42 (.BL(BL42),.BLN(BLN42),.WL(WL80));
sram_cell_6t_5 inst_cell_80_43 (.BL(BL43),.BLN(BLN43),.WL(WL80));
sram_cell_6t_5 inst_cell_80_44 (.BL(BL44),.BLN(BLN44),.WL(WL80));
sram_cell_6t_5 inst_cell_80_45 (.BL(BL45),.BLN(BLN45),.WL(WL80));
sram_cell_6t_5 inst_cell_80_46 (.BL(BL46),.BLN(BLN46),.WL(WL80));
sram_cell_6t_5 inst_cell_80_47 (.BL(BL47),.BLN(BLN47),.WL(WL80));
sram_cell_6t_5 inst_cell_80_48 (.BL(BL48),.BLN(BLN48),.WL(WL80));
sram_cell_6t_5 inst_cell_80_49 (.BL(BL49),.BLN(BLN49),.WL(WL80));
sram_cell_6t_5 inst_cell_80_50 (.BL(BL50),.BLN(BLN50),.WL(WL80));
sram_cell_6t_5 inst_cell_80_51 (.BL(BL51),.BLN(BLN51),.WL(WL80));
sram_cell_6t_5 inst_cell_80_52 (.BL(BL52),.BLN(BLN52),.WL(WL80));
sram_cell_6t_5 inst_cell_80_53 (.BL(BL53),.BLN(BLN53),.WL(WL80));
sram_cell_6t_5 inst_cell_80_54 (.BL(BL54),.BLN(BLN54),.WL(WL80));
sram_cell_6t_5 inst_cell_80_55 (.BL(BL55),.BLN(BLN55),.WL(WL80));
sram_cell_6t_5 inst_cell_80_56 (.BL(BL56),.BLN(BLN56),.WL(WL80));
sram_cell_6t_5 inst_cell_80_57 (.BL(BL57),.BLN(BLN57),.WL(WL80));
sram_cell_6t_5 inst_cell_80_58 (.BL(BL58),.BLN(BLN58),.WL(WL80));
sram_cell_6t_5 inst_cell_80_59 (.BL(BL59),.BLN(BLN59),.WL(WL80));
sram_cell_6t_5 inst_cell_80_60 (.BL(BL60),.BLN(BLN60),.WL(WL80));
sram_cell_6t_5 inst_cell_80_61 (.BL(BL61),.BLN(BLN61),.WL(WL80));
sram_cell_6t_5 inst_cell_80_62 (.BL(BL62),.BLN(BLN62),.WL(WL80));
sram_cell_6t_5 inst_cell_80_63 (.BL(BL63),.BLN(BLN63),.WL(WL80));
sram_cell_6t_5 inst_cell_80_64 (.BL(BL64),.BLN(BLN64),.WL(WL80));
sram_cell_6t_5 inst_cell_80_65 (.BL(BL65),.BLN(BLN65),.WL(WL80));
sram_cell_6t_5 inst_cell_80_66 (.BL(BL66),.BLN(BLN66),.WL(WL80));
sram_cell_6t_5 inst_cell_80_67 (.BL(BL67),.BLN(BLN67),.WL(WL80));
sram_cell_6t_5 inst_cell_80_68 (.BL(BL68),.BLN(BLN68),.WL(WL80));
sram_cell_6t_5 inst_cell_80_69 (.BL(BL69),.BLN(BLN69),.WL(WL80));
sram_cell_6t_5 inst_cell_80_70 (.BL(BL70),.BLN(BLN70),.WL(WL80));
sram_cell_6t_5 inst_cell_80_71 (.BL(BL71),.BLN(BLN71),.WL(WL80));
sram_cell_6t_5 inst_cell_80_72 (.BL(BL72),.BLN(BLN72),.WL(WL80));
sram_cell_6t_5 inst_cell_80_73 (.BL(BL73),.BLN(BLN73),.WL(WL80));
sram_cell_6t_5 inst_cell_80_74 (.BL(BL74),.BLN(BLN74),.WL(WL80));
sram_cell_6t_5 inst_cell_80_75 (.BL(BL75),.BLN(BLN75),.WL(WL80));
sram_cell_6t_5 inst_cell_80_76 (.BL(BL76),.BLN(BLN76),.WL(WL80));
sram_cell_6t_5 inst_cell_80_77 (.BL(BL77),.BLN(BLN77),.WL(WL80));
sram_cell_6t_5 inst_cell_80_78 (.BL(BL78),.BLN(BLN78),.WL(WL80));
sram_cell_6t_5 inst_cell_80_79 (.BL(BL79),.BLN(BLN79),.WL(WL80));
sram_cell_6t_5 inst_cell_80_80 (.BL(BL80),.BLN(BLN80),.WL(WL80));
sram_cell_6t_5 inst_cell_80_81 (.BL(BL81),.BLN(BLN81),.WL(WL80));
sram_cell_6t_5 inst_cell_80_82 (.BL(BL82),.BLN(BLN82),.WL(WL80));
sram_cell_6t_5 inst_cell_80_83 (.BL(BL83),.BLN(BLN83),.WL(WL80));
sram_cell_6t_5 inst_cell_80_84 (.BL(BL84),.BLN(BLN84),.WL(WL80));
sram_cell_6t_5 inst_cell_80_85 (.BL(BL85),.BLN(BLN85),.WL(WL80));
sram_cell_6t_5 inst_cell_80_86 (.BL(BL86),.BLN(BLN86),.WL(WL80));
sram_cell_6t_5 inst_cell_80_87 (.BL(BL87),.BLN(BLN87),.WL(WL80));
sram_cell_6t_5 inst_cell_80_88 (.BL(BL88),.BLN(BLN88),.WL(WL80));
sram_cell_6t_5 inst_cell_80_89 (.BL(BL89),.BLN(BLN89),.WL(WL80));
sram_cell_6t_5 inst_cell_80_90 (.BL(BL90),.BLN(BLN90),.WL(WL80));
sram_cell_6t_5 inst_cell_80_91 (.BL(BL91),.BLN(BLN91),.WL(WL80));
sram_cell_6t_5 inst_cell_80_92 (.BL(BL92),.BLN(BLN92),.WL(WL80));
sram_cell_6t_5 inst_cell_80_93 (.BL(BL93),.BLN(BLN93),.WL(WL80));
sram_cell_6t_5 inst_cell_80_94 (.BL(BL94),.BLN(BLN94),.WL(WL80));
sram_cell_6t_5 inst_cell_80_95 (.BL(BL95),.BLN(BLN95),.WL(WL80));
sram_cell_6t_5 inst_cell_80_96 (.BL(BL96),.BLN(BLN96),.WL(WL80));
sram_cell_6t_5 inst_cell_80_97 (.BL(BL97),.BLN(BLN97),.WL(WL80));
sram_cell_6t_5 inst_cell_80_98 (.BL(BL98),.BLN(BLN98),.WL(WL80));
sram_cell_6t_5 inst_cell_80_99 (.BL(BL99),.BLN(BLN99),.WL(WL80));
sram_cell_6t_5 inst_cell_80_100 (.BL(BL100),.BLN(BLN100),.WL(WL80));
sram_cell_6t_5 inst_cell_80_101 (.BL(BL101),.BLN(BLN101),.WL(WL80));
sram_cell_6t_5 inst_cell_80_102 (.BL(BL102),.BLN(BLN102),.WL(WL80));
sram_cell_6t_5 inst_cell_80_103 (.BL(BL103),.BLN(BLN103),.WL(WL80));
sram_cell_6t_5 inst_cell_80_104 (.BL(BL104),.BLN(BLN104),.WL(WL80));
sram_cell_6t_5 inst_cell_80_105 (.BL(BL105),.BLN(BLN105),.WL(WL80));
sram_cell_6t_5 inst_cell_80_106 (.BL(BL106),.BLN(BLN106),.WL(WL80));
sram_cell_6t_5 inst_cell_80_107 (.BL(BL107),.BLN(BLN107),.WL(WL80));
sram_cell_6t_5 inst_cell_80_108 (.BL(BL108),.BLN(BLN108),.WL(WL80));
sram_cell_6t_5 inst_cell_80_109 (.BL(BL109),.BLN(BLN109),.WL(WL80));
sram_cell_6t_5 inst_cell_80_110 (.BL(BL110),.BLN(BLN110),.WL(WL80));
sram_cell_6t_5 inst_cell_80_111 (.BL(BL111),.BLN(BLN111),.WL(WL80));
sram_cell_6t_5 inst_cell_80_112 (.BL(BL112),.BLN(BLN112),.WL(WL80));
sram_cell_6t_5 inst_cell_80_113 (.BL(BL113),.BLN(BLN113),.WL(WL80));
sram_cell_6t_5 inst_cell_80_114 (.BL(BL114),.BLN(BLN114),.WL(WL80));
sram_cell_6t_5 inst_cell_80_115 (.BL(BL115),.BLN(BLN115),.WL(WL80));
sram_cell_6t_5 inst_cell_80_116 (.BL(BL116),.BLN(BLN116),.WL(WL80));
sram_cell_6t_5 inst_cell_80_117 (.BL(BL117),.BLN(BLN117),.WL(WL80));
sram_cell_6t_5 inst_cell_80_118 (.BL(BL118),.BLN(BLN118),.WL(WL80));
sram_cell_6t_5 inst_cell_80_119 (.BL(BL119),.BLN(BLN119),.WL(WL80));
sram_cell_6t_5 inst_cell_80_120 (.BL(BL120),.BLN(BLN120),.WL(WL80));
sram_cell_6t_5 inst_cell_80_121 (.BL(BL121),.BLN(BLN121),.WL(WL80));
sram_cell_6t_5 inst_cell_80_122 (.BL(BL122),.BLN(BLN122),.WL(WL80));
sram_cell_6t_5 inst_cell_80_123 (.BL(BL123),.BLN(BLN123),.WL(WL80));
sram_cell_6t_5 inst_cell_80_124 (.BL(BL124),.BLN(BLN124),.WL(WL80));
sram_cell_6t_5 inst_cell_80_125 (.BL(BL125),.BLN(BLN125),.WL(WL80));
sram_cell_6t_5 inst_cell_80_126 (.BL(BL126),.BLN(BLN126),.WL(WL80));
sram_cell_6t_5 inst_cell_80_127 (.BL(BL127),.BLN(BLN127),.WL(WL80));
sram_cell_6t_5 inst_cell_81_0 (.BL(BL0),.BLN(BLN0),.WL(WL81));
sram_cell_6t_5 inst_cell_81_1 (.BL(BL1),.BLN(BLN1),.WL(WL81));
sram_cell_6t_5 inst_cell_81_2 (.BL(BL2),.BLN(BLN2),.WL(WL81));
sram_cell_6t_5 inst_cell_81_3 (.BL(BL3),.BLN(BLN3),.WL(WL81));
sram_cell_6t_5 inst_cell_81_4 (.BL(BL4),.BLN(BLN4),.WL(WL81));
sram_cell_6t_5 inst_cell_81_5 (.BL(BL5),.BLN(BLN5),.WL(WL81));
sram_cell_6t_5 inst_cell_81_6 (.BL(BL6),.BLN(BLN6),.WL(WL81));
sram_cell_6t_5 inst_cell_81_7 (.BL(BL7),.BLN(BLN7),.WL(WL81));
sram_cell_6t_5 inst_cell_81_8 (.BL(BL8),.BLN(BLN8),.WL(WL81));
sram_cell_6t_5 inst_cell_81_9 (.BL(BL9),.BLN(BLN9),.WL(WL81));
sram_cell_6t_5 inst_cell_81_10 (.BL(BL10),.BLN(BLN10),.WL(WL81));
sram_cell_6t_5 inst_cell_81_11 (.BL(BL11),.BLN(BLN11),.WL(WL81));
sram_cell_6t_5 inst_cell_81_12 (.BL(BL12),.BLN(BLN12),.WL(WL81));
sram_cell_6t_5 inst_cell_81_13 (.BL(BL13),.BLN(BLN13),.WL(WL81));
sram_cell_6t_5 inst_cell_81_14 (.BL(BL14),.BLN(BLN14),.WL(WL81));
sram_cell_6t_5 inst_cell_81_15 (.BL(BL15),.BLN(BLN15),.WL(WL81));
sram_cell_6t_5 inst_cell_81_16 (.BL(BL16),.BLN(BLN16),.WL(WL81));
sram_cell_6t_5 inst_cell_81_17 (.BL(BL17),.BLN(BLN17),.WL(WL81));
sram_cell_6t_5 inst_cell_81_18 (.BL(BL18),.BLN(BLN18),.WL(WL81));
sram_cell_6t_5 inst_cell_81_19 (.BL(BL19),.BLN(BLN19),.WL(WL81));
sram_cell_6t_5 inst_cell_81_20 (.BL(BL20),.BLN(BLN20),.WL(WL81));
sram_cell_6t_5 inst_cell_81_21 (.BL(BL21),.BLN(BLN21),.WL(WL81));
sram_cell_6t_5 inst_cell_81_22 (.BL(BL22),.BLN(BLN22),.WL(WL81));
sram_cell_6t_5 inst_cell_81_23 (.BL(BL23),.BLN(BLN23),.WL(WL81));
sram_cell_6t_5 inst_cell_81_24 (.BL(BL24),.BLN(BLN24),.WL(WL81));
sram_cell_6t_5 inst_cell_81_25 (.BL(BL25),.BLN(BLN25),.WL(WL81));
sram_cell_6t_5 inst_cell_81_26 (.BL(BL26),.BLN(BLN26),.WL(WL81));
sram_cell_6t_5 inst_cell_81_27 (.BL(BL27),.BLN(BLN27),.WL(WL81));
sram_cell_6t_5 inst_cell_81_28 (.BL(BL28),.BLN(BLN28),.WL(WL81));
sram_cell_6t_5 inst_cell_81_29 (.BL(BL29),.BLN(BLN29),.WL(WL81));
sram_cell_6t_5 inst_cell_81_30 (.BL(BL30),.BLN(BLN30),.WL(WL81));
sram_cell_6t_5 inst_cell_81_31 (.BL(BL31),.BLN(BLN31),.WL(WL81));
sram_cell_6t_5 inst_cell_81_32 (.BL(BL32),.BLN(BLN32),.WL(WL81));
sram_cell_6t_5 inst_cell_81_33 (.BL(BL33),.BLN(BLN33),.WL(WL81));
sram_cell_6t_5 inst_cell_81_34 (.BL(BL34),.BLN(BLN34),.WL(WL81));
sram_cell_6t_5 inst_cell_81_35 (.BL(BL35),.BLN(BLN35),.WL(WL81));
sram_cell_6t_5 inst_cell_81_36 (.BL(BL36),.BLN(BLN36),.WL(WL81));
sram_cell_6t_5 inst_cell_81_37 (.BL(BL37),.BLN(BLN37),.WL(WL81));
sram_cell_6t_5 inst_cell_81_38 (.BL(BL38),.BLN(BLN38),.WL(WL81));
sram_cell_6t_5 inst_cell_81_39 (.BL(BL39),.BLN(BLN39),.WL(WL81));
sram_cell_6t_5 inst_cell_81_40 (.BL(BL40),.BLN(BLN40),.WL(WL81));
sram_cell_6t_5 inst_cell_81_41 (.BL(BL41),.BLN(BLN41),.WL(WL81));
sram_cell_6t_5 inst_cell_81_42 (.BL(BL42),.BLN(BLN42),.WL(WL81));
sram_cell_6t_5 inst_cell_81_43 (.BL(BL43),.BLN(BLN43),.WL(WL81));
sram_cell_6t_5 inst_cell_81_44 (.BL(BL44),.BLN(BLN44),.WL(WL81));
sram_cell_6t_5 inst_cell_81_45 (.BL(BL45),.BLN(BLN45),.WL(WL81));
sram_cell_6t_5 inst_cell_81_46 (.BL(BL46),.BLN(BLN46),.WL(WL81));
sram_cell_6t_5 inst_cell_81_47 (.BL(BL47),.BLN(BLN47),.WL(WL81));
sram_cell_6t_5 inst_cell_81_48 (.BL(BL48),.BLN(BLN48),.WL(WL81));
sram_cell_6t_5 inst_cell_81_49 (.BL(BL49),.BLN(BLN49),.WL(WL81));
sram_cell_6t_5 inst_cell_81_50 (.BL(BL50),.BLN(BLN50),.WL(WL81));
sram_cell_6t_5 inst_cell_81_51 (.BL(BL51),.BLN(BLN51),.WL(WL81));
sram_cell_6t_5 inst_cell_81_52 (.BL(BL52),.BLN(BLN52),.WL(WL81));
sram_cell_6t_5 inst_cell_81_53 (.BL(BL53),.BLN(BLN53),.WL(WL81));
sram_cell_6t_5 inst_cell_81_54 (.BL(BL54),.BLN(BLN54),.WL(WL81));
sram_cell_6t_5 inst_cell_81_55 (.BL(BL55),.BLN(BLN55),.WL(WL81));
sram_cell_6t_5 inst_cell_81_56 (.BL(BL56),.BLN(BLN56),.WL(WL81));
sram_cell_6t_5 inst_cell_81_57 (.BL(BL57),.BLN(BLN57),.WL(WL81));
sram_cell_6t_5 inst_cell_81_58 (.BL(BL58),.BLN(BLN58),.WL(WL81));
sram_cell_6t_5 inst_cell_81_59 (.BL(BL59),.BLN(BLN59),.WL(WL81));
sram_cell_6t_5 inst_cell_81_60 (.BL(BL60),.BLN(BLN60),.WL(WL81));
sram_cell_6t_5 inst_cell_81_61 (.BL(BL61),.BLN(BLN61),.WL(WL81));
sram_cell_6t_5 inst_cell_81_62 (.BL(BL62),.BLN(BLN62),.WL(WL81));
sram_cell_6t_5 inst_cell_81_63 (.BL(BL63),.BLN(BLN63),.WL(WL81));
sram_cell_6t_5 inst_cell_81_64 (.BL(BL64),.BLN(BLN64),.WL(WL81));
sram_cell_6t_5 inst_cell_81_65 (.BL(BL65),.BLN(BLN65),.WL(WL81));
sram_cell_6t_5 inst_cell_81_66 (.BL(BL66),.BLN(BLN66),.WL(WL81));
sram_cell_6t_5 inst_cell_81_67 (.BL(BL67),.BLN(BLN67),.WL(WL81));
sram_cell_6t_5 inst_cell_81_68 (.BL(BL68),.BLN(BLN68),.WL(WL81));
sram_cell_6t_5 inst_cell_81_69 (.BL(BL69),.BLN(BLN69),.WL(WL81));
sram_cell_6t_5 inst_cell_81_70 (.BL(BL70),.BLN(BLN70),.WL(WL81));
sram_cell_6t_5 inst_cell_81_71 (.BL(BL71),.BLN(BLN71),.WL(WL81));
sram_cell_6t_5 inst_cell_81_72 (.BL(BL72),.BLN(BLN72),.WL(WL81));
sram_cell_6t_5 inst_cell_81_73 (.BL(BL73),.BLN(BLN73),.WL(WL81));
sram_cell_6t_5 inst_cell_81_74 (.BL(BL74),.BLN(BLN74),.WL(WL81));
sram_cell_6t_5 inst_cell_81_75 (.BL(BL75),.BLN(BLN75),.WL(WL81));
sram_cell_6t_5 inst_cell_81_76 (.BL(BL76),.BLN(BLN76),.WL(WL81));
sram_cell_6t_5 inst_cell_81_77 (.BL(BL77),.BLN(BLN77),.WL(WL81));
sram_cell_6t_5 inst_cell_81_78 (.BL(BL78),.BLN(BLN78),.WL(WL81));
sram_cell_6t_5 inst_cell_81_79 (.BL(BL79),.BLN(BLN79),.WL(WL81));
sram_cell_6t_5 inst_cell_81_80 (.BL(BL80),.BLN(BLN80),.WL(WL81));
sram_cell_6t_5 inst_cell_81_81 (.BL(BL81),.BLN(BLN81),.WL(WL81));
sram_cell_6t_5 inst_cell_81_82 (.BL(BL82),.BLN(BLN82),.WL(WL81));
sram_cell_6t_5 inst_cell_81_83 (.BL(BL83),.BLN(BLN83),.WL(WL81));
sram_cell_6t_5 inst_cell_81_84 (.BL(BL84),.BLN(BLN84),.WL(WL81));
sram_cell_6t_5 inst_cell_81_85 (.BL(BL85),.BLN(BLN85),.WL(WL81));
sram_cell_6t_5 inst_cell_81_86 (.BL(BL86),.BLN(BLN86),.WL(WL81));
sram_cell_6t_5 inst_cell_81_87 (.BL(BL87),.BLN(BLN87),.WL(WL81));
sram_cell_6t_5 inst_cell_81_88 (.BL(BL88),.BLN(BLN88),.WL(WL81));
sram_cell_6t_5 inst_cell_81_89 (.BL(BL89),.BLN(BLN89),.WL(WL81));
sram_cell_6t_5 inst_cell_81_90 (.BL(BL90),.BLN(BLN90),.WL(WL81));
sram_cell_6t_5 inst_cell_81_91 (.BL(BL91),.BLN(BLN91),.WL(WL81));
sram_cell_6t_5 inst_cell_81_92 (.BL(BL92),.BLN(BLN92),.WL(WL81));
sram_cell_6t_5 inst_cell_81_93 (.BL(BL93),.BLN(BLN93),.WL(WL81));
sram_cell_6t_5 inst_cell_81_94 (.BL(BL94),.BLN(BLN94),.WL(WL81));
sram_cell_6t_5 inst_cell_81_95 (.BL(BL95),.BLN(BLN95),.WL(WL81));
sram_cell_6t_5 inst_cell_81_96 (.BL(BL96),.BLN(BLN96),.WL(WL81));
sram_cell_6t_5 inst_cell_81_97 (.BL(BL97),.BLN(BLN97),.WL(WL81));
sram_cell_6t_5 inst_cell_81_98 (.BL(BL98),.BLN(BLN98),.WL(WL81));
sram_cell_6t_5 inst_cell_81_99 (.BL(BL99),.BLN(BLN99),.WL(WL81));
sram_cell_6t_5 inst_cell_81_100 (.BL(BL100),.BLN(BLN100),.WL(WL81));
sram_cell_6t_5 inst_cell_81_101 (.BL(BL101),.BLN(BLN101),.WL(WL81));
sram_cell_6t_5 inst_cell_81_102 (.BL(BL102),.BLN(BLN102),.WL(WL81));
sram_cell_6t_5 inst_cell_81_103 (.BL(BL103),.BLN(BLN103),.WL(WL81));
sram_cell_6t_5 inst_cell_81_104 (.BL(BL104),.BLN(BLN104),.WL(WL81));
sram_cell_6t_5 inst_cell_81_105 (.BL(BL105),.BLN(BLN105),.WL(WL81));
sram_cell_6t_5 inst_cell_81_106 (.BL(BL106),.BLN(BLN106),.WL(WL81));
sram_cell_6t_5 inst_cell_81_107 (.BL(BL107),.BLN(BLN107),.WL(WL81));
sram_cell_6t_5 inst_cell_81_108 (.BL(BL108),.BLN(BLN108),.WL(WL81));
sram_cell_6t_5 inst_cell_81_109 (.BL(BL109),.BLN(BLN109),.WL(WL81));
sram_cell_6t_5 inst_cell_81_110 (.BL(BL110),.BLN(BLN110),.WL(WL81));
sram_cell_6t_5 inst_cell_81_111 (.BL(BL111),.BLN(BLN111),.WL(WL81));
sram_cell_6t_5 inst_cell_81_112 (.BL(BL112),.BLN(BLN112),.WL(WL81));
sram_cell_6t_5 inst_cell_81_113 (.BL(BL113),.BLN(BLN113),.WL(WL81));
sram_cell_6t_5 inst_cell_81_114 (.BL(BL114),.BLN(BLN114),.WL(WL81));
sram_cell_6t_5 inst_cell_81_115 (.BL(BL115),.BLN(BLN115),.WL(WL81));
sram_cell_6t_5 inst_cell_81_116 (.BL(BL116),.BLN(BLN116),.WL(WL81));
sram_cell_6t_5 inst_cell_81_117 (.BL(BL117),.BLN(BLN117),.WL(WL81));
sram_cell_6t_5 inst_cell_81_118 (.BL(BL118),.BLN(BLN118),.WL(WL81));
sram_cell_6t_5 inst_cell_81_119 (.BL(BL119),.BLN(BLN119),.WL(WL81));
sram_cell_6t_5 inst_cell_81_120 (.BL(BL120),.BLN(BLN120),.WL(WL81));
sram_cell_6t_5 inst_cell_81_121 (.BL(BL121),.BLN(BLN121),.WL(WL81));
sram_cell_6t_5 inst_cell_81_122 (.BL(BL122),.BLN(BLN122),.WL(WL81));
sram_cell_6t_5 inst_cell_81_123 (.BL(BL123),.BLN(BLN123),.WL(WL81));
sram_cell_6t_5 inst_cell_81_124 (.BL(BL124),.BLN(BLN124),.WL(WL81));
sram_cell_6t_5 inst_cell_81_125 (.BL(BL125),.BLN(BLN125),.WL(WL81));
sram_cell_6t_5 inst_cell_81_126 (.BL(BL126),.BLN(BLN126),.WL(WL81));
sram_cell_6t_5 inst_cell_81_127 (.BL(BL127),.BLN(BLN127),.WL(WL81));
sram_cell_6t_5 inst_cell_82_0 (.BL(BL0),.BLN(BLN0),.WL(WL82));
sram_cell_6t_5 inst_cell_82_1 (.BL(BL1),.BLN(BLN1),.WL(WL82));
sram_cell_6t_5 inst_cell_82_2 (.BL(BL2),.BLN(BLN2),.WL(WL82));
sram_cell_6t_5 inst_cell_82_3 (.BL(BL3),.BLN(BLN3),.WL(WL82));
sram_cell_6t_5 inst_cell_82_4 (.BL(BL4),.BLN(BLN4),.WL(WL82));
sram_cell_6t_5 inst_cell_82_5 (.BL(BL5),.BLN(BLN5),.WL(WL82));
sram_cell_6t_5 inst_cell_82_6 (.BL(BL6),.BLN(BLN6),.WL(WL82));
sram_cell_6t_5 inst_cell_82_7 (.BL(BL7),.BLN(BLN7),.WL(WL82));
sram_cell_6t_5 inst_cell_82_8 (.BL(BL8),.BLN(BLN8),.WL(WL82));
sram_cell_6t_5 inst_cell_82_9 (.BL(BL9),.BLN(BLN9),.WL(WL82));
sram_cell_6t_5 inst_cell_82_10 (.BL(BL10),.BLN(BLN10),.WL(WL82));
sram_cell_6t_5 inst_cell_82_11 (.BL(BL11),.BLN(BLN11),.WL(WL82));
sram_cell_6t_5 inst_cell_82_12 (.BL(BL12),.BLN(BLN12),.WL(WL82));
sram_cell_6t_5 inst_cell_82_13 (.BL(BL13),.BLN(BLN13),.WL(WL82));
sram_cell_6t_5 inst_cell_82_14 (.BL(BL14),.BLN(BLN14),.WL(WL82));
sram_cell_6t_5 inst_cell_82_15 (.BL(BL15),.BLN(BLN15),.WL(WL82));
sram_cell_6t_5 inst_cell_82_16 (.BL(BL16),.BLN(BLN16),.WL(WL82));
sram_cell_6t_5 inst_cell_82_17 (.BL(BL17),.BLN(BLN17),.WL(WL82));
sram_cell_6t_5 inst_cell_82_18 (.BL(BL18),.BLN(BLN18),.WL(WL82));
sram_cell_6t_5 inst_cell_82_19 (.BL(BL19),.BLN(BLN19),.WL(WL82));
sram_cell_6t_5 inst_cell_82_20 (.BL(BL20),.BLN(BLN20),.WL(WL82));
sram_cell_6t_5 inst_cell_82_21 (.BL(BL21),.BLN(BLN21),.WL(WL82));
sram_cell_6t_5 inst_cell_82_22 (.BL(BL22),.BLN(BLN22),.WL(WL82));
sram_cell_6t_5 inst_cell_82_23 (.BL(BL23),.BLN(BLN23),.WL(WL82));
sram_cell_6t_5 inst_cell_82_24 (.BL(BL24),.BLN(BLN24),.WL(WL82));
sram_cell_6t_5 inst_cell_82_25 (.BL(BL25),.BLN(BLN25),.WL(WL82));
sram_cell_6t_5 inst_cell_82_26 (.BL(BL26),.BLN(BLN26),.WL(WL82));
sram_cell_6t_5 inst_cell_82_27 (.BL(BL27),.BLN(BLN27),.WL(WL82));
sram_cell_6t_5 inst_cell_82_28 (.BL(BL28),.BLN(BLN28),.WL(WL82));
sram_cell_6t_5 inst_cell_82_29 (.BL(BL29),.BLN(BLN29),.WL(WL82));
sram_cell_6t_5 inst_cell_82_30 (.BL(BL30),.BLN(BLN30),.WL(WL82));
sram_cell_6t_5 inst_cell_82_31 (.BL(BL31),.BLN(BLN31),.WL(WL82));
sram_cell_6t_5 inst_cell_82_32 (.BL(BL32),.BLN(BLN32),.WL(WL82));
sram_cell_6t_5 inst_cell_82_33 (.BL(BL33),.BLN(BLN33),.WL(WL82));
sram_cell_6t_5 inst_cell_82_34 (.BL(BL34),.BLN(BLN34),.WL(WL82));
sram_cell_6t_5 inst_cell_82_35 (.BL(BL35),.BLN(BLN35),.WL(WL82));
sram_cell_6t_5 inst_cell_82_36 (.BL(BL36),.BLN(BLN36),.WL(WL82));
sram_cell_6t_5 inst_cell_82_37 (.BL(BL37),.BLN(BLN37),.WL(WL82));
sram_cell_6t_5 inst_cell_82_38 (.BL(BL38),.BLN(BLN38),.WL(WL82));
sram_cell_6t_5 inst_cell_82_39 (.BL(BL39),.BLN(BLN39),.WL(WL82));
sram_cell_6t_5 inst_cell_82_40 (.BL(BL40),.BLN(BLN40),.WL(WL82));
sram_cell_6t_5 inst_cell_82_41 (.BL(BL41),.BLN(BLN41),.WL(WL82));
sram_cell_6t_5 inst_cell_82_42 (.BL(BL42),.BLN(BLN42),.WL(WL82));
sram_cell_6t_5 inst_cell_82_43 (.BL(BL43),.BLN(BLN43),.WL(WL82));
sram_cell_6t_5 inst_cell_82_44 (.BL(BL44),.BLN(BLN44),.WL(WL82));
sram_cell_6t_5 inst_cell_82_45 (.BL(BL45),.BLN(BLN45),.WL(WL82));
sram_cell_6t_5 inst_cell_82_46 (.BL(BL46),.BLN(BLN46),.WL(WL82));
sram_cell_6t_5 inst_cell_82_47 (.BL(BL47),.BLN(BLN47),.WL(WL82));
sram_cell_6t_5 inst_cell_82_48 (.BL(BL48),.BLN(BLN48),.WL(WL82));
sram_cell_6t_5 inst_cell_82_49 (.BL(BL49),.BLN(BLN49),.WL(WL82));
sram_cell_6t_5 inst_cell_82_50 (.BL(BL50),.BLN(BLN50),.WL(WL82));
sram_cell_6t_5 inst_cell_82_51 (.BL(BL51),.BLN(BLN51),.WL(WL82));
sram_cell_6t_5 inst_cell_82_52 (.BL(BL52),.BLN(BLN52),.WL(WL82));
sram_cell_6t_5 inst_cell_82_53 (.BL(BL53),.BLN(BLN53),.WL(WL82));
sram_cell_6t_5 inst_cell_82_54 (.BL(BL54),.BLN(BLN54),.WL(WL82));
sram_cell_6t_5 inst_cell_82_55 (.BL(BL55),.BLN(BLN55),.WL(WL82));
sram_cell_6t_5 inst_cell_82_56 (.BL(BL56),.BLN(BLN56),.WL(WL82));
sram_cell_6t_5 inst_cell_82_57 (.BL(BL57),.BLN(BLN57),.WL(WL82));
sram_cell_6t_5 inst_cell_82_58 (.BL(BL58),.BLN(BLN58),.WL(WL82));
sram_cell_6t_5 inst_cell_82_59 (.BL(BL59),.BLN(BLN59),.WL(WL82));
sram_cell_6t_5 inst_cell_82_60 (.BL(BL60),.BLN(BLN60),.WL(WL82));
sram_cell_6t_5 inst_cell_82_61 (.BL(BL61),.BLN(BLN61),.WL(WL82));
sram_cell_6t_5 inst_cell_82_62 (.BL(BL62),.BLN(BLN62),.WL(WL82));
sram_cell_6t_5 inst_cell_82_63 (.BL(BL63),.BLN(BLN63),.WL(WL82));
sram_cell_6t_5 inst_cell_82_64 (.BL(BL64),.BLN(BLN64),.WL(WL82));
sram_cell_6t_5 inst_cell_82_65 (.BL(BL65),.BLN(BLN65),.WL(WL82));
sram_cell_6t_5 inst_cell_82_66 (.BL(BL66),.BLN(BLN66),.WL(WL82));
sram_cell_6t_5 inst_cell_82_67 (.BL(BL67),.BLN(BLN67),.WL(WL82));
sram_cell_6t_5 inst_cell_82_68 (.BL(BL68),.BLN(BLN68),.WL(WL82));
sram_cell_6t_5 inst_cell_82_69 (.BL(BL69),.BLN(BLN69),.WL(WL82));
sram_cell_6t_5 inst_cell_82_70 (.BL(BL70),.BLN(BLN70),.WL(WL82));
sram_cell_6t_5 inst_cell_82_71 (.BL(BL71),.BLN(BLN71),.WL(WL82));
sram_cell_6t_5 inst_cell_82_72 (.BL(BL72),.BLN(BLN72),.WL(WL82));
sram_cell_6t_5 inst_cell_82_73 (.BL(BL73),.BLN(BLN73),.WL(WL82));
sram_cell_6t_5 inst_cell_82_74 (.BL(BL74),.BLN(BLN74),.WL(WL82));
sram_cell_6t_5 inst_cell_82_75 (.BL(BL75),.BLN(BLN75),.WL(WL82));
sram_cell_6t_5 inst_cell_82_76 (.BL(BL76),.BLN(BLN76),.WL(WL82));
sram_cell_6t_5 inst_cell_82_77 (.BL(BL77),.BLN(BLN77),.WL(WL82));
sram_cell_6t_5 inst_cell_82_78 (.BL(BL78),.BLN(BLN78),.WL(WL82));
sram_cell_6t_5 inst_cell_82_79 (.BL(BL79),.BLN(BLN79),.WL(WL82));
sram_cell_6t_5 inst_cell_82_80 (.BL(BL80),.BLN(BLN80),.WL(WL82));
sram_cell_6t_5 inst_cell_82_81 (.BL(BL81),.BLN(BLN81),.WL(WL82));
sram_cell_6t_5 inst_cell_82_82 (.BL(BL82),.BLN(BLN82),.WL(WL82));
sram_cell_6t_5 inst_cell_82_83 (.BL(BL83),.BLN(BLN83),.WL(WL82));
sram_cell_6t_5 inst_cell_82_84 (.BL(BL84),.BLN(BLN84),.WL(WL82));
sram_cell_6t_5 inst_cell_82_85 (.BL(BL85),.BLN(BLN85),.WL(WL82));
sram_cell_6t_5 inst_cell_82_86 (.BL(BL86),.BLN(BLN86),.WL(WL82));
sram_cell_6t_5 inst_cell_82_87 (.BL(BL87),.BLN(BLN87),.WL(WL82));
sram_cell_6t_5 inst_cell_82_88 (.BL(BL88),.BLN(BLN88),.WL(WL82));
sram_cell_6t_5 inst_cell_82_89 (.BL(BL89),.BLN(BLN89),.WL(WL82));
sram_cell_6t_5 inst_cell_82_90 (.BL(BL90),.BLN(BLN90),.WL(WL82));
sram_cell_6t_5 inst_cell_82_91 (.BL(BL91),.BLN(BLN91),.WL(WL82));
sram_cell_6t_5 inst_cell_82_92 (.BL(BL92),.BLN(BLN92),.WL(WL82));
sram_cell_6t_5 inst_cell_82_93 (.BL(BL93),.BLN(BLN93),.WL(WL82));
sram_cell_6t_5 inst_cell_82_94 (.BL(BL94),.BLN(BLN94),.WL(WL82));
sram_cell_6t_5 inst_cell_82_95 (.BL(BL95),.BLN(BLN95),.WL(WL82));
sram_cell_6t_5 inst_cell_82_96 (.BL(BL96),.BLN(BLN96),.WL(WL82));
sram_cell_6t_5 inst_cell_82_97 (.BL(BL97),.BLN(BLN97),.WL(WL82));
sram_cell_6t_5 inst_cell_82_98 (.BL(BL98),.BLN(BLN98),.WL(WL82));
sram_cell_6t_5 inst_cell_82_99 (.BL(BL99),.BLN(BLN99),.WL(WL82));
sram_cell_6t_5 inst_cell_82_100 (.BL(BL100),.BLN(BLN100),.WL(WL82));
sram_cell_6t_5 inst_cell_82_101 (.BL(BL101),.BLN(BLN101),.WL(WL82));
sram_cell_6t_5 inst_cell_82_102 (.BL(BL102),.BLN(BLN102),.WL(WL82));
sram_cell_6t_5 inst_cell_82_103 (.BL(BL103),.BLN(BLN103),.WL(WL82));
sram_cell_6t_5 inst_cell_82_104 (.BL(BL104),.BLN(BLN104),.WL(WL82));
sram_cell_6t_5 inst_cell_82_105 (.BL(BL105),.BLN(BLN105),.WL(WL82));
sram_cell_6t_5 inst_cell_82_106 (.BL(BL106),.BLN(BLN106),.WL(WL82));
sram_cell_6t_5 inst_cell_82_107 (.BL(BL107),.BLN(BLN107),.WL(WL82));
sram_cell_6t_5 inst_cell_82_108 (.BL(BL108),.BLN(BLN108),.WL(WL82));
sram_cell_6t_5 inst_cell_82_109 (.BL(BL109),.BLN(BLN109),.WL(WL82));
sram_cell_6t_5 inst_cell_82_110 (.BL(BL110),.BLN(BLN110),.WL(WL82));
sram_cell_6t_5 inst_cell_82_111 (.BL(BL111),.BLN(BLN111),.WL(WL82));
sram_cell_6t_5 inst_cell_82_112 (.BL(BL112),.BLN(BLN112),.WL(WL82));
sram_cell_6t_5 inst_cell_82_113 (.BL(BL113),.BLN(BLN113),.WL(WL82));
sram_cell_6t_5 inst_cell_82_114 (.BL(BL114),.BLN(BLN114),.WL(WL82));
sram_cell_6t_5 inst_cell_82_115 (.BL(BL115),.BLN(BLN115),.WL(WL82));
sram_cell_6t_5 inst_cell_82_116 (.BL(BL116),.BLN(BLN116),.WL(WL82));
sram_cell_6t_5 inst_cell_82_117 (.BL(BL117),.BLN(BLN117),.WL(WL82));
sram_cell_6t_5 inst_cell_82_118 (.BL(BL118),.BLN(BLN118),.WL(WL82));
sram_cell_6t_5 inst_cell_82_119 (.BL(BL119),.BLN(BLN119),.WL(WL82));
sram_cell_6t_5 inst_cell_82_120 (.BL(BL120),.BLN(BLN120),.WL(WL82));
sram_cell_6t_5 inst_cell_82_121 (.BL(BL121),.BLN(BLN121),.WL(WL82));
sram_cell_6t_5 inst_cell_82_122 (.BL(BL122),.BLN(BLN122),.WL(WL82));
sram_cell_6t_5 inst_cell_82_123 (.BL(BL123),.BLN(BLN123),.WL(WL82));
sram_cell_6t_5 inst_cell_82_124 (.BL(BL124),.BLN(BLN124),.WL(WL82));
sram_cell_6t_5 inst_cell_82_125 (.BL(BL125),.BLN(BLN125),.WL(WL82));
sram_cell_6t_5 inst_cell_82_126 (.BL(BL126),.BLN(BLN126),.WL(WL82));
sram_cell_6t_5 inst_cell_82_127 (.BL(BL127),.BLN(BLN127),.WL(WL82));
sram_cell_6t_5 inst_cell_83_0 (.BL(BL0),.BLN(BLN0),.WL(WL83));
sram_cell_6t_5 inst_cell_83_1 (.BL(BL1),.BLN(BLN1),.WL(WL83));
sram_cell_6t_5 inst_cell_83_2 (.BL(BL2),.BLN(BLN2),.WL(WL83));
sram_cell_6t_5 inst_cell_83_3 (.BL(BL3),.BLN(BLN3),.WL(WL83));
sram_cell_6t_5 inst_cell_83_4 (.BL(BL4),.BLN(BLN4),.WL(WL83));
sram_cell_6t_5 inst_cell_83_5 (.BL(BL5),.BLN(BLN5),.WL(WL83));
sram_cell_6t_5 inst_cell_83_6 (.BL(BL6),.BLN(BLN6),.WL(WL83));
sram_cell_6t_5 inst_cell_83_7 (.BL(BL7),.BLN(BLN7),.WL(WL83));
sram_cell_6t_5 inst_cell_83_8 (.BL(BL8),.BLN(BLN8),.WL(WL83));
sram_cell_6t_5 inst_cell_83_9 (.BL(BL9),.BLN(BLN9),.WL(WL83));
sram_cell_6t_5 inst_cell_83_10 (.BL(BL10),.BLN(BLN10),.WL(WL83));
sram_cell_6t_5 inst_cell_83_11 (.BL(BL11),.BLN(BLN11),.WL(WL83));
sram_cell_6t_5 inst_cell_83_12 (.BL(BL12),.BLN(BLN12),.WL(WL83));
sram_cell_6t_5 inst_cell_83_13 (.BL(BL13),.BLN(BLN13),.WL(WL83));
sram_cell_6t_5 inst_cell_83_14 (.BL(BL14),.BLN(BLN14),.WL(WL83));
sram_cell_6t_5 inst_cell_83_15 (.BL(BL15),.BLN(BLN15),.WL(WL83));
sram_cell_6t_5 inst_cell_83_16 (.BL(BL16),.BLN(BLN16),.WL(WL83));
sram_cell_6t_5 inst_cell_83_17 (.BL(BL17),.BLN(BLN17),.WL(WL83));
sram_cell_6t_5 inst_cell_83_18 (.BL(BL18),.BLN(BLN18),.WL(WL83));
sram_cell_6t_5 inst_cell_83_19 (.BL(BL19),.BLN(BLN19),.WL(WL83));
sram_cell_6t_5 inst_cell_83_20 (.BL(BL20),.BLN(BLN20),.WL(WL83));
sram_cell_6t_5 inst_cell_83_21 (.BL(BL21),.BLN(BLN21),.WL(WL83));
sram_cell_6t_5 inst_cell_83_22 (.BL(BL22),.BLN(BLN22),.WL(WL83));
sram_cell_6t_5 inst_cell_83_23 (.BL(BL23),.BLN(BLN23),.WL(WL83));
sram_cell_6t_5 inst_cell_83_24 (.BL(BL24),.BLN(BLN24),.WL(WL83));
sram_cell_6t_5 inst_cell_83_25 (.BL(BL25),.BLN(BLN25),.WL(WL83));
sram_cell_6t_5 inst_cell_83_26 (.BL(BL26),.BLN(BLN26),.WL(WL83));
sram_cell_6t_5 inst_cell_83_27 (.BL(BL27),.BLN(BLN27),.WL(WL83));
sram_cell_6t_5 inst_cell_83_28 (.BL(BL28),.BLN(BLN28),.WL(WL83));
sram_cell_6t_5 inst_cell_83_29 (.BL(BL29),.BLN(BLN29),.WL(WL83));
sram_cell_6t_5 inst_cell_83_30 (.BL(BL30),.BLN(BLN30),.WL(WL83));
sram_cell_6t_5 inst_cell_83_31 (.BL(BL31),.BLN(BLN31),.WL(WL83));
sram_cell_6t_5 inst_cell_83_32 (.BL(BL32),.BLN(BLN32),.WL(WL83));
sram_cell_6t_5 inst_cell_83_33 (.BL(BL33),.BLN(BLN33),.WL(WL83));
sram_cell_6t_5 inst_cell_83_34 (.BL(BL34),.BLN(BLN34),.WL(WL83));
sram_cell_6t_5 inst_cell_83_35 (.BL(BL35),.BLN(BLN35),.WL(WL83));
sram_cell_6t_5 inst_cell_83_36 (.BL(BL36),.BLN(BLN36),.WL(WL83));
sram_cell_6t_5 inst_cell_83_37 (.BL(BL37),.BLN(BLN37),.WL(WL83));
sram_cell_6t_5 inst_cell_83_38 (.BL(BL38),.BLN(BLN38),.WL(WL83));
sram_cell_6t_5 inst_cell_83_39 (.BL(BL39),.BLN(BLN39),.WL(WL83));
sram_cell_6t_5 inst_cell_83_40 (.BL(BL40),.BLN(BLN40),.WL(WL83));
sram_cell_6t_5 inst_cell_83_41 (.BL(BL41),.BLN(BLN41),.WL(WL83));
sram_cell_6t_5 inst_cell_83_42 (.BL(BL42),.BLN(BLN42),.WL(WL83));
sram_cell_6t_5 inst_cell_83_43 (.BL(BL43),.BLN(BLN43),.WL(WL83));
sram_cell_6t_5 inst_cell_83_44 (.BL(BL44),.BLN(BLN44),.WL(WL83));
sram_cell_6t_5 inst_cell_83_45 (.BL(BL45),.BLN(BLN45),.WL(WL83));
sram_cell_6t_5 inst_cell_83_46 (.BL(BL46),.BLN(BLN46),.WL(WL83));
sram_cell_6t_5 inst_cell_83_47 (.BL(BL47),.BLN(BLN47),.WL(WL83));
sram_cell_6t_5 inst_cell_83_48 (.BL(BL48),.BLN(BLN48),.WL(WL83));
sram_cell_6t_5 inst_cell_83_49 (.BL(BL49),.BLN(BLN49),.WL(WL83));
sram_cell_6t_5 inst_cell_83_50 (.BL(BL50),.BLN(BLN50),.WL(WL83));
sram_cell_6t_5 inst_cell_83_51 (.BL(BL51),.BLN(BLN51),.WL(WL83));
sram_cell_6t_5 inst_cell_83_52 (.BL(BL52),.BLN(BLN52),.WL(WL83));
sram_cell_6t_5 inst_cell_83_53 (.BL(BL53),.BLN(BLN53),.WL(WL83));
sram_cell_6t_5 inst_cell_83_54 (.BL(BL54),.BLN(BLN54),.WL(WL83));
sram_cell_6t_5 inst_cell_83_55 (.BL(BL55),.BLN(BLN55),.WL(WL83));
sram_cell_6t_5 inst_cell_83_56 (.BL(BL56),.BLN(BLN56),.WL(WL83));
sram_cell_6t_5 inst_cell_83_57 (.BL(BL57),.BLN(BLN57),.WL(WL83));
sram_cell_6t_5 inst_cell_83_58 (.BL(BL58),.BLN(BLN58),.WL(WL83));
sram_cell_6t_5 inst_cell_83_59 (.BL(BL59),.BLN(BLN59),.WL(WL83));
sram_cell_6t_5 inst_cell_83_60 (.BL(BL60),.BLN(BLN60),.WL(WL83));
sram_cell_6t_5 inst_cell_83_61 (.BL(BL61),.BLN(BLN61),.WL(WL83));
sram_cell_6t_5 inst_cell_83_62 (.BL(BL62),.BLN(BLN62),.WL(WL83));
sram_cell_6t_5 inst_cell_83_63 (.BL(BL63),.BLN(BLN63),.WL(WL83));
sram_cell_6t_5 inst_cell_83_64 (.BL(BL64),.BLN(BLN64),.WL(WL83));
sram_cell_6t_5 inst_cell_83_65 (.BL(BL65),.BLN(BLN65),.WL(WL83));
sram_cell_6t_5 inst_cell_83_66 (.BL(BL66),.BLN(BLN66),.WL(WL83));
sram_cell_6t_5 inst_cell_83_67 (.BL(BL67),.BLN(BLN67),.WL(WL83));
sram_cell_6t_5 inst_cell_83_68 (.BL(BL68),.BLN(BLN68),.WL(WL83));
sram_cell_6t_5 inst_cell_83_69 (.BL(BL69),.BLN(BLN69),.WL(WL83));
sram_cell_6t_5 inst_cell_83_70 (.BL(BL70),.BLN(BLN70),.WL(WL83));
sram_cell_6t_5 inst_cell_83_71 (.BL(BL71),.BLN(BLN71),.WL(WL83));
sram_cell_6t_5 inst_cell_83_72 (.BL(BL72),.BLN(BLN72),.WL(WL83));
sram_cell_6t_5 inst_cell_83_73 (.BL(BL73),.BLN(BLN73),.WL(WL83));
sram_cell_6t_5 inst_cell_83_74 (.BL(BL74),.BLN(BLN74),.WL(WL83));
sram_cell_6t_5 inst_cell_83_75 (.BL(BL75),.BLN(BLN75),.WL(WL83));
sram_cell_6t_5 inst_cell_83_76 (.BL(BL76),.BLN(BLN76),.WL(WL83));
sram_cell_6t_5 inst_cell_83_77 (.BL(BL77),.BLN(BLN77),.WL(WL83));
sram_cell_6t_5 inst_cell_83_78 (.BL(BL78),.BLN(BLN78),.WL(WL83));
sram_cell_6t_5 inst_cell_83_79 (.BL(BL79),.BLN(BLN79),.WL(WL83));
sram_cell_6t_5 inst_cell_83_80 (.BL(BL80),.BLN(BLN80),.WL(WL83));
sram_cell_6t_5 inst_cell_83_81 (.BL(BL81),.BLN(BLN81),.WL(WL83));
sram_cell_6t_5 inst_cell_83_82 (.BL(BL82),.BLN(BLN82),.WL(WL83));
sram_cell_6t_5 inst_cell_83_83 (.BL(BL83),.BLN(BLN83),.WL(WL83));
sram_cell_6t_5 inst_cell_83_84 (.BL(BL84),.BLN(BLN84),.WL(WL83));
sram_cell_6t_5 inst_cell_83_85 (.BL(BL85),.BLN(BLN85),.WL(WL83));
sram_cell_6t_5 inst_cell_83_86 (.BL(BL86),.BLN(BLN86),.WL(WL83));
sram_cell_6t_5 inst_cell_83_87 (.BL(BL87),.BLN(BLN87),.WL(WL83));
sram_cell_6t_5 inst_cell_83_88 (.BL(BL88),.BLN(BLN88),.WL(WL83));
sram_cell_6t_5 inst_cell_83_89 (.BL(BL89),.BLN(BLN89),.WL(WL83));
sram_cell_6t_5 inst_cell_83_90 (.BL(BL90),.BLN(BLN90),.WL(WL83));
sram_cell_6t_5 inst_cell_83_91 (.BL(BL91),.BLN(BLN91),.WL(WL83));
sram_cell_6t_5 inst_cell_83_92 (.BL(BL92),.BLN(BLN92),.WL(WL83));
sram_cell_6t_5 inst_cell_83_93 (.BL(BL93),.BLN(BLN93),.WL(WL83));
sram_cell_6t_5 inst_cell_83_94 (.BL(BL94),.BLN(BLN94),.WL(WL83));
sram_cell_6t_5 inst_cell_83_95 (.BL(BL95),.BLN(BLN95),.WL(WL83));
sram_cell_6t_5 inst_cell_83_96 (.BL(BL96),.BLN(BLN96),.WL(WL83));
sram_cell_6t_5 inst_cell_83_97 (.BL(BL97),.BLN(BLN97),.WL(WL83));
sram_cell_6t_5 inst_cell_83_98 (.BL(BL98),.BLN(BLN98),.WL(WL83));
sram_cell_6t_5 inst_cell_83_99 (.BL(BL99),.BLN(BLN99),.WL(WL83));
sram_cell_6t_5 inst_cell_83_100 (.BL(BL100),.BLN(BLN100),.WL(WL83));
sram_cell_6t_5 inst_cell_83_101 (.BL(BL101),.BLN(BLN101),.WL(WL83));
sram_cell_6t_5 inst_cell_83_102 (.BL(BL102),.BLN(BLN102),.WL(WL83));
sram_cell_6t_5 inst_cell_83_103 (.BL(BL103),.BLN(BLN103),.WL(WL83));
sram_cell_6t_5 inst_cell_83_104 (.BL(BL104),.BLN(BLN104),.WL(WL83));
sram_cell_6t_5 inst_cell_83_105 (.BL(BL105),.BLN(BLN105),.WL(WL83));
sram_cell_6t_5 inst_cell_83_106 (.BL(BL106),.BLN(BLN106),.WL(WL83));
sram_cell_6t_5 inst_cell_83_107 (.BL(BL107),.BLN(BLN107),.WL(WL83));
sram_cell_6t_5 inst_cell_83_108 (.BL(BL108),.BLN(BLN108),.WL(WL83));
sram_cell_6t_5 inst_cell_83_109 (.BL(BL109),.BLN(BLN109),.WL(WL83));
sram_cell_6t_5 inst_cell_83_110 (.BL(BL110),.BLN(BLN110),.WL(WL83));
sram_cell_6t_5 inst_cell_83_111 (.BL(BL111),.BLN(BLN111),.WL(WL83));
sram_cell_6t_5 inst_cell_83_112 (.BL(BL112),.BLN(BLN112),.WL(WL83));
sram_cell_6t_5 inst_cell_83_113 (.BL(BL113),.BLN(BLN113),.WL(WL83));
sram_cell_6t_5 inst_cell_83_114 (.BL(BL114),.BLN(BLN114),.WL(WL83));
sram_cell_6t_5 inst_cell_83_115 (.BL(BL115),.BLN(BLN115),.WL(WL83));
sram_cell_6t_5 inst_cell_83_116 (.BL(BL116),.BLN(BLN116),.WL(WL83));
sram_cell_6t_5 inst_cell_83_117 (.BL(BL117),.BLN(BLN117),.WL(WL83));
sram_cell_6t_5 inst_cell_83_118 (.BL(BL118),.BLN(BLN118),.WL(WL83));
sram_cell_6t_5 inst_cell_83_119 (.BL(BL119),.BLN(BLN119),.WL(WL83));
sram_cell_6t_5 inst_cell_83_120 (.BL(BL120),.BLN(BLN120),.WL(WL83));
sram_cell_6t_5 inst_cell_83_121 (.BL(BL121),.BLN(BLN121),.WL(WL83));
sram_cell_6t_5 inst_cell_83_122 (.BL(BL122),.BLN(BLN122),.WL(WL83));
sram_cell_6t_5 inst_cell_83_123 (.BL(BL123),.BLN(BLN123),.WL(WL83));
sram_cell_6t_5 inst_cell_83_124 (.BL(BL124),.BLN(BLN124),.WL(WL83));
sram_cell_6t_5 inst_cell_83_125 (.BL(BL125),.BLN(BLN125),.WL(WL83));
sram_cell_6t_5 inst_cell_83_126 (.BL(BL126),.BLN(BLN126),.WL(WL83));
sram_cell_6t_5 inst_cell_83_127 (.BL(BL127),.BLN(BLN127),.WL(WL83));
sram_cell_6t_5 inst_cell_84_0 (.BL(BL0),.BLN(BLN0),.WL(WL84));
sram_cell_6t_5 inst_cell_84_1 (.BL(BL1),.BLN(BLN1),.WL(WL84));
sram_cell_6t_5 inst_cell_84_2 (.BL(BL2),.BLN(BLN2),.WL(WL84));
sram_cell_6t_5 inst_cell_84_3 (.BL(BL3),.BLN(BLN3),.WL(WL84));
sram_cell_6t_5 inst_cell_84_4 (.BL(BL4),.BLN(BLN4),.WL(WL84));
sram_cell_6t_5 inst_cell_84_5 (.BL(BL5),.BLN(BLN5),.WL(WL84));
sram_cell_6t_5 inst_cell_84_6 (.BL(BL6),.BLN(BLN6),.WL(WL84));
sram_cell_6t_5 inst_cell_84_7 (.BL(BL7),.BLN(BLN7),.WL(WL84));
sram_cell_6t_5 inst_cell_84_8 (.BL(BL8),.BLN(BLN8),.WL(WL84));
sram_cell_6t_5 inst_cell_84_9 (.BL(BL9),.BLN(BLN9),.WL(WL84));
sram_cell_6t_5 inst_cell_84_10 (.BL(BL10),.BLN(BLN10),.WL(WL84));
sram_cell_6t_5 inst_cell_84_11 (.BL(BL11),.BLN(BLN11),.WL(WL84));
sram_cell_6t_5 inst_cell_84_12 (.BL(BL12),.BLN(BLN12),.WL(WL84));
sram_cell_6t_5 inst_cell_84_13 (.BL(BL13),.BLN(BLN13),.WL(WL84));
sram_cell_6t_5 inst_cell_84_14 (.BL(BL14),.BLN(BLN14),.WL(WL84));
sram_cell_6t_5 inst_cell_84_15 (.BL(BL15),.BLN(BLN15),.WL(WL84));
sram_cell_6t_5 inst_cell_84_16 (.BL(BL16),.BLN(BLN16),.WL(WL84));
sram_cell_6t_5 inst_cell_84_17 (.BL(BL17),.BLN(BLN17),.WL(WL84));
sram_cell_6t_5 inst_cell_84_18 (.BL(BL18),.BLN(BLN18),.WL(WL84));
sram_cell_6t_5 inst_cell_84_19 (.BL(BL19),.BLN(BLN19),.WL(WL84));
sram_cell_6t_5 inst_cell_84_20 (.BL(BL20),.BLN(BLN20),.WL(WL84));
sram_cell_6t_5 inst_cell_84_21 (.BL(BL21),.BLN(BLN21),.WL(WL84));
sram_cell_6t_5 inst_cell_84_22 (.BL(BL22),.BLN(BLN22),.WL(WL84));
sram_cell_6t_5 inst_cell_84_23 (.BL(BL23),.BLN(BLN23),.WL(WL84));
sram_cell_6t_5 inst_cell_84_24 (.BL(BL24),.BLN(BLN24),.WL(WL84));
sram_cell_6t_5 inst_cell_84_25 (.BL(BL25),.BLN(BLN25),.WL(WL84));
sram_cell_6t_5 inst_cell_84_26 (.BL(BL26),.BLN(BLN26),.WL(WL84));
sram_cell_6t_5 inst_cell_84_27 (.BL(BL27),.BLN(BLN27),.WL(WL84));
sram_cell_6t_5 inst_cell_84_28 (.BL(BL28),.BLN(BLN28),.WL(WL84));
sram_cell_6t_5 inst_cell_84_29 (.BL(BL29),.BLN(BLN29),.WL(WL84));
sram_cell_6t_5 inst_cell_84_30 (.BL(BL30),.BLN(BLN30),.WL(WL84));
sram_cell_6t_5 inst_cell_84_31 (.BL(BL31),.BLN(BLN31),.WL(WL84));
sram_cell_6t_5 inst_cell_84_32 (.BL(BL32),.BLN(BLN32),.WL(WL84));
sram_cell_6t_5 inst_cell_84_33 (.BL(BL33),.BLN(BLN33),.WL(WL84));
sram_cell_6t_5 inst_cell_84_34 (.BL(BL34),.BLN(BLN34),.WL(WL84));
sram_cell_6t_5 inst_cell_84_35 (.BL(BL35),.BLN(BLN35),.WL(WL84));
sram_cell_6t_5 inst_cell_84_36 (.BL(BL36),.BLN(BLN36),.WL(WL84));
sram_cell_6t_5 inst_cell_84_37 (.BL(BL37),.BLN(BLN37),.WL(WL84));
sram_cell_6t_5 inst_cell_84_38 (.BL(BL38),.BLN(BLN38),.WL(WL84));
sram_cell_6t_5 inst_cell_84_39 (.BL(BL39),.BLN(BLN39),.WL(WL84));
sram_cell_6t_5 inst_cell_84_40 (.BL(BL40),.BLN(BLN40),.WL(WL84));
sram_cell_6t_5 inst_cell_84_41 (.BL(BL41),.BLN(BLN41),.WL(WL84));
sram_cell_6t_5 inst_cell_84_42 (.BL(BL42),.BLN(BLN42),.WL(WL84));
sram_cell_6t_5 inst_cell_84_43 (.BL(BL43),.BLN(BLN43),.WL(WL84));
sram_cell_6t_5 inst_cell_84_44 (.BL(BL44),.BLN(BLN44),.WL(WL84));
sram_cell_6t_5 inst_cell_84_45 (.BL(BL45),.BLN(BLN45),.WL(WL84));
sram_cell_6t_5 inst_cell_84_46 (.BL(BL46),.BLN(BLN46),.WL(WL84));
sram_cell_6t_5 inst_cell_84_47 (.BL(BL47),.BLN(BLN47),.WL(WL84));
sram_cell_6t_5 inst_cell_84_48 (.BL(BL48),.BLN(BLN48),.WL(WL84));
sram_cell_6t_5 inst_cell_84_49 (.BL(BL49),.BLN(BLN49),.WL(WL84));
sram_cell_6t_5 inst_cell_84_50 (.BL(BL50),.BLN(BLN50),.WL(WL84));
sram_cell_6t_5 inst_cell_84_51 (.BL(BL51),.BLN(BLN51),.WL(WL84));
sram_cell_6t_5 inst_cell_84_52 (.BL(BL52),.BLN(BLN52),.WL(WL84));
sram_cell_6t_5 inst_cell_84_53 (.BL(BL53),.BLN(BLN53),.WL(WL84));
sram_cell_6t_5 inst_cell_84_54 (.BL(BL54),.BLN(BLN54),.WL(WL84));
sram_cell_6t_5 inst_cell_84_55 (.BL(BL55),.BLN(BLN55),.WL(WL84));
sram_cell_6t_5 inst_cell_84_56 (.BL(BL56),.BLN(BLN56),.WL(WL84));
sram_cell_6t_5 inst_cell_84_57 (.BL(BL57),.BLN(BLN57),.WL(WL84));
sram_cell_6t_5 inst_cell_84_58 (.BL(BL58),.BLN(BLN58),.WL(WL84));
sram_cell_6t_5 inst_cell_84_59 (.BL(BL59),.BLN(BLN59),.WL(WL84));
sram_cell_6t_5 inst_cell_84_60 (.BL(BL60),.BLN(BLN60),.WL(WL84));
sram_cell_6t_5 inst_cell_84_61 (.BL(BL61),.BLN(BLN61),.WL(WL84));
sram_cell_6t_5 inst_cell_84_62 (.BL(BL62),.BLN(BLN62),.WL(WL84));
sram_cell_6t_5 inst_cell_84_63 (.BL(BL63),.BLN(BLN63),.WL(WL84));
sram_cell_6t_5 inst_cell_84_64 (.BL(BL64),.BLN(BLN64),.WL(WL84));
sram_cell_6t_5 inst_cell_84_65 (.BL(BL65),.BLN(BLN65),.WL(WL84));
sram_cell_6t_5 inst_cell_84_66 (.BL(BL66),.BLN(BLN66),.WL(WL84));
sram_cell_6t_5 inst_cell_84_67 (.BL(BL67),.BLN(BLN67),.WL(WL84));
sram_cell_6t_5 inst_cell_84_68 (.BL(BL68),.BLN(BLN68),.WL(WL84));
sram_cell_6t_5 inst_cell_84_69 (.BL(BL69),.BLN(BLN69),.WL(WL84));
sram_cell_6t_5 inst_cell_84_70 (.BL(BL70),.BLN(BLN70),.WL(WL84));
sram_cell_6t_5 inst_cell_84_71 (.BL(BL71),.BLN(BLN71),.WL(WL84));
sram_cell_6t_5 inst_cell_84_72 (.BL(BL72),.BLN(BLN72),.WL(WL84));
sram_cell_6t_5 inst_cell_84_73 (.BL(BL73),.BLN(BLN73),.WL(WL84));
sram_cell_6t_5 inst_cell_84_74 (.BL(BL74),.BLN(BLN74),.WL(WL84));
sram_cell_6t_5 inst_cell_84_75 (.BL(BL75),.BLN(BLN75),.WL(WL84));
sram_cell_6t_5 inst_cell_84_76 (.BL(BL76),.BLN(BLN76),.WL(WL84));
sram_cell_6t_5 inst_cell_84_77 (.BL(BL77),.BLN(BLN77),.WL(WL84));
sram_cell_6t_5 inst_cell_84_78 (.BL(BL78),.BLN(BLN78),.WL(WL84));
sram_cell_6t_5 inst_cell_84_79 (.BL(BL79),.BLN(BLN79),.WL(WL84));
sram_cell_6t_5 inst_cell_84_80 (.BL(BL80),.BLN(BLN80),.WL(WL84));
sram_cell_6t_5 inst_cell_84_81 (.BL(BL81),.BLN(BLN81),.WL(WL84));
sram_cell_6t_5 inst_cell_84_82 (.BL(BL82),.BLN(BLN82),.WL(WL84));
sram_cell_6t_5 inst_cell_84_83 (.BL(BL83),.BLN(BLN83),.WL(WL84));
sram_cell_6t_5 inst_cell_84_84 (.BL(BL84),.BLN(BLN84),.WL(WL84));
sram_cell_6t_5 inst_cell_84_85 (.BL(BL85),.BLN(BLN85),.WL(WL84));
sram_cell_6t_5 inst_cell_84_86 (.BL(BL86),.BLN(BLN86),.WL(WL84));
sram_cell_6t_5 inst_cell_84_87 (.BL(BL87),.BLN(BLN87),.WL(WL84));
sram_cell_6t_5 inst_cell_84_88 (.BL(BL88),.BLN(BLN88),.WL(WL84));
sram_cell_6t_5 inst_cell_84_89 (.BL(BL89),.BLN(BLN89),.WL(WL84));
sram_cell_6t_5 inst_cell_84_90 (.BL(BL90),.BLN(BLN90),.WL(WL84));
sram_cell_6t_5 inst_cell_84_91 (.BL(BL91),.BLN(BLN91),.WL(WL84));
sram_cell_6t_5 inst_cell_84_92 (.BL(BL92),.BLN(BLN92),.WL(WL84));
sram_cell_6t_5 inst_cell_84_93 (.BL(BL93),.BLN(BLN93),.WL(WL84));
sram_cell_6t_5 inst_cell_84_94 (.BL(BL94),.BLN(BLN94),.WL(WL84));
sram_cell_6t_5 inst_cell_84_95 (.BL(BL95),.BLN(BLN95),.WL(WL84));
sram_cell_6t_5 inst_cell_84_96 (.BL(BL96),.BLN(BLN96),.WL(WL84));
sram_cell_6t_5 inst_cell_84_97 (.BL(BL97),.BLN(BLN97),.WL(WL84));
sram_cell_6t_5 inst_cell_84_98 (.BL(BL98),.BLN(BLN98),.WL(WL84));
sram_cell_6t_5 inst_cell_84_99 (.BL(BL99),.BLN(BLN99),.WL(WL84));
sram_cell_6t_5 inst_cell_84_100 (.BL(BL100),.BLN(BLN100),.WL(WL84));
sram_cell_6t_5 inst_cell_84_101 (.BL(BL101),.BLN(BLN101),.WL(WL84));
sram_cell_6t_5 inst_cell_84_102 (.BL(BL102),.BLN(BLN102),.WL(WL84));
sram_cell_6t_5 inst_cell_84_103 (.BL(BL103),.BLN(BLN103),.WL(WL84));
sram_cell_6t_5 inst_cell_84_104 (.BL(BL104),.BLN(BLN104),.WL(WL84));
sram_cell_6t_5 inst_cell_84_105 (.BL(BL105),.BLN(BLN105),.WL(WL84));
sram_cell_6t_5 inst_cell_84_106 (.BL(BL106),.BLN(BLN106),.WL(WL84));
sram_cell_6t_5 inst_cell_84_107 (.BL(BL107),.BLN(BLN107),.WL(WL84));
sram_cell_6t_5 inst_cell_84_108 (.BL(BL108),.BLN(BLN108),.WL(WL84));
sram_cell_6t_5 inst_cell_84_109 (.BL(BL109),.BLN(BLN109),.WL(WL84));
sram_cell_6t_5 inst_cell_84_110 (.BL(BL110),.BLN(BLN110),.WL(WL84));
sram_cell_6t_5 inst_cell_84_111 (.BL(BL111),.BLN(BLN111),.WL(WL84));
sram_cell_6t_5 inst_cell_84_112 (.BL(BL112),.BLN(BLN112),.WL(WL84));
sram_cell_6t_5 inst_cell_84_113 (.BL(BL113),.BLN(BLN113),.WL(WL84));
sram_cell_6t_5 inst_cell_84_114 (.BL(BL114),.BLN(BLN114),.WL(WL84));
sram_cell_6t_5 inst_cell_84_115 (.BL(BL115),.BLN(BLN115),.WL(WL84));
sram_cell_6t_5 inst_cell_84_116 (.BL(BL116),.BLN(BLN116),.WL(WL84));
sram_cell_6t_5 inst_cell_84_117 (.BL(BL117),.BLN(BLN117),.WL(WL84));
sram_cell_6t_5 inst_cell_84_118 (.BL(BL118),.BLN(BLN118),.WL(WL84));
sram_cell_6t_5 inst_cell_84_119 (.BL(BL119),.BLN(BLN119),.WL(WL84));
sram_cell_6t_5 inst_cell_84_120 (.BL(BL120),.BLN(BLN120),.WL(WL84));
sram_cell_6t_5 inst_cell_84_121 (.BL(BL121),.BLN(BLN121),.WL(WL84));
sram_cell_6t_5 inst_cell_84_122 (.BL(BL122),.BLN(BLN122),.WL(WL84));
sram_cell_6t_5 inst_cell_84_123 (.BL(BL123),.BLN(BLN123),.WL(WL84));
sram_cell_6t_5 inst_cell_84_124 (.BL(BL124),.BLN(BLN124),.WL(WL84));
sram_cell_6t_5 inst_cell_84_125 (.BL(BL125),.BLN(BLN125),.WL(WL84));
sram_cell_6t_5 inst_cell_84_126 (.BL(BL126),.BLN(BLN126),.WL(WL84));
sram_cell_6t_5 inst_cell_84_127 (.BL(BL127),.BLN(BLN127),.WL(WL84));
sram_cell_6t_5 inst_cell_85_0 (.BL(BL0),.BLN(BLN0),.WL(WL85));
sram_cell_6t_5 inst_cell_85_1 (.BL(BL1),.BLN(BLN1),.WL(WL85));
sram_cell_6t_5 inst_cell_85_2 (.BL(BL2),.BLN(BLN2),.WL(WL85));
sram_cell_6t_5 inst_cell_85_3 (.BL(BL3),.BLN(BLN3),.WL(WL85));
sram_cell_6t_5 inst_cell_85_4 (.BL(BL4),.BLN(BLN4),.WL(WL85));
sram_cell_6t_5 inst_cell_85_5 (.BL(BL5),.BLN(BLN5),.WL(WL85));
sram_cell_6t_5 inst_cell_85_6 (.BL(BL6),.BLN(BLN6),.WL(WL85));
sram_cell_6t_5 inst_cell_85_7 (.BL(BL7),.BLN(BLN7),.WL(WL85));
sram_cell_6t_5 inst_cell_85_8 (.BL(BL8),.BLN(BLN8),.WL(WL85));
sram_cell_6t_5 inst_cell_85_9 (.BL(BL9),.BLN(BLN9),.WL(WL85));
sram_cell_6t_5 inst_cell_85_10 (.BL(BL10),.BLN(BLN10),.WL(WL85));
sram_cell_6t_5 inst_cell_85_11 (.BL(BL11),.BLN(BLN11),.WL(WL85));
sram_cell_6t_5 inst_cell_85_12 (.BL(BL12),.BLN(BLN12),.WL(WL85));
sram_cell_6t_5 inst_cell_85_13 (.BL(BL13),.BLN(BLN13),.WL(WL85));
sram_cell_6t_5 inst_cell_85_14 (.BL(BL14),.BLN(BLN14),.WL(WL85));
sram_cell_6t_5 inst_cell_85_15 (.BL(BL15),.BLN(BLN15),.WL(WL85));
sram_cell_6t_5 inst_cell_85_16 (.BL(BL16),.BLN(BLN16),.WL(WL85));
sram_cell_6t_5 inst_cell_85_17 (.BL(BL17),.BLN(BLN17),.WL(WL85));
sram_cell_6t_5 inst_cell_85_18 (.BL(BL18),.BLN(BLN18),.WL(WL85));
sram_cell_6t_5 inst_cell_85_19 (.BL(BL19),.BLN(BLN19),.WL(WL85));
sram_cell_6t_5 inst_cell_85_20 (.BL(BL20),.BLN(BLN20),.WL(WL85));
sram_cell_6t_5 inst_cell_85_21 (.BL(BL21),.BLN(BLN21),.WL(WL85));
sram_cell_6t_5 inst_cell_85_22 (.BL(BL22),.BLN(BLN22),.WL(WL85));
sram_cell_6t_5 inst_cell_85_23 (.BL(BL23),.BLN(BLN23),.WL(WL85));
sram_cell_6t_5 inst_cell_85_24 (.BL(BL24),.BLN(BLN24),.WL(WL85));
sram_cell_6t_5 inst_cell_85_25 (.BL(BL25),.BLN(BLN25),.WL(WL85));
sram_cell_6t_5 inst_cell_85_26 (.BL(BL26),.BLN(BLN26),.WL(WL85));
sram_cell_6t_5 inst_cell_85_27 (.BL(BL27),.BLN(BLN27),.WL(WL85));
sram_cell_6t_5 inst_cell_85_28 (.BL(BL28),.BLN(BLN28),.WL(WL85));
sram_cell_6t_5 inst_cell_85_29 (.BL(BL29),.BLN(BLN29),.WL(WL85));
sram_cell_6t_5 inst_cell_85_30 (.BL(BL30),.BLN(BLN30),.WL(WL85));
sram_cell_6t_5 inst_cell_85_31 (.BL(BL31),.BLN(BLN31),.WL(WL85));
sram_cell_6t_5 inst_cell_85_32 (.BL(BL32),.BLN(BLN32),.WL(WL85));
sram_cell_6t_5 inst_cell_85_33 (.BL(BL33),.BLN(BLN33),.WL(WL85));
sram_cell_6t_5 inst_cell_85_34 (.BL(BL34),.BLN(BLN34),.WL(WL85));
sram_cell_6t_5 inst_cell_85_35 (.BL(BL35),.BLN(BLN35),.WL(WL85));
sram_cell_6t_5 inst_cell_85_36 (.BL(BL36),.BLN(BLN36),.WL(WL85));
sram_cell_6t_5 inst_cell_85_37 (.BL(BL37),.BLN(BLN37),.WL(WL85));
sram_cell_6t_5 inst_cell_85_38 (.BL(BL38),.BLN(BLN38),.WL(WL85));
sram_cell_6t_5 inst_cell_85_39 (.BL(BL39),.BLN(BLN39),.WL(WL85));
sram_cell_6t_5 inst_cell_85_40 (.BL(BL40),.BLN(BLN40),.WL(WL85));
sram_cell_6t_5 inst_cell_85_41 (.BL(BL41),.BLN(BLN41),.WL(WL85));
sram_cell_6t_5 inst_cell_85_42 (.BL(BL42),.BLN(BLN42),.WL(WL85));
sram_cell_6t_5 inst_cell_85_43 (.BL(BL43),.BLN(BLN43),.WL(WL85));
sram_cell_6t_5 inst_cell_85_44 (.BL(BL44),.BLN(BLN44),.WL(WL85));
sram_cell_6t_5 inst_cell_85_45 (.BL(BL45),.BLN(BLN45),.WL(WL85));
sram_cell_6t_5 inst_cell_85_46 (.BL(BL46),.BLN(BLN46),.WL(WL85));
sram_cell_6t_5 inst_cell_85_47 (.BL(BL47),.BLN(BLN47),.WL(WL85));
sram_cell_6t_5 inst_cell_85_48 (.BL(BL48),.BLN(BLN48),.WL(WL85));
sram_cell_6t_5 inst_cell_85_49 (.BL(BL49),.BLN(BLN49),.WL(WL85));
sram_cell_6t_5 inst_cell_85_50 (.BL(BL50),.BLN(BLN50),.WL(WL85));
sram_cell_6t_5 inst_cell_85_51 (.BL(BL51),.BLN(BLN51),.WL(WL85));
sram_cell_6t_5 inst_cell_85_52 (.BL(BL52),.BLN(BLN52),.WL(WL85));
sram_cell_6t_5 inst_cell_85_53 (.BL(BL53),.BLN(BLN53),.WL(WL85));
sram_cell_6t_5 inst_cell_85_54 (.BL(BL54),.BLN(BLN54),.WL(WL85));
sram_cell_6t_5 inst_cell_85_55 (.BL(BL55),.BLN(BLN55),.WL(WL85));
sram_cell_6t_5 inst_cell_85_56 (.BL(BL56),.BLN(BLN56),.WL(WL85));
sram_cell_6t_5 inst_cell_85_57 (.BL(BL57),.BLN(BLN57),.WL(WL85));
sram_cell_6t_5 inst_cell_85_58 (.BL(BL58),.BLN(BLN58),.WL(WL85));
sram_cell_6t_5 inst_cell_85_59 (.BL(BL59),.BLN(BLN59),.WL(WL85));
sram_cell_6t_5 inst_cell_85_60 (.BL(BL60),.BLN(BLN60),.WL(WL85));
sram_cell_6t_5 inst_cell_85_61 (.BL(BL61),.BLN(BLN61),.WL(WL85));
sram_cell_6t_5 inst_cell_85_62 (.BL(BL62),.BLN(BLN62),.WL(WL85));
sram_cell_6t_5 inst_cell_85_63 (.BL(BL63),.BLN(BLN63),.WL(WL85));
sram_cell_6t_5 inst_cell_85_64 (.BL(BL64),.BLN(BLN64),.WL(WL85));
sram_cell_6t_5 inst_cell_85_65 (.BL(BL65),.BLN(BLN65),.WL(WL85));
sram_cell_6t_5 inst_cell_85_66 (.BL(BL66),.BLN(BLN66),.WL(WL85));
sram_cell_6t_5 inst_cell_85_67 (.BL(BL67),.BLN(BLN67),.WL(WL85));
sram_cell_6t_5 inst_cell_85_68 (.BL(BL68),.BLN(BLN68),.WL(WL85));
sram_cell_6t_5 inst_cell_85_69 (.BL(BL69),.BLN(BLN69),.WL(WL85));
sram_cell_6t_5 inst_cell_85_70 (.BL(BL70),.BLN(BLN70),.WL(WL85));
sram_cell_6t_5 inst_cell_85_71 (.BL(BL71),.BLN(BLN71),.WL(WL85));
sram_cell_6t_5 inst_cell_85_72 (.BL(BL72),.BLN(BLN72),.WL(WL85));
sram_cell_6t_5 inst_cell_85_73 (.BL(BL73),.BLN(BLN73),.WL(WL85));
sram_cell_6t_5 inst_cell_85_74 (.BL(BL74),.BLN(BLN74),.WL(WL85));
sram_cell_6t_5 inst_cell_85_75 (.BL(BL75),.BLN(BLN75),.WL(WL85));
sram_cell_6t_5 inst_cell_85_76 (.BL(BL76),.BLN(BLN76),.WL(WL85));
sram_cell_6t_5 inst_cell_85_77 (.BL(BL77),.BLN(BLN77),.WL(WL85));
sram_cell_6t_5 inst_cell_85_78 (.BL(BL78),.BLN(BLN78),.WL(WL85));
sram_cell_6t_5 inst_cell_85_79 (.BL(BL79),.BLN(BLN79),.WL(WL85));
sram_cell_6t_5 inst_cell_85_80 (.BL(BL80),.BLN(BLN80),.WL(WL85));
sram_cell_6t_5 inst_cell_85_81 (.BL(BL81),.BLN(BLN81),.WL(WL85));
sram_cell_6t_5 inst_cell_85_82 (.BL(BL82),.BLN(BLN82),.WL(WL85));
sram_cell_6t_5 inst_cell_85_83 (.BL(BL83),.BLN(BLN83),.WL(WL85));
sram_cell_6t_5 inst_cell_85_84 (.BL(BL84),.BLN(BLN84),.WL(WL85));
sram_cell_6t_5 inst_cell_85_85 (.BL(BL85),.BLN(BLN85),.WL(WL85));
sram_cell_6t_5 inst_cell_85_86 (.BL(BL86),.BLN(BLN86),.WL(WL85));
sram_cell_6t_5 inst_cell_85_87 (.BL(BL87),.BLN(BLN87),.WL(WL85));
sram_cell_6t_5 inst_cell_85_88 (.BL(BL88),.BLN(BLN88),.WL(WL85));
sram_cell_6t_5 inst_cell_85_89 (.BL(BL89),.BLN(BLN89),.WL(WL85));
sram_cell_6t_5 inst_cell_85_90 (.BL(BL90),.BLN(BLN90),.WL(WL85));
sram_cell_6t_5 inst_cell_85_91 (.BL(BL91),.BLN(BLN91),.WL(WL85));
sram_cell_6t_5 inst_cell_85_92 (.BL(BL92),.BLN(BLN92),.WL(WL85));
sram_cell_6t_5 inst_cell_85_93 (.BL(BL93),.BLN(BLN93),.WL(WL85));
sram_cell_6t_5 inst_cell_85_94 (.BL(BL94),.BLN(BLN94),.WL(WL85));
sram_cell_6t_5 inst_cell_85_95 (.BL(BL95),.BLN(BLN95),.WL(WL85));
sram_cell_6t_5 inst_cell_85_96 (.BL(BL96),.BLN(BLN96),.WL(WL85));
sram_cell_6t_5 inst_cell_85_97 (.BL(BL97),.BLN(BLN97),.WL(WL85));
sram_cell_6t_5 inst_cell_85_98 (.BL(BL98),.BLN(BLN98),.WL(WL85));
sram_cell_6t_5 inst_cell_85_99 (.BL(BL99),.BLN(BLN99),.WL(WL85));
sram_cell_6t_5 inst_cell_85_100 (.BL(BL100),.BLN(BLN100),.WL(WL85));
sram_cell_6t_5 inst_cell_85_101 (.BL(BL101),.BLN(BLN101),.WL(WL85));
sram_cell_6t_5 inst_cell_85_102 (.BL(BL102),.BLN(BLN102),.WL(WL85));
sram_cell_6t_5 inst_cell_85_103 (.BL(BL103),.BLN(BLN103),.WL(WL85));
sram_cell_6t_5 inst_cell_85_104 (.BL(BL104),.BLN(BLN104),.WL(WL85));
sram_cell_6t_5 inst_cell_85_105 (.BL(BL105),.BLN(BLN105),.WL(WL85));
sram_cell_6t_5 inst_cell_85_106 (.BL(BL106),.BLN(BLN106),.WL(WL85));
sram_cell_6t_5 inst_cell_85_107 (.BL(BL107),.BLN(BLN107),.WL(WL85));
sram_cell_6t_5 inst_cell_85_108 (.BL(BL108),.BLN(BLN108),.WL(WL85));
sram_cell_6t_5 inst_cell_85_109 (.BL(BL109),.BLN(BLN109),.WL(WL85));
sram_cell_6t_5 inst_cell_85_110 (.BL(BL110),.BLN(BLN110),.WL(WL85));
sram_cell_6t_5 inst_cell_85_111 (.BL(BL111),.BLN(BLN111),.WL(WL85));
sram_cell_6t_5 inst_cell_85_112 (.BL(BL112),.BLN(BLN112),.WL(WL85));
sram_cell_6t_5 inst_cell_85_113 (.BL(BL113),.BLN(BLN113),.WL(WL85));
sram_cell_6t_5 inst_cell_85_114 (.BL(BL114),.BLN(BLN114),.WL(WL85));
sram_cell_6t_5 inst_cell_85_115 (.BL(BL115),.BLN(BLN115),.WL(WL85));
sram_cell_6t_5 inst_cell_85_116 (.BL(BL116),.BLN(BLN116),.WL(WL85));
sram_cell_6t_5 inst_cell_85_117 (.BL(BL117),.BLN(BLN117),.WL(WL85));
sram_cell_6t_5 inst_cell_85_118 (.BL(BL118),.BLN(BLN118),.WL(WL85));
sram_cell_6t_5 inst_cell_85_119 (.BL(BL119),.BLN(BLN119),.WL(WL85));
sram_cell_6t_5 inst_cell_85_120 (.BL(BL120),.BLN(BLN120),.WL(WL85));
sram_cell_6t_5 inst_cell_85_121 (.BL(BL121),.BLN(BLN121),.WL(WL85));
sram_cell_6t_5 inst_cell_85_122 (.BL(BL122),.BLN(BLN122),.WL(WL85));
sram_cell_6t_5 inst_cell_85_123 (.BL(BL123),.BLN(BLN123),.WL(WL85));
sram_cell_6t_5 inst_cell_85_124 (.BL(BL124),.BLN(BLN124),.WL(WL85));
sram_cell_6t_5 inst_cell_85_125 (.BL(BL125),.BLN(BLN125),.WL(WL85));
sram_cell_6t_5 inst_cell_85_126 (.BL(BL126),.BLN(BLN126),.WL(WL85));
sram_cell_6t_5 inst_cell_85_127 (.BL(BL127),.BLN(BLN127),.WL(WL85));
sram_cell_6t_5 inst_cell_86_0 (.BL(BL0),.BLN(BLN0),.WL(WL86));
sram_cell_6t_5 inst_cell_86_1 (.BL(BL1),.BLN(BLN1),.WL(WL86));
sram_cell_6t_5 inst_cell_86_2 (.BL(BL2),.BLN(BLN2),.WL(WL86));
sram_cell_6t_5 inst_cell_86_3 (.BL(BL3),.BLN(BLN3),.WL(WL86));
sram_cell_6t_5 inst_cell_86_4 (.BL(BL4),.BLN(BLN4),.WL(WL86));
sram_cell_6t_5 inst_cell_86_5 (.BL(BL5),.BLN(BLN5),.WL(WL86));
sram_cell_6t_5 inst_cell_86_6 (.BL(BL6),.BLN(BLN6),.WL(WL86));
sram_cell_6t_5 inst_cell_86_7 (.BL(BL7),.BLN(BLN7),.WL(WL86));
sram_cell_6t_5 inst_cell_86_8 (.BL(BL8),.BLN(BLN8),.WL(WL86));
sram_cell_6t_5 inst_cell_86_9 (.BL(BL9),.BLN(BLN9),.WL(WL86));
sram_cell_6t_5 inst_cell_86_10 (.BL(BL10),.BLN(BLN10),.WL(WL86));
sram_cell_6t_5 inst_cell_86_11 (.BL(BL11),.BLN(BLN11),.WL(WL86));
sram_cell_6t_5 inst_cell_86_12 (.BL(BL12),.BLN(BLN12),.WL(WL86));
sram_cell_6t_5 inst_cell_86_13 (.BL(BL13),.BLN(BLN13),.WL(WL86));
sram_cell_6t_5 inst_cell_86_14 (.BL(BL14),.BLN(BLN14),.WL(WL86));
sram_cell_6t_5 inst_cell_86_15 (.BL(BL15),.BLN(BLN15),.WL(WL86));
sram_cell_6t_5 inst_cell_86_16 (.BL(BL16),.BLN(BLN16),.WL(WL86));
sram_cell_6t_5 inst_cell_86_17 (.BL(BL17),.BLN(BLN17),.WL(WL86));
sram_cell_6t_5 inst_cell_86_18 (.BL(BL18),.BLN(BLN18),.WL(WL86));
sram_cell_6t_5 inst_cell_86_19 (.BL(BL19),.BLN(BLN19),.WL(WL86));
sram_cell_6t_5 inst_cell_86_20 (.BL(BL20),.BLN(BLN20),.WL(WL86));
sram_cell_6t_5 inst_cell_86_21 (.BL(BL21),.BLN(BLN21),.WL(WL86));
sram_cell_6t_5 inst_cell_86_22 (.BL(BL22),.BLN(BLN22),.WL(WL86));
sram_cell_6t_5 inst_cell_86_23 (.BL(BL23),.BLN(BLN23),.WL(WL86));
sram_cell_6t_5 inst_cell_86_24 (.BL(BL24),.BLN(BLN24),.WL(WL86));
sram_cell_6t_5 inst_cell_86_25 (.BL(BL25),.BLN(BLN25),.WL(WL86));
sram_cell_6t_5 inst_cell_86_26 (.BL(BL26),.BLN(BLN26),.WL(WL86));
sram_cell_6t_5 inst_cell_86_27 (.BL(BL27),.BLN(BLN27),.WL(WL86));
sram_cell_6t_5 inst_cell_86_28 (.BL(BL28),.BLN(BLN28),.WL(WL86));
sram_cell_6t_5 inst_cell_86_29 (.BL(BL29),.BLN(BLN29),.WL(WL86));
sram_cell_6t_5 inst_cell_86_30 (.BL(BL30),.BLN(BLN30),.WL(WL86));
sram_cell_6t_5 inst_cell_86_31 (.BL(BL31),.BLN(BLN31),.WL(WL86));
sram_cell_6t_5 inst_cell_86_32 (.BL(BL32),.BLN(BLN32),.WL(WL86));
sram_cell_6t_5 inst_cell_86_33 (.BL(BL33),.BLN(BLN33),.WL(WL86));
sram_cell_6t_5 inst_cell_86_34 (.BL(BL34),.BLN(BLN34),.WL(WL86));
sram_cell_6t_5 inst_cell_86_35 (.BL(BL35),.BLN(BLN35),.WL(WL86));
sram_cell_6t_5 inst_cell_86_36 (.BL(BL36),.BLN(BLN36),.WL(WL86));
sram_cell_6t_5 inst_cell_86_37 (.BL(BL37),.BLN(BLN37),.WL(WL86));
sram_cell_6t_5 inst_cell_86_38 (.BL(BL38),.BLN(BLN38),.WL(WL86));
sram_cell_6t_5 inst_cell_86_39 (.BL(BL39),.BLN(BLN39),.WL(WL86));
sram_cell_6t_5 inst_cell_86_40 (.BL(BL40),.BLN(BLN40),.WL(WL86));
sram_cell_6t_5 inst_cell_86_41 (.BL(BL41),.BLN(BLN41),.WL(WL86));
sram_cell_6t_5 inst_cell_86_42 (.BL(BL42),.BLN(BLN42),.WL(WL86));
sram_cell_6t_5 inst_cell_86_43 (.BL(BL43),.BLN(BLN43),.WL(WL86));
sram_cell_6t_5 inst_cell_86_44 (.BL(BL44),.BLN(BLN44),.WL(WL86));
sram_cell_6t_5 inst_cell_86_45 (.BL(BL45),.BLN(BLN45),.WL(WL86));
sram_cell_6t_5 inst_cell_86_46 (.BL(BL46),.BLN(BLN46),.WL(WL86));
sram_cell_6t_5 inst_cell_86_47 (.BL(BL47),.BLN(BLN47),.WL(WL86));
sram_cell_6t_5 inst_cell_86_48 (.BL(BL48),.BLN(BLN48),.WL(WL86));
sram_cell_6t_5 inst_cell_86_49 (.BL(BL49),.BLN(BLN49),.WL(WL86));
sram_cell_6t_5 inst_cell_86_50 (.BL(BL50),.BLN(BLN50),.WL(WL86));
sram_cell_6t_5 inst_cell_86_51 (.BL(BL51),.BLN(BLN51),.WL(WL86));
sram_cell_6t_5 inst_cell_86_52 (.BL(BL52),.BLN(BLN52),.WL(WL86));
sram_cell_6t_5 inst_cell_86_53 (.BL(BL53),.BLN(BLN53),.WL(WL86));
sram_cell_6t_5 inst_cell_86_54 (.BL(BL54),.BLN(BLN54),.WL(WL86));
sram_cell_6t_5 inst_cell_86_55 (.BL(BL55),.BLN(BLN55),.WL(WL86));
sram_cell_6t_5 inst_cell_86_56 (.BL(BL56),.BLN(BLN56),.WL(WL86));
sram_cell_6t_5 inst_cell_86_57 (.BL(BL57),.BLN(BLN57),.WL(WL86));
sram_cell_6t_5 inst_cell_86_58 (.BL(BL58),.BLN(BLN58),.WL(WL86));
sram_cell_6t_5 inst_cell_86_59 (.BL(BL59),.BLN(BLN59),.WL(WL86));
sram_cell_6t_5 inst_cell_86_60 (.BL(BL60),.BLN(BLN60),.WL(WL86));
sram_cell_6t_5 inst_cell_86_61 (.BL(BL61),.BLN(BLN61),.WL(WL86));
sram_cell_6t_5 inst_cell_86_62 (.BL(BL62),.BLN(BLN62),.WL(WL86));
sram_cell_6t_5 inst_cell_86_63 (.BL(BL63),.BLN(BLN63),.WL(WL86));
sram_cell_6t_5 inst_cell_86_64 (.BL(BL64),.BLN(BLN64),.WL(WL86));
sram_cell_6t_5 inst_cell_86_65 (.BL(BL65),.BLN(BLN65),.WL(WL86));
sram_cell_6t_5 inst_cell_86_66 (.BL(BL66),.BLN(BLN66),.WL(WL86));
sram_cell_6t_5 inst_cell_86_67 (.BL(BL67),.BLN(BLN67),.WL(WL86));
sram_cell_6t_5 inst_cell_86_68 (.BL(BL68),.BLN(BLN68),.WL(WL86));
sram_cell_6t_5 inst_cell_86_69 (.BL(BL69),.BLN(BLN69),.WL(WL86));
sram_cell_6t_5 inst_cell_86_70 (.BL(BL70),.BLN(BLN70),.WL(WL86));
sram_cell_6t_5 inst_cell_86_71 (.BL(BL71),.BLN(BLN71),.WL(WL86));
sram_cell_6t_5 inst_cell_86_72 (.BL(BL72),.BLN(BLN72),.WL(WL86));
sram_cell_6t_5 inst_cell_86_73 (.BL(BL73),.BLN(BLN73),.WL(WL86));
sram_cell_6t_5 inst_cell_86_74 (.BL(BL74),.BLN(BLN74),.WL(WL86));
sram_cell_6t_5 inst_cell_86_75 (.BL(BL75),.BLN(BLN75),.WL(WL86));
sram_cell_6t_5 inst_cell_86_76 (.BL(BL76),.BLN(BLN76),.WL(WL86));
sram_cell_6t_5 inst_cell_86_77 (.BL(BL77),.BLN(BLN77),.WL(WL86));
sram_cell_6t_5 inst_cell_86_78 (.BL(BL78),.BLN(BLN78),.WL(WL86));
sram_cell_6t_5 inst_cell_86_79 (.BL(BL79),.BLN(BLN79),.WL(WL86));
sram_cell_6t_5 inst_cell_86_80 (.BL(BL80),.BLN(BLN80),.WL(WL86));
sram_cell_6t_5 inst_cell_86_81 (.BL(BL81),.BLN(BLN81),.WL(WL86));
sram_cell_6t_5 inst_cell_86_82 (.BL(BL82),.BLN(BLN82),.WL(WL86));
sram_cell_6t_5 inst_cell_86_83 (.BL(BL83),.BLN(BLN83),.WL(WL86));
sram_cell_6t_5 inst_cell_86_84 (.BL(BL84),.BLN(BLN84),.WL(WL86));
sram_cell_6t_5 inst_cell_86_85 (.BL(BL85),.BLN(BLN85),.WL(WL86));
sram_cell_6t_5 inst_cell_86_86 (.BL(BL86),.BLN(BLN86),.WL(WL86));
sram_cell_6t_5 inst_cell_86_87 (.BL(BL87),.BLN(BLN87),.WL(WL86));
sram_cell_6t_5 inst_cell_86_88 (.BL(BL88),.BLN(BLN88),.WL(WL86));
sram_cell_6t_5 inst_cell_86_89 (.BL(BL89),.BLN(BLN89),.WL(WL86));
sram_cell_6t_5 inst_cell_86_90 (.BL(BL90),.BLN(BLN90),.WL(WL86));
sram_cell_6t_5 inst_cell_86_91 (.BL(BL91),.BLN(BLN91),.WL(WL86));
sram_cell_6t_5 inst_cell_86_92 (.BL(BL92),.BLN(BLN92),.WL(WL86));
sram_cell_6t_5 inst_cell_86_93 (.BL(BL93),.BLN(BLN93),.WL(WL86));
sram_cell_6t_5 inst_cell_86_94 (.BL(BL94),.BLN(BLN94),.WL(WL86));
sram_cell_6t_5 inst_cell_86_95 (.BL(BL95),.BLN(BLN95),.WL(WL86));
sram_cell_6t_5 inst_cell_86_96 (.BL(BL96),.BLN(BLN96),.WL(WL86));
sram_cell_6t_5 inst_cell_86_97 (.BL(BL97),.BLN(BLN97),.WL(WL86));
sram_cell_6t_5 inst_cell_86_98 (.BL(BL98),.BLN(BLN98),.WL(WL86));
sram_cell_6t_5 inst_cell_86_99 (.BL(BL99),.BLN(BLN99),.WL(WL86));
sram_cell_6t_5 inst_cell_86_100 (.BL(BL100),.BLN(BLN100),.WL(WL86));
sram_cell_6t_5 inst_cell_86_101 (.BL(BL101),.BLN(BLN101),.WL(WL86));
sram_cell_6t_5 inst_cell_86_102 (.BL(BL102),.BLN(BLN102),.WL(WL86));
sram_cell_6t_5 inst_cell_86_103 (.BL(BL103),.BLN(BLN103),.WL(WL86));
sram_cell_6t_5 inst_cell_86_104 (.BL(BL104),.BLN(BLN104),.WL(WL86));
sram_cell_6t_5 inst_cell_86_105 (.BL(BL105),.BLN(BLN105),.WL(WL86));
sram_cell_6t_5 inst_cell_86_106 (.BL(BL106),.BLN(BLN106),.WL(WL86));
sram_cell_6t_5 inst_cell_86_107 (.BL(BL107),.BLN(BLN107),.WL(WL86));
sram_cell_6t_5 inst_cell_86_108 (.BL(BL108),.BLN(BLN108),.WL(WL86));
sram_cell_6t_5 inst_cell_86_109 (.BL(BL109),.BLN(BLN109),.WL(WL86));
sram_cell_6t_5 inst_cell_86_110 (.BL(BL110),.BLN(BLN110),.WL(WL86));
sram_cell_6t_5 inst_cell_86_111 (.BL(BL111),.BLN(BLN111),.WL(WL86));
sram_cell_6t_5 inst_cell_86_112 (.BL(BL112),.BLN(BLN112),.WL(WL86));
sram_cell_6t_5 inst_cell_86_113 (.BL(BL113),.BLN(BLN113),.WL(WL86));
sram_cell_6t_5 inst_cell_86_114 (.BL(BL114),.BLN(BLN114),.WL(WL86));
sram_cell_6t_5 inst_cell_86_115 (.BL(BL115),.BLN(BLN115),.WL(WL86));
sram_cell_6t_5 inst_cell_86_116 (.BL(BL116),.BLN(BLN116),.WL(WL86));
sram_cell_6t_5 inst_cell_86_117 (.BL(BL117),.BLN(BLN117),.WL(WL86));
sram_cell_6t_5 inst_cell_86_118 (.BL(BL118),.BLN(BLN118),.WL(WL86));
sram_cell_6t_5 inst_cell_86_119 (.BL(BL119),.BLN(BLN119),.WL(WL86));
sram_cell_6t_5 inst_cell_86_120 (.BL(BL120),.BLN(BLN120),.WL(WL86));
sram_cell_6t_5 inst_cell_86_121 (.BL(BL121),.BLN(BLN121),.WL(WL86));
sram_cell_6t_5 inst_cell_86_122 (.BL(BL122),.BLN(BLN122),.WL(WL86));
sram_cell_6t_5 inst_cell_86_123 (.BL(BL123),.BLN(BLN123),.WL(WL86));
sram_cell_6t_5 inst_cell_86_124 (.BL(BL124),.BLN(BLN124),.WL(WL86));
sram_cell_6t_5 inst_cell_86_125 (.BL(BL125),.BLN(BLN125),.WL(WL86));
sram_cell_6t_5 inst_cell_86_126 (.BL(BL126),.BLN(BLN126),.WL(WL86));
sram_cell_6t_5 inst_cell_86_127 (.BL(BL127),.BLN(BLN127),.WL(WL86));
sram_cell_6t_5 inst_cell_87_0 (.BL(BL0),.BLN(BLN0),.WL(WL87));
sram_cell_6t_5 inst_cell_87_1 (.BL(BL1),.BLN(BLN1),.WL(WL87));
sram_cell_6t_5 inst_cell_87_2 (.BL(BL2),.BLN(BLN2),.WL(WL87));
sram_cell_6t_5 inst_cell_87_3 (.BL(BL3),.BLN(BLN3),.WL(WL87));
sram_cell_6t_5 inst_cell_87_4 (.BL(BL4),.BLN(BLN4),.WL(WL87));
sram_cell_6t_5 inst_cell_87_5 (.BL(BL5),.BLN(BLN5),.WL(WL87));
sram_cell_6t_5 inst_cell_87_6 (.BL(BL6),.BLN(BLN6),.WL(WL87));
sram_cell_6t_5 inst_cell_87_7 (.BL(BL7),.BLN(BLN7),.WL(WL87));
sram_cell_6t_5 inst_cell_87_8 (.BL(BL8),.BLN(BLN8),.WL(WL87));
sram_cell_6t_5 inst_cell_87_9 (.BL(BL9),.BLN(BLN9),.WL(WL87));
sram_cell_6t_5 inst_cell_87_10 (.BL(BL10),.BLN(BLN10),.WL(WL87));
sram_cell_6t_5 inst_cell_87_11 (.BL(BL11),.BLN(BLN11),.WL(WL87));
sram_cell_6t_5 inst_cell_87_12 (.BL(BL12),.BLN(BLN12),.WL(WL87));
sram_cell_6t_5 inst_cell_87_13 (.BL(BL13),.BLN(BLN13),.WL(WL87));
sram_cell_6t_5 inst_cell_87_14 (.BL(BL14),.BLN(BLN14),.WL(WL87));
sram_cell_6t_5 inst_cell_87_15 (.BL(BL15),.BLN(BLN15),.WL(WL87));
sram_cell_6t_5 inst_cell_87_16 (.BL(BL16),.BLN(BLN16),.WL(WL87));
sram_cell_6t_5 inst_cell_87_17 (.BL(BL17),.BLN(BLN17),.WL(WL87));
sram_cell_6t_5 inst_cell_87_18 (.BL(BL18),.BLN(BLN18),.WL(WL87));
sram_cell_6t_5 inst_cell_87_19 (.BL(BL19),.BLN(BLN19),.WL(WL87));
sram_cell_6t_5 inst_cell_87_20 (.BL(BL20),.BLN(BLN20),.WL(WL87));
sram_cell_6t_5 inst_cell_87_21 (.BL(BL21),.BLN(BLN21),.WL(WL87));
sram_cell_6t_5 inst_cell_87_22 (.BL(BL22),.BLN(BLN22),.WL(WL87));
sram_cell_6t_5 inst_cell_87_23 (.BL(BL23),.BLN(BLN23),.WL(WL87));
sram_cell_6t_5 inst_cell_87_24 (.BL(BL24),.BLN(BLN24),.WL(WL87));
sram_cell_6t_5 inst_cell_87_25 (.BL(BL25),.BLN(BLN25),.WL(WL87));
sram_cell_6t_5 inst_cell_87_26 (.BL(BL26),.BLN(BLN26),.WL(WL87));
sram_cell_6t_5 inst_cell_87_27 (.BL(BL27),.BLN(BLN27),.WL(WL87));
sram_cell_6t_5 inst_cell_87_28 (.BL(BL28),.BLN(BLN28),.WL(WL87));
sram_cell_6t_5 inst_cell_87_29 (.BL(BL29),.BLN(BLN29),.WL(WL87));
sram_cell_6t_5 inst_cell_87_30 (.BL(BL30),.BLN(BLN30),.WL(WL87));
sram_cell_6t_5 inst_cell_87_31 (.BL(BL31),.BLN(BLN31),.WL(WL87));
sram_cell_6t_5 inst_cell_87_32 (.BL(BL32),.BLN(BLN32),.WL(WL87));
sram_cell_6t_5 inst_cell_87_33 (.BL(BL33),.BLN(BLN33),.WL(WL87));
sram_cell_6t_5 inst_cell_87_34 (.BL(BL34),.BLN(BLN34),.WL(WL87));
sram_cell_6t_5 inst_cell_87_35 (.BL(BL35),.BLN(BLN35),.WL(WL87));
sram_cell_6t_5 inst_cell_87_36 (.BL(BL36),.BLN(BLN36),.WL(WL87));
sram_cell_6t_5 inst_cell_87_37 (.BL(BL37),.BLN(BLN37),.WL(WL87));
sram_cell_6t_5 inst_cell_87_38 (.BL(BL38),.BLN(BLN38),.WL(WL87));
sram_cell_6t_5 inst_cell_87_39 (.BL(BL39),.BLN(BLN39),.WL(WL87));
sram_cell_6t_5 inst_cell_87_40 (.BL(BL40),.BLN(BLN40),.WL(WL87));
sram_cell_6t_5 inst_cell_87_41 (.BL(BL41),.BLN(BLN41),.WL(WL87));
sram_cell_6t_5 inst_cell_87_42 (.BL(BL42),.BLN(BLN42),.WL(WL87));
sram_cell_6t_5 inst_cell_87_43 (.BL(BL43),.BLN(BLN43),.WL(WL87));
sram_cell_6t_5 inst_cell_87_44 (.BL(BL44),.BLN(BLN44),.WL(WL87));
sram_cell_6t_5 inst_cell_87_45 (.BL(BL45),.BLN(BLN45),.WL(WL87));
sram_cell_6t_5 inst_cell_87_46 (.BL(BL46),.BLN(BLN46),.WL(WL87));
sram_cell_6t_5 inst_cell_87_47 (.BL(BL47),.BLN(BLN47),.WL(WL87));
sram_cell_6t_5 inst_cell_87_48 (.BL(BL48),.BLN(BLN48),.WL(WL87));
sram_cell_6t_5 inst_cell_87_49 (.BL(BL49),.BLN(BLN49),.WL(WL87));
sram_cell_6t_5 inst_cell_87_50 (.BL(BL50),.BLN(BLN50),.WL(WL87));
sram_cell_6t_5 inst_cell_87_51 (.BL(BL51),.BLN(BLN51),.WL(WL87));
sram_cell_6t_5 inst_cell_87_52 (.BL(BL52),.BLN(BLN52),.WL(WL87));
sram_cell_6t_5 inst_cell_87_53 (.BL(BL53),.BLN(BLN53),.WL(WL87));
sram_cell_6t_5 inst_cell_87_54 (.BL(BL54),.BLN(BLN54),.WL(WL87));
sram_cell_6t_5 inst_cell_87_55 (.BL(BL55),.BLN(BLN55),.WL(WL87));
sram_cell_6t_5 inst_cell_87_56 (.BL(BL56),.BLN(BLN56),.WL(WL87));
sram_cell_6t_5 inst_cell_87_57 (.BL(BL57),.BLN(BLN57),.WL(WL87));
sram_cell_6t_5 inst_cell_87_58 (.BL(BL58),.BLN(BLN58),.WL(WL87));
sram_cell_6t_5 inst_cell_87_59 (.BL(BL59),.BLN(BLN59),.WL(WL87));
sram_cell_6t_5 inst_cell_87_60 (.BL(BL60),.BLN(BLN60),.WL(WL87));
sram_cell_6t_5 inst_cell_87_61 (.BL(BL61),.BLN(BLN61),.WL(WL87));
sram_cell_6t_5 inst_cell_87_62 (.BL(BL62),.BLN(BLN62),.WL(WL87));
sram_cell_6t_5 inst_cell_87_63 (.BL(BL63),.BLN(BLN63),.WL(WL87));
sram_cell_6t_5 inst_cell_87_64 (.BL(BL64),.BLN(BLN64),.WL(WL87));
sram_cell_6t_5 inst_cell_87_65 (.BL(BL65),.BLN(BLN65),.WL(WL87));
sram_cell_6t_5 inst_cell_87_66 (.BL(BL66),.BLN(BLN66),.WL(WL87));
sram_cell_6t_5 inst_cell_87_67 (.BL(BL67),.BLN(BLN67),.WL(WL87));
sram_cell_6t_5 inst_cell_87_68 (.BL(BL68),.BLN(BLN68),.WL(WL87));
sram_cell_6t_5 inst_cell_87_69 (.BL(BL69),.BLN(BLN69),.WL(WL87));
sram_cell_6t_5 inst_cell_87_70 (.BL(BL70),.BLN(BLN70),.WL(WL87));
sram_cell_6t_5 inst_cell_87_71 (.BL(BL71),.BLN(BLN71),.WL(WL87));
sram_cell_6t_5 inst_cell_87_72 (.BL(BL72),.BLN(BLN72),.WL(WL87));
sram_cell_6t_5 inst_cell_87_73 (.BL(BL73),.BLN(BLN73),.WL(WL87));
sram_cell_6t_5 inst_cell_87_74 (.BL(BL74),.BLN(BLN74),.WL(WL87));
sram_cell_6t_5 inst_cell_87_75 (.BL(BL75),.BLN(BLN75),.WL(WL87));
sram_cell_6t_5 inst_cell_87_76 (.BL(BL76),.BLN(BLN76),.WL(WL87));
sram_cell_6t_5 inst_cell_87_77 (.BL(BL77),.BLN(BLN77),.WL(WL87));
sram_cell_6t_5 inst_cell_87_78 (.BL(BL78),.BLN(BLN78),.WL(WL87));
sram_cell_6t_5 inst_cell_87_79 (.BL(BL79),.BLN(BLN79),.WL(WL87));
sram_cell_6t_5 inst_cell_87_80 (.BL(BL80),.BLN(BLN80),.WL(WL87));
sram_cell_6t_5 inst_cell_87_81 (.BL(BL81),.BLN(BLN81),.WL(WL87));
sram_cell_6t_5 inst_cell_87_82 (.BL(BL82),.BLN(BLN82),.WL(WL87));
sram_cell_6t_5 inst_cell_87_83 (.BL(BL83),.BLN(BLN83),.WL(WL87));
sram_cell_6t_5 inst_cell_87_84 (.BL(BL84),.BLN(BLN84),.WL(WL87));
sram_cell_6t_5 inst_cell_87_85 (.BL(BL85),.BLN(BLN85),.WL(WL87));
sram_cell_6t_5 inst_cell_87_86 (.BL(BL86),.BLN(BLN86),.WL(WL87));
sram_cell_6t_5 inst_cell_87_87 (.BL(BL87),.BLN(BLN87),.WL(WL87));
sram_cell_6t_5 inst_cell_87_88 (.BL(BL88),.BLN(BLN88),.WL(WL87));
sram_cell_6t_5 inst_cell_87_89 (.BL(BL89),.BLN(BLN89),.WL(WL87));
sram_cell_6t_5 inst_cell_87_90 (.BL(BL90),.BLN(BLN90),.WL(WL87));
sram_cell_6t_5 inst_cell_87_91 (.BL(BL91),.BLN(BLN91),.WL(WL87));
sram_cell_6t_5 inst_cell_87_92 (.BL(BL92),.BLN(BLN92),.WL(WL87));
sram_cell_6t_5 inst_cell_87_93 (.BL(BL93),.BLN(BLN93),.WL(WL87));
sram_cell_6t_5 inst_cell_87_94 (.BL(BL94),.BLN(BLN94),.WL(WL87));
sram_cell_6t_5 inst_cell_87_95 (.BL(BL95),.BLN(BLN95),.WL(WL87));
sram_cell_6t_5 inst_cell_87_96 (.BL(BL96),.BLN(BLN96),.WL(WL87));
sram_cell_6t_5 inst_cell_87_97 (.BL(BL97),.BLN(BLN97),.WL(WL87));
sram_cell_6t_5 inst_cell_87_98 (.BL(BL98),.BLN(BLN98),.WL(WL87));
sram_cell_6t_5 inst_cell_87_99 (.BL(BL99),.BLN(BLN99),.WL(WL87));
sram_cell_6t_5 inst_cell_87_100 (.BL(BL100),.BLN(BLN100),.WL(WL87));
sram_cell_6t_5 inst_cell_87_101 (.BL(BL101),.BLN(BLN101),.WL(WL87));
sram_cell_6t_5 inst_cell_87_102 (.BL(BL102),.BLN(BLN102),.WL(WL87));
sram_cell_6t_5 inst_cell_87_103 (.BL(BL103),.BLN(BLN103),.WL(WL87));
sram_cell_6t_5 inst_cell_87_104 (.BL(BL104),.BLN(BLN104),.WL(WL87));
sram_cell_6t_5 inst_cell_87_105 (.BL(BL105),.BLN(BLN105),.WL(WL87));
sram_cell_6t_5 inst_cell_87_106 (.BL(BL106),.BLN(BLN106),.WL(WL87));
sram_cell_6t_5 inst_cell_87_107 (.BL(BL107),.BLN(BLN107),.WL(WL87));
sram_cell_6t_5 inst_cell_87_108 (.BL(BL108),.BLN(BLN108),.WL(WL87));
sram_cell_6t_5 inst_cell_87_109 (.BL(BL109),.BLN(BLN109),.WL(WL87));
sram_cell_6t_5 inst_cell_87_110 (.BL(BL110),.BLN(BLN110),.WL(WL87));
sram_cell_6t_5 inst_cell_87_111 (.BL(BL111),.BLN(BLN111),.WL(WL87));
sram_cell_6t_5 inst_cell_87_112 (.BL(BL112),.BLN(BLN112),.WL(WL87));
sram_cell_6t_5 inst_cell_87_113 (.BL(BL113),.BLN(BLN113),.WL(WL87));
sram_cell_6t_5 inst_cell_87_114 (.BL(BL114),.BLN(BLN114),.WL(WL87));
sram_cell_6t_5 inst_cell_87_115 (.BL(BL115),.BLN(BLN115),.WL(WL87));
sram_cell_6t_5 inst_cell_87_116 (.BL(BL116),.BLN(BLN116),.WL(WL87));
sram_cell_6t_5 inst_cell_87_117 (.BL(BL117),.BLN(BLN117),.WL(WL87));
sram_cell_6t_5 inst_cell_87_118 (.BL(BL118),.BLN(BLN118),.WL(WL87));
sram_cell_6t_5 inst_cell_87_119 (.BL(BL119),.BLN(BLN119),.WL(WL87));
sram_cell_6t_5 inst_cell_87_120 (.BL(BL120),.BLN(BLN120),.WL(WL87));
sram_cell_6t_5 inst_cell_87_121 (.BL(BL121),.BLN(BLN121),.WL(WL87));
sram_cell_6t_5 inst_cell_87_122 (.BL(BL122),.BLN(BLN122),.WL(WL87));
sram_cell_6t_5 inst_cell_87_123 (.BL(BL123),.BLN(BLN123),.WL(WL87));
sram_cell_6t_5 inst_cell_87_124 (.BL(BL124),.BLN(BLN124),.WL(WL87));
sram_cell_6t_5 inst_cell_87_125 (.BL(BL125),.BLN(BLN125),.WL(WL87));
sram_cell_6t_5 inst_cell_87_126 (.BL(BL126),.BLN(BLN126),.WL(WL87));
sram_cell_6t_5 inst_cell_87_127 (.BL(BL127),.BLN(BLN127),.WL(WL87));
sram_cell_6t_5 inst_cell_88_0 (.BL(BL0),.BLN(BLN0),.WL(WL88));
sram_cell_6t_5 inst_cell_88_1 (.BL(BL1),.BLN(BLN1),.WL(WL88));
sram_cell_6t_5 inst_cell_88_2 (.BL(BL2),.BLN(BLN2),.WL(WL88));
sram_cell_6t_5 inst_cell_88_3 (.BL(BL3),.BLN(BLN3),.WL(WL88));
sram_cell_6t_5 inst_cell_88_4 (.BL(BL4),.BLN(BLN4),.WL(WL88));
sram_cell_6t_5 inst_cell_88_5 (.BL(BL5),.BLN(BLN5),.WL(WL88));
sram_cell_6t_5 inst_cell_88_6 (.BL(BL6),.BLN(BLN6),.WL(WL88));
sram_cell_6t_5 inst_cell_88_7 (.BL(BL7),.BLN(BLN7),.WL(WL88));
sram_cell_6t_5 inst_cell_88_8 (.BL(BL8),.BLN(BLN8),.WL(WL88));
sram_cell_6t_5 inst_cell_88_9 (.BL(BL9),.BLN(BLN9),.WL(WL88));
sram_cell_6t_5 inst_cell_88_10 (.BL(BL10),.BLN(BLN10),.WL(WL88));
sram_cell_6t_5 inst_cell_88_11 (.BL(BL11),.BLN(BLN11),.WL(WL88));
sram_cell_6t_5 inst_cell_88_12 (.BL(BL12),.BLN(BLN12),.WL(WL88));
sram_cell_6t_5 inst_cell_88_13 (.BL(BL13),.BLN(BLN13),.WL(WL88));
sram_cell_6t_5 inst_cell_88_14 (.BL(BL14),.BLN(BLN14),.WL(WL88));
sram_cell_6t_5 inst_cell_88_15 (.BL(BL15),.BLN(BLN15),.WL(WL88));
sram_cell_6t_5 inst_cell_88_16 (.BL(BL16),.BLN(BLN16),.WL(WL88));
sram_cell_6t_5 inst_cell_88_17 (.BL(BL17),.BLN(BLN17),.WL(WL88));
sram_cell_6t_5 inst_cell_88_18 (.BL(BL18),.BLN(BLN18),.WL(WL88));
sram_cell_6t_5 inst_cell_88_19 (.BL(BL19),.BLN(BLN19),.WL(WL88));
sram_cell_6t_5 inst_cell_88_20 (.BL(BL20),.BLN(BLN20),.WL(WL88));
sram_cell_6t_5 inst_cell_88_21 (.BL(BL21),.BLN(BLN21),.WL(WL88));
sram_cell_6t_5 inst_cell_88_22 (.BL(BL22),.BLN(BLN22),.WL(WL88));
sram_cell_6t_5 inst_cell_88_23 (.BL(BL23),.BLN(BLN23),.WL(WL88));
sram_cell_6t_5 inst_cell_88_24 (.BL(BL24),.BLN(BLN24),.WL(WL88));
sram_cell_6t_5 inst_cell_88_25 (.BL(BL25),.BLN(BLN25),.WL(WL88));
sram_cell_6t_5 inst_cell_88_26 (.BL(BL26),.BLN(BLN26),.WL(WL88));
sram_cell_6t_5 inst_cell_88_27 (.BL(BL27),.BLN(BLN27),.WL(WL88));
sram_cell_6t_5 inst_cell_88_28 (.BL(BL28),.BLN(BLN28),.WL(WL88));
sram_cell_6t_5 inst_cell_88_29 (.BL(BL29),.BLN(BLN29),.WL(WL88));
sram_cell_6t_5 inst_cell_88_30 (.BL(BL30),.BLN(BLN30),.WL(WL88));
sram_cell_6t_5 inst_cell_88_31 (.BL(BL31),.BLN(BLN31),.WL(WL88));
sram_cell_6t_5 inst_cell_88_32 (.BL(BL32),.BLN(BLN32),.WL(WL88));
sram_cell_6t_5 inst_cell_88_33 (.BL(BL33),.BLN(BLN33),.WL(WL88));
sram_cell_6t_5 inst_cell_88_34 (.BL(BL34),.BLN(BLN34),.WL(WL88));
sram_cell_6t_5 inst_cell_88_35 (.BL(BL35),.BLN(BLN35),.WL(WL88));
sram_cell_6t_5 inst_cell_88_36 (.BL(BL36),.BLN(BLN36),.WL(WL88));
sram_cell_6t_5 inst_cell_88_37 (.BL(BL37),.BLN(BLN37),.WL(WL88));
sram_cell_6t_5 inst_cell_88_38 (.BL(BL38),.BLN(BLN38),.WL(WL88));
sram_cell_6t_5 inst_cell_88_39 (.BL(BL39),.BLN(BLN39),.WL(WL88));
sram_cell_6t_5 inst_cell_88_40 (.BL(BL40),.BLN(BLN40),.WL(WL88));
sram_cell_6t_5 inst_cell_88_41 (.BL(BL41),.BLN(BLN41),.WL(WL88));
sram_cell_6t_5 inst_cell_88_42 (.BL(BL42),.BLN(BLN42),.WL(WL88));
sram_cell_6t_5 inst_cell_88_43 (.BL(BL43),.BLN(BLN43),.WL(WL88));
sram_cell_6t_5 inst_cell_88_44 (.BL(BL44),.BLN(BLN44),.WL(WL88));
sram_cell_6t_5 inst_cell_88_45 (.BL(BL45),.BLN(BLN45),.WL(WL88));
sram_cell_6t_5 inst_cell_88_46 (.BL(BL46),.BLN(BLN46),.WL(WL88));
sram_cell_6t_5 inst_cell_88_47 (.BL(BL47),.BLN(BLN47),.WL(WL88));
sram_cell_6t_5 inst_cell_88_48 (.BL(BL48),.BLN(BLN48),.WL(WL88));
sram_cell_6t_5 inst_cell_88_49 (.BL(BL49),.BLN(BLN49),.WL(WL88));
sram_cell_6t_5 inst_cell_88_50 (.BL(BL50),.BLN(BLN50),.WL(WL88));
sram_cell_6t_5 inst_cell_88_51 (.BL(BL51),.BLN(BLN51),.WL(WL88));
sram_cell_6t_5 inst_cell_88_52 (.BL(BL52),.BLN(BLN52),.WL(WL88));
sram_cell_6t_5 inst_cell_88_53 (.BL(BL53),.BLN(BLN53),.WL(WL88));
sram_cell_6t_5 inst_cell_88_54 (.BL(BL54),.BLN(BLN54),.WL(WL88));
sram_cell_6t_5 inst_cell_88_55 (.BL(BL55),.BLN(BLN55),.WL(WL88));
sram_cell_6t_5 inst_cell_88_56 (.BL(BL56),.BLN(BLN56),.WL(WL88));
sram_cell_6t_5 inst_cell_88_57 (.BL(BL57),.BLN(BLN57),.WL(WL88));
sram_cell_6t_5 inst_cell_88_58 (.BL(BL58),.BLN(BLN58),.WL(WL88));
sram_cell_6t_5 inst_cell_88_59 (.BL(BL59),.BLN(BLN59),.WL(WL88));
sram_cell_6t_5 inst_cell_88_60 (.BL(BL60),.BLN(BLN60),.WL(WL88));
sram_cell_6t_5 inst_cell_88_61 (.BL(BL61),.BLN(BLN61),.WL(WL88));
sram_cell_6t_5 inst_cell_88_62 (.BL(BL62),.BLN(BLN62),.WL(WL88));
sram_cell_6t_5 inst_cell_88_63 (.BL(BL63),.BLN(BLN63),.WL(WL88));
sram_cell_6t_5 inst_cell_88_64 (.BL(BL64),.BLN(BLN64),.WL(WL88));
sram_cell_6t_5 inst_cell_88_65 (.BL(BL65),.BLN(BLN65),.WL(WL88));
sram_cell_6t_5 inst_cell_88_66 (.BL(BL66),.BLN(BLN66),.WL(WL88));
sram_cell_6t_5 inst_cell_88_67 (.BL(BL67),.BLN(BLN67),.WL(WL88));
sram_cell_6t_5 inst_cell_88_68 (.BL(BL68),.BLN(BLN68),.WL(WL88));
sram_cell_6t_5 inst_cell_88_69 (.BL(BL69),.BLN(BLN69),.WL(WL88));
sram_cell_6t_5 inst_cell_88_70 (.BL(BL70),.BLN(BLN70),.WL(WL88));
sram_cell_6t_5 inst_cell_88_71 (.BL(BL71),.BLN(BLN71),.WL(WL88));
sram_cell_6t_5 inst_cell_88_72 (.BL(BL72),.BLN(BLN72),.WL(WL88));
sram_cell_6t_5 inst_cell_88_73 (.BL(BL73),.BLN(BLN73),.WL(WL88));
sram_cell_6t_5 inst_cell_88_74 (.BL(BL74),.BLN(BLN74),.WL(WL88));
sram_cell_6t_5 inst_cell_88_75 (.BL(BL75),.BLN(BLN75),.WL(WL88));
sram_cell_6t_5 inst_cell_88_76 (.BL(BL76),.BLN(BLN76),.WL(WL88));
sram_cell_6t_5 inst_cell_88_77 (.BL(BL77),.BLN(BLN77),.WL(WL88));
sram_cell_6t_5 inst_cell_88_78 (.BL(BL78),.BLN(BLN78),.WL(WL88));
sram_cell_6t_5 inst_cell_88_79 (.BL(BL79),.BLN(BLN79),.WL(WL88));
sram_cell_6t_5 inst_cell_88_80 (.BL(BL80),.BLN(BLN80),.WL(WL88));
sram_cell_6t_5 inst_cell_88_81 (.BL(BL81),.BLN(BLN81),.WL(WL88));
sram_cell_6t_5 inst_cell_88_82 (.BL(BL82),.BLN(BLN82),.WL(WL88));
sram_cell_6t_5 inst_cell_88_83 (.BL(BL83),.BLN(BLN83),.WL(WL88));
sram_cell_6t_5 inst_cell_88_84 (.BL(BL84),.BLN(BLN84),.WL(WL88));
sram_cell_6t_5 inst_cell_88_85 (.BL(BL85),.BLN(BLN85),.WL(WL88));
sram_cell_6t_5 inst_cell_88_86 (.BL(BL86),.BLN(BLN86),.WL(WL88));
sram_cell_6t_5 inst_cell_88_87 (.BL(BL87),.BLN(BLN87),.WL(WL88));
sram_cell_6t_5 inst_cell_88_88 (.BL(BL88),.BLN(BLN88),.WL(WL88));
sram_cell_6t_5 inst_cell_88_89 (.BL(BL89),.BLN(BLN89),.WL(WL88));
sram_cell_6t_5 inst_cell_88_90 (.BL(BL90),.BLN(BLN90),.WL(WL88));
sram_cell_6t_5 inst_cell_88_91 (.BL(BL91),.BLN(BLN91),.WL(WL88));
sram_cell_6t_5 inst_cell_88_92 (.BL(BL92),.BLN(BLN92),.WL(WL88));
sram_cell_6t_5 inst_cell_88_93 (.BL(BL93),.BLN(BLN93),.WL(WL88));
sram_cell_6t_5 inst_cell_88_94 (.BL(BL94),.BLN(BLN94),.WL(WL88));
sram_cell_6t_5 inst_cell_88_95 (.BL(BL95),.BLN(BLN95),.WL(WL88));
sram_cell_6t_5 inst_cell_88_96 (.BL(BL96),.BLN(BLN96),.WL(WL88));
sram_cell_6t_5 inst_cell_88_97 (.BL(BL97),.BLN(BLN97),.WL(WL88));
sram_cell_6t_5 inst_cell_88_98 (.BL(BL98),.BLN(BLN98),.WL(WL88));
sram_cell_6t_5 inst_cell_88_99 (.BL(BL99),.BLN(BLN99),.WL(WL88));
sram_cell_6t_5 inst_cell_88_100 (.BL(BL100),.BLN(BLN100),.WL(WL88));
sram_cell_6t_5 inst_cell_88_101 (.BL(BL101),.BLN(BLN101),.WL(WL88));
sram_cell_6t_5 inst_cell_88_102 (.BL(BL102),.BLN(BLN102),.WL(WL88));
sram_cell_6t_5 inst_cell_88_103 (.BL(BL103),.BLN(BLN103),.WL(WL88));
sram_cell_6t_5 inst_cell_88_104 (.BL(BL104),.BLN(BLN104),.WL(WL88));
sram_cell_6t_5 inst_cell_88_105 (.BL(BL105),.BLN(BLN105),.WL(WL88));
sram_cell_6t_5 inst_cell_88_106 (.BL(BL106),.BLN(BLN106),.WL(WL88));
sram_cell_6t_5 inst_cell_88_107 (.BL(BL107),.BLN(BLN107),.WL(WL88));
sram_cell_6t_5 inst_cell_88_108 (.BL(BL108),.BLN(BLN108),.WL(WL88));
sram_cell_6t_5 inst_cell_88_109 (.BL(BL109),.BLN(BLN109),.WL(WL88));
sram_cell_6t_5 inst_cell_88_110 (.BL(BL110),.BLN(BLN110),.WL(WL88));
sram_cell_6t_5 inst_cell_88_111 (.BL(BL111),.BLN(BLN111),.WL(WL88));
sram_cell_6t_5 inst_cell_88_112 (.BL(BL112),.BLN(BLN112),.WL(WL88));
sram_cell_6t_5 inst_cell_88_113 (.BL(BL113),.BLN(BLN113),.WL(WL88));
sram_cell_6t_5 inst_cell_88_114 (.BL(BL114),.BLN(BLN114),.WL(WL88));
sram_cell_6t_5 inst_cell_88_115 (.BL(BL115),.BLN(BLN115),.WL(WL88));
sram_cell_6t_5 inst_cell_88_116 (.BL(BL116),.BLN(BLN116),.WL(WL88));
sram_cell_6t_5 inst_cell_88_117 (.BL(BL117),.BLN(BLN117),.WL(WL88));
sram_cell_6t_5 inst_cell_88_118 (.BL(BL118),.BLN(BLN118),.WL(WL88));
sram_cell_6t_5 inst_cell_88_119 (.BL(BL119),.BLN(BLN119),.WL(WL88));
sram_cell_6t_5 inst_cell_88_120 (.BL(BL120),.BLN(BLN120),.WL(WL88));
sram_cell_6t_5 inst_cell_88_121 (.BL(BL121),.BLN(BLN121),.WL(WL88));
sram_cell_6t_5 inst_cell_88_122 (.BL(BL122),.BLN(BLN122),.WL(WL88));
sram_cell_6t_5 inst_cell_88_123 (.BL(BL123),.BLN(BLN123),.WL(WL88));
sram_cell_6t_5 inst_cell_88_124 (.BL(BL124),.BLN(BLN124),.WL(WL88));
sram_cell_6t_5 inst_cell_88_125 (.BL(BL125),.BLN(BLN125),.WL(WL88));
sram_cell_6t_5 inst_cell_88_126 (.BL(BL126),.BLN(BLN126),.WL(WL88));
sram_cell_6t_5 inst_cell_88_127 (.BL(BL127),.BLN(BLN127),.WL(WL88));
sram_cell_6t_5 inst_cell_89_0 (.BL(BL0),.BLN(BLN0),.WL(WL89));
sram_cell_6t_5 inst_cell_89_1 (.BL(BL1),.BLN(BLN1),.WL(WL89));
sram_cell_6t_5 inst_cell_89_2 (.BL(BL2),.BLN(BLN2),.WL(WL89));
sram_cell_6t_5 inst_cell_89_3 (.BL(BL3),.BLN(BLN3),.WL(WL89));
sram_cell_6t_5 inst_cell_89_4 (.BL(BL4),.BLN(BLN4),.WL(WL89));
sram_cell_6t_5 inst_cell_89_5 (.BL(BL5),.BLN(BLN5),.WL(WL89));
sram_cell_6t_5 inst_cell_89_6 (.BL(BL6),.BLN(BLN6),.WL(WL89));
sram_cell_6t_5 inst_cell_89_7 (.BL(BL7),.BLN(BLN7),.WL(WL89));
sram_cell_6t_5 inst_cell_89_8 (.BL(BL8),.BLN(BLN8),.WL(WL89));
sram_cell_6t_5 inst_cell_89_9 (.BL(BL9),.BLN(BLN9),.WL(WL89));
sram_cell_6t_5 inst_cell_89_10 (.BL(BL10),.BLN(BLN10),.WL(WL89));
sram_cell_6t_5 inst_cell_89_11 (.BL(BL11),.BLN(BLN11),.WL(WL89));
sram_cell_6t_5 inst_cell_89_12 (.BL(BL12),.BLN(BLN12),.WL(WL89));
sram_cell_6t_5 inst_cell_89_13 (.BL(BL13),.BLN(BLN13),.WL(WL89));
sram_cell_6t_5 inst_cell_89_14 (.BL(BL14),.BLN(BLN14),.WL(WL89));
sram_cell_6t_5 inst_cell_89_15 (.BL(BL15),.BLN(BLN15),.WL(WL89));
sram_cell_6t_5 inst_cell_89_16 (.BL(BL16),.BLN(BLN16),.WL(WL89));
sram_cell_6t_5 inst_cell_89_17 (.BL(BL17),.BLN(BLN17),.WL(WL89));
sram_cell_6t_5 inst_cell_89_18 (.BL(BL18),.BLN(BLN18),.WL(WL89));
sram_cell_6t_5 inst_cell_89_19 (.BL(BL19),.BLN(BLN19),.WL(WL89));
sram_cell_6t_5 inst_cell_89_20 (.BL(BL20),.BLN(BLN20),.WL(WL89));
sram_cell_6t_5 inst_cell_89_21 (.BL(BL21),.BLN(BLN21),.WL(WL89));
sram_cell_6t_5 inst_cell_89_22 (.BL(BL22),.BLN(BLN22),.WL(WL89));
sram_cell_6t_5 inst_cell_89_23 (.BL(BL23),.BLN(BLN23),.WL(WL89));
sram_cell_6t_5 inst_cell_89_24 (.BL(BL24),.BLN(BLN24),.WL(WL89));
sram_cell_6t_5 inst_cell_89_25 (.BL(BL25),.BLN(BLN25),.WL(WL89));
sram_cell_6t_5 inst_cell_89_26 (.BL(BL26),.BLN(BLN26),.WL(WL89));
sram_cell_6t_5 inst_cell_89_27 (.BL(BL27),.BLN(BLN27),.WL(WL89));
sram_cell_6t_5 inst_cell_89_28 (.BL(BL28),.BLN(BLN28),.WL(WL89));
sram_cell_6t_5 inst_cell_89_29 (.BL(BL29),.BLN(BLN29),.WL(WL89));
sram_cell_6t_5 inst_cell_89_30 (.BL(BL30),.BLN(BLN30),.WL(WL89));
sram_cell_6t_5 inst_cell_89_31 (.BL(BL31),.BLN(BLN31),.WL(WL89));
sram_cell_6t_5 inst_cell_89_32 (.BL(BL32),.BLN(BLN32),.WL(WL89));
sram_cell_6t_5 inst_cell_89_33 (.BL(BL33),.BLN(BLN33),.WL(WL89));
sram_cell_6t_5 inst_cell_89_34 (.BL(BL34),.BLN(BLN34),.WL(WL89));
sram_cell_6t_5 inst_cell_89_35 (.BL(BL35),.BLN(BLN35),.WL(WL89));
sram_cell_6t_5 inst_cell_89_36 (.BL(BL36),.BLN(BLN36),.WL(WL89));
sram_cell_6t_5 inst_cell_89_37 (.BL(BL37),.BLN(BLN37),.WL(WL89));
sram_cell_6t_5 inst_cell_89_38 (.BL(BL38),.BLN(BLN38),.WL(WL89));
sram_cell_6t_5 inst_cell_89_39 (.BL(BL39),.BLN(BLN39),.WL(WL89));
sram_cell_6t_5 inst_cell_89_40 (.BL(BL40),.BLN(BLN40),.WL(WL89));
sram_cell_6t_5 inst_cell_89_41 (.BL(BL41),.BLN(BLN41),.WL(WL89));
sram_cell_6t_5 inst_cell_89_42 (.BL(BL42),.BLN(BLN42),.WL(WL89));
sram_cell_6t_5 inst_cell_89_43 (.BL(BL43),.BLN(BLN43),.WL(WL89));
sram_cell_6t_5 inst_cell_89_44 (.BL(BL44),.BLN(BLN44),.WL(WL89));
sram_cell_6t_5 inst_cell_89_45 (.BL(BL45),.BLN(BLN45),.WL(WL89));
sram_cell_6t_5 inst_cell_89_46 (.BL(BL46),.BLN(BLN46),.WL(WL89));
sram_cell_6t_5 inst_cell_89_47 (.BL(BL47),.BLN(BLN47),.WL(WL89));
sram_cell_6t_5 inst_cell_89_48 (.BL(BL48),.BLN(BLN48),.WL(WL89));
sram_cell_6t_5 inst_cell_89_49 (.BL(BL49),.BLN(BLN49),.WL(WL89));
sram_cell_6t_5 inst_cell_89_50 (.BL(BL50),.BLN(BLN50),.WL(WL89));
sram_cell_6t_5 inst_cell_89_51 (.BL(BL51),.BLN(BLN51),.WL(WL89));
sram_cell_6t_5 inst_cell_89_52 (.BL(BL52),.BLN(BLN52),.WL(WL89));
sram_cell_6t_5 inst_cell_89_53 (.BL(BL53),.BLN(BLN53),.WL(WL89));
sram_cell_6t_5 inst_cell_89_54 (.BL(BL54),.BLN(BLN54),.WL(WL89));
sram_cell_6t_5 inst_cell_89_55 (.BL(BL55),.BLN(BLN55),.WL(WL89));
sram_cell_6t_5 inst_cell_89_56 (.BL(BL56),.BLN(BLN56),.WL(WL89));
sram_cell_6t_5 inst_cell_89_57 (.BL(BL57),.BLN(BLN57),.WL(WL89));
sram_cell_6t_5 inst_cell_89_58 (.BL(BL58),.BLN(BLN58),.WL(WL89));
sram_cell_6t_5 inst_cell_89_59 (.BL(BL59),.BLN(BLN59),.WL(WL89));
sram_cell_6t_5 inst_cell_89_60 (.BL(BL60),.BLN(BLN60),.WL(WL89));
sram_cell_6t_5 inst_cell_89_61 (.BL(BL61),.BLN(BLN61),.WL(WL89));
sram_cell_6t_5 inst_cell_89_62 (.BL(BL62),.BLN(BLN62),.WL(WL89));
sram_cell_6t_5 inst_cell_89_63 (.BL(BL63),.BLN(BLN63),.WL(WL89));
sram_cell_6t_5 inst_cell_89_64 (.BL(BL64),.BLN(BLN64),.WL(WL89));
sram_cell_6t_5 inst_cell_89_65 (.BL(BL65),.BLN(BLN65),.WL(WL89));
sram_cell_6t_5 inst_cell_89_66 (.BL(BL66),.BLN(BLN66),.WL(WL89));
sram_cell_6t_5 inst_cell_89_67 (.BL(BL67),.BLN(BLN67),.WL(WL89));
sram_cell_6t_5 inst_cell_89_68 (.BL(BL68),.BLN(BLN68),.WL(WL89));
sram_cell_6t_5 inst_cell_89_69 (.BL(BL69),.BLN(BLN69),.WL(WL89));
sram_cell_6t_5 inst_cell_89_70 (.BL(BL70),.BLN(BLN70),.WL(WL89));
sram_cell_6t_5 inst_cell_89_71 (.BL(BL71),.BLN(BLN71),.WL(WL89));
sram_cell_6t_5 inst_cell_89_72 (.BL(BL72),.BLN(BLN72),.WL(WL89));
sram_cell_6t_5 inst_cell_89_73 (.BL(BL73),.BLN(BLN73),.WL(WL89));
sram_cell_6t_5 inst_cell_89_74 (.BL(BL74),.BLN(BLN74),.WL(WL89));
sram_cell_6t_5 inst_cell_89_75 (.BL(BL75),.BLN(BLN75),.WL(WL89));
sram_cell_6t_5 inst_cell_89_76 (.BL(BL76),.BLN(BLN76),.WL(WL89));
sram_cell_6t_5 inst_cell_89_77 (.BL(BL77),.BLN(BLN77),.WL(WL89));
sram_cell_6t_5 inst_cell_89_78 (.BL(BL78),.BLN(BLN78),.WL(WL89));
sram_cell_6t_5 inst_cell_89_79 (.BL(BL79),.BLN(BLN79),.WL(WL89));
sram_cell_6t_5 inst_cell_89_80 (.BL(BL80),.BLN(BLN80),.WL(WL89));
sram_cell_6t_5 inst_cell_89_81 (.BL(BL81),.BLN(BLN81),.WL(WL89));
sram_cell_6t_5 inst_cell_89_82 (.BL(BL82),.BLN(BLN82),.WL(WL89));
sram_cell_6t_5 inst_cell_89_83 (.BL(BL83),.BLN(BLN83),.WL(WL89));
sram_cell_6t_5 inst_cell_89_84 (.BL(BL84),.BLN(BLN84),.WL(WL89));
sram_cell_6t_5 inst_cell_89_85 (.BL(BL85),.BLN(BLN85),.WL(WL89));
sram_cell_6t_5 inst_cell_89_86 (.BL(BL86),.BLN(BLN86),.WL(WL89));
sram_cell_6t_5 inst_cell_89_87 (.BL(BL87),.BLN(BLN87),.WL(WL89));
sram_cell_6t_5 inst_cell_89_88 (.BL(BL88),.BLN(BLN88),.WL(WL89));
sram_cell_6t_5 inst_cell_89_89 (.BL(BL89),.BLN(BLN89),.WL(WL89));
sram_cell_6t_5 inst_cell_89_90 (.BL(BL90),.BLN(BLN90),.WL(WL89));
sram_cell_6t_5 inst_cell_89_91 (.BL(BL91),.BLN(BLN91),.WL(WL89));
sram_cell_6t_5 inst_cell_89_92 (.BL(BL92),.BLN(BLN92),.WL(WL89));
sram_cell_6t_5 inst_cell_89_93 (.BL(BL93),.BLN(BLN93),.WL(WL89));
sram_cell_6t_5 inst_cell_89_94 (.BL(BL94),.BLN(BLN94),.WL(WL89));
sram_cell_6t_5 inst_cell_89_95 (.BL(BL95),.BLN(BLN95),.WL(WL89));
sram_cell_6t_5 inst_cell_89_96 (.BL(BL96),.BLN(BLN96),.WL(WL89));
sram_cell_6t_5 inst_cell_89_97 (.BL(BL97),.BLN(BLN97),.WL(WL89));
sram_cell_6t_5 inst_cell_89_98 (.BL(BL98),.BLN(BLN98),.WL(WL89));
sram_cell_6t_5 inst_cell_89_99 (.BL(BL99),.BLN(BLN99),.WL(WL89));
sram_cell_6t_5 inst_cell_89_100 (.BL(BL100),.BLN(BLN100),.WL(WL89));
sram_cell_6t_5 inst_cell_89_101 (.BL(BL101),.BLN(BLN101),.WL(WL89));
sram_cell_6t_5 inst_cell_89_102 (.BL(BL102),.BLN(BLN102),.WL(WL89));
sram_cell_6t_5 inst_cell_89_103 (.BL(BL103),.BLN(BLN103),.WL(WL89));
sram_cell_6t_5 inst_cell_89_104 (.BL(BL104),.BLN(BLN104),.WL(WL89));
sram_cell_6t_5 inst_cell_89_105 (.BL(BL105),.BLN(BLN105),.WL(WL89));
sram_cell_6t_5 inst_cell_89_106 (.BL(BL106),.BLN(BLN106),.WL(WL89));
sram_cell_6t_5 inst_cell_89_107 (.BL(BL107),.BLN(BLN107),.WL(WL89));
sram_cell_6t_5 inst_cell_89_108 (.BL(BL108),.BLN(BLN108),.WL(WL89));
sram_cell_6t_5 inst_cell_89_109 (.BL(BL109),.BLN(BLN109),.WL(WL89));
sram_cell_6t_5 inst_cell_89_110 (.BL(BL110),.BLN(BLN110),.WL(WL89));
sram_cell_6t_5 inst_cell_89_111 (.BL(BL111),.BLN(BLN111),.WL(WL89));
sram_cell_6t_5 inst_cell_89_112 (.BL(BL112),.BLN(BLN112),.WL(WL89));
sram_cell_6t_5 inst_cell_89_113 (.BL(BL113),.BLN(BLN113),.WL(WL89));
sram_cell_6t_5 inst_cell_89_114 (.BL(BL114),.BLN(BLN114),.WL(WL89));
sram_cell_6t_5 inst_cell_89_115 (.BL(BL115),.BLN(BLN115),.WL(WL89));
sram_cell_6t_5 inst_cell_89_116 (.BL(BL116),.BLN(BLN116),.WL(WL89));
sram_cell_6t_5 inst_cell_89_117 (.BL(BL117),.BLN(BLN117),.WL(WL89));
sram_cell_6t_5 inst_cell_89_118 (.BL(BL118),.BLN(BLN118),.WL(WL89));
sram_cell_6t_5 inst_cell_89_119 (.BL(BL119),.BLN(BLN119),.WL(WL89));
sram_cell_6t_5 inst_cell_89_120 (.BL(BL120),.BLN(BLN120),.WL(WL89));
sram_cell_6t_5 inst_cell_89_121 (.BL(BL121),.BLN(BLN121),.WL(WL89));
sram_cell_6t_5 inst_cell_89_122 (.BL(BL122),.BLN(BLN122),.WL(WL89));
sram_cell_6t_5 inst_cell_89_123 (.BL(BL123),.BLN(BLN123),.WL(WL89));
sram_cell_6t_5 inst_cell_89_124 (.BL(BL124),.BLN(BLN124),.WL(WL89));
sram_cell_6t_5 inst_cell_89_125 (.BL(BL125),.BLN(BLN125),.WL(WL89));
sram_cell_6t_5 inst_cell_89_126 (.BL(BL126),.BLN(BLN126),.WL(WL89));
sram_cell_6t_5 inst_cell_89_127 (.BL(BL127),.BLN(BLN127),.WL(WL89));
sram_cell_6t_5 inst_cell_90_0 (.BL(BL0),.BLN(BLN0),.WL(WL90));
sram_cell_6t_5 inst_cell_90_1 (.BL(BL1),.BLN(BLN1),.WL(WL90));
sram_cell_6t_5 inst_cell_90_2 (.BL(BL2),.BLN(BLN2),.WL(WL90));
sram_cell_6t_5 inst_cell_90_3 (.BL(BL3),.BLN(BLN3),.WL(WL90));
sram_cell_6t_5 inst_cell_90_4 (.BL(BL4),.BLN(BLN4),.WL(WL90));
sram_cell_6t_5 inst_cell_90_5 (.BL(BL5),.BLN(BLN5),.WL(WL90));
sram_cell_6t_5 inst_cell_90_6 (.BL(BL6),.BLN(BLN6),.WL(WL90));
sram_cell_6t_5 inst_cell_90_7 (.BL(BL7),.BLN(BLN7),.WL(WL90));
sram_cell_6t_5 inst_cell_90_8 (.BL(BL8),.BLN(BLN8),.WL(WL90));
sram_cell_6t_5 inst_cell_90_9 (.BL(BL9),.BLN(BLN9),.WL(WL90));
sram_cell_6t_5 inst_cell_90_10 (.BL(BL10),.BLN(BLN10),.WL(WL90));
sram_cell_6t_5 inst_cell_90_11 (.BL(BL11),.BLN(BLN11),.WL(WL90));
sram_cell_6t_5 inst_cell_90_12 (.BL(BL12),.BLN(BLN12),.WL(WL90));
sram_cell_6t_5 inst_cell_90_13 (.BL(BL13),.BLN(BLN13),.WL(WL90));
sram_cell_6t_5 inst_cell_90_14 (.BL(BL14),.BLN(BLN14),.WL(WL90));
sram_cell_6t_5 inst_cell_90_15 (.BL(BL15),.BLN(BLN15),.WL(WL90));
sram_cell_6t_5 inst_cell_90_16 (.BL(BL16),.BLN(BLN16),.WL(WL90));
sram_cell_6t_5 inst_cell_90_17 (.BL(BL17),.BLN(BLN17),.WL(WL90));
sram_cell_6t_5 inst_cell_90_18 (.BL(BL18),.BLN(BLN18),.WL(WL90));
sram_cell_6t_5 inst_cell_90_19 (.BL(BL19),.BLN(BLN19),.WL(WL90));
sram_cell_6t_5 inst_cell_90_20 (.BL(BL20),.BLN(BLN20),.WL(WL90));
sram_cell_6t_5 inst_cell_90_21 (.BL(BL21),.BLN(BLN21),.WL(WL90));
sram_cell_6t_5 inst_cell_90_22 (.BL(BL22),.BLN(BLN22),.WL(WL90));
sram_cell_6t_5 inst_cell_90_23 (.BL(BL23),.BLN(BLN23),.WL(WL90));
sram_cell_6t_5 inst_cell_90_24 (.BL(BL24),.BLN(BLN24),.WL(WL90));
sram_cell_6t_5 inst_cell_90_25 (.BL(BL25),.BLN(BLN25),.WL(WL90));
sram_cell_6t_5 inst_cell_90_26 (.BL(BL26),.BLN(BLN26),.WL(WL90));
sram_cell_6t_5 inst_cell_90_27 (.BL(BL27),.BLN(BLN27),.WL(WL90));
sram_cell_6t_5 inst_cell_90_28 (.BL(BL28),.BLN(BLN28),.WL(WL90));
sram_cell_6t_5 inst_cell_90_29 (.BL(BL29),.BLN(BLN29),.WL(WL90));
sram_cell_6t_5 inst_cell_90_30 (.BL(BL30),.BLN(BLN30),.WL(WL90));
sram_cell_6t_5 inst_cell_90_31 (.BL(BL31),.BLN(BLN31),.WL(WL90));
sram_cell_6t_5 inst_cell_90_32 (.BL(BL32),.BLN(BLN32),.WL(WL90));
sram_cell_6t_5 inst_cell_90_33 (.BL(BL33),.BLN(BLN33),.WL(WL90));
sram_cell_6t_5 inst_cell_90_34 (.BL(BL34),.BLN(BLN34),.WL(WL90));
sram_cell_6t_5 inst_cell_90_35 (.BL(BL35),.BLN(BLN35),.WL(WL90));
sram_cell_6t_5 inst_cell_90_36 (.BL(BL36),.BLN(BLN36),.WL(WL90));
sram_cell_6t_5 inst_cell_90_37 (.BL(BL37),.BLN(BLN37),.WL(WL90));
sram_cell_6t_5 inst_cell_90_38 (.BL(BL38),.BLN(BLN38),.WL(WL90));
sram_cell_6t_5 inst_cell_90_39 (.BL(BL39),.BLN(BLN39),.WL(WL90));
sram_cell_6t_5 inst_cell_90_40 (.BL(BL40),.BLN(BLN40),.WL(WL90));
sram_cell_6t_5 inst_cell_90_41 (.BL(BL41),.BLN(BLN41),.WL(WL90));
sram_cell_6t_5 inst_cell_90_42 (.BL(BL42),.BLN(BLN42),.WL(WL90));
sram_cell_6t_5 inst_cell_90_43 (.BL(BL43),.BLN(BLN43),.WL(WL90));
sram_cell_6t_5 inst_cell_90_44 (.BL(BL44),.BLN(BLN44),.WL(WL90));
sram_cell_6t_5 inst_cell_90_45 (.BL(BL45),.BLN(BLN45),.WL(WL90));
sram_cell_6t_5 inst_cell_90_46 (.BL(BL46),.BLN(BLN46),.WL(WL90));
sram_cell_6t_5 inst_cell_90_47 (.BL(BL47),.BLN(BLN47),.WL(WL90));
sram_cell_6t_5 inst_cell_90_48 (.BL(BL48),.BLN(BLN48),.WL(WL90));
sram_cell_6t_5 inst_cell_90_49 (.BL(BL49),.BLN(BLN49),.WL(WL90));
sram_cell_6t_5 inst_cell_90_50 (.BL(BL50),.BLN(BLN50),.WL(WL90));
sram_cell_6t_5 inst_cell_90_51 (.BL(BL51),.BLN(BLN51),.WL(WL90));
sram_cell_6t_5 inst_cell_90_52 (.BL(BL52),.BLN(BLN52),.WL(WL90));
sram_cell_6t_5 inst_cell_90_53 (.BL(BL53),.BLN(BLN53),.WL(WL90));
sram_cell_6t_5 inst_cell_90_54 (.BL(BL54),.BLN(BLN54),.WL(WL90));
sram_cell_6t_5 inst_cell_90_55 (.BL(BL55),.BLN(BLN55),.WL(WL90));
sram_cell_6t_5 inst_cell_90_56 (.BL(BL56),.BLN(BLN56),.WL(WL90));
sram_cell_6t_5 inst_cell_90_57 (.BL(BL57),.BLN(BLN57),.WL(WL90));
sram_cell_6t_5 inst_cell_90_58 (.BL(BL58),.BLN(BLN58),.WL(WL90));
sram_cell_6t_5 inst_cell_90_59 (.BL(BL59),.BLN(BLN59),.WL(WL90));
sram_cell_6t_5 inst_cell_90_60 (.BL(BL60),.BLN(BLN60),.WL(WL90));
sram_cell_6t_5 inst_cell_90_61 (.BL(BL61),.BLN(BLN61),.WL(WL90));
sram_cell_6t_5 inst_cell_90_62 (.BL(BL62),.BLN(BLN62),.WL(WL90));
sram_cell_6t_5 inst_cell_90_63 (.BL(BL63),.BLN(BLN63),.WL(WL90));
sram_cell_6t_5 inst_cell_90_64 (.BL(BL64),.BLN(BLN64),.WL(WL90));
sram_cell_6t_5 inst_cell_90_65 (.BL(BL65),.BLN(BLN65),.WL(WL90));
sram_cell_6t_5 inst_cell_90_66 (.BL(BL66),.BLN(BLN66),.WL(WL90));
sram_cell_6t_5 inst_cell_90_67 (.BL(BL67),.BLN(BLN67),.WL(WL90));
sram_cell_6t_5 inst_cell_90_68 (.BL(BL68),.BLN(BLN68),.WL(WL90));
sram_cell_6t_5 inst_cell_90_69 (.BL(BL69),.BLN(BLN69),.WL(WL90));
sram_cell_6t_5 inst_cell_90_70 (.BL(BL70),.BLN(BLN70),.WL(WL90));
sram_cell_6t_5 inst_cell_90_71 (.BL(BL71),.BLN(BLN71),.WL(WL90));
sram_cell_6t_5 inst_cell_90_72 (.BL(BL72),.BLN(BLN72),.WL(WL90));
sram_cell_6t_5 inst_cell_90_73 (.BL(BL73),.BLN(BLN73),.WL(WL90));
sram_cell_6t_5 inst_cell_90_74 (.BL(BL74),.BLN(BLN74),.WL(WL90));
sram_cell_6t_5 inst_cell_90_75 (.BL(BL75),.BLN(BLN75),.WL(WL90));
sram_cell_6t_5 inst_cell_90_76 (.BL(BL76),.BLN(BLN76),.WL(WL90));
sram_cell_6t_5 inst_cell_90_77 (.BL(BL77),.BLN(BLN77),.WL(WL90));
sram_cell_6t_5 inst_cell_90_78 (.BL(BL78),.BLN(BLN78),.WL(WL90));
sram_cell_6t_5 inst_cell_90_79 (.BL(BL79),.BLN(BLN79),.WL(WL90));
sram_cell_6t_5 inst_cell_90_80 (.BL(BL80),.BLN(BLN80),.WL(WL90));
sram_cell_6t_5 inst_cell_90_81 (.BL(BL81),.BLN(BLN81),.WL(WL90));
sram_cell_6t_5 inst_cell_90_82 (.BL(BL82),.BLN(BLN82),.WL(WL90));
sram_cell_6t_5 inst_cell_90_83 (.BL(BL83),.BLN(BLN83),.WL(WL90));
sram_cell_6t_5 inst_cell_90_84 (.BL(BL84),.BLN(BLN84),.WL(WL90));
sram_cell_6t_5 inst_cell_90_85 (.BL(BL85),.BLN(BLN85),.WL(WL90));
sram_cell_6t_5 inst_cell_90_86 (.BL(BL86),.BLN(BLN86),.WL(WL90));
sram_cell_6t_5 inst_cell_90_87 (.BL(BL87),.BLN(BLN87),.WL(WL90));
sram_cell_6t_5 inst_cell_90_88 (.BL(BL88),.BLN(BLN88),.WL(WL90));
sram_cell_6t_5 inst_cell_90_89 (.BL(BL89),.BLN(BLN89),.WL(WL90));
sram_cell_6t_5 inst_cell_90_90 (.BL(BL90),.BLN(BLN90),.WL(WL90));
sram_cell_6t_5 inst_cell_90_91 (.BL(BL91),.BLN(BLN91),.WL(WL90));
sram_cell_6t_5 inst_cell_90_92 (.BL(BL92),.BLN(BLN92),.WL(WL90));
sram_cell_6t_5 inst_cell_90_93 (.BL(BL93),.BLN(BLN93),.WL(WL90));
sram_cell_6t_5 inst_cell_90_94 (.BL(BL94),.BLN(BLN94),.WL(WL90));
sram_cell_6t_5 inst_cell_90_95 (.BL(BL95),.BLN(BLN95),.WL(WL90));
sram_cell_6t_5 inst_cell_90_96 (.BL(BL96),.BLN(BLN96),.WL(WL90));
sram_cell_6t_5 inst_cell_90_97 (.BL(BL97),.BLN(BLN97),.WL(WL90));
sram_cell_6t_5 inst_cell_90_98 (.BL(BL98),.BLN(BLN98),.WL(WL90));
sram_cell_6t_5 inst_cell_90_99 (.BL(BL99),.BLN(BLN99),.WL(WL90));
sram_cell_6t_5 inst_cell_90_100 (.BL(BL100),.BLN(BLN100),.WL(WL90));
sram_cell_6t_5 inst_cell_90_101 (.BL(BL101),.BLN(BLN101),.WL(WL90));
sram_cell_6t_5 inst_cell_90_102 (.BL(BL102),.BLN(BLN102),.WL(WL90));
sram_cell_6t_5 inst_cell_90_103 (.BL(BL103),.BLN(BLN103),.WL(WL90));
sram_cell_6t_5 inst_cell_90_104 (.BL(BL104),.BLN(BLN104),.WL(WL90));
sram_cell_6t_5 inst_cell_90_105 (.BL(BL105),.BLN(BLN105),.WL(WL90));
sram_cell_6t_5 inst_cell_90_106 (.BL(BL106),.BLN(BLN106),.WL(WL90));
sram_cell_6t_5 inst_cell_90_107 (.BL(BL107),.BLN(BLN107),.WL(WL90));
sram_cell_6t_5 inst_cell_90_108 (.BL(BL108),.BLN(BLN108),.WL(WL90));
sram_cell_6t_5 inst_cell_90_109 (.BL(BL109),.BLN(BLN109),.WL(WL90));
sram_cell_6t_5 inst_cell_90_110 (.BL(BL110),.BLN(BLN110),.WL(WL90));
sram_cell_6t_5 inst_cell_90_111 (.BL(BL111),.BLN(BLN111),.WL(WL90));
sram_cell_6t_5 inst_cell_90_112 (.BL(BL112),.BLN(BLN112),.WL(WL90));
sram_cell_6t_5 inst_cell_90_113 (.BL(BL113),.BLN(BLN113),.WL(WL90));
sram_cell_6t_5 inst_cell_90_114 (.BL(BL114),.BLN(BLN114),.WL(WL90));
sram_cell_6t_5 inst_cell_90_115 (.BL(BL115),.BLN(BLN115),.WL(WL90));
sram_cell_6t_5 inst_cell_90_116 (.BL(BL116),.BLN(BLN116),.WL(WL90));
sram_cell_6t_5 inst_cell_90_117 (.BL(BL117),.BLN(BLN117),.WL(WL90));
sram_cell_6t_5 inst_cell_90_118 (.BL(BL118),.BLN(BLN118),.WL(WL90));
sram_cell_6t_5 inst_cell_90_119 (.BL(BL119),.BLN(BLN119),.WL(WL90));
sram_cell_6t_5 inst_cell_90_120 (.BL(BL120),.BLN(BLN120),.WL(WL90));
sram_cell_6t_5 inst_cell_90_121 (.BL(BL121),.BLN(BLN121),.WL(WL90));
sram_cell_6t_5 inst_cell_90_122 (.BL(BL122),.BLN(BLN122),.WL(WL90));
sram_cell_6t_5 inst_cell_90_123 (.BL(BL123),.BLN(BLN123),.WL(WL90));
sram_cell_6t_5 inst_cell_90_124 (.BL(BL124),.BLN(BLN124),.WL(WL90));
sram_cell_6t_5 inst_cell_90_125 (.BL(BL125),.BLN(BLN125),.WL(WL90));
sram_cell_6t_5 inst_cell_90_126 (.BL(BL126),.BLN(BLN126),.WL(WL90));
sram_cell_6t_5 inst_cell_90_127 (.BL(BL127),.BLN(BLN127),.WL(WL90));
sram_cell_6t_5 inst_cell_91_0 (.BL(BL0),.BLN(BLN0),.WL(WL91));
sram_cell_6t_5 inst_cell_91_1 (.BL(BL1),.BLN(BLN1),.WL(WL91));
sram_cell_6t_5 inst_cell_91_2 (.BL(BL2),.BLN(BLN2),.WL(WL91));
sram_cell_6t_5 inst_cell_91_3 (.BL(BL3),.BLN(BLN3),.WL(WL91));
sram_cell_6t_5 inst_cell_91_4 (.BL(BL4),.BLN(BLN4),.WL(WL91));
sram_cell_6t_5 inst_cell_91_5 (.BL(BL5),.BLN(BLN5),.WL(WL91));
sram_cell_6t_5 inst_cell_91_6 (.BL(BL6),.BLN(BLN6),.WL(WL91));
sram_cell_6t_5 inst_cell_91_7 (.BL(BL7),.BLN(BLN7),.WL(WL91));
sram_cell_6t_5 inst_cell_91_8 (.BL(BL8),.BLN(BLN8),.WL(WL91));
sram_cell_6t_5 inst_cell_91_9 (.BL(BL9),.BLN(BLN9),.WL(WL91));
sram_cell_6t_5 inst_cell_91_10 (.BL(BL10),.BLN(BLN10),.WL(WL91));
sram_cell_6t_5 inst_cell_91_11 (.BL(BL11),.BLN(BLN11),.WL(WL91));
sram_cell_6t_5 inst_cell_91_12 (.BL(BL12),.BLN(BLN12),.WL(WL91));
sram_cell_6t_5 inst_cell_91_13 (.BL(BL13),.BLN(BLN13),.WL(WL91));
sram_cell_6t_5 inst_cell_91_14 (.BL(BL14),.BLN(BLN14),.WL(WL91));
sram_cell_6t_5 inst_cell_91_15 (.BL(BL15),.BLN(BLN15),.WL(WL91));
sram_cell_6t_5 inst_cell_91_16 (.BL(BL16),.BLN(BLN16),.WL(WL91));
sram_cell_6t_5 inst_cell_91_17 (.BL(BL17),.BLN(BLN17),.WL(WL91));
sram_cell_6t_5 inst_cell_91_18 (.BL(BL18),.BLN(BLN18),.WL(WL91));
sram_cell_6t_5 inst_cell_91_19 (.BL(BL19),.BLN(BLN19),.WL(WL91));
sram_cell_6t_5 inst_cell_91_20 (.BL(BL20),.BLN(BLN20),.WL(WL91));
sram_cell_6t_5 inst_cell_91_21 (.BL(BL21),.BLN(BLN21),.WL(WL91));
sram_cell_6t_5 inst_cell_91_22 (.BL(BL22),.BLN(BLN22),.WL(WL91));
sram_cell_6t_5 inst_cell_91_23 (.BL(BL23),.BLN(BLN23),.WL(WL91));
sram_cell_6t_5 inst_cell_91_24 (.BL(BL24),.BLN(BLN24),.WL(WL91));
sram_cell_6t_5 inst_cell_91_25 (.BL(BL25),.BLN(BLN25),.WL(WL91));
sram_cell_6t_5 inst_cell_91_26 (.BL(BL26),.BLN(BLN26),.WL(WL91));
sram_cell_6t_5 inst_cell_91_27 (.BL(BL27),.BLN(BLN27),.WL(WL91));
sram_cell_6t_5 inst_cell_91_28 (.BL(BL28),.BLN(BLN28),.WL(WL91));
sram_cell_6t_5 inst_cell_91_29 (.BL(BL29),.BLN(BLN29),.WL(WL91));
sram_cell_6t_5 inst_cell_91_30 (.BL(BL30),.BLN(BLN30),.WL(WL91));
sram_cell_6t_5 inst_cell_91_31 (.BL(BL31),.BLN(BLN31),.WL(WL91));
sram_cell_6t_5 inst_cell_91_32 (.BL(BL32),.BLN(BLN32),.WL(WL91));
sram_cell_6t_5 inst_cell_91_33 (.BL(BL33),.BLN(BLN33),.WL(WL91));
sram_cell_6t_5 inst_cell_91_34 (.BL(BL34),.BLN(BLN34),.WL(WL91));
sram_cell_6t_5 inst_cell_91_35 (.BL(BL35),.BLN(BLN35),.WL(WL91));
sram_cell_6t_5 inst_cell_91_36 (.BL(BL36),.BLN(BLN36),.WL(WL91));
sram_cell_6t_5 inst_cell_91_37 (.BL(BL37),.BLN(BLN37),.WL(WL91));
sram_cell_6t_5 inst_cell_91_38 (.BL(BL38),.BLN(BLN38),.WL(WL91));
sram_cell_6t_5 inst_cell_91_39 (.BL(BL39),.BLN(BLN39),.WL(WL91));
sram_cell_6t_5 inst_cell_91_40 (.BL(BL40),.BLN(BLN40),.WL(WL91));
sram_cell_6t_5 inst_cell_91_41 (.BL(BL41),.BLN(BLN41),.WL(WL91));
sram_cell_6t_5 inst_cell_91_42 (.BL(BL42),.BLN(BLN42),.WL(WL91));
sram_cell_6t_5 inst_cell_91_43 (.BL(BL43),.BLN(BLN43),.WL(WL91));
sram_cell_6t_5 inst_cell_91_44 (.BL(BL44),.BLN(BLN44),.WL(WL91));
sram_cell_6t_5 inst_cell_91_45 (.BL(BL45),.BLN(BLN45),.WL(WL91));
sram_cell_6t_5 inst_cell_91_46 (.BL(BL46),.BLN(BLN46),.WL(WL91));
sram_cell_6t_5 inst_cell_91_47 (.BL(BL47),.BLN(BLN47),.WL(WL91));
sram_cell_6t_5 inst_cell_91_48 (.BL(BL48),.BLN(BLN48),.WL(WL91));
sram_cell_6t_5 inst_cell_91_49 (.BL(BL49),.BLN(BLN49),.WL(WL91));
sram_cell_6t_5 inst_cell_91_50 (.BL(BL50),.BLN(BLN50),.WL(WL91));
sram_cell_6t_5 inst_cell_91_51 (.BL(BL51),.BLN(BLN51),.WL(WL91));
sram_cell_6t_5 inst_cell_91_52 (.BL(BL52),.BLN(BLN52),.WL(WL91));
sram_cell_6t_5 inst_cell_91_53 (.BL(BL53),.BLN(BLN53),.WL(WL91));
sram_cell_6t_5 inst_cell_91_54 (.BL(BL54),.BLN(BLN54),.WL(WL91));
sram_cell_6t_5 inst_cell_91_55 (.BL(BL55),.BLN(BLN55),.WL(WL91));
sram_cell_6t_5 inst_cell_91_56 (.BL(BL56),.BLN(BLN56),.WL(WL91));
sram_cell_6t_5 inst_cell_91_57 (.BL(BL57),.BLN(BLN57),.WL(WL91));
sram_cell_6t_5 inst_cell_91_58 (.BL(BL58),.BLN(BLN58),.WL(WL91));
sram_cell_6t_5 inst_cell_91_59 (.BL(BL59),.BLN(BLN59),.WL(WL91));
sram_cell_6t_5 inst_cell_91_60 (.BL(BL60),.BLN(BLN60),.WL(WL91));
sram_cell_6t_5 inst_cell_91_61 (.BL(BL61),.BLN(BLN61),.WL(WL91));
sram_cell_6t_5 inst_cell_91_62 (.BL(BL62),.BLN(BLN62),.WL(WL91));
sram_cell_6t_5 inst_cell_91_63 (.BL(BL63),.BLN(BLN63),.WL(WL91));
sram_cell_6t_5 inst_cell_91_64 (.BL(BL64),.BLN(BLN64),.WL(WL91));
sram_cell_6t_5 inst_cell_91_65 (.BL(BL65),.BLN(BLN65),.WL(WL91));
sram_cell_6t_5 inst_cell_91_66 (.BL(BL66),.BLN(BLN66),.WL(WL91));
sram_cell_6t_5 inst_cell_91_67 (.BL(BL67),.BLN(BLN67),.WL(WL91));
sram_cell_6t_5 inst_cell_91_68 (.BL(BL68),.BLN(BLN68),.WL(WL91));
sram_cell_6t_5 inst_cell_91_69 (.BL(BL69),.BLN(BLN69),.WL(WL91));
sram_cell_6t_5 inst_cell_91_70 (.BL(BL70),.BLN(BLN70),.WL(WL91));
sram_cell_6t_5 inst_cell_91_71 (.BL(BL71),.BLN(BLN71),.WL(WL91));
sram_cell_6t_5 inst_cell_91_72 (.BL(BL72),.BLN(BLN72),.WL(WL91));
sram_cell_6t_5 inst_cell_91_73 (.BL(BL73),.BLN(BLN73),.WL(WL91));
sram_cell_6t_5 inst_cell_91_74 (.BL(BL74),.BLN(BLN74),.WL(WL91));
sram_cell_6t_5 inst_cell_91_75 (.BL(BL75),.BLN(BLN75),.WL(WL91));
sram_cell_6t_5 inst_cell_91_76 (.BL(BL76),.BLN(BLN76),.WL(WL91));
sram_cell_6t_5 inst_cell_91_77 (.BL(BL77),.BLN(BLN77),.WL(WL91));
sram_cell_6t_5 inst_cell_91_78 (.BL(BL78),.BLN(BLN78),.WL(WL91));
sram_cell_6t_5 inst_cell_91_79 (.BL(BL79),.BLN(BLN79),.WL(WL91));
sram_cell_6t_5 inst_cell_91_80 (.BL(BL80),.BLN(BLN80),.WL(WL91));
sram_cell_6t_5 inst_cell_91_81 (.BL(BL81),.BLN(BLN81),.WL(WL91));
sram_cell_6t_5 inst_cell_91_82 (.BL(BL82),.BLN(BLN82),.WL(WL91));
sram_cell_6t_5 inst_cell_91_83 (.BL(BL83),.BLN(BLN83),.WL(WL91));
sram_cell_6t_5 inst_cell_91_84 (.BL(BL84),.BLN(BLN84),.WL(WL91));
sram_cell_6t_5 inst_cell_91_85 (.BL(BL85),.BLN(BLN85),.WL(WL91));
sram_cell_6t_5 inst_cell_91_86 (.BL(BL86),.BLN(BLN86),.WL(WL91));
sram_cell_6t_5 inst_cell_91_87 (.BL(BL87),.BLN(BLN87),.WL(WL91));
sram_cell_6t_5 inst_cell_91_88 (.BL(BL88),.BLN(BLN88),.WL(WL91));
sram_cell_6t_5 inst_cell_91_89 (.BL(BL89),.BLN(BLN89),.WL(WL91));
sram_cell_6t_5 inst_cell_91_90 (.BL(BL90),.BLN(BLN90),.WL(WL91));
sram_cell_6t_5 inst_cell_91_91 (.BL(BL91),.BLN(BLN91),.WL(WL91));
sram_cell_6t_5 inst_cell_91_92 (.BL(BL92),.BLN(BLN92),.WL(WL91));
sram_cell_6t_5 inst_cell_91_93 (.BL(BL93),.BLN(BLN93),.WL(WL91));
sram_cell_6t_5 inst_cell_91_94 (.BL(BL94),.BLN(BLN94),.WL(WL91));
sram_cell_6t_5 inst_cell_91_95 (.BL(BL95),.BLN(BLN95),.WL(WL91));
sram_cell_6t_5 inst_cell_91_96 (.BL(BL96),.BLN(BLN96),.WL(WL91));
sram_cell_6t_5 inst_cell_91_97 (.BL(BL97),.BLN(BLN97),.WL(WL91));
sram_cell_6t_5 inst_cell_91_98 (.BL(BL98),.BLN(BLN98),.WL(WL91));
sram_cell_6t_5 inst_cell_91_99 (.BL(BL99),.BLN(BLN99),.WL(WL91));
sram_cell_6t_5 inst_cell_91_100 (.BL(BL100),.BLN(BLN100),.WL(WL91));
sram_cell_6t_5 inst_cell_91_101 (.BL(BL101),.BLN(BLN101),.WL(WL91));
sram_cell_6t_5 inst_cell_91_102 (.BL(BL102),.BLN(BLN102),.WL(WL91));
sram_cell_6t_5 inst_cell_91_103 (.BL(BL103),.BLN(BLN103),.WL(WL91));
sram_cell_6t_5 inst_cell_91_104 (.BL(BL104),.BLN(BLN104),.WL(WL91));
sram_cell_6t_5 inst_cell_91_105 (.BL(BL105),.BLN(BLN105),.WL(WL91));
sram_cell_6t_5 inst_cell_91_106 (.BL(BL106),.BLN(BLN106),.WL(WL91));
sram_cell_6t_5 inst_cell_91_107 (.BL(BL107),.BLN(BLN107),.WL(WL91));
sram_cell_6t_5 inst_cell_91_108 (.BL(BL108),.BLN(BLN108),.WL(WL91));
sram_cell_6t_5 inst_cell_91_109 (.BL(BL109),.BLN(BLN109),.WL(WL91));
sram_cell_6t_5 inst_cell_91_110 (.BL(BL110),.BLN(BLN110),.WL(WL91));
sram_cell_6t_5 inst_cell_91_111 (.BL(BL111),.BLN(BLN111),.WL(WL91));
sram_cell_6t_5 inst_cell_91_112 (.BL(BL112),.BLN(BLN112),.WL(WL91));
sram_cell_6t_5 inst_cell_91_113 (.BL(BL113),.BLN(BLN113),.WL(WL91));
sram_cell_6t_5 inst_cell_91_114 (.BL(BL114),.BLN(BLN114),.WL(WL91));
sram_cell_6t_5 inst_cell_91_115 (.BL(BL115),.BLN(BLN115),.WL(WL91));
sram_cell_6t_5 inst_cell_91_116 (.BL(BL116),.BLN(BLN116),.WL(WL91));
sram_cell_6t_5 inst_cell_91_117 (.BL(BL117),.BLN(BLN117),.WL(WL91));
sram_cell_6t_5 inst_cell_91_118 (.BL(BL118),.BLN(BLN118),.WL(WL91));
sram_cell_6t_5 inst_cell_91_119 (.BL(BL119),.BLN(BLN119),.WL(WL91));
sram_cell_6t_5 inst_cell_91_120 (.BL(BL120),.BLN(BLN120),.WL(WL91));
sram_cell_6t_5 inst_cell_91_121 (.BL(BL121),.BLN(BLN121),.WL(WL91));
sram_cell_6t_5 inst_cell_91_122 (.BL(BL122),.BLN(BLN122),.WL(WL91));
sram_cell_6t_5 inst_cell_91_123 (.BL(BL123),.BLN(BLN123),.WL(WL91));
sram_cell_6t_5 inst_cell_91_124 (.BL(BL124),.BLN(BLN124),.WL(WL91));
sram_cell_6t_5 inst_cell_91_125 (.BL(BL125),.BLN(BLN125),.WL(WL91));
sram_cell_6t_5 inst_cell_91_126 (.BL(BL126),.BLN(BLN126),.WL(WL91));
sram_cell_6t_5 inst_cell_91_127 (.BL(BL127),.BLN(BLN127),.WL(WL91));
sram_cell_6t_5 inst_cell_92_0 (.BL(BL0),.BLN(BLN0),.WL(WL92));
sram_cell_6t_5 inst_cell_92_1 (.BL(BL1),.BLN(BLN1),.WL(WL92));
sram_cell_6t_5 inst_cell_92_2 (.BL(BL2),.BLN(BLN2),.WL(WL92));
sram_cell_6t_5 inst_cell_92_3 (.BL(BL3),.BLN(BLN3),.WL(WL92));
sram_cell_6t_5 inst_cell_92_4 (.BL(BL4),.BLN(BLN4),.WL(WL92));
sram_cell_6t_5 inst_cell_92_5 (.BL(BL5),.BLN(BLN5),.WL(WL92));
sram_cell_6t_5 inst_cell_92_6 (.BL(BL6),.BLN(BLN6),.WL(WL92));
sram_cell_6t_5 inst_cell_92_7 (.BL(BL7),.BLN(BLN7),.WL(WL92));
sram_cell_6t_5 inst_cell_92_8 (.BL(BL8),.BLN(BLN8),.WL(WL92));
sram_cell_6t_5 inst_cell_92_9 (.BL(BL9),.BLN(BLN9),.WL(WL92));
sram_cell_6t_5 inst_cell_92_10 (.BL(BL10),.BLN(BLN10),.WL(WL92));
sram_cell_6t_5 inst_cell_92_11 (.BL(BL11),.BLN(BLN11),.WL(WL92));
sram_cell_6t_5 inst_cell_92_12 (.BL(BL12),.BLN(BLN12),.WL(WL92));
sram_cell_6t_5 inst_cell_92_13 (.BL(BL13),.BLN(BLN13),.WL(WL92));
sram_cell_6t_5 inst_cell_92_14 (.BL(BL14),.BLN(BLN14),.WL(WL92));
sram_cell_6t_5 inst_cell_92_15 (.BL(BL15),.BLN(BLN15),.WL(WL92));
sram_cell_6t_5 inst_cell_92_16 (.BL(BL16),.BLN(BLN16),.WL(WL92));
sram_cell_6t_5 inst_cell_92_17 (.BL(BL17),.BLN(BLN17),.WL(WL92));
sram_cell_6t_5 inst_cell_92_18 (.BL(BL18),.BLN(BLN18),.WL(WL92));
sram_cell_6t_5 inst_cell_92_19 (.BL(BL19),.BLN(BLN19),.WL(WL92));
sram_cell_6t_5 inst_cell_92_20 (.BL(BL20),.BLN(BLN20),.WL(WL92));
sram_cell_6t_5 inst_cell_92_21 (.BL(BL21),.BLN(BLN21),.WL(WL92));
sram_cell_6t_5 inst_cell_92_22 (.BL(BL22),.BLN(BLN22),.WL(WL92));
sram_cell_6t_5 inst_cell_92_23 (.BL(BL23),.BLN(BLN23),.WL(WL92));
sram_cell_6t_5 inst_cell_92_24 (.BL(BL24),.BLN(BLN24),.WL(WL92));
sram_cell_6t_5 inst_cell_92_25 (.BL(BL25),.BLN(BLN25),.WL(WL92));
sram_cell_6t_5 inst_cell_92_26 (.BL(BL26),.BLN(BLN26),.WL(WL92));
sram_cell_6t_5 inst_cell_92_27 (.BL(BL27),.BLN(BLN27),.WL(WL92));
sram_cell_6t_5 inst_cell_92_28 (.BL(BL28),.BLN(BLN28),.WL(WL92));
sram_cell_6t_5 inst_cell_92_29 (.BL(BL29),.BLN(BLN29),.WL(WL92));
sram_cell_6t_5 inst_cell_92_30 (.BL(BL30),.BLN(BLN30),.WL(WL92));
sram_cell_6t_5 inst_cell_92_31 (.BL(BL31),.BLN(BLN31),.WL(WL92));
sram_cell_6t_5 inst_cell_92_32 (.BL(BL32),.BLN(BLN32),.WL(WL92));
sram_cell_6t_5 inst_cell_92_33 (.BL(BL33),.BLN(BLN33),.WL(WL92));
sram_cell_6t_5 inst_cell_92_34 (.BL(BL34),.BLN(BLN34),.WL(WL92));
sram_cell_6t_5 inst_cell_92_35 (.BL(BL35),.BLN(BLN35),.WL(WL92));
sram_cell_6t_5 inst_cell_92_36 (.BL(BL36),.BLN(BLN36),.WL(WL92));
sram_cell_6t_5 inst_cell_92_37 (.BL(BL37),.BLN(BLN37),.WL(WL92));
sram_cell_6t_5 inst_cell_92_38 (.BL(BL38),.BLN(BLN38),.WL(WL92));
sram_cell_6t_5 inst_cell_92_39 (.BL(BL39),.BLN(BLN39),.WL(WL92));
sram_cell_6t_5 inst_cell_92_40 (.BL(BL40),.BLN(BLN40),.WL(WL92));
sram_cell_6t_5 inst_cell_92_41 (.BL(BL41),.BLN(BLN41),.WL(WL92));
sram_cell_6t_5 inst_cell_92_42 (.BL(BL42),.BLN(BLN42),.WL(WL92));
sram_cell_6t_5 inst_cell_92_43 (.BL(BL43),.BLN(BLN43),.WL(WL92));
sram_cell_6t_5 inst_cell_92_44 (.BL(BL44),.BLN(BLN44),.WL(WL92));
sram_cell_6t_5 inst_cell_92_45 (.BL(BL45),.BLN(BLN45),.WL(WL92));
sram_cell_6t_5 inst_cell_92_46 (.BL(BL46),.BLN(BLN46),.WL(WL92));
sram_cell_6t_5 inst_cell_92_47 (.BL(BL47),.BLN(BLN47),.WL(WL92));
sram_cell_6t_5 inst_cell_92_48 (.BL(BL48),.BLN(BLN48),.WL(WL92));
sram_cell_6t_5 inst_cell_92_49 (.BL(BL49),.BLN(BLN49),.WL(WL92));
sram_cell_6t_5 inst_cell_92_50 (.BL(BL50),.BLN(BLN50),.WL(WL92));
sram_cell_6t_5 inst_cell_92_51 (.BL(BL51),.BLN(BLN51),.WL(WL92));
sram_cell_6t_5 inst_cell_92_52 (.BL(BL52),.BLN(BLN52),.WL(WL92));
sram_cell_6t_5 inst_cell_92_53 (.BL(BL53),.BLN(BLN53),.WL(WL92));
sram_cell_6t_5 inst_cell_92_54 (.BL(BL54),.BLN(BLN54),.WL(WL92));
sram_cell_6t_5 inst_cell_92_55 (.BL(BL55),.BLN(BLN55),.WL(WL92));
sram_cell_6t_5 inst_cell_92_56 (.BL(BL56),.BLN(BLN56),.WL(WL92));
sram_cell_6t_5 inst_cell_92_57 (.BL(BL57),.BLN(BLN57),.WL(WL92));
sram_cell_6t_5 inst_cell_92_58 (.BL(BL58),.BLN(BLN58),.WL(WL92));
sram_cell_6t_5 inst_cell_92_59 (.BL(BL59),.BLN(BLN59),.WL(WL92));
sram_cell_6t_5 inst_cell_92_60 (.BL(BL60),.BLN(BLN60),.WL(WL92));
sram_cell_6t_5 inst_cell_92_61 (.BL(BL61),.BLN(BLN61),.WL(WL92));
sram_cell_6t_5 inst_cell_92_62 (.BL(BL62),.BLN(BLN62),.WL(WL92));
sram_cell_6t_5 inst_cell_92_63 (.BL(BL63),.BLN(BLN63),.WL(WL92));
sram_cell_6t_5 inst_cell_92_64 (.BL(BL64),.BLN(BLN64),.WL(WL92));
sram_cell_6t_5 inst_cell_92_65 (.BL(BL65),.BLN(BLN65),.WL(WL92));
sram_cell_6t_5 inst_cell_92_66 (.BL(BL66),.BLN(BLN66),.WL(WL92));
sram_cell_6t_5 inst_cell_92_67 (.BL(BL67),.BLN(BLN67),.WL(WL92));
sram_cell_6t_5 inst_cell_92_68 (.BL(BL68),.BLN(BLN68),.WL(WL92));
sram_cell_6t_5 inst_cell_92_69 (.BL(BL69),.BLN(BLN69),.WL(WL92));
sram_cell_6t_5 inst_cell_92_70 (.BL(BL70),.BLN(BLN70),.WL(WL92));
sram_cell_6t_5 inst_cell_92_71 (.BL(BL71),.BLN(BLN71),.WL(WL92));
sram_cell_6t_5 inst_cell_92_72 (.BL(BL72),.BLN(BLN72),.WL(WL92));
sram_cell_6t_5 inst_cell_92_73 (.BL(BL73),.BLN(BLN73),.WL(WL92));
sram_cell_6t_5 inst_cell_92_74 (.BL(BL74),.BLN(BLN74),.WL(WL92));
sram_cell_6t_5 inst_cell_92_75 (.BL(BL75),.BLN(BLN75),.WL(WL92));
sram_cell_6t_5 inst_cell_92_76 (.BL(BL76),.BLN(BLN76),.WL(WL92));
sram_cell_6t_5 inst_cell_92_77 (.BL(BL77),.BLN(BLN77),.WL(WL92));
sram_cell_6t_5 inst_cell_92_78 (.BL(BL78),.BLN(BLN78),.WL(WL92));
sram_cell_6t_5 inst_cell_92_79 (.BL(BL79),.BLN(BLN79),.WL(WL92));
sram_cell_6t_5 inst_cell_92_80 (.BL(BL80),.BLN(BLN80),.WL(WL92));
sram_cell_6t_5 inst_cell_92_81 (.BL(BL81),.BLN(BLN81),.WL(WL92));
sram_cell_6t_5 inst_cell_92_82 (.BL(BL82),.BLN(BLN82),.WL(WL92));
sram_cell_6t_5 inst_cell_92_83 (.BL(BL83),.BLN(BLN83),.WL(WL92));
sram_cell_6t_5 inst_cell_92_84 (.BL(BL84),.BLN(BLN84),.WL(WL92));
sram_cell_6t_5 inst_cell_92_85 (.BL(BL85),.BLN(BLN85),.WL(WL92));
sram_cell_6t_5 inst_cell_92_86 (.BL(BL86),.BLN(BLN86),.WL(WL92));
sram_cell_6t_5 inst_cell_92_87 (.BL(BL87),.BLN(BLN87),.WL(WL92));
sram_cell_6t_5 inst_cell_92_88 (.BL(BL88),.BLN(BLN88),.WL(WL92));
sram_cell_6t_5 inst_cell_92_89 (.BL(BL89),.BLN(BLN89),.WL(WL92));
sram_cell_6t_5 inst_cell_92_90 (.BL(BL90),.BLN(BLN90),.WL(WL92));
sram_cell_6t_5 inst_cell_92_91 (.BL(BL91),.BLN(BLN91),.WL(WL92));
sram_cell_6t_5 inst_cell_92_92 (.BL(BL92),.BLN(BLN92),.WL(WL92));
sram_cell_6t_5 inst_cell_92_93 (.BL(BL93),.BLN(BLN93),.WL(WL92));
sram_cell_6t_5 inst_cell_92_94 (.BL(BL94),.BLN(BLN94),.WL(WL92));
sram_cell_6t_5 inst_cell_92_95 (.BL(BL95),.BLN(BLN95),.WL(WL92));
sram_cell_6t_5 inst_cell_92_96 (.BL(BL96),.BLN(BLN96),.WL(WL92));
sram_cell_6t_5 inst_cell_92_97 (.BL(BL97),.BLN(BLN97),.WL(WL92));
sram_cell_6t_5 inst_cell_92_98 (.BL(BL98),.BLN(BLN98),.WL(WL92));
sram_cell_6t_5 inst_cell_92_99 (.BL(BL99),.BLN(BLN99),.WL(WL92));
sram_cell_6t_5 inst_cell_92_100 (.BL(BL100),.BLN(BLN100),.WL(WL92));
sram_cell_6t_5 inst_cell_92_101 (.BL(BL101),.BLN(BLN101),.WL(WL92));
sram_cell_6t_5 inst_cell_92_102 (.BL(BL102),.BLN(BLN102),.WL(WL92));
sram_cell_6t_5 inst_cell_92_103 (.BL(BL103),.BLN(BLN103),.WL(WL92));
sram_cell_6t_5 inst_cell_92_104 (.BL(BL104),.BLN(BLN104),.WL(WL92));
sram_cell_6t_5 inst_cell_92_105 (.BL(BL105),.BLN(BLN105),.WL(WL92));
sram_cell_6t_5 inst_cell_92_106 (.BL(BL106),.BLN(BLN106),.WL(WL92));
sram_cell_6t_5 inst_cell_92_107 (.BL(BL107),.BLN(BLN107),.WL(WL92));
sram_cell_6t_5 inst_cell_92_108 (.BL(BL108),.BLN(BLN108),.WL(WL92));
sram_cell_6t_5 inst_cell_92_109 (.BL(BL109),.BLN(BLN109),.WL(WL92));
sram_cell_6t_5 inst_cell_92_110 (.BL(BL110),.BLN(BLN110),.WL(WL92));
sram_cell_6t_5 inst_cell_92_111 (.BL(BL111),.BLN(BLN111),.WL(WL92));
sram_cell_6t_5 inst_cell_92_112 (.BL(BL112),.BLN(BLN112),.WL(WL92));
sram_cell_6t_5 inst_cell_92_113 (.BL(BL113),.BLN(BLN113),.WL(WL92));
sram_cell_6t_5 inst_cell_92_114 (.BL(BL114),.BLN(BLN114),.WL(WL92));
sram_cell_6t_5 inst_cell_92_115 (.BL(BL115),.BLN(BLN115),.WL(WL92));
sram_cell_6t_5 inst_cell_92_116 (.BL(BL116),.BLN(BLN116),.WL(WL92));
sram_cell_6t_5 inst_cell_92_117 (.BL(BL117),.BLN(BLN117),.WL(WL92));
sram_cell_6t_5 inst_cell_92_118 (.BL(BL118),.BLN(BLN118),.WL(WL92));
sram_cell_6t_5 inst_cell_92_119 (.BL(BL119),.BLN(BLN119),.WL(WL92));
sram_cell_6t_5 inst_cell_92_120 (.BL(BL120),.BLN(BLN120),.WL(WL92));
sram_cell_6t_5 inst_cell_92_121 (.BL(BL121),.BLN(BLN121),.WL(WL92));
sram_cell_6t_5 inst_cell_92_122 (.BL(BL122),.BLN(BLN122),.WL(WL92));
sram_cell_6t_5 inst_cell_92_123 (.BL(BL123),.BLN(BLN123),.WL(WL92));
sram_cell_6t_5 inst_cell_92_124 (.BL(BL124),.BLN(BLN124),.WL(WL92));
sram_cell_6t_5 inst_cell_92_125 (.BL(BL125),.BLN(BLN125),.WL(WL92));
sram_cell_6t_5 inst_cell_92_126 (.BL(BL126),.BLN(BLN126),.WL(WL92));
sram_cell_6t_5 inst_cell_92_127 (.BL(BL127),.BLN(BLN127),.WL(WL92));
sram_cell_6t_5 inst_cell_93_0 (.BL(BL0),.BLN(BLN0),.WL(WL93));
sram_cell_6t_5 inst_cell_93_1 (.BL(BL1),.BLN(BLN1),.WL(WL93));
sram_cell_6t_5 inst_cell_93_2 (.BL(BL2),.BLN(BLN2),.WL(WL93));
sram_cell_6t_5 inst_cell_93_3 (.BL(BL3),.BLN(BLN3),.WL(WL93));
sram_cell_6t_5 inst_cell_93_4 (.BL(BL4),.BLN(BLN4),.WL(WL93));
sram_cell_6t_5 inst_cell_93_5 (.BL(BL5),.BLN(BLN5),.WL(WL93));
sram_cell_6t_5 inst_cell_93_6 (.BL(BL6),.BLN(BLN6),.WL(WL93));
sram_cell_6t_5 inst_cell_93_7 (.BL(BL7),.BLN(BLN7),.WL(WL93));
sram_cell_6t_5 inst_cell_93_8 (.BL(BL8),.BLN(BLN8),.WL(WL93));
sram_cell_6t_5 inst_cell_93_9 (.BL(BL9),.BLN(BLN9),.WL(WL93));
sram_cell_6t_5 inst_cell_93_10 (.BL(BL10),.BLN(BLN10),.WL(WL93));
sram_cell_6t_5 inst_cell_93_11 (.BL(BL11),.BLN(BLN11),.WL(WL93));
sram_cell_6t_5 inst_cell_93_12 (.BL(BL12),.BLN(BLN12),.WL(WL93));
sram_cell_6t_5 inst_cell_93_13 (.BL(BL13),.BLN(BLN13),.WL(WL93));
sram_cell_6t_5 inst_cell_93_14 (.BL(BL14),.BLN(BLN14),.WL(WL93));
sram_cell_6t_5 inst_cell_93_15 (.BL(BL15),.BLN(BLN15),.WL(WL93));
sram_cell_6t_5 inst_cell_93_16 (.BL(BL16),.BLN(BLN16),.WL(WL93));
sram_cell_6t_5 inst_cell_93_17 (.BL(BL17),.BLN(BLN17),.WL(WL93));
sram_cell_6t_5 inst_cell_93_18 (.BL(BL18),.BLN(BLN18),.WL(WL93));
sram_cell_6t_5 inst_cell_93_19 (.BL(BL19),.BLN(BLN19),.WL(WL93));
sram_cell_6t_5 inst_cell_93_20 (.BL(BL20),.BLN(BLN20),.WL(WL93));
sram_cell_6t_5 inst_cell_93_21 (.BL(BL21),.BLN(BLN21),.WL(WL93));
sram_cell_6t_5 inst_cell_93_22 (.BL(BL22),.BLN(BLN22),.WL(WL93));
sram_cell_6t_5 inst_cell_93_23 (.BL(BL23),.BLN(BLN23),.WL(WL93));
sram_cell_6t_5 inst_cell_93_24 (.BL(BL24),.BLN(BLN24),.WL(WL93));
sram_cell_6t_5 inst_cell_93_25 (.BL(BL25),.BLN(BLN25),.WL(WL93));
sram_cell_6t_5 inst_cell_93_26 (.BL(BL26),.BLN(BLN26),.WL(WL93));
sram_cell_6t_5 inst_cell_93_27 (.BL(BL27),.BLN(BLN27),.WL(WL93));
sram_cell_6t_5 inst_cell_93_28 (.BL(BL28),.BLN(BLN28),.WL(WL93));
sram_cell_6t_5 inst_cell_93_29 (.BL(BL29),.BLN(BLN29),.WL(WL93));
sram_cell_6t_5 inst_cell_93_30 (.BL(BL30),.BLN(BLN30),.WL(WL93));
sram_cell_6t_5 inst_cell_93_31 (.BL(BL31),.BLN(BLN31),.WL(WL93));
sram_cell_6t_5 inst_cell_93_32 (.BL(BL32),.BLN(BLN32),.WL(WL93));
sram_cell_6t_5 inst_cell_93_33 (.BL(BL33),.BLN(BLN33),.WL(WL93));
sram_cell_6t_5 inst_cell_93_34 (.BL(BL34),.BLN(BLN34),.WL(WL93));
sram_cell_6t_5 inst_cell_93_35 (.BL(BL35),.BLN(BLN35),.WL(WL93));
sram_cell_6t_5 inst_cell_93_36 (.BL(BL36),.BLN(BLN36),.WL(WL93));
sram_cell_6t_5 inst_cell_93_37 (.BL(BL37),.BLN(BLN37),.WL(WL93));
sram_cell_6t_5 inst_cell_93_38 (.BL(BL38),.BLN(BLN38),.WL(WL93));
sram_cell_6t_5 inst_cell_93_39 (.BL(BL39),.BLN(BLN39),.WL(WL93));
sram_cell_6t_5 inst_cell_93_40 (.BL(BL40),.BLN(BLN40),.WL(WL93));
sram_cell_6t_5 inst_cell_93_41 (.BL(BL41),.BLN(BLN41),.WL(WL93));
sram_cell_6t_5 inst_cell_93_42 (.BL(BL42),.BLN(BLN42),.WL(WL93));
sram_cell_6t_5 inst_cell_93_43 (.BL(BL43),.BLN(BLN43),.WL(WL93));
sram_cell_6t_5 inst_cell_93_44 (.BL(BL44),.BLN(BLN44),.WL(WL93));
sram_cell_6t_5 inst_cell_93_45 (.BL(BL45),.BLN(BLN45),.WL(WL93));
sram_cell_6t_5 inst_cell_93_46 (.BL(BL46),.BLN(BLN46),.WL(WL93));
sram_cell_6t_5 inst_cell_93_47 (.BL(BL47),.BLN(BLN47),.WL(WL93));
sram_cell_6t_5 inst_cell_93_48 (.BL(BL48),.BLN(BLN48),.WL(WL93));
sram_cell_6t_5 inst_cell_93_49 (.BL(BL49),.BLN(BLN49),.WL(WL93));
sram_cell_6t_5 inst_cell_93_50 (.BL(BL50),.BLN(BLN50),.WL(WL93));
sram_cell_6t_5 inst_cell_93_51 (.BL(BL51),.BLN(BLN51),.WL(WL93));
sram_cell_6t_5 inst_cell_93_52 (.BL(BL52),.BLN(BLN52),.WL(WL93));
sram_cell_6t_5 inst_cell_93_53 (.BL(BL53),.BLN(BLN53),.WL(WL93));
sram_cell_6t_5 inst_cell_93_54 (.BL(BL54),.BLN(BLN54),.WL(WL93));
sram_cell_6t_5 inst_cell_93_55 (.BL(BL55),.BLN(BLN55),.WL(WL93));
sram_cell_6t_5 inst_cell_93_56 (.BL(BL56),.BLN(BLN56),.WL(WL93));
sram_cell_6t_5 inst_cell_93_57 (.BL(BL57),.BLN(BLN57),.WL(WL93));
sram_cell_6t_5 inst_cell_93_58 (.BL(BL58),.BLN(BLN58),.WL(WL93));
sram_cell_6t_5 inst_cell_93_59 (.BL(BL59),.BLN(BLN59),.WL(WL93));
sram_cell_6t_5 inst_cell_93_60 (.BL(BL60),.BLN(BLN60),.WL(WL93));
sram_cell_6t_5 inst_cell_93_61 (.BL(BL61),.BLN(BLN61),.WL(WL93));
sram_cell_6t_5 inst_cell_93_62 (.BL(BL62),.BLN(BLN62),.WL(WL93));
sram_cell_6t_5 inst_cell_93_63 (.BL(BL63),.BLN(BLN63),.WL(WL93));
sram_cell_6t_5 inst_cell_93_64 (.BL(BL64),.BLN(BLN64),.WL(WL93));
sram_cell_6t_5 inst_cell_93_65 (.BL(BL65),.BLN(BLN65),.WL(WL93));
sram_cell_6t_5 inst_cell_93_66 (.BL(BL66),.BLN(BLN66),.WL(WL93));
sram_cell_6t_5 inst_cell_93_67 (.BL(BL67),.BLN(BLN67),.WL(WL93));
sram_cell_6t_5 inst_cell_93_68 (.BL(BL68),.BLN(BLN68),.WL(WL93));
sram_cell_6t_5 inst_cell_93_69 (.BL(BL69),.BLN(BLN69),.WL(WL93));
sram_cell_6t_5 inst_cell_93_70 (.BL(BL70),.BLN(BLN70),.WL(WL93));
sram_cell_6t_5 inst_cell_93_71 (.BL(BL71),.BLN(BLN71),.WL(WL93));
sram_cell_6t_5 inst_cell_93_72 (.BL(BL72),.BLN(BLN72),.WL(WL93));
sram_cell_6t_5 inst_cell_93_73 (.BL(BL73),.BLN(BLN73),.WL(WL93));
sram_cell_6t_5 inst_cell_93_74 (.BL(BL74),.BLN(BLN74),.WL(WL93));
sram_cell_6t_5 inst_cell_93_75 (.BL(BL75),.BLN(BLN75),.WL(WL93));
sram_cell_6t_5 inst_cell_93_76 (.BL(BL76),.BLN(BLN76),.WL(WL93));
sram_cell_6t_5 inst_cell_93_77 (.BL(BL77),.BLN(BLN77),.WL(WL93));
sram_cell_6t_5 inst_cell_93_78 (.BL(BL78),.BLN(BLN78),.WL(WL93));
sram_cell_6t_5 inst_cell_93_79 (.BL(BL79),.BLN(BLN79),.WL(WL93));
sram_cell_6t_5 inst_cell_93_80 (.BL(BL80),.BLN(BLN80),.WL(WL93));
sram_cell_6t_5 inst_cell_93_81 (.BL(BL81),.BLN(BLN81),.WL(WL93));
sram_cell_6t_5 inst_cell_93_82 (.BL(BL82),.BLN(BLN82),.WL(WL93));
sram_cell_6t_5 inst_cell_93_83 (.BL(BL83),.BLN(BLN83),.WL(WL93));
sram_cell_6t_5 inst_cell_93_84 (.BL(BL84),.BLN(BLN84),.WL(WL93));
sram_cell_6t_5 inst_cell_93_85 (.BL(BL85),.BLN(BLN85),.WL(WL93));
sram_cell_6t_5 inst_cell_93_86 (.BL(BL86),.BLN(BLN86),.WL(WL93));
sram_cell_6t_5 inst_cell_93_87 (.BL(BL87),.BLN(BLN87),.WL(WL93));
sram_cell_6t_5 inst_cell_93_88 (.BL(BL88),.BLN(BLN88),.WL(WL93));
sram_cell_6t_5 inst_cell_93_89 (.BL(BL89),.BLN(BLN89),.WL(WL93));
sram_cell_6t_5 inst_cell_93_90 (.BL(BL90),.BLN(BLN90),.WL(WL93));
sram_cell_6t_5 inst_cell_93_91 (.BL(BL91),.BLN(BLN91),.WL(WL93));
sram_cell_6t_5 inst_cell_93_92 (.BL(BL92),.BLN(BLN92),.WL(WL93));
sram_cell_6t_5 inst_cell_93_93 (.BL(BL93),.BLN(BLN93),.WL(WL93));
sram_cell_6t_5 inst_cell_93_94 (.BL(BL94),.BLN(BLN94),.WL(WL93));
sram_cell_6t_5 inst_cell_93_95 (.BL(BL95),.BLN(BLN95),.WL(WL93));
sram_cell_6t_5 inst_cell_93_96 (.BL(BL96),.BLN(BLN96),.WL(WL93));
sram_cell_6t_5 inst_cell_93_97 (.BL(BL97),.BLN(BLN97),.WL(WL93));
sram_cell_6t_5 inst_cell_93_98 (.BL(BL98),.BLN(BLN98),.WL(WL93));
sram_cell_6t_5 inst_cell_93_99 (.BL(BL99),.BLN(BLN99),.WL(WL93));
sram_cell_6t_5 inst_cell_93_100 (.BL(BL100),.BLN(BLN100),.WL(WL93));
sram_cell_6t_5 inst_cell_93_101 (.BL(BL101),.BLN(BLN101),.WL(WL93));
sram_cell_6t_5 inst_cell_93_102 (.BL(BL102),.BLN(BLN102),.WL(WL93));
sram_cell_6t_5 inst_cell_93_103 (.BL(BL103),.BLN(BLN103),.WL(WL93));
sram_cell_6t_5 inst_cell_93_104 (.BL(BL104),.BLN(BLN104),.WL(WL93));
sram_cell_6t_5 inst_cell_93_105 (.BL(BL105),.BLN(BLN105),.WL(WL93));
sram_cell_6t_5 inst_cell_93_106 (.BL(BL106),.BLN(BLN106),.WL(WL93));
sram_cell_6t_5 inst_cell_93_107 (.BL(BL107),.BLN(BLN107),.WL(WL93));
sram_cell_6t_5 inst_cell_93_108 (.BL(BL108),.BLN(BLN108),.WL(WL93));
sram_cell_6t_5 inst_cell_93_109 (.BL(BL109),.BLN(BLN109),.WL(WL93));
sram_cell_6t_5 inst_cell_93_110 (.BL(BL110),.BLN(BLN110),.WL(WL93));
sram_cell_6t_5 inst_cell_93_111 (.BL(BL111),.BLN(BLN111),.WL(WL93));
sram_cell_6t_5 inst_cell_93_112 (.BL(BL112),.BLN(BLN112),.WL(WL93));
sram_cell_6t_5 inst_cell_93_113 (.BL(BL113),.BLN(BLN113),.WL(WL93));
sram_cell_6t_5 inst_cell_93_114 (.BL(BL114),.BLN(BLN114),.WL(WL93));
sram_cell_6t_5 inst_cell_93_115 (.BL(BL115),.BLN(BLN115),.WL(WL93));
sram_cell_6t_5 inst_cell_93_116 (.BL(BL116),.BLN(BLN116),.WL(WL93));
sram_cell_6t_5 inst_cell_93_117 (.BL(BL117),.BLN(BLN117),.WL(WL93));
sram_cell_6t_5 inst_cell_93_118 (.BL(BL118),.BLN(BLN118),.WL(WL93));
sram_cell_6t_5 inst_cell_93_119 (.BL(BL119),.BLN(BLN119),.WL(WL93));
sram_cell_6t_5 inst_cell_93_120 (.BL(BL120),.BLN(BLN120),.WL(WL93));
sram_cell_6t_5 inst_cell_93_121 (.BL(BL121),.BLN(BLN121),.WL(WL93));
sram_cell_6t_5 inst_cell_93_122 (.BL(BL122),.BLN(BLN122),.WL(WL93));
sram_cell_6t_5 inst_cell_93_123 (.BL(BL123),.BLN(BLN123),.WL(WL93));
sram_cell_6t_5 inst_cell_93_124 (.BL(BL124),.BLN(BLN124),.WL(WL93));
sram_cell_6t_5 inst_cell_93_125 (.BL(BL125),.BLN(BLN125),.WL(WL93));
sram_cell_6t_5 inst_cell_93_126 (.BL(BL126),.BLN(BLN126),.WL(WL93));
sram_cell_6t_5 inst_cell_93_127 (.BL(BL127),.BLN(BLN127),.WL(WL93));
sram_cell_6t_5 inst_cell_94_0 (.BL(BL0),.BLN(BLN0),.WL(WL94));
sram_cell_6t_5 inst_cell_94_1 (.BL(BL1),.BLN(BLN1),.WL(WL94));
sram_cell_6t_5 inst_cell_94_2 (.BL(BL2),.BLN(BLN2),.WL(WL94));
sram_cell_6t_5 inst_cell_94_3 (.BL(BL3),.BLN(BLN3),.WL(WL94));
sram_cell_6t_5 inst_cell_94_4 (.BL(BL4),.BLN(BLN4),.WL(WL94));
sram_cell_6t_5 inst_cell_94_5 (.BL(BL5),.BLN(BLN5),.WL(WL94));
sram_cell_6t_5 inst_cell_94_6 (.BL(BL6),.BLN(BLN6),.WL(WL94));
sram_cell_6t_5 inst_cell_94_7 (.BL(BL7),.BLN(BLN7),.WL(WL94));
sram_cell_6t_5 inst_cell_94_8 (.BL(BL8),.BLN(BLN8),.WL(WL94));
sram_cell_6t_5 inst_cell_94_9 (.BL(BL9),.BLN(BLN9),.WL(WL94));
sram_cell_6t_5 inst_cell_94_10 (.BL(BL10),.BLN(BLN10),.WL(WL94));
sram_cell_6t_5 inst_cell_94_11 (.BL(BL11),.BLN(BLN11),.WL(WL94));
sram_cell_6t_5 inst_cell_94_12 (.BL(BL12),.BLN(BLN12),.WL(WL94));
sram_cell_6t_5 inst_cell_94_13 (.BL(BL13),.BLN(BLN13),.WL(WL94));
sram_cell_6t_5 inst_cell_94_14 (.BL(BL14),.BLN(BLN14),.WL(WL94));
sram_cell_6t_5 inst_cell_94_15 (.BL(BL15),.BLN(BLN15),.WL(WL94));
sram_cell_6t_5 inst_cell_94_16 (.BL(BL16),.BLN(BLN16),.WL(WL94));
sram_cell_6t_5 inst_cell_94_17 (.BL(BL17),.BLN(BLN17),.WL(WL94));
sram_cell_6t_5 inst_cell_94_18 (.BL(BL18),.BLN(BLN18),.WL(WL94));
sram_cell_6t_5 inst_cell_94_19 (.BL(BL19),.BLN(BLN19),.WL(WL94));
sram_cell_6t_5 inst_cell_94_20 (.BL(BL20),.BLN(BLN20),.WL(WL94));
sram_cell_6t_5 inst_cell_94_21 (.BL(BL21),.BLN(BLN21),.WL(WL94));
sram_cell_6t_5 inst_cell_94_22 (.BL(BL22),.BLN(BLN22),.WL(WL94));
sram_cell_6t_5 inst_cell_94_23 (.BL(BL23),.BLN(BLN23),.WL(WL94));
sram_cell_6t_5 inst_cell_94_24 (.BL(BL24),.BLN(BLN24),.WL(WL94));
sram_cell_6t_5 inst_cell_94_25 (.BL(BL25),.BLN(BLN25),.WL(WL94));
sram_cell_6t_5 inst_cell_94_26 (.BL(BL26),.BLN(BLN26),.WL(WL94));
sram_cell_6t_5 inst_cell_94_27 (.BL(BL27),.BLN(BLN27),.WL(WL94));
sram_cell_6t_5 inst_cell_94_28 (.BL(BL28),.BLN(BLN28),.WL(WL94));
sram_cell_6t_5 inst_cell_94_29 (.BL(BL29),.BLN(BLN29),.WL(WL94));
sram_cell_6t_5 inst_cell_94_30 (.BL(BL30),.BLN(BLN30),.WL(WL94));
sram_cell_6t_5 inst_cell_94_31 (.BL(BL31),.BLN(BLN31),.WL(WL94));
sram_cell_6t_5 inst_cell_94_32 (.BL(BL32),.BLN(BLN32),.WL(WL94));
sram_cell_6t_5 inst_cell_94_33 (.BL(BL33),.BLN(BLN33),.WL(WL94));
sram_cell_6t_5 inst_cell_94_34 (.BL(BL34),.BLN(BLN34),.WL(WL94));
sram_cell_6t_5 inst_cell_94_35 (.BL(BL35),.BLN(BLN35),.WL(WL94));
sram_cell_6t_5 inst_cell_94_36 (.BL(BL36),.BLN(BLN36),.WL(WL94));
sram_cell_6t_5 inst_cell_94_37 (.BL(BL37),.BLN(BLN37),.WL(WL94));
sram_cell_6t_5 inst_cell_94_38 (.BL(BL38),.BLN(BLN38),.WL(WL94));
sram_cell_6t_5 inst_cell_94_39 (.BL(BL39),.BLN(BLN39),.WL(WL94));
sram_cell_6t_5 inst_cell_94_40 (.BL(BL40),.BLN(BLN40),.WL(WL94));
sram_cell_6t_5 inst_cell_94_41 (.BL(BL41),.BLN(BLN41),.WL(WL94));
sram_cell_6t_5 inst_cell_94_42 (.BL(BL42),.BLN(BLN42),.WL(WL94));
sram_cell_6t_5 inst_cell_94_43 (.BL(BL43),.BLN(BLN43),.WL(WL94));
sram_cell_6t_5 inst_cell_94_44 (.BL(BL44),.BLN(BLN44),.WL(WL94));
sram_cell_6t_5 inst_cell_94_45 (.BL(BL45),.BLN(BLN45),.WL(WL94));
sram_cell_6t_5 inst_cell_94_46 (.BL(BL46),.BLN(BLN46),.WL(WL94));
sram_cell_6t_5 inst_cell_94_47 (.BL(BL47),.BLN(BLN47),.WL(WL94));
sram_cell_6t_5 inst_cell_94_48 (.BL(BL48),.BLN(BLN48),.WL(WL94));
sram_cell_6t_5 inst_cell_94_49 (.BL(BL49),.BLN(BLN49),.WL(WL94));
sram_cell_6t_5 inst_cell_94_50 (.BL(BL50),.BLN(BLN50),.WL(WL94));
sram_cell_6t_5 inst_cell_94_51 (.BL(BL51),.BLN(BLN51),.WL(WL94));
sram_cell_6t_5 inst_cell_94_52 (.BL(BL52),.BLN(BLN52),.WL(WL94));
sram_cell_6t_5 inst_cell_94_53 (.BL(BL53),.BLN(BLN53),.WL(WL94));
sram_cell_6t_5 inst_cell_94_54 (.BL(BL54),.BLN(BLN54),.WL(WL94));
sram_cell_6t_5 inst_cell_94_55 (.BL(BL55),.BLN(BLN55),.WL(WL94));
sram_cell_6t_5 inst_cell_94_56 (.BL(BL56),.BLN(BLN56),.WL(WL94));
sram_cell_6t_5 inst_cell_94_57 (.BL(BL57),.BLN(BLN57),.WL(WL94));
sram_cell_6t_5 inst_cell_94_58 (.BL(BL58),.BLN(BLN58),.WL(WL94));
sram_cell_6t_5 inst_cell_94_59 (.BL(BL59),.BLN(BLN59),.WL(WL94));
sram_cell_6t_5 inst_cell_94_60 (.BL(BL60),.BLN(BLN60),.WL(WL94));
sram_cell_6t_5 inst_cell_94_61 (.BL(BL61),.BLN(BLN61),.WL(WL94));
sram_cell_6t_5 inst_cell_94_62 (.BL(BL62),.BLN(BLN62),.WL(WL94));
sram_cell_6t_5 inst_cell_94_63 (.BL(BL63),.BLN(BLN63),.WL(WL94));
sram_cell_6t_5 inst_cell_94_64 (.BL(BL64),.BLN(BLN64),.WL(WL94));
sram_cell_6t_5 inst_cell_94_65 (.BL(BL65),.BLN(BLN65),.WL(WL94));
sram_cell_6t_5 inst_cell_94_66 (.BL(BL66),.BLN(BLN66),.WL(WL94));
sram_cell_6t_5 inst_cell_94_67 (.BL(BL67),.BLN(BLN67),.WL(WL94));
sram_cell_6t_5 inst_cell_94_68 (.BL(BL68),.BLN(BLN68),.WL(WL94));
sram_cell_6t_5 inst_cell_94_69 (.BL(BL69),.BLN(BLN69),.WL(WL94));
sram_cell_6t_5 inst_cell_94_70 (.BL(BL70),.BLN(BLN70),.WL(WL94));
sram_cell_6t_5 inst_cell_94_71 (.BL(BL71),.BLN(BLN71),.WL(WL94));
sram_cell_6t_5 inst_cell_94_72 (.BL(BL72),.BLN(BLN72),.WL(WL94));
sram_cell_6t_5 inst_cell_94_73 (.BL(BL73),.BLN(BLN73),.WL(WL94));
sram_cell_6t_5 inst_cell_94_74 (.BL(BL74),.BLN(BLN74),.WL(WL94));
sram_cell_6t_5 inst_cell_94_75 (.BL(BL75),.BLN(BLN75),.WL(WL94));
sram_cell_6t_5 inst_cell_94_76 (.BL(BL76),.BLN(BLN76),.WL(WL94));
sram_cell_6t_5 inst_cell_94_77 (.BL(BL77),.BLN(BLN77),.WL(WL94));
sram_cell_6t_5 inst_cell_94_78 (.BL(BL78),.BLN(BLN78),.WL(WL94));
sram_cell_6t_5 inst_cell_94_79 (.BL(BL79),.BLN(BLN79),.WL(WL94));
sram_cell_6t_5 inst_cell_94_80 (.BL(BL80),.BLN(BLN80),.WL(WL94));
sram_cell_6t_5 inst_cell_94_81 (.BL(BL81),.BLN(BLN81),.WL(WL94));
sram_cell_6t_5 inst_cell_94_82 (.BL(BL82),.BLN(BLN82),.WL(WL94));
sram_cell_6t_5 inst_cell_94_83 (.BL(BL83),.BLN(BLN83),.WL(WL94));
sram_cell_6t_5 inst_cell_94_84 (.BL(BL84),.BLN(BLN84),.WL(WL94));
sram_cell_6t_5 inst_cell_94_85 (.BL(BL85),.BLN(BLN85),.WL(WL94));
sram_cell_6t_5 inst_cell_94_86 (.BL(BL86),.BLN(BLN86),.WL(WL94));
sram_cell_6t_5 inst_cell_94_87 (.BL(BL87),.BLN(BLN87),.WL(WL94));
sram_cell_6t_5 inst_cell_94_88 (.BL(BL88),.BLN(BLN88),.WL(WL94));
sram_cell_6t_5 inst_cell_94_89 (.BL(BL89),.BLN(BLN89),.WL(WL94));
sram_cell_6t_5 inst_cell_94_90 (.BL(BL90),.BLN(BLN90),.WL(WL94));
sram_cell_6t_5 inst_cell_94_91 (.BL(BL91),.BLN(BLN91),.WL(WL94));
sram_cell_6t_5 inst_cell_94_92 (.BL(BL92),.BLN(BLN92),.WL(WL94));
sram_cell_6t_5 inst_cell_94_93 (.BL(BL93),.BLN(BLN93),.WL(WL94));
sram_cell_6t_5 inst_cell_94_94 (.BL(BL94),.BLN(BLN94),.WL(WL94));
sram_cell_6t_5 inst_cell_94_95 (.BL(BL95),.BLN(BLN95),.WL(WL94));
sram_cell_6t_5 inst_cell_94_96 (.BL(BL96),.BLN(BLN96),.WL(WL94));
sram_cell_6t_5 inst_cell_94_97 (.BL(BL97),.BLN(BLN97),.WL(WL94));
sram_cell_6t_5 inst_cell_94_98 (.BL(BL98),.BLN(BLN98),.WL(WL94));
sram_cell_6t_5 inst_cell_94_99 (.BL(BL99),.BLN(BLN99),.WL(WL94));
sram_cell_6t_5 inst_cell_94_100 (.BL(BL100),.BLN(BLN100),.WL(WL94));
sram_cell_6t_5 inst_cell_94_101 (.BL(BL101),.BLN(BLN101),.WL(WL94));
sram_cell_6t_5 inst_cell_94_102 (.BL(BL102),.BLN(BLN102),.WL(WL94));
sram_cell_6t_5 inst_cell_94_103 (.BL(BL103),.BLN(BLN103),.WL(WL94));
sram_cell_6t_5 inst_cell_94_104 (.BL(BL104),.BLN(BLN104),.WL(WL94));
sram_cell_6t_5 inst_cell_94_105 (.BL(BL105),.BLN(BLN105),.WL(WL94));
sram_cell_6t_5 inst_cell_94_106 (.BL(BL106),.BLN(BLN106),.WL(WL94));
sram_cell_6t_5 inst_cell_94_107 (.BL(BL107),.BLN(BLN107),.WL(WL94));
sram_cell_6t_5 inst_cell_94_108 (.BL(BL108),.BLN(BLN108),.WL(WL94));
sram_cell_6t_5 inst_cell_94_109 (.BL(BL109),.BLN(BLN109),.WL(WL94));
sram_cell_6t_5 inst_cell_94_110 (.BL(BL110),.BLN(BLN110),.WL(WL94));
sram_cell_6t_5 inst_cell_94_111 (.BL(BL111),.BLN(BLN111),.WL(WL94));
sram_cell_6t_5 inst_cell_94_112 (.BL(BL112),.BLN(BLN112),.WL(WL94));
sram_cell_6t_5 inst_cell_94_113 (.BL(BL113),.BLN(BLN113),.WL(WL94));
sram_cell_6t_5 inst_cell_94_114 (.BL(BL114),.BLN(BLN114),.WL(WL94));
sram_cell_6t_5 inst_cell_94_115 (.BL(BL115),.BLN(BLN115),.WL(WL94));
sram_cell_6t_5 inst_cell_94_116 (.BL(BL116),.BLN(BLN116),.WL(WL94));
sram_cell_6t_5 inst_cell_94_117 (.BL(BL117),.BLN(BLN117),.WL(WL94));
sram_cell_6t_5 inst_cell_94_118 (.BL(BL118),.BLN(BLN118),.WL(WL94));
sram_cell_6t_5 inst_cell_94_119 (.BL(BL119),.BLN(BLN119),.WL(WL94));
sram_cell_6t_5 inst_cell_94_120 (.BL(BL120),.BLN(BLN120),.WL(WL94));
sram_cell_6t_5 inst_cell_94_121 (.BL(BL121),.BLN(BLN121),.WL(WL94));
sram_cell_6t_5 inst_cell_94_122 (.BL(BL122),.BLN(BLN122),.WL(WL94));
sram_cell_6t_5 inst_cell_94_123 (.BL(BL123),.BLN(BLN123),.WL(WL94));
sram_cell_6t_5 inst_cell_94_124 (.BL(BL124),.BLN(BLN124),.WL(WL94));
sram_cell_6t_5 inst_cell_94_125 (.BL(BL125),.BLN(BLN125),.WL(WL94));
sram_cell_6t_5 inst_cell_94_126 (.BL(BL126),.BLN(BLN126),.WL(WL94));
sram_cell_6t_5 inst_cell_94_127 (.BL(BL127),.BLN(BLN127),.WL(WL94));
sram_cell_6t_5 inst_cell_95_0 (.BL(BL0),.BLN(BLN0),.WL(WL95));
sram_cell_6t_5 inst_cell_95_1 (.BL(BL1),.BLN(BLN1),.WL(WL95));
sram_cell_6t_5 inst_cell_95_2 (.BL(BL2),.BLN(BLN2),.WL(WL95));
sram_cell_6t_5 inst_cell_95_3 (.BL(BL3),.BLN(BLN3),.WL(WL95));
sram_cell_6t_5 inst_cell_95_4 (.BL(BL4),.BLN(BLN4),.WL(WL95));
sram_cell_6t_5 inst_cell_95_5 (.BL(BL5),.BLN(BLN5),.WL(WL95));
sram_cell_6t_5 inst_cell_95_6 (.BL(BL6),.BLN(BLN6),.WL(WL95));
sram_cell_6t_5 inst_cell_95_7 (.BL(BL7),.BLN(BLN7),.WL(WL95));
sram_cell_6t_5 inst_cell_95_8 (.BL(BL8),.BLN(BLN8),.WL(WL95));
sram_cell_6t_5 inst_cell_95_9 (.BL(BL9),.BLN(BLN9),.WL(WL95));
sram_cell_6t_5 inst_cell_95_10 (.BL(BL10),.BLN(BLN10),.WL(WL95));
sram_cell_6t_5 inst_cell_95_11 (.BL(BL11),.BLN(BLN11),.WL(WL95));
sram_cell_6t_5 inst_cell_95_12 (.BL(BL12),.BLN(BLN12),.WL(WL95));
sram_cell_6t_5 inst_cell_95_13 (.BL(BL13),.BLN(BLN13),.WL(WL95));
sram_cell_6t_5 inst_cell_95_14 (.BL(BL14),.BLN(BLN14),.WL(WL95));
sram_cell_6t_5 inst_cell_95_15 (.BL(BL15),.BLN(BLN15),.WL(WL95));
sram_cell_6t_5 inst_cell_95_16 (.BL(BL16),.BLN(BLN16),.WL(WL95));
sram_cell_6t_5 inst_cell_95_17 (.BL(BL17),.BLN(BLN17),.WL(WL95));
sram_cell_6t_5 inst_cell_95_18 (.BL(BL18),.BLN(BLN18),.WL(WL95));
sram_cell_6t_5 inst_cell_95_19 (.BL(BL19),.BLN(BLN19),.WL(WL95));
sram_cell_6t_5 inst_cell_95_20 (.BL(BL20),.BLN(BLN20),.WL(WL95));
sram_cell_6t_5 inst_cell_95_21 (.BL(BL21),.BLN(BLN21),.WL(WL95));
sram_cell_6t_5 inst_cell_95_22 (.BL(BL22),.BLN(BLN22),.WL(WL95));
sram_cell_6t_5 inst_cell_95_23 (.BL(BL23),.BLN(BLN23),.WL(WL95));
sram_cell_6t_5 inst_cell_95_24 (.BL(BL24),.BLN(BLN24),.WL(WL95));
sram_cell_6t_5 inst_cell_95_25 (.BL(BL25),.BLN(BLN25),.WL(WL95));
sram_cell_6t_5 inst_cell_95_26 (.BL(BL26),.BLN(BLN26),.WL(WL95));
sram_cell_6t_5 inst_cell_95_27 (.BL(BL27),.BLN(BLN27),.WL(WL95));
sram_cell_6t_5 inst_cell_95_28 (.BL(BL28),.BLN(BLN28),.WL(WL95));
sram_cell_6t_5 inst_cell_95_29 (.BL(BL29),.BLN(BLN29),.WL(WL95));
sram_cell_6t_5 inst_cell_95_30 (.BL(BL30),.BLN(BLN30),.WL(WL95));
sram_cell_6t_5 inst_cell_95_31 (.BL(BL31),.BLN(BLN31),.WL(WL95));
sram_cell_6t_5 inst_cell_95_32 (.BL(BL32),.BLN(BLN32),.WL(WL95));
sram_cell_6t_5 inst_cell_95_33 (.BL(BL33),.BLN(BLN33),.WL(WL95));
sram_cell_6t_5 inst_cell_95_34 (.BL(BL34),.BLN(BLN34),.WL(WL95));
sram_cell_6t_5 inst_cell_95_35 (.BL(BL35),.BLN(BLN35),.WL(WL95));
sram_cell_6t_5 inst_cell_95_36 (.BL(BL36),.BLN(BLN36),.WL(WL95));
sram_cell_6t_5 inst_cell_95_37 (.BL(BL37),.BLN(BLN37),.WL(WL95));
sram_cell_6t_5 inst_cell_95_38 (.BL(BL38),.BLN(BLN38),.WL(WL95));
sram_cell_6t_5 inst_cell_95_39 (.BL(BL39),.BLN(BLN39),.WL(WL95));
sram_cell_6t_5 inst_cell_95_40 (.BL(BL40),.BLN(BLN40),.WL(WL95));
sram_cell_6t_5 inst_cell_95_41 (.BL(BL41),.BLN(BLN41),.WL(WL95));
sram_cell_6t_5 inst_cell_95_42 (.BL(BL42),.BLN(BLN42),.WL(WL95));
sram_cell_6t_5 inst_cell_95_43 (.BL(BL43),.BLN(BLN43),.WL(WL95));
sram_cell_6t_5 inst_cell_95_44 (.BL(BL44),.BLN(BLN44),.WL(WL95));
sram_cell_6t_5 inst_cell_95_45 (.BL(BL45),.BLN(BLN45),.WL(WL95));
sram_cell_6t_5 inst_cell_95_46 (.BL(BL46),.BLN(BLN46),.WL(WL95));
sram_cell_6t_5 inst_cell_95_47 (.BL(BL47),.BLN(BLN47),.WL(WL95));
sram_cell_6t_5 inst_cell_95_48 (.BL(BL48),.BLN(BLN48),.WL(WL95));
sram_cell_6t_5 inst_cell_95_49 (.BL(BL49),.BLN(BLN49),.WL(WL95));
sram_cell_6t_5 inst_cell_95_50 (.BL(BL50),.BLN(BLN50),.WL(WL95));
sram_cell_6t_5 inst_cell_95_51 (.BL(BL51),.BLN(BLN51),.WL(WL95));
sram_cell_6t_5 inst_cell_95_52 (.BL(BL52),.BLN(BLN52),.WL(WL95));
sram_cell_6t_5 inst_cell_95_53 (.BL(BL53),.BLN(BLN53),.WL(WL95));
sram_cell_6t_5 inst_cell_95_54 (.BL(BL54),.BLN(BLN54),.WL(WL95));
sram_cell_6t_5 inst_cell_95_55 (.BL(BL55),.BLN(BLN55),.WL(WL95));
sram_cell_6t_5 inst_cell_95_56 (.BL(BL56),.BLN(BLN56),.WL(WL95));
sram_cell_6t_5 inst_cell_95_57 (.BL(BL57),.BLN(BLN57),.WL(WL95));
sram_cell_6t_5 inst_cell_95_58 (.BL(BL58),.BLN(BLN58),.WL(WL95));
sram_cell_6t_5 inst_cell_95_59 (.BL(BL59),.BLN(BLN59),.WL(WL95));
sram_cell_6t_5 inst_cell_95_60 (.BL(BL60),.BLN(BLN60),.WL(WL95));
sram_cell_6t_5 inst_cell_95_61 (.BL(BL61),.BLN(BLN61),.WL(WL95));
sram_cell_6t_5 inst_cell_95_62 (.BL(BL62),.BLN(BLN62),.WL(WL95));
sram_cell_6t_5 inst_cell_95_63 (.BL(BL63),.BLN(BLN63),.WL(WL95));
sram_cell_6t_5 inst_cell_95_64 (.BL(BL64),.BLN(BLN64),.WL(WL95));
sram_cell_6t_5 inst_cell_95_65 (.BL(BL65),.BLN(BLN65),.WL(WL95));
sram_cell_6t_5 inst_cell_95_66 (.BL(BL66),.BLN(BLN66),.WL(WL95));
sram_cell_6t_5 inst_cell_95_67 (.BL(BL67),.BLN(BLN67),.WL(WL95));
sram_cell_6t_5 inst_cell_95_68 (.BL(BL68),.BLN(BLN68),.WL(WL95));
sram_cell_6t_5 inst_cell_95_69 (.BL(BL69),.BLN(BLN69),.WL(WL95));
sram_cell_6t_5 inst_cell_95_70 (.BL(BL70),.BLN(BLN70),.WL(WL95));
sram_cell_6t_5 inst_cell_95_71 (.BL(BL71),.BLN(BLN71),.WL(WL95));
sram_cell_6t_5 inst_cell_95_72 (.BL(BL72),.BLN(BLN72),.WL(WL95));
sram_cell_6t_5 inst_cell_95_73 (.BL(BL73),.BLN(BLN73),.WL(WL95));
sram_cell_6t_5 inst_cell_95_74 (.BL(BL74),.BLN(BLN74),.WL(WL95));
sram_cell_6t_5 inst_cell_95_75 (.BL(BL75),.BLN(BLN75),.WL(WL95));
sram_cell_6t_5 inst_cell_95_76 (.BL(BL76),.BLN(BLN76),.WL(WL95));
sram_cell_6t_5 inst_cell_95_77 (.BL(BL77),.BLN(BLN77),.WL(WL95));
sram_cell_6t_5 inst_cell_95_78 (.BL(BL78),.BLN(BLN78),.WL(WL95));
sram_cell_6t_5 inst_cell_95_79 (.BL(BL79),.BLN(BLN79),.WL(WL95));
sram_cell_6t_5 inst_cell_95_80 (.BL(BL80),.BLN(BLN80),.WL(WL95));
sram_cell_6t_5 inst_cell_95_81 (.BL(BL81),.BLN(BLN81),.WL(WL95));
sram_cell_6t_5 inst_cell_95_82 (.BL(BL82),.BLN(BLN82),.WL(WL95));
sram_cell_6t_5 inst_cell_95_83 (.BL(BL83),.BLN(BLN83),.WL(WL95));
sram_cell_6t_5 inst_cell_95_84 (.BL(BL84),.BLN(BLN84),.WL(WL95));
sram_cell_6t_5 inst_cell_95_85 (.BL(BL85),.BLN(BLN85),.WL(WL95));
sram_cell_6t_5 inst_cell_95_86 (.BL(BL86),.BLN(BLN86),.WL(WL95));
sram_cell_6t_5 inst_cell_95_87 (.BL(BL87),.BLN(BLN87),.WL(WL95));
sram_cell_6t_5 inst_cell_95_88 (.BL(BL88),.BLN(BLN88),.WL(WL95));
sram_cell_6t_5 inst_cell_95_89 (.BL(BL89),.BLN(BLN89),.WL(WL95));
sram_cell_6t_5 inst_cell_95_90 (.BL(BL90),.BLN(BLN90),.WL(WL95));
sram_cell_6t_5 inst_cell_95_91 (.BL(BL91),.BLN(BLN91),.WL(WL95));
sram_cell_6t_5 inst_cell_95_92 (.BL(BL92),.BLN(BLN92),.WL(WL95));
sram_cell_6t_5 inst_cell_95_93 (.BL(BL93),.BLN(BLN93),.WL(WL95));
sram_cell_6t_5 inst_cell_95_94 (.BL(BL94),.BLN(BLN94),.WL(WL95));
sram_cell_6t_5 inst_cell_95_95 (.BL(BL95),.BLN(BLN95),.WL(WL95));
sram_cell_6t_5 inst_cell_95_96 (.BL(BL96),.BLN(BLN96),.WL(WL95));
sram_cell_6t_5 inst_cell_95_97 (.BL(BL97),.BLN(BLN97),.WL(WL95));
sram_cell_6t_5 inst_cell_95_98 (.BL(BL98),.BLN(BLN98),.WL(WL95));
sram_cell_6t_5 inst_cell_95_99 (.BL(BL99),.BLN(BLN99),.WL(WL95));
sram_cell_6t_5 inst_cell_95_100 (.BL(BL100),.BLN(BLN100),.WL(WL95));
sram_cell_6t_5 inst_cell_95_101 (.BL(BL101),.BLN(BLN101),.WL(WL95));
sram_cell_6t_5 inst_cell_95_102 (.BL(BL102),.BLN(BLN102),.WL(WL95));
sram_cell_6t_5 inst_cell_95_103 (.BL(BL103),.BLN(BLN103),.WL(WL95));
sram_cell_6t_5 inst_cell_95_104 (.BL(BL104),.BLN(BLN104),.WL(WL95));
sram_cell_6t_5 inst_cell_95_105 (.BL(BL105),.BLN(BLN105),.WL(WL95));
sram_cell_6t_5 inst_cell_95_106 (.BL(BL106),.BLN(BLN106),.WL(WL95));
sram_cell_6t_5 inst_cell_95_107 (.BL(BL107),.BLN(BLN107),.WL(WL95));
sram_cell_6t_5 inst_cell_95_108 (.BL(BL108),.BLN(BLN108),.WL(WL95));
sram_cell_6t_5 inst_cell_95_109 (.BL(BL109),.BLN(BLN109),.WL(WL95));
sram_cell_6t_5 inst_cell_95_110 (.BL(BL110),.BLN(BLN110),.WL(WL95));
sram_cell_6t_5 inst_cell_95_111 (.BL(BL111),.BLN(BLN111),.WL(WL95));
sram_cell_6t_5 inst_cell_95_112 (.BL(BL112),.BLN(BLN112),.WL(WL95));
sram_cell_6t_5 inst_cell_95_113 (.BL(BL113),.BLN(BLN113),.WL(WL95));
sram_cell_6t_5 inst_cell_95_114 (.BL(BL114),.BLN(BLN114),.WL(WL95));
sram_cell_6t_5 inst_cell_95_115 (.BL(BL115),.BLN(BLN115),.WL(WL95));
sram_cell_6t_5 inst_cell_95_116 (.BL(BL116),.BLN(BLN116),.WL(WL95));
sram_cell_6t_5 inst_cell_95_117 (.BL(BL117),.BLN(BLN117),.WL(WL95));
sram_cell_6t_5 inst_cell_95_118 (.BL(BL118),.BLN(BLN118),.WL(WL95));
sram_cell_6t_5 inst_cell_95_119 (.BL(BL119),.BLN(BLN119),.WL(WL95));
sram_cell_6t_5 inst_cell_95_120 (.BL(BL120),.BLN(BLN120),.WL(WL95));
sram_cell_6t_5 inst_cell_95_121 (.BL(BL121),.BLN(BLN121),.WL(WL95));
sram_cell_6t_5 inst_cell_95_122 (.BL(BL122),.BLN(BLN122),.WL(WL95));
sram_cell_6t_5 inst_cell_95_123 (.BL(BL123),.BLN(BLN123),.WL(WL95));
sram_cell_6t_5 inst_cell_95_124 (.BL(BL124),.BLN(BLN124),.WL(WL95));
sram_cell_6t_5 inst_cell_95_125 (.BL(BL125),.BLN(BLN125),.WL(WL95));
sram_cell_6t_5 inst_cell_95_126 (.BL(BL126),.BLN(BLN126),.WL(WL95));
sram_cell_6t_5 inst_cell_95_127 (.BL(BL127),.BLN(BLN127),.WL(WL95));
sram_cell_6t_5 inst_cell_96_0 (.BL(BL0),.BLN(BLN0),.WL(WL96));
sram_cell_6t_5 inst_cell_96_1 (.BL(BL1),.BLN(BLN1),.WL(WL96));
sram_cell_6t_5 inst_cell_96_2 (.BL(BL2),.BLN(BLN2),.WL(WL96));
sram_cell_6t_5 inst_cell_96_3 (.BL(BL3),.BLN(BLN3),.WL(WL96));
sram_cell_6t_5 inst_cell_96_4 (.BL(BL4),.BLN(BLN4),.WL(WL96));
sram_cell_6t_5 inst_cell_96_5 (.BL(BL5),.BLN(BLN5),.WL(WL96));
sram_cell_6t_5 inst_cell_96_6 (.BL(BL6),.BLN(BLN6),.WL(WL96));
sram_cell_6t_5 inst_cell_96_7 (.BL(BL7),.BLN(BLN7),.WL(WL96));
sram_cell_6t_5 inst_cell_96_8 (.BL(BL8),.BLN(BLN8),.WL(WL96));
sram_cell_6t_5 inst_cell_96_9 (.BL(BL9),.BLN(BLN9),.WL(WL96));
sram_cell_6t_5 inst_cell_96_10 (.BL(BL10),.BLN(BLN10),.WL(WL96));
sram_cell_6t_5 inst_cell_96_11 (.BL(BL11),.BLN(BLN11),.WL(WL96));
sram_cell_6t_5 inst_cell_96_12 (.BL(BL12),.BLN(BLN12),.WL(WL96));
sram_cell_6t_5 inst_cell_96_13 (.BL(BL13),.BLN(BLN13),.WL(WL96));
sram_cell_6t_5 inst_cell_96_14 (.BL(BL14),.BLN(BLN14),.WL(WL96));
sram_cell_6t_5 inst_cell_96_15 (.BL(BL15),.BLN(BLN15),.WL(WL96));
sram_cell_6t_5 inst_cell_96_16 (.BL(BL16),.BLN(BLN16),.WL(WL96));
sram_cell_6t_5 inst_cell_96_17 (.BL(BL17),.BLN(BLN17),.WL(WL96));
sram_cell_6t_5 inst_cell_96_18 (.BL(BL18),.BLN(BLN18),.WL(WL96));
sram_cell_6t_5 inst_cell_96_19 (.BL(BL19),.BLN(BLN19),.WL(WL96));
sram_cell_6t_5 inst_cell_96_20 (.BL(BL20),.BLN(BLN20),.WL(WL96));
sram_cell_6t_5 inst_cell_96_21 (.BL(BL21),.BLN(BLN21),.WL(WL96));
sram_cell_6t_5 inst_cell_96_22 (.BL(BL22),.BLN(BLN22),.WL(WL96));
sram_cell_6t_5 inst_cell_96_23 (.BL(BL23),.BLN(BLN23),.WL(WL96));
sram_cell_6t_5 inst_cell_96_24 (.BL(BL24),.BLN(BLN24),.WL(WL96));
sram_cell_6t_5 inst_cell_96_25 (.BL(BL25),.BLN(BLN25),.WL(WL96));
sram_cell_6t_5 inst_cell_96_26 (.BL(BL26),.BLN(BLN26),.WL(WL96));
sram_cell_6t_5 inst_cell_96_27 (.BL(BL27),.BLN(BLN27),.WL(WL96));
sram_cell_6t_5 inst_cell_96_28 (.BL(BL28),.BLN(BLN28),.WL(WL96));
sram_cell_6t_5 inst_cell_96_29 (.BL(BL29),.BLN(BLN29),.WL(WL96));
sram_cell_6t_5 inst_cell_96_30 (.BL(BL30),.BLN(BLN30),.WL(WL96));
sram_cell_6t_5 inst_cell_96_31 (.BL(BL31),.BLN(BLN31),.WL(WL96));
sram_cell_6t_5 inst_cell_96_32 (.BL(BL32),.BLN(BLN32),.WL(WL96));
sram_cell_6t_5 inst_cell_96_33 (.BL(BL33),.BLN(BLN33),.WL(WL96));
sram_cell_6t_5 inst_cell_96_34 (.BL(BL34),.BLN(BLN34),.WL(WL96));
sram_cell_6t_5 inst_cell_96_35 (.BL(BL35),.BLN(BLN35),.WL(WL96));
sram_cell_6t_5 inst_cell_96_36 (.BL(BL36),.BLN(BLN36),.WL(WL96));
sram_cell_6t_5 inst_cell_96_37 (.BL(BL37),.BLN(BLN37),.WL(WL96));
sram_cell_6t_5 inst_cell_96_38 (.BL(BL38),.BLN(BLN38),.WL(WL96));
sram_cell_6t_5 inst_cell_96_39 (.BL(BL39),.BLN(BLN39),.WL(WL96));
sram_cell_6t_5 inst_cell_96_40 (.BL(BL40),.BLN(BLN40),.WL(WL96));
sram_cell_6t_5 inst_cell_96_41 (.BL(BL41),.BLN(BLN41),.WL(WL96));
sram_cell_6t_5 inst_cell_96_42 (.BL(BL42),.BLN(BLN42),.WL(WL96));
sram_cell_6t_5 inst_cell_96_43 (.BL(BL43),.BLN(BLN43),.WL(WL96));
sram_cell_6t_5 inst_cell_96_44 (.BL(BL44),.BLN(BLN44),.WL(WL96));
sram_cell_6t_5 inst_cell_96_45 (.BL(BL45),.BLN(BLN45),.WL(WL96));
sram_cell_6t_5 inst_cell_96_46 (.BL(BL46),.BLN(BLN46),.WL(WL96));
sram_cell_6t_5 inst_cell_96_47 (.BL(BL47),.BLN(BLN47),.WL(WL96));
sram_cell_6t_5 inst_cell_96_48 (.BL(BL48),.BLN(BLN48),.WL(WL96));
sram_cell_6t_5 inst_cell_96_49 (.BL(BL49),.BLN(BLN49),.WL(WL96));
sram_cell_6t_5 inst_cell_96_50 (.BL(BL50),.BLN(BLN50),.WL(WL96));
sram_cell_6t_5 inst_cell_96_51 (.BL(BL51),.BLN(BLN51),.WL(WL96));
sram_cell_6t_5 inst_cell_96_52 (.BL(BL52),.BLN(BLN52),.WL(WL96));
sram_cell_6t_5 inst_cell_96_53 (.BL(BL53),.BLN(BLN53),.WL(WL96));
sram_cell_6t_5 inst_cell_96_54 (.BL(BL54),.BLN(BLN54),.WL(WL96));
sram_cell_6t_5 inst_cell_96_55 (.BL(BL55),.BLN(BLN55),.WL(WL96));
sram_cell_6t_5 inst_cell_96_56 (.BL(BL56),.BLN(BLN56),.WL(WL96));
sram_cell_6t_5 inst_cell_96_57 (.BL(BL57),.BLN(BLN57),.WL(WL96));
sram_cell_6t_5 inst_cell_96_58 (.BL(BL58),.BLN(BLN58),.WL(WL96));
sram_cell_6t_5 inst_cell_96_59 (.BL(BL59),.BLN(BLN59),.WL(WL96));
sram_cell_6t_5 inst_cell_96_60 (.BL(BL60),.BLN(BLN60),.WL(WL96));
sram_cell_6t_5 inst_cell_96_61 (.BL(BL61),.BLN(BLN61),.WL(WL96));
sram_cell_6t_5 inst_cell_96_62 (.BL(BL62),.BLN(BLN62),.WL(WL96));
sram_cell_6t_5 inst_cell_96_63 (.BL(BL63),.BLN(BLN63),.WL(WL96));
sram_cell_6t_5 inst_cell_96_64 (.BL(BL64),.BLN(BLN64),.WL(WL96));
sram_cell_6t_5 inst_cell_96_65 (.BL(BL65),.BLN(BLN65),.WL(WL96));
sram_cell_6t_5 inst_cell_96_66 (.BL(BL66),.BLN(BLN66),.WL(WL96));
sram_cell_6t_5 inst_cell_96_67 (.BL(BL67),.BLN(BLN67),.WL(WL96));
sram_cell_6t_5 inst_cell_96_68 (.BL(BL68),.BLN(BLN68),.WL(WL96));
sram_cell_6t_5 inst_cell_96_69 (.BL(BL69),.BLN(BLN69),.WL(WL96));
sram_cell_6t_5 inst_cell_96_70 (.BL(BL70),.BLN(BLN70),.WL(WL96));
sram_cell_6t_5 inst_cell_96_71 (.BL(BL71),.BLN(BLN71),.WL(WL96));
sram_cell_6t_5 inst_cell_96_72 (.BL(BL72),.BLN(BLN72),.WL(WL96));
sram_cell_6t_5 inst_cell_96_73 (.BL(BL73),.BLN(BLN73),.WL(WL96));
sram_cell_6t_5 inst_cell_96_74 (.BL(BL74),.BLN(BLN74),.WL(WL96));
sram_cell_6t_5 inst_cell_96_75 (.BL(BL75),.BLN(BLN75),.WL(WL96));
sram_cell_6t_5 inst_cell_96_76 (.BL(BL76),.BLN(BLN76),.WL(WL96));
sram_cell_6t_5 inst_cell_96_77 (.BL(BL77),.BLN(BLN77),.WL(WL96));
sram_cell_6t_5 inst_cell_96_78 (.BL(BL78),.BLN(BLN78),.WL(WL96));
sram_cell_6t_5 inst_cell_96_79 (.BL(BL79),.BLN(BLN79),.WL(WL96));
sram_cell_6t_5 inst_cell_96_80 (.BL(BL80),.BLN(BLN80),.WL(WL96));
sram_cell_6t_5 inst_cell_96_81 (.BL(BL81),.BLN(BLN81),.WL(WL96));
sram_cell_6t_5 inst_cell_96_82 (.BL(BL82),.BLN(BLN82),.WL(WL96));
sram_cell_6t_5 inst_cell_96_83 (.BL(BL83),.BLN(BLN83),.WL(WL96));
sram_cell_6t_5 inst_cell_96_84 (.BL(BL84),.BLN(BLN84),.WL(WL96));
sram_cell_6t_5 inst_cell_96_85 (.BL(BL85),.BLN(BLN85),.WL(WL96));
sram_cell_6t_5 inst_cell_96_86 (.BL(BL86),.BLN(BLN86),.WL(WL96));
sram_cell_6t_5 inst_cell_96_87 (.BL(BL87),.BLN(BLN87),.WL(WL96));
sram_cell_6t_5 inst_cell_96_88 (.BL(BL88),.BLN(BLN88),.WL(WL96));
sram_cell_6t_5 inst_cell_96_89 (.BL(BL89),.BLN(BLN89),.WL(WL96));
sram_cell_6t_5 inst_cell_96_90 (.BL(BL90),.BLN(BLN90),.WL(WL96));
sram_cell_6t_5 inst_cell_96_91 (.BL(BL91),.BLN(BLN91),.WL(WL96));
sram_cell_6t_5 inst_cell_96_92 (.BL(BL92),.BLN(BLN92),.WL(WL96));
sram_cell_6t_5 inst_cell_96_93 (.BL(BL93),.BLN(BLN93),.WL(WL96));
sram_cell_6t_5 inst_cell_96_94 (.BL(BL94),.BLN(BLN94),.WL(WL96));
sram_cell_6t_5 inst_cell_96_95 (.BL(BL95),.BLN(BLN95),.WL(WL96));
sram_cell_6t_5 inst_cell_96_96 (.BL(BL96),.BLN(BLN96),.WL(WL96));
sram_cell_6t_5 inst_cell_96_97 (.BL(BL97),.BLN(BLN97),.WL(WL96));
sram_cell_6t_5 inst_cell_96_98 (.BL(BL98),.BLN(BLN98),.WL(WL96));
sram_cell_6t_5 inst_cell_96_99 (.BL(BL99),.BLN(BLN99),.WL(WL96));
sram_cell_6t_5 inst_cell_96_100 (.BL(BL100),.BLN(BLN100),.WL(WL96));
sram_cell_6t_5 inst_cell_96_101 (.BL(BL101),.BLN(BLN101),.WL(WL96));
sram_cell_6t_5 inst_cell_96_102 (.BL(BL102),.BLN(BLN102),.WL(WL96));
sram_cell_6t_5 inst_cell_96_103 (.BL(BL103),.BLN(BLN103),.WL(WL96));
sram_cell_6t_5 inst_cell_96_104 (.BL(BL104),.BLN(BLN104),.WL(WL96));
sram_cell_6t_5 inst_cell_96_105 (.BL(BL105),.BLN(BLN105),.WL(WL96));
sram_cell_6t_5 inst_cell_96_106 (.BL(BL106),.BLN(BLN106),.WL(WL96));
sram_cell_6t_5 inst_cell_96_107 (.BL(BL107),.BLN(BLN107),.WL(WL96));
sram_cell_6t_5 inst_cell_96_108 (.BL(BL108),.BLN(BLN108),.WL(WL96));
sram_cell_6t_5 inst_cell_96_109 (.BL(BL109),.BLN(BLN109),.WL(WL96));
sram_cell_6t_5 inst_cell_96_110 (.BL(BL110),.BLN(BLN110),.WL(WL96));
sram_cell_6t_5 inst_cell_96_111 (.BL(BL111),.BLN(BLN111),.WL(WL96));
sram_cell_6t_5 inst_cell_96_112 (.BL(BL112),.BLN(BLN112),.WL(WL96));
sram_cell_6t_5 inst_cell_96_113 (.BL(BL113),.BLN(BLN113),.WL(WL96));
sram_cell_6t_5 inst_cell_96_114 (.BL(BL114),.BLN(BLN114),.WL(WL96));
sram_cell_6t_5 inst_cell_96_115 (.BL(BL115),.BLN(BLN115),.WL(WL96));
sram_cell_6t_5 inst_cell_96_116 (.BL(BL116),.BLN(BLN116),.WL(WL96));
sram_cell_6t_5 inst_cell_96_117 (.BL(BL117),.BLN(BLN117),.WL(WL96));
sram_cell_6t_5 inst_cell_96_118 (.BL(BL118),.BLN(BLN118),.WL(WL96));
sram_cell_6t_5 inst_cell_96_119 (.BL(BL119),.BLN(BLN119),.WL(WL96));
sram_cell_6t_5 inst_cell_96_120 (.BL(BL120),.BLN(BLN120),.WL(WL96));
sram_cell_6t_5 inst_cell_96_121 (.BL(BL121),.BLN(BLN121),.WL(WL96));
sram_cell_6t_5 inst_cell_96_122 (.BL(BL122),.BLN(BLN122),.WL(WL96));
sram_cell_6t_5 inst_cell_96_123 (.BL(BL123),.BLN(BLN123),.WL(WL96));
sram_cell_6t_5 inst_cell_96_124 (.BL(BL124),.BLN(BLN124),.WL(WL96));
sram_cell_6t_5 inst_cell_96_125 (.BL(BL125),.BLN(BLN125),.WL(WL96));
sram_cell_6t_5 inst_cell_96_126 (.BL(BL126),.BLN(BLN126),.WL(WL96));
sram_cell_6t_5 inst_cell_96_127 (.BL(BL127),.BLN(BLN127),.WL(WL96));
sram_cell_6t_5 inst_cell_97_0 (.BL(BL0),.BLN(BLN0),.WL(WL97));
sram_cell_6t_5 inst_cell_97_1 (.BL(BL1),.BLN(BLN1),.WL(WL97));
sram_cell_6t_5 inst_cell_97_2 (.BL(BL2),.BLN(BLN2),.WL(WL97));
sram_cell_6t_5 inst_cell_97_3 (.BL(BL3),.BLN(BLN3),.WL(WL97));
sram_cell_6t_5 inst_cell_97_4 (.BL(BL4),.BLN(BLN4),.WL(WL97));
sram_cell_6t_5 inst_cell_97_5 (.BL(BL5),.BLN(BLN5),.WL(WL97));
sram_cell_6t_5 inst_cell_97_6 (.BL(BL6),.BLN(BLN6),.WL(WL97));
sram_cell_6t_5 inst_cell_97_7 (.BL(BL7),.BLN(BLN7),.WL(WL97));
sram_cell_6t_5 inst_cell_97_8 (.BL(BL8),.BLN(BLN8),.WL(WL97));
sram_cell_6t_5 inst_cell_97_9 (.BL(BL9),.BLN(BLN9),.WL(WL97));
sram_cell_6t_5 inst_cell_97_10 (.BL(BL10),.BLN(BLN10),.WL(WL97));
sram_cell_6t_5 inst_cell_97_11 (.BL(BL11),.BLN(BLN11),.WL(WL97));
sram_cell_6t_5 inst_cell_97_12 (.BL(BL12),.BLN(BLN12),.WL(WL97));
sram_cell_6t_5 inst_cell_97_13 (.BL(BL13),.BLN(BLN13),.WL(WL97));
sram_cell_6t_5 inst_cell_97_14 (.BL(BL14),.BLN(BLN14),.WL(WL97));
sram_cell_6t_5 inst_cell_97_15 (.BL(BL15),.BLN(BLN15),.WL(WL97));
sram_cell_6t_5 inst_cell_97_16 (.BL(BL16),.BLN(BLN16),.WL(WL97));
sram_cell_6t_5 inst_cell_97_17 (.BL(BL17),.BLN(BLN17),.WL(WL97));
sram_cell_6t_5 inst_cell_97_18 (.BL(BL18),.BLN(BLN18),.WL(WL97));
sram_cell_6t_5 inst_cell_97_19 (.BL(BL19),.BLN(BLN19),.WL(WL97));
sram_cell_6t_5 inst_cell_97_20 (.BL(BL20),.BLN(BLN20),.WL(WL97));
sram_cell_6t_5 inst_cell_97_21 (.BL(BL21),.BLN(BLN21),.WL(WL97));
sram_cell_6t_5 inst_cell_97_22 (.BL(BL22),.BLN(BLN22),.WL(WL97));
sram_cell_6t_5 inst_cell_97_23 (.BL(BL23),.BLN(BLN23),.WL(WL97));
sram_cell_6t_5 inst_cell_97_24 (.BL(BL24),.BLN(BLN24),.WL(WL97));
sram_cell_6t_5 inst_cell_97_25 (.BL(BL25),.BLN(BLN25),.WL(WL97));
sram_cell_6t_5 inst_cell_97_26 (.BL(BL26),.BLN(BLN26),.WL(WL97));
sram_cell_6t_5 inst_cell_97_27 (.BL(BL27),.BLN(BLN27),.WL(WL97));
sram_cell_6t_5 inst_cell_97_28 (.BL(BL28),.BLN(BLN28),.WL(WL97));
sram_cell_6t_5 inst_cell_97_29 (.BL(BL29),.BLN(BLN29),.WL(WL97));
sram_cell_6t_5 inst_cell_97_30 (.BL(BL30),.BLN(BLN30),.WL(WL97));
sram_cell_6t_5 inst_cell_97_31 (.BL(BL31),.BLN(BLN31),.WL(WL97));
sram_cell_6t_5 inst_cell_97_32 (.BL(BL32),.BLN(BLN32),.WL(WL97));
sram_cell_6t_5 inst_cell_97_33 (.BL(BL33),.BLN(BLN33),.WL(WL97));
sram_cell_6t_5 inst_cell_97_34 (.BL(BL34),.BLN(BLN34),.WL(WL97));
sram_cell_6t_5 inst_cell_97_35 (.BL(BL35),.BLN(BLN35),.WL(WL97));
sram_cell_6t_5 inst_cell_97_36 (.BL(BL36),.BLN(BLN36),.WL(WL97));
sram_cell_6t_5 inst_cell_97_37 (.BL(BL37),.BLN(BLN37),.WL(WL97));
sram_cell_6t_5 inst_cell_97_38 (.BL(BL38),.BLN(BLN38),.WL(WL97));
sram_cell_6t_5 inst_cell_97_39 (.BL(BL39),.BLN(BLN39),.WL(WL97));
sram_cell_6t_5 inst_cell_97_40 (.BL(BL40),.BLN(BLN40),.WL(WL97));
sram_cell_6t_5 inst_cell_97_41 (.BL(BL41),.BLN(BLN41),.WL(WL97));
sram_cell_6t_5 inst_cell_97_42 (.BL(BL42),.BLN(BLN42),.WL(WL97));
sram_cell_6t_5 inst_cell_97_43 (.BL(BL43),.BLN(BLN43),.WL(WL97));
sram_cell_6t_5 inst_cell_97_44 (.BL(BL44),.BLN(BLN44),.WL(WL97));
sram_cell_6t_5 inst_cell_97_45 (.BL(BL45),.BLN(BLN45),.WL(WL97));
sram_cell_6t_5 inst_cell_97_46 (.BL(BL46),.BLN(BLN46),.WL(WL97));
sram_cell_6t_5 inst_cell_97_47 (.BL(BL47),.BLN(BLN47),.WL(WL97));
sram_cell_6t_5 inst_cell_97_48 (.BL(BL48),.BLN(BLN48),.WL(WL97));
sram_cell_6t_5 inst_cell_97_49 (.BL(BL49),.BLN(BLN49),.WL(WL97));
sram_cell_6t_5 inst_cell_97_50 (.BL(BL50),.BLN(BLN50),.WL(WL97));
sram_cell_6t_5 inst_cell_97_51 (.BL(BL51),.BLN(BLN51),.WL(WL97));
sram_cell_6t_5 inst_cell_97_52 (.BL(BL52),.BLN(BLN52),.WL(WL97));
sram_cell_6t_5 inst_cell_97_53 (.BL(BL53),.BLN(BLN53),.WL(WL97));
sram_cell_6t_5 inst_cell_97_54 (.BL(BL54),.BLN(BLN54),.WL(WL97));
sram_cell_6t_5 inst_cell_97_55 (.BL(BL55),.BLN(BLN55),.WL(WL97));
sram_cell_6t_5 inst_cell_97_56 (.BL(BL56),.BLN(BLN56),.WL(WL97));
sram_cell_6t_5 inst_cell_97_57 (.BL(BL57),.BLN(BLN57),.WL(WL97));
sram_cell_6t_5 inst_cell_97_58 (.BL(BL58),.BLN(BLN58),.WL(WL97));
sram_cell_6t_5 inst_cell_97_59 (.BL(BL59),.BLN(BLN59),.WL(WL97));
sram_cell_6t_5 inst_cell_97_60 (.BL(BL60),.BLN(BLN60),.WL(WL97));
sram_cell_6t_5 inst_cell_97_61 (.BL(BL61),.BLN(BLN61),.WL(WL97));
sram_cell_6t_5 inst_cell_97_62 (.BL(BL62),.BLN(BLN62),.WL(WL97));
sram_cell_6t_5 inst_cell_97_63 (.BL(BL63),.BLN(BLN63),.WL(WL97));
sram_cell_6t_5 inst_cell_97_64 (.BL(BL64),.BLN(BLN64),.WL(WL97));
sram_cell_6t_5 inst_cell_97_65 (.BL(BL65),.BLN(BLN65),.WL(WL97));
sram_cell_6t_5 inst_cell_97_66 (.BL(BL66),.BLN(BLN66),.WL(WL97));
sram_cell_6t_5 inst_cell_97_67 (.BL(BL67),.BLN(BLN67),.WL(WL97));
sram_cell_6t_5 inst_cell_97_68 (.BL(BL68),.BLN(BLN68),.WL(WL97));
sram_cell_6t_5 inst_cell_97_69 (.BL(BL69),.BLN(BLN69),.WL(WL97));
sram_cell_6t_5 inst_cell_97_70 (.BL(BL70),.BLN(BLN70),.WL(WL97));
sram_cell_6t_5 inst_cell_97_71 (.BL(BL71),.BLN(BLN71),.WL(WL97));
sram_cell_6t_5 inst_cell_97_72 (.BL(BL72),.BLN(BLN72),.WL(WL97));
sram_cell_6t_5 inst_cell_97_73 (.BL(BL73),.BLN(BLN73),.WL(WL97));
sram_cell_6t_5 inst_cell_97_74 (.BL(BL74),.BLN(BLN74),.WL(WL97));
sram_cell_6t_5 inst_cell_97_75 (.BL(BL75),.BLN(BLN75),.WL(WL97));
sram_cell_6t_5 inst_cell_97_76 (.BL(BL76),.BLN(BLN76),.WL(WL97));
sram_cell_6t_5 inst_cell_97_77 (.BL(BL77),.BLN(BLN77),.WL(WL97));
sram_cell_6t_5 inst_cell_97_78 (.BL(BL78),.BLN(BLN78),.WL(WL97));
sram_cell_6t_5 inst_cell_97_79 (.BL(BL79),.BLN(BLN79),.WL(WL97));
sram_cell_6t_5 inst_cell_97_80 (.BL(BL80),.BLN(BLN80),.WL(WL97));
sram_cell_6t_5 inst_cell_97_81 (.BL(BL81),.BLN(BLN81),.WL(WL97));
sram_cell_6t_5 inst_cell_97_82 (.BL(BL82),.BLN(BLN82),.WL(WL97));
sram_cell_6t_5 inst_cell_97_83 (.BL(BL83),.BLN(BLN83),.WL(WL97));
sram_cell_6t_5 inst_cell_97_84 (.BL(BL84),.BLN(BLN84),.WL(WL97));
sram_cell_6t_5 inst_cell_97_85 (.BL(BL85),.BLN(BLN85),.WL(WL97));
sram_cell_6t_5 inst_cell_97_86 (.BL(BL86),.BLN(BLN86),.WL(WL97));
sram_cell_6t_5 inst_cell_97_87 (.BL(BL87),.BLN(BLN87),.WL(WL97));
sram_cell_6t_5 inst_cell_97_88 (.BL(BL88),.BLN(BLN88),.WL(WL97));
sram_cell_6t_5 inst_cell_97_89 (.BL(BL89),.BLN(BLN89),.WL(WL97));
sram_cell_6t_5 inst_cell_97_90 (.BL(BL90),.BLN(BLN90),.WL(WL97));
sram_cell_6t_5 inst_cell_97_91 (.BL(BL91),.BLN(BLN91),.WL(WL97));
sram_cell_6t_5 inst_cell_97_92 (.BL(BL92),.BLN(BLN92),.WL(WL97));
sram_cell_6t_5 inst_cell_97_93 (.BL(BL93),.BLN(BLN93),.WL(WL97));
sram_cell_6t_5 inst_cell_97_94 (.BL(BL94),.BLN(BLN94),.WL(WL97));
sram_cell_6t_5 inst_cell_97_95 (.BL(BL95),.BLN(BLN95),.WL(WL97));
sram_cell_6t_5 inst_cell_97_96 (.BL(BL96),.BLN(BLN96),.WL(WL97));
sram_cell_6t_5 inst_cell_97_97 (.BL(BL97),.BLN(BLN97),.WL(WL97));
sram_cell_6t_5 inst_cell_97_98 (.BL(BL98),.BLN(BLN98),.WL(WL97));
sram_cell_6t_5 inst_cell_97_99 (.BL(BL99),.BLN(BLN99),.WL(WL97));
sram_cell_6t_5 inst_cell_97_100 (.BL(BL100),.BLN(BLN100),.WL(WL97));
sram_cell_6t_5 inst_cell_97_101 (.BL(BL101),.BLN(BLN101),.WL(WL97));
sram_cell_6t_5 inst_cell_97_102 (.BL(BL102),.BLN(BLN102),.WL(WL97));
sram_cell_6t_5 inst_cell_97_103 (.BL(BL103),.BLN(BLN103),.WL(WL97));
sram_cell_6t_5 inst_cell_97_104 (.BL(BL104),.BLN(BLN104),.WL(WL97));
sram_cell_6t_5 inst_cell_97_105 (.BL(BL105),.BLN(BLN105),.WL(WL97));
sram_cell_6t_5 inst_cell_97_106 (.BL(BL106),.BLN(BLN106),.WL(WL97));
sram_cell_6t_5 inst_cell_97_107 (.BL(BL107),.BLN(BLN107),.WL(WL97));
sram_cell_6t_5 inst_cell_97_108 (.BL(BL108),.BLN(BLN108),.WL(WL97));
sram_cell_6t_5 inst_cell_97_109 (.BL(BL109),.BLN(BLN109),.WL(WL97));
sram_cell_6t_5 inst_cell_97_110 (.BL(BL110),.BLN(BLN110),.WL(WL97));
sram_cell_6t_5 inst_cell_97_111 (.BL(BL111),.BLN(BLN111),.WL(WL97));
sram_cell_6t_5 inst_cell_97_112 (.BL(BL112),.BLN(BLN112),.WL(WL97));
sram_cell_6t_5 inst_cell_97_113 (.BL(BL113),.BLN(BLN113),.WL(WL97));
sram_cell_6t_5 inst_cell_97_114 (.BL(BL114),.BLN(BLN114),.WL(WL97));
sram_cell_6t_5 inst_cell_97_115 (.BL(BL115),.BLN(BLN115),.WL(WL97));
sram_cell_6t_5 inst_cell_97_116 (.BL(BL116),.BLN(BLN116),.WL(WL97));
sram_cell_6t_5 inst_cell_97_117 (.BL(BL117),.BLN(BLN117),.WL(WL97));
sram_cell_6t_5 inst_cell_97_118 (.BL(BL118),.BLN(BLN118),.WL(WL97));
sram_cell_6t_5 inst_cell_97_119 (.BL(BL119),.BLN(BLN119),.WL(WL97));
sram_cell_6t_5 inst_cell_97_120 (.BL(BL120),.BLN(BLN120),.WL(WL97));
sram_cell_6t_5 inst_cell_97_121 (.BL(BL121),.BLN(BLN121),.WL(WL97));
sram_cell_6t_5 inst_cell_97_122 (.BL(BL122),.BLN(BLN122),.WL(WL97));
sram_cell_6t_5 inst_cell_97_123 (.BL(BL123),.BLN(BLN123),.WL(WL97));
sram_cell_6t_5 inst_cell_97_124 (.BL(BL124),.BLN(BLN124),.WL(WL97));
sram_cell_6t_5 inst_cell_97_125 (.BL(BL125),.BLN(BLN125),.WL(WL97));
sram_cell_6t_5 inst_cell_97_126 (.BL(BL126),.BLN(BLN126),.WL(WL97));
sram_cell_6t_5 inst_cell_97_127 (.BL(BL127),.BLN(BLN127),.WL(WL97));
sram_cell_6t_5 inst_cell_98_0 (.BL(BL0),.BLN(BLN0),.WL(WL98));
sram_cell_6t_5 inst_cell_98_1 (.BL(BL1),.BLN(BLN1),.WL(WL98));
sram_cell_6t_5 inst_cell_98_2 (.BL(BL2),.BLN(BLN2),.WL(WL98));
sram_cell_6t_5 inst_cell_98_3 (.BL(BL3),.BLN(BLN3),.WL(WL98));
sram_cell_6t_5 inst_cell_98_4 (.BL(BL4),.BLN(BLN4),.WL(WL98));
sram_cell_6t_5 inst_cell_98_5 (.BL(BL5),.BLN(BLN5),.WL(WL98));
sram_cell_6t_5 inst_cell_98_6 (.BL(BL6),.BLN(BLN6),.WL(WL98));
sram_cell_6t_5 inst_cell_98_7 (.BL(BL7),.BLN(BLN7),.WL(WL98));
sram_cell_6t_5 inst_cell_98_8 (.BL(BL8),.BLN(BLN8),.WL(WL98));
sram_cell_6t_5 inst_cell_98_9 (.BL(BL9),.BLN(BLN9),.WL(WL98));
sram_cell_6t_5 inst_cell_98_10 (.BL(BL10),.BLN(BLN10),.WL(WL98));
sram_cell_6t_5 inst_cell_98_11 (.BL(BL11),.BLN(BLN11),.WL(WL98));
sram_cell_6t_5 inst_cell_98_12 (.BL(BL12),.BLN(BLN12),.WL(WL98));
sram_cell_6t_5 inst_cell_98_13 (.BL(BL13),.BLN(BLN13),.WL(WL98));
sram_cell_6t_5 inst_cell_98_14 (.BL(BL14),.BLN(BLN14),.WL(WL98));
sram_cell_6t_5 inst_cell_98_15 (.BL(BL15),.BLN(BLN15),.WL(WL98));
sram_cell_6t_5 inst_cell_98_16 (.BL(BL16),.BLN(BLN16),.WL(WL98));
sram_cell_6t_5 inst_cell_98_17 (.BL(BL17),.BLN(BLN17),.WL(WL98));
sram_cell_6t_5 inst_cell_98_18 (.BL(BL18),.BLN(BLN18),.WL(WL98));
sram_cell_6t_5 inst_cell_98_19 (.BL(BL19),.BLN(BLN19),.WL(WL98));
sram_cell_6t_5 inst_cell_98_20 (.BL(BL20),.BLN(BLN20),.WL(WL98));
sram_cell_6t_5 inst_cell_98_21 (.BL(BL21),.BLN(BLN21),.WL(WL98));
sram_cell_6t_5 inst_cell_98_22 (.BL(BL22),.BLN(BLN22),.WL(WL98));
sram_cell_6t_5 inst_cell_98_23 (.BL(BL23),.BLN(BLN23),.WL(WL98));
sram_cell_6t_5 inst_cell_98_24 (.BL(BL24),.BLN(BLN24),.WL(WL98));
sram_cell_6t_5 inst_cell_98_25 (.BL(BL25),.BLN(BLN25),.WL(WL98));
sram_cell_6t_5 inst_cell_98_26 (.BL(BL26),.BLN(BLN26),.WL(WL98));
sram_cell_6t_5 inst_cell_98_27 (.BL(BL27),.BLN(BLN27),.WL(WL98));
sram_cell_6t_5 inst_cell_98_28 (.BL(BL28),.BLN(BLN28),.WL(WL98));
sram_cell_6t_5 inst_cell_98_29 (.BL(BL29),.BLN(BLN29),.WL(WL98));
sram_cell_6t_5 inst_cell_98_30 (.BL(BL30),.BLN(BLN30),.WL(WL98));
sram_cell_6t_5 inst_cell_98_31 (.BL(BL31),.BLN(BLN31),.WL(WL98));
sram_cell_6t_5 inst_cell_98_32 (.BL(BL32),.BLN(BLN32),.WL(WL98));
sram_cell_6t_5 inst_cell_98_33 (.BL(BL33),.BLN(BLN33),.WL(WL98));
sram_cell_6t_5 inst_cell_98_34 (.BL(BL34),.BLN(BLN34),.WL(WL98));
sram_cell_6t_5 inst_cell_98_35 (.BL(BL35),.BLN(BLN35),.WL(WL98));
sram_cell_6t_5 inst_cell_98_36 (.BL(BL36),.BLN(BLN36),.WL(WL98));
sram_cell_6t_5 inst_cell_98_37 (.BL(BL37),.BLN(BLN37),.WL(WL98));
sram_cell_6t_5 inst_cell_98_38 (.BL(BL38),.BLN(BLN38),.WL(WL98));
sram_cell_6t_5 inst_cell_98_39 (.BL(BL39),.BLN(BLN39),.WL(WL98));
sram_cell_6t_5 inst_cell_98_40 (.BL(BL40),.BLN(BLN40),.WL(WL98));
sram_cell_6t_5 inst_cell_98_41 (.BL(BL41),.BLN(BLN41),.WL(WL98));
sram_cell_6t_5 inst_cell_98_42 (.BL(BL42),.BLN(BLN42),.WL(WL98));
sram_cell_6t_5 inst_cell_98_43 (.BL(BL43),.BLN(BLN43),.WL(WL98));
sram_cell_6t_5 inst_cell_98_44 (.BL(BL44),.BLN(BLN44),.WL(WL98));
sram_cell_6t_5 inst_cell_98_45 (.BL(BL45),.BLN(BLN45),.WL(WL98));
sram_cell_6t_5 inst_cell_98_46 (.BL(BL46),.BLN(BLN46),.WL(WL98));
sram_cell_6t_5 inst_cell_98_47 (.BL(BL47),.BLN(BLN47),.WL(WL98));
sram_cell_6t_5 inst_cell_98_48 (.BL(BL48),.BLN(BLN48),.WL(WL98));
sram_cell_6t_5 inst_cell_98_49 (.BL(BL49),.BLN(BLN49),.WL(WL98));
sram_cell_6t_5 inst_cell_98_50 (.BL(BL50),.BLN(BLN50),.WL(WL98));
sram_cell_6t_5 inst_cell_98_51 (.BL(BL51),.BLN(BLN51),.WL(WL98));
sram_cell_6t_5 inst_cell_98_52 (.BL(BL52),.BLN(BLN52),.WL(WL98));
sram_cell_6t_5 inst_cell_98_53 (.BL(BL53),.BLN(BLN53),.WL(WL98));
sram_cell_6t_5 inst_cell_98_54 (.BL(BL54),.BLN(BLN54),.WL(WL98));
sram_cell_6t_5 inst_cell_98_55 (.BL(BL55),.BLN(BLN55),.WL(WL98));
sram_cell_6t_5 inst_cell_98_56 (.BL(BL56),.BLN(BLN56),.WL(WL98));
sram_cell_6t_5 inst_cell_98_57 (.BL(BL57),.BLN(BLN57),.WL(WL98));
sram_cell_6t_5 inst_cell_98_58 (.BL(BL58),.BLN(BLN58),.WL(WL98));
sram_cell_6t_5 inst_cell_98_59 (.BL(BL59),.BLN(BLN59),.WL(WL98));
sram_cell_6t_5 inst_cell_98_60 (.BL(BL60),.BLN(BLN60),.WL(WL98));
sram_cell_6t_5 inst_cell_98_61 (.BL(BL61),.BLN(BLN61),.WL(WL98));
sram_cell_6t_5 inst_cell_98_62 (.BL(BL62),.BLN(BLN62),.WL(WL98));
sram_cell_6t_5 inst_cell_98_63 (.BL(BL63),.BLN(BLN63),.WL(WL98));
sram_cell_6t_5 inst_cell_98_64 (.BL(BL64),.BLN(BLN64),.WL(WL98));
sram_cell_6t_5 inst_cell_98_65 (.BL(BL65),.BLN(BLN65),.WL(WL98));
sram_cell_6t_5 inst_cell_98_66 (.BL(BL66),.BLN(BLN66),.WL(WL98));
sram_cell_6t_5 inst_cell_98_67 (.BL(BL67),.BLN(BLN67),.WL(WL98));
sram_cell_6t_5 inst_cell_98_68 (.BL(BL68),.BLN(BLN68),.WL(WL98));
sram_cell_6t_5 inst_cell_98_69 (.BL(BL69),.BLN(BLN69),.WL(WL98));
sram_cell_6t_5 inst_cell_98_70 (.BL(BL70),.BLN(BLN70),.WL(WL98));
sram_cell_6t_5 inst_cell_98_71 (.BL(BL71),.BLN(BLN71),.WL(WL98));
sram_cell_6t_5 inst_cell_98_72 (.BL(BL72),.BLN(BLN72),.WL(WL98));
sram_cell_6t_5 inst_cell_98_73 (.BL(BL73),.BLN(BLN73),.WL(WL98));
sram_cell_6t_5 inst_cell_98_74 (.BL(BL74),.BLN(BLN74),.WL(WL98));
sram_cell_6t_5 inst_cell_98_75 (.BL(BL75),.BLN(BLN75),.WL(WL98));
sram_cell_6t_5 inst_cell_98_76 (.BL(BL76),.BLN(BLN76),.WL(WL98));
sram_cell_6t_5 inst_cell_98_77 (.BL(BL77),.BLN(BLN77),.WL(WL98));
sram_cell_6t_5 inst_cell_98_78 (.BL(BL78),.BLN(BLN78),.WL(WL98));
sram_cell_6t_5 inst_cell_98_79 (.BL(BL79),.BLN(BLN79),.WL(WL98));
sram_cell_6t_5 inst_cell_98_80 (.BL(BL80),.BLN(BLN80),.WL(WL98));
sram_cell_6t_5 inst_cell_98_81 (.BL(BL81),.BLN(BLN81),.WL(WL98));
sram_cell_6t_5 inst_cell_98_82 (.BL(BL82),.BLN(BLN82),.WL(WL98));
sram_cell_6t_5 inst_cell_98_83 (.BL(BL83),.BLN(BLN83),.WL(WL98));
sram_cell_6t_5 inst_cell_98_84 (.BL(BL84),.BLN(BLN84),.WL(WL98));
sram_cell_6t_5 inst_cell_98_85 (.BL(BL85),.BLN(BLN85),.WL(WL98));
sram_cell_6t_5 inst_cell_98_86 (.BL(BL86),.BLN(BLN86),.WL(WL98));
sram_cell_6t_5 inst_cell_98_87 (.BL(BL87),.BLN(BLN87),.WL(WL98));
sram_cell_6t_5 inst_cell_98_88 (.BL(BL88),.BLN(BLN88),.WL(WL98));
sram_cell_6t_5 inst_cell_98_89 (.BL(BL89),.BLN(BLN89),.WL(WL98));
sram_cell_6t_5 inst_cell_98_90 (.BL(BL90),.BLN(BLN90),.WL(WL98));
sram_cell_6t_5 inst_cell_98_91 (.BL(BL91),.BLN(BLN91),.WL(WL98));
sram_cell_6t_5 inst_cell_98_92 (.BL(BL92),.BLN(BLN92),.WL(WL98));
sram_cell_6t_5 inst_cell_98_93 (.BL(BL93),.BLN(BLN93),.WL(WL98));
sram_cell_6t_5 inst_cell_98_94 (.BL(BL94),.BLN(BLN94),.WL(WL98));
sram_cell_6t_5 inst_cell_98_95 (.BL(BL95),.BLN(BLN95),.WL(WL98));
sram_cell_6t_5 inst_cell_98_96 (.BL(BL96),.BLN(BLN96),.WL(WL98));
sram_cell_6t_5 inst_cell_98_97 (.BL(BL97),.BLN(BLN97),.WL(WL98));
sram_cell_6t_5 inst_cell_98_98 (.BL(BL98),.BLN(BLN98),.WL(WL98));
sram_cell_6t_5 inst_cell_98_99 (.BL(BL99),.BLN(BLN99),.WL(WL98));
sram_cell_6t_5 inst_cell_98_100 (.BL(BL100),.BLN(BLN100),.WL(WL98));
sram_cell_6t_5 inst_cell_98_101 (.BL(BL101),.BLN(BLN101),.WL(WL98));
sram_cell_6t_5 inst_cell_98_102 (.BL(BL102),.BLN(BLN102),.WL(WL98));
sram_cell_6t_5 inst_cell_98_103 (.BL(BL103),.BLN(BLN103),.WL(WL98));
sram_cell_6t_5 inst_cell_98_104 (.BL(BL104),.BLN(BLN104),.WL(WL98));
sram_cell_6t_5 inst_cell_98_105 (.BL(BL105),.BLN(BLN105),.WL(WL98));
sram_cell_6t_5 inst_cell_98_106 (.BL(BL106),.BLN(BLN106),.WL(WL98));
sram_cell_6t_5 inst_cell_98_107 (.BL(BL107),.BLN(BLN107),.WL(WL98));
sram_cell_6t_5 inst_cell_98_108 (.BL(BL108),.BLN(BLN108),.WL(WL98));
sram_cell_6t_5 inst_cell_98_109 (.BL(BL109),.BLN(BLN109),.WL(WL98));
sram_cell_6t_5 inst_cell_98_110 (.BL(BL110),.BLN(BLN110),.WL(WL98));
sram_cell_6t_5 inst_cell_98_111 (.BL(BL111),.BLN(BLN111),.WL(WL98));
sram_cell_6t_5 inst_cell_98_112 (.BL(BL112),.BLN(BLN112),.WL(WL98));
sram_cell_6t_5 inst_cell_98_113 (.BL(BL113),.BLN(BLN113),.WL(WL98));
sram_cell_6t_5 inst_cell_98_114 (.BL(BL114),.BLN(BLN114),.WL(WL98));
sram_cell_6t_5 inst_cell_98_115 (.BL(BL115),.BLN(BLN115),.WL(WL98));
sram_cell_6t_5 inst_cell_98_116 (.BL(BL116),.BLN(BLN116),.WL(WL98));
sram_cell_6t_5 inst_cell_98_117 (.BL(BL117),.BLN(BLN117),.WL(WL98));
sram_cell_6t_5 inst_cell_98_118 (.BL(BL118),.BLN(BLN118),.WL(WL98));
sram_cell_6t_5 inst_cell_98_119 (.BL(BL119),.BLN(BLN119),.WL(WL98));
sram_cell_6t_5 inst_cell_98_120 (.BL(BL120),.BLN(BLN120),.WL(WL98));
sram_cell_6t_5 inst_cell_98_121 (.BL(BL121),.BLN(BLN121),.WL(WL98));
sram_cell_6t_5 inst_cell_98_122 (.BL(BL122),.BLN(BLN122),.WL(WL98));
sram_cell_6t_5 inst_cell_98_123 (.BL(BL123),.BLN(BLN123),.WL(WL98));
sram_cell_6t_5 inst_cell_98_124 (.BL(BL124),.BLN(BLN124),.WL(WL98));
sram_cell_6t_5 inst_cell_98_125 (.BL(BL125),.BLN(BLN125),.WL(WL98));
sram_cell_6t_5 inst_cell_98_126 (.BL(BL126),.BLN(BLN126),.WL(WL98));
sram_cell_6t_5 inst_cell_98_127 (.BL(BL127),.BLN(BLN127),.WL(WL98));
sram_cell_6t_5 inst_cell_99_0 (.BL(BL0),.BLN(BLN0),.WL(WL99));
sram_cell_6t_5 inst_cell_99_1 (.BL(BL1),.BLN(BLN1),.WL(WL99));
sram_cell_6t_5 inst_cell_99_2 (.BL(BL2),.BLN(BLN2),.WL(WL99));
sram_cell_6t_5 inst_cell_99_3 (.BL(BL3),.BLN(BLN3),.WL(WL99));
sram_cell_6t_5 inst_cell_99_4 (.BL(BL4),.BLN(BLN4),.WL(WL99));
sram_cell_6t_5 inst_cell_99_5 (.BL(BL5),.BLN(BLN5),.WL(WL99));
sram_cell_6t_5 inst_cell_99_6 (.BL(BL6),.BLN(BLN6),.WL(WL99));
sram_cell_6t_5 inst_cell_99_7 (.BL(BL7),.BLN(BLN7),.WL(WL99));
sram_cell_6t_5 inst_cell_99_8 (.BL(BL8),.BLN(BLN8),.WL(WL99));
sram_cell_6t_5 inst_cell_99_9 (.BL(BL9),.BLN(BLN9),.WL(WL99));
sram_cell_6t_5 inst_cell_99_10 (.BL(BL10),.BLN(BLN10),.WL(WL99));
sram_cell_6t_5 inst_cell_99_11 (.BL(BL11),.BLN(BLN11),.WL(WL99));
sram_cell_6t_5 inst_cell_99_12 (.BL(BL12),.BLN(BLN12),.WL(WL99));
sram_cell_6t_5 inst_cell_99_13 (.BL(BL13),.BLN(BLN13),.WL(WL99));
sram_cell_6t_5 inst_cell_99_14 (.BL(BL14),.BLN(BLN14),.WL(WL99));
sram_cell_6t_5 inst_cell_99_15 (.BL(BL15),.BLN(BLN15),.WL(WL99));
sram_cell_6t_5 inst_cell_99_16 (.BL(BL16),.BLN(BLN16),.WL(WL99));
sram_cell_6t_5 inst_cell_99_17 (.BL(BL17),.BLN(BLN17),.WL(WL99));
sram_cell_6t_5 inst_cell_99_18 (.BL(BL18),.BLN(BLN18),.WL(WL99));
sram_cell_6t_5 inst_cell_99_19 (.BL(BL19),.BLN(BLN19),.WL(WL99));
sram_cell_6t_5 inst_cell_99_20 (.BL(BL20),.BLN(BLN20),.WL(WL99));
sram_cell_6t_5 inst_cell_99_21 (.BL(BL21),.BLN(BLN21),.WL(WL99));
sram_cell_6t_5 inst_cell_99_22 (.BL(BL22),.BLN(BLN22),.WL(WL99));
sram_cell_6t_5 inst_cell_99_23 (.BL(BL23),.BLN(BLN23),.WL(WL99));
sram_cell_6t_5 inst_cell_99_24 (.BL(BL24),.BLN(BLN24),.WL(WL99));
sram_cell_6t_5 inst_cell_99_25 (.BL(BL25),.BLN(BLN25),.WL(WL99));
sram_cell_6t_5 inst_cell_99_26 (.BL(BL26),.BLN(BLN26),.WL(WL99));
sram_cell_6t_5 inst_cell_99_27 (.BL(BL27),.BLN(BLN27),.WL(WL99));
sram_cell_6t_5 inst_cell_99_28 (.BL(BL28),.BLN(BLN28),.WL(WL99));
sram_cell_6t_5 inst_cell_99_29 (.BL(BL29),.BLN(BLN29),.WL(WL99));
sram_cell_6t_5 inst_cell_99_30 (.BL(BL30),.BLN(BLN30),.WL(WL99));
sram_cell_6t_5 inst_cell_99_31 (.BL(BL31),.BLN(BLN31),.WL(WL99));
sram_cell_6t_5 inst_cell_99_32 (.BL(BL32),.BLN(BLN32),.WL(WL99));
sram_cell_6t_5 inst_cell_99_33 (.BL(BL33),.BLN(BLN33),.WL(WL99));
sram_cell_6t_5 inst_cell_99_34 (.BL(BL34),.BLN(BLN34),.WL(WL99));
sram_cell_6t_5 inst_cell_99_35 (.BL(BL35),.BLN(BLN35),.WL(WL99));
sram_cell_6t_5 inst_cell_99_36 (.BL(BL36),.BLN(BLN36),.WL(WL99));
sram_cell_6t_5 inst_cell_99_37 (.BL(BL37),.BLN(BLN37),.WL(WL99));
sram_cell_6t_5 inst_cell_99_38 (.BL(BL38),.BLN(BLN38),.WL(WL99));
sram_cell_6t_5 inst_cell_99_39 (.BL(BL39),.BLN(BLN39),.WL(WL99));
sram_cell_6t_5 inst_cell_99_40 (.BL(BL40),.BLN(BLN40),.WL(WL99));
sram_cell_6t_5 inst_cell_99_41 (.BL(BL41),.BLN(BLN41),.WL(WL99));
sram_cell_6t_5 inst_cell_99_42 (.BL(BL42),.BLN(BLN42),.WL(WL99));
sram_cell_6t_5 inst_cell_99_43 (.BL(BL43),.BLN(BLN43),.WL(WL99));
sram_cell_6t_5 inst_cell_99_44 (.BL(BL44),.BLN(BLN44),.WL(WL99));
sram_cell_6t_5 inst_cell_99_45 (.BL(BL45),.BLN(BLN45),.WL(WL99));
sram_cell_6t_5 inst_cell_99_46 (.BL(BL46),.BLN(BLN46),.WL(WL99));
sram_cell_6t_5 inst_cell_99_47 (.BL(BL47),.BLN(BLN47),.WL(WL99));
sram_cell_6t_5 inst_cell_99_48 (.BL(BL48),.BLN(BLN48),.WL(WL99));
sram_cell_6t_5 inst_cell_99_49 (.BL(BL49),.BLN(BLN49),.WL(WL99));
sram_cell_6t_5 inst_cell_99_50 (.BL(BL50),.BLN(BLN50),.WL(WL99));
sram_cell_6t_5 inst_cell_99_51 (.BL(BL51),.BLN(BLN51),.WL(WL99));
sram_cell_6t_5 inst_cell_99_52 (.BL(BL52),.BLN(BLN52),.WL(WL99));
sram_cell_6t_5 inst_cell_99_53 (.BL(BL53),.BLN(BLN53),.WL(WL99));
sram_cell_6t_5 inst_cell_99_54 (.BL(BL54),.BLN(BLN54),.WL(WL99));
sram_cell_6t_5 inst_cell_99_55 (.BL(BL55),.BLN(BLN55),.WL(WL99));
sram_cell_6t_5 inst_cell_99_56 (.BL(BL56),.BLN(BLN56),.WL(WL99));
sram_cell_6t_5 inst_cell_99_57 (.BL(BL57),.BLN(BLN57),.WL(WL99));
sram_cell_6t_5 inst_cell_99_58 (.BL(BL58),.BLN(BLN58),.WL(WL99));
sram_cell_6t_5 inst_cell_99_59 (.BL(BL59),.BLN(BLN59),.WL(WL99));
sram_cell_6t_5 inst_cell_99_60 (.BL(BL60),.BLN(BLN60),.WL(WL99));
sram_cell_6t_5 inst_cell_99_61 (.BL(BL61),.BLN(BLN61),.WL(WL99));
sram_cell_6t_5 inst_cell_99_62 (.BL(BL62),.BLN(BLN62),.WL(WL99));
sram_cell_6t_5 inst_cell_99_63 (.BL(BL63),.BLN(BLN63),.WL(WL99));
sram_cell_6t_5 inst_cell_99_64 (.BL(BL64),.BLN(BLN64),.WL(WL99));
sram_cell_6t_5 inst_cell_99_65 (.BL(BL65),.BLN(BLN65),.WL(WL99));
sram_cell_6t_5 inst_cell_99_66 (.BL(BL66),.BLN(BLN66),.WL(WL99));
sram_cell_6t_5 inst_cell_99_67 (.BL(BL67),.BLN(BLN67),.WL(WL99));
sram_cell_6t_5 inst_cell_99_68 (.BL(BL68),.BLN(BLN68),.WL(WL99));
sram_cell_6t_5 inst_cell_99_69 (.BL(BL69),.BLN(BLN69),.WL(WL99));
sram_cell_6t_5 inst_cell_99_70 (.BL(BL70),.BLN(BLN70),.WL(WL99));
sram_cell_6t_5 inst_cell_99_71 (.BL(BL71),.BLN(BLN71),.WL(WL99));
sram_cell_6t_5 inst_cell_99_72 (.BL(BL72),.BLN(BLN72),.WL(WL99));
sram_cell_6t_5 inst_cell_99_73 (.BL(BL73),.BLN(BLN73),.WL(WL99));
sram_cell_6t_5 inst_cell_99_74 (.BL(BL74),.BLN(BLN74),.WL(WL99));
sram_cell_6t_5 inst_cell_99_75 (.BL(BL75),.BLN(BLN75),.WL(WL99));
sram_cell_6t_5 inst_cell_99_76 (.BL(BL76),.BLN(BLN76),.WL(WL99));
sram_cell_6t_5 inst_cell_99_77 (.BL(BL77),.BLN(BLN77),.WL(WL99));
sram_cell_6t_5 inst_cell_99_78 (.BL(BL78),.BLN(BLN78),.WL(WL99));
sram_cell_6t_5 inst_cell_99_79 (.BL(BL79),.BLN(BLN79),.WL(WL99));
sram_cell_6t_5 inst_cell_99_80 (.BL(BL80),.BLN(BLN80),.WL(WL99));
sram_cell_6t_5 inst_cell_99_81 (.BL(BL81),.BLN(BLN81),.WL(WL99));
sram_cell_6t_5 inst_cell_99_82 (.BL(BL82),.BLN(BLN82),.WL(WL99));
sram_cell_6t_5 inst_cell_99_83 (.BL(BL83),.BLN(BLN83),.WL(WL99));
sram_cell_6t_5 inst_cell_99_84 (.BL(BL84),.BLN(BLN84),.WL(WL99));
sram_cell_6t_5 inst_cell_99_85 (.BL(BL85),.BLN(BLN85),.WL(WL99));
sram_cell_6t_5 inst_cell_99_86 (.BL(BL86),.BLN(BLN86),.WL(WL99));
sram_cell_6t_5 inst_cell_99_87 (.BL(BL87),.BLN(BLN87),.WL(WL99));
sram_cell_6t_5 inst_cell_99_88 (.BL(BL88),.BLN(BLN88),.WL(WL99));
sram_cell_6t_5 inst_cell_99_89 (.BL(BL89),.BLN(BLN89),.WL(WL99));
sram_cell_6t_5 inst_cell_99_90 (.BL(BL90),.BLN(BLN90),.WL(WL99));
sram_cell_6t_5 inst_cell_99_91 (.BL(BL91),.BLN(BLN91),.WL(WL99));
sram_cell_6t_5 inst_cell_99_92 (.BL(BL92),.BLN(BLN92),.WL(WL99));
sram_cell_6t_5 inst_cell_99_93 (.BL(BL93),.BLN(BLN93),.WL(WL99));
sram_cell_6t_5 inst_cell_99_94 (.BL(BL94),.BLN(BLN94),.WL(WL99));
sram_cell_6t_5 inst_cell_99_95 (.BL(BL95),.BLN(BLN95),.WL(WL99));
sram_cell_6t_5 inst_cell_99_96 (.BL(BL96),.BLN(BLN96),.WL(WL99));
sram_cell_6t_5 inst_cell_99_97 (.BL(BL97),.BLN(BLN97),.WL(WL99));
sram_cell_6t_5 inst_cell_99_98 (.BL(BL98),.BLN(BLN98),.WL(WL99));
sram_cell_6t_5 inst_cell_99_99 (.BL(BL99),.BLN(BLN99),.WL(WL99));
sram_cell_6t_5 inst_cell_99_100 (.BL(BL100),.BLN(BLN100),.WL(WL99));
sram_cell_6t_5 inst_cell_99_101 (.BL(BL101),.BLN(BLN101),.WL(WL99));
sram_cell_6t_5 inst_cell_99_102 (.BL(BL102),.BLN(BLN102),.WL(WL99));
sram_cell_6t_5 inst_cell_99_103 (.BL(BL103),.BLN(BLN103),.WL(WL99));
sram_cell_6t_5 inst_cell_99_104 (.BL(BL104),.BLN(BLN104),.WL(WL99));
sram_cell_6t_5 inst_cell_99_105 (.BL(BL105),.BLN(BLN105),.WL(WL99));
sram_cell_6t_5 inst_cell_99_106 (.BL(BL106),.BLN(BLN106),.WL(WL99));
sram_cell_6t_5 inst_cell_99_107 (.BL(BL107),.BLN(BLN107),.WL(WL99));
sram_cell_6t_5 inst_cell_99_108 (.BL(BL108),.BLN(BLN108),.WL(WL99));
sram_cell_6t_5 inst_cell_99_109 (.BL(BL109),.BLN(BLN109),.WL(WL99));
sram_cell_6t_5 inst_cell_99_110 (.BL(BL110),.BLN(BLN110),.WL(WL99));
sram_cell_6t_5 inst_cell_99_111 (.BL(BL111),.BLN(BLN111),.WL(WL99));
sram_cell_6t_5 inst_cell_99_112 (.BL(BL112),.BLN(BLN112),.WL(WL99));
sram_cell_6t_5 inst_cell_99_113 (.BL(BL113),.BLN(BLN113),.WL(WL99));
sram_cell_6t_5 inst_cell_99_114 (.BL(BL114),.BLN(BLN114),.WL(WL99));
sram_cell_6t_5 inst_cell_99_115 (.BL(BL115),.BLN(BLN115),.WL(WL99));
sram_cell_6t_5 inst_cell_99_116 (.BL(BL116),.BLN(BLN116),.WL(WL99));
sram_cell_6t_5 inst_cell_99_117 (.BL(BL117),.BLN(BLN117),.WL(WL99));
sram_cell_6t_5 inst_cell_99_118 (.BL(BL118),.BLN(BLN118),.WL(WL99));
sram_cell_6t_5 inst_cell_99_119 (.BL(BL119),.BLN(BLN119),.WL(WL99));
sram_cell_6t_5 inst_cell_99_120 (.BL(BL120),.BLN(BLN120),.WL(WL99));
sram_cell_6t_5 inst_cell_99_121 (.BL(BL121),.BLN(BLN121),.WL(WL99));
sram_cell_6t_5 inst_cell_99_122 (.BL(BL122),.BLN(BLN122),.WL(WL99));
sram_cell_6t_5 inst_cell_99_123 (.BL(BL123),.BLN(BLN123),.WL(WL99));
sram_cell_6t_5 inst_cell_99_124 (.BL(BL124),.BLN(BLN124),.WL(WL99));
sram_cell_6t_5 inst_cell_99_125 (.BL(BL125),.BLN(BLN125),.WL(WL99));
sram_cell_6t_5 inst_cell_99_126 (.BL(BL126),.BLN(BLN126),.WL(WL99));
sram_cell_6t_5 inst_cell_99_127 (.BL(BL127),.BLN(BLN127),.WL(WL99));
sram_cell_6t_5 inst_cell_100_0 (.BL(BL0),.BLN(BLN0),.WL(WL100));
sram_cell_6t_5 inst_cell_100_1 (.BL(BL1),.BLN(BLN1),.WL(WL100));
sram_cell_6t_5 inst_cell_100_2 (.BL(BL2),.BLN(BLN2),.WL(WL100));
sram_cell_6t_5 inst_cell_100_3 (.BL(BL3),.BLN(BLN3),.WL(WL100));
sram_cell_6t_5 inst_cell_100_4 (.BL(BL4),.BLN(BLN4),.WL(WL100));
sram_cell_6t_5 inst_cell_100_5 (.BL(BL5),.BLN(BLN5),.WL(WL100));
sram_cell_6t_5 inst_cell_100_6 (.BL(BL6),.BLN(BLN6),.WL(WL100));
sram_cell_6t_5 inst_cell_100_7 (.BL(BL7),.BLN(BLN7),.WL(WL100));
sram_cell_6t_5 inst_cell_100_8 (.BL(BL8),.BLN(BLN8),.WL(WL100));
sram_cell_6t_5 inst_cell_100_9 (.BL(BL9),.BLN(BLN9),.WL(WL100));
sram_cell_6t_5 inst_cell_100_10 (.BL(BL10),.BLN(BLN10),.WL(WL100));
sram_cell_6t_5 inst_cell_100_11 (.BL(BL11),.BLN(BLN11),.WL(WL100));
sram_cell_6t_5 inst_cell_100_12 (.BL(BL12),.BLN(BLN12),.WL(WL100));
sram_cell_6t_5 inst_cell_100_13 (.BL(BL13),.BLN(BLN13),.WL(WL100));
sram_cell_6t_5 inst_cell_100_14 (.BL(BL14),.BLN(BLN14),.WL(WL100));
sram_cell_6t_5 inst_cell_100_15 (.BL(BL15),.BLN(BLN15),.WL(WL100));
sram_cell_6t_5 inst_cell_100_16 (.BL(BL16),.BLN(BLN16),.WL(WL100));
sram_cell_6t_5 inst_cell_100_17 (.BL(BL17),.BLN(BLN17),.WL(WL100));
sram_cell_6t_5 inst_cell_100_18 (.BL(BL18),.BLN(BLN18),.WL(WL100));
sram_cell_6t_5 inst_cell_100_19 (.BL(BL19),.BLN(BLN19),.WL(WL100));
sram_cell_6t_5 inst_cell_100_20 (.BL(BL20),.BLN(BLN20),.WL(WL100));
sram_cell_6t_5 inst_cell_100_21 (.BL(BL21),.BLN(BLN21),.WL(WL100));
sram_cell_6t_5 inst_cell_100_22 (.BL(BL22),.BLN(BLN22),.WL(WL100));
sram_cell_6t_5 inst_cell_100_23 (.BL(BL23),.BLN(BLN23),.WL(WL100));
sram_cell_6t_5 inst_cell_100_24 (.BL(BL24),.BLN(BLN24),.WL(WL100));
sram_cell_6t_5 inst_cell_100_25 (.BL(BL25),.BLN(BLN25),.WL(WL100));
sram_cell_6t_5 inst_cell_100_26 (.BL(BL26),.BLN(BLN26),.WL(WL100));
sram_cell_6t_5 inst_cell_100_27 (.BL(BL27),.BLN(BLN27),.WL(WL100));
sram_cell_6t_5 inst_cell_100_28 (.BL(BL28),.BLN(BLN28),.WL(WL100));
sram_cell_6t_5 inst_cell_100_29 (.BL(BL29),.BLN(BLN29),.WL(WL100));
sram_cell_6t_5 inst_cell_100_30 (.BL(BL30),.BLN(BLN30),.WL(WL100));
sram_cell_6t_5 inst_cell_100_31 (.BL(BL31),.BLN(BLN31),.WL(WL100));
sram_cell_6t_5 inst_cell_100_32 (.BL(BL32),.BLN(BLN32),.WL(WL100));
sram_cell_6t_5 inst_cell_100_33 (.BL(BL33),.BLN(BLN33),.WL(WL100));
sram_cell_6t_5 inst_cell_100_34 (.BL(BL34),.BLN(BLN34),.WL(WL100));
sram_cell_6t_5 inst_cell_100_35 (.BL(BL35),.BLN(BLN35),.WL(WL100));
sram_cell_6t_5 inst_cell_100_36 (.BL(BL36),.BLN(BLN36),.WL(WL100));
sram_cell_6t_5 inst_cell_100_37 (.BL(BL37),.BLN(BLN37),.WL(WL100));
sram_cell_6t_5 inst_cell_100_38 (.BL(BL38),.BLN(BLN38),.WL(WL100));
sram_cell_6t_5 inst_cell_100_39 (.BL(BL39),.BLN(BLN39),.WL(WL100));
sram_cell_6t_5 inst_cell_100_40 (.BL(BL40),.BLN(BLN40),.WL(WL100));
sram_cell_6t_5 inst_cell_100_41 (.BL(BL41),.BLN(BLN41),.WL(WL100));
sram_cell_6t_5 inst_cell_100_42 (.BL(BL42),.BLN(BLN42),.WL(WL100));
sram_cell_6t_5 inst_cell_100_43 (.BL(BL43),.BLN(BLN43),.WL(WL100));
sram_cell_6t_5 inst_cell_100_44 (.BL(BL44),.BLN(BLN44),.WL(WL100));
sram_cell_6t_5 inst_cell_100_45 (.BL(BL45),.BLN(BLN45),.WL(WL100));
sram_cell_6t_5 inst_cell_100_46 (.BL(BL46),.BLN(BLN46),.WL(WL100));
sram_cell_6t_5 inst_cell_100_47 (.BL(BL47),.BLN(BLN47),.WL(WL100));
sram_cell_6t_5 inst_cell_100_48 (.BL(BL48),.BLN(BLN48),.WL(WL100));
sram_cell_6t_5 inst_cell_100_49 (.BL(BL49),.BLN(BLN49),.WL(WL100));
sram_cell_6t_5 inst_cell_100_50 (.BL(BL50),.BLN(BLN50),.WL(WL100));
sram_cell_6t_5 inst_cell_100_51 (.BL(BL51),.BLN(BLN51),.WL(WL100));
sram_cell_6t_5 inst_cell_100_52 (.BL(BL52),.BLN(BLN52),.WL(WL100));
sram_cell_6t_5 inst_cell_100_53 (.BL(BL53),.BLN(BLN53),.WL(WL100));
sram_cell_6t_5 inst_cell_100_54 (.BL(BL54),.BLN(BLN54),.WL(WL100));
sram_cell_6t_5 inst_cell_100_55 (.BL(BL55),.BLN(BLN55),.WL(WL100));
sram_cell_6t_5 inst_cell_100_56 (.BL(BL56),.BLN(BLN56),.WL(WL100));
sram_cell_6t_5 inst_cell_100_57 (.BL(BL57),.BLN(BLN57),.WL(WL100));
sram_cell_6t_5 inst_cell_100_58 (.BL(BL58),.BLN(BLN58),.WL(WL100));
sram_cell_6t_5 inst_cell_100_59 (.BL(BL59),.BLN(BLN59),.WL(WL100));
sram_cell_6t_5 inst_cell_100_60 (.BL(BL60),.BLN(BLN60),.WL(WL100));
sram_cell_6t_5 inst_cell_100_61 (.BL(BL61),.BLN(BLN61),.WL(WL100));
sram_cell_6t_5 inst_cell_100_62 (.BL(BL62),.BLN(BLN62),.WL(WL100));
sram_cell_6t_5 inst_cell_100_63 (.BL(BL63),.BLN(BLN63),.WL(WL100));
sram_cell_6t_5 inst_cell_100_64 (.BL(BL64),.BLN(BLN64),.WL(WL100));
sram_cell_6t_5 inst_cell_100_65 (.BL(BL65),.BLN(BLN65),.WL(WL100));
sram_cell_6t_5 inst_cell_100_66 (.BL(BL66),.BLN(BLN66),.WL(WL100));
sram_cell_6t_5 inst_cell_100_67 (.BL(BL67),.BLN(BLN67),.WL(WL100));
sram_cell_6t_5 inst_cell_100_68 (.BL(BL68),.BLN(BLN68),.WL(WL100));
sram_cell_6t_5 inst_cell_100_69 (.BL(BL69),.BLN(BLN69),.WL(WL100));
sram_cell_6t_5 inst_cell_100_70 (.BL(BL70),.BLN(BLN70),.WL(WL100));
sram_cell_6t_5 inst_cell_100_71 (.BL(BL71),.BLN(BLN71),.WL(WL100));
sram_cell_6t_5 inst_cell_100_72 (.BL(BL72),.BLN(BLN72),.WL(WL100));
sram_cell_6t_5 inst_cell_100_73 (.BL(BL73),.BLN(BLN73),.WL(WL100));
sram_cell_6t_5 inst_cell_100_74 (.BL(BL74),.BLN(BLN74),.WL(WL100));
sram_cell_6t_5 inst_cell_100_75 (.BL(BL75),.BLN(BLN75),.WL(WL100));
sram_cell_6t_5 inst_cell_100_76 (.BL(BL76),.BLN(BLN76),.WL(WL100));
sram_cell_6t_5 inst_cell_100_77 (.BL(BL77),.BLN(BLN77),.WL(WL100));
sram_cell_6t_5 inst_cell_100_78 (.BL(BL78),.BLN(BLN78),.WL(WL100));
sram_cell_6t_5 inst_cell_100_79 (.BL(BL79),.BLN(BLN79),.WL(WL100));
sram_cell_6t_5 inst_cell_100_80 (.BL(BL80),.BLN(BLN80),.WL(WL100));
sram_cell_6t_5 inst_cell_100_81 (.BL(BL81),.BLN(BLN81),.WL(WL100));
sram_cell_6t_5 inst_cell_100_82 (.BL(BL82),.BLN(BLN82),.WL(WL100));
sram_cell_6t_5 inst_cell_100_83 (.BL(BL83),.BLN(BLN83),.WL(WL100));
sram_cell_6t_5 inst_cell_100_84 (.BL(BL84),.BLN(BLN84),.WL(WL100));
sram_cell_6t_5 inst_cell_100_85 (.BL(BL85),.BLN(BLN85),.WL(WL100));
sram_cell_6t_5 inst_cell_100_86 (.BL(BL86),.BLN(BLN86),.WL(WL100));
sram_cell_6t_5 inst_cell_100_87 (.BL(BL87),.BLN(BLN87),.WL(WL100));
sram_cell_6t_5 inst_cell_100_88 (.BL(BL88),.BLN(BLN88),.WL(WL100));
sram_cell_6t_5 inst_cell_100_89 (.BL(BL89),.BLN(BLN89),.WL(WL100));
sram_cell_6t_5 inst_cell_100_90 (.BL(BL90),.BLN(BLN90),.WL(WL100));
sram_cell_6t_5 inst_cell_100_91 (.BL(BL91),.BLN(BLN91),.WL(WL100));
sram_cell_6t_5 inst_cell_100_92 (.BL(BL92),.BLN(BLN92),.WL(WL100));
sram_cell_6t_5 inst_cell_100_93 (.BL(BL93),.BLN(BLN93),.WL(WL100));
sram_cell_6t_5 inst_cell_100_94 (.BL(BL94),.BLN(BLN94),.WL(WL100));
sram_cell_6t_5 inst_cell_100_95 (.BL(BL95),.BLN(BLN95),.WL(WL100));
sram_cell_6t_5 inst_cell_100_96 (.BL(BL96),.BLN(BLN96),.WL(WL100));
sram_cell_6t_5 inst_cell_100_97 (.BL(BL97),.BLN(BLN97),.WL(WL100));
sram_cell_6t_5 inst_cell_100_98 (.BL(BL98),.BLN(BLN98),.WL(WL100));
sram_cell_6t_5 inst_cell_100_99 (.BL(BL99),.BLN(BLN99),.WL(WL100));
sram_cell_6t_5 inst_cell_100_100 (.BL(BL100),.BLN(BLN100),.WL(WL100));
sram_cell_6t_5 inst_cell_100_101 (.BL(BL101),.BLN(BLN101),.WL(WL100));
sram_cell_6t_5 inst_cell_100_102 (.BL(BL102),.BLN(BLN102),.WL(WL100));
sram_cell_6t_5 inst_cell_100_103 (.BL(BL103),.BLN(BLN103),.WL(WL100));
sram_cell_6t_5 inst_cell_100_104 (.BL(BL104),.BLN(BLN104),.WL(WL100));
sram_cell_6t_5 inst_cell_100_105 (.BL(BL105),.BLN(BLN105),.WL(WL100));
sram_cell_6t_5 inst_cell_100_106 (.BL(BL106),.BLN(BLN106),.WL(WL100));
sram_cell_6t_5 inst_cell_100_107 (.BL(BL107),.BLN(BLN107),.WL(WL100));
sram_cell_6t_5 inst_cell_100_108 (.BL(BL108),.BLN(BLN108),.WL(WL100));
sram_cell_6t_5 inst_cell_100_109 (.BL(BL109),.BLN(BLN109),.WL(WL100));
sram_cell_6t_5 inst_cell_100_110 (.BL(BL110),.BLN(BLN110),.WL(WL100));
sram_cell_6t_5 inst_cell_100_111 (.BL(BL111),.BLN(BLN111),.WL(WL100));
sram_cell_6t_5 inst_cell_100_112 (.BL(BL112),.BLN(BLN112),.WL(WL100));
sram_cell_6t_5 inst_cell_100_113 (.BL(BL113),.BLN(BLN113),.WL(WL100));
sram_cell_6t_5 inst_cell_100_114 (.BL(BL114),.BLN(BLN114),.WL(WL100));
sram_cell_6t_5 inst_cell_100_115 (.BL(BL115),.BLN(BLN115),.WL(WL100));
sram_cell_6t_5 inst_cell_100_116 (.BL(BL116),.BLN(BLN116),.WL(WL100));
sram_cell_6t_5 inst_cell_100_117 (.BL(BL117),.BLN(BLN117),.WL(WL100));
sram_cell_6t_5 inst_cell_100_118 (.BL(BL118),.BLN(BLN118),.WL(WL100));
sram_cell_6t_5 inst_cell_100_119 (.BL(BL119),.BLN(BLN119),.WL(WL100));
sram_cell_6t_5 inst_cell_100_120 (.BL(BL120),.BLN(BLN120),.WL(WL100));
sram_cell_6t_5 inst_cell_100_121 (.BL(BL121),.BLN(BLN121),.WL(WL100));
sram_cell_6t_5 inst_cell_100_122 (.BL(BL122),.BLN(BLN122),.WL(WL100));
sram_cell_6t_5 inst_cell_100_123 (.BL(BL123),.BLN(BLN123),.WL(WL100));
sram_cell_6t_5 inst_cell_100_124 (.BL(BL124),.BLN(BLN124),.WL(WL100));
sram_cell_6t_5 inst_cell_100_125 (.BL(BL125),.BLN(BLN125),.WL(WL100));
sram_cell_6t_5 inst_cell_100_126 (.BL(BL126),.BLN(BLN126),.WL(WL100));
sram_cell_6t_5 inst_cell_100_127 (.BL(BL127),.BLN(BLN127),.WL(WL100));
sram_cell_6t_5 inst_cell_101_0 (.BL(BL0),.BLN(BLN0),.WL(WL101));
sram_cell_6t_5 inst_cell_101_1 (.BL(BL1),.BLN(BLN1),.WL(WL101));
sram_cell_6t_5 inst_cell_101_2 (.BL(BL2),.BLN(BLN2),.WL(WL101));
sram_cell_6t_5 inst_cell_101_3 (.BL(BL3),.BLN(BLN3),.WL(WL101));
sram_cell_6t_5 inst_cell_101_4 (.BL(BL4),.BLN(BLN4),.WL(WL101));
sram_cell_6t_5 inst_cell_101_5 (.BL(BL5),.BLN(BLN5),.WL(WL101));
sram_cell_6t_5 inst_cell_101_6 (.BL(BL6),.BLN(BLN6),.WL(WL101));
sram_cell_6t_5 inst_cell_101_7 (.BL(BL7),.BLN(BLN7),.WL(WL101));
sram_cell_6t_5 inst_cell_101_8 (.BL(BL8),.BLN(BLN8),.WL(WL101));
sram_cell_6t_5 inst_cell_101_9 (.BL(BL9),.BLN(BLN9),.WL(WL101));
sram_cell_6t_5 inst_cell_101_10 (.BL(BL10),.BLN(BLN10),.WL(WL101));
sram_cell_6t_5 inst_cell_101_11 (.BL(BL11),.BLN(BLN11),.WL(WL101));
sram_cell_6t_5 inst_cell_101_12 (.BL(BL12),.BLN(BLN12),.WL(WL101));
sram_cell_6t_5 inst_cell_101_13 (.BL(BL13),.BLN(BLN13),.WL(WL101));
sram_cell_6t_5 inst_cell_101_14 (.BL(BL14),.BLN(BLN14),.WL(WL101));
sram_cell_6t_5 inst_cell_101_15 (.BL(BL15),.BLN(BLN15),.WL(WL101));
sram_cell_6t_5 inst_cell_101_16 (.BL(BL16),.BLN(BLN16),.WL(WL101));
sram_cell_6t_5 inst_cell_101_17 (.BL(BL17),.BLN(BLN17),.WL(WL101));
sram_cell_6t_5 inst_cell_101_18 (.BL(BL18),.BLN(BLN18),.WL(WL101));
sram_cell_6t_5 inst_cell_101_19 (.BL(BL19),.BLN(BLN19),.WL(WL101));
sram_cell_6t_5 inst_cell_101_20 (.BL(BL20),.BLN(BLN20),.WL(WL101));
sram_cell_6t_5 inst_cell_101_21 (.BL(BL21),.BLN(BLN21),.WL(WL101));
sram_cell_6t_5 inst_cell_101_22 (.BL(BL22),.BLN(BLN22),.WL(WL101));
sram_cell_6t_5 inst_cell_101_23 (.BL(BL23),.BLN(BLN23),.WL(WL101));
sram_cell_6t_5 inst_cell_101_24 (.BL(BL24),.BLN(BLN24),.WL(WL101));
sram_cell_6t_5 inst_cell_101_25 (.BL(BL25),.BLN(BLN25),.WL(WL101));
sram_cell_6t_5 inst_cell_101_26 (.BL(BL26),.BLN(BLN26),.WL(WL101));
sram_cell_6t_5 inst_cell_101_27 (.BL(BL27),.BLN(BLN27),.WL(WL101));
sram_cell_6t_5 inst_cell_101_28 (.BL(BL28),.BLN(BLN28),.WL(WL101));
sram_cell_6t_5 inst_cell_101_29 (.BL(BL29),.BLN(BLN29),.WL(WL101));
sram_cell_6t_5 inst_cell_101_30 (.BL(BL30),.BLN(BLN30),.WL(WL101));
sram_cell_6t_5 inst_cell_101_31 (.BL(BL31),.BLN(BLN31),.WL(WL101));
sram_cell_6t_5 inst_cell_101_32 (.BL(BL32),.BLN(BLN32),.WL(WL101));
sram_cell_6t_5 inst_cell_101_33 (.BL(BL33),.BLN(BLN33),.WL(WL101));
sram_cell_6t_5 inst_cell_101_34 (.BL(BL34),.BLN(BLN34),.WL(WL101));
sram_cell_6t_5 inst_cell_101_35 (.BL(BL35),.BLN(BLN35),.WL(WL101));
sram_cell_6t_5 inst_cell_101_36 (.BL(BL36),.BLN(BLN36),.WL(WL101));
sram_cell_6t_5 inst_cell_101_37 (.BL(BL37),.BLN(BLN37),.WL(WL101));
sram_cell_6t_5 inst_cell_101_38 (.BL(BL38),.BLN(BLN38),.WL(WL101));
sram_cell_6t_5 inst_cell_101_39 (.BL(BL39),.BLN(BLN39),.WL(WL101));
sram_cell_6t_5 inst_cell_101_40 (.BL(BL40),.BLN(BLN40),.WL(WL101));
sram_cell_6t_5 inst_cell_101_41 (.BL(BL41),.BLN(BLN41),.WL(WL101));
sram_cell_6t_5 inst_cell_101_42 (.BL(BL42),.BLN(BLN42),.WL(WL101));
sram_cell_6t_5 inst_cell_101_43 (.BL(BL43),.BLN(BLN43),.WL(WL101));
sram_cell_6t_5 inst_cell_101_44 (.BL(BL44),.BLN(BLN44),.WL(WL101));
sram_cell_6t_5 inst_cell_101_45 (.BL(BL45),.BLN(BLN45),.WL(WL101));
sram_cell_6t_5 inst_cell_101_46 (.BL(BL46),.BLN(BLN46),.WL(WL101));
sram_cell_6t_5 inst_cell_101_47 (.BL(BL47),.BLN(BLN47),.WL(WL101));
sram_cell_6t_5 inst_cell_101_48 (.BL(BL48),.BLN(BLN48),.WL(WL101));
sram_cell_6t_5 inst_cell_101_49 (.BL(BL49),.BLN(BLN49),.WL(WL101));
sram_cell_6t_5 inst_cell_101_50 (.BL(BL50),.BLN(BLN50),.WL(WL101));
sram_cell_6t_5 inst_cell_101_51 (.BL(BL51),.BLN(BLN51),.WL(WL101));
sram_cell_6t_5 inst_cell_101_52 (.BL(BL52),.BLN(BLN52),.WL(WL101));
sram_cell_6t_5 inst_cell_101_53 (.BL(BL53),.BLN(BLN53),.WL(WL101));
sram_cell_6t_5 inst_cell_101_54 (.BL(BL54),.BLN(BLN54),.WL(WL101));
sram_cell_6t_5 inst_cell_101_55 (.BL(BL55),.BLN(BLN55),.WL(WL101));
sram_cell_6t_5 inst_cell_101_56 (.BL(BL56),.BLN(BLN56),.WL(WL101));
sram_cell_6t_5 inst_cell_101_57 (.BL(BL57),.BLN(BLN57),.WL(WL101));
sram_cell_6t_5 inst_cell_101_58 (.BL(BL58),.BLN(BLN58),.WL(WL101));
sram_cell_6t_5 inst_cell_101_59 (.BL(BL59),.BLN(BLN59),.WL(WL101));
sram_cell_6t_5 inst_cell_101_60 (.BL(BL60),.BLN(BLN60),.WL(WL101));
sram_cell_6t_5 inst_cell_101_61 (.BL(BL61),.BLN(BLN61),.WL(WL101));
sram_cell_6t_5 inst_cell_101_62 (.BL(BL62),.BLN(BLN62),.WL(WL101));
sram_cell_6t_5 inst_cell_101_63 (.BL(BL63),.BLN(BLN63),.WL(WL101));
sram_cell_6t_5 inst_cell_101_64 (.BL(BL64),.BLN(BLN64),.WL(WL101));
sram_cell_6t_5 inst_cell_101_65 (.BL(BL65),.BLN(BLN65),.WL(WL101));
sram_cell_6t_5 inst_cell_101_66 (.BL(BL66),.BLN(BLN66),.WL(WL101));
sram_cell_6t_5 inst_cell_101_67 (.BL(BL67),.BLN(BLN67),.WL(WL101));
sram_cell_6t_5 inst_cell_101_68 (.BL(BL68),.BLN(BLN68),.WL(WL101));
sram_cell_6t_5 inst_cell_101_69 (.BL(BL69),.BLN(BLN69),.WL(WL101));
sram_cell_6t_5 inst_cell_101_70 (.BL(BL70),.BLN(BLN70),.WL(WL101));
sram_cell_6t_5 inst_cell_101_71 (.BL(BL71),.BLN(BLN71),.WL(WL101));
sram_cell_6t_5 inst_cell_101_72 (.BL(BL72),.BLN(BLN72),.WL(WL101));
sram_cell_6t_5 inst_cell_101_73 (.BL(BL73),.BLN(BLN73),.WL(WL101));
sram_cell_6t_5 inst_cell_101_74 (.BL(BL74),.BLN(BLN74),.WL(WL101));
sram_cell_6t_5 inst_cell_101_75 (.BL(BL75),.BLN(BLN75),.WL(WL101));
sram_cell_6t_5 inst_cell_101_76 (.BL(BL76),.BLN(BLN76),.WL(WL101));
sram_cell_6t_5 inst_cell_101_77 (.BL(BL77),.BLN(BLN77),.WL(WL101));
sram_cell_6t_5 inst_cell_101_78 (.BL(BL78),.BLN(BLN78),.WL(WL101));
sram_cell_6t_5 inst_cell_101_79 (.BL(BL79),.BLN(BLN79),.WL(WL101));
sram_cell_6t_5 inst_cell_101_80 (.BL(BL80),.BLN(BLN80),.WL(WL101));
sram_cell_6t_5 inst_cell_101_81 (.BL(BL81),.BLN(BLN81),.WL(WL101));
sram_cell_6t_5 inst_cell_101_82 (.BL(BL82),.BLN(BLN82),.WL(WL101));
sram_cell_6t_5 inst_cell_101_83 (.BL(BL83),.BLN(BLN83),.WL(WL101));
sram_cell_6t_5 inst_cell_101_84 (.BL(BL84),.BLN(BLN84),.WL(WL101));
sram_cell_6t_5 inst_cell_101_85 (.BL(BL85),.BLN(BLN85),.WL(WL101));
sram_cell_6t_5 inst_cell_101_86 (.BL(BL86),.BLN(BLN86),.WL(WL101));
sram_cell_6t_5 inst_cell_101_87 (.BL(BL87),.BLN(BLN87),.WL(WL101));
sram_cell_6t_5 inst_cell_101_88 (.BL(BL88),.BLN(BLN88),.WL(WL101));
sram_cell_6t_5 inst_cell_101_89 (.BL(BL89),.BLN(BLN89),.WL(WL101));
sram_cell_6t_5 inst_cell_101_90 (.BL(BL90),.BLN(BLN90),.WL(WL101));
sram_cell_6t_5 inst_cell_101_91 (.BL(BL91),.BLN(BLN91),.WL(WL101));
sram_cell_6t_5 inst_cell_101_92 (.BL(BL92),.BLN(BLN92),.WL(WL101));
sram_cell_6t_5 inst_cell_101_93 (.BL(BL93),.BLN(BLN93),.WL(WL101));
sram_cell_6t_5 inst_cell_101_94 (.BL(BL94),.BLN(BLN94),.WL(WL101));
sram_cell_6t_5 inst_cell_101_95 (.BL(BL95),.BLN(BLN95),.WL(WL101));
sram_cell_6t_5 inst_cell_101_96 (.BL(BL96),.BLN(BLN96),.WL(WL101));
sram_cell_6t_5 inst_cell_101_97 (.BL(BL97),.BLN(BLN97),.WL(WL101));
sram_cell_6t_5 inst_cell_101_98 (.BL(BL98),.BLN(BLN98),.WL(WL101));
sram_cell_6t_5 inst_cell_101_99 (.BL(BL99),.BLN(BLN99),.WL(WL101));
sram_cell_6t_5 inst_cell_101_100 (.BL(BL100),.BLN(BLN100),.WL(WL101));
sram_cell_6t_5 inst_cell_101_101 (.BL(BL101),.BLN(BLN101),.WL(WL101));
sram_cell_6t_5 inst_cell_101_102 (.BL(BL102),.BLN(BLN102),.WL(WL101));
sram_cell_6t_5 inst_cell_101_103 (.BL(BL103),.BLN(BLN103),.WL(WL101));
sram_cell_6t_5 inst_cell_101_104 (.BL(BL104),.BLN(BLN104),.WL(WL101));
sram_cell_6t_5 inst_cell_101_105 (.BL(BL105),.BLN(BLN105),.WL(WL101));
sram_cell_6t_5 inst_cell_101_106 (.BL(BL106),.BLN(BLN106),.WL(WL101));
sram_cell_6t_5 inst_cell_101_107 (.BL(BL107),.BLN(BLN107),.WL(WL101));
sram_cell_6t_5 inst_cell_101_108 (.BL(BL108),.BLN(BLN108),.WL(WL101));
sram_cell_6t_5 inst_cell_101_109 (.BL(BL109),.BLN(BLN109),.WL(WL101));
sram_cell_6t_5 inst_cell_101_110 (.BL(BL110),.BLN(BLN110),.WL(WL101));
sram_cell_6t_5 inst_cell_101_111 (.BL(BL111),.BLN(BLN111),.WL(WL101));
sram_cell_6t_5 inst_cell_101_112 (.BL(BL112),.BLN(BLN112),.WL(WL101));
sram_cell_6t_5 inst_cell_101_113 (.BL(BL113),.BLN(BLN113),.WL(WL101));
sram_cell_6t_5 inst_cell_101_114 (.BL(BL114),.BLN(BLN114),.WL(WL101));
sram_cell_6t_5 inst_cell_101_115 (.BL(BL115),.BLN(BLN115),.WL(WL101));
sram_cell_6t_5 inst_cell_101_116 (.BL(BL116),.BLN(BLN116),.WL(WL101));
sram_cell_6t_5 inst_cell_101_117 (.BL(BL117),.BLN(BLN117),.WL(WL101));
sram_cell_6t_5 inst_cell_101_118 (.BL(BL118),.BLN(BLN118),.WL(WL101));
sram_cell_6t_5 inst_cell_101_119 (.BL(BL119),.BLN(BLN119),.WL(WL101));
sram_cell_6t_5 inst_cell_101_120 (.BL(BL120),.BLN(BLN120),.WL(WL101));
sram_cell_6t_5 inst_cell_101_121 (.BL(BL121),.BLN(BLN121),.WL(WL101));
sram_cell_6t_5 inst_cell_101_122 (.BL(BL122),.BLN(BLN122),.WL(WL101));
sram_cell_6t_5 inst_cell_101_123 (.BL(BL123),.BLN(BLN123),.WL(WL101));
sram_cell_6t_5 inst_cell_101_124 (.BL(BL124),.BLN(BLN124),.WL(WL101));
sram_cell_6t_5 inst_cell_101_125 (.BL(BL125),.BLN(BLN125),.WL(WL101));
sram_cell_6t_5 inst_cell_101_126 (.BL(BL126),.BLN(BLN126),.WL(WL101));
sram_cell_6t_5 inst_cell_101_127 (.BL(BL127),.BLN(BLN127),.WL(WL101));
sram_cell_6t_5 inst_cell_102_0 (.BL(BL0),.BLN(BLN0),.WL(WL102));
sram_cell_6t_5 inst_cell_102_1 (.BL(BL1),.BLN(BLN1),.WL(WL102));
sram_cell_6t_5 inst_cell_102_2 (.BL(BL2),.BLN(BLN2),.WL(WL102));
sram_cell_6t_5 inst_cell_102_3 (.BL(BL3),.BLN(BLN3),.WL(WL102));
sram_cell_6t_5 inst_cell_102_4 (.BL(BL4),.BLN(BLN4),.WL(WL102));
sram_cell_6t_5 inst_cell_102_5 (.BL(BL5),.BLN(BLN5),.WL(WL102));
sram_cell_6t_5 inst_cell_102_6 (.BL(BL6),.BLN(BLN6),.WL(WL102));
sram_cell_6t_5 inst_cell_102_7 (.BL(BL7),.BLN(BLN7),.WL(WL102));
sram_cell_6t_5 inst_cell_102_8 (.BL(BL8),.BLN(BLN8),.WL(WL102));
sram_cell_6t_5 inst_cell_102_9 (.BL(BL9),.BLN(BLN9),.WL(WL102));
sram_cell_6t_5 inst_cell_102_10 (.BL(BL10),.BLN(BLN10),.WL(WL102));
sram_cell_6t_5 inst_cell_102_11 (.BL(BL11),.BLN(BLN11),.WL(WL102));
sram_cell_6t_5 inst_cell_102_12 (.BL(BL12),.BLN(BLN12),.WL(WL102));
sram_cell_6t_5 inst_cell_102_13 (.BL(BL13),.BLN(BLN13),.WL(WL102));
sram_cell_6t_5 inst_cell_102_14 (.BL(BL14),.BLN(BLN14),.WL(WL102));
sram_cell_6t_5 inst_cell_102_15 (.BL(BL15),.BLN(BLN15),.WL(WL102));
sram_cell_6t_5 inst_cell_102_16 (.BL(BL16),.BLN(BLN16),.WL(WL102));
sram_cell_6t_5 inst_cell_102_17 (.BL(BL17),.BLN(BLN17),.WL(WL102));
sram_cell_6t_5 inst_cell_102_18 (.BL(BL18),.BLN(BLN18),.WL(WL102));
sram_cell_6t_5 inst_cell_102_19 (.BL(BL19),.BLN(BLN19),.WL(WL102));
sram_cell_6t_5 inst_cell_102_20 (.BL(BL20),.BLN(BLN20),.WL(WL102));
sram_cell_6t_5 inst_cell_102_21 (.BL(BL21),.BLN(BLN21),.WL(WL102));
sram_cell_6t_5 inst_cell_102_22 (.BL(BL22),.BLN(BLN22),.WL(WL102));
sram_cell_6t_5 inst_cell_102_23 (.BL(BL23),.BLN(BLN23),.WL(WL102));
sram_cell_6t_5 inst_cell_102_24 (.BL(BL24),.BLN(BLN24),.WL(WL102));
sram_cell_6t_5 inst_cell_102_25 (.BL(BL25),.BLN(BLN25),.WL(WL102));
sram_cell_6t_5 inst_cell_102_26 (.BL(BL26),.BLN(BLN26),.WL(WL102));
sram_cell_6t_5 inst_cell_102_27 (.BL(BL27),.BLN(BLN27),.WL(WL102));
sram_cell_6t_5 inst_cell_102_28 (.BL(BL28),.BLN(BLN28),.WL(WL102));
sram_cell_6t_5 inst_cell_102_29 (.BL(BL29),.BLN(BLN29),.WL(WL102));
sram_cell_6t_5 inst_cell_102_30 (.BL(BL30),.BLN(BLN30),.WL(WL102));
sram_cell_6t_5 inst_cell_102_31 (.BL(BL31),.BLN(BLN31),.WL(WL102));
sram_cell_6t_5 inst_cell_102_32 (.BL(BL32),.BLN(BLN32),.WL(WL102));
sram_cell_6t_5 inst_cell_102_33 (.BL(BL33),.BLN(BLN33),.WL(WL102));
sram_cell_6t_5 inst_cell_102_34 (.BL(BL34),.BLN(BLN34),.WL(WL102));
sram_cell_6t_5 inst_cell_102_35 (.BL(BL35),.BLN(BLN35),.WL(WL102));
sram_cell_6t_5 inst_cell_102_36 (.BL(BL36),.BLN(BLN36),.WL(WL102));
sram_cell_6t_5 inst_cell_102_37 (.BL(BL37),.BLN(BLN37),.WL(WL102));
sram_cell_6t_5 inst_cell_102_38 (.BL(BL38),.BLN(BLN38),.WL(WL102));
sram_cell_6t_5 inst_cell_102_39 (.BL(BL39),.BLN(BLN39),.WL(WL102));
sram_cell_6t_5 inst_cell_102_40 (.BL(BL40),.BLN(BLN40),.WL(WL102));
sram_cell_6t_5 inst_cell_102_41 (.BL(BL41),.BLN(BLN41),.WL(WL102));
sram_cell_6t_5 inst_cell_102_42 (.BL(BL42),.BLN(BLN42),.WL(WL102));
sram_cell_6t_5 inst_cell_102_43 (.BL(BL43),.BLN(BLN43),.WL(WL102));
sram_cell_6t_5 inst_cell_102_44 (.BL(BL44),.BLN(BLN44),.WL(WL102));
sram_cell_6t_5 inst_cell_102_45 (.BL(BL45),.BLN(BLN45),.WL(WL102));
sram_cell_6t_5 inst_cell_102_46 (.BL(BL46),.BLN(BLN46),.WL(WL102));
sram_cell_6t_5 inst_cell_102_47 (.BL(BL47),.BLN(BLN47),.WL(WL102));
sram_cell_6t_5 inst_cell_102_48 (.BL(BL48),.BLN(BLN48),.WL(WL102));
sram_cell_6t_5 inst_cell_102_49 (.BL(BL49),.BLN(BLN49),.WL(WL102));
sram_cell_6t_5 inst_cell_102_50 (.BL(BL50),.BLN(BLN50),.WL(WL102));
sram_cell_6t_5 inst_cell_102_51 (.BL(BL51),.BLN(BLN51),.WL(WL102));
sram_cell_6t_5 inst_cell_102_52 (.BL(BL52),.BLN(BLN52),.WL(WL102));
sram_cell_6t_5 inst_cell_102_53 (.BL(BL53),.BLN(BLN53),.WL(WL102));
sram_cell_6t_5 inst_cell_102_54 (.BL(BL54),.BLN(BLN54),.WL(WL102));
sram_cell_6t_5 inst_cell_102_55 (.BL(BL55),.BLN(BLN55),.WL(WL102));
sram_cell_6t_5 inst_cell_102_56 (.BL(BL56),.BLN(BLN56),.WL(WL102));
sram_cell_6t_5 inst_cell_102_57 (.BL(BL57),.BLN(BLN57),.WL(WL102));
sram_cell_6t_5 inst_cell_102_58 (.BL(BL58),.BLN(BLN58),.WL(WL102));
sram_cell_6t_5 inst_cell_102_59 (.BL(BL59),.BLN(BLN59),.WL(WL102));
sram_cell_6t_5 inst_cell_102_60 (.BL(BL60),.BLN(BLN60),.WL(WL102));
sram_cell_6t_5 inst_cell_102_61 (.BL(BL61),.BLN(BLN61),.WL(WL102));
sram_cell_6t_5 inst_cell_102_62 (.BL(BL62),.BLN(BLN62),.WL(WL102));
sram_cell_6t_5 inst_cell_102_63 (.BL(BL63),.BLN(BLN63),.WL(WL102));
sram_cell_6t_5 inst_cell_102_64 (.BL(BL64),.BLN(BLN64),.WL(WL102));
sram_cell_6t_5 inst_cell_102_65 (.BL(BL65),.BLN(BLN65),.WL(WL102));
sram_cell_6t_5 inst_cell_102_66 (.BL(BL66),.BLN(BLN66),.WL(WL102));
sram_cell_6t_5 inst_cell_102_67 (.BL(BL67),.BLN(BLN67),.WL(WL102));
sram_cell_6t_5 inst_cell_102_68 (.BL(BL68),.BLN(BLN68),.WL(WL102));
sram_cell_6t_5 inst_cell_102_69 (.BL(BL69),.BLN(BLN69),.WL(WL102));
sram_cell_6t_5 inst_cell_102_70 (.BL(BL70),.BLN(BLN70),.WL(WL102));
sram_cell_6t_5 inst_cell_102_71 (.BL(BL71),.BLN(BLN71),.WL(WL102));
sram_cell_6t_5 inst_cell_102_72 (.BL(BL72),.BLN(BLN72),.WL(WL102));
sram_cell_6t_5 inst_cell_102_73 (.BL(BL73),.BLN(BLN73),.WL(WL102));
sram_cell_6t_5 inst_cell_102_74 (.BL(BL74),.BLN(BLN74),.WL(WL102));
sram_cell_6t_5 inst_cell_102_75 (.BL(BL75),.BLN(BLN75),.WL(WL102));
sram_cell_6t_5 inst_cell_102_76 (.BL(BL76),.BLN(BLN76),.WL(WL102));
sram_cell_6t_5 inst_cell_102_77 (.BL(BL77),.BLN(BLN77),.WL(WL102));
sram_cell_6t_5 inst_cell_102_78 (.BL(BL78),.BLN(BLN78),.WL(WL102));
sram_cell_6t_5 inst_cell_102_79 (.BL(BL79),.BLN(BLN79),.WL(WL102));
sram_cell_6t_5 inst_cell_102_80 (.BL(BL80),.BLN(BLN80),.WL(WL102));
sram_cell_6t_5 inst_cell_102_81 (.BL(BL81),.BLN(BLN81),.WL(WL102));
sram_cell_6t_5 inst_cell_102_82 (.BL(BL82),.BLN(BLN82),.WL(WL102));
sram_cell_6t_5 inst_cell_102_83 (.BL(BL83),.BLN(BLN83),.WL(WL102));
sram_cell_6t_5 inst_cell_102_84 (.BL(BL84),.BLN(BLN84),.WL(WL102));
sram_cell_6t_5 inst_cell_102_85 (.BL(BL85),.BLN(BLN85),.WL(WL102));
sram_cell_6t_5 inst_cell_102_86 (.BL(BL86),.BLN(BLN86),.WL(WL102));
sram_cell_6t_5 inst_cell_102_87 (.BL(BL87),.BLN(BLN87),.WL(WL102));
sram_cell_6t_5 inst_cell_102_88 (.BL(BL88),.BLN(BLN88),.WL(WL102));
sram_cell_6t_5 inst_cell_102_89 (.BL(BL89),.BLN(BLN89),.WL(WL102));
sram_cell_6t_5 inst_cell_102_90 (.BL(BL90),.BLN(BLN90),.WL(WL102));
sram_cell_6t_5 inst_cell_102_91 (.BL(BL91),.BLN(BLN91),.WL(WL102));
sram_cell_6t_5 inst_cell_102_92 (.BL(BL92),.BLN(BLN92),.WL(WL102));
sram_cell_6t_5 inst_cell_102_93 (.BL(BL93),.BLN(BLN93),.WL(WL102));
sram_cell_6t_5 inst_cell_102_94 (.BL(BL94),.BLN(BLN94),.WL(WL102));
sram_cell_6t_5 inst_cell_102_95 (.BL(BL95),.BLN(BLN95),.WL(WL102));
sram_cell_6t_5 inst_cell_102_96 (.BL(BL96),.BLN(BLN96),.WL(WL102));
sram_cell_6t_5 inst_cell_102_97 (.BL(BL97),.BLN(BLN97),.WL(WL102));
sram_cell_6t_5 inst_cell_102_98 (.BL(BL98),.BLN(BLN98),.WL(WL102));
sram_cell_6t_5 inst_cell_102_99 (.BL(BL99),.BLN(BLN99),.WL(WL102));
sram_cell_6t_5 inst_cell_102_100 (.BL(BL100),.BLN(BLN100),.WL(WL102));
sram_cell_6t_5 inst_cell_102_101 (.BL(BL101),.BLN(BLN101),.WL(WL102));
sram_cell_6t_5 inst_cell_102_102 (.BL(BL102),.BLN(BLN102),.WL(WL102));
sram_cell_6t_5 inst_cell_102_103 (.BL(BL103),.BLN(BLN103),.WL(WL102));
sram_cell_6t_5 inst_cell_102_104 (.BL(BL104),.BLN(BLN104),.WL(WL102));
sram_cell_6t_5 inst_cell_102_105 (.BL(BL105),.BLN(BLN105),.WL(WL102));
sram_cell_6t_5 inst_cell_102_106 (.BL(BL106),.BLN(BLN106),.WL(WL102));
sram_cell_6t_5 inst_cell_102_107 (.BL(BL107),.BLN(BLN107),.WL(WL102));
sram_cell_6t_5 inst_cell_102_108 (.BL(BL108),.BLN(BLN108),.WL(WL102));
sram_cell_6t_5 inst_cell_102_109 (.BL(BL109),.BLN(BLN109),.WL(WL102));
sram_cell_6t_5 inst_cell_102_110 (.BL(BL110),.BLN(BLN110),.WL(WL102));
sram_cell_6t_5 inst_cell_102_111 (.BL(BL111),.BLN(BLN111),.WL(WL102));
sram_cell_6t_5 inst_cell_102_112 (.BL(BL112),.BLN(BLN112),.WL(WL102));
sram_cell_6t_5 inst_cell_102_113 (.BL(BL113),.BLN(BLN113),.WL(WL102));
sram_cell_6t_5 inst_cell_102_114 (.BL(BL114),.BLN(BLN114),.WL(WL102));
sram_cell_6t_5 inst_cell_102_115 (.BL(BL115),.BLN(BLN115),.WL(WL102));
sram_cell_6t_5 inst_cell_102_116 (.BL(BL116),.BLN(BLN116),.WL(WL102));
sram_cell_6t_5 inst_cell_102_117 (.BL(BL117),.BLN(BLN117),.WL(WL102));
sram_cell_6t_5 inst_cell_102_118 (.BL(BL118),.BLN(BLN118),.WL(WL102));
sram_cell_6t_5 inst_cell_102_119 (.BL(BL119),.BLN(BLN119),.WL(WL102));
sram_cell_6t_5 inst_cell_102_120 (.BL(BL120),.BLN(BLN120),.WL(WL102));
sram_cell_6t_5 inst_cell_102_121 (.BL(BL121),.BLN(BLN121),.WL(WL102));
sram_cell_6t_5 inst_cell_102_122 (.BL(BL122),.BLN(BLN122),.WL(WL102));
sram_cell_6t_5 inst_cell_102_123 (.BL(BL123),.BLN(BLN123),.WL(WL102));
sram_cell_6t_5 inst_cell_102_124 (.BL(BL124),.BLN(BLN124),.WL(WL102));
sram_cell_6t_5 inst_cell_102_125 (.BL(BL125),.BLN(BLN125),.WL(WL102));
sram_cell_6t_5 inst_cell_102_126 (.BL(BL126),.BLN(BLN126),.WL(WL102));
sram_cell_6t_5 inst_cell_102_127 (.BL(BL127),.BLN(BLN127),.WL(WL102));
sram_cell_6t_5 inst_cell_103_0 (.BL(BL0),.BLN(BLN0),.WL(WL103));
sram_cell_6t_5 inst_cell_103_1 (.BL(BL1),.BLN(BLN1),.WL(WL103));
sram_cell_6t_5 inst_cell_103_2 (.BL(BL2),.BLN(BLN2),.WL(WL103));
sram_cell_6t_5 inst_cell_103_3 (.BL(BL3),.BLN(BLN3),.WL(WL103));
sram_cell_6t_5 inst_cell_103_4 (.BL(BL4),.BLN(BLN4),.WL(WL103));
sram_cell_6t_5 inst_cell_103_5 (.BL(BL5),.BLN(BLN5),.WL(WL103));
sram_cell_6t_5 inst_cell_103_6 (.BL(BL6),.BLN(BLN6),.WL(WL103));
sram_cell_6t_5 inst_cell_103_7 (.BL(BL7),.BLN(BLN7),.WL(WL103));
sram_cell_6t_5 inst_cell_103_8 (.BL(BL8),.BLN(BLN8),.WL(WL103));
sram_cell_6t_5 inst_cell_103_9 (.BL(BL9),.BLN(BLN9),.WL(WL103));
sram_cell_6t_5 inst_cell_103_10 (.BL(BL10),.BLN(BLN10),.WL(WL103));
sram_cell_6t_5 inst_cell_103_11 (.BL(BL11),.BLN(BLN11),.WL(WL103));
sram_cell_6t_5 inst_cell_103_12 (.BL(BL12),.BLN(BLN12),.WL(WL103));
sram_cell_6t_5 inst_cell_103_13 (.BL(BL13),.BLN(BLN13),.WL(WL103));
sram_cell_6t_5 inst_cell_103_14 (.BL(BL14),.BLN(BLN14),.WL(WL103));
sram_cell_6t_5 inst_cell_103_15 (.BL(BL15),.BLN(BLN15),.WL(WL103));
sram_cell_6t_5 inst_cell_103_16 (.BL(BL16),.BLN(BLN16),.WL(WL103));
sram_cell_6t_5 inst_cell_103_17 (.BL(BL17),.BLN(BLN17),.WL(WL103));
sram_cell_6t_5 inst_cell_103_18 (.BL(BL18),.BLN(BLN18),.WL(WL103));
sram_cell_6t_5 inst_cell_103_19 (.BL(BL19),.BLN(BLN19),.WL(WL103));
sram_cell_6t_5 inst_cell_103_20 (.BL(BL20),.BLN(BLN20),.WL(WL103));
sram_cell_6t_5 inst_cell_103_21 (.BL(BL21),.BLN(BLN21),.WL(WL103));
sram_cell_6t_5 inst_cell_103_22 (.BL(BL22),.BLN(BLN22),.WL(WL103));
sram_cell_6t_5 inst_cell_103_23 (.BL(BL23),.BLN(BLN23),.WL(WL103));
sram_cell_6t_5 inst_cell_103_24 (.BL(BL24),.BLN(BLN24),.WL(WL103));
sram_cell_6t_5 inst_cell_103_25 (.BL(BL25),.BLN(BLN25),.WL(WL103));
sram_cell_6t_5 inst_cell_103_26 (.BL(BL26),.BLN(BLN26),.WL(WL103));
sram_cell_6t_5 inst_cell_103_27 (.BL(BL27),.BLN(BLN27),.WL(WL103));
sram_cell_6t_5 inst_cell_103_28 (.BL(BL28),.BLN(BLN28),.WL(WL103));
sram_cell_6t_5 inst_cell_103_29 (.BL(BL29),.BLN(BLN29),.WL(WL103));
sram_cell_6t_5 inst_cell_103_30 (.BL(BL30),.BLN(BLN30),.WL(WL103));
sram_cell_6t_5 inst_cell_103_31 (.BL(BL31),.BLN(BLN31),.WL(WL103));
sram_cell_6t_5 inst_cell_103_32 (.BL(BL32),.BLN(BLN32),.WL(WL103));
sram_cell_6t_5 inst_cell_103_33 (.BL(BL33),.BLN(BLN33),.WL(WL103));
sram_cell_6t_5 inst_cell_103_34 (.BL(BL34),.BLN(BLN34),.WL(WL103));
sram_cell_6t_5 inst_cell_103_35 (.BL(BL35),.BLN(BLN35),.WL(WL103));
sram_cell_6t_5 inst_cell_103_36 (.BL(BL36),.BLN(BLN36),.WL(WL103));
sram_cell_6t_5 inst_cell_103_37 (.BL(BL37),.BLN(BLN37),.WL(WL103));
sram_cell_6t_5 inst_cell_103_38 (.BL(BL38),.BLN(BLN38),.WL(WL103));
sram_cell_6t_5 inst_cell_103_39 (.BL(BL39),.BLN(BLN39),.WL(WL103));
sram_cell_6t_5 inst_cell_103_40 (.BL(BL40),.BLN(BLN40),.WL(WL103));
sram_cell_6t_5 inst_cell_103_41 (.BL(BL41),.BLN(BLN41),.WL(WL103));
sram_cell_6t_5 inst_cell_103_42 (.BL(BL42),.BLN(BLN42),.WL(WL103));
sram_cell_6t_5 inst_cell_103_43 (.BL(BL43),.BLN(BLN43),.WL(WL103));
sram_cell_6t_5 inst_cell_103_44 (.BL(BL44),.BLN(BLN44),.WL(WL103));
sram_cell_6t_5 inst_cell_103_45 (.BL(BL45),.BLN(BLN45),.WL(WL103));
sram_cell_6t_5 inst_cell_103_46 (.BL(BL46),.BLN(BLN46),.WL(WL103));
sram_cell_6t_5 inst_cell_103_47 (.BL(BL47),.BLN(BLN47),.WL(WL103));
sram_cell_6t_5 inst_cell_103_48 (.BL(BL48),.BLN(BLN48),.WL(WL103));
sram_cell_6t_5 inst_cell_103_49 (.BL(BL49),.BLN(BLN49),.WL(WL103));
sram_cell_6t_5 inst_cell_103_50 (.BL(BL50),.BLN(BLN50),.WL(WL103));
sram_cell_6t_5 inst_cell_103_51 (.BL(BL51),.BLN(BLN51),.WL(WL103));
sram_cell_6t_5 inst_cell_103_52 (.BL(BL52),.BLN(BLN52),.WL(WL103));
sram_cell_6t_5 inst_cell_103_53 (.BL(BL53),.BLN(BLN53),.WL(WL103));
sram_cell_6t_5 inst_cell_103_54 (.BL(BL54),.BLN(BLN54),.WL(WL103));
sram_cell_6t_5 inst_cell_103_55 (.BL(BL55),.BLN(BLN55),.WL(WL103));
sram_cell_6t_5 inst_cell_103_56 (.BL(BL56),.BLN(BLN56),.WL(WL103));
sram_cell_6t_5 inst_cell_103_57 (.BL(BL57),.BLN(BLN57),.WL(WL103));
sram_cell_6t_5 inst_cell_103_58 (.BL(BL58),.BLN(BLN58),.WL(WL103));
sram_cell_6t_5 inst_cell_103_59 (.BL(BL59),.BLN(BLN59),.WL(WL103));
sram_cell_6t_5 inst_cell_103_60 (.BL(BL60),.BLN(BLN60),.WL(WL103));
sram_cell_6t_5 inst_cell_103_61 (.BL(BL61),.BLN(BLN61),.WL(WL103));
sram_cell_6t_5 inst_cell_103_62 (.BL(BL62),.BLN(BLN62),.WL(WL103));
sram_cell_6t_5 inst_cell_103_63 (.BL(BL63),.BLN(BLN63),.WL(WL103));
sram_cell_6t_5 inst_cell_103_64 (.BL(BL64),.BLN(BLN64),.WL(WL103));
sram_cell_6t_5 inst_cell_103_65 (.BL(BL65),.BLN(BLN65),.WL(WL103));
sram_cell_6t_5 inst_cell_103_66 (.BL(BL66),.BLN(BLN66),.WL(WL103));
sram_cell_6t_5 inst_cell_103_67 (.BL(BL67),.BLN(BLN67),.WL(WL103));
sram_cell_6t_5 inst_cell_103_68 (.BL(BL68),.BLN(BLN68),.WL(WL103));
sram_cell_6t_5 inst_cell_103_69 (.BL(BL69),.BLN(BLN69),.WL(WL103));
sram_cell_6t_5 inst_cell_103_70 (.BL(BL70),.BLN(BLN70),.WL(WL103));
sram_cell_6t_5 inst_cell_103_71 (.BL(BL71),.BLN(BLN71),.WL(WL103));
sram_cell_6t_5 inst_cell_103_72 (.BL(BL72),.BLN(BLN72),.WL(WL103));
sram_cell_6t_5 inst_cell_103_73 (.BL(BL73),.BLN(BLN73),.WL(WL103));
sram_cell_6t_5 inst_cell_103_74 (.BL(BL74),.BLN(BLN74),.WL(WL103));
sram_cell_6t_5 inst_cell_103_75 (.BL(BL75),.BLN(BLN75),.WL(WL103));
sram_cell_6t_5 inst_cell_103_76 (.BL(BL76),.BLN(BLN76),.WL(WL103));
sram_cell_6t_5 inst_cell_103_77 (.BL(BL77),.BLN(BLN77),.WL(WL103));
sram_cell_6t_5 inst_cell_103_78 (.BL(BL78),.BLN(BLN78),.WL(WL103));
sram_cell_6t_5 inst_cell_103_79 (.BL(BL79),.BLN(BLN79),.WL(WL103));
sram_cell_6t_5 inst_cell_103_80 (.BL(BL80),.BLN(BLN80),.WL(WL103));
sram_cell_6t_5 inst_cell_103_81 (.BL(BL81),.BLN(BLN81),.WL(WL103));
sram_cell_6t_5 inst_cell_103_82 (.BL(BL82),.BLN(BLN82),.WL(WL103));
sram_cell_6t_5 inst_cell_103_83 (.BL(BL83),.BLN(BLN83),.WL(WL103));
sram_cell_6t_5 inst_cell_103_84 (.BL(BL84),.BLN(BLN84),.WL(WL103));
sram_cell_6t_5 inst_cell_103_85 (.BL(BL85),.BLN(BLN85),.WL(WL103));
sram_cell_6t_5 inst_cell_103_86 (.BL(BL86),.BLN(BLN86),.WL(WL103));
sram_cell_6t_5 inst_cell_103_87 (.BL(BL87),.BLN(BLN87),.WL(WL103));
sram_cell_6t_5 inst_cell_103_88 (.BL(BL88),.BLN(BLN88),.WL(WL103));
sram_cell_6t_5 inst_cell_103_89 (.BL(BL89),.BLN(BLN89),.WL(WL103));
sram_cell_6t_5 inst_cell_103_90 (.BL(BL90),.BLN(BLN90),.WL(WL103));
sram_cell_6t_5 inst_cell_103_91 (.BL(BL91),.BLN(BLN91),.WL(WL103));
sram_cell_6t_5 inst_cell_103_92 (.BL(BL92),.BLN(BLN92),.WL(WL103));
sram_cell_6t_5 inst_cell_103_93 (.BL(BL93),.BLN(BLN93),.WL(WL103));
sram_cell_6t_5 inst_cell_103_94 (.BL(BL94),.BLN(BLN94),.WL(WL103));
sram_cell_6t_5 inst_cell_103_95 (.BL(BL95),.BLN(BLN95),.WL(WL103));
sram_cell_6t_5 inst_cell_103_96 (.BL(BL96),.BLN(BLN96),.WL(WL103));
sram_cell_6t_5 inst_cell_103_97 (.BL(BL97),.BLN(BLN97),.WL(WL103));
sram_cell_6t_5 inst_cell_103_98 (.BL(BL98),.BLN(BLN98),.WL(WL103));
sram_cell_6t_5 inst_cell_103_99 (.BL(BL99),.BLN(BLN99),.WL(WL103));
sram_cell_6t_5 inst_cell_103_100 (.BL(BL100),.BLN(BLN100),.WL(WL103));
sram_cell_6t_5 inst_cell_103_101 (.BL(BL101),.BLN(BLN101),.WL(WL103));
sram_cell_6t_5 inst_cell_103_102 (.BL(BL102),.BLN(BLN102),.WL(WL103));
sram_cell_6t_5 inst_cell_103_103 (.BL(BL103),.BLN(BLN103),.WL(WL103));
sram_cell_6t_5 inst_cell_103_104 (.BL(BL104),.BLN(BLN104),.WL(WL103));
sram_cell_6t_5 inst_cell_103_105 (.BL(BL105),.BLN(BLN105),.WL(WL103));
sram_cell_6t_5 inst_cell_103_106 (.BL(BL106),.BLN(BLN106),.WL(WL103));
sram_cell_6t_5 inst_cell_103_107 (.BL(BL107),.BLN(BLN107),.WL(WL103));
sram_cell_6t_5 inst_cell_103_108 (.BL(BL108),.BLN(BLN108),.WL(WL103));
sram_cell_6t_5 inst_cell_103_109 (.BL(BL109),.BLN(BLN109),.WL(WL103));
sram_cell_6t_5 inst_cell_103_110 (.BL(BL110),.BLN(BLN110),.WL(WL103));
sram_cell_6t_5 inst_cell_103_111 (.BL(BL111),.BLN(BLN111),.WL(WL103));
sram_cell_6t_5 inst_cell_103_112 (.BL(BL112),.BLN(BLN112),.WL(WL103));
sram_cell_6t_5 inst_cell_103_113 (.BL(BL113),.BLN(BLN113),.WL(WL103));
sram_cell_6t_5 inst_cell_103_114 (.BL(BL114),.BLN(BLN114),.WL(WL103));
sram_cell_6t_5 inst_cell_103_115 (.BL(BL115),.BLN(BLN115),.WL(WL103));
sram_cell_6t_5 inst_cell_103_116 (.BL(BL116),.BLN(BLN116),.WL(WL103));
sram_cell_6t_5 inst_cell_103_117 (.BL(BL117),.BLN(BLN117),.WL(WL103));
sram_cell_6t_5 inst_cell_103_118 (.BL(BL118),.BLN(BLN118),.WL(WL103));
sram_cell_6t_5 inst_cell_103_119 (.BL(BL119),.BLN(BLN119),.WL(WL103));
sram_cell_6t_5 inst_cell_103_120 (.BL(BL120),.BLN(BLN120),.WL(WL103));
sram_cell_6t_5 inst_cell_103_121 (.BL(BL121),.BLN(BLN121),.WL(WL103));
sram_cell_6t_5 inst_cell_103_122 (.BL(BL122),.BLN(BLN122),.WL(WL103));
sram_cell_6t_5 inst_cell_103_123 (.BL(BL123),.BLN(BLN123),.WL(WL103));
sram_cell_6t_5 inst_cell_103_124 (.BL(BL124),.BLN(BLN124),.WL(WL103));
sram_cell_6t_5 inst_cell_103_125 (.BL(BL125),.BLN(BLN125),.WL(WL103));
sram_cell_6t_5 inst_cell_103_126 (.BL(BL126),.BLN(BLN126),.WL(WL103));
sram_cell_6t_5 inst_cell_103_127 (.BL(BL127),.BLN(BLN127),.WL(WL103));
sram_cell_6t_5 inst_cell_104_0 (.BL(BL0),.BLN(BLN0),.WL(WL104));
sram_cell_6t_5 inst_cell_104_1 (.BL(BL1),.BLN(BLN1),.WL(WL104));
sram_cell_6t_5 inst_cell_104_2 (.BL(BL2),.BLN(BLN2),.WL(WL104));
sram_cell_6t_5 inst_cell_104_3 (.BL(BL3),.BLN(BLN3),.WL(WL104));
sram_cell_6t_5 inst_cell_104_4 (.BL(BL4),.BLN(BLN4),.WL(WL104));
sram_cell_6t_5 inst_cell_104_5 (.BL(BL5),.BLN(BLN5),.WL(WL104));
sram_cell_6t_5 inst_cell_104_6 (.BL(BL6),.BLN(BLN6),.WL(WL104));
sram_cell_6t_5 inst_cell_104_7 (.BL(BL7),.BLN(BLN7),.WL(WL104));
sram_cell_6t_5 inst_cell_104_8 (.BL(BL8),.BLN(BLN8),.WL(WL104));
sram_cell_6t_5 inst_cell_104_9 (.BL(BL9),.BLN(BLN9),.WL(WL104));
sram_cell_6t_5 inst_cell_104_10 (.BL(BL10),.BLN(BLN10),.WL(WL104));
sram_cell_6t_5 inst_cell_104_11 (.BL(BL11),.BLN(BLN11),.WL(WL104));
sram_cell_6t_5 inst_cell_104_12 (.BL(BL12),.BLN(BLN12),.WL(WL104));
sram_cell_6t_5 inst_cell_104_13 (.BL(BL13),.BLN(BLN13),.WL(WL104));
sram_cell_6t_5 inst_cell_104_14 (.BL(BL14),.BLN(BLN14),.WL(WL104));
sram_cell_6t_5 inst_cell_104_15 (.BL(BL15),.BLN(BLN15),.WL(WL104));
sram_cell_6t_5 inst_cell_104_16 (.BL(BL16),.BLN(BLN16),.WL(WL104));
sram_cell_6t_5 inst_cell_104_17 (.BL(BL17),.BLN(BLN17),.WL(WL104));
sram_cell_6t_5 inst_cell_104_18 (.BL(BL18),.BLN(BLN18),.WL(WL104));
sram_cell_6t_5 inst_cell_104_19 (.BL(BL19),.BLN(BLN19),.WL(WL104));
sram_cell_6t_5 inst_cell_104_20 (.BL(BL20),.BLN(BLN20),.WL(WL104));
sram_cell_6t_5 inst_cell_104_21 (.BL(BL21),.BLN(BLN21),.WL(WL104));
sram_cell_6t_5 inst_cell_104_22 (.BL(BL22),.BLN(BLN22),.WL(WL104));
sram_cell_6t_5 inst_cell_104_23 (.BL(BL23),.BLN(BLN23),.WL(WL104));
sram_cell_6t_5 inst_cell_104_24 (.BL(BL24),.BLN(BLN24),.WL(WL104));
sram_cell_6t_5 inst_cell_104_25 (.BL(BL25),.BLN(BLN25),.WL(WL104));
sram_cell_6t_5 inst_cell_104_26 (.BL(BL26),.BLN(BLN26),.WL(WL104));
sram_cell_6t_5 inst_cell_104_27 (.BL(BL27),.BLN(BLN27),.WL(WL104));
sram_cell_6t_5 inst_cell_104_28 (.BL(BL28),.BLN(BLN28),.WL(WL104));
sram_cell_6t_5 inst_cell_104_29 (.BL(BL29),.BLN(BLN29),.WL(WL104));
sram_cell_6t_5 inst_cell_104_30 (.BL(BL30),.BLN(BLN30),.WL(WL104));
sram_cell_6t_5 inst_cell_104_31 (.BL(BL31),.BLN(BLN31),.WL(WL104));
sram_cell_6t_5 inst_cell_104_32 (.BL(BL32),.BLN(BLN32),.WL(WL104));
sram_cell_6t_5 inst_cell_104_33 (.BL(BL33),.BLN(BLN33),.WL(WL104));
sram_cell_6t_5 inst_cell_104_34 (.BL(BL34),.BLN(BLN34),.WL(WL104));
sram_cell_6t_5 inst_cell_104_35 (.BL(BL35),.BLN(BLN35),.WL(WL104));
sram_cell_6t_5 inst_cell_104_36 (.BL(BL36),.BLN(BLN36),.WL(WL104));
sram_cell_6t_5 inst_cell_104_37 (.BL(BL37),.BLN(BLN37),.WL(WL104));
sram_cell_6t_5 inst_cell_104_38 (.BL(BL38),.BLN(BLN38),.WL(WL104));
sram_cell_6t_5 inst_cell_104_39 (.BL(BL39),.BLN(BLN39),.WL(WL104));
sram_cell_6t_5 inst_cell_104_40 (.BL(BL40),.BLN(BLN40),.WL(WL104));
sram_cell_6t_5 inst_cell_104_41 (.BL(BL41),.BLN(BLN41),.WL(WL104));
sram_cell_6t_5 inst_cell_104_42 (.BL(BL42),.BLN(BLN42),.WL(WL104));
sram_cell_6t_5 inst_cell_104_43 (.BL(BL43),.BLN(BLN43),.WL(WL104));
sram_cell_6t_5 inst_cell_104_44 (.BL(BL44),.BLN(BLN44),.WL(WL104));
sram_cell_6t_5 inst_cell_104_45 (.BL(BL45),.BLN(BLN45),.WL(WL104));
sram_cell_6t_5 inst_cell_104_46 (.BL(BL46),.BLN(BLN46),.WL(WL104));
sram_cell_6t_5 inst_cell_104_47 (.BL(BL47),.BLN(BLN47),.WL(WL104));
sram_cell_6t_5 inst_cell_104_48 (.BL(BL48),.BLN(BLN48),.WL(WL104));
sram_cell_6t_5 inst_cell_104_49 (.BL(BL49),.BLN(BLN49),.WL(WL104));
sram_cell_6t_5 inst_cell_104_50 (.BL(BL50),.BLN(BLN50),.WL(WL104));
sram_cell_6t_5 inst_cell_104_51 (.BL(BL51),.BLN(BLN51),.WL(WL104));
sram_cell_6t_5 inst_cell_104_52 (.BL(BL52),.BLN(BLN52),.WL(WL104));
sram_cell_6t_5 inst_cell_104_53 (.BL(BL53),.BLN(BLN53),.WL(WL104));
sram_cell_6t_5 inst_cell_104_54 (.BL(BL54),.BLN(BLN54),.WL(WL104));
sram_cell_6t_5 inst_cell_104_55 (.BL(BL55),.BLN(BLN55),.WL(WL104));
sram_cell_6t_5 inst_cell_104_56 (.BL(BL56),.BLN(BLN56),.WL(WL104));
sram_cell_6t_5 inst_cell_104_57 (.BL(BL57),.BLN(BLN57),.WL(WL104));
sram_cell_6t_5 inst_cell_104_58 (.BL(BL58),.BLN(BLN58),.WL(WL104));
sram_cell_6t_5 inst_cell_104_59 (.BL(BL59),.BLN(BLN59),.WL(WL104));
sram_cell_6t_5 inst_cell_104_60 (.BL(BL60),.BLN(BLN60),.WL(WL104));
sram_cell_6t_5 inst_cell_104_61 (.BL(BL61),.BLN(BLN61),.WL(WL104));
sram_cell_6t_5 inst_cell_104_62 (.BL(BL62),.BLN(BLN62),.WL(WL104));
sram_cell_6t_5 inst_cell_104_63 (.BL(BL63),.BLN(BLN63),.WL(WL104));
sram_cell_6t_5 inst_cell_104_64 (.BL(BL64),.BLN(BLN64),.WL(WL104));
sram_cell_6t_5 inst_cell_104_65 (.BL(BL65),.BLN(BLN65),.WL(WL104));
sram_cell_6t_5 inst_cell_104_66 (.BL(BL66),.BLN(BLN66),.WL(WL104));
sram_cell_6t_5 inst_cell_104_67 (.BL(BL67),.BLN(BLN67),.WL(WL104));
sram_cell_6t_5 inst_cell_104_68 (.BL(BL68),.BLN(BLN68),.WL(WL104));
sram_cell_6t_5 inst_cell_104_69 (.BL(BL69),.BLN(BLN69),.WL(WL104));
sram_cell_6t_5 inst_cell_104_70 (.BL(BL70),.BLN(BLN70),.WL(WL104));
sram_cell_6t_5 inst_cell_104_71 (.BL(BL71),.BLN(BLN71),.WL(WL104));
sram_cell_6t_5 inst_cell_104_72 (.BL(BL72),.BLN(BLN72),.WL(WL104));
sram_cell_6t_5 inst_cell_104_73 (.BL(BL73),.BLN(BLN73),.WL(WL104));
sram_cell_6t_5 inst_cell_104_74 (.BL(BL74),.BLN(BLN74),.WL(WL104));
sram_cell_6t_5 inst_cell_104_75 (.BL(BL75),.BLN(BLN75),.WL(WL104));
sram_cell_6t_5 inst_cell_104_76 (.BL(BL76),.BLN(BLN76),.WL(WL104));
sram_cell_6t_5 inst_cell_104_77 (.BL(BL77),.BLN(BLN77),.WL(WL104));
sram_cell_6t_5 inst_cell_104_78 (.BL(BL78),.BLN(BLN78),.WL(WL104));
sram_cell_6t_5 inst_cell_104_79 (.BL(BL79),.BLN(BLN79),.WL(WL104));
sram_cell_6t_5 inst_cell_104_80 (.BL(BL80),.BLN(BLN80),.WL(WL104));
sram_cell_6t_5 inst_cell_104_81 (.BL(BL81),.BLN(BLN81),.WL(WL104));
sram_cell_6t_5 inst_cell_104_82 (.BL(BL82),.BLN(BLN82),.WL(WL104));
sram_cell_6t_5 inst_cell_104_83 (.BL(BL83),.BLN(BLN83),.WL(WL104));
sram_cell_6t_5 inst_cell_104_84 (.BL(BL84),.BLN(BLN84),.WL(WL104));
sram_cell_6t_5 inst_cell_104_85 (.BL(BL85),.BLN(BLN85),.WL(WL104));
sram_cell_6t_5 inst_cell_104_86 (.BL(BL86),.BLN(BLN86),.WL(WL104));
sram_cell_6t_5 inst_cell_104_87 (.BL(BL87),.BLN(BLN87),.WL(WL104));
sram_cell_6t_5 inst_cell_104_88 (.BL(BL88),.BLN(BLN88),.WL(WL104));
sram_cell_6t_5 inst_cell_104_89 (.BL(BL89),.BLN(BLN89),.WL(WL104));
sram_cell_6t_5 inst_cell_104_90 (.BL(BL90),.BLN(BLN90),.WL(WL104));
sram_cell_6t_5 inst_cell_104_91 (.BL(BL91),.BLN(BLN91),.WL(WL104));
sram_cell_6t_5 inst_cell_104_92 (.BL(BL92),.BLN(BLN92),.WL(WL104));
sram_cell_6t_5 inst_cell_104_93 (.BL(BL93),.BLN(BLN93),.WL(WL104));
sram_cell_6t_5 inst_cell_104_94 (.BL(BL94),.BLN(BLN94),.WL(WL104));
sram_cell_6t_5 inst_cell_104_95 (.BL(BL95),.BLN(BLN95),.WL(WL104));
sram_cell_6t_5 inst_cell_104_96 (.BL(BL96),.BLN(BLN96),.WL(WL104));
sram_cell_6t_5 inst_cell_104_97 (.BL(BL97),.BLN(BLN97),.WL(WL104));
sram_cell_6t_5 inst_cell_104_98 (.BL(BL98),.BLN(BLN98),.WL(WL104));
sram_cell_6t_5 inst_cell_104_99 (.BL(BL99),.BLN(BLN99),.WL(WL104));
sram_cell_6t_5 inst_cell_104_100 (.BL(BL100),.BLN(BLN100),.WL(WL104));
sram_cell_6t_5 inst_cell_104_101 (.BL(BL101),.BLN(BLN101),.WL(WL104));
sram_cell_6t_5 inst_cell_104_102 (.BL(BL102),.BLN(BLN102),.WL(WL104));
sram_cell_6t_5 inst_cell_104_103 (.BL(BL103),.BLN(BLN103),.WL(WL104));
sram_cell_6t_5 inst_cell_104_104 (.BL(BL104),.BLN(BLN104),.WL(WL104));
sram_cell_6t_5 inst_cell_104_105 (.BL(BL105),.BLN(BLN105),.WL(WL104));
sram_cell_6t_5 inst_cell_104_106 (.BL(BL106),.BLN(BLN106),.WL(WL104));
sram_cell_6t_5 inst_cell_104_107 (.BL(BL107),.BLN(BLN107),.WL(WL104));
sram_cell_6t_5 inst_cell_104_108 (.BL(BL108),.BLN(BLN108),.WL(WL104));
sram_cell_6t_5 inst_cell_104_109 (.BL(BL109),.BLN(BLN109),.WL(WL104));
sram_cell_6t_5 inst_cell_104_110 (.BL(BL110),.BLN(BLN110),.WL(WL104));
sram_cell_6t_5 inst_cell_104_111 (.BL(BL111),.BLN(BLN111),.WL(WL104));
sram_cell_6t_5 inst_cell_104_112 (.BL(BL112),.BLN(BLN112),.WL(WL104));
sram_cell_6t_5 inst_cell_104_113 (.BL(BL113),.BLN(BLN113),.WL(WL104));
sram_cell_6t_5 inst_cell_104_114 (.BL(BL114),.BLN(BLN114),.WL(WL104));
sram_cell_6t_5 inst_cell_104_115 (.BL(BL115),.BLN(BLN115),.WL(WL104));
sram_cell_6t_5 inst_cell_104_116 (.BL(BL116),.BLN(BLN116),.WL(WL104));
sram_cell_6t_5 inst_cell_104_117 (.BL(BL117),.BLN(BLN117),.WL(WL104));
sram_cell_6t_5 inst_cell_104_118 (.BL(BL118),.BLN(BLN118),.WL(WL104));
sram_cell_6t_5 inst_cell_104_119 (.BL(BL119),.BLN(BLN119),.WL(WL104));
sram_cell_6t_5 inst_cell_104_120 (.BL(BL120),.BLN(BLN120),.WL(WL104));
sram_cell_6t_5 inst_cell_104_121 (.BL(BL121),.BLN(BLN121),.WL(WL104));
sram_cell_6t_5 inst_cell_104_122 (.BL(BL122),.BLN(BLN122),.WL(WL104));
sram_cell_6t_5 inst_cell_104_123 (.BL(BL123),.BLN(BLN123),.WL(WL104));
sram_cell_6t_5 inst_cell_104_124 (.BL(BL124),.BLN(BLN124),.WL(WL104));
sram_cell_6t_5 inst_cell_104_125 (.BL(BL125),.BLN(BLN125),.WL(WL104));
sram_cell_6t_5 inst_cell_104_126 (.BL(BL126),.BLN(BLN126),.WL(WL104));
sram_cell_6t_5 inst_cell_104_127 (.BL(BL127),.BLN(BLN127),.WL(WL104));
sram_cell_6t_5 inst_cell_105_0 (.BL(BL0),.BLN(BLN0),.WL(WL105));
sram_cell_6t_5 inst_cell_105_1 (.BL(BL1),.BLN(BLN1),.WL(WL105));
sram_cell_6t_5 inst_cell_105_2 (.BL(BL2),.BLN(BLN2),.WL(WL105));
sram_cell_6t_5 inst_cell_105_3 (.BL(BL3),.BLN(BLN3),.WL(WL105));
sram_cell_6t_5 inst_cell_105_4 (.BL(BL4),.BLN(BLN4),.WL(WL105));
sram_cell_6t_5 inst_cell_105_5 (.BL(BL5),.BLN(BLN5),.WL(WL105));
sram_cell_6t_5 inst_cell_105_6 (.BL(BL6),.BLN(BLN6),.WL(WL105));
sram_cell_6t_5 inst_cell_105_7 (.BL(BL7),.BLN(BLN7),.WL(WL105));
sram_cell_6t_5 inst_cell_105_8 (.BL(BL8),.BLN(BLN8),.WL(WL105));
sram_cell_6t_5 inst_cell_105_9 (.BL(BL9),.BLN(BLN9),.WL(WL105));
sram_cell_6t_5 inst_cell_105_10 (.BL(BL10),.BLN(BLN10),.WL(WL105));
sram_cell_6t_5 inst_cell_105_11 (.BL(BL11),.BLN(BLN11),.WL(WL105));
sram_cell_6t_5 inst_cell_105_12 (.BL(BL12),.BLN(BLN12),.WL(WL105));
sram_cell_6t_5 inst_cell_105_13 (.BL(BL13),.BLN(BLN13),.WL(WL105));
sram_cell_6t_5 inst_cell_105_14 (.BL(BL14),.BLN(BLN14),.WL(WL105));
sram_cell_6t_5 inst_cell_105_15 (.BL(BL15),.BLN(BLN15),.WL(WL105));
sram_cell_6t_5 inst_cell_105_16 (.BL(BL16),.BLN(BLN16),.WL(WL105));
sram_cell_6t_5 inst_cell_105_17 (.BL(BL17),.BLN(BLN17),.WL(WL105));
sram_cell_6t_5 inst_cell_105_18 (.BL(BL18),.BLN(BLN18),.WL(WL105));
sram_cell_6t_5 inst_cell_105_19 (.BL(BL19),.BLN(BLN19),.WL(WL105));
sram_cell_6t_5 inst_cell_105_20 (.BL(BL20),.BLN(BLN20),.WL(WL105));
sram_cell_6t_5 inst_cell_105_21 (.BL(BL21),.BLN(BLN21),.WL(WL105));
sram_cell_6t_5 inst_cell_105_22 (.BL(BL22),.BLN(BLN22),.WL(WL105));
sram_cell_6t_5 inst_cell_105_23 (.BL(BL23),.BLN(BLN23),.WL(WL105));
sram_cell_6t_5 inst_cell_105_24 (.BL(BL24),.BLN(BLN24),.WL(WL105));
sram_cell_6t_5 inst_cell_105_25 (.BL(BL25),.BLN(BLN25),.WL(WL105));
sram_cell_6t_5 inst_cell_105_26 (.BL(BL26),.BLN(BLN26),.WL(WL105));
sram_cell_6t_5 inst_cell_105_27 (.BL(BL27),.BLN(BLN27),.WL(WL105));
sram_cell_6t_5 inst_cell_105_28 (.BL(BL28),.BLN(BLN28),.WL(WL105));
sram_cell_6t_5 inst_cell_105_29 (.BL(BL29),.BLN(BLN29),.WL(WL105));
sram_cell_6t_5 inst_cell_105_30 (.BL(BL30),.BLN(BLN30),.WL(WL105));
sram_cell_6t_5 inst_cell_105_31 (.BL(BL31),.BLN(BLN31),.WL(WL105));
sram_cell_6t_5 inst_cell_105_32 (.BL(BL32),.BLN(BLN32),.WL(WL105));
sram_cell_6t_5 inst_cell_105_33 (.BL(BL33),.BLN(BLN33),.WL(WL105));
sram_cell_6t_5 inst_cell_105_34 (.BL(BL34),.BLN(BLN34),.WL(WL105));
sram_cell_6t_5 inst_cell_105_35 (.BL(BL35),.BLN(BLN35),.WL(WL105));
sram_cell_6t_5 inst_cell_105_36 (.BL(BL36),.BLN(BLN36),.WL(WL105));
sram_cell_6t_5 inst_cell_105_37 (.BL(BL37),.BLN(BLN37),.WL(WL105));
sram_cell_6t_5 inst_cell_105_38 (.BL(BL38),.BLN(BLN38),.WL(WL105));
sram_cell_6t_5 inst_cell_105_39 (.BL(BL39),.BLN(BLN39),.WL(WL105));
sram_cell_6t_5 inst_cell_105_40 (.BL(BL40),.BLN(BLN40),.WL(WL105));
sram_cell_6t_5 inst_cell_105_41 (.BL(BL41),.BLN(BLN41),.WL(WL105));
sram_cell_6t_5 inst_cell_105_42 (.BL(BL42),.BLN(BLN42),.WL(WL105));
sram_cell_6t_5 inst_cell_105_43 (.BL(BL43),.BLN(BLN43),.WL(WL105));
sram_cell_6t_5 inst_cell_105_44 (.BL(BL44),.BLN(BLN44),.WL(WL105));
sram_cell_6t_5 inst_cell_105_45 (.BL(BL45),.BLN(BLN45),.WL(WL105));
sram_cell_6t_5 inst_cell_105_46 (.BL(BL46),.BLN(BLN46),.WL(WL105));
sram_cell_6t_5 inst_cell_105_47 (.BL(BL47),.BLN(BLN47),.WL(WL105));
sram_cell_6t_5 inst_cell_105_48 (.BL(BL48),.BLN(BLN48),.WL(WL105));
sram_cell_6t_5 inst_cell_105_49 (.BL(BL49),.BLN(BLN49),.WL(WL105));
sram_cell_6t_5 inst_cell_105_50 (.BL(BL50),.BLN(BLN50),.WL(WL105));
sram_cell_6t_5 inst_cell_105_51 (.BL(BL51),.BLN(BLN51),.WL(WL105));
sram_cell_6t_5 inst_cell_105_52 (.BL(BL52),.BLN(BLN52),.WL(WL105));
sram_cell_6t_5 inst_cell_105_53 (.BL(BL53),.BLN(BLN53),.WL(WL105));
sram_cell_6t_5 inst_cell_105_54 (.BL(BL54),.BLN(BLN54),.WL(WL105));
sram_cell_6t_5 inst_cell_105_55 (.BL(BL55),.BLN(BLN55),.WL(WL105));
sram_cell_6t_5 inst_cell_105_56 (.BL(BL56),.BLN(BLN56),.WL(WL105));
sram_cell_6t_5 inst_cell_105_57 (.BL(BL57),.BLN(BLN57),.WL(WL105));
sram_cell_6t_5 inst_cell_105_58 (.BL(BL58),.BLN(BLN58),.WL(WL105));
sram_cell_6t_5 inst_cell_105_59 (.BL(BL59),.BLN(BLN59),.WL(WL105));
sram_cell_6t_5 inst_cell_105_60 (.BL(BL60),.BLN(BLN60),.WL(WL105));
sram_cell_6t_5 inst_cell_105_61 (.BL(BL61),.BLN(BLN61),.WL(WL105));
sram_cell_6t_5 inst_cell_105_62 (.BL(BL62),.BLN(BLN62),.WL(WL105));
sram_cell_6t_5 inst_cell_105_63 (.BL(BL63),.BLN(BLN63),.WL(WL105));
sram_cell_6t_5 inst_cell_105_64 (.BL(BL64),.BLN(BLN64),.WL(WL105));
sram_cell_6t_5 inst_cell_105_65 (.BL(BL65),.BLN(BLN65),.WL(WL105));
sram_cell_6t_5 inst_cell_105_66 (.BL(BL66),.BLN(BLN66),.WL(WL105));
sram_cell_6t_5 inst_cell_105_67 (.BL(BL67),.BLN(BLN67),.WL(WL105));
sram_cell_6t_5 inst_cell_105_68 (.BL(BL68),.BLN(BLN68),.WL(WL105));
sram_cell_6t_5 inst_cell_105_69 (.BL(BL69),.BLN(BLN69),.WL(WL105));
sram_cell_6t_5 inst_cell_105_70 (.BL(BL70),.BLN(BLN70),.WL(WL105));
sram_cell_6t_5 inst_cell_105_71 (.BL(BL71),.BLN(BLN71),.WL(WL105));
sram_cell_6t_5 inst_cell_105_72 (.BL(BL72),.BLN(BLN72),.WL(WL105));
sram_cell_6t_5 inst_cell_105_73 (.BL(BL73),.BLN(BLN73),.WL(WL105));
sram_cell_6t_5 inst_cell_105_74 (.BL(BL74),.BLN(BLN74),.WL(WL105));
sram_cell_6t_5 inst_cell_105_75 (.BL(BL75),.BLN(BLN75),.WL(WL105));
sram_cell_6t_5 inst_cell_105_76 (.BL(BL76),.BLN(BLN76),.WL(WL105));
sram_cell_6t_5 inst_cell_105_77 (.BL(BL77),.BLN(BLN77),.WL(WL105));
sram_cell_6t_5 inst_cell_105_78 (.BL(BL78),.BLN(BLN78),.WL(WL105));
sram_cell_6t_5 inst_cell_105_79 (.BL(BL79),.BLN(BLN79),.WL(WL105));
sram_cell_6t_5 inst_cell_105_80 (.BL(BL80),.BLN(BLN80),.WL(WL105));
sram_cell_6t_5 inst_cell_105_81 (.BL(BL81),.BLN(BLN81),.WL(WL105));
sram_cell_6t_5 inst_cell_105_82 (.BL(BL82),.BLN(BLN82),.WL(WL105));
sram_cell_6t_5 inst_cell_105_83 (.BL(BL83),.BLN(BLN83),.WL(WL105));
sram_cell_6t_5 inst_cell_105_84 (.BL(BL84),.BLN(BLN84),.WL(WL105));
sram_cell_6t_5 inst_cell_105_85 (.BL(BL85),.BLN(BLN85),.WL(WL105));
sram_cell_6t_5 inst_cell_105_86 (.BL(BL86),.BLN(BLN86),.WL(WL105));
sram_cell_6t_5 inst_cell_105_87 (.BL(BL87),.BLN(BLN87),.WL(WL105));
sram_cell_6t_5 inst_cell_105_88 (.BL(BL88),.BLN(BLN88),.WL(WL105));
sram_cell_6t_5 inst_cell_105_89 (.BL(BL89),.BLN(BLN89),.WL(WL105));
sram_cell_6t_5 inst_cell_105_90 (.BL(BL90),.BLN(BLN90),.WL(WL105));
sram_cell_6t_5 inst_cell_105_91 (.BL(BL91),.BLN(BLN91),.WL(WL105));
sram_cell_6t_5 inst_cell_105_92 (.BL(BL92),.BLN(BLN92),.WL(WL105));
sram_cell_6t_5 inst_cell_105_93 (.BL(BL93),.BLN(BLN93),.WL(WL105));
sram_cell_6t_5 inst_cell_105_94 (.BL(BL94),.BLN(BLN94),.WL(WL105));
sram_cell_6t_5 inst_cell_105_95 (.BL(BL95),.BLN(BLN95),.WL(WL105));
sram_cell_6t_5 inst_cell_105_96 (.BL(BL96),.BLN(BLN96),.WL(WL105));
sram_cell_6t_5 inst_cell_105_97 (.BL(BL97),.BLN(BLN97),.WL(WL105));
sram_cell_6t_5 inst_cell_105_98 (.BL(BL98),.BLN(BLN98),.WL(WL105));
sram_cell_6t_5 inst_cell_105_99 (.BL(BL99),.BLN(BLN99),.WL(WL105));
sram_cell_6t_5 inst_cell_105_100 (.BL(BL100),.BLN(BLN100),.WL(WL105));
sram_cell_6t_5 inst_cell_105_101 (.BL(BL101),.BLN(BLN101),.WL(WL105));
sram_cell_6t_5 inst_cell_105_102 (.BL(BL102),.BLN(BLN102),.WL(WL105));
sram_cell_6t_5 inst_cell_105_103 (.BL(BL103),.BLN(BLN103),.WL(WL105));
sram_cell_6t_5 inst_cell_105_104 (.BL(BL104),.BLN(BLN104),.WL(WL105));
sram_cell_6t_5 inst_cell_105_105 (.BL(BL105),.BLN(BLN105),.WL(WL105));
sram_cell_6t_5 inst_cell_105_106 (.BL(BL106),.BLN(BLN106),.WL(WL105));
sram_cell_6t_5 inst_cell_105_107 (.BL(BL107),.BLN(BLN107),.WL(WL105));
sram_cell_6t_5 inst_cell_105_108 (.BL(BL108),.BLN(BLN108),.WL(WL105));
sram_cell_6t_5 inst_cell_105_109 (.BL(BL109),.BLN(BLN109),.WL(WL105));
sram_cell_6t_5 inst_cell_105_110 (.BL(BL110),.BLN(BLN110),.WL(WL105));
sram_cell_6t_5 inst_cell_105_111 (.BL(BL111),.BLN(BLN111),.WL(WL105));
sram_cell_6t_5 inst_cell_105_112 (.BL(BL112),.BLN(BLN112),.WL(WL105));
sram_cell_6t_5 inst_cell_105_113 (.BL(BL113),.BLN(BLN113),.WL(WL105));
sram_cell_6t_5 inst_cell_105_114 (.BL(BL114),.BLN(BLN114),.WL(WL105));
sram_cell_6t_5 inst_cell_105_115 (.BL(BL115),.BLN(BLN115),.WL(WL105));
sram_cell_6t_5 inst_cell_105_116 (.BL(BL116),.BLN(BLN116),.WL(WL105));
sram_cell_6t_5 inst_cell_105_117 (.BL(BL117),.BLN(BLN117),.WL(WL105));
sram_cell_6t_5 inst_cell_105_118 (.BL(BL118),.BLN(BLN118),.WL(WL105));
sram_cell_6t_5 inst_cell_105_119 (.BL(BL119),.BLN(BLN119),.WL(WL105));
sram_cell_6t_5 inst_cell_105_120 (.BL(BL120),.BLN(BLN120),.WL(WL105));
sram_cell_6t_5 inst_cell_105_121 (.BL(BL121),.BLN(BLN121),.WL(WL105));
sram_cell_6t_5 inst_cell_105_122 (.BL(BL122),.BLN(BLN122),.WL(WL105));
sram_cell_6t_5 inst_cell_105_123 (.BL(BL123),.BLN(BLN123),.WL(WL105));
sram_cell_6t_5 inst_cell_105_124 (.BL(BL124),.BLN(BLN124),.WL(WL105));
sram_cell_6t_5 inst_cell_105_125 (.BL(BL125),.BLN(BLN125),.WL(WL105));
sram_cell_6t_5 inst_cell_105_126 (.BL(BL126),.BLN(BLN126),.WL(WL105));
sram_cell_6t_5 inst_cell_105_127 (.BL(BL127),.BLN(BLN127),.WL(WL105));
sram_cell_6t_5 inst_cell_106_0 (.BL(BL0),.BLN(BLN0),.WL(WL106));
sram_cell_6t_5 inst_cell_106_1 (.BL(BL1),.BLN(BLN1),.WL(WL106));
sram_cell_6t_5 inst_cell_106_2 (.BL(BL2),.BLN(BLN2),.WL(WL106));
sram_cell_6t_5 inst_cell_106_3 (.BL(BL3),.BLN(BLN3),.WL(WL106));
sram_cell_6t_5 inst_cell_106_4 (.BL(BL4),.BLN(BLN4),.WL(WL106));
sram_cell_6t_5 inst_cell_106_5 (.BL(BL5),.BLN(BLN5),.WL(WL106));
sram_cell_6t_5 inst_cell_106_6 (.BL(BL6),.BLN(BLN6),.WL(WL106));
sram_cell_6t_5 inst_cell_106_7 (.BL(BL7),.BLN(BLN7),.WL(WL106));
sram_cell_6t_5 inst_cell_106_8 (.BL(BL8),.BLN(BLN8),.WL(WL106));
sram_cell_6t_5 inst_cell_106_9 (.BL(BL9),.BLN(BLN9),.WL(WL106));
sram_cell_6t_5 inst_cell_106_10 (.BL(BL10),.BLN(BLN10),.WL(WL106));
sram_cell_6t_5 inst_cell_106_11 (.BL(BL11),.BLN(BLN11),.WL(WL106));
sram_cell_6t_5 inst_cell_106_12 (.BL(BL12),.BLN(BLN12),.WL(WL106));
sram_cell_6t_5 inst_cell_106_13 (.BL(BL13),.BLN(BLN13),.WL(WL106));
sram_cell_6t_5 inst_cell_106_14 (.BL(BL14),.BLN(BLN14),.WL(WL106));
sram_cell_6t_5 inst_cell_106_15 (.BL(BL15),.BLN(BLN15),.WL(WL106));
sram_cell_6t_5 inst_cell_106_16 (.BL(BL16),.BLN(BLN16),.WL(WL106));
sram_cell_6t_5 inst_cell_106_17 (.BL(BL17),.BLN(BLN17),.WL(WL106));
sram_cell_6t_5 inst_cell_106_18 (.BL(BL18),.BLN(BLN18),.WL(WL106));
sram_cell_6t_5 inst_cell_106_19 (.BL(BL19),.BLN(BLN19),.WL(WL106));
sram_cell_6t_5 inst_cell_106_20 (.BL(BL20),.BLN(BLN20),.WL(WL106));
sram_cell_6t_5 inst_cell_106_21 (.BL(BL21),.BLN(BLN21),.WL(WL106));
sram_cell_6t_5 inst_cell_106_22 (.BL(BL22),.BLN(BLN22),.WL(WL106));
sram_cell_6t_5 inst_cell_106_23 (.BL(BL23),.BLN(BLN23),.WL(WL106));
sram_cell_6t_5 inst_cell_106_24 (.BL(BL24),.BLN(BLN24),.WL(WL106));
sram_cell_6t_5 inst_cell_106_25 (.BL(BL25),.BLN(BLN25),.WL(WL106));
sram_cell_6t_5 inst_cell_106_26 (.BL(BL26),.BLN(BLN26),.WL(WL106));
sram_cell_6t_5 inst_cell_106_27 (.BL(BL27),.BLN(BLN27),.WL(WL106));
sram_cell_6t_5 inst_cell_106_28 (.BL(BL28),.BLN(BLN28),.WL(WL106));
sram_cell_6t_5 inst_cell_106_29 (.BL(BL29),.BLN(BLN29),.WL(WL106));
sram_cell_6t_5 inst_cell_106_30 (.BL(BL30),.BLN(BLN30),.WL(WL106));
sram_cell_6t_5 inst_cell_106_31 (.BL(BL31),.BLN(BLN31),.WL(WL106));
sram_cell_6t_5 inst_cell_106_32 (.BL(BL32),.BLN(BLN32),.WL(WL106));
sram_cell_6t_5 inst_cell_106_33 (.BL(BL33),.BLN(BLN33),.WL(WL106));
sram_cell_6t_5 inst_cell_106_34 (.BL(BL34),.BLN(BLN34),.WL(WL106));
sram_cell_6t_5 inst_cell_106_35 (.BL(BL35),.BLN(BLN35),.WL(WL106));
sram_cell_6t_5 inst_cell_106_36 (.BL(BL36),.BLN(BLN36),.WL(WL106));
sram_cell_6t_5 inst_cell_106_37 (.BL(BL37),.BLN(BLN37),.WL(WL106));
sram_cell_6t_5 inst_cell_106_38 (.BL(BL38),.BLN(BLN38),.WL(WL106));
sram_cell_6t_5 inst_cell_106_39 (.BL(BL39),.BLN(BLN39),.WL(WL106));
sram_cell_6t_5 inst_cell_106_40 (.BL(BL40),.BLN(BLN40),.WL(WL106));
sram_cell_6t_5 inst_cell_106_41 (.BL(BL41),.BLN(BLN41),.WL(WL106));
sram_cell_6t_5 inst_cell_106_42 (.BL(BL42),.BLN(BLN42),.WL(WL106));
sram_cell_6t_5 inst_cell_106_43 (.BL(BL43),.BLN(BLN43),.WL(WL106));
sram_cell_6t_5 inst_cell_106_44 (.BL(BL44),.BLN(BLN44),.WL(WL106));
sram_cell_6t_5 inst_cell_106_45 (.BL(BL45),.BLN(BLN45),.WL(WL106));
sram_cell_6t_5 inst_cell_106_46 (.BL(BL46),.BLN(BLN46),.WL(WL106));
sram_cell_6t_5 inst_cell_106_47 (.BL(BL47),.BLN(BLN47),.WL(WL106));
sram_cell_6t_5 inst_cell_106_48 (.BL(BL48),.BLN(BLN48),.WL(WL106));
sram_cell_6t_5 inst_cell_106_49 (.BL(BL49),.BLN(BLN49),.WL(WL106));
sram_cell_6t_5 inst_cell_106_50 (.BL(BL50),.BLN(BLN50),.WL(WL106));
sram_cell_6t_5 inst_cell_106_51 (.BL(BL51),.BLN(BLN51),.WL(WL106));
sram_cell_6t_5 inst_cell_106_52 (.BL(BL52),.BLN(BLN52),.WL(WL106));
sram_cell_6t_5 inst_cell_106_53 (.BL(BL53),.BLN(BLN53),.WL(WL106));
sram_cell_6t_5 inst_cell_106_54 (.BL(BL54),.BLN(BLN54),.WL(WL106));
sram_cell_6t_5 inst_cell_106_55 (.BL(BL55),.BLN(BLN55),.WL(WL106));
sram_cell_6t_5 inst_cell_106_56 (.BL(BL56),.BLN(BLN56),.WL(WL106));
sram_cell_6t_5 inst_cell_106_57 (.BL(BL57),.BLN(BLN57),.WL(WL106));
sram_cell_6t_5 inst_cell_106_58 (.BL(BL58),.BLN(BLN58),.WL(WL106));
sram_cell_6t_5 inst_cell_106_59 (.BL(BL59),.BLN(BLN59),.WL(WL106));
sram_cell_6t_5 inst_cell_106_60 (.BL(BL60),.BLN(BLN60),.WL(WL106));
sram_cell_6t_5 inst_cell_106_61 (.BL(BL61),.BLN(BLN61),.WL(WL106));
sram_cell_6t_5 inst_cell_106_62 (.BL(BL62),.BLN(BLN62),.WL(WL106));
sram_cell_6t_5 inst_cell_106_63 (.BL(BL63),.BLN(BLN63),.WL(WL106));
sram_cell_6t_5 inst_cell_106_64 (.BL(BL64),.BLN(BLN64),.WL(WL106));
sram_cell_6t_5 inst_cell_106_65 (.BL(BL65),.BLN(BLN65),.WL(WL106));
sram_cell_6t_5 inst_cell_106_66 (.BL(BL66),.BLN(BLN66),.WL(WL106));
sram_cell_6t_5 inst_cell_106_67 (.BL(BL67),.BLN(BLN67),.WL(WL106));
sram_cell_6t_5 inst_cell_106_68 (.BL(BL68),.BLN(BLN68),.WL(WL106));
sram_cell_6t_5 inst_cell_106_69 (.BL(BL69),.BLN(BLN69),.WL(WL106));
sram_cell_6t_5 inst_cell_106_70 (.BL(BL70),.BLN(BLN70),.WL(WL106));
sram_cell_6t_5 inst_cell_106_71 (.BL(BL71),.BLN(BLN71),.WL(WL106));
sram_cell_6t_5 inst_cell_106_72 (.BL(BL72),.BLN(BLN72),.WL(WL106));
sram_cell_6t_5 inst_cell_106_73 (.BL(BL73),.BLN(BLN73),.WL(WL106));
sram_cell_6t_5 inst_cell_106_74 (.BL(BL74),.BLN(BLN74),.WL(WL106));
sram_cell_6t_5 inst_cell_106_75 (.BL(BL75),.BLN(BLN75),.WL(WL106));
sram_cell_6t_5 inst_cell_106_76 (.BL(BL76),.BLN(BLN76),.WL(WL106));
sram_cell_6t_5 inst_cell_106_77 (.BL(BL77),.BLN(BLN77),.WL(WL106));
sram_cell_6t_5 inst_cell_106_78 (.BL(BL78),.BLN(BLN78),.WL(WL106));
sram_cell_6t_5 inst_cell_106_79 (.BL(BL79),.BLN(BLN79),.WL(WL106));
sram_cell_6t_5 inst_cell_106_80 (.BL(BL80),.BLN(BLN80),.WL(WL106));
sram_cell_6t_5 inst_cell_106_81 (.BL(BL81),.BLN(BLN81),.WL(WL106));
sram_cell_6t_5 inst_cell_106_82 (.BL(BL82),.BLN(BLN82),.WL(WL106));
sram_cell_6t_5 inst_cell_106_83 (.BL(BL83),.BLN(BLN83),.WL(WL106));
sram_cell_6t_5 inst_cell_106_84 (.BL(BL84),.BLN(BLN84),.WL(WL106));
sram_cell_6t_5 inst_cell_106_85 (.BL(BL85),.BLN(BLN85),.WL(WL106));
sram_cell_6t_5 inst_cell_106_86 (.BL(BL86),.BLN(BLN86),.WL(WL106));
sram_cell_6t_5 inst_cell_106_87 (.BL(BL87),.BLN(BLN87),.WL(WL106));
sram_cell_6t_5 inst_cell_106_88 (.BL(BL88),.BLN(BLN88),.WL(WL106));
sram_cell_6t_5 inst_cell_106_89 (.BL(BL89),.BLN(BLN89),.WL(WL106));
sram_cell_6t_5 inst_cell_106_90 (.BL(BL90),.BLN(BLN90),.WL(WL106));
sram_cell_6t_5 inst_cell_106_91 (.BL(BL91),.BLN(BLN91),.WL(WL106));
sram_cell_6t_5 inst_cell_106_92 (.BL(BL92),.BLN(BLN92),.WL(WL106));
sram_cell_6t_5 inst_cell_106_93 (.BL(BL93),.BLN(BLN93),.WL(WL106));
sram_cell_6t_5 inst_cell_106_94 (.BL(BL94),.BLN(BLN94),.WL(WL106));
sram_cell_6t_5 inst_cell_106_95 (.BL(BL95),.BLN(BLN95),.WL(WL106));
sram_cell_6t_5 inst_cell_106_96 (.BL(BL96),.BLN(BLN96),.WL(WL106));
sram_cell_6t_5 inst_cell_106_97 (.BL(BL97),.BLN(BLN97),.WL(WL106));
sram_cell_6t_5 inst_cell_106_98 (.BL(BL98),.BLN(BLN98),.WL(WL106));
sram_cell_6t_5 inst_cell_106_99 (.BL(BL99),.BLN(BLN99),.WL(WL106));
sram_cell_6t_5 inst_cell_106_100 (.BL(BL100),.BLN(BLN100),.WL(WL106));
sram_cell_6t_5 inst_cell_106_101 (.BL(BL101),.BLN(BLN101),.WL(WL106));
sram_cell_6t_5 inst_cell_106_102 (.BL(BL102),.BLN(BLN102),.WL(WL106));
sram_cell_6t_5 inst_cell_106_103 (.BL(BL103),.BLN(BLN103),.WL(WL106));
sram_cell_6t_5 inst_cell_106_104 (.BL(BL104),.BLN(BLN104),.WL(WL106));
sram_cell_6t_5 inst_cell_106_105 (.BL(BL105),.BLN(BLN105),.WL(WL106));
sram_cell_6t_5 inst_cell_106_106 (.BL(BL106),.BLN(BLN106),.WL(WL106));
sram_cell_6t_5 inst_cell_106_107 (.BL(BL107),.BLN(BLN107),.WL(WL106));
sram_cell_6t_5 inst_cell_106_108 (.BL(BL108),.BLN(BLN108),.WL(WL106));
sram_cell_6t_5 inst_cell_106_109 (.BL(BL109),.BLN(BLN109),.WL(WL106));
sram_cell_6t_5 inst_cell_106_110 (.BL(BL110),.BLN(BLN110),.WL(WL106));
sram_cell_6t_5 inst_cell_106_111 (.BL(BL111),.BLN(BLN111),.WL(WL106));
sram_cell_6t_5 inst_cell_106_112 (.BL(BL112),.BLN(BLN112),.WL(WL106));
sram_cell_6t_5 inst_cell_106_113 (.BL(BL113),.BLN(BLN113),.WL(WL106));
sram_cell_6t_5 inst_cell_106_114 (.BL(BL114),.BLN(BLN114),.WL(WL106));
sram_cell_6t_5 inst_cell_106_115 (.BL(BL115),.BLN(BLN115),.WL(WL106));
sram_cell_6t_5 inst_cell_106_116 (.BL(BL116),.BLN(BLN116),.WL(WL106));
sram_cell_6t_5 inst_cell_106_117 (.BL(BL117),.BLN(BLN117),.WL(WL106));
sram_cell_6t_5 inst_cell_106_118 (.BL(BL118),.BLN(BLN118),.WL(WL106));
sram_cell_6t_5 inst_cell_106_119 (.BL(BL119),.BLN(BLN119),.WL(WL106));
sram_cell_6t_5 inst_cell_106_120 (.BL(BL120),.BLN(BLN120),.WL(WL106));
sram_cell_6t_5 inst_cell_106_121 (.BL(BL121),.BLN(BLN121),.WL(WL106));
sram_cell_6t_5 inst_cell_106_122 (.BL(BL122),.BLN(BLN122),.WL(WL106));
sram_cell_6t_5 inst_cell_106_123 (.BL(BL123),.BLN(BLN123),.WL(WL106));
sram_cell_6t_5 inst_cell_106_124 (.BL(BL124),.BLN(BLN124),.WL(WL106));
sram_cell_6t_5 inst_cell_106_125 (.BL(BL125),.BLN(BLN125),.WL(WL106));
sram_cell_6t_5 inst_cell_106_126 (.BL(BL126),.BLN(BLN126),.WL(WL106));
sram_cell_6t_5 inst_cell_106_127 (.BL(BL127),.BLN(BLN127),.WL(WL106));
sram_cell_6t_5 inst_cell_107_0 (.BL(BL0),.BLN(BLN0),.WL(WL107));
sram_cell_6t_5 inst_cell_107_1 (.BL(BL1),.BLN(BLN1),.WL(WL107));
sram_cell_6t_5 inst_cell_107_2 (.BL(BL2),.BLN(BLN2),.WL(WL107));
sram_cell_6t_5 inst_cell_107_3 (.BL(BL3),.BLN(BLN3),.WL(WL107));
sram_cell_6t_5 inst_cell_107_4 (.BL(BL4),.BLN(BLN4),.WL(WL107));
sram_cell_6t_5 inst_cell_107_5 (.BL(BL5),.BLN(BLN5),.WL(WL107));
sram_cell_6t_5 inst_cell_107_6 (.BL(BL6),.BLN(BLN6),.WL(WL107));
sram_cell_6t_5 inst_cell_107_7 (.BL(BL7),.BLN(BLN7),.WL(WL107));
sram_cell_6t_5 inst_cell_107_8 (.BL(BL8),.BLN(BLN8),.WL(WL107));
sram_cell_6t_5 inst_cell_107_9 (.BL(BL9),.BLN(BLN9),.WL(WL107));
sram_cell_6t_5 inst_cell_107_10 (.BL(BL10),.BLN(BLN10),.WL(WL107));
sram_cell_6t_5 inst_cell_107_11 (.BL(BL11),.BLN(BLN11),.WL(WL107));
sram_cell_6t_5 inst_cell_107_12 (.BL(BL12),.BLN(BLN12),.WL(WL107));
sram_cell_6t_5 inst_cell_107_13 (.BL(BL13),.BLN(BLN13),.WL(WL107));
sram_cell_6t_5 inst_cell_107_14 (.BL(BL14),.BLN(BLN14),.WL(WL107));
sram_cell_6t_5 inst_cell_107_15 (.BL(BL15),.BLN(BLN15),.WL(WL107));
sram_cell_6t_5 inst_cell_107_16 (.BL(BL16),.BLN(BLN16),.WL(WL107));
sram_cell_6t_5 inst_cell_107_17 (.BL(BL17),.BLN(BLN17),.WL(WL107));
sram_cell_6t_5 inst_cell_107_18 (.BL(BL18),.BLN(BLN18),.WL(WL107));
sram_cell_6t_5 inst_cell_107_19 (.BL(BL19),.BLN(BLN19),.WL(WL107));
sram_cell_6t_5 inst_cell_107_20 (.BL(BL20),.BLN(BLN20),.WL(WL107));
sram_cell_6t_5 inst_cell_107_21 (.BL(BL21),.BLN(BLN21),.WL(WL107));
sram_cell_6t_5 inst_cell_107_22 (.BL(BL22),.BLN(BLN22),.WL(WL107));
sram_cell_6t_5 inst_cell_107_23 (.BL(BL23),.BLN(BLN23),.WL(WL107));
sram_cell_6t_5 inst_cell_107_24 (.BL(BL24),.BLN(BLN24),.WL(WL107));
sram_cell_6t_5 inst_cell_107_25 (.BL(BL25),.BLN(BLN25),.WL(WL107));
sram_cell_6t_5 inst_cell_107_26 (.BL(BL26),.BLN(BLN26),.WL(WL107));
sram_cell_6t_5 inst_cell_107_27 (.BL(BL27),.BLN(BLN27),.WL(WL107));
sram_cell_6t_5 inst_cell_107_28 (.BL(BL28),.BLN(BLN28),.WL(WL107));
sram_cell_6t_5 inst_cell_107_29 (.BL(BL29),.BLN(BLN29),.WL(WL107));
sram_cell_6t_5 inst_cell_107_30 (.BL(BL30),.BLN(BLN30),.WL(WL107));
sram_cell_6t_5 inst_cell_107_31 (.BL(BL31),.BLN(BLN31),.WL(WL107));
sram_cell_6t_5 inst_cell_107_32 (.BL(BL32),.BLN(BLN32),.WL(WL107));
sram_cell_6t_5 inst_cell_107_33 (.BL(BL33),.BLN(BLN33),.WL(WL107));
sram_cell_6t_5 inst_cell_107_34 (.BL(BL34),.BLN(BLN34),.WL(WL107));
sram_cell_6t_5 inst_cell_107_35 (.BL(BL35),.BLN(BLN35),.WL(WL107));
sram_cell_6t_5 inst_cell_107_36 (.BL(BL36),.BLN(BLN36),.WL(WL107));
sram_cell_6t_5 inst_cell_107_37 (.BL(BL37),.BLN(BLN37),.WL(WL107));
sram_cell_6t_5 inst_cell_107_38 (.BL(BL38),.BLN(BLN38),.WL(WL107));
sram_cell_6t_5 inst_cell_107_39 (.BL(BL39),.BLN(BLN39),.WL(WL107));
sram_cell_6t_5 inst_cell_107_40 (.BL(BL40),.BLN(BLN40),.WL(WL107));
sram_cell_6t_5 inst_cell_107_41 (.BL(BL41),.BLN(BLN41),.WL(WL107));
sram_cell_6t_5 inst_cell_107_42 (.BL(BL42),.BLN(BLN42),.WL(WL107));
sram_cell_6t_5 inst_cell_107_43 (.BL(BL43),.BLN(BLN43),.WL(WL107));
sram_cell_6t_5 inst_cell_107_44 (.BL(BL44),.BLN(BLN44),.WL(WL107));
sram_cell_6t_5 inst_cell_107_45 (.BL(BL45),.BLN(BLN45),.WL(WL107));
sram_cell_6t_5 inst_cell_107_46 (.BL(BL46),.BLN(BLN46),.WL(WL107));
sram_cell_6t_5 inst_cell_107_47 (.BL(BL47),.BLN(BLN47),.WL(WL107));
sram_cell_6t_5 inst_cell_107_48 (.BL(BL48),.BLN(BLN48),.WL(WL107));
sram_cell_6t_5 inst_cell_107_49 (.BL(BL49),.BLN(BLN49),.WL(WL107));
sram_cell_6t_5 inst_cell_107_50 (.BL(BL50),.BLN(BLN50),.WL(WL107));
sram_cell_6t_5 inst_cell_107_51 (.BL(BL51),.BLN(BLN51),.WL(WL107));
sram_cell_6t_5 inst_cell_107_52 (.BL(BL52),.BLN(BLN52),.WL(WL107));
sram_cell_6t_5 inst_cell_107_53 (.BL(BL53),.BLN(BLN53),.WL(WL107));
sram_cell_6t_5 inst_cell_107_54 (.BL(BL54),.BLN(BLN54),.WL(WL107));
sram_cell_6t_5 inst_cell_107_55 (.BL(BL55),.BLN(BLN55),.WL(WL107));
sram_cell_6t_5 inst_cell_107_56 (.BL(BL56),.BLN(BLN56),.WL(WL107));
sram_cell_6t_5 inst_cell_107_57 (.BL(BL57),.BLN(BLN57),.WL(WL107));
sram_cell_6t_5 inst_cell_107_58 (.BL(BL58),.BLN(BLN58),.WL(WL107));
sram_cell_6t_5 inst_cell_107_59 (.BL(BL59),.BLN(BLN59),.WL(WL107));
sram_cell_6t_5 inst_cell_107_60 (.BL(BL60),.BLN(BLN60),.WL(WL107));
sram_cell_6t_5 inst_cell_107_61 (.BL(BL61),.BLN(BLN61),.WL(WL107));
sram_cell_6t_5 inst_cell_107_62 (.BL(BL62),.BLN(BLN62),.WL(WL107));
sram_cell_6t_5 inst_cell_107_63 (.BL(BL63),.BLN(BLN63),.WL(WL107));
sram_cell_6t_5 inst_cell_107_64 (.BL(BL64),.BLN(BLN64),.WL(WL107));
sram_cell_6t_5 inst_cell_107_65 (.BL(BL65),.BLN(BLN65),.WL(WL107));
sram_cell_6t_5 inst_cell_107_66 (.BL(BL66),.BLN(BLN66),.WL(WL107));
sram_cell_6t_5 inst_cell_107_67 (.BL(BL67),.BLN(BLN67),.WL(WL107));
sram_cell_6t_5 inst_cell_107_68 (.BL(BL68),.BLN(BLN68),.WL(WL107));
sram_cell_6t_5 inst_cell_107_69 (.BL(BL69),.BLN(BLN69),.WL(WL107));
sram_cell_6t_5 inst_cell_107_70 (.BL(BL70),.BLN(BLN70),.WL(WL107));
sram_cell_6t_5 inst_cell_107_71 (.BL(BL71),.BLN(BLN71),.WL(WL107));
sram_cell_6t_5 inst_cell_107_72 (.BL(BL72),.BLN(BLN72),.WL(WL107));
sram_cell_6t_5 inst_cell_107_73 (.BL(BL73),.BLN(BLN73),.WL(WL107));
sram_cell_6t_5 inst_cell_107_74 (.BL(BL74),.BLN(BLN74),.WL(WL107));
sram_cell_6t_5 inst_cell_107_75 (.BL(BL75),.BLN(BLN75),.WL(WL107));
sram_cell_6t_5 inst_cell_107_76 (.BL(BL76),.BLN(BLN76),.WL(WL107));
sram_cell_6t_5 inst_cell_107_77 (.BL(BL77),.BLN(BLN77),.WL(WL107));
sram_cell_6t_5 inst_cell_107_78 (.BL(BL78),.BLN(BLN78),.WL(WL107));
sram_cell_6t_5 inst_cell_107_79 (.BL(BL79),.BLN(BLN79),.WL(WL107));
sram_cell_6t_5 inst_cell_107_80 (.BL(BL80),.BLN(BLN80),.WL(WL107));
sram_cell_6t_5 inst_cell_107_81 (.BL(BL81),.BLN(BLN81),.WL(WL107));
sram_cell_6t_5 inst_cell_107_82 (.BL(BL82),.BLN(BLN82),.WL(WL107));
sram_cell_6t_5 inst_cell_107_83 (.BL(BL83),.BLN(BLN83),.WL(WL107));
sram_cell_6t_5 inst_cell_107_84 (.BL(BL84),.BLN(BLN84),.WL(WL107));
sram_cell_6t_5 inst_cell_107_85 (.BL(BL85),.BLN(BLN85),.WL(WL107));
sram_cell_6t_5 inst_cell_107_86 (.BL(BL86),.BLN(BLN86),.WL(WL107));
sram_cell_6t_5 inst_cell_107_87 (.BL(BL87),.BLN(BLN87),.WL(WL107));
sram_cell_6t_5 inst_cell_107_88 (.BL(BL88),.BLN(BLN88),.WL(WL107));
sram_cell_6t_5 inst_cell_107_89 (.BL(BL89),.BLN(BLN89),.WL(WL107));
sram_cell_6t_5 inst_cell_107_90 (.BL(BL90),.BLN(BLN90),.WL(WL107));
sram_cell_6t_5 inst_cell_107_91 (.BL(BL91),.BLN(BLN91),.WL(WL107));
sram_cell_6t_5 inst_cell_107_92 (.BL(BL92),.BLN(BLN92),.WL(WL107));
sram_cell_6t_5 inst_cell_107_93 (.BL(BL93),.BLN(BLN93),.WL(WL107));
sram_cell_6t_5 inst_cell_107_94 (.BL(BL94),.BLN(BLN94),.WL(WL107));
sram_cell_6t_5 inst_cell_107_95 (.BL(BL95),.BLN(BLN95),.WL(WL107));
sram_cell_6t_5 inst_cell_107_96 (.BL(BL96),.BLN(BLN96),.WL(WL107));
sram_cell_6t_5 inst_cell_107_97 (.BL(BL97),.BLN(BLN97),.WL(WL107));
sram_cell_6t_5 inst_cell_107_98 (.BL(BL98),.BLN(BLN98),.WL(WL107));
sram_cell_6t_5 inst_cell_107_99 (.BL(BL99),.BLN(BLN99),.WL(WL107));
sram_cell_6t_5 inst_cell_107_100 (.BL(BL100),.BLN(BLN100),.WL(WL107));
sram_cell_6t_5 inst_cell_107_101 (.BL(BL101),.BLN(BLN101),.WL(WL107));
sram_cell_6t_5 inst_cell_107_102 (.BL(BL102),.BLN(BLN102),.WL(WL107));
sram_cell_6t_5 inst_cell_107_103 (.BL(BL103),.BLN(BLN103),.WL(WL107));
sram_cell_6t_5 inst_cell_107_104 (.BL(BL104),.BLN(BLN104),.WL(WL107));
sram_cell_6t_5 inst_cell_107_105 (.BL(BL105),.BLN(BLN105),.WL(WL107));
sram_cell_6t_5 inst_cell_107_106 (.BL(BL106),.BLN(BLN106),.WL(WL107));
sram_cell_6t_5 inst_cell_107_107 (.BL(BL107),.BLN(BLN107),.WL(WL107));
sram_cell_6t_5 inst_cell_107_108 (.BL(BL108),.BLN(BLN108),.WL(WL107));
sram_cell_6t_5 inst_cell_107_109 (.BL(BL109),.BLN(BLN109),.WL(WL107));
sram_cell_6t_5 inst_cell_107_110 (.BL(BL110),.BLN(BLN110),.WL(WL107));
sram_cell_6t_5 inst_cell_107_111 (.BL(BL111),.BLN(BLN111),.WL(WL107));
sram_cell_6t_5 inst_cell_107_112 (.BL(BL112),.BLN(BLN112),.WL(WL107));
sram_cell_6t_5 inst_cell_107_113 (.BL(BL113),.BLN(BLN113),.WL(WL107));
sram_cell_6t_5 inst_cell_107_114 (.BL(BL114),.BLN(BLN114),.WL(WL107));
sram_cell_6t_5 inst_cell_107_115 (.BL(BL115),.BLN(BLN115),.WL(WL107));
sram_cell_6t_5 inst_cell_107_116 (.BL(BL116),.BLN(BLN116),.WL(WL107));
sram_cell_6t_5 inst_cell_107_117 (.BL(BL117),.BLN(BLN117),.WL(WL107));
sram_cell_6t_5 inst_cell_107_118 (.BL(BL118),.BLN(BLN118),.WL(WL107));
sram_cell_6t_5 inst_cell_107_119 (.BL(BL119),.BLN(BLN119),.WL(WL107));
sram_cell_6t_5 inst_cell_107_120 (.BL(BL120),.BLN(BLN120),.WL(WL107));
sram_cell_6t_5 inst_cell_107_121 (.BL(BL121),.BLN(BLN121),.WL(WL107));
sram_cell_6t_5 inst_cell_107_122 (.BL(BL122),.BLN(BLN122),.WL(WL107));
sram_cell_6t_5 inst_cell_107_123 (.BL(BL123),.BLN(BLN123),.WL(WL107));
sram_cell_6t_5 inst_cell_107_124 (.BL(BL124),.BLN(BLN124),.WL(WL107));
sram_cell_6t_5 inst_cell_107_125 (.BL(BL125),.BLN(BLN125),.WL(WL107));
sram_cell_6t_5 inst_cell_107_126 (.BL(BL126),.BLN(BLN126),.WL(WL107));
sram_cell_6t_5 inst_cell_107_127 (.BL(BL127),.BLN(BLN127),.WL(WL107));
sram_cell_6t_5 inst_cell_108_0 (.BL(BL0),.BLN(BLN0),.WL(WL108));
sram_cell_6t_5 inst_cell_108_1 (.BL(BL1),.BLN(BLN1),.WL(WL108));
sram_cell_6t_5 inst_cell_108_2 (.BL(BL2),.BLN(BLN2),.WL(WL108));
sram_cell_6t_5 inst_cell_108_3 (.BL(BL3),.BLN(BLN3),.WL(WL108));
sram_cell_6t_5 inst_cell_108_4 (.BL(BL4),.BLN(BLN4),.WL(WL108));
sram_cell_6t_5 inst_cell_108_5 (.BL(BL5),.BLN(BLN5),.WL(WL108));
sram_cell_6t_5 inst_cell_108_6 (.BL(BL6),.BLN(BLN6),.WL(WL108));
sram_cell_6t_5 inst_cell_108_7 (.BL(BL7),.BLN(BLN7),.WL(WL108));
sram_cell_6t_5 inst_cell_108_8 (.BL(BL8),.BLN(BLN8),.WL(WL108));
sram_cell_6t_5 inst_cell_108_9 (.BL(BL9),.BLN(BLN9),.WL(WL108));
sram_cell_6t_5 inst_cell_108_10 (.BL(BL10),.BLN(BLN10),.WL(WL108));
sram_cell_6t_5 inst_cell_108_11 (.BL(BL11),.BLN(BLN11),.WL(WL108));
sram_cell_6t_5 inst_cell_108_12 (.BL(BL12),.BLN(BLN12),.WL(WL108));
sram_cell_6t_5 inst_cell_108_13 (.BL(BL13),.BLN(BLN13),.WL(WL108));
sram_cell_6t_5 inst_cell_108_14 (.BL(BL14),.BLN(BLN14),.WL(WL108));
sram_cell_6t_5 inst_cell_108_15 (.BL(BL15),.BLN(BLN15),.WL(WL108));
sram_cell_6t_5 inst_cell_108_16 (.BL(BL16),.BLN(BLN16),.WL(WL108));
sram_cell_6t_5 inst_cell_108_17 (.BL(BL17),.BLN(BLN17),.WL(WL108));
sram_cell_6t_5 inst_cell_108_18 (.BL(BL18),.BLN(BLN18),.WL(WL108));
sram_cell_6t_5 inst_cell_108_19 (.BL(BL19),.BLN(BLN19),.WL(WL108));
sram_cell_6t_5 inst_cell_108_20 (.BL(BL20),.BLN(BLN20),.WL(WL108));
sram_cell_6t_5 inst_cell_108_21 (.BL(BL21),.BLN(BLN21),.WL(WL108));
sram_cell_6t_5 inst_cell_108_22 (.BL(BL22),.BLN(BLN22),.WL(WL108));
sram_cell_6t_5 inst_cell_108_23 (.BL(BL23),.BLN(BLN23),.WL(WL108));
sram_cell_6t_5 inst_cell_108_24 (.BL(BL24),.BLN(BLN24),.WL(WL108));
sram_cell_6t_5 inst_cell_108_25 (.BL(BL25),.BLN(BLN25),.WL(WL108));
sram_cell_6t_5 inst_cell_108_26 (.BL(BL26),.BLN(BLN26),.WL(WL108));
sram_cell_6t_5 inst_cell_108_27 (.BL(BL27),.BLN(BLN27),.WL(WL108));
sram_cell_6t_5 inst_cell_108_28 (.BL(BL28),.BLN(BLN28),.WL(WL108));
sram_cell_6t_5 inst_cell_108_29 (.BL(BL29),.BLN(BLN29),.WL(WL108));
sram_cell_6t_5 inst_cell_108_30 (.BL(BL30),.BLN(BLN30),.WL(WL108));
sram_cell_6t_5 inst_cell_108_31 (.BL(BL31),.BLN(BLN31),.WL(WL108));
sram_cell_6t_5 inst_cell_108_32 (.BL(BL32),.BLN(BLN32),.WL(WL108));
sram_cell_6t_5 inst_cell_108_33 (.BL(BL33),.BLN(BLN33),.WL(WL108));
sram_cell_6t_5 inst_cell_108_34 (.BL(BL34),.BLN(BLN34),.WL(WL108));
sram_cell_6t_5 inst_cell_108_35 (.BL(BL35),.BLN(BLN35),.WL(WL108));
sram_cell_6t_5 inst_cell_108_36 (.BL(BL36),.BLN(BLN36),.WL(WL108));
sram_cell_6t_5 inst_cell_108_37 (.BL(BL37),.BLN(BLN37),.WL(WL108));
sram_cell_6t_5 inst_cell_108_38 (.BL(BL38),.BLN(BLN38),.WL(WL108));
sram_cell_6t_5 inst_cell_108_39 (.BL(BL39),.BLN(BLN39),.WL(WL108));
sram_cell_6t_5 inst_cell_108_40 (.BL(BL40),.BLN(BLN40),.WL(WL108));
sram_cell_6t_5 inst_cell_108_41 (.BL(BL41),.BLN(BLN41),.WL(WL108));
sram_cell_6t_5 inst_cell_108_42 (.BL(BL42),.BLN(BLN42),.WL(WL108));
sram_cell_6t_5 inst_cell_108_43 (.BL(BL43),.BLN(BLN43),.WL(WL108));
sram_cell_6t_5 inst_cell_108_44 (.BL(BL44),.BLN(BLN44),.WL(WL108));
sram_cell_6t_5 inst_cell_108_45 (.BL(BL45),.BLN(BLN45),.WL(WL108));
sram_cell_6t_5 inst_cell_108_46 (.BL(BL46),.BLN(BLN46),.WL(WL108));
sram_cell_6t_5 inst_cell_108_47 (.BL(BL47),.BLN(BLN47),.WL(WL108));
sram_cell_6t_5 inst_cell_108_48 (.BL(BL48),.BLN(BLN48),.WL(WL108));
sram_cell_6t_5 inst_cell_108_49 (.BL(BL49),.BLN(BLN49),.WL(WL108));
sram_cell_6t_5 inst_cell_108_50 (.BL(BL50),.BLN(BLN50),.WL(WL108));
sram_cell_6t_5 inst_cell_108_51 (.BL(BL51),.BLN(BLN51),.WL(WL108));
sram_cell_6t_5 inst_cell_108_52 (.BL(BL52),.BLN(BLN52),.WL(WL108));
sram_cell_6t_5 inst_cell_108_53 (.BL(BL53),.BLN(BLN53),.WL(WL108));
sram_cell_6t_5 inst_cell_108_54 (.BL(BL54),.BLN(BLN54),.WL(WL108));
sram_cell_6t_5 inst_cell_108_55 (.BL(BL55),.BLN(BLN55),.WL(WL108));
sram_cell_6t_5 inst_cell_108_56 (.BL(BL56),.BLN(BLN56),.WL(WL108));
sram_cell_6t_5 inst_cell_108_57 (.BL(BL57),.BLN(BLN57),.WL(WL108));
sram_cell_6t_5 inst_cell_108_58 (.BL(BL58),.BLN(BLN58),.WL(WL108));
sram_cell_6t_5 inst_cell_108_59 (.BL(BL59),.BLN(BLN59),.WL(WL108));
sram_cell_6t_5 inst_cell_108_60 (.BL(BL60),.BLN(BLN60),.WL(WL108));
sram_cell_6t_5 inst_cell_108_61 (.BL(BL61),.BLN(BLN61),.WL(WL108));
sram_cell_6t_5 inst_cell_108_62 (.BL(BL62),.BLN(BLN62),.WL(WL108));
sram_cell_6t_5 inst_cell_108_63 (.BL(BL63),.BLN(BLN63),.WL(WL108));
sram_cell_6t_5 inst_cell_108_64 (.BL(BL64),.BLN(BLN64),.WL(WL108));
sram_cell_6t_5 inst_cell_108_65 (.BL(BL65),.BLN(BLN65),.WL(WL108));
sram_cell_6t_5 inst_cell_108_66 (.BL(BL66),.BLN(BLN66),.WL(WL108));
sram_cell_6t_5 inst_cell_108_67 (.BL(BL67),.BLN(BLN67),.WL(WL108));
sram_cell_6t_5 inst_cell_108_68 (.BL(BL68),.BLN(BLN68),.WL(WL108));
sram_cell_6t_5 inst_cell_108_69 (.BL(BL69),.BLN(BLN69),.WL(WL108));
sram_cell_6t_5 inst_cell_108_70 (.BL(BL70),.BLN(BLN70),.WL(WL108));
sram_cell_6t_5 inst_cell_108_71 (.BL(BL71),.BLN(BLN71),.WL(WL108));
sram_cell_6t_5 inst_cell_108_72 (.BL(BL72),.BLN(BLN72),.WL(WL108));
sram_cell_6t_5 inst_cell_108_73 (.BL(BL73),.BLN(BLN73),.WL(WL108));
sram_cell_6t_5 inst_cell_108_74 (.BL(BL74),.BLN(BLN74),.WL(WL108));
sram_cell_6t_5 inst_cell_108_75 (.BL(BL75),.BLN(BLN75),.WL(WL108));
sram_cell_6t_5 inst_cell_108_76 (.BL(BL76),.BLN(BLN76),.WL(WL108));
sram_cell_6t_5 inst_cell_108_77 (.BL(BL77),.BLN(BLN77),.WL(WL108));
sram_cell_6t_5 inst_cell_108_78 (.BL(BL78),.BLN(BLN78),.WL(WL108));
sram_cell_6t_5 inst_cell_108_79 (.BL(BL79),.BLN(BLN79),.WL(WL108));
sram_cell_6t_5 inst_cell_108_80 (.BL(BL80),.BLN(BLN80),.WL(WL108));
sram_cell_6t_5 inst_cell_108_81 (.BL(BL81),.BLN(BLN81),.WL(WL108));
sram_cell_6t_5 inst_cell_108_82 (.BL(BL82),.BLN(BLN82),.WL(WL108));
sram_cell_6t_5 inst_cell_108_83 (.BL(BL83),.BLN(BLN83),.WL(WL108));
sram_cell_6t_5 inst_cell_108_84 (.BL(BL84),.BLN(BLN84),.WL(WL108));
sram_cell_6t_5 inst_cell_108_85 (.BL(BL85),.BLN(BLN85),.WL(WL108));
sram_cell_6t_5 inst_cell_108_86 (.BL(BL86),.BLN(BLN86),.WL(WL108));
sram_cell_6t_5 inst_cell_108_87 (.BL(BL87),.BLN(BLN87),.WL(WL108));
sram_cell_6t_5 inst_cell_108_88 (.BL(BL88),.BLN(BLN88),.WL(WL108));
sram_cell_6t_5 inst_cell_108_89 (.BL(BL89),.BLN(BLN89),.WL(WL108));
sram_cell_6t_5 inst_cell_108_90 (.BL(BL90),.BLN(BLN90),.WL(WL108));
sram_cell_6t_5 inst_cell_108_91 (.BL(BL91),.BLN(BLN91),.WL(WL108));
sram_cell_6t_5 inst_cell_108_92 (.BL(BL92),.BLN(BLN92),.WL(WL108));
sram_cell_6t_5 inst_cell_108_93 (.BL(BL93),.BLN(BLN93),.WL(WL108));
sram_cell_6t_5 inst_cell_108_94 (.BL(BL94),.BLN(BLN94),.WL(WL108));
sram_cell_6t_5 inst_cell_108_95 (.BL(BL95),.BLN(BLN95),.WL(WL108));
sram_cell_6t_5 inst_cell_108_96 (.BL(BL96),.BLN(BLN96),.WL(WL108));
sram_cell_6t_5 inst_cell_108_97 (.BL(BL97),.BLN(BLN97),.WL(WL108));
sram_cell_6t_5 inst_cell_108_98 (.BL(BL98),.BLN(BLN98),.WL(WL108));
sram_cell_6t_5 inst_cell_108_99 (.BL(BL99),.BLN(BLN99),.WL(WL108));
sram_cell_6t_5 inst_cell_108_100 (.BL(BL100),.BLN(BLN100),.WL(WL108));
sram_cell_6t_5 inst_cell_108_101 (.BL(BL101),.BLN(BLN101),.WL(WL108));
sram_cell_6t_5 inst_cell_108_102 (.BL(BL102),.BLN(BLN102),.WL(WL108));
sram_cell_6t_5 inst_cell_108_103 (.BL(BL103),.BLN(BLN103),.WL(WL108));
sram_cell_6t_5 inst_cell_108_104 (.BL(BL104),.BLN(BLN104),.WL(WL108));
sram_cell_6t_5 inst_cell_108_105 (.BL(BL105),.BLN(BLN105),.WL(WL108));
sram_cell_6t_5 inst_cell_108_106 (.BL(BL106),.BLN(BLN106),.WL(WL108));
sram_cell_6t_5 inst_cell_108_107 (.BL(BL107),.BLN(BLN107),.WL(WL108));
sram_cell_6t_5 inst_cell_108_108 (.BL(BL108),.BLN(BLN108),.WL(WL108));
sram_cell_6t_5 inst_cell_108_109 (.BL(BL109),.BLN(BLN109),.WL(WL108));
sram_cell_6t_5 inst_cell_108_110 (.BL(BL110),.BLN(BLN110),.WL(WL108));
sram_cell_6t_5 inst_cell_108_111 (.BL(BL111),.BLN(BLN111),.WL(WL108));
sram_cell_6t_5 inst_cell_108_112 (.BL(BL112),.BLN(BLN112),.WL(WL108));
sram_cell_6t_5 inst_cell_108_113 (.BL(BL113),.BLN(BLN113),.WL(WL108));
sram_cell_6t_5 inst_cell_108_114 (.BL(BL114),.BLN(BLN114),.WL(WL108));
sram_cell_6t_5 inst_cell_108_115 (.BL(BL115),.BLN(BLN115),.WL(WL108));
sram_cell_6t_5 inst_cell_108_116 (.BL(BL116),.BLN(BLN116),.WL(WL108));
sram_cell_6t_5 inst_cell_108_117 (.BL(BL117),.BLN(BLN117),.WL(WL108));
sram_cell_6t_5 inst_cell_108_118 (.BL(BL118),.BLN(BLN118),.WL(WL108));
sram_cell_6t_5 inst_cell_108_119 (.BL(BL119),.BLN(BLN119),.WL(WL108));
sram_cell_6t_5 inst_cell_108_120 (.BL(BL120),.BLN(BLN120),.WL(WL108));
sram_cell_6t_5 inst_cell_108_121 (.BL(BL121),.BLN(BLN121),.WL(WL108));
sram_cell_6t_5 inst_cell_108_122 (.BL(BL122),.BLN(BLN122),.WL(WL108));
sram_cell_6t_5 inst_cell_108_123 (.BL(BL123),.BLN(BLN123),.WL(WL108));
sram_cell_6t_5 inst_cell_108_124 (.BL(BL124),.BLN(BLN124),.WL(WL108));
sram_cell_6t_5 inst_cell_108_125 (.BL(BL125),.BLN(BLN125),.WL(WL108));
sram_cell_6t_5 inst_cell_108_126 (.BL(BL126),.BLN(BLN126),.WL(WL108));
sram_cell_6t_5 inst_cell_108_127 (.BL(BL127),.BLN(BLN127),.WL(WL108));
sram_cell_6t_5 inst_cell_109_0 (.BL(BL0),.BLN(BLN0),.WL(WL109));
sram_cell_6t_5 inst_cell_109_1 (.BL(BL1),.BLN(BLN1),.WL(WL109));
sram_cell_6t_5 inst_cell_109_2 (.BL(BL2),.BLN(BLN2),.WL(WL109));
sram_cell_6t_5 inst_cell_109_3 (.BL(BL3),.BLN(BLN3),.WL(WL109));
sram_cell_6t_5 inst_cell_109_4 (.BL(BL4),.BLN(BLN4),.WL(WL109));
sram_cell_6t_5 inst_cell_109_5 (.BL(BL5),.BLN(BLN5),.WL(WL109));
sram_cell_6t_5 inst_cell_109_6 (.BL(BL6),.BLN(BLN6),.WL(WL109));
sram_cell_6t_5 inst_cell_109_7 (.BL(BL7),.BLN(BLN7),.WL(WL109));
sram_cell_6t_5 inst_cell_109_8 (.BL(BL8),.BLN(BLN8),.WL(WL109));
sram_cell_6t_5 inst_cell_109_9 (.BL(BL9),.BLN(BLN9),.WL(WL109));
sram_cell_6t_5 inst_cell_109_10 (.BL(BL10),.BLN(BLN10),.WL(WL109));
sram_cell_6t_5 inst_cell_109_11 (.BL(BL11),.BLN(BLN11),.WL(WL109));
sram_cell_6t_5 inst_cell_109_12 (.BL(BL12),.BLN(BLN12),.WL(WL109));
sram_cell_6t_5 inst_cell_109_13 (.BL(BL13),.BLN(BLN13),.WL(WL109));
sram_cell_6t_5 inst_cell_109_14 (.BL(BL14),.BLN(BLN14),.WL(WL109));
sram_cell_6t_5 inst_cell_109_15 (.BL(BL15),.BLN(BLN15),.WL(WL109));
sram_cell_6t_5 inst_cell_109_16 (.BL(BL16),.BLN(BLN16),.WL(WL109));
sram_cell_6t_5 inst_cell_109_17 (.BL(BL17),.BLN(BLN17),.WL(WL109));
sram_cell_6t_5 inst_cell_109_18 (.BL(BL18),.BLN(BLN18),.WL(WL109));
sram_cell_6t_5 inst_cell_109_19 (.BL(BL19),.BLN(BLN19),.WL(WL109));
sram_cell_6t_5 inst_cell_109_20 (.BL(BL20),.BLN(BLN20),.WL(WL109));
sram_cell_6t_5 inst_cell_109_21 (.BL(BL21),.BLN(BLN21),.WL(WL109));
sram_cell_6t_5 inst_cell_109_22 (.BL(BL22),.BLN(BLN22),.WL(WL109));
sram_cell_6t_5 inst_cell_109_23 (.BL(BL23),.BLN(BLN23),.WL(WL109));
sram_cell_6t_5 inst_cell_109_24 (.BL(BL24),.BLN(BLN24),.WL(WL109));
sram_cell_6t_5 inst_cell_109_25 (.BL(BL25),.BLN(BLN25),.WL(WL109));
sram_cell_6t_5 inst_cell_109_26 (.BL(BL26),.BLN(BLN26),.WL(WL109));
sram_cell_6t_5 inst_cell_109_27 (.BL(BL27),.BLN(BLN27),.WL(WL109));
sram_cell_6t_5 inst_cell_109_28 (.BL(BL28),.BLN(BLN28),.WL(WL109));
sram_cell_6t_5 inst_cell_109_29 (.BL(BL29),.BLN(BLN29),.WL(WL109));
sram_cell_6t_5 inst_cell_109_30 (.BL(BL30),.BLN(BLN30),.WL(WL109));
sram_cell_6t_5 inst_cell_109_31 (.BL(BL31),.BLN(BLN31),.WL(WL109));
sram_cell_6t_5 inst_cell_109_32 (.BL(BL32),.BLN(BLN32),.WL(WL109));
sram_cell_6t_5 inst_cell_109_33 (.BL(BL33),.BLN(BLN33),.WL(WL109));
sram_cell_6t_5 inst_cell_109_34 (.BL(BL34),.BLN(BLN34),.WL(WL109));
sram_cell_6t_5 inst_cell_109_35 (.BL(BL35),.BLN(BLN35),.WL(WL109));
sram_cell_6t_5 inst_cell_109_36 (.BL(BL36),.BLN(BLN36),.WL(WL109));
sram_cell_6t_5 inst_cell_109_37 (.BL(BL37),.BLN(BLN37),.WL(WL109));
sram_cell_6t_5 inst_cell_109_38 (.BL(BL38),.BLN(BLN38),.WL(WL109));
sram_cell_6t_5 inst_cell_109_39 (.BL(BL39),.BLN(BLN39),.WL(WL109));
sram_cell_6t_5 inst_cell_109_40 (.BL(BL40),.BLN(BLN40),.WL(WL109));
sram_cell_6t_5 inst_cell_109_41 (.BL(BL41),.BLN(BLN41),.WL(WL109));
sram_cell_6t_5 inst_cell_109_42 (.BL(BL42),.BLN(BLN42),.WL(WL109));
sram_cell_6t_5 inst_cell_109_43 (.BL(BL43),.BLN(BLN43),.WL(WL109));
sram_cell_6t_5 inst_cell_109_44 (.BL(BL44),.BLN(BLN44),.WL(WL109));
sram_cell_6t_5 inst_cell_109_45 (.BL(BL45),.BLN(BLN45),.WL(WL109));
sram_cell_6t_5 inst_cell_109_46 (.BL(BL46),.BLN(BLN46),.WL(WL109));
sram_cell_6t_5 inst_cell_109_47 (.BL(BL47),.BLN(BLN47),.WL(WL109));
sram_cell_6t_5 inst_cell_109_48 (.BL(BL48),.BLN(BLN48),.WL(WL109));
sram_cell_6t_5 inst_cell_109_49 (.BL(BL49),.BLN(BLN49),.WL(WL109));
sram_cell_6t_5 inst_cell_109_50 (.BL(BL50),.BLN(BLN50),.WL(WL109));
sram_cell_6t_5 inst_cell_109_51 (.BL(BL51),.BLN(BLN51),.WL(WL109));
sram_cell_6t_5 inst_cell_109_52 (.BL(BL52),.BLN(BLN52),.WL(WL109));
sram_cell_6t_5 inst_cell_109_53 (.BL(BL53),.BLN(BLN53),.WL(WL109));
sram_cell_6t_5 inst_cell_109_54 (.BL(BL54),.BLN(BLN54),.WL(WL109));
sram_cell_6t_5 inst_cell_109_55 (.BL(BL55),.BLN(BLN55),.WL(WL109));
sram_cell_6t_5 inst_cell_109_56 (.BL(BL56),.BLN(BLN56),.WL(WL109));
sram_cell_6t_5 inst_cell_109_57 (.BL(BL57),.BLN(BLN57),.WL(WL109));
sram_cell_6t_5 inst_cell_109_58 (.BL(BL58),.BLN(BLN58),.WL(WL109));
sram_cell_6t_5 inst_cell_109_59 (.BL(BL59),.BLN(BLN59),.WL(WL109));
sram_cell_6t_5 inst_cell_109_60 (.BL(BL60),.BLN(BLN60),.WL(WL109));
sram_cell_6t_5 inst_cell_109_61 (.BL(BL61),.BLN(BLN61),.WL(WL109));
sram_cell_6t_5 inst_cell_109_62 (.BL(BL62),.BLN(BLN62),.WL(WL109));
sram_cell_6t_5 inst_cell_109_63 (.BL(BL63),.BLN(BLN63),.WL(WL109));
sram_cell_6t_5 inst_cell_109_64 (.BL(BL64),.BLN(BLN64),.WL(WL109));
sram_cell_6t_5 inst_cell_109_65 (.BL(BL65),.BLN(BLN65),.WL(WL109));
sram_cell_6t_5 inst_cell_109_66 (.BL(BL66),.BLN(BLN66),.WL(WL109));
sram_cell_6t_5 inst_cell_109_67 (.BL(BL67),.BLN(BLN67),.WL(WL109));
sram_cell_6t_5 inst_cell_109_68 (.BL(BL68),.BLN(BLN68),.WL(WL109));
sram_cell_6t_5 inst_cell_109_69 (.BL(BL69),.BLN(BLN69),.WL(WL109));
sram_cell_6t_5 inst_cell_109_70 (.BL(BL70),.BLN(BLN70),.WL(WL109));
sram_cell_6t_5 inst_cell_109_71 (.BL(BL71),.BLN(BLN71),.WL(WL109));
sram_cell_6t_5 inst_cell_109_72 (.BL(BL72),.BLN(BLN72),.WL(WL109));
sram_cell_6t_5 inst_cell_109_73 (.BL(BL73),.BLN(BLN73),.WL(WL109));
sram_cell_6t_5 inst_cell_109_74 (.BL(BL74),.BLN(BLN74),.WL(WL109));
sram_cell_6t_5 inst_cell_109_75 (.BL(BL75),.BLN(BLN75),.WL(WL109));
sram_cell_6t_5 inst_cell_109_76 (.BL(BL76),.BLN(BLN76),.WL(WL109));
sram_cell_6t_5 inst_cell_109_77 (.BL(BL77),.BLN(BLN77),.WL(WL109));
sram_cell_6t_5 inst_cell_109_78 (.BL(BL78),.BLN(BLN78),.WL(WL109));
sram_cell_6t_5 inst_cell_109_79 (.BL(BL79),.BLN(BLN79),.WL(WL109));
sram_cell_6t_5 inst_cell_109_80 (.BL(BL80),.BLN(BLN80),.WL(WL109));
sram_cell_6t_5 inst_cell_109_81 (.BL(BL81),.BLN(BLN81),.WL(WL109));
sram_cell_6t_5 inst_cell_109_82 (.BL(BL82),.BLN(BLN82),.WL(WL109));
sram_cell_6t_5 inst_cell_109_83 (.BL(BL83),.BLN(BLN83),.WL(WL109));
sram_cell_6t_5 inst_cell_109_84 (.BL(BL84),.BLN(BLN84),.WL(WL109));
sram_cell_6t_5 inst_cell_109_85 (.BL(BL85),.BLN(BLN85),.WL(WL109));
sram_cell_6t_5 inst_cell_109_86 (.BL(BL86),.BLN(BLN86),.WL(WL109));
sram_cell_6t_5 inst_cell_109_87 (.BL(BL87),.BLN(BLN87),.WL(WL109));
sram_cell_6t_5 inst_cell_109_88 (.BL(BL88),.BLN(BLN88),.WL(WL109));
sram_cell_6t_5 inst_cell_109_89 (.BL(BL89),.BLN(BLN89),.WL(WL109));
sram_cell_6t_5 inst_cell_109_90 (.BL(BL90),.BLN(BLN90),.WL(WL109));
sram_cell_6t_5 inst_cell_109_91 (.BL(BL91),.BLN(BLN91),.WL(WL109));
sram_cell_6t_5 inst_cell_109_92 (.BL(BL92),.BLN(BLN92),.WL(WL109));
sram_cell_6t_5 inst_cell_109_93 (.BL(BL93),.BLN(BLN93),.WL(WL109));
sram_cell_6t_5 inst_cell_109_94 (.BL(BL94),.BLN(BLN94),.WL(WL109));
sram_cell_6t_5 inst_cell_109_95 (.BL(BL95),.BLN(BLN95),.WL(WL109));
sram_cell_6t_5 inst_cell_109_96 (.BL(BL96),.BLN(BLN96),.WL(WL109));
sram_cell_6t_5 inst_cell_109_97 (.BL(BL97),.BLN(BLN97),.WL(WL109));
sram_cell_6t_5 inst_cell_109_98 (.BL(BL98),.BLN(BLN98),.WL(WL109));
sram_cell_6t_5 inst_cell_109_99 (.BL(BL99),.BLN(BLN99),.WL(WL109));
sram_cell_6t_5 inst_cell_109_100 (.BL(BL100),.BLN(BLN100),.WL(WL109));
sram_cell_6t_5 inst_cell_109_101 (.BL(BL101),.BLN(BLN101),.WL(WL109));
sram_cell_6t_5 inst_cell_109_102 (.BL(BL102),.BLN(BLN102),.WL(WL109));
sram_cell_6t_5 inst_cell_109_103 (.BL(BL103),.BLN(BLN103),.WL(WL109));
sram_cell_6t_5 inst_cell_109_104 (.BL(BL104),.BLN(BLN104),.WL(WL109));
sram_cell_6t_5 inst_cell_109_105 (.BL(BL105),.BLN(BLN105),.WL(WL109));
sram_cell_6t_5 inst_cell_109_106 (.BL(BL106),.BLN(BLN106),.WL(WL109));
sram_cell_6t_5 inst_cell_109_107 (.BL(BL107),.BLN(BLN107),.WL(WL109));
sram_cell_6t_5 inst_cell_109_108 (.BL(BL108),.BLN(BLN108),.WL(WL109));
sram_cell_6t_5 inst_cell_109_109 (.BL(BL109),.BLN(BLN109),.WL(WL109));
sram_cell_6t_5 inst_cell_109_110 (.BL(BL110),.BLN(BLN110),.WL(WL109));
sram_cell_6t_5 inst_cell_109_111 (.BL(BL111),.BLN(BLN111),.WL(WL109));
sram_cell_6t_5 inst_cell_109_112 (.BL(BL112),.BLN(BLN112),.WL(WL109));
sram_cell_6t_5 inst_cell_109_113 (.BL(BL113),.BLN(BLN113),.WL(WL109));
sram_cell_6t_5 inst_cell_109_114 (.BL(BL114),.BLN(BLN114),.WL(WL109));
sram_cell_6t_5 inst_cell_109_115 (.BL(BL115),.BLN(BLN115),.WL(WL109));
sram_cell_6t_5 inst_cell_109_116 (.BL(BL116),.BLN(BLN116),.WL(WL109));
sram_cell_6t_5 inst_cell_109_117 (.BL(BL117),.BLN(BLN117),.WL(WL109));
sram_cell_6t_5 inst_cell_109_118 (.BL(BL118),.BLN(BLN118),.WL(WL109));
sram_cell_6t_5 inst_cell_109_119 (.BL(BL119),.BLN(BLN119),.WL(WL109));
sram_cell_6t_5 inst_cell_109_120 (.BL(BL120),.BLN(BLN120),.WL(WL109));
sram_cell_6t_5 inst_cell_109_121 (.BL(BL121),.BLN(BLN121),.WL(WL109));
sram_cell_6t_5 inst_cell_109_122 (.BL(BL122),.BLN(BLN122),.WL(WL109));
sram_cell_6t_5 inst_cell_109_123 (.BL(BL123),.BLN(BLN123),.WL(WL109));
sram_cell_6t_5 inst_cell_109_124 (.BL(BL124),.BLN(BLN124),.WL(WL109));
sram_cell_6t_5 inst_cell_109_125 (.BL(BL125),.BLN(BLN125),.WL(WL109));
sram_cell_6t_5 inst_cell_109_126 (.BL(BL126),.BLN(BLN126),.WL(WL109));
sram_cell_6t_5 inst_cell_109_127 (.BL(BL127),.BLN(BLN127),.WL(WL109));
sram_cell_6t_5 inst_cell_110_0 (.BL(BL0),.BLN(BLN0),.WL(WL110));
sram_cell_6t_5 inst_cell_110_1 (.BL(BL1),.BLN(BLN1),.WL(WL110));
sram_cell_6t_5 inst_cell_110_2 (.BL(BL2),.BLN(BLN2),.WL(WL110));
sram_cell_6t_5 inst_cell_110_3 (.BL(BL3),.BLN(BLN3),.WL(WL110));
sram_cell_6t_5 inst_cell_110_4 (.BL(BL4),.BLN(BLN4),.WL(WL110));
sram_cell_6t_5 inst_cell_110_5 (.BL(BL5),.BLN(BLN5),.WL(WL110));
sram_cell_6t_5 inst_cell_110_6 (.BL(BL6),.BLN(BLN6),.WL(WL110));
sram_cell_6t_5 inst_cell_110_7 (.BL(BL7),.BLN(BLN7),.WL(WL110));
sram_cell_6t_5 inst_cell_110_8 (.BL(BL8),.BLN(BLN8),.WL(WL110));
sram_cell_6t_5 inst_cell_110_9 (.BL(BL9),.BLN(BLN9),.WL(WL110));
sram_cell_6t_5 inst_cell_110_10 (.BL(BL10),.BLN(BLN10),.WL(WL110));
sram_cell_6t_5 inst_cell_110_11 (.BL(BL11),.BLN(BLN11),.WL(WL110));
sram_cell_6t_5 inst_cell_110_12 (.BL(BL12),.BLN(BLN12),.WL(WL110));
sram_cell_6t_5 inst_cell_110_13 (.BL(BL13),.BLN(BLN13),.WL(WL110));
sram_cell_6t_5 inst_cell_110_14 (.BL(BL14),.BLN(BLN14),.WL(WL110));
sram_cell_6t_5 inst_cell_110_15 (.BL(BL15),.BLN(BLN15),.WL(WL110));
sram_cell_6t_5 inst_cell_110_16 (.BL(BL16),.BLN(BLN16),.WL(WL110));
sram_cell_6t_5 inst_cell_110_17 (.BL(BL17),.BLN(BLN17),.WL(WL110));
sram_cell_6t_5 inst_cell_110_18 (.BL(BL18),.BLN(BLN18),.WL(WL110));
sram_cell_6t_5 inst_cell_110_19 (.BL(BL19),.BLN(BLN19),.WL(WL110));
sram_cell_6t_5 inst_cell_110_20 (.BL(BL20),.BLN(BLN20),.WL(WL110));
sram_cell_6t_5 inst_cell_110_21 (.BL(BL21),.BLN(BLN21),.WL(WL110));
sram_cell_6t_5 inst_cell_110_22 (.BL(BL22),.BLN(BLN22),.WL(WL110));
sram_cell_6t_5 inst_cell_110_23 (.BL(BL23),.BLN(BLN23),.WL(WL110));
sram_cell_6t_5 inst_cell_110_24 (.BL(BL24),.BLN(BLN24),.WL(WL110));
sram_cell_6t_5 inst_cell_110_25 (.BL(BL25),.BLN(BLN25),.WL(WL110));
sram_cell_6t_5 inst_cell_110_26 (.BL(BL26),.BLN(BLN26),.WL(WL110));
sram_cell_6t_5 inst_cell_110_27 (.BL(BL27),.BLN(BLN27),.WL(WL110));
sram_cell_6t_5 inst_cell_110_28 (.BL(BL28),.BLN(BLN28),.WL(WL110));
sram_cell_6t_5 inst_cell_110_29 (.BL(BL29),.BLN(BLN29),.WL(WL110));
sram_cell_6t_5 inst_cell_110_30 (.BL(BL30),.BLN(BLN30),.WL(WL110));
sram_cell_6t_5 inst_cell_110_31 (.BL(BL31),.BLN(BLN31),.WL(WL110));
sram_cell_6t_5 inst_cell_110_32 (.BL(BL32),.BLN(BLN32),.WL(WL110));
sram_cell_6t_5 inst_cell_110_33 (.BL(BL33),.BLN(BLN33),.WL(WL110));
sram_cell_6t_5 inst_cell_110_34 (.BL(BL34),.BLN(BLN34),.WL(WL110));
sram_cell_6t_5 inst_cell_110_35 (.BL(BL35),.BLN(BLN35),.WL(WL110));
sram_cell_6t_5 inst_cell_110_36 (.BL(BL36),.BLN(BLN36),.WL(WL110));
sram_cell_6t_5 inst_cell_110_37 (.BL(BL37),.BLN(BLN37),.WL(WL110));
sram_cell_6t_5 inst_cell_110_38 (.BL(BL38),.BLN(BLN38),.WL(WL110));
sram_cell_6t_5 inst_cell_110_39 (.BL(BL39),.BLN(BLN39),.WL(WL110));
sram_cell_6t_5 inst_cell_110_40 (.BL(BL40),.BLN(BLN40),.WL(WL110));
sram_cell_6t_5 inst_cell_110_41 (.BL(BL41),.BLN(BLN41),.WL(WL110));
sram_cell_6t_5 inst_cell_110_42 (.BL(BL42),.BLN(BLN42),.WL(WL110));
sram_cell_6t_5 inst_cell_110_43 (.BL(BL43),.BLN(BLN43),.WL(WL110));
sram_cell_6t_5 inst_cell_110_44 (.BL(BL44),.BLN(BLN44),.WL(WL110));
sram_cell_6t_5 inst_cell_110_45 (.BL(BL45),.BLN(BLN45),.WL(WL110));
sram_cell_6t_5 inst_cell_110_46 (.BL(BL46),.BLN(BLN46),.WL(WL110));
sram_cell_6t_5 inst_cell_110_47 (.BL(BL47),.BLN(BLN47),.WL(WL110));
sram_cell_6t_5 inst_cell_110_48 (.BL(BL48),.BLN(BLN48),.WL(WL110));
sram_cell_6t_5 inst_cell_110_49 (.BL(BL49),.BLN(BLN49),.WL(WL110));
sram_cell_6t_5 inst_cell_110_50 (.BL(BL50),.BLN(BLN50),.WL(WL110));
sram_cell_6t_5 inst_cell_110_51 (.BL(BL51),.BLN(BLN51),.WL(WL110));
sram_cell_6t_5 inst_cell_110_52 (.BL(BL52),.BLN(BLN52),.WL(WL110));
sram_cell_6t_5 inst_cell_110_53 (.BL(BL53),.BLN(BLN53),.WL(WL110));
sram_cell_6t_5 inst_cell_110_54 (.BL(BL54),.BLN(BLN54),.WL(WL110));
sram_cell_6t_5 inst_cell_110_55 (.BL(BL55),.BLN(BLN55),.WL(WL110));
sram_cell_6t_5 inst_cell_110_56 (.BL(BL56),.BLN(BLN56),.WL(WL110));
sram_cell_6t_5 inst_cell_110_57 (.BL(BL57),.BLN(BLN57),.WL(WL110));
sram_cell_6t_5 inst_cell_110_58 (.BL(BL58),.BLN(BLN58),.WL(WL110));
sram_cell_6t_5 inst_cell_110_59 (.BL(BL59),.BLN(BLN59),.WL(WL110));
sram_cell_6t_5 inst_cell_110_60 (.BL(BL60),.BLN(BLN60),.WL(WL110));
sram_cell_6t_5 inst_cell_110_61 (.BL(BL61),.BLN(BLN61),.WL(WL110));
sram_cell_6t_5 inst_cell_110_62 (.BL(BL62),.BLN(BLN62),.WL(WL110));
sram_cell_6t_5 inst_cell_110_63 (.BL(BL63),.BLN(BLN63),.WL(WL110));
sram_cell_6t_5 inst_cell_110_64 (.BL(BL64),.BLN(BLN64),.WL(WL110));
sram_cell_6t_5 inst_cell_110_65 (.BL(BL65),.BLN(BLN65),.WL(WL110));
sram_cell_6t_5 inst_cell_110_66 (.BL(BL66),.BLN(BLN66),.WL(WL110));
sram_cell_6t_5 inst_cell_110_67 (.BL(BL67),.BLN(BLN67),.WL(WL110));
sram_cell_6t_5 inst_cell_110_68 (.BL(BL68),.BLN(BLN68),.WL(WL110));
sram_cell_6t_5 inst_cell_110_69 (.BL(BL69),.BLN(BLN69),.WL(WL110));
sram_cell_6t_5 inst_cell_110_70 (.BL(BL70),.BLN(BLN70),.WL(WL110));
sram_cell_6t_5 inst_cell_110_71 (.BL(BL71),.BLN(BLN71),.WL(WL110));
sram_cell_6t_5 inst_cell_110_72 (.BL(BL72),.BLN(BLN72),.WL(WL110));
sram_cell_6t_5 inst_cell_110_73 (.BL(BL73),.BLN(BLN73),.WL(WL110));
sram_cell_6t_5 inst_cell_110_74 (.BL(BL74),.BLN(BLN74),.WL(WL110));
sram_cell_6t_5 inst_cell_110_75 (.BL(BL75),.BLN(BLN75),.WL(WL110));
sram_cell_6t_5 inst_cell_110_76 (.BL(BL76),.BLN(BLN76),.WL(WL110));
sram_cell_6t_5 inst_cell_110_77 (.BL(BL77),.BLN(BLN77),.WL(WL110));
sram_cell_6t_5 inst_cell_110_78 (.BL(BL78),.BLN(BLN78),.WL(WL110));
sram_cell_6t_5 inst_cell_110_79 (.BL(BL79),.BLN(BLN79),.WL(WL110));
sram_cell_6t_5 inst_cell_110_80 (.BL(BL80),.BLN(BLN80),.WL(WL110));
sram_cell_6t_5 inst_cell_110_81 (.BL(BL81),.BLN(BLN81),.WL(WL110));
sram_cell_6t_5 inst_cell_110_82 (.BL(BL82),.BLN(BLN82),.WL(WL110));
sram_cell_6t_5 inst_cell_110_83 (.BL(BL83),.BLN(BLN83),.WL(WL110));
sram_cell_6t_5 inst_cell_110_84 (.BL(BL84),.BLN(BLN84),.WL(WL110));
sram_cell_6t_5 inst_cell_110_85 (.BL(BL85),.BLN(BLN85),.WL(WL110));
sram_cell_6t_5 inst_cell_110_86 (.BL(BL86),.BLN(BLN86),.WL(WL110));
sram_cell_6t_5 inst_cell_110_87 (.BL(BL87),.BLN(BLN87),.WL(WL110));
sram_cell_6t_5 inst_cell_110_88 (.BL(BL88),.BLN(BLN88),.WL(WL110));
sram_cell_6t_5 inst_cell_110_89 (.BL(BL89),.BLN(BLN89),.WL(WL110));
sram_cell_6t_5 inst_cell_110_90 (.BL(BL90),.BLN(BLN90),.WL(WL110));
sram_cell_6t_5 inst_cell_110_91 (.BL(BL91),.BLN(BLN91),.WL(WL110));
sram_cell_6t_5 inst_cell_110_92 (.BL(BL92),.BLN(BLN92),.WL(WL110));
sram_cell_6t_5 inst_cell_110_93 (.BL(BL93),.BLN(BLN93),.WL(WL110));
sram_cell_6t_5 inst_cell_110_94 (.BL(BL94),.BLN(BLN94),.WL(WL110));
sram_cell_6t_5 inst_cell_110_95 (.BL(BL95),.BLN(BLN95),.WL(WL110));
sram_cell_6t_5 inst_cell_110_96 (.BL(BL96),.BLN(BLN96),.WL(WL110));
sram_cell_6t_5 inst_cell_110_97 (.BL(BL97),.BLN(BLN97),.WL(WL110));
sram_cell_6t_5 inst_cell_110_98 (.BL(BL98),.BLN(BLN98),.WL(WL110));
sram_cell_6t_5 inst_cell_110_99 (.BL(BL99),.BLN(BLN99),.WL(WL110));
sram_cell_6t_5 inst_cell_110_100 (.BL(BL100),.BLN(BLN100),.WL(WL110));
sram_cell_6t_5 inst_cell_110_101 (.BL(BL101),.BLN(BLN101),.WL(WL110));
sram_cell_6t_5 inst_cell_110_102 (.BL(BL102),.BLN(BLN102),.WL(WL110));
sram_cell_6t_5 inst_cell_110_103 (.BL(BL103),.BLN(BLN103),.WL(WL110));
sram_cell_6t_5 inst_cell_110_104 (.BL(BL104),.BLN(BLN104),.WL(WL110));
sram_cell_6t_5 inst_cell_110_105 (.BL(BL105),.BLN(BLN105),.WL(WL110));
sram_cell_6t_5 inst_cell_110_106 (.BL(BL106),.BLN(BLN106),.WL(WL110));
sram_cell_6t_5 inst_cell_110_107 (.BL(BL107),.BLN(BLN107),.WL(WL110));
sram_cell_6t_5 inst_cell_110_108 (.BL(BL108),.BLN(BLN108),.WL(WL110));
sram_cell_6t_5 inst_cell_110_109 (.BL(BL109),.BLN(BLN109),.WL(WL110));
sram_cell_6t_5 inst_cell_110_110 (.BL(BL110),.BLN(BLN110),.WL(WL110));
sram_cell_6t_5 inst_cell_110_111 (.BL(BL111),.BLN(BLN111),.WL(WL110));
sram_cell_6t_5 inst_cell_110_112 (.BL(BL112),.BLN(BLN112),.WL(WL110));
sram_cell_6t_5 inst_cell_110_113 (.BL(BL113),.BLN(BLN113),.WL(WL110));
sram_cell_6t_5 inst_cell_110_114 (.BL(BL114),.BLN(BLN114),.WL(WL110));
sram_cell_6t_5 inst_cell_110_115 (.BL(BL115),.BLN(BLN115),.WL(WL110));
sram_cell_6t_5 inst_cell_110_116 (.BL(BL116),.BLN(BLN116),.WL(WL110));
sram_cell_6t_5 inst_cell_110_117 (.BL(BL117),.BLN(BLN117),.WL(WL110));
sram_cell_6t_5 inst_cell_110_118 (.BL(BL118),.BLN(BLN118),.WL(WL110));
sram_cell_6t_5 inst_cell_110_119 (.BL(BL119),.BLN(BLN119),.WL(WL110));
sram_cell_6t_5 inst_cell_110_120 (.BL(BL120),.BLN(BLN120),.WL(WL110));
sram_cell_6t_5 inst_cell_110_121 (.BL(BL121),.BLN(BLN121),.WL(WL110));
sram_cell_6t_5 inst_cell_110_122 (.BL(BL122),.BLN(BLN122),.WL(WL110));
sram_cell_6t_5 inst_cell_110_123 (.BL(BL123),.BLN(BLN123),.WL(WL110));
sram_cell_6t_5 inst_cell_110_124 (.BL(BL124),.BLN(BLN124),.WL(WL110));
sram_cell_6t_5 inst_cell_110_125 (.BL(BL125),.BLN(BLN125),.WL(WL110));
sram_cell_6t_5 inst_cell_110_126 (.BL(BL126),.BLN(BLN126),.WL(WL110));
sram_cell_6t_5 inst_cell_110_127 (.BL(BL127),.BLN(BLN127),.WL(WL110));
sram_cell_6t_5 inst_cell_111_0 (.BL(BL0),.BLN(BLN0),.WL(WL111));
sram_cell_6t_5 inst_cell_111_1 (.BL(BL1),.BLN(BLN1),.WL(WL111));
sram_cell_6t_5 inst_cell_111_2 (.BL(BL2),.BLN(BLN2),.WL(WL111));
sram_cell_6t_5 inst_cell_111_3 (.BL(BL3),.BLN(BLN3),.WL(WL111));
sram_cell_6t_5 inst_cell_111_4 (.BL(BL4),.BLN(BLN4),.WL(WL111));
sram_cell_6t_5 inst_cell_111_5 (.BL(BL5),.BLN(BLN5),.WL(WL111));
sram_cell_6t_5 inst_cell_111_6 (.BL(BL6),.BLN(BLN6),.WL(WL111));
sram_cell_6t_5 inst_cell_111_7 (.BL(BL7),.BLN(BLN7),.WL(WL111));
sram_cell_6t_5 inst_cell_111_8 (.BL(BL8),.BLN(BLN8),.WL(WL111));
sram_cell_6t_5 inst_cell_111_9 (.BL(BL9),.BLN(BLN9),.WL(WL111));
sram_cell_6t_5 inst_cell_111_10 (.BL(BL10),.BLN(BLN10),.WL(WL111));
sram_cell_6t_5 inst_cell_111_11 (.BL(BL11),.BLN(BLN11),.WL(WL111));
sram_cell_6t_5 inst_cell_111_12 (.BL(BL12),.BLN(BLN12),.WL(WL111));
sram_cell_6t_5 inst_cell_111_13 (.BL(BL13),.BLN(BLN13),.WL(WL111));
sram_cell_6t_5 inst_cell_111_14 (.BL(BL14),.BLN(BLN14),.WL(WL111));
sram_cell_6t_5 inst_cell_111_15 (.BL(BL15),.BLN(BLN15),.WL(WL111));
sram_cell_6t_5 inst_cell_111_16 (.BL(BL16),.BLN(BLN16),.WL(WL111));
sram_cell_6t_5 inst_cell_111_17 (.BL(BL17),.BLN(BLN17),.WL(WL111));
sram_cell_6t_5 inst_cell_111_18 (.BL(BL18),.BLN(BLN18),.WL(WL111));
sram_cell_6t_5 inst_cell_111_19 (.BL(BL19),.BLN(BLN19),.WL(WL111));
sram_cell_6t_5 inst_cell_111_20 (.BL(BL20),.BLN(BLN20),.WL(WL111));
sram_cell_6t_5 inst_cell_111_21 (.BL(BL21),.BLN(BLN21),.WL(WL111));
sram_cell_6t_5 inst_cell_111_22 (.BL(BL22),.BLN(BLN22),.WL(WL111));
sram_cell_6t_5 inst_cell_111_23 (.BL(BL23),.BLN(BLN23),.WL(WL111));
sram_cell_6t_5 inst_cell_111_24 (.BL(BL24),.BLN(BLN24),.WL(WL111));
sram_cell_6t_5 inst_cell_111_25 (.BL(BL25),.BLN(BLN25),.WL(WL111));
sram_cell_6t_5 inst_cell_111_26 (.BL(BL26),.BLN(BLN26),.WL(WL111));
sram_cell_6t_5 inst_cell_111_27 (.BL(BL27),.BLN(BLN27),.WL(WL111));
sram_cell_6t_5 inst_cell_111_28 (.BL(BL28),.BLN(BLN28),.WL(WL111));
sram_cell_6t_5 inst_cell_111_29 (.BL(BL29),.BLN(BLN29),.WL(WL111));
sram_cell_6t_5 inst_cell_111_30 (.BL(BL30),.BLN(BLN30),.WL(WL111));
sram_cell_6t_5 inst_cell_111_31 (.BL(BL31),.BLN(BLN31),.WL(WL111));
sram_cell_6t_5 inst_cell_111_32 (.BL(BL32),.BLN(BLN32),.WL(WL111));
sram_cell_6t_5 inst_cell_111_33 (.BL(BL33),.BLN(BLN33),.WL(WL111));
sram_cell_6t_5 inst_cell_111_34 (.BL(BL34),.BLN(BLN34),.WL(WL111));
sram_cell_6t_5 inst_cell_111_35 (.BL(BL35),.BLN(BLN35),.WL(WL111));
sram_cell_6t_5 inst_cell_111_36 (.BL(BL36),.BLN(BLN36),.WL(WL111));
sram_cell_6t_5 inst_cell_111_37 (.BL(BL37),.BLN(BLN37),.WL(WL111));
sram_cell_6t_5 inst_cell_111_38 (.BL(BL38),.BLN(BLN38),.WL(WL111));
sram_cell_6t_5 inst_cell_111_39 (.BL(BL39),.BLN(BLN39),.WL(WL111));
sram_cell_6t_5 inst_cell_111_40 (.BL(BL40),.BLN(BLN40),.WL(WL111));
sram_cell_6t_5 inst_cell_111_41 (.BL(BL41),.BLN(BLN41),.WL(WL111));
sram_cell_6t_5 inst_cell_111_42 (.BL(BL42),.BLN(BLN42),.WL(WL111));
sram_cell_6t_5 inst_cell_111_43 (.BL(BL43),.BLN(BLN43),.WL(WL111));
sram_cell_6t_5 inst_cell_111_44 (.BL(BL44),.BLN(BLN44),.WL(WL111));
sram_cell_6t_5 inst_cell_111_45 (.BL(BL45),.BLN(BLN45),.WL(WL111));
sram_cell_6t_5 inst_cell_111_46 (.BL(BL46),.BLN(BLN46),.WL(WL111));
sram_cell_6t_5 inst_cell_111_47 (.BL(BL47),.BLN(BLN47),.WL(WL111));
sram_cell_6t_5 inst_cell_111_48 (.BL(BL48),.BLN(BLN48),.WL(WL111));
sram_cell_6t_5 inst_cell_111_49 (.BL(BL49),.BLN(BLN49),.WL(WL111));
sram_cell_6t_5 inst_cell_111_50 (.BL(BL50),.BLN(BLN50),.WL(WL111));
sram_cell_6t_5 inst_cell_111_51 (.BL(BL51),.BLN(BLN51),.WL(WL111));
sram_cell_6t_5 inst_cell_111_52 (.BL(BL52),.BLN(BLN52),.WL(WL111));
sram_cell_6t_5 inst_cell_111_53 (.BL(BL53),.BLN(BLN53),.WL(WL111));
sram_cell_6t_5 inst_cell_111_54 (.BL(BL54),.BLN(BLN54),.WL(WL111));
sram_cell_6t_5 inst_cell_111_55 (.BL(BL55),.BLN(BLN55),.WL(WL111));
sram_cell_6t_5 inst_cell_111_56 (.BL(BL56),.BLN(BLN56),.WL(WL111));
sram_cell_6t_5 inst_cell_111_57 (.BL(BL57),.BLN(BLN57),.WL(WL111));
sram_cell_6t_5 inst_cell_111_58 (.BL(BL58),.BLN(BLN58),.WL(WL111));
sram_cell_6t_5 inst_cell_111_59 (.BL(BL59),.BLN(BLN59),.WL(WL111));
sram_cell_6t_5 inst_cell_111_60 (.BL(BL60),.BLN(BLN60),.WL(WL111));
sram_cell_6t_5 inst_cell_111_61 (.BL(BL61),.BLN(BLN61),.WL(WL111));
sram_cell_6t_5 inst_cell_111_62 (.BL(BL62),.BLN(BLN62),.WL(WL111));
sram_cell_6t_5 inst_cell_111_63 (.BL(BL63),.BLN(BLN63),.WL(WL111));
sram_cell_6t_5 inst_cell_111_64 (.BL(BL64),.BLN(BLN64),.WL(WL111));
sram_cell_6t_5 inst_cell_111_65 (.BL(BL65),.BLN(BLN65),.WL(WL111));
sram_cell_6t_5 inst_cell_111_66 (.BL(BL66),.BLN(BLN66),.WL(WL111));
sram_cell_6t_5 inst_cell_111_67 (.BL(BL67),.BLN(BLN67),.WL(WL111));
sram_cell_6t_5 inst_cell_111_68 (.BL(BL68),.BLN(BLN68),.WL(WL111));
sram_cell_6t_5 inst_cell_111_69 (.BL(BL69),.BLN(BLN69),.WL(WL111));
sram_cell_6t_5 inst_cell_111_70 (.BL(BL70),.BLN(BLN70),.WL(WL111));
sram_cell_6t_5 inst_cell_111_71 (.BL(BL71),.BLN(BLN71),.WL(WL111));
sram_cell_6t_5 inst_cell_111_72 (.BL(BL72),.BLN(BLN72),.WL(WL111));
sram_cell_6t_5 inst_cell_111_73 (.BL(BL73),.BLN(BLN73),.WL(WL111));
sram_cell_6t_5 inst_cell_111_74 (.BL(BL74),.BLN(BLN74),.WL(WL111));
sram_cell_6t_5 inst_cell_111_75 (.BL(BL75),.BLN(BLN75),.WL(WL111));
sram_cell_6t_5 inst_cell_111_76 (.BL(BL76),.BLN(BLN76),.WL(WL111));
sram_cell_6t_5 inst_cell_111_77 (.BL(BL77),.BLN(BLN77),.WL(WL111));
sram_cell_6t_5 inst_cell_111_78 (.BL(BL78),.BLN(BLN78),.WL(WL111));
sram_cell_6t_5 inst_cell_111_79 (.BL(BL79),.BLN(BLN79),.WL(WL111));
sram_cell_6t_5 inst_cell_111_80 (.BL(BL80),.BLN(BLN80),.WL(WL111));
sram_cell_6t_5 inst_cell_111_81 (.BL(BL81),.BLN(BLN81),.WL(WL111));
sram_cell_6t_5 inst_cell_111_82 (.BL(BL82),.BLN(BLN82),.WL(WL111));
sram_cell_6t_5 inst_cell_111_83 (.BL(BL83),.BLN(BLN83),.WL(WL111));
sram_cell_6t_5 inst_cell_111_84 (.BL(BL84),.BLN(BLN84),.WL(WL111));
sram_cell_6t_5 inst_cell_111_85 (.BL(BL85),.BLN(BLN85),.WL(WL111));
sram_cell_6t_5 inst_cell_111_86 (.BL(BL86),.BLN(BLN86),.WL(WL111));
sram_cell_6t_5 inst_cell_111_87 (.BL(BL87),.BLN(BLN87),.WL(WL111));
sram_cell_6t_5 inst_cell_111_88 (.BL(BL88),.BLN(BLN88),.WL(WL111));
sram_cell_6t_5 inst_cell_111_89 (.BL(BL89),.BLN(BLN89),.WL(WL111));
sram_cell_6t_5 inst_cell_111_90 (.BL(BL90),.BLN(BLN90),.WL(WL111));
sram_cell_6t_5 inst_cell_111_91 (.BL(BL91),.BLN(BLN91),.WL(WL111));
sram_cell_6t_5 inst_cell_111_92 (.BL(BL92),.BLN(BLN92),.WL(WL111));
sram_cell_6t_5 inst_cell_111_93 (.BL(BL93),.BLN(BLN93),.WL(WL111));
sram_cell_6t_5 inst_cell_111_94 (.BL(BL94),.BLN(BLN94),.WL(WL111));
sram_cell_6t_5 inst_cell_111_95 (.BL(BL95),.BLN(BLN95),.WL(WL111));
sram_cell_6t_5 inst_cell_111_96 (.BL(BL96),.BLN(BLN96),.WL(WL111));
sram_cell_6t_5 inst_cell_111_97 (.BL(BL97),.BLN(BLN97),.WL(WL111));
sram_cell_6t_5 inst_cell_111_98 (.BL(BL98),.BLN(BLN98),.WL(WL111));
sram_cell_6t_5 inst_cell_111_99 (.BL(BL99),.BLN(BLN99),.WL(WL111));
sram_cell_6t_5 inst_cell_111_100 (.BL(BL100),.BLN(BLN100),.WL(WL111));
sram_cell_6t_5 inst_cell_111_101 (.BL(BL101),.BLN(BLN101),.WL(WL111));
sram_cell_6t_5 inst_cell_111_102 (.BL(BL102),.BLN(BLN102),.WL(WL111));
sram_cell_6t_5 inst_cell_111_103 (.BL(BL103),.BLN(BLN103),.WL(WL111));
sram_cell_6t_5 inst_cell_111_104 (.BL(BL104),.BLN(BLN104),.WL(WL111));
sram_cell_6t_5 inst_cell_111_105 (.BL(BL105),.BLN(BLN105),.WL(WL111));
sram_cell_6t_5 inst_cell_111_106 (.BL(BL106),.BLN(BLN106),.WL(WL111));
sram_cell_6t_5 inst_cell_111_107 (.BL(BL107),.BLN(BLN107),.WL(WL111));
sram_cell_6t_5 inst_cell_111_108 (.BL(BL108),.BLN(BLN108),.WL(WL111));
sram_cell_6t_5 inst_cell_111_109 (.BL(BL109),.BLN(BLN109),.WL(WL111));
sram_cell_6t_5 inst_cell_111_110 (.BL(BL110),.BLN(BLN110),.WL(WL111));
sram_cell_6t_5 inst_cell_111_111 (.BL(BL111),.BLN(BLN111),.WL(WL111));
sram_cell_6t_5 inst_cell_111_112 (.BL(BL112),.BLN(BLN112),.WL(WL111));
sram_cell_6t_5 inst_cell_111_113 (.BL(BL113),.BLN(BLN113),.WL(WL111));
sram_cell_6t_5 inst_cell_111_114 (.BL(BL114),.BLN(BLN114),.WL(WL111));
sram_cell_6t_5 inst_cell_111_115 (.BL(BL115),.BLN(BLN115),.WL(WL111));
sram_cell_6t_5 inst_cell_111_116 (.BL(BL116),.BLN(BLN116),.WL(WL111));
sram_cell_6t_5 inst_cell_111_117 (.BL(BL117),.BLN(BLN117),.WL(WL111));
sram_cell_6t_5 inst_cell_111_118 (.BL(BL118),.BLN(BLN118),.WL(WL111));
sram_cell_6t_5 inst_cell_111_119 (.BL(BL119),.BLN(BLN119),.WL(WL111));
sram_cell_6t_5 inst_cell_111_120 (.BL(BL120),.BLN(BLN120),.WL(WL111));
sram_cell_6t_5 inst_cell_111_121 (.BL(BL121),.BLN(BLN121),.WL(WL111));
sram_cell_6t_5 inst_cell_111_122 (.BL(BL122),.BLN(BLN122),.WL(WL111));
sram_cell_6t_5 inst_cell_111_123 (.BL(BL123),.BLN(BLN123),.WL(WL111));
sram_cell_6t_5 inst_cell_111_124 (.BL(BL124),.BLN(BLN124),.WL(WL111));
sram_cell_6t_5 inst_cell_111_125 (.BL(BL125),.BLN(BLN125),.WL(WL111));
sram_cell_6t_5 inst_cell_111_126 (.BL(BL126),.BLN(BLN126),.WL(WL111));
sram_cell_6t_5 inst_cell_111_127 (.BL(BL127),.BLN(BLN127),.WL(WL111));
sram_cell_6t_5 inst_cell_112_0 (.BL(BL0),.BLN(BLN0),.WL(WL112));
sram_cell_6t_5 inst_cell_112_1 (.BL(BL1),.BLN(BLN1),.WL(WL112));
sram_cell_6t_5 inst_cell_112_2 (.BL(BL2),.BLN(BLN2),.WL(WL112));
sram_cell_6t_5 inst_cell_112_3 (.BL(BL3),.BLN(BLN3),.WL(WL112));
sram_cell_6t_5 inst_cell_112_4 (.BL(BL4),.BLN(BLN4),.WL(WL112));
sram_cell_6t_5 inst_cell_112_5 (.BL(BL5),.BLN(BLN5),.WL(WL112));
sram_cell_6t_5 inst_cell_112_6 (.BL(BL6),.BLN(BLN6),.WL(WL112));
sram_cell_6t_5 inst_cell_112_7 (.BL(BL7),.BLN(BLN7),.WL(WL112));
sram_cell_6t_5 inst_cell_112_8 (.BL(BL8),.BLN(BLN8),.WL(WL112));
sram_cell_6t_5 inst_cell_112_9 (.BL(BL9),.BLN(BLN9),.WL(WL112));
sram_cell_6t_5 inst_cell_112_10 (.BL(BL10),.BLN(BLN10),.WL(WL112));
sram_cell_6t_5 inst_cell_112_11 (.BL(BL11),.BLN(BLN11),.WL(WL112));
sram_cell_6t_5 inst_cell_112_12 (.BL(BL12),.BLN(BLN12),.WL(WL112));
sram_cell_6t_5 inst_cell_112_13 (.BL(BL13),.BLN(BLN13),.WL(WL112));
sram_cell_6t_5 inst_cell_112_14 (.BL(BL14),.BLN(BLN14),.WL(WL112));
sram_cell_6t_5 inst_cell_112_15 (.BL(BL15),.BLN(BLN15),.WL(WL112));
sram_cell_6t_5 inst_cell_112_16 (.BL(BL16),.BLN(BLN16),.WL(WL112));
sram_cell_6t_5 inst_cell_112_17 (.BL(BL17),.BLN(BLN17),.WL(WL112));
sram_cell_6t_5 inst_cell_112_18 (.BL(BL18),.BLN(BLN18),.WL(WL112));
sram_cell_6t_5 inst_cell_112_19 (.BL(BL19),.BLN(BLN19),.WL(WL112));
sram_cell_6t_5 inst_cell_112_20 (.BL(BL20),.BLN(BLN20),.WL(WL112));
sram_cell_6t_5 inst_cell_112_21 (.BL(BL21),.BLN(BLN21),.WL(WL112));
sram_cell_6t_5 inst_cell_112_22 (.BL(BL22),.BLN(BLN22),.WL(WL112));
sram_cell_6t_5 inst_cell_112_23 (.BL(BL23),.BLN(BLN23),.WL(WL112));
sram_cell_6t_5 inst_cell_112_24 (.BL(BL24),.BLN(BLN24),.WL(WL112));
sram_cell_6t_5 inst_cell_112_25 (.BL(BL25),.BLN(BLN25),.WL(WL112));
sram_cell_6t_5 inst_cell_112_26 (.BL(BL26),.BLN(BLN26),.WL(WL112));
sram_cell_6t_5 inst_cell_112_27 (.BL(BL27),.BLN(BLN27),.WL(WL112));
sram_cell_6t_5 inst_cell_112_28 (.BL(BL28),.BLN(BLN28),.WL(WL112));
sram_cell_6t_5 inst_cell_112_29 (.BL(BL29),.BLN(BLN29),.WL(WL112));
sram_cell_6t_5 inst_cell_112_30 (.BL(BL30),.BLN(BLN30),.WL(WL112));
sram_cell_6t_5 inst_cell_112_31 (.BL(BL31),.BLN(BLN31),.WL(WL112));
sram_cell_6t_5 inst_cell_112_32 (.BL(BL32),.BLN(BLN32),.WL(WL112));
sram_cell_6t_5 inst_cell_112_33 (.BL(BL33),.BLN(BLN33),.WL(WL112));
sram_cell_6t_5 inst_cell_112_34 (.BL(BL34),.BLN(BLN34),.WL(WL112));
sram_cell_6t_5 inst_cell_112_35 (.BL(BL35),.BLN(BLN35),.WL(WL112));
sram_cell_6t_5 inst_cell_112_36 (.BL(BL36),.BLN(BLN36),.WL(WL112));
sram_cell_6t_5 inst_cell_112_37 (.BL(BL37),.BLN(BLN37),.WL(WL112));
sram_cell_6t_5 inst_cell_112_38 (.BL(BL38),.BLN(BLN38),.WL(WL112));
sram_cell_6t_5 inst_cell_112_39 (.BL(BL39),.BLN(BLN39),.WL(WL112));
sram_cell_6t_5 inst_cell_112_40 (.BL(BL40),.BLN(BLN40),.WL(WL112));
sram_cell_6t_5 inst_cell_112_41 (.BL(BL41),.BLN(BLN41),.WL(WL112));
sram_cell_6t_5 inst_cell_112_42 (.BL(BL42),.BLN(BLN42),.WL(WL112));
sram_cell_6t_5 inst_cell_112_43 (.BL(BL43),.BLN(BLN43),.WL(WL112));
sram_cell_6t_5 inst_cell_112_44 (.BL(BL44),.BLN(BLN44),.WL(WL112));
sram_cell_6t_5 inst_cell_112_45 (.BL(BL45),.BLN(BLN45),.WL(WL112));
sram_cell_6t_5 inst_cell_112_46 (.BL(BL46),.BLN(BLN46),.WL(WL112));
sram_cell_6t_5 inst_cell_112_47 (.BL(BL47),.BLN(BLN47),.WL(WL112));
sram_cell_6t_5 inst_cell_112_48 (.BL(BL48),.BLN(BLN48),.WL(WL112));
sram_cell_6t_5 inst_cell_112_49 (.BL(BL49),.BLN(BLN49),.WL(WL112));
sram_cell_6t_5 inst_cell_112_50 (.BL(BL50),.BLN(BLN50),.WL(WL112));
sram_cell_6t_5 inst_cell_112_51 (.BL(BL51),.BLN(BLN51),.WL(WL112));
sram_cell_6t_5 inst_cell_112_52 (.BL(BL52),.BLN(BLN52),.WL(WL112));
sram_cell_6t_5 inst_cell_112_53 (.BL(BL53),.BLN(BLN53),.WL(WL112));
sram_cell_6t_5 inst_cell_112_54 (.BL(BL54),.BLN(BLN54),.WL(WL112));
sram_cell_6t_5 inst_cell_112_55 (.BL(BL55),.BLN(BLN55),.WL(WL112));
sram_cell_6t_5 inst_cell_112_56 (.BL(BL56),.BLN(BLN56),.WL(WL112));
sram_cell_6t_5 inst_cell_112_57 (.BL(BL57),.BLN(BLN57),.WL(WL112));
sram_cell_6t_5 inst_cell_112_58 (.BL(BL58),.BLN(BLN58),.WL(WL112));
sram_cell_6t_5 inst_cell_112_59 (.BL(BL59),.BLN(BLN59),.WL(WL112));
sram_cell_6t_5 inst_cell_112_60 (.BL(BL60),.BLN(BLN60),.WL(WL112));
sram_cell_6t_5 inst_cell_112_61 (.BL(BL61),.BLN(BLN61),.WL(WL112));
sram_cell_6t_5 inst_cell_112_62 (.BL(BL62),.BLN(BLN62),.WL(WL112));
sram_cell_6t_5 inst_cell_112_63 (.BL(BL63),.BLN(BLN63),.WL(WL112));
sram_cell_6t_5 inst_cell_112_64 (.BL(BL64),.BLN(BLN64),.WL(WL112));
sram_cell_6t_5 inst_cell_112_65 (.BL(BL65),.BLN(BLN65),.WL(WL112));
sram_cell_6t_5 inst_cell_112_66 (.BL(BL66),.BLN(BLN66),.WL(WL112));
sram_cell_6t_5 inst_cell_112_67 (.BL(BL67),.BLN(BLN67),.WL(WL112));
sram_cell_6t_5 inst_cell_112_68 (.BL(BL68),.BLN(BLN68),.WL(WL112));
sram_cell_6t_5 inst_cell_112_69 (.BL(BL69),.BLN(BLN69),.WL(WL112));
sram_cell_6t_5 inst_cell_112_70 (.BL(BL70),.BLN(BLN70),.WL(WL112));
sram_cell_6t_5 inst_cell_112_71 (.BL(BL71),.BLN(BLN71),.WL(WL112));
sram_cell_6t_5 inst_cell_112_72 (.BL(BL72),.BLN(BLN72),.WL(WL112));
sram_cell_6t_5 inst_cell_112_73 (.BL(BL73),.BLN(BLN73),.WL(WL112));
sram_cell_6t_5 inst_cell_112_74 (.BL(BL74),.BLN(BLN74),.WL(WL112));
sram_cell_6t_5 inst_cell_112_75 (.BL(BL75),.BLN(BLN75),.WL(WL112));
sram_cell_6t_5 inst_cell_112_76 (.BL(BL76),.BLN(BLN76),.WL(WL112));
sram_cell_6t_5 inst_cell_112_77 (.BL(BL77),.BLN(BLN77),.WL(WL112));
sram_cell_6t_5 inst_cell_112_78 (.BL(BL78),.BLN(BLN78),.WL(WL112));
sram_cell_6t_5 inst_cell_112_79 (.BL(BL79),.BLN(BLN79),.WL(WL112));
sram_cell_6t_5 inst_cell_112_80 (.BL(BL80),.BLN(BLN80),.WL(WL112));
sram_cell_6t_5 inst_cell_112_81 (.BL(BL81),.BLN(BLN81),.WL(WL112));
sram_cell_6t_5 inst_cell_112_82 (.BL(BL82),.BLN(BLN82),.WL(WL112));
sram_cell_6t_5 inst_cell_112_83 (.BL(BL83),.BLN(BLN83),.WL(WL112));
sram_cell_6t_5 inst_cell_112_84 (.BL(BL84),.BLN(BLN84),.WL(WL112));
sram_cell_6t_5 inst_cell_112_85 (.BL(BL85),.BLN(BLN85),.WL(WL112));
sram_cell_6t_5 inst_cell_112_86 (.BL(BL86),.BLN(BLN86),.WL(WL112));
sram_cell_6t_5 inst_cell_112_87 (.BL(BL87),.BLN(BLN87),.WL(WL112));
sram_cell_6t_5 inst_cell_112_88 (.BL(BL88),.BLN(BLN88),.WL(WL112));
sram_cell_6t_5 inst_cell_112_89 (.BL(BL89),.BLN(BLN89),.WL(WL112));
sram_cell_6t_5 inst_cell_112_90 (.BL(BL90),.BLN(BLN90),.WL(WL112));
sram_cell_6t_5 inst_cell_112_91 (.BL(BL91),.BLN(BLN91),.WL(WL112));
sram_cell_6t_5 inst_cell_112_92 (.BL(BL92),.BLN(BLN92),.WL(WL112));
sram_cell_6t_5 inst_cell_112_93 (.BL(BL93),.BLN(BLN93),.WL(WL112));
sram_cell_6t_5 inst_cell_112_94 (.BL(BL94),.BLN(BLN94),.WL(WL112));
sram_cell_6t_5 inst_cell_112_95 (.BL(BL95),.BLN(BLN95),.WL(WL112));
sram_cell_6t_5 inst_cell_112_96 (.BL(BL96),.BLN(BLN96),.WL(WL112));
sram_cell_6t_5 inst_cell_112_97 (.BL(BL97),.BLN(BLN97),.WL(WL112));
sram_cell_6t_5 inst_cell_112_98 (.BL(BL98),.BLN(BLN98),.WL(WL112));
sram_cell_6t_5 inst_cell_112_99 (.BL(BL99),.BLN(BLN99),.WL(WL112));
sram_cell_6t_5 inst_cell_112_100 (.BL(BL100),.BLN(BLN100),.WL(WL112));
sram_cell_6t_5 inst_cell_112_101 (.BL(BL101),.BLN(BLN101),.WL(WL112));
sram_cell_6t_5 inst_cell_112_102 (.BL(BL102),.BLN(BLN102),.WL(WL112));
sram_cell_6t_5 inst_cell_112_103 (.BL(BL103),.BLN(BLN103),.WL(WL112));
sram_cell_6t_5 inst_cell_112_104 (.BL(BL104),.BLN(BLN104),.WL(WL112));
sram_cell_6t_5 inst_cell_112_105 (.BL(BL105),.BLN(BLN105),.WL(WL112));
sram_cell_6t_5 inst_cell_112_106 (.BL(BL106),.BLN(BLN106),.WL(WL112));
sram_cell_6t_5 inst_cell_112_107 (.BL(BL107),.BLN(BLN107),.WL(WL112));
sram_cell_6t_5 inst_cell_112_108 (.BL(BL108),.BLN(BLN108),.WL(WL112));
sram_cell_6t_5 inst_cell_112_109 (.BL(BL109),.BLN(BLN109),.WL(WL112));
sram_cell_6t_5 inst_cell_112_110 (.BL(BL110),.BLN(BLN110),.WL(WL112));
sram_cell_6t_5 inst_cell_112_111 (.BL(BL111),.BLN(BLN111),.WL(WL112));
sram_cell_6t_5 inst_cell_112_112 (.BL(BL112),.BLN(BLN112),.WL(WL112));
sram_cell_6t_5 inst_cell_112_113 (.BL(BL113),.BLN(BLN113),.WL(WL112));
sram_cell_6t_5 inst_cell_112_114 (.BL(BL114),.BLN(BLN114),.WL(WL112));
sram_cell_6t_5 inst_cell_112_115 (.BL(BL115),.BLN(BLN115),.WL(WL112));
sram_cell_6t_5 inst_cell_112_116 (.BL(BL116),.BLN(BLN116),.WL(WL112));
sram_cell_6t_5 inst_cell_112_117 (.BL(BL117),.BLN(BLN117),.WL(WL112));
sram_cell_6t_5 inst_cell_112_118 (.BL(BL118),.BLN(BLN118),.WL(WL112));
sram_cell_6t_5 inst_cell_112_119 (.BL(BL119),.BLN(BLN119),.WL(WL112));
sram_cell_6t_5 inst_cell_112_120 (.BL(BL120),.BLN(BLN120),.WL(WL112));
sram_cell_6t_5 inst_cell_112_121 (.BL(BL121),.BLN(BLN121),.WL(WL112));
sram_cell_6t_5 inst_cell_112_122 (.BL(BL122),.BLN(BLN122),.WL(WL112));
sram_cell_6t_5 inst_cell_112_123 (.BL(BL123),.BLN(BLN123),.WL(WL112));
sram_cell_6t_5 inst_cell_112_124 (.BL(BL124),.BLN(BLN124),.WL(WL112));
sram_cell_6t_5 inst_cell_112_125 (.BL(BL125),.BLN(BLN125),.WL(WL112));
sram_cell_6t_5 inst_cell_112_126 (.BL(BL126),.BLN(BLN126),.WL(WL112));
sram_cell_6t_5 inst_cell_112_127 (.BL(BL127),.BLN(BLN127),.WL(WL112));
sram_cell_6t_5 inst_cell_113_0 (.BL(BL0),.BLN(BLN0),.WL(WL113));
sram_cell_6t_5 inst_cell_113_1 (.BL(BL1),.BLN(BLN1),.WL(WL113));
sram_cell_6t_5 inst_cell_113_2 (.BL(BL2),.BLN(BLN2),.WL(WL113));
sram_cell_6t_5 inst_cell_113_3 (.BL(BL3),.BLN(BLN3),.WL(WL113));
sram_cell_6t_5 inst_cell_113_4 (.BL(BL4),.BLN(BLN4),.WL(WL113));
sram_cell_6t_5 inst_cell_113_5 (.BL(BL5),.BLN(BLN5),.WL(WL113));
sram_cell_6t_5 inst_cell_113_6 (.BL(BL6),.BLN(BLN6),.WL(WL113));
sram_cell_6t_5 inst_cell_113_7 (.BL(BL7),.BLN(BLN7),.WL(WL113));
sram_cell_6t_5 inst_cell_113_8 (.BL(BL8),.BLN(BLN8),.WL(WL113));
sram_cell_6t_5 inst_cell_113_9 (.BL(BL9),.BLN(BLN9),.WL(WL113));
sram_cell_6t_5 inst_cell_113_10 (.BL(BL10),.BLN(BLN10),.WL(WL113));
sram_cell_6t_5 inst_cell_113_11 (.BL(BL11),.BLN(BLN11),.WL(WL113));
sram_cell_6t_5 inst_cell_113_12 (.BL(BL12),.BLN(BLN12),.WL(WL113));
sram_cell_6t_5 inst_cell_113_13 (.BL(BL13),.BLN(BLN13),.WL(WL113));
sram_cell_6t_5 inst_cell_113_14 (.BL(BL14),.BLN(BLN14),.WL(WL113));
sram_cell_6t_5 inst_cell_113_15 (.BL(BL15),.BLN(BLN15),.WL(WL113));
sram_cell_6t_5 inst_cell_113_16 (.BL(BL16),.BLN(BLN16),.WL(WL113));
sram_cell_6t_5 inst_cell_113_17 (.BL(BL17),.BLN(BLN17),.WL(WL113));
sram_cell_6t_5 inst_cell_113_18 (.BL(BL18),.BLN(BLN18),.WL(WL113));
sram_cell_6t_5 inst_cell_113_19 (.BL(BL19),.BLN(BLN19),.WL(WL113));
sram_cell_6t_5 inst_cell_113_20 (.BL(BL20),.BLN(BLN20),.WL(WL113));
sram_cell_6t_5 inst_cell_113_21 (.BL(BL21),.BLN(BLN21),.WL(WL113));
sram_cell_6t_5 inst_cell_113_22 (.BL(BL22),.BLN(BLN22),.WL(WL113));
sram_cell_6t_5 inst_cell_113_23 (.BL(BL23),.BLN(BLN23),.WL(WL113));
sram_cell_6t_5 inst_cell_113_24 (.BL(BL24),.BLN(BLN24),.WL(WL113));
sram_cell_6t_5 inst_cell_113_25 (.BL(BL25),.BLN(BLN25),.WL(WL113));
sram_cell_6t_5 inst_cell_113_26 (.BL(BL26),.BLN(BLN26),.WL(WL113));
sram_cell_6t_5 inst_cell_113_27 (.BL(BL27),.BLN(BLN27),.WL(WL113));
sram_cell_6t_5 inst_cell_113_28 (.BL(BL28),.BLN(BLN28),.WL(WL113));
sram_cell_6t_5 inst_cell_113_29 (.BL(BL29),.BLN(BLN29),.WL(WL113));
sram_cell_6t_5 inst_cell_113_30 (.BL(BL30),.BLN(BLN30),.WL(WL113));
sram_cell_6t_5 inst_cell_113_31 (.BL(BL31),.BLN(BLN31),.WL(WL113));
sram_cell_6t_5 inst_cell_113_32 (.BL(BL32),.BLN(BLN32),.WL(WL113));
sram_cell_6t_5 inst_cell_113_33 (.BL(BL33),.BLN(BLN33),.WL(WL113));
sram_cell_6t_5 inst_cell_113_34 (.BL(BL34),.BLN(BLN34),.WL(WL113));
sram_cell_6t_5 inst_cell_113_35 (.BL(BL35),.BLN(BLN35),.WL(WL113));
sram_cell_6t_5 inst_cell_113_36 (.BL(BL36),.BLN(BLN36),.WL(WL113));
sram_cell_6t_5 inst_cell_113_37 (.BL(BL37),.BLN(BLN37),.WL(WL113));
sram_cell_6t_5 inst_cell_113_38 (.BL(BL38),.BLN(BLN38),.WL(WL113));
sram_cell_6t_5 inst_cell_113_39 (.BL(BL39),.BLN(BLN39),.WL(WL113));
sram_cell_6t_5 inst_cell_113_40 (.BL(BL40),.BLN(BLN40),.WL(WL113));
sram_cell_6t_5 inst_cell_113_41 (.BL(BL41),.BLN(BLN41),.WL(WL113));
sram_cell_6t_5 inst_cell_113_42 (.BL(BL42),.BLN(BLN42),.WL(WL113));
sram_cell_6t_5 inst_cell_113_43 (.BL(BL43),.BLN(BLN43),.WL(WL113));
sram_cell_6t_5 inst_cell_113_44 (.BL(BL44),.BLN(BLN44),.WL(WL113));
sram_cell_6t_5 inst_cell_113_45 (.BL(BL45),.BLN(BLN45),.WL(WL113));
sram_cell_6t_5 inst_cell_113_46 (.BL(BL46),.BLN(BLN46),.WL(WL113));
sram_cell_6t_5 inst_cell_113_47 (.BL(BL47),.BLN(BLN47),.WL(WL113));
sram_cell_6t_5 inst_cell_113_48 (.BL(BL48),.BLN(BLN48),.WL(WL113));
sram_cell_6t_5 inst_cell_113_49 (.BL(BL49),.BLN(BLN49),.WL(WL113));
sram_cell_6t_5 inst_cell_113_50 (.BL(BL50),.BLN(BLN50),.WL(WL113));
sram_cell_6t_5 inst_cell_113_51 (.BL(BL51),.BLN(BLN51),.WL(WL113));
sram_cell_6t_5 inst_cell_113_52 (.BL(BL52),.BLN(BLN52),.WL(WL113));
sram_cell_6t_5 inst_cell_113_53 (.BL(BL53),.BLN(BLN53),.WL(WL113));
sram_cell_6t_5 inst_cell_113_54 (.BL(BL54),.BLN(BLN54),.WL(WL113));
sram_cell_6t_5 inst_cell_113_55 (.BL(BL55),.BLN(BLN55),.WL(WL113));
sram_cell_6t_5 inst_cell_113_56 (.BL(BL56),.BLN(BLN56),.WL(WL113));
sram_cell_6t_5 inst_cell_113_57 (.BL(BL57),.BLN(BLN57),.WL(WL113));
sram_cell_6t_5 inst_cell_113_58 (.BL(BL58),.BLN(BLN58),.WL(WL113));
sram_cell_6t_5 inst_cell_113_59 (.BL(BL59),.BLN(BLN59),.WL(WL113));
sram_cell_6t_5 inst_cell_113_60 (.BL(BL60),.BLN(BLN60),.WL(WL113));
sram_cell_6t_5 inst_cell_113_61 (.BL(BL61),.BLN(BLN61),.WL(WL113));
sram_cell_6t_5 inst_cell_113_62 (.BL(BL62),.BLN(BLN62),.WL(WL113));
sram_cell_6t_5 inst_cell_113_63 (.BL(BL63),.BLN(BLN63),.WL(WL113));
sram_cell_6t_5 inst_cell_113_64 (.BL(BL64),.BLN(BLN64),.WL(WL113));
sram_cell_6t_5 inst_cell_113_65 (.BL(BL65),.BLN(BLN65),.WL(WL113));
sram_cell_6t_5 inst_cell_113_66 (.BL(BL66),.BLN(BLN66),.WL(WL113));
sram_cell_6t_5 inst_cell_113_67 (.BL(BL67),.BLN(BLN67),.WL(WL113));
sram_cell_6t_5 inst_cell_113_68 (.BL(BL68),.BLN(BLN68),.WL(WL113));
sram_cell_6t_5 inst_cell_113_69 (.BL(BL69),.BLN(BLN69),.WL(WL113));
sram_cell_6t_5 inst_cell_113_70 (.BL(BL70),.BLN(BLN70),.WL(WL113));
sram_cell_6t_5 inst_cell_113_71 (.BL(BL71),.BLN(BLN71),.WL(WL113));
sram_cell_6t_5 inst_cell_113_72 (.BL(BL72),.BLN(BLN72),.WL(WL113));
sram_cell_6t_5 inst_cell_113_73 (.BL(BL73),.BLN(BLN73),.WL(WL113));
sram_cell_6t_5 inst_cell_113_74 (.BL(BL74),.BLN(BLN74),.WL(WL113));
sram_cell_6t_5 inst_cell_113_75 (.BL(BL75),.BLN(BLN75),.WL(WL113));
sram_cell_6t_5 inst_cell_113_76 (.BL(BL76),.BLN(BLN76),.WL(WL113));
sram_cell_6t_5 inst_cell_113_77 (.BL(BL77),.BLN(BLN77),.WL(WL113));
sram_cell_6t_5 inst_cell_113_78 (.BL(BL78),.BLN(BLN78),.WL(WL113));
sram_cell_6t_5 inst_cell_113_79 (.BL(BL79),.BLN(BLN79),.WL(WL113));
sram_cell_6t_5 inst_cell_113_80 (.BL(BL80),.BLN(BLN80),.WL(WL113));
sram_cell_6t_5 inst_cell_113_81 (.BL(BL81),.BLN(BLN81),.WL(WL113));
sram_cell_6t_5 inst_cell_113_82 (.BL(BL82),.BLN(BLN82),.WL(WL113));
sram_cell_6t_5 inst_cell_113_83 (.BL(BL83),.BLN(BLN83),.WL(WL113));
sram_cell_6t_5 inst_cell_113_84 (.BL(BL84),.BLN(BLN84),.WL(WL113));
sram_cell_6t_5 inst_cell_113_85 (.BL(BL85),.BLN(BLN85),.WL(WL113));
sram_cell_6t_5 inst_cell_113_86 (.BL(BL86),.BLN(BLN86),.WL(WL113));
sram_cell_6t_5 inst_cell_113_87 (.BL(BL87),.BLN(BLN87),.WL(WL113));
sram_cell_6t_5 inst_cell_113_88 (.BL(BL88),.BLN(BLN88),.WL(WL113));
sram_cell_6t_5 inst_cell_113_89 (.BL(BL89),.BLN(BLN89),.WL(WL113));
sram_cell_6t_5 inst_cell_113_90 (.BL(BL90),.BLN(BLN90),.WL(WL113));
sram_cell_6t_5 inst_cell_113_91 (.BL(BL91),.BLN(BLN91),.WL(WL113));
sram_cell_6t_5 inst_cell_113_92 (.BL(BL92),.BLN(BLN92),.WL(WL113));
sram_cell_6t_5 inst_cell_113_93 (.BL(BL93),.BLN(BLN93),.WL(WL113));
sram_cell_6t_5 inst_cell_113_94 (.BL(BL94),.BLN(BLN94),.WL(WL113));
sram_cell_6t_5 inst_cell_113_95 (.BL(BL95),.BLN(BLN95),.WL(WL113));
sram_cell_6t_5 inst_cell_113_96 (.BL(BL96),.BLN(BLN96),.WL(WL113));
sram_cell_6t_5 inst_cell_113_97 (.BL(BL97),.BLN(BLN97),.WL(WL113));
sram_cell_6t_5 inst_cell_113_98 (.BL(BL98),.BLN(BLN98),.WL(WL113));
sram_cell_6t_5 inst_cell_113_99 (.BL(BL99),.BLN(BLN99),.WL(WL113));
sram_cell_6t_5 inst_cell_113_100 (.BL(BL100),.BLN(BLN100),.WL(WL113));
sram_cell_6t_5 inst_cell_113_101 (.BL(BL101),.BLN(BLN101),.WL(WL113));
sram_cell_6t_5 inst_cell_113_102 (.BL(BL102),.BLN(BLN102),.WL(WL113));
sram_cell_6t_5 inst_cell_113_103 (.BL(BL103),.BLN(BLN103),.WL(WL113));
sram_cell_6t_5 inst_cell_113_104 (.BL(BL104),.BLN(BLN104),.WL(WL113));
sram_cell_6t_5 inst_cell_113_105 (.BL(BL105),.BLN(BLN105),.WL(WL113));
sram_cell_6t_5 inst_cell_113_106 (.BL(BL106),.BLN(BLN106),.WL(WL113));
sram_cell_6t_5 inst_cell_113_107 (.BL(BL107),.BLN(BLN107),.WL(WL113));
sram_cell_6t_5 inst_cell_113_108 (.BL(BL108),.BLN(BLN108),.WL(WL113));
sram_cell_6t_5 inst_cell_113_109 (.BL(BL109),.BLN(BLN109),.WL(WL113));
sram_cell_6t_5 inst_cell_113_110 (.BL(BL110),.BLN(BLN110),.WL(WL113));
sram_cell_6t_5 inst_cell_113_111 (.BL(BL111),.BLN(BLN111),.WL(WL113));
sram_cell_6t_5 inst_cell_113_112 (.BL(BL112),.BLN(BLN112),.WL(WL113));
sram_cell_6t_5 inst_cell_113_113 (.BL(BL113),.BLN(BLN113),.WL(WL113));
sram_cell_6t_5 inst_cell_113_114 (.BL(BL114),.BLN(BLN114),.WL(WL113));
sram_cell_6t_5 inst_cell_113_115 (.BL(BL115),.BLN(BLN115),.WL(WL113));
sram_cell_6t_5 inst_cell_113_116 (.BL(BL116),.BLN(BLN116),.WL(WL113));
sram_cell_6t_5 inst_cell_113_117 (.BL(BL117),.BLN(BLN117),.WL(WL113));
sram_cell_6t_5 inst_cell_113_118 (.BL(BL118),.BLN(BLN118),.WL(WL113));
sram_cell_6t_5 inst_cell_113_119 (.BL(BL119),.BLN(BLN119),.WL(WL113));
sram_cell_6t_5 inst_cell_113_120 (.BL(BL120),.BLN(BLN120),.WL(WL113));
sram_cell_6t_5 inst_cell_113_121 (.BL(BL121),.BLN(BLN121),.WL(WL113));
sram_cell_6t_5 inst_cell_113_122 (.BL(BL122),.BLN(BLN122),.WL(WL113));
sram_cell_6t_5 inst_cell_113_123 (.BL(BL123),.BLN(BLN123),.WL(WL113));
sram_cell_6t_5 inst_cell_113_124 (.BL(BL124),.BLN(BLN124),.WL(WL113));
sram_cell_6t_5 inst_cell_113_125 (.BL(BL125),.BLN(BLN125),.WL(WL113));
sram_cell_6t_5 inst_cell_113_126 (.BL(BL126),.BLN(BLN126),.WL(WL113));
sram_cell_6t_5 inst_cell_113_127 (.BL(BL127),.BLN(BLN127),.WL(WL113));
sram_cell_6t_5 inst_cell_114_0 (.BL(BL0),.BLN(BLN0),.WL(WL114));
sram_cell_6t_5 inst_cell_114_1 (.BL(BL1),.BLN(BLN1),.WL(WL114));
sram_cell_6t_5 inst_cell_114_2 (.BL(BL2),.BLN(BLN2),.WL(WL114));
sram_cell_6t_5 inst_cell_114_3 (.BL(BL3),.BLN(BLN3),.WL(WL114));
sram_cell_6t_5 inst_cell_114_4 (.BL(BL4),.BLN(BLN4),.WL(WL114));
sram_cell_6t_5 inst_cell_114_5 (.BL(BL5),.BLN(BLN5),.WL(WL114));
sram_cell_6t_5 inst_cell_114_6 (.BL(BL6),.BLN(BLN6),.WL(WL114));
sram_cell_6t_5 inst_cell_114_7 (.BL(BL7),.BLN(BLN7),.WL(WL114));
sram_cell_6t_5 inst_cell_114_8 (.BL(BL8),.BLN(BLN8),.WL(WL114));
sram_cell_6t_5 inst_cell_114_9 (.BL(BL9),.BLN(BLN9),.WL(WL114));
sram_cell_6t_5 inst_cell_114_10 (.BL(BL10),.BLN(BLN10),.WL(WL114));
sram_cell_6t_5 inst_cell_114_11 (.BL(BL11),.BLN(BLN11),.WL(WL114));
sram_cell_6t_5 inst_cell_114_12 (.BL(BL12),.BLN(BLN12),.WL(WL114));
sram_cell_6t_5 inst_cell_114_13 (.BL(BL13),.BLN(BLN13),.WL(WL114));
sram_cell_6t_5 inst_cell_114_14 (.BL(BL14),.BLN(BLN14),.WL(WL114));
sram_cell_6t_5 inst_cell_114_15 (.BL(BL15),.BLN(BLN15),.WL(WL114));
sram_cell_6t_5 inst_cell_114_16 (.BL(BL16),.BLN(BLN16),.WL(WL114));
sram_cell_6t_5 inst_cell_114_17 (.BL(BL17),.BLN(BLN17),.WL(WL114));
sram_cell_6t_5 inst_cell_114_18 (.BL(BL18),.BLN(BLN18),.WL(WL114));
sram_cell_6t_5 inst_cell_114_19 (.BL(BL19),.BLN(BLN19),.WL(WL114));
sram_cell_6t_5 inst_cell_114_20 (.BL(BL20),.BLN(BLN20),.WL(WL114));
sram_cell_6t_5 inst_cell_114_21 (.BL(BL21),.BLN(BLN21),.WL(WL114));
sram_cell_6t_5 inst_cell_114_22 (.BL(BL22),.BLN(BLN22),.WL(WL114));
sram_cell_6t_5 inst_cell_114_23 (.BL(BL23),.BLN(BLN23),.WL(WL114));
sram_cell_6t_5 inst_cell_114_24 (.BL(BL24),.BLN(BLN24),.WL(WL114));
sram_cell_6t_5 inst_cell_114_25 (.BL(BL25),.BLN(BLN25),.WL(WL114));
sram_cell_6t_5 inst_cell_114_26 (.BL(BL26),.BLN(BLN26),.WL(WL114));
sram_cell_6t_5 inst_cell_114_27 (.BL(BL27),.BLN(BLN27),.WL(WL114));
sram_cell_6t_5 inst_cell_114_28 (.BL(BL28),.BLN(BLN28),.WL(WL114));
sram_cell_6t_5 inst_cell_114_29 (.BL(BL29),.BLN(BLN29),.WL(WL114));
sram_cell_6t_5 inst_cell_114_30 (.BL(BL30),.BLN(BLN30),.WL(WL114));
sram_cell_6t_5 inst_cell_114_31 (.BL(BL31),.BLN(BLN31),.WL(WL114));
sram_cell_6t_5 inst_cell_114_32 (.BL(BL32),.BLN(BLN32),.WL(WL114));
sram_cell_6t_5 inst_cell_114_33 (.BL(BL33),.BLN(BLN33),.WL(WL114));
sram_cell_6t_5 inst_cell_114_34 (.BL(BL34),.BLN(BLN34),.WL(WL114));
sram_cell_6t_5 inst_cell_114_35 (.BL(BL35),.BLN(BLN35),.WL(WL114));
sram_cell_6t_5 inst_cell_114_36 (.BL(BL36),.BLN(BLN36),.WL(WL114));
sram_cell_6t_5 inst_cell_114_37 (.BL(BL37),.BLN(BLN37),.WL(WL114));
sram_cell_6t_5 inst_cell_114_38 (.BL(BL38),.BLN(BLN38),.WL(WL114));
sram_cell_6t_5 inst_cell_114_39 (.BL(BL39),.BLN(BLN39),.WL(WL114));
sram_cell_6t_5 inst_cell_114_40 (.BL(BL40),.BLN(BLN40),.WL(WL114));
sram_cell_6t_5 inst_cell_114_41 (.BL(BL41),.BLN(BLN41),.WL(WL114));
sram_cell_6t_5 inst_cell_114_42 (.BL(BL42),.BLN(BLN42),.WL(WL114));
sram_cell_6t_5 inst_cell_114_43 (.BL(BL43),.BLN(BLN43),.WL(WL114));
sram_cell_6t_5 inst_cell_114_44 (.BL(BL44),.BLN(BLN44),.WL(WL114));
sram_cell_6t_5 inst_cell_114_45 (.BL(BL45),.BLN(BLN45),.WL(WL114));
sram_cell_6t_5 inst_cell_114_46 (.BL(BL46),.BLN(BLN46),.WL(WL114));
sram_cell_6t_5 inst_cell_114_47 (.BL(BL47),.BLN(BLN47),.WL(WL114));
sram_cell_6t_5 inst_cell_114_48 (.BL(BL48),.BLN(BLN48),.WL(WL114));
sram_cell_6t_5 inst_cell_114_49 (.BL(BL49),.BLN(BLN49),.WL(WL114));
sram_cell_6t_5 inst_cell_114_50 (.BL(BL50),.BLN(BLN50),.WL(WL114));
sram_cell_6t_5 inst_cell_114_51 (.BL(BL51),.BLN(BLN51),.WL(WL114));
sram_cell_6t_5 inst_cell_114_52 (.BL(BL52),.BLN(BLN52),.WL(WL114));
sram_cell_6t_5 inst_cell_114_53 (.BL(BL53),.BLN(BLN53),.WL(WL114));
sram_cell_6t_5 inst_cell_114_54 (.BL(BL54),.BLN(BLN54),.WL(WL114));
sram_cell_6t_5 inst_cell_114_55 (.BL(BL55),.BLN(BLN55),.WL(WL114));
sram_cell_6t_5 inst_cell_114_56 (.BL(BL56),.BLN(BLN56),.WL(WL114));
sram_cell_6t_5 inst_cell_114_57 (.BL(BL57),.BLN(BLN57),.WL(WL114));
sram_cell_6t_5 inst_cell_114_58 (.BL(BL58),.BLN(BLN58),.WL(WL114));
sram_cell_6t_5 inst_cell_114_59 (.BL(BL59),.BLN(BLN59),.WL(WL114));
sram_cell_6t_5 inst_cell_114_60 (.BL(BL60),.BLN(BLN60),.WL(WL114));
sram_cell_6t_5 inst_cell_114_61 (.BL(BL61),.BLN(BLN61),.WL(WL114));
sram_cell_6t_5 inst_cell_114_62 (.BL(BL62),.BLN(BLN62),.WL(WL114));
sram_cell_6t_5 inst_cell_114_63 (.BL(BL63),.BLN(BLN63),.WL(WL114));
sram_cell_6t_5 inst_cell_114_64 (.BL(BL64),.BLN(BLN64),.WL(WL114));
sram_cell_6t_5 inst_cell_114_65 (.BL(BL65),.BLN(BLN65),.WL(WL114));
sram_cell_6t_5 inst_cell_114_66 (.BL(BL66),.BLN(BLN66),.WL(WL114));
sram_cell_6t_5 inst_cell_114_67 (.BL(BL67),.BLN(BLN67),.WL(WL114));
sram_cell_6t_5 inst_cell_114_68 (.BL(BL68),.BLN(BLN68),.WL(WL114));
sram_cell_6t_5 inst_cell_114_69 (.BL(BL69),.BLN(BLN69),.WL(WL114));
sram_cell_6t_5 inst_cell_114_70 (.BL(BL70),.BLN(BLN70),.WL(WL114));
sram_cell_6t_5 inst_cell_114_71 (.BL(BL71),.BLN(BLN71),.WL(WL114));
sram_cell_6t_5 inst_cell_114_72 (.BL(BL72),.BLN(BLN72),.WL(WL114));
sram_cell_6t_5 inst_cell_114_73 (.BL(BL73),.BLN(BLN73),.WL(WL114));
sram_cell_6t_5 inst_cell_114_74 (.BL(BL74),.BLN(BLN74),.WL(WL114));
sram_cell_6t_5 inst_cell_114_75 (.BL(BL75),.BLN(BLN75),.WL(WL114));
sram_cell_6t_5 inst_cell_114_76 (.BL(BL76),.BLN(BLN76),.WL(WL114));
sram_cell_6t_5 inst_cell_114_77 (.BL(BL77),.BLN(BLN77),.WL(WL114));
sram_cell_6t_5 inst_cell_114_78 (.BL(BL78),.BLN(BLN78),.WL(WL114));
sram_cell_6t_5 inst_cell_114_79 (.BL(BL79),.BLN(BLN79),.WL(WL114));
sram_cell_6t_5 inst_cell_114_80 (.BL(BL80),.BLN(BLN80),.WL(WL114));
sram_cell_6t_5 inst_cell_114_81 (.BL(BL81),.BLN(BLN81),.WL(WL114));
sram_cell_6t_5 inst_cell_114_82 (.BL(BL82),.BLN(BLN82),.WL(WL114));
sram_cell_6t_5 inst_cell_114_83 (.BL(BL83),.BLN(BLN83),.WL(WL114));
sram_cell_6t_5 inst_cell_114_84 (.BL(BL84),.BLN(BLN84),.WL(WL114));
sram_cell_6t_5 inst_cell_114_85 (.BL(BL85),.BLN(BLN85),.WL(WL114));
sram_cell_6t_5 inst_cell_114_86 (.BL(BL86),.BLN(BLN86),.WL(WL114));
sram_cell_6t_5 inst_cell_114_87 (.BL(BL87),.BLN(BLN87),.WL(WL114));
sram_cell_6t_5 inst_cell_114_88 (.BL(BL88),.BLN(BLN88),.WL(WL114));
sram_cell_6t_5 inst_cell_114_89 (.BL(BL89),.BLN(BLN89),.WL(WL114));
sram_cell_6t_5 inst_cell_114_90 (.BL(BL90),.BLN(BLN90),.WL(WL114));
sram_cell_6t_5 inst_cell_114_91 (.BL(BL91),.BLN(BLN91),.WL(WL114));
sram_cell_6t_5 inst_cell_114_92 (.BL(BL92),.BLN(BLN92),.WL(WL114));
sram_cell_6t_5 inst_cell_114_93 (.BL(BL93),.BLN(BLN93),.WL(WL114));
sram_cell_6t_5 inst_cell_114_94 (.BL(BL94),.BLN(BLN94),.WL(WL114));
sram_cell_6t_5 inst_cell_114_95 (.BL(BL95),.BLN(BLN95),.WL(WL114));
sram_cell_6t_5 inst_cell_114_96 (.BL(BL96),.BLN(BLN96),.WL(WL114));
sram_cell_6t_5 inst_cell_114_97 (.BL(BL97),.BLN(BLN97),.WL(WL114));
sram_cell_6t_5 inst_cell_114_98 (.BL(BL98),.BLN(BLN98),.WL(WL114));
sram_cell_6t_5 inst_cell_114_99 (.BL(BL99),.BLN(BLN99),.WL(WL114));
sram_cell_6t_5 inst_cell_114_100 (.BL(BL100),.BLN(BLN100),.WL(WL114));
sram_cell_6t_5 inst_cell_114_101 (.BL(BL101),.BLN(BLN101),.WL(WL114));
sram_cell_6t_5 inst_cell_114_102 (.BL(BL102),.BLN(BLN102),.WL(WL114));
sram_cell_6t_5 inst_cell_114_103 (.BL(BL103),.BLN(BLN103),.WL(WL114));
sram_cell_6t_5 inst_cell_114_104 (.BL(BL104),.BLN(BLN104),.WL(WL114));
sram_cell_6t_5 inst_cell_114_105 (.BL(BL105),.BLN(BLN105),.WL(WL114));
sram_cell_6t_5 inst_cell_114_106 (.BL(BL106),.BLN(BLN106),.WL(WL114));
sram_cell_6t_5 inst_cell_114_107 (.BL(BL107),.BLN(BLN107),.WL(WL114));
sram_cell_6t_5 inst_cell_114_108 (.BL(BL108),.BLN(BLN108),.WL(WL114));
sram_cell_6t_5 inst_cell_114_109 (.BL(BL109),.BLN(BLN109),.WL(WL114));
sram_cell_6t_5 inst_cell_114_110 (.BL(BL110),.BLN(BLN110),.WL(WL114));
sram_cell_6t_5 inst_cell_114_111 (.BL(BL111),.BLN(BLN111),.WL(WL114));
sram_cell_6t_5 inst_cell_114_112 (.BL(BL112),.BLN(BLN112),.WL(WL114));
sram_cell_6t_5 inst_cell_114_113 (.BL(BL113),.BLN(BLN113),.WL(WL114));
sram_cell_6t_5 inst_cell_114_114 (.BL(BL114),.BLN(BLN114),.WL(WL114));
sram_cell_6t_5 inst_cell_114_115 (.BL(BL115),.BLN(BLN115),.WL(WL114));
sram_cell_6t_5 inst_cell_114_116 (.BL(BL116),.BLN(BLN116),.WL(WL114));
sram_cell_6t_5 inst_cell_114_117 (.BL(BL117),.BLN(BLN117),.WL(WL114));
sram_cell_6t_5 inst_cell_114_118 (.BL(BL118),.BLN(BLN118),.WL(WL114));
sram_cell_6t_5 inst_cell_114_119 (.BL(BL119),.BLN(BLN119),.WL(WL114));
sram_cell_6t_5 inst_cell_114_120 (.BL(BL120),.BLN(BLN120),.WL(WL114));
sram_cell_6t_5 inst_cell_114_121 (.BL(BL121),.BLN(BLN121),.WL(WL114));
sram_cell_6t_5 inst_cell_114_122 (.BL(BL122),.BLN(BLN122),.WL(WL114));
sram_cell_6t_5 inst_cell_114_123 (.BL(BL123),.BLN(BLN123),.WL(WL114));
sram_cell_6t_5 inst_cell_114_124 (.BL(BL124),.BLN(BLN124),.WL(WL114));
sram_cell_6t_5 inst_cell_114_125 (.BL(BL125),.BLN(BLN125),.WL(WL114));
sram_cell_6t_5 inst_cell_114_126 (.BL(BL126),.BLN(BLN126),.WL(WL114));
sram_cell_6t_5 inst_cell_114_127 (.BL(BL127),.BLN(BLN127),.WL(WL114));
sram_cell_6t_5 inst_cell_115_0 (.BL(BL0),.BLN(BLN0),.WL(WL115));
sram_cell_6t_5 inst_cell_115_1 (.BL(BL1),.BLN(BLN1),.WL(WL115));
sram_cell_6t_5 inst_cell_115_2 (.BL(BL2),.BLN(BLN2),.WL(WL115));
sram_cell_6t_5 inst_cell_115_3 (.BL(BL3),.BLN(BLN3),.WL(WL115));
sram_cell_6t_5 inst_cell_115_4 (.BL(BL4),.BLN(BLN4),.WL(WL115));
sram_cell_6t_5 inst_cell_115_5 (.BL(BL5),.BLN(BLN5),.WL(WL115));
sram_cell_6t_5 inst_cell_115_6 (.BL(BL6),.BLN(BLN6),.WL(WL115));
sram_cell_6t_5 inst_cell_115_7 (.BL(BL7),.BLN(BLN7),.WL(WL115));
sram_cell_6t_5 inst_cell_115_8 (.BL(BL8),.BLN(BLN8),.WL(WL115));
sram_cell_6t_5 inst_cell_115_9 (.BL(BL9),.BLN(BLN9),.WL(WL115));
sram_cell_6t_5 inst_cell_115_10 (.BL(BL10),.BLN(BLN10),.WL(WL115));
sram_cell_6t_5 inst_cell_115_11 (.BL(BL11),.BLN(BLN11),.WL(WL115));
sram_cell_6t_5 inst_cell_115_12 (.BL(BL12),.BLN(BLN12),.WL(WL115));
sram_cell_6t_5 inst_cell_115_13 (.BL(BL13),.BLN(BLN13),.WL(WL115));
sram_cell_6t_5 inst_cell_115_14 (.BL(BL14),.BLN(BLN14),.WL(WL115));
sram_cell_6t_5 inst_cell_115_15 (.BL(BL15),.BLN(BLN15),.WL(WL115));
sram_cell_6t_5 inst_cell_115_16 (.BL(BL16),.BLN(BLN16),.WL(WL115));
sram_cell_6t_5 inst_cell_115_17 (.BL(BL17),.BLN(BLN17),.WL(WL115));
sram_cell_6t_5 inst_cell_115_18 (.BL(BL18),.BLN(BLN18),.WL(WL115));
sram_cell_6t_5 inst_cell_115_19 (.BL(BL19),.BLN(BLN19),.WL(WL115));
sram_cell_6t_5 inst_cell_115_20 (.BL(BL20),.BLN(BLN20),.WL(WL115));
sram_cell_6t_5 inst_cell_115_21 (.BL(BL21),.BLN(BLN21),.WL(WL115));
sram_cell_6t_5 inst_cell_115_22 (.BL(BL22),.BLN(BLN22),.WL(WL115));
sram_cell_6t_5 inst_cell_115_23 (.BL(BL23),.BLN(BLN23),.WL(WL115));
sram_cell_6t_5 inst_cell_115_24 (.BL(BL24),.BLN(BLN24),.WL(WL115));
sram_cell_6t_5 inst_cell_115_25 (.BL(BL25),.BLN(BLN25),.WL(WL115));
sram_cell_6t_5 inst_cell_115_26 (.BL(BL26),.BLN(BLN26),.WL(WL115));
sram_cell_6t_5 inst_cell_115_27 (.BL(BL27),.BLN(BLN27),.WL(WL115));
sram_cell_6t_5 inst_cell_115_28 (.BL(BL28),.BLN(BLN28),.WL(WL115));
sram_cell_6t_5 inst_cell_115_29 (.BL(BL29),.BLN(BLN29),.WL(WL115));
sram_cell_6t_5 inst_cell_115_30 (.BL(BL30),.BLN(BLN30),.WL(WL115));
sram_cell_6t_5 inst_cell_115_31 (.BL(BL31),.BLN(BLN31),.WL(WL115));
sram_cell_6t_5 inst_cell_115_32 (.BL(BL32),.BLN(BLN32),.WL(WL115));
sram_cell_6t_5 inst_cell_115_33 (.BL(BL33),.BLN(BLN33),.WL(WL115));
sram_cell_6t_5 inst_cell_115_34 (.BL(BL34),.BLN(BLN34),.WL(WL115));
sram_cell_6t_5 inst_cell_115_35 (.BL(BL35),.BLN(BLN35),.WL(WL115));
sram_cell_6t_5 inst_cell_115_36 (.BL(BL36),.BLN(BLN36),.WL(WL115));
sram_cell_6t_5 inst_cell_115_37 (.BL(BL37),.BLN(BLN37),.WL(WL115));
sram_cell_6t_5 inst_cell_115_38 (.BL(BL38),.BLN(BLN38),.WL(WL115));
sram_cell_6t_5 inst_cell_115_39 (.BL(BL39),.BLN(BLN39),.WL(WL115));
sram_cell_6t_5 inst_cell_115_40 (.BL(BL40),.BLN(BLN40),.WL(WL115));
sram_cell_6t_5 inst_cell_115_41 (.BL(BL41),.BLN(BLN41),.WL(WL115));
sram_cell_6t_5 inst_cell_115_42 (.BL(BL42),.BLN(BLN42),.WL(WL115));
sram_cell_6t_5 inst_cell_115_43 (.BL(BL43),.BLN(BLN43),.WL(WL115));
sram_cell_6t_5 inst_cell_115_44 (.BL(BL44),.BLN(BLN44),.WL(WL115));
sram_cell_6t_5 inst_cell_115_45 (.BL(BL45),.BLN(BLN45),.WL(WL115));
sram_cell_6t_5 inst_cell_115_46 (.BL(BL46),.BLN(BLN46),.WL(WL115));
sram_cell_6t_5 inst_cell_115_47 (.BL(BL47),.BLN(BLN47),.WL(WL115));
sram_cell_6t_5 inst_cell_115_48 (.BL(BL48),.BLN(BLN48),.WL(WL115));
sram_cell_6t_5 inst_cell_115_49 (.BL(BL49),.BLN(BLN49),.WL(WL115));
sram_cell_6t_5 inst_cell_115_50 (.BL(BL50),.BLN(BLN50),.WL(WL115));
sram_cell_6t_5 inst_cell_115_51 (.BL(BL51),.BLN(BLN51),.WL(WL115));
sram_cell_6t_5 inst_cell_115_52 (.BL(BL52),.BLN(BLN52),.WL(WL115));
sram_cell_6t_5 inst_cell_115_53 (.BL(BL53),.BLN(BLN53),.WL(WL115));
sram_cell_6t_5 inst_cell_115_54 (.BL(BL54),.BLN(BLN54),.WL(WL115));
sram_cell_6t_5 inst_cell_115_55 (.BL(BL55),.BLN(BLN55),.WL(WL115));
sram_cell_6t_5 inst_cell_115_56 (.BL(BL56),.BLN(BLN56),.WL(WL115));
sram_cell_6t_5 inst_cell_115_57 (.BL(BL57),.BLN(BLN57),.WL(WL115));
sram_cell_6t_5 inst_cell_115_58 (.BL(BL58),.BLN(BLN58),.WL(WL115));
sram_cell_6t_5 inst_cell_115_59 (.BL(BL59),.BLN(BLN59),.WL(WL115));
sram_cell_6t_5 inst_cell_115_60 (.BL(BL60),.BLN(BLN60),.WL(WL115));
sram_cell_6t_5 inst_cell_115_61 (.BL(BL61),.BLN(BLN61),.WL(WL115));
sram_cell_6t_5 inst_cell_115_62 (.BL(BL62),.BLN(BLN62),.WL(WL115));
sram_cell_6t_5 inst_cell_115_63 (.BL(BL63),.BLN(BLN63),.WL(WL115));
sram_cell_6t_5 inst_cell_115_64 (.BL(BL64),.BLN(BLN64),.WL(WL115));
sram_cell_6t_5 inst_cell_115_65 (.BL(BL65),.BLN(BLN65),.WL(WL115));
sram_cell_6t_5 inst_cell_115_66 (.BL(BL66),.BLN(BLN66),.WL(WL115));
sram_cell_6t_5 inst_cell_115_67 (.BL(BL67),.BLN(BLN67),.WL(WL115));
sram_cell_6t_5 inst_cell_115_68 (.BL(BL68),.BLN(BLN68),.WL(WL115));
sram_cell_6t_5 inst_cell_115_69 (.BL(BL69),.BLN(BLN69),.WL(WL115));
sram_cell_6t_5 inst_cell_115_70 (.BL(BL70),.BLN(BLN70),.WL(WL115));
sram_cell_6t_5 inst_cell_115_71 (.BL(BL71),.BLN(BLN71),.WL(WL115));
sram_cell_6t_5 inst_cell_115_72 (.BL(BL72),.BLN(BLN72),.WL(WL115));
sram_cell_6t_5 inst_cell_115_73 (.BL(BL73),.BLN(BLN73),.WL(WL115));
sram_cell_6t_5 inst_cell_115_74 (.BL(BL74),.BLN(BLN74),.WL(WL115));
sram_cell_6t_5 inst_cell_115_75 (.BL(BL75),.BLN(BLN75),.WL(WL115));
sram_cell_6t_5 inst_cell_115_76 (.BL(BL76),.BLN(BLN76),.WL(WL115));
sram_cell_6t_5 inst_cell_115_77 (.BL(BL77),.BLN(BLN77),.WL(WL115));
sram_cell_6t_5 inst_cell_115_78 (.BL(BL78),.BLN(BLN78),.WL(WL115));
sram_cell_6t_5 inst_cell_115_79 (.BL(BL79),.BLN(BLN79),.WL(WL115));
sram_cell_6t_5 inst_cell_115_80 (.BL(BL80),.BLN(BLN80),.WL(WL115));
sram_cell_6t_5 inst_cell_115_81 (.BL(BL81),.BLN(BLN81),.WL(WL115));
sram_cell_6t_5 inst_cell_115_82 (.BL(BL82),.BLN(BLN82),.WL(WL115));
sram_cell_6t_5 inst_cell_115_83 (.BL(BL83),.BLN(BLN83),.WL(WL115));
sram_cell_6t_5 inst_cell_115_84 (.BL(BL84),.BLN(BLN84),.WL(WL115));
sram_cell_6t_5 inst_cell_115_85 (.BL(BL85),.BLN(BLN85),.WL(WL115));
sram_cell_6t_5 inst_cell_115_86 (.BL(BL86),.BLN(BLN86),.WL(WL115));
sram_cell_6t_5 inst_cell_115_87 (.BL(BL87),.BLN(BLN87),.WL(WL115));
sram_cell_6t_5 inst_cell_115_88 (.BL(BL88),.BLN(BLN88),.WL(WL115));
sram_cell_6t_5 inst_cell_115_89 (.BL(BL89),.BLN(BLN89),.WL(WL115));
sram_cell_6t_5 inst_cell_115_90 (.BL(BL90),.BLN(BLN90),.WL(WL115));
sram_cell_6t_5 inst_cell_115_91 (.BL(BL91),.BLN(BLN91),.WL(WL115));
sram_cell_6t_5 inst_cell_115_92 (.BL(BL92),.BLN(BLN92),.WL(WL115));
sram_cell_6t_5 inst_cell_115_93 (.BL(BL93),.BLN(BLN93),.WL(WL115));
sram_cell_6t_5 inst_cell_115_94 (.BL(BL94),.BLN(BLN94),.WL(WL115));
sram_cell_6t_5 inst_cell_115_95 (.BL(BL95),.BLN(BLN95),.WL(WL115));
sram_cell_6t_5 inst_cell_115_96 (.BL(BL96),.BLN(BLN96),.WL(WL115));
sram_cell_6t_5 inst_cell_115_97 (.BL(BL97),.BLN(BLN97),.WL(WL115));
sram_cell_6t_5 inst_cell_115_98 (.BL(BL98),.BLN(BLN98),.WL(WL115));
sram_cell_6t_5 inst_cell_115_99 (.BL(BL99),.BLN(BLN99),.WL(WL115));
sram_cell_6t_5 inst_cell_115_100 (.BL(BL100),.BLN(BLN100),.WL(WL115));
sram_cell_6t_5 inst_cell_115_101 (.BL(BL101),.BLN(BLN101),.WL(WL115));
sram_cell_6t_5 inst_cell_115_102 (.BL(BL102),.BLN(BLN102),.WL(WL115));
sram_cell_6t_5 inst_cell_115_103 (.BL(BL103),.BLN(BLN103),.WL(WL115));
sram_cell_6t_5 inst_cell_115_104 (.BL(BL104),.BLN(BLN104),.WL(WL115));
sram_cell_6t_5 inst_cell_115_105 (.BL(BL105),.BLN(BLN105),.WL(WL115));
sram_cell_6t_5 inst_cell_115_106 (.BL(BL106),.BLN(BLN106),.WL(WL115));
sram_cell_6t_5 inst_cell_115_107 (.BL(BL107),.BLN(BLN107),.WL(WL115));
sram_cell_6t_5 inst_cell_115_108 (.BL(BL108),.BLN(BLN108),.WL(WL115));
sram_cell_6t_5 inst_cell_115_109 (.BL(BL109),.BLN(BLN109),.WL(WL115));
sram_cell_6t_5 inst_cell_115_110 (.BL(BL110),.BLN(BLN110),.WL(WL115));
sram_cell_6t_5 inst_cell_115_111 (.BL(BL111),.BLN(BLN111),.WL(WL115));
sram_cell_6t_5 inst_cell_115_112 (.BL(BL112),.BLN(BLN112),.WL(WL115));
sram_cell_6t_5 inst_cell_115_113 (.BL(BL113),.BLN(BLN113),.WL(WL115));
sram_cell_6t_5 inst_cell_115_114 (.BL(BL114),.BLN(BLN114),.WL(WL115));
sram_cell_6t_5 inst_cell_115_115 (.BL(BL115),.BLN(BLN115),.WL(WL115));
sram_cell_6t_5 inst_cell_115_116 (.BL(BL116),.BLN(BLN116),.WL(WL115));
sram_cell_6t_5 inst_cell_115_117 (.BL(BL117),.BLN(BLN117),.WL(WL115));
sram_cell_6t_5 inst_cell_115_118 (.BL(BL118),.BLN(BLN118),.WL(WL115));
sram_cell_6t_5 inst_cell_115_119 (.BL(BL119),.BLN(BLN119),.WL(WL115));
sram_cell_6t_5 inst_cell_115_120 (.BL(BL120),.BLN(BLN120),.WL(WL115));
sram_cell_6t_5 inst_cell_115_121 (.BL(BL121),.BLN(BLN121),.WL(WL115));
sram_cell_6t_5 inst_cell_115_122 (.BL(BL122),.BLN(BLN122),.WL(WL115));
sram_cell_6t_5 inst_cell_115_123 (.BL(BL123),.BLN(BLN123),.WL(WL115));
sram_cell_6t_5 inst_cell_115_124 (.BL(BL124),.BLN(BLN124),.WL(WL115));
sram_cell_6t_5 inst_cell_115_125 (.BL(BL125),.BLN(BLN125),.WL(WL115));
sram_cell_6t_5 inst_cell_115_126 (.BL(BL126),.BLN(BLN126),.WL(WL115));
sram_cell_6t_5 inst_cell_115_127 (.BL(BL127),.BLN(BLN127),.WL(WL115));
sram_cell_6t_5 inst_cell_116_0 (.BL(BL0),.BLN(BLN0),.WL(WL116));
sram_cell_6t_5 inst_cell_116_1 (.BL(BL1),.BLN(BLN1),.WL(WL116));
sram_cell_6t_5 inst_cell_116_2 (.BL(BL2),.BLN(BLN2),.WL(WL116));
sram_cell_6t_5 inst_cell_116_3 (.BL(BL3),.BLN(BLN3),.WL(WL116));
sram_cell_6t_5 inst_cell_116_4 (.BL(BL4),.BLN(BLN4),.WL(WL116));
sram_cell_6t_5 inst_cell_116_5 (.BL(BL5),.BLN(BLN5),.WL(WL116));
sram_cell_6t_5 inst_cell_116_6 (.BL(BL6),.BLN(BLN6),.WL(WL116));
sram_cell_6t_5 inst_cell_116_7 (.BL(BL7),.BLN(BLN7),.WL(WL116));
sram_cell_6t_5 inst_cell_116_8 (.BL(BL8),.BLN(BLN8),.WL(WL116));
sram_cell_6t_5 inst_cell_116_9 (.BL(BL9),.BLN(BLN9),.WL(WL116));
sram_cell_6t_5 inst_cell_116_10 (.BL(BL10),.BLN(BLN10),.WL(WL116));
sram_cell_6t_5 inst_cell_116_11 (.BL(BL11),.BLN(BLN11),.WL(WL116));
sram_cell_6t_5 inst_cell_116_12 (.BL(BL12),.BLN(BLN12),.WL(WL116));
sram_cell_6t_5 inst_cell_116_13 (.BL(BL13),.BLN(BLN13),.WL(WL116));
sram_cell_6t_5 inst_cell_116_14 (.BL(BL14),.BLN(BLN14),.WL(WL116));
sram_cell_6t_5 inst_cell_116_15 (.BL(BL15),.BLN(BLN15),.WL(WL116));
sram_cell_6t_5 inst_cell_116_16 (.BL(BL16),.BLN(BLN16),.WL(WL116));
sram_cell_6t_5 inst_cell_116_17 (.BL(BL17),.BLN(BLN17),.WL(WL116));
sram_cell_6t_5 inst_cell_116_18 (.BL(BL18),.BLN(BLN18),.WL(WL116));
sram_cell_6t_5 inst_cell_116_19 (.BL(BL19),.BLN(BLN19),.WL(WL116));
sram_cell_6t_5 inst_cell_116_20 (.BL(BL20),.BLN(BLN20),.WL(WL116));
sram_cell_6t_5 inst_cell_116_21 (.BL(BL21),.BLN(BLN21),.WL(WL116));
sram_cell_6t_5 inst_cell_116_22 (.BL(BL22),.BLN(BLN22),.WL(WL116));
sram_cell_6t_5 inst_cell_116_23 (.BL(BL23),.BLN(BLN23),.WL(WL116));
sram_cell_6t_5 inst_cell_116_24 (.BL(BL24),.BLN(BLN24),.WL(WL116));
sram_cell_6t_5 inst_cell_116_25 (.BL(BL25),.BLN(BLN25),.WL(WL116));
sram_cell_6t_5 inst_cell_116_26 (.BL(BL26),.BLN(BLN26),.WL(WL116));
sram_cell_6t_5 inst_cell_116_27 (.BL(BL27),.BLN(BLN27),.WL(WL116));
sram_cell_6t_5 inst_cell_116_28 (.BL(BL28),.BLN(BLN28),.WL(WL116));
sram_cell_6t_5 inst_cell_116_29 (.BL(BL29),.BLN(BLN29),.WL(WL116));
sram_cell_6t_5 inst_cell_116_30 (.BL(BL30),.BLN(BLN30),.WL(WL116));
sram_cell_6t_5 inst_cell_116_31 (.BL(BL31),.BLN(BLN31),.WL(WL116));
sram_cell_6t_5 inst_cell_116_32 (.BL(BL32),.BLN(BLN32),.WL(WL116));
sram_cell_6t_5 inst_cell_116_33 (.BL(BL33),.BLN(BLN33),.WL(WL116));
sram_cell_6t_5 inst_cell_116_34 (.BL(BL34),.BLN(BLN34),.WL(WL116));
sram_cell_6t_5 inst_cell_116_35 (.BL(BL35),.BLN(BLN35),.WL(WL116));
sram_cell_6t_5 inst_cell_116_36 (.BL(BL36),.BLN(BLN36),.WL(WL116));
sram_cell_6t_5 inst_cell_116_37 (.BL(BL37),.BLN(BLN37),.WL(WL116));
sram_cell_6t_5 inst_cell_116_38 (.BL(BL38),.BLN(BLN38),.WL(WL116));
sram_cell_6t_5 inst_cell_116_39 (.BL(BL39),.BLN(BLN39),.WL(WL116));
sram_cell_6t_5 inst_cell_116_40 (.BL(BL40),.BLN(BLN40),.WL(WL116));
sram_cell_6t_5 inst_cell_116_41 (.BL(BL41),.BLN(BLN41),.WL(WL116));
sram_cell_6t_5 inst_cell_116_42 (.BL(BL42),.BLN(BLN42),.WL(WL116));
sram_cell_6t_5 inst_cell_116_43 (.BL(BL43),.BLN(BLN43),.WL(WL116));
sram_cell_6t_5 inst_cell_116_44 (.BL(BL44),.BLN(BLN44),.WL(WL116));
sram_cell_6t_5 inst_cell_116_45 (.BL(BL45),.BLN(BLN45),.WL(WL116));
sram_cell_6t_5 inst_cell_116_46 (.BL(BL46),.BLN(BLN46),.WL(WL116));
sram_cell_6t_5 inst_cell_116_47 (.BL(BL47),.BLN(BLN47),.WL(WL116));
sram_cell_6t_5 inst_cell_116_48 (.BL(BL48),.BLN(BLN48),.WL(WL116));
sram_cell_6t_5 inst_cell_116_49 (.BL(BL49),.BLN(BLN49),.WL(WL116));
sram_cell_6t_5 inst_cell_116_50 (.BL(BL50),.BLN(BLN50),.WL(WL116));
sram_cell_6t_5 inst_cell_116_51 (.BL(BL51),.BLN(BLN51),.WL(WL116));
sram_cell_6t_5 inst_cell_116_52 (.BL(BL52),.BLN(BLN52),.WL(WL116));
sram_cell_6t_5 inst_cell_116_53 (.BL(BL53),.BLN(BLN53),.WL(WL116));
sram_cell_6t_5 inst_cell_116_54 (.BL(BL54),.BLN(BLN54),.WL(WL116));
sram_cell_6t_5 inst_cell_116_55 (.BL(BL55),.BLN(BLN55),.WL(WL116));
sram_cell_6t_5 inst_cell_116_56 (.BL(BL56),.BLN(BLN56),.WL(WL116));
sram_cell_6t_5 inst_cell_116_57 (.BL(BL57),.BLN(BLN57),.WL(WL116));
sram_cell_6t_5 inst_cell_116_58 (.BL(BL58),.BLN(BLN58),.WL(WL116));
sram_cell_6t_5 inst_cell_116_59 (.BL(BL59),.BLN(BLN59),.WL(WL116));
sram_cell_6t_5 inst_cell_116_60 (.BL(BL60),.BLN(BLN60),.WL(WL116));
sram_cell_6t_5 inst_cell_116_61 (.BL(BL61),.BLN(BLN61),.WL(WL116));
sram_cell_6t_5 inst_cell_116_62 (.BL(BL62),.BLN(BLN62),.WL(WL116));
sram_cell_6t_5 inst_cell_116_63 (.BL(BL63),.BLN(BLN63),.WL(WL116));
sram_cell_6t_5 inst_cell_116_64 (.BL(BL64),.BLN(BLN64),.WL(WL116));
sram_cell_6t_5 inst_cell_116_65 (.BL(BL65),.BLN(BLN65),.WL(WL116));
sram_cell_6t_5 inst_cell_116_66 (.BL(BL66),.BLN(BLN66),.WL(WL116));
sram_cell_6t_5 inst_cell_116_67 (.BL(BL67),.BLN(BLN67),.WL(WL116));
sram_cell_6t_5 inst_cell_116_68 (.BL(BL68),.BLN(BLN68),.WL(WL116));
sram_cell_6t_5 inst_cell_116_69 (.BL(BL69),.BLN(BLN69),.WL(WL116));
sram_cell_6t_5 inst_cell_116_70 (.BL(BL70),.BLN(BLN70),.WL(WL116));
sram_cell_6t_5 inst_cell_116_71 (.BL(BL71),.BLN(BLN71),.WL(WL116));
sram_cell_6t_5 inst_cell_116_72 (.BL(BL72),.BLN(BLN72),.WL(WL116));
sram_cell_6t_5 inst_cell_116_73 (.BL(BL73),.BLN(BLN73),.WL(WL116));
sram_cell_6t_5 inst_cell_116_74 (.BL(BL74),.BLN(BLN74),.WL(WL116));
sram_cell_6t_5 inst_cell_116_75 (.BL(BL75),.BLN(BLN75),.WL(WL116));
sram_cell_6t_5 inst_cell_116_76 (.BL(BL76),.BLN(BLN76),.WL(WL116));
sram_cell_6t_5 inst_cell_116_77 (.BL(BL77),.BLN(BLN77),.WL(WL116));
sram_cell_6t_5 inst_cell_116_78 (.BL(BL78),.BLN(BLN78),.WL(WL116));
sram_cell_6t_5 inst_cell_116_79 (.BL(BL79),.BLN(BLN79),.WL(WL116));
sram_cell_6t_5 inst_cell_116_80 (.BL(BL80),.BLN(BLN80),.WL(WL116));
sram_cell_6t_5 inst_cell_116_81 (.BL(BL81),.BLN(BLN81),.WL(WL116));
sram_cell_6t_5 inst_cell_116_82 (.BL(BL82),.BLN(BLN82),.WL(WL116));
sram_cell_6t_5 inst_cell_116_83 (.BL(BL83),.BLN(BLN83),.WL(WL116));
sram_cell_6t_5 inst_cell_116_84 (.BL(BL84),.BLN(BLN84),.WL(WL116));
sram_cell_6t_5 inst_cell_116_85 (.BL(BL85),.BLN(BLN85),.WL(WL116));
sram_cell_6t_5 inst_cell_116_86 (.BL(BL86),.BLN(BLN86),.WL(WL116));
sram_cell_6t_5 inst_cell_116_87 (.BL(BL87),.BLN(BLN87),.WL(WL116));
sram_cell_6t_5 inst_cell_116_88 (.BL(BL88),.BLN(BLN88),.WL(WL116));
sram_cell_6t_5 inst_cell_116_89 (.BL(BL89),.BLN(BLN89),.WL(WL116));
sram_cell_6t_5 inst_cell_116_90 (.BL(BL90),.BLN(BLN90),.WL(WL116));
sram_cell_6t_5 inst_cell_116_91 (.BL(BL91),.BLN(BLN91),.WL(WL116));
sram_cell_6t_5 inst_cell_116_92 (.BL(BL92),.BLN(BLN92),.WL(WL116));
sram_cell_6t_5 inst_cell_116_93 (.BL(BL93),.BLN(BLN93),.WL(WL116));
sram_cell_6t_5 inst_cell_116_94 (.BL(BL94),.BLN(BLN94),.WL(WL116));
sram_cell_6t_5 inst_cell_116_95 (.BL(BL95),.BLN(BLN95),.WL(WL116));
sram_cell_6t_5 inst_cell_116_96 (.BL(BL96),.BLN(BLN96),.WL(WL116));
sram_cell_6t_5 inst_cell_116_97 (.BL(BL97),.BLN(BLN97),.WL(WL116));
sram_cell_6t_5 inst_cell_116_98 (.BL(BL98),.BLN(BLN98),.WL(WL116));
sram_cell_6t_5 inst_cell_116_99 (.BL(BL99),.BLN(BLN99),.WL(WL116));
sram_cell_6t_5 inst_cell_116_100 (.BL(BL100),.BLN(BLN100),.WL(WL116));
sram_cell_6t_5 inst_cell_116_101 (.BL(BL101),.BLN(BLN101),.WL(WL116));
sram_cell_6t_5 inst_cell_116_102 (.BL(BL102),.BLN(BLN102),.WL(WL116));
sram_cell_6t_5 inst_cell_116_103 (.BL(BL103),.BLN(BLN103),.WL(WL116));
sram_cell_6t_5 inst_cell_116_104 (.BL(BL104),.BLN(BLN104),.WL(WL116));
sram_cell_6t_5 inst_cell_116_105 (.BL(BL105),.BLN(BLN105),.WL(WL116));
sram_cell_6t_5 inst_cell_116_106 (.BL(BL106),.BLN(BLN106),.WL(WL116));
sram_cell_6t_5 inst_cell_116_107 (.BL(BL107),.BLN(BLN107),.WL(WL116));
sram_cell_6t_5 inst_cell_116_108 (.BL(BL108),.BLN(BLN108),.WL(WL116));
sram_cell_6t_5 inst_cell_116_109 (.BL(BL109),.BLN(BLN109),.WL(WL116));
sram_cell_6t_5 inst_cell_116_110 (.BL(BL110),.BLN(BLN110),.WL(WL116));
sram_cell_6t_5 inst_cell_116_111 (.BL(BL111),.BLN(BLN111),.WL(WL116));
sram_cell_6t_5 inst_cell_116_112 (.BL(BL112),.BLN(BLN112),.WL(WL116));
sram_cell_6t_5 inst_cell_116_113 (.BL(BL113),.BLN(BLN113),.WL(WL116));
sram_cell_6t_5 inst_cell_116_114 (.BL(BL114),.BLN(BLN114),.WL(WL116));
sram_cell_6t_5 inst_cell_116_115 (.BL(BL115),.BLN(BLN115),.WL(WL116));
sram_cell_6t_5 inst_cell_116_116 (.BL(BL116),.BLN(BLN116),.WL(WL116));
sram_cell_6t_5 inst_cell_116_117 (.BL(BL117),.BLN(BLN117),.WL(WL116));
sram_cell_6t_5 inst_cell_116_118 (.BL(BL118),.BLN(BLN118),.WL(WL116));
sram_cell_6t_5 inst_cell_116_119 (.BL(BL119),.BLN(BLN119),.WL(WL116));
sram_cell_6t_5 inst_cell_116_120 (.BL(BL120),.BLN(BLN120),.WL(WL116));
sram_cell_6t_5 inst_cell_116_121 (.BL(BL121),.BLN(BLN121),.WL(WL116));
sram_cell_6t_5 inst_cell_116_122 (.BL(BL122),.BLN(BLN122),.WL(WL116));
sram_cell_6t_5 inst_cell_116_123 (.BL(BL123),.BLN(BLN123),.WL(WL116));
sram_cell_6t_5 inst_cell_116_124 (.BL(BL124),.BLN(BLN124),.WL(WL116));
sram_cell_6t_5 inst_cell_116_125 (.BL(BL125),.BLN(BLN125),.WL(WL116));
sram_cell_6t_5 inst_cell_116_126 (.BL(BL126),.BLN(BLN126),.WL(WL116));
sram_cell_6t_5 inst_cell_116_127 (.BL(BL127),.BLN(BLN127),.WL(WL116));
sram_cell_6t_5 inst_cell_117_0 (.BL(BL0),.BLN(BLN0),.WL(WL117));
sram_cell_6t_5 inst_cell_117_1 (.BL(BL1),.BLN(BLN1),.WL(WL117));
sram_cell_6t_5 inst_cell_117_2 (.BL(BL2),.BLN(BLN2),.WL(WL117));
sram_cell_6t_5 inst_cell_117_3 (.BL(BL3),.BLN(BLN3),.WL(WL117));
sram_cell_6t_5 inst_cell_117_4 (.BL(BL4),.BLN(BLN4),.WL(WL117));
sram_cell_6t_5 inst_cell_117_5 (.BL(BL5),.BLN(BLN5),.WL(WL117));
sram_cell_6t_5 inst_cell_117_6 (.BL(BL6),.BLN(BLN6),.WL(WL117));
sram_cell_6t_5 inst_cell_117_7 (.BL(BL7),.BLN(BLN7),.WL(WL117));
sram_cell_6t_5 inst_cell_117_8 (.BL(BL8),.BLN(BLN8),.WL(WL117));
sram_cell_6t_5 inst_cell_117_9 (.BL(BL9),.BLN(BLN9),.WL(WL117));
sram_cell_6t_5 inst_cell_117_10 (.BL(BL10),.BLN(BLN10),.WL(WL117));
sram_cell_6t_5 inst_cell_117_11 (.BL(BL11),.BLN(BLN11),.WL(WL117));
sram_cell_6t_5 inst_cell_117_12 (.BL(BL12),.BLN(BLN12),.WL(WL117));
sram_cell_6t_5 inst_cell_117_13 (.BL(BL13),.BLN(BLN13),.WL(WL117));
sram_cell_6t_5 inst_cell_117_14 (.BL(BL14),.BLN(BLN14),.WL(WL117));
sram_cell_6t_5 inst_cell_117_15 (.BL(BL15),.BLN(BLN15),.WL(WL117));
sram_cell_6t_5 inst_cell_117_16 (.BL(BL16),.BLN(BLN16),.WL(WL117));
sram_cell_6t_5 inst_cell_117_17 (.BL(BL17),.BLN(BLN17),.WL(WL117));
sram_cell_6t_5 inst_cell_117_18 (.BL(BL18),.BLN(BLN18),.WL(WL117));
sram_cell_6t_5 inst_cell_117_19 (.BL(BL19),.BLN(BLN19),.WL(WL117));
sram_cell_6t_5 inst_cell_117_20 (.BL(BL20),.BLN(BLN20),.WL(WL117));
sram_cell_6t_5 inst_cell_117_21 (.BL(BL21),.BLN(BLN21),.WL(WL117));
sram_cell_6t_5 inst_cell_117_22 (.BL(BL22),.BLN(BLN22),.WL(WL117));
sram_cell_6t_5 inst_cell_117_23 (.BL(BL23),.BLN(BLN23),.WL(WL117));
sram_cell_6t_5 inst_cell_117_24 (.BL(BL24),.BLN(BLN24),.WL(WL117));
sram_cell_6t_5 inst_cell_117_25 (.BL(BL25),.BLN(BLN25),.WL(WL117));
sram_cell_6t_5 inst_cell_117_26 (.BL(BL26),.BLN(BLN26),.WL(WL117));
sram_cell_6t_5 inst_cell_117_27 (.BL(BL27),.BLN(BLN27),.WL(WL117));
sram_cell_6t_5 inst_cell_117_28 (.BL(BL28),.BLN(BLN28),.WL(WL117));
sram_cell_6t_5 inst_cell_117_29 (.BL(BL29),.BLN(BLN29),.WL(WL117));
sram_cell_6t_5 inst_cell_117_30 (.BL(BL30),.BLN(BLN30),.WL(WL117));
sram_cell_6t_5 inst_cell_117_31 (.BL(BL31),.BLN(BLN31),.WL(WL117));
sram_cell_6t_5 inst_cell_117_32 (.BL(BL32),.BLN(BLN32),.WL(WL117));
sram_cell_6t_5 inst_cell_117_33 (.BL(BL33),.BLN(BLN33),.WL(WL117));
sram_cell_6t_5 inst_cell_117_34 (.BL(BL34),.BLN(BLN34),.WL(WL117));
sram_cell_6t_5 inst_cell_117_35 (.BL(BL35),.BLN(BLN35),.WL(WL117));
sram_cell_6t_5 inst_cell_117_36 (.BL(BL36),.BLN(BLN36),.WL(WL117));
sram_cell_6t_5 inst_cell_117_37 (.BL(BL37),.BLN(BLN37),.WL(WL117));
sram_cell_6t_5 inst_cell_117_38 (.BL(BL38),.BLN(BLN38),.WL(WL117));
sram_cell_6t_5 inst_cell_117_39 (.BL(BL39),.BLN(BLN39),.WL(WL117));
sram_cell_6t_5 inst_cell_117_40 (.BL(BL40),.BLN(BLN40),.WL(WL117));
sram_cell_6t_5 inst_cell_117_41 (.BL(BL41),.BLN(BLN41),.WL(WL117));
sram_cell_6t_5 inst_cell_117_42 (.BL(BL42),.BLN(BLN42),.WL(WL117));
sram_cell_6t_5 inst_cell_117_43 (.BL(BL43),.BLN(BLN43),.WL(WL117));
sram_cell_6t_5 inst_cell_117_44 (.BL(BL44),.BLN(BLN44),.WL(WL117));
sram_cell_6t_5 inst_cell_117_45 (.BL(BL45),.BLN(BLN45),.WL(WL117));
sram_cell_6t_5 inst_cell_117_46 (.BL(BL46),.BLN(BLN46),.WL(WL117));
sram_cell_6t_5 inst_cell_117_47 (.BL(BL47),.BLN(BLN47),.WL(WL117));
sram_cell_6t_5 inst_cell_117_48 (.BL(BL48),.BLN(BLN48),.WL(WL117));
sram_cell_6t_5 inst_cell_117_49 (.BL(BL49),.BLN(BLN49),.WL(WL117));
sram_cell_6t_5 inst_cell_117_50 (.BL(BL50),.BLN(BLN50),.WL(WL117));
sram_cell_6t_5 inst_cell_117_51 (.BL(BL51),.BLN(BLN51),.WL(WL117));
sram_cell_6t_5 inst_cell_117_52 (.BL(BL52),.BLN(BLN52),.WL(WL117));
sram_cell_6t_5 inst_cell_117_53 (.BL(BL53),.BLN(BLN53),.WL(WL117));
sram_cell_6t_5 inst_cell_117_54 (.BL(BL54),.BLN(BLN54),.WL(WL117));
sram_cell_6t_5 inst_cell_117_55 (.BL(BL55),.BLN(BLN55),.WL(WL117));
sram_cell_6t_5 inst_cell_117_56 (.BL(BL56),.BLN(BLN56),.WL(WL117));
sram_cell_6t_5 inst_cell_117_57 (.BL(BL57),.BLN(BLN57),.WL(WL117));
sram_cell_6t_5 inst_cell_117_58 (.BL(BL58),.BLN(BLN58),.WL(WL117));
sram_cell_6t_5 inst_cell_117_59 (.BL(BL59),.BLN(BLN59),.WL(WL117));
sram_cell_6t_5 inst_cell_117_60 (.BL(BL60),.BLN(BLN60),.WL(WL117));
sram_cell_6t_5 inst_cell_117_61 (.BL(BL61),.BLN(BLN61),.WL(WL117));
sram_cell_6t_5 inst_cell_117_62 (.BL(BL62),.BLN(BLN62),.WL(WL117));
sram_cell_6t_5 inst_cell_117_63 (.BL(BL63),.BLN(BLN63),.WL(WL117));
sram_cell_6t_5 inst_cell_117_64 (.BL(BL64),.BLN(BLN64),.WL(WL117));
sram_cell_6t_5 inst_cell_117_65 (.BL(BL65),.BLN(BLN65),.WL(WL117));
sram_cell_6t_5 inst_cell_117_66 (.BL(BL66),.BLN(BLN66),.WL(WL117));
sram_cell_6t_5 inst_cell_117_67 (.BL(BL67),.BLN(BLN67),.WL(WL117));
sram_cell_6t_5 inst_cell_117_68 (.BL(BL68),.BLN(BLN68),.WL(WL117));
sram_cell_6t_5 inst_cell_117_69 (.BL(BL69),.BLN(BLN69),.WL(WL117));
sram_cell_6t_5 inst_cell_117_70 (.BL(BL70),.BLN(BLN70),.WL(WL117));
sram_cell_6t_5 inst_cell_117_71 (.BL(BL71),.BLN(BLN71),.WL(WL117));
sram_cell_6t_5 inst_cell_117_72 (.BL(BL72),.BLN(BLN72),.WL(WL117));
sram_cell_6t_5 inst_cell_117_73 (.BL(BL73),.BLN(BLN73),.WL(WL117));
sram_cell_6t_5 inst_cell_117_74 (.BL(BL74),.BLN(BLN74),.WL(WL117));
sram_cell_6t_5 inst_cell_117_75 (.BL(BL75),.BLN(BLN75),.WL(WL117));
sram_cell_6t_5 inst_cell_117_76 (.BL(BL76),.BLN(BLN76),.WL(WL117));
sram_cell_6t_5 inst_cell_117_77 (.BL(BL77),.BLN(BLN77),.WL(WL117));
sram_cell_6t_5 inst_cell_117_78 (.BL(BL78),.BLN(BLN78),.WL(WL117));
sram_cell_6t_5 inst_cell_117_79 (.BL(BL79),.BLN(BLN79),.WL(WL117));
sram_cell_6t_5 inst_cell_117_80 (.BL(BL80),.BLN(BLN80),.WL(WL117));
sram_cell_6t_5 inst_cell_117_81 (.BL(BL81),.BLN(BLN81),.WL(WL117));
sram_cell_6t_5 inst_cell_117_82 (.BL(BL82),.BLN(BLN82),.WL(WL117));
sram_cell_6t_5 inst_cell_117_83 (.BL(BL83),.BLN(BLN83),.WL(WL117));
sram_cell_6t_5 inst_cell_117_84 (.BL(BL84),.BLN(BLN84),.WL(WL117));
sram_cell_6t_5 inst_cell_117_85 (.BL(BL85),.BLN(BLN85),.WL(WL117));
sram_cell_6t_5 inst_cell_117_86 (.BL(BL86),.BLN(BLN86),.WL(WL117));
sram_cell_6t_5 inst_cell_117_87 (.BL(BL87),.BLN(BLN87),.WL(WL117));
sram_cell_6t_5 inst_cell_117_88 (.BL(BL88),.BLN(BLN88),.WL(WL117));
sram_cell_6t_5 inst_cell_117_89 (.BL(BL89),.BLN(BLN89),.WL(WL117));
sram_cell_6t_5 inst_cell_117_90 (.BL(BL90),.BLN(BLN90),.WL(WL117));
sram_cell_6t_5 inst_cell_117_91 (.BL(BL91),.BLN(BLN91),.WL(WL117));
sram_cell_6t_5 inst_cell_117_92 (.BL(BL92),.BLN(BLN92),.WL(WL117));
sram_cell_6t_5 inst_cell_117_93 (.BL(BL93),.BLN(BLN93),.WL(WL117));
sram_cell_6t_5 inst_cell_117_94 (.BL(BL94),.BLN(BLN94),.WL(WL117));
sram_cell_6t_5 inst_cell_117_95 (.BL(BL95),.BLN(BLN95),.WL(WL117));
sram_cell_6t_5 inst_cell_117_96 (.BL(BL96),.BLN(BLN96),.WL(WL117));
sram_cell_6t_5 inst_cell_117_97 (.BL(BL97),.BLN(BLN97),.WL(WL117));
sram_cell_6t_5 inst_cell_117_98 (.BL(BL98),.BLN(BLN98),.WL(WL117));
sram_cell_6t_5 inst_cell_117_99 (.BL(BL99),.BLN(BLN99),.WL(WL117));
sram_cell_6t_5 inst_cell_117_100 (.BL(BL100),.BLN(BLN100),.WL(WL117));
sram_cell_6t_5 inst_cell_117_101 (.BL(BL101),.BLN(BLN101),.WL(WL117));
sram_cell_6t_5 inst_cell_117_102 (.BL(BL102),.BLN(BLN102),.WL(WL117));
sram_cell_6t_5 inst_cell_117_103 (.BL(BL103),.BLN(BLN103),.WL(WL117));
sram_cell_6t_5 inst_cell_117_104 (.BL(BL104),.BLN(BLN104),.WL(WL117));
sram_cell_6t_5 inst_cell_117_105 (.BL(BL105),.BLN(BLN105),.WL(WL117));
sram_cell_6t_5 inst_cell_117_106 (.BL(BL106),.BLN(BLN106),.WL(WL117));
sram_cell_6t_5 inst_cell_117_107 (.BL(BL107),.BLN(BLN107),.WL(WL117));
sram_cell_6t_5 inst_cell_117_108 (.BL(BL108),.BLN(BLN108),.WL(WL117));
sram_cell_6t_5 inst_cell_117_109 (.BL(BL109),.BLN(BLN109),.WL(WL117));
sram_cell_6t_5 inst_cell_117_110 (.BL(BL110),.BLN(BLN110),.WL(WL117));
sram_cell_6t_5 inst_cell_117_111 (.BL(BL111),.BLN(BLN111),.WL(WL117));
sram_cell_6t_5 inst_cell_117_112 (.BL(BL112),.BLN(BLN112),.WL(WL117));
sram_cell_6t_5 inst_cell_117_113 (.BL(BL113),.BLN(BLN113),.WL(WL117));
sram_cell_6t_5 inst_cell_117_114 (.BL(BL114),.BLN(BLN114),.WL(WL117));
sram_cell_6t_5 inst_cell_117_115 (.BL(BL115),.BLN(BLN115),.WL(WL117));
sram_cell_6t_5 inst_cell_117_116 (.BL(BL116),.BLN(BLN116),.WL(WL117));
sram_cell_6t_5 inst_cell_117_117 (.BL(BL117),.BLN(BLN117),.WL(WL117));
sram_cell_6t_5 inst_cell_117_118 (.BL(BL118),.BLN(BLN118),.WL(WL117));
sram_cell_6t_5 inst_cell_117_119 (.BL(BL119),.BLN(BLN119),.WL(WL117));
sram_cell_6t_5 inst_cell_117_120 (.BL(BL120),.BLN(BLN120),.WL(WL117));
sram_cell_6t_5 inst_cell_117_121 (.BL(BL121),.BLN(BLN121),.WL(WL117));
sram_cell_6t_5 inst_cell_117_122 (.BL(BL122),.BLN(BLN122),.WL(WL117));
sram_cell_6t_5 inst_cell_117_123 (.BL(BL123),.BLN(BLN123),.WL(WL117));
sram_cell_6t_5 inst_cell_117_124 (.BL(BL124),.BLN(BLN124),.WL(WL117));
sram_cell_6t_5 inst_cell_117_125 (.BL(BL125),.BLN(BLN125),.WL(WL117));
sram_cell_6t_5 inst_cell_117_126 (.BL(BL126),.BLN(BLN126),.WL(WL117));
sram_cell_6t_5 inst_cell_117_127 (.BL(BL127),.BLN(BLN127),.WL(WL117));
sram_cell_6t_5 inst_cell_118_0 (.BL(BL0),.BLN(BLN0),.WL(WL118));
sram_cell_6t_5 inst_cell_118_1 (.BL(BL1),.BLN(BLN1),.WL(WL118));
sram_cell_6t_5 inst_cell_118_2 (.BL(BL2),.BLN(BLN2),.WL(WL118));
sram_cell_6t_5 inst_cell_118_3 (.BL(BL3),.BLN(BLN3),.WL(WL118));
sram_cell_6t_5 inst_cell_118_4 (.BL(BL4),.BLN(BLN4),.WL(WL118));
sram_cell_6t_5 inst_cell_118_5 (.BL(BL5),.BLN(BLN5),.WL(WL118));
sram_cell_6t_5 inst_cell_118_6 (.BL(BL6),.BLN(BLN6),.WL(WL118));
sram_cell_6t_5 inst_cell_118_7 (.BL(BL7),.BLN(BLN7),.WL(WL118));
sram_cell_6t_5 inst_cell_118_8 (.BL(BL8),.BLN(BLN8),.WL(WL118));
sram_cell_6t_5 inst_cell_118_9 (.BL(BL9),.BLN(BLN9),.WL(WL118));
sram_cell_6t_5 inst_cell_118_10 (.BL(BL10),.BLN(BLN10),.WL(WL118));
sram_cell_6t_5 inst_cell_118_11 (.BL(BL11),.BLN(BLN11),.WL(WL118));
sram_cell_6t_5 inst_cell_118_12 (.BL(BL12),.BLN(BLN12),.WL(WL118));
sram_cell_6t_5 inst_cell_118_13 (.BL(BL13),.BLN(BLN13),.WL(WL118));
sram_cell_6t_5 inst_cell_118_14 (.BL(BL14),.BLN(BLN14),.WL(WL118));
sram_cell_6t_5 inst_cell_118_15 (.BL(BL15),.BLN(BLN15),.WL(WL118));
sram_cell_6t_5 inst_cell_118_16 (.BL(BL16),.BLN(BLN16),.WL(WL118));
sram_cell_6t_5 inst_cell_118_17 (.BL(BL17),.BLN(BLN17),.WL(WL118));
sram_cell_6t_5 inst_cell_118_18 (.BL(BL18),.BLN(BLN18),.WL(WL118));
sram_cell_6t_5 inst_cell_118_19 (.BL(BL19),.BLN(BLN19),.WL(WL118));
sram_cell_6t_5 inst_cell_118_20 (.BL(BL20),.BLN(BLN20),.WL(WL118));
sram_cell_6t_5 inst_cell_118_21 (.BL(BL21),.BLN(BLN21),.WL(WL118));
sram_cell_6t_5 inst_cell_118_22 (.BL(BL22),.BLN(BLN22),.WL(WL118));
sram_cell_6t_5 inst_cell_118_23 (.BL(BL23),.BLN(BLN23),.WL(WL118));
sram_cell_6t_5 inst_cell_118_24 (.BL(BL24),.BLN(BLN24),.WL(WL118));
sram_cell_6t_5 inst_cell_118_25 (.BL(BL25),.BLN(BLN25),.WL(WL118));
sram_cell_6t_5 inst_cell_118_26 (.BL(BL26),.BLN(BLN26),.WL(WL118));
sram_cell_6t_5 inst_cell_118_27 (.BL(BL27),.BLN(BLN27),.WL(WL118));
sram_cell_6t_5 inst_cell_118_28 (.BL(BL28),.BLN(BLN28),.WL(WL118));
sram_cell_6t_5 inst_cell_118_29 (.BL(BL29),.BLN(BLN29),.WL(WL118));
sram_cell_6t_5 inst_cell_118_30 (.BL(BL30),.BLN(BLN30),.WL(WL118));
sram_cell_6t_5 inst_cell_118_31 (.BL(BL31),.BLN(BLN31),.WL(WL118));
sram_cell_6t_5 inst_cell_118_32 (.BL(BL32),.BLN(BLN32),.WL(WL118));
sram_cell_6t_5 inst_cell_118_33 (.BL(BL33),.BLN(BLN33),.WL(WL118));
sram_cell_6t_5 inst_cell_118_34 (.BL(BL34),.BLN(BLN34),.WL(WL118));
sram_cell_6t_5 inst_cell_118_35 (.BL(BL35),.BLN(BLN35),.WL(WL118));
sram_cell_6t_5 inst_cell_118_36 (.BL(BL36),.BLN(BLN36),.WL(WL118));
sram_cell_6t_5 inst_cell_118_37 (.BL(BL37),.BLN(BLN37),.WL(WL118));
sram_cell_6t_5 inst_cell_118_38 (.BL(BL38),.BLN(BLN38),.WL(WL118));
sram_cell_6t_5 inst_cell_118_39 (.BL(BL39),.BLN(BLN39),.WL(WL118));
sram_cell_6t_5 inst_cell_118_40 (.BL(BL40),.BLN(BLN40),.WL(WL118));
sram_cell_6t_5 inst_cell_118_41 (.BL(BL41),.BLN(BLN41),.WL(WL118));
sram_cell_6t_5 inst_cell_118_42 (.BL(BL42),.BLN(BLN42),.WL(WL118));
sram_cell_6t_5 inst_cell_118_43 (.BL(BL43),.BLN(BLN43),.WL(WL118));
sram_cell_6t_5 inst_cell_118_44 (.BL(BL44),.BLN(BLN44),.WL(WL118));
sram_cell_6t_5 inst_cell_118_45 (.BL(BL45),.BLN(BLN45),.WL(WL118));
sram_cell_6t_5 inst_cell_118_46 (.BL(BL46),.BLN(BLN46),.WL(WL118));
sram_cell_6t_5 inst_cell_118_47 (.BL(BL47),.BLN(BLN47),.WL(WL118));
sram_cell_6t_5 inst_cell_118_48 (.BL(BL48),.BLN(BLN48),.WL(WL118));
sram_cell_6t_5 inst_cell_118_49 (.BL(BL49),.BLN(BLN49),.WL(WL118));
sram_cell_6t_5 inst_cell_118_50 (.BL(BL50),.BLN(BLN50),.WL(WL118));
sram_cell_6t_5 inst_cell_118_51 (.BL(BL51),.BLN(BLN51),.WL(WL118));
sram_cell_6t_5 inst_cell_118_52 (.BL(BL52),.BLN(BLN52),.WL(WL118));
sram_cell_6t_5 inst_cell_118_53 (.BL(BL53),.BLN(BLN53),.WL(WL118));
sram_cell_6t_5 inst_cell_118_54 (.BL(BL54),.BLN(BLN54),.WL(WL118));
sram_cell_6t_5 inst_cell_118_55 (.BL(BL55),.BLN(BLN55),.WL(WL118));
sram_cell_6t_5 inst_cell_118_56 (.BL(BL56),.BLN(BLN56),.WL(WL118));
sram_cell_6t_5 inst_cell_118_57 (.BL(BL57),.BLN(BLN57),.WL(WL118));
sram_cell_6t_5 inst_cell_118_58 (.BL(BL58),.BLN(BLN58),.WL(WL118));
sram_cell_6t_5 inst_cell_118_59 (.BL(BL59),.BLN(BLN59),.WL(WL118));
sram_cell_6t_5 inst_cell_118_60 (.BL(BL60),.BLN(BLN60),.WL(WL118));
sram_cell_6t_5 inst_cell_118_61 (.BL(BL61),.BLN(BLN61),.WL(WL118));
sram_cell_6t_5 inst_cell_118_62 (.BL(BL62),.BLN(BLN62),.WL(WL118));
sram_cell_6t_5 inst_cell_118_63 (.BL(BL63),.BLN(BLN63),.WL(WL118));
sram_cell_6t_5 inst_cell_118_64 (.BL(BL64),.BLN(BLN64),.WL(WL118));
sram_cell_6t_5 inst_cell_118_65 (.BL(BL65),.BLN(BLN65),.WL(WL118));
sram_cell_6t_5 inst_cell_118_66 (.BL(BL66),.BLN(BLN66),.WL(WL118));
sram_cell_6t_5 inst_cell_118_67 (.BL(BL67),.BLN(BLN67),.WL(WL118));
sram_cell_6t_5 inst_cell_118_68 (.BL(BL68),.BLN(BLN68),.WL(WL118));
sram_cell_6t_5 inst_cell_118_69 (.BL(BL69),.BLN(BLN69),.WL(WL118));
sram_cell_6t_5 inst_cell_118_70 (.BL(BL70),.BLN(BLN70),.WL(WL118));
sram_cell_6t_5 inst_cell_118_71 (.BL(BL71),.BLN(BLN71),.WL(WL118));
sram_cell_6t_5 inst_cell_118_72 (.BL(BL72),.BLN(BLN72),.WL(WL118));
sram_cell_6t_5 inst_cell_118_73 (.BL(BL73),.BLN(BLN73),.WL(WL118));
sram_cell_6t_5 inst_cell_118_74 (.BL(BL74),.BLN(BLN74),.WL(WL118));
sram_cell_6t_5 inst_cell_118_75 (.BL(BL75),.BLN(BLN75),.WL(WL118));
sram_cell_6t_5 inst_cell_118_76 (.BL(BL76),.BLN(BLN76),.WL(WL118));
sram_cell_6t_5 inst_cell_118_77 (.BL(BL77),.BLN(BLN77),.WL(WL118));
sram_cell_6t_5 inst_cell_118_78 (.BL(BL78),.BLN(BLN78),.WL(WL118));
sram_cell_6t_5 inst_cell_118_79 (.BL(BL79),.BLN(BLN79),.WL(WL118));
sram_cell_6t_5 inst_cell_118_80 (.BL(BL80),.BLN(BLN80),.WL(WL118));
sram_cell_6t_5 inst_cell_118_81 (.BL(BL81),.BLN(BLN81),.WL(WL118));
sram_cell_6t_5 inst_cell_118_82 (.BL(BL82),.BLN(BLN82),.WL(WL118));
sram_cell_6t_5 inst_cell_118_83 (.BL(BL83),.BLN(BLN83),.WL(WL118));
sram_cell_6t_5 inst_cell_118_84 (.BL(BL84),.BLN(BLN84),.WL(WL118));
sram_cell_6t_5 inst_cell_118_85 (.BL(BL85),.BLN(BLN85),.WL(WL118));
sram_cell_6t_5 inst_cell_118_86 (.BL(BL86),.BLN(BLN86),.WL(WL118));
sram_cell_6t_5 inst_cell_118_87 (.BL(BL87),.BLN(BLN87),.WL(WL118));
sram_cell_6t_5 inst_cell_118_88 (.BL(BL88),.BLN(BLN88),.WL(WL118));
sram_cell_6t_5 inst_cell_118_89 (.BL(BL89),.BLN(BLN89),.WL(WL118));
sram_cell_6t_5 inst_cell_118_90 (.BL(BL90),.BLN(BLN90),.WL(WL118));
sram_cell_6t_5 inst_cell_118_91 (.BL(BL91),.BLN(BLN91),.WL(WL118));
sram_cell_6t_5 inst_cell_118_92 (.BL(BL92),.BLN(BLN92),.WL(WL118));
sram_cell_6t_5 inst_cell_118_93 (.BL(BL93),.BLN(BLN93),.WL(WL118));
sram_cell_6t_5 inst_cell_118_94 (.BL(BL94),.BLN(BLN94),.WL(WL118));
sram_cell_6t_5 inst_cell_118_95 (.BL(BL95),.BLN(BLN95),.WL(WL118));
sram_cell_6t_5 inst_cell_118_96 (.BL(BL96),.BLN(BLN96),.WL(WL118));
sram_cell_6t_5 inst_cell_118_97 (.BL(BL97),.BLN(BLN97),.WL(WL118));
sram_cell_6t_5 inst_cell_118_98 (.BL(BL98),.BLN(BLN98),.WL(WL118));
sram_cell_6t_5 inst_cell_118_99 (.BL(BL99),.BLN(BLN99),.WL(WL118));
sram_cell_6t_5 inst_cell_118_100 (.BL(BL100),.BLN(BLN100),.WL(WL118));
sram_cell_6t_5 inst_cell_118_101 (.BL(BL101),.BLN(BLN101),.WL(WL118));
sram_cell_6t_5 inst_cell_118_102 (.BL(BL102),.BLN(BLN102),.WL(WL118));
sram_cell_6t_5 inst_cell_118_103 (.BL(BL103),.BLN(BLN103),.WL(WL118));
sram_cell_6t_5 inst_cell_118_104 (.BL(BL104),.BLN(BLN104),.WL(WL118));
sram_cell_6t_5 inst_cell_118_105 (.BL(BL105),.BLN(BLN105),.WL(WL118));
sram_cell_6t_5 inst_cell_118_106 (.BL(BL106),.BLN(BLN106),.WL(WL118));
sram_cell_6t_5 inst_cell_118_107 (.BL(BL107),.BLN(BLN107),.WL(WL118));
sram_cell_6t_5 inst_cell_118_108 (.BL(BL108),.BLN(BLN108),.WL(WL118));
sram_cell_6t_5 inst_cell_118_109 (.BL(BL109),.BLN(BLN109),.WL(WL118));
sram_cell_6t_5 inst_cell_118_110 (.BL(BL110),.BLN(BLN110),.WL(WL118));
sram_cell_6t_5 inst_cell_118_111 (.BL(BL111),.BLN(BLN111),.WL(WL118));
sram_cell_6t_5 inst_cell_118_112 (.BL(BL112),.BLN(BLN112),.WL(WL118));
sram_cell_6t_5 inst_cell_118_113 (.BL(BL113),.BLN(BLN113),.WL(WL118));
sram_cell_6t_5 inst_cell_118_114 (.BL(BL114),.BLN(BLN114),.WL(WL118));
sram_cell_6t_5 inst_cell_118_115 (.BL(BL115),.BLN(BLN115),.WL(WL118));
sram_cell_6t_5 inst_cell_118_116 (.BL(BL116),.BLN(BLN116),.WL(WL118));
sram_cell_6t_5 inst_cell_118_117 (.BL(BL117),.BLN(BLN117),.WL(WL118));
sram_cell_6t_5 inst_cell_118_118 (.BL(BL118),.BLN(BLN118),.WL(WL118));
sram_cell_6t_5 inst_cell_118_119 (.BL(BL119),.BLN(BLN119),.WL(WL118));
sram_cell_6t_5 inst_cell_118_120 (.BL(BL120),.BLN(BLN120),.WL(WL118));
sram_cell_6t_5 inst_cell_118_121 (.BL(BL121),.BLN(BLN121),.WL(WL118));
sram_cell_6t_5 inst_cell_118_122 (.BL(BL122),.BLN(BLN122),.WL(WL118));
sram_cell_6t_5 inst_cell_118_123 (.BL(BL123),.BLN(BLN123),.WL(WL118));
sram_cell_6t_5 inst_cell_118_124 (.BL(BL124),.BLN(BLN124),.WL(WL118));
sram_cell_6t_5 inst_cell_118_125 (.BL(BL125),.BLN(BLN125),.WL(WL118));
sram_cell_6t_5 inst_cell_118_126 (.BL(BL126),.BLN(BLN126),.WL(WL118));
sram_cell_6t_5 inst_cell_118_127 (.BL(BL127),.BLN(BLN127),.WL(WL118));
sram_cell_6t_5 inst_cell_119_0 (.BL(BL0),.BLN(BLN0),.WL(WL119));
sram_cell_6t_5 inst_cell_119_1 (.BL(BL1),.BLN(BLN1),.WL(WL119));
sram_cell_6t_5 inst_cell_119_2 (.BL(BL2),.BLN(BLN2),.WL(WL119));
sram_cell_6t_5 inst_cell_119_3 (.BL(BL3),.BLN(BLN3),.WL(WL119));
sram_cell_6t_5 inst_cell_119_4 (.BL(BL4),.BLN(BLN4),.WL(WL119));
sram_cell_6t_5 inst_cell_119_5 (.BL(BL5),.BLN(BLN5),.WL(WL119));
sram_cell_6t_5 inst_cell_119_6 (.BL(BL6),.BLN(BLN6),.WL(WL119));
sram_cell_6t_5 inst_cell_119_7 (.BL(BL7),.BLN(BLN7),.WL(WL119));
sram_cell_6t_5 inst_cell_119_8 (.BL(BL8),.BLN(BLN8),.WL(WL119));
sram_cell_6t_5 inst_cell_119_9 (.BL(BL9),.BLN(BLN9),.WL(WL119));
sram_cell_6t_5 inst_cell_119_10 (.BL(BL10),.BLN(BLN10),.WL(WL119));
sram_cell_6t_5 inst_cell_119_11 (.BL(BL11),.BLN(BLN11),.WL(WL119));
sram_cell_6t_5 inst_cell_119_12 (.BL(BL12),.BLN(BLN12),.WL(WL119));
sram_cell_6t_5 inst_cell_119_13 (.BL(BL13),.BLN(BLN13),.WL(WL119));
sram_cell_6t_5 inst_cell_119_14 (.BL(BL14),.BLN(BLN14),.WL(WL119));
sram_cell_6t_5 inst_cell_119_15 (.BL(BL15),.BLN(BLN15),.WL(WL119));
sram_cell_6t_5 inst_cell_119_16 (.BL(BL16),.BLN(BLN16),.WL(WL119));
sram_cell_6t_5 inst_cell_119_17 (.BL(BL17),.BLN(BLN17),.WL(WL119));
sram_cell_6t_5 inst_cell_119_18 (.BL(BL18),.BLN(BLN18),.WL(WL119));
sram_cell_6t_5 inst_cell_119_19 (.BL(BL19),.BLN(BLN19),.WL(WL119));
sram_cell_6t_5 inst_cell_119_20 (.BL(BL20),.BLN(BLN20),.WL(WL119));
sram_cell_6t_5 inst_cell_119_21 (.BL(BL21),.BLN(BLN21),.WL(WL119));
sram_cell_6t_5 inst_cell_119_22 (.BL(BL22),.BLN(BLN22),.WL(WL119));
sram_cell_6t_5 inst_cell_119_23 (.BL(BL23),.BLN(BLN23),.WL(WL119));
sram_cell_6t_5 inst_cell_119_24 (.BL(BL24),.BLN(BLN24),.WL(WL119));
sram_cell_6t_5 inst_cell_119_25 (.BL(BL25),.BLN(BLN25),.WL(WL119));
sram_cell_6t_5 inst_cell_119_26 (.BL(BL26),.BLN(BLN26),.WL(WL119));
sram_cell_6t_5 inst_cell_119_27 (.BL(BL27),.BLN(BLN27),.WL(WL119));
sram_cell_6t_5 inst_cell_119_28 (.BL(BL28),.BLN(BLN28),.WL(WL119));
sram_cell_6t_5 inst_cell_119_29 (.BL(BL29),.BLN(BLN29),.WL(WL119));
sram_cell_6t_5 inst_cell_119_30 (.BL(BL30),.BLN(BLN30),.WL(WL119));
sram_cell_6t_5 inst_cell_119_31 (.BL(BL31),.BLN(BLN31),.WL(WL119));
sram_cell_6t_5 inst_cell_119_32 (.BL(BL32),.BLN(BLN32),.WL(WL119));
sram_cell_6t_5 inst_cell_119_33 (.BL(BL33),.BLN(BLN33),.WL(WL119));
sram_cell_6t_5 inst_cell_119_34 (.BL(BL34),.BLN(BLN34),.WL(WL119));
sram_cell_6t_5 inst_cell_119_35 (.BL(BL35),.BLN(BLN35),.WL(WL119));
sram_cell_6t_5 inst_cell_119_36 (.BL(BL36),.BLN(BLN36),.WL(WL119));
sram_cell_6t_5 inst_cell_119_37 (.BL(BL37),.BLN(BLN37),.WL(WL119));
sram_cell_6t_5 inst_cell_119_38 (.BL(BL38),.BLN(BLN38),.WL(WL119));
sram_cell_6t_5 inst_cell_119_39 (.BL(BL39),.BLN(BLN39),.WL(WL119));
sram_cell_6t_5 inst_cell_119_40 (.BL(BL40),.BLN(BLN40),.WL(WL119));
sram_cell_6t_5 inst_cell_119_41 (.BL(BL41),.BLN(BLN41),.WL(WL119));
sram_cell_6t_5 inst_cell_119_42 (.BL(BL42),.BLN(BLN42),.WL(WL119));
sram_cell_6t_5 inst_cell_119_43 (.BL(BL43),.BLN(BLN43),.WL(WL119));
sram_cell_6t_5 inst_cell_119_44 (.BL(BL44),.BLN(BLN44),.WL(WL119));
sram_cell_6t_5 inst_cell_119_45 (.BL(BL45),.BLN(BLN45),.WL(WL119));
sram_cell_6t_5 inst_cell_119_46 (.BL(BL46),.BLN(BLN46),.WL(WL119));
sram_cell_6t_5 inst_cell_119_47 (.BL(BL47),.BLN(BLN47),.WL(WL119));
sram_cell_6t_5 inst_cell_119_48 (.BL(BL48),.BLN(BLN48),.WL(WL119));
sram_cell_6t_5 inst_cell_119_49 (.BL(BL49),.BLN(BLN49),.WL(WL119));
sram_cell_6t_5 inst_cell_119_50 (.BL(BL50),.BLN(BLN50),.WL(WL119));
sram_cell_6t_5 inst_cell_119_51 (.BL(BL51),.BLN(BLN51),.WL(WL119));
sram_cell_6t_5 inst_cell_119_52 (.BL(BL52),.BLN(BLN52),.WL(WL119));
sram_cell_6t_5 inst_cell_119_53 (.BL(BL53),.BLN(BLN53),.WL(WL119));
sram_cell_6t_5 inst_cell_119_54 (.BL(BL54),.BLN(BLN54),.WL(WL119));
sram_cell_6t_5 inst_cell_119_55 (.BL(BL55),.BLN(BLN55),.WL(WL119));
sram_cell_6t_5 inst_cell_119_56 (.BL(BL56),.BLN(BLN56),.WL(WL119));
sram_cell_6t_5 inst_cell_119_57 (.BL(BL57),.BLN(BLN57),.WL(WL119));
sram_cell_6t_5 inst_cell_119_58 (.BL(BL58),.BLN(BLN58),.WL(WL119));
sram_cell_6t_5 inst_cell_119_59 (.BL(BL59),.BLN(BLN59),.WL(WL119));
sram_cell_6t_5 inst_cell_119_60 (.BL(BL60),.BLN(BLN60),.WL(WL119));
sram_cell_6t_5 inst_cell_119_61 (.BL(BL61),.BLN(BLN61),.WL(WL119));
sram_cell_6t_5 inst_cell_119_62 (.BL(BL62),.BLN(BLN62),.WL(WL119));
sram_cell_6t_5 inst_cell_119_63 (.BL(BL63),.BLN(BLN63),.WL(WL119));
sram_cell_6t_5 inst_cell_119_64 (.BL(BL64),.BLN(BLN64),.WL(WL119));
sram_cell_6t_5 inst_cell_119_65 (.BL(BL65),.BLN(BLN65),.WL(WL119));
sram_cell_6t_5 inst_cell_119_66 (.BL(BL66),.BLN(BLN66),.WL(WL119));
sram_cell_6t_5 inst_cell_119_67 (.BL(BL67),.BLN(BLN67),.WL(WL119));
sram_cell_6t_5 inst_cell_119_68 (.BL(BL68),.BLN(BLN68),.WL(WL119));
sram_cell_6t_5 inst_cell_119_69 (.BL(BL69),.BLN(BLN69),.WL(WL119));
sram_cell_6t_5 inst_cell_119_70 (.BL(BL70),.BLN(BLN70),.WL(WL119));
sram_cell_6t_5 inst_cell_119_71 (.BL(BL71),.BLN(BLN71),.WL(WL119));
sram_cell_6t_5 inst_cell_119_72 (.BL(BL72),.BLN(BLN72),.WL(WL119));
sram_cell_6t_5 inst_cell_119_73 (.BL(BL73),.BLN(BLN73),.WL(WL119));
sram_cell_6t_5 inst_cell_119_74 (.BL(BL74),.BLN(BLN74),.WL(WL119));
sram_cell_6t_5 inst_cell_119_75 (.BL(BL75),.BLN(BLN75),.WL(WL119));
sram_cell_6t_5 inst_cell_119_76 (.BL(BL76),.BLN(BLN76),.WL(WL119));
sram_cell_6t_5 inst_cell_119_77 (.BL(BL77),.BLN(BLN77),.WL(WL119));
sram_cell_6t_5 inst_cell_119_78 (.BL(BL78),.BLN(BLN78),.WL(WL119));
sram_cell_6t_5 inst_cell_119_79 (.BL(BL79),.BLN(BLN79),.WL(WL119));
sram_cell_6t_5 inst_cell_119_80 (.BL(BL80),.BLN(BLN80),.WL(WL119));
sram_cell_6t_5 inst_cell_119_81 (.BL(BL81),.BLN(BLN81),.WL(WL119));
sram_cell_6t_5 inst_cell_119_82 (.BL(BL82),.BLN(BLN82),.WL(WL119));
sram_cell_6t_5 inst_cell_119_83 (.BL(BL83),.BLN(BLN83),.WL(WL119));
sram_cell_6t_5 inst_cell_119_84 (.BL(BL84),.BLN(BLN84),.WL(WL119));
sram_cell_6t_5 inst_cell_119_85 (.BL(BL85),.BLN(BLN85),.WL(WL119));
sram_cell_6t_5 inst_cell_119_86 (.BL(BL86),.BLN(BLN86),.WL(WL119));
sram_cell_6t_5 inst_cell_119_87 (.BL(BL87),.BLN(BLN87),.WL(WL119));
sram_cell_6t_5 inst_cell_119_88 (.BL(BL88),.BLN(BLN88),.WL(WL119));
sram_cell_6t_5 inst_cell_119_89 (.BL(BL89),.BLN(BLN89),.WL(WL119));
sram_cell_6t_5 inst_cell_119_90 (.BL(BL90),.BLN(BLN90),.WL(WL119));
sram_cell_6t_5 inst_cell_119_91 (.BL(BL91),.BLN(BLN91),.WL(WL119));
sram_cell_6t_5 inst_cell_119_92 (.BL(BL92),.BLN(BLN92),.WL(WL119));
sram_cell_6t_5 inst_cell_119_93 (.BL(BL93),.BLN(BLN93),.WL(WL119));
sram_cell_6t_5 inst_cell_119_94 (.BL(BL94),.BLN(BLN94),.WL(WL119));
sram_cell_6t_5 inst_cell_119_95 (.BL(BL95),.BLN(BLN95),.WL(WL119));
sram_cell_6t_5 inst_cell_119_96 (.BL(BL96),.BLN(BLN96),.WL(WL119));
sram_cell_6t_5 inst_cell_119_97 (.BL(BL97),.BLN(BLN97),.WL(WL119));
sram_cell_6t_5 inst_cell_119_98 (.BL(BL98),.BLN(BLN98),.WL(WL119));
sram_cell_6t_5 inst_cell_119_99 (.BL(BL99),.BLN(BLN99),.WL(WL119));
sram_cell_6t_5 inst_cell_119_100 (.BL(BL100),.BLN(BLN100),.WL(WL119));
sram_cell_6t_5 inst_cell_119_101 (.BL(BL101),.BLN(BLN101),.WL(WL119));
sram_cell_6t_5 inst_cell_119_102 (.BL(BL102),.BLN(BLN102),.WL(WL119));
sram_cell_6t_5 inst_cell_119_103 (.BL(BL103),.BLN(BLN103),.WL(WL119));
sram_cell_6t_5 inst_cell_119_104 (.BL(BL104),.BLN(BLN104),.WL(WL119));
sram_cell_6t_5 inst_cell_119_105 (.BL(BL105),.BLN(BLN105),.WL(WL119));
sram_cell_6t_5 inst_cell_119_106 (.BL(BL106),.BLN(BLN106),.WL(WL119));
sram_cell_6t_5 inst_cell_119_107 (.BL(BL107),.BLN(BLN107),.WL(WL119));
sram_cell_6t_5 inst_cell_119_108 (.BL(BL108),.BLN(BLN108),.WL(WL119));
sram_cell_6t_5 inst_cell_119_109 (.BL(BL109),.BLN(BLN109),.WL(WL119));
sram_cell_6t_5 inst_cell_119_110 (.BL(BL110),.BLN(BLN110),.WL(WL119));
sram_cell_6t_5 inst_cell_119_111 (.BL(BL111),.BLN(BLN111),.WL(WL119));
sram_cell_6t_5 inst_cell_119_112 (.BL(BL112),.BLN(BLN112),.WL(WL119));
sram_cell_6t_5 inst_cell_119_113 (.BL(BL113),.BLN(BLN113),.WL(WL119));
sram_cell_6t_5 inst_cell_119_114 (.BL(BL114),.BLN(BLN114),.WL(WL119));
sram_cell_6t_5 inst_cell_119_115 (.BL(BL115),.BLN(BLN115),.WL(WL119));
sram_cell_6t_5 inst_cell_119_116 (.BL(BL116),.BLN(BLN116),.WL(WL119));
sram_cell_6t_5 inst_cell_119_117 (.BL(BL117),.BLN(BLN117),.WL(WL119));
sram_cell_6t_5 inst_cell_119_118 (.BL(BL118),.BLN(BLN118),.WL(WL119));
sram_cell_6t_5 inst_cell_119_119 (.BL(BL119),.BLN(BLN119),.WL(WL119));
sram_cell_6t_5 inst_cell_119_120 (.BL(BL120),.BLN(BLN120),.WL(WL119));
sram_cell_6t_5 inst_cell_119_121 (.BL(BL121),.BLN(BLN121),.WL(WL119));
sram_cell_6t_5 inst_cell_119_122 (.BL(BL122),.BLN(BLN122),.WL(WL119));
sram_cell_6t_5 inst_cell_119_123 (.BL(BL123),.BLN(BLN123),.WL(WL119));
sram_cell_6t_5 inst_cell_119_124 (.BL(BL124),.BLN(BLN124),.WL(WL119));
sram_cell_6t_5 inst_cell_119_125 (.BL(BL125),.BLN(BLN125),.WL(WL119));
sram_cell_6t_5 inst_cell_119_126 (.BL(BL126),.BLN(BLN126),.WL(WL119));
sram_cell_6t_5 inst_cell_119_127 (.BL(BL127),.BLN(BLN127),.WL(WL119));
sram_cell_6t_5 inst_cell_120_0 (.BL(BL0),.BLN(BLN0),.WL(WL120));
sram_cell_6t_5 inst_cell_120_1 (.BL(BL1),.BLN(BLN1),.WL(WL120));
sram_cell_6t_5 inst_cell_120_2 (.BL(BL2),.BLN(BLN2),.WL(WL120));
sram_cell_6t_5 inst_cell_120_3 (.BL(BL3),.BLN(BLN3),.WL(WL120));
sram_cell_6t_5 inst_cell_120_4 (.BL(BL4),.BLN(BLN4),.WL(WL120));
sram_cell_6t_5 inst_cell_120_5 (.BL(BL5),.BLN(BLN5),.WL(WL120));
sram_cell_6t_5 inst_cell_120_6 (.BL(BL6),.BLN(BLN6),.WL(WL120));
sram_cell_6t_5 inst_cell_120_7 (.BL(BL7),.BLN(BLN7),.WL(WL120));
sram_cell_6t_5 inst_cell_120_8 (.BL(BL8),.BLN(BLN8),.WL(WL120));
sram_cell_6t_5 inst_cell_120_9 (.BL(BL9),.BLN(BLN9),.WL(WL120));
sram_cell_6t_5 inst_cell_120_10 (.BL(BL10),.BLN(BLN10),.WL(WL120));
sram_cell_6t_5 inst_cell_120_11 (.BL(BL11),.BLN(BLN11),.WL(WL120));
sram_cell_6t_5 inst_cell_120_12 (.BL(BL12),.BLN(BLN12),.WL(WL120));
sram_cell_6t_5 inst_cell_120_13 (.BL(BL13),.BLN(BLN13),.WL(WL120));
sram_cell_6t_5 inst_cell_120_14 (.BL(BL14),.BLN(BLN14),.WL(WL120));
sram_cell_6t_5 inst_cell_120_15 (.BL(BL15),.BLN(BLN15),.WL(WL120));
sram_cell_6t_5 inst_cell_120_16 (.BL(BL16),.BLN(BLN16),.WL(WL120));
sram_cell_6t_5 inst_cell_120_17 (.BL(BL17),.BLN(BLN17),.WL(WL120));
sram_cell_6t_5 inst_cell_120_18 (.BL(BL18),.BLN(BLN18),.WL(WL120));
sram_cell_6t_5 inst_cell_120_19 (.BL(BL19),.BLN(BLN19),.WL(WL120));
sram_cell_6t_5 inst_cell_120_20 (.BL(BL20),.BLN(BLN20),.WL(WL120));
sram_cell_6t_5 inst_cell_120_21 (.BL(BL21),.BLN(BLN21),.WL(WL120));
sram_cell_6t_5 inst_cell_120_22 (.BL(BL22),.BLN(BLN22),.WL(WL120));
sram_cell_6t_5 inst_cell_120_23 (.BL(BL23),.BLN(BLN23),.WL(WL120));
sram_cell_6t_5 inst_cell_120_24 (.BL(BL24),.BLN(BLN24),.WL(WL120));
sram_cell_6t_5 inst_cell_120_25 (.BL(BL25),.BLN(BLN25),.WL(WL120));
sram_cell_6t_5 inst_cell_120_26 (.BL(BL26),.BLN(BLN26),.WL(WL120));
sram_cell_6t_5 inst_cell_120_27 (.BL(BL27),.BLN(BLN27),.WL(WL120));
sram_cell_6t_5 inst_cell_120_28 (.BL(BL28),.BLN(BLN28),.WL(WL120));
sram_cell_6t_5 inst_cell_120_29 (.BL(BL29),.BLN(BLN29),.WL(WL120));
sram_cell_6t_5 inst_cell_120_30 (.BL(BL30),.BLN(BLN30),.WL(WL120));
sram_cell_6t_5 inst_cell_120_31 (.BL(BL31),.BLN(BLN31),.WL(WL120));
sram_cell_6t_5 inst_cell_120_32 (.BL(BL32),.BLN(BLN32),.WL(WL120));
sram_cell_6t_5 inst_cell_120_33 (.BL(BL33),.BLN(BLN33),.WL(WL120));
sram_cell_6t_5 inst_cell_120_34 (.BL(BL34),.BLN(BLN34),.WL(WL120));
sram_cell_6t_5 inst_cell_120_35 (.BL(BL35),.BLN(BLN35),.WL(WL120));
sram_cell_6t_5 inst_cell_120_36 (.BL(BL36),.BLN(BLN36),.WL(WL120));
sram_cell_6t_5 inst_cell_120_37 (.BL(BL37),.BLN(BLN37),.WL(WL120));
sram_cell_6t_5 inst_cell_120_38 (.BL(BL38),.BLN(BLN38),.WL(WL120));
sram_cell_6t_5 inst_cell_120_39 (.BL(BL39),.BLN(BLN39),.WL(WL120));
sram_cell_6t_5 inst_cell_120_40 (.BL(BL40),.BLN(BLN40),.WL(WL120));
sram_cell_6t_5 inst_cell_120_41 (.BL(BL41),.BLN(BLN41),.WL(WL120));
sram_cell_6t_5 inst_cell_120_42 (.BL(BL42),.BLN(BLN42),.WL(WL120));
sram_cell_6t_5 inst_cell_120_43 (.BL(BL43),.BLN(BLN43),.WL(WL120));
sram_cell_6t_5 inst_cell_120_44 (.BL(BL44),.BLN(BLN44),.WL(WL120));
sram_cell_6t_5 inst_cell_120_45 (.BL(BL45),.BLN(BLN45),.WL(WL120));
sram_cell_6t_5 inst_cell_120_46 (.BL(BL46),.BLN(BLN46),.WL(WL120));
sram_cell_6t_5 inst_cell_120_47 (.BL(BL47),.BLN(BLN47),.WL(WL120));
sram_cell_6t_5 inst_cell_120_48 (.BL(BL48),.BLN(BLN48),.WL(WL120));
sram_cell_6t_5 inst_cell_120_49 (.BL(BL49),.BLN(BLN49),.WL(WL120));
sram_cell_6t_5 inst_cell_120_50 (.BL(BL50),.BLN(BLN50),.WL(WL120));
sram_cell_6t_5 inst_cell_120_51 (.BL(BL51),.BLN(BLN51),.WL(WL120));
sram_cell_6t_5 inst_cell_120_52 (.BL(BL52),.BLN(BLN52),.WL(WL120));
sram_cell_6t_5 inst_cell_120_53 (.BL(BL53),.BLN(BLN53),.WL(WL120));
sram_cell_6t_5 inst_cell_120_54 (.BL(BL54),.BLN(BLN54),.WL(WL120));
sram_cell_6t_5 inst_cell_120_55 (.BL(BL55),.BLN(BLN55),.WL(WL120));
sram_cell_6t_5 inst_cell_120_56 (.BL(BL56),.BLN(BLN56),.WL(WL120));
sram_cell_6t_5 inst_cell_120_57 (.BL(BL57),.BLN(BLN57),.WL(WL120));
sram_cell_6t_5 inst_cell_120_58 (.BL(BL58),.BLN(BLN58),.WL(WL120));
sram_cell_6t_5 inst_cell_120_59 (.BL(BL59),.BLN(BLN59),.WL(WL120));
sram_cell_6t_5 inst_cell_120_60 (.BL(BL60),.BLN(BLN60),.WL(WL120));
sram_cell_6t_5 inst_cell_120_61 (.BL(BL61),.BLN(BLN61),.WL(WL120));
sram_cell_6t_5 inst_cell_120_62 (.BL(BL62),.BLN(BLN62),.WL(WL120));
sram_cell_6t_5 inst_cell_120_63 (.BL(BL63),.BLN(BLN63),.WL(WL120));
sram_cell_6t_5 inst_cell_120_64 (.BL(BL64),.BLN(BLN64),.WL(WL120));
sram_cell_6t_5 inst_cell_120_65 (.BL(BL65),.BLN(BLN65),.WL(WL120));
sram_cell_6t_5 inst_cell_120_66 (.BL(BL66),.BLN(BLN66),.WL(WL120));
sram_cell_6t_5 inst_cell_120_67 (.BL(BL67),.BLN(BLN67),.WL(WL120));
sram_cell_6t_5 inst_cell_120_68 (.BL(BL68),.BLN(BLN68),.WL(WL120));
sram_cell_6t_5 inst_cell_120_69 (.BL(BL69),.BLN(BLN69),.WL(WL120));
sram_cell_6t_5 inst_cell_120_70 (.BL(BL70),.BLN(BLN70),.WL(WL120));
sram_cell_6t_5 inst_cell_120_71 (.BL(BL71),.BLN(BLN71),.WL(WL120));
sram_cell_6t_5 inst_cell_120_72 (.BL(BL72),.BLN(BLN72),.WL(WL120));
sram_cell_6t_5 inst_cell_120_73 (.BL(BL73),.BLN(BLN73),.WL(WL120));
sram_cell_6t_5 inst_cell_120_74 (.BL(BL74),.BLN(BLN74),.WL(WL120));
sram_cell_6t_5 inst_cell_120_75 (.BL(BL75),.BLN(BLN75),.WL(WL120));
sram_cell_6t_5 inst_cell_120_76 (.BL(BL76),.BLN(BLN76),.WL(WL120));
sram_cell_6t_5 inst_cell_120_77 (.BL(BL77),.BLN(BLN77),.WL(WL120));
sram_cell_6t_5 inst_cell_120_78 (.BL(BL78),.BLN(BLN78),.WL(WL120));
sram_cell_6t_5 inst_cell_120_79 (.BL(BL79),.BLN(BLN79),.WL(WL120));
sram_cell_6t_5 inst_cell_120_80 (.BL(BL80),.BLN(BLN80),.WL(WL120));
sram_cell_6t_5 inst_cell_120_81 (.BL(BL81),.BLN(BLN81),.WL(WL120));
sram_cell_6t_5 inst_cell_120_82 (.BL(BL82),.BLN(BLN82),.WL(WL120));
sram_cell_6t_5 inst_cell_120_83 (.BL(BL83),.BLN(BLN83),.WL(WL120));
sram_cell_6t_5 inst_cell_120_84 (.BL(BL84),.BLN(BLN84),.WL(WL120));
sram_cell_6t_5 inst_cell_120_85 (.BL(BL85),.BLN(BLN85),.WL(WL120));
sram_cell_6t_5 inst_cell_120_86 (.BL(BL86),.BLN(BLN86),.WL(WL120));
sram_cell_6t_5 inst_cell_120_87 (.BL(BL87),.BLN(BLN87),.WL(WL120));
sram_cell_6t_5 inst_cell_120_88 (.BL(BL88),.BLN(BLN88),.WL(WL120));
sram_cell_6t_5 inst_cell_120_89 (.BL(BL89),.BLN(BLN89),.WL(WL120));
sram_cell_6t_5 inst_cell_120_90 (.BL(BL90),.BLN(BLN90),.WL(WL120));
sram_cell_6t_5 inst_cell_120_91 (.BL(BL91),.BLN(BLN91),.WL(WL120));
sram_cell_6t_5 inst_cell_120_92 (.BL(BL92),.BLN(BLN92),.WL(WL120));
sram_cell_6t_5 inst_cell_120_93 (.BL(BL93),.BLN(BLN93),.WL(WL120));
sram_cell_6t_5 inst_cell_120_94 (.BL(BL94),.BLN(BLN94),.WL(WL120));
sram_cell_6t_5 inst_cell_120_95 (.BL(BL95),.BLN(BLN95),.WL(WL120));
sram_cell_6t_5 inst_cell_120_96 (.BL(BL96),.BLN(BLN96),.WL(WL120));
sram_cell_6t_5 inst_cell_120_97 (.BL(BL97),.BLN(BLN97),.WL(WL120));
sram_cell_6t_5 inst_cell_120_98 (.BL(BL98),.BLN(BLN98),.WL(WL120));
sram_cell_6t_5 inst_cell_120_99 (.BL(BL99),.BLN(BLN99),.WL(WL120));
sram_cell_6t_5 inst_cell_120_100 (.BL(BL100),.BLN(BLN100),.WL(WL120));
sram_cell_6t_5 inst_cell_120_101 (.BL(BL101),.BLN(BLN101),.WL(WL120));
sram_cell_6t_5 inst_cell_120_102 (.BL(BL102),.BLN(BLN102),.WL(WL120));
sram_cell_6t_5 inst_cell_120_103 (.BL(BL103),.BLN(BLN103),.WL(WL120));
sram_cell_6t_5 inst_cell_120_104 (.BL(BL104),.BLN(BLN104),.WL(WL120));
sram_cell_6t_5 inst_cell_120_105 (.BL(BL105),.BLN(BLN105),.WL(WL120));
sram_cell_6t_5 inst_cell_120_106 (.BL(BL106),.BLN(BLN106),.WL(WL120));
sram_cell_6t_5 inst_cell_120_107 (.BL(BL107),.BLN(BLN107),.WL(WL120));
sram_cell_6t_5 inst_cell_120_108 (.BL(BL108),.BLN(BLN108),.WL(WL120));
sram_cell_6t_5 inst_cell_120_109 (.BL(BL109),.BLN(BLN109),.WL(WL120));
sram_cell_6t_5 inst_cell_120_110 (.BL(BL110),.BLN(BLN110),.WL(WL120));
sram_cell_6t_5 inst_cell_120_111 (.BL(BL111),.BLN(BLN111),.WL(WL120));
sram_cell_6t_5 inst_cell_120_112 (.BL(BL112),.BLN(BLN112),.WL(WL120));
sram_cell_6t_5 inst_cell_120_113 (.BL(BL113),.BLN(BLN113),.WL(WL120));
sram_cell_6t_5 inst_cell_120_114 (.BL(BL114),.BLN(BLN114),.WL(WL120));
sram_cell_6t_5 inst_cell_120_115 (.BL(BL115),.BLN(BLN115),.WL(WL120));
sram_cell_6t_5 inst_cell_120_116 (.BL(BL116),.BLN(BLN116),.WL(WL120));
sram_cell_6t_5 inst_cell_120_117 (.BL(BL117),.BLN(BLN117),.WL(WL120));
sram_cell_6t_5 inst_cell_120_118 (.BL(BL118),.BLN(BLN118),.WL(WL120));
sram_cell_6t_5 inst_cell_120_119 (.BL(BL119),.BLN(BLN119),.WL(WL120));
sram_cell_6t_5 inst_cell_120_120 (.BL(BL120),.BLN(BLN120),.WL(WL120));
sram_cell_6t_5 inst_cell_120_121 (.BL(BL121),.BLN(BLN121),.WL(WL120));
sram_cell_6t_5 inst_cell_120_122 (.BL(BL122),.BLN(BLN122),.WL(WL120));
sram_cell_6t_5 inst_cell_120_123 (.BL(BL123),.BLN(BLN123),.WL(WL120));
sram_cell_6t_5 inst_cell_120_124 (.BL(BL124),.BLN(BLN124),.WL(WL120));
sram_cell_6t_5 inst_cell_120_125 (.BL(BL125),.BLN(BLN125),.WL(WL120));
sram_cell_6t_5 inst_cell_120_126 (.BL(BL126),.BLN(BLN126),.WL(WL120));
sram_cell_6t_5 inst_cell_120_127 (.BL(BL127),.BLN(BLN127),.WL(WL120));
sram_cell_6t_5 inst_cell_121_0 (.BL(BL0),.BLN(BLN0),.WL(WL121));
sram_cell_6t_5 inst_cell_121_1 (.BL(BL1),.BLN(BLN1),.WL(WL121));
sram_cell_6t_5 inst_cell_121_2 (.BL(BL2),.BLN(BLN2),.WL(WL121));
sram_cell_6t_5 inst_cell_121_3 (.BL(BL3),.BLN(BLN3),.WL(WL121));
sram_cell_6t_5 inst_cell_121_4 (.BL(BL4),.BLN(BLN4),.WL(WL121));
sram_cell_6t_5 inst_cell_121_5 (.BL(BL5),.BLN(BLN5),.WL(WL121));
sram_cell_6t_5 inst_cell_121_6 (.BL(BL6),.BLN(BLN6),.WL(WL121));
sram_cell_6t_5 inst_cell_121_7 (.BL(BL7),.BLN(BLN7),.WL(WL121));
sram_cell_6t_5 inst_cell_121_8 (.BL(BL8),.BLN(BLN8),.WL(WL121));
sram_cell_6t_5 inst_cell_121_9 (.BL(BL9),.BLN(BLN9),.WL(WL121));
sram_cell_6t_5 inst_cell_121_10 (.BL(BL10),.BLN(BLN10),.WL(WL121));
sram_cell_6t_5 inst_cell_121_11 (.BL(BL11),.BLN(BLN11),.WL(WL121));
sram_cell_6t_5 inst_cell_121_12 (.BL(BL12),.BLN(BLN12),.WL(WL121));
sram_cell_6t_5 inst_cell_121_13 (.BL(BL13),.BLN(BLN13),.WL(WL121));
sram_cell_6t_5 inst_cell_121_14 (.BL(BL14),.BLN(BLN14),.WL(WL121));
sram_cell_6t_5 inst_cell_121_15 (.BL(BL15),.BLN(BLN15),.WL(WL121));
sram_cell_6t_5 inst_cell_121_16 (.BL(BL16),.BLN(BLN16),.WL(WL121));
sram_cell_6t_5 inst_cell_121_17 (.BL(BL17),.BLN(BLN17),.WL(WL121));
sram_cell_6t_5 inst_cell_121_18 (.BL(BL18),.BLN(BLN18),.WL(WL121));
sram_cell_6t_5 inst_cell_121_19 (.BL(BL19),.BLN(BLN19),.WL(WL121));
sram_cell_6t_5 inst_cell_121_20 (.BL(BL20),.BLN(BLN20),.WL(WL121));
sram_cell_6t_5 inst_cell_121_21 (.BL(BL21),.BLN(BLN21),.WL(WL121));
sram_cell_6t_5 inst_cell_121_22 (.BL(BL22),.BLN(BLN22),.WL(WL121));
sram_cell_6t_5 inst_cell_121_23 (.BL(BL23),.BLN(BLN23),.WL(WL121));
sram_cell_6t_5 inst_cell_121_24 (.BL(BL24),.BLN(BLN24),.WL(WL121));
sram_cell_6t_5 inst_cell_121_25 (.BL(BL25),.BLN(BLN25),.WL(WL121));
sram_cell_6t_5 inst_cell_121_26 (.BL(BL26),.BLN(BLN26),.WL(WL121));
sram_cell_6t_5 inst_cell_121_27 (.BL(BL27),.BLN(BLN27),.WL(WL121));
sram_cell_6t_5 inst_cell_121_28 (.BL(BL28),.BLN(BLN28),.WL(WL121));
sram_cell_6t_5 inst_cell_121_29 (.BL(BL29),.BLN(BLN29),.WL(WL121));
sram_cell_6t_5 inst_cell_121_30 (.BL(BL30),.BLN(BLN30),.WL(WL121));
sram_cell_6t_5 inst_cell_121_31 (.BL(BL31),.BLN(BLN31),.WL(WL121));
sram_cell_6t_5 inst_cell_121_32 (.BL(BL32),.BLN(BLN32),.WL(WL121));
sram_cell_6t_5 inst_cell_121_33 (.BL(BL33),.BLN(BLN33),.WL(WL121));
sram_cell_6t_5 inst_cell_121_34 (.BL(BL34),.BLN(BLN34),.WL(WL121));
sram_cell_6t_5 inst_cell_121_35 (.BL(BL35),.BLN(BLN35),.WL(WL121));
sram_cell_6t_5 inst_cell_121_36 (.BL(BL36),.BLN(BLN36),.WL(WL121));
sram_cell_6t_5 inst_cell_121_37 (.BL(BL37),.BLN(BLN37),.WL(WL121));
sram_cell_6t_5 inst_cell_121_38 (.BL(BL38),.BLN(BLN38),.WL(WL121));
sram_cell_6t_5 inst_cell_121_39 (.BL(BL39),.BLN(BLN39),.WL(WL121));
sram_cell_6t_5 inst_cell_121_40 (.BL(BL40),.BLN(BLN40),.WL(WL121));
sram_cell_6t_5 inst_cell_121_41 (.BL(BL41),.BLN(BLN41),.WL(WL121));
sram_cell_6t_5 inst_cell_121_42 (.BL(BL42),.BLN(BLN42),.WL(WL121));
sram_cell_6t_5 inst_cell_121_43 (.BL(BL43),.BLN(BLN43),.WL(WL121));
sram_cell_6t_5 inst_cell_121_44 (.BL(BL44),.BLN(BLN44),.WL(WL121));
sram_cell_6t_5 inst_cell_121_45 (.BL(BL45),.BLN(BLN45),.WL(WL121));
sram_cell_6t_5 inst_cell_121_46 (.BL(BL46),.BLN(BLN46),.WL(WL121));
sram_cell_6t_5 inst_cell_121_47 (.BL(BL47),.BLN(BLN47),.WL(WL121));
sram_cell_6t_5 inst_cell_121_48 (.BL(BL48),.BLN(BLN48),.WL(WL121));
sram_cell_6t_5 inst_cell_121_49 (.BL(BL49),.BLN(BLN49),.WL(WL121));
sram_cell_6t_5 inst_cell_121_50 (.BL(BL50),.BLN(BLN50),.WL(WL121));
sram_cell_6t_5 inst_cell_121_51 (.BL(BL51),.BLN(BLN51),.WL(WL121));
sram_cell_6t_5 inst_cell_121_52 (.BL(BL52),.BLN(BLN52),.WL(WL121));
sram_cell_6t_5 inst_cell_121_53 (.BL(BL53),.BLN(BLN53),.WL(WL121));
sram_cell_6t_5 inst_cell_121_54 (.BL(BL54),.BLN(BLN54),.WL(WL121));
sram_cell_6t_5 inst_cell_121_55 (.BL(BL55),.BLN(BLN55),.WL(WL121));
sram_cell_6t_5 inst_cell_121_56 (.BL(BL56),.BLN(BLN56),.WL(WL121));
sram_cell_6t_5 inst_cell_121_57 (.BL(BL57),.BLN(BLN57),.WL(WL121));
sram_cell_6t_5 inst_cell_121_58 (.BL(BL58),.BLN(BLN58),.WL(WL121));
sram_cell_6t_5 inst_cell_121_59 (.BL(BL59),.BLN(BLN59),.WL(WL121));
sram_cell_6t_5 inst_cell_121_60 (.BL(BL60),.BLN(BLN60),.WL(WL121));
sram_cell_6t_5 inst_cell_121_61 (.BL(BL61),.BLN(BLN61),.WL(WL121));
sram_cell_6t_5 inst_cell_121_62 (.BL(BL62),.BLN(BLN62),.WL(WL121));
sram_cell_6t_5 inst_cell_121_63 (.BL(BL63),.BLN(BLN63),.WL(WL121));
sram_cell_6t_5 inst_cell_121_64 (.BL(BL64),.BLN(BLN64),.WL(WL121));
sram_cell_6t_5 inst_cell_121_65 (.BL(BL65),.BLN(BLN65),.WL(WL121));
sram_cell_6t_5 inst_cell_121_66 (.BL(BL66),.BLN(BLN66),.WL(WL121));
sram_cell_6t_5 inst_cell_121_67 (.BL(BL67),.BLN(BLN67),.WL(WL121));
sram_cell_6t_5 inst_cell_121_68 (.BL(BL68),.BLN(BLN68),.WL(WL121));
sram_cell_6t_5 inst_cell_121_69 (.BL(BL69),.BLN(BLN69),.WL(WL121));
sram_cell_6t_5 inst_cell_121_70 (.BL(BL70),.BLN(BLN70),.WL(WL121));
sram_cell_6t_5 inst_cell_121_71 (.BL(BL71),.BLN(BLN71),.WL(WL121));
sram_cell_6t_5 inst_cell_121_72 (.BL(BL72),.BLN(BLN72),.WL(WL121));
sram_cell_6t_5 inst_cell_121_73 (.BL(BL73),.BLN(BLN73),.WL(WL121));
sram_cell_6t_5 inst_cell_121_74 (.BL(BL74),.BLN(BLN74),.WL(WL121));
sram_cell_6t_5 inst_cell_121_75 (.BL(BL75),.BLN(BLN75),.WL(WL121));
sram_cell_6t_5 inst_cell_121_76 (.BL(BL76),.BLN(BLN76),.WL(WL121));
sram_cell_6t_5 inst_cell_121_77 (.BL(BL77),.BLN(BLN77),.WL(WL121));
sram_cell_6t_5 inst_cell_121_78 (.BL(BL78),.BLN(BLN78),.WL(WL121));
sram_cell_6t_5 inst_cell_121_79 (.BL(BL79),.BLN(BLN79),.WL(WL121));
sram_cell_6t_5 inst_cell_121_80 (.BL(BL80),.BLN(BLN80),.WL(WL121));
sram_cell_6t_5 inst_cell_121_81 (.BL(BL81),.BLN(BLN81),.WL(WL121));
sram_cell_6t_5 inst_cell_121_82 (.BL(BL82),.BLN(BLN82),.WL(WL121));
sram_cell_6t_5 inst_cell_121_83 (.BL(BL83),.BLN(BLN83),.WL(WL121));
sram_cell_6t_5 inst_cell_121_84 (.BL(BL84),.BLN(BLN84),.WL(WL121));
sram_cell_6t_5 inst_cell_121_85 (.BL(BL85),.BLN(BLN85),.WL(WL121));
sram_cell_6t_5 inst_cell_121_86 (.BL(BL86),.BLN(BLN86),.WL(WL121));
sram_cell_6t_5 inst_cell_121_87 (.BL(BL87),.BLN(BLN87),.WL(WL121));
sram_cell_6t_5 inst_cell_121_88 (.BL(BL88),.BLN(BLN88),.WL(WL121));
sram_cell_6t_5 inst_cell_121_89 (.BL(BL89),.BLN(BLN89),.WL(WL121));
sram_cell_6t_5 inst_cell_121_90 (.BL(BL90),.BLN(BLN90),.WL(WL121));
sram_cell_6t_5 inst_cell_121_91 (.BL(BL91),.BLN(BLN91),.WL(WL121));
sram_cell_6t_5 inst_cell_121_92 (.BL(BL92),.BLN(BLN92),.WL(WL121));
sram_cell_6t_5 inst_cell_121_93 (.BL(BL93),.BLN(BLN93),.WL(WL121));
sram_cell_6t_5 inst_cell_121_94 (.BL(BL94),.BLN(BLN94),.WL(WL121));
sram_cell_6t_5 inst_cell_121_95 (.BL(BL95),.BLN(BLN95),.WL(WL121));
sram_cell_6t_5 inst_cell_121_96 (.BL(BL96),.BLN(BLN96),.WL(WL121));
sram_cell_6t_5 inst_cell_121_97 (.BL(BL97),.BLN(BLN97),.WL(WL121));
sram_cell_6t_5 inst_cell_121_98 (.BL(BL98),.BLN(BLN98),.WL(WL121));
sram_cell_6t_5 inst_cell_121_99 (.BL(BL99),.BLN(BLN99),.WL(WL121));
sram_cell_6t_5 inst_cell_121_100 (.BL(BL100),.BLN(BLN100),.WL(WL121));
sram_cell_6t_5 inst_cell_121_101 (.BL(BL101),.BLN(BLN101),.WL(WL121));
sram_cell_6t_5 inst_cell_121_102 (.BL(BL102),.BLN(BLN102),.WL(WL121));
sram_cell_6t_5 inst_cell_121_103 (.BL(BL103),.BLN(BLN103),.WL(WL121));
sram_cell_6t_5 inst_cell_121_104 (.BL(BL104),.BLN(BLN104),.WL(WL121));
sram_cell_6t_5 inst_cell_121_105 (.BL(BL105),.BLN(BLN105),.WL(WL121));
sram_cell_6t_5 inst_cell_121_106 (.BL(BL106),.BLN(BLN106),.WL(WL121));
sram_cell_6t_5 inst_cell_121_107 (.BL(BL107),.BLN(BLN107),.WL(WL121));
sram_cell_6t_5 inst_cell_121_108 (.BL(BL108),.BLN(BLN108),.WL(WL121));
sram_cell_6t_5 inst_cell_121_109 (.BL(BL109),.BLN(BLN109),.WL(WL121));
sram_cell_6t_5 inst_cell_121_110 (.BL(BL110),.BLN(BLN110),.WL(WL121));
sram_cell_6t_5 inst_cell_121_111 (.BL(BL111),.BLN(BLN111),.WL(WL121));
sram_cell_6t_5 inst_cell_121_112 (.BL(BL112),.BLN(BLN112),.WL(WL121));
sram_cell_6t_5 inst_cell_121_113 (.BL(BL113),.BLN(BLN113),.WL(WL121));
sram_cell_6t_5 inst_cell_121_114 (.BL(BL114),.BLN(BLN114),.WL(WL121));
sram_cell_6t_5 inst_cell_121_115 (.BL(BL115),.BLN(BLN115),.WL(WL121));
sram_cell_6t_5 inst_cell_121_116 (.BL(BL116),.BLN(BLN116),.WL(WL121));
sram_cell_6t_5 inst_cell_121_117 (.BL(BL117),.BLN(BLN117),.WL(WL121));
sram_cell_6t_5 inst_cell_121_118 (.BL(BL118),.BLN(BLN118),.WL(WL121));
sram_cell_6t_5 inst_cell_121_119 (.BL(BL119),.BLN(BLN119),.WL(WL121));
sram_cell_6t_5 inst_cell_121_120 (.BL(BL120),.BLN(BLN120),.WL(WL121));
sram_cell_6t_5 inst_cell_121_121 (.BL(BL121),.BLN(BLN121),.WL(WL121));
sram_cell_6t_5 inst_cell_121_122 (.BL(BL122),.BLN(BLN122),.WL(WL121));
sram_cell_6t_5 inst_cell_121_123 (.BL(BL123),.BLN(BLN123),.WL(WL121));
sram_cell_6t_5 inst_cell_121_124 (.BL(BL124),.BLN(BLN124),.WL(WL121));
sram_cell_6t_5 inst_cell_121_125 (.BL(BL125),.BLN(BLN125),.WL(WL121));
sram_cell_6t_5 inst_cell_121_126 (.BL(BL126),.BLN(BLN126),.WL(WL121));
sram_cell_6t_5 inst_cell_121_127 (.BL(BL127),.BLN(BLN127),.WL(WL121));
sram_cell_6t_5 inst_cell_122_0 (.BL(BL0),.BLN(BLN0),.WL(WL122));
sram_cell_6t_5 inst_cell_122_1 (.BL(BL1),.BLN(BLN1),.WL(WL122));
sram_cell_6t_5 inst_cell_122_2 (.BL(BL2),.BLN(BLN2),.WL(WL122));
sram_cell_6t_5 inst_cell_122_3 (.BL(BL3),.BLN(BLN3),.WL(WL122));
sram_cell_6t_5 inst_cell_122_4 (.BL(BL4),.BLN(BLN4),.WL(WL122));
sram_cell_6t_5 inst_cell_122_5 (.BL(BL5),.BLN(BLN5),.WL(WL122));
sram_cell_6t_5 inst_cell_122_6 (.BL(BL6),.BLN(BLN6),.WL(WL122));
sram_cell_6t_5 inst_cell_122_7 (.BL(BL7),.BLN(BLN7),.WL(WL122));
sram_cell_6t_5 inst_cell_122_8 (.BL(BL8),.BLN(BLN8),.WL(WL122));
sram_cell_6t_5 inst_cell_122_9 (.BL(BL9),.BLN(BLN9),.WL(WL122));
sram_cell_6t_5 inst_cell_122_10 (.BL(BL10),.BLN(BLN10),.WL(WL122));
sram_cell_6t_5 inst_cell_122_11 (.BL(BL11),.BLN(BLN11),.WL(WL122));
sram_cell_6t_5 inst_cell_122_12 (.BL(BL12),.BLN(BLN12),.WL(WL122));
sram_cell_6t_5 inst_cell_122_13 (.BL(BL13),.BLN(BLN13),.WL(WL122));
sram_cell_6t_5 inst_cell_122_14 (.BL(BL14),.BLN(BLN14),.WL(WL122));
sram_cell_6t_5 inst_cell_122_15 (.BL(BL15),.BLN(BLN15),.WL(WL122));
sram_cell_6t_5 inst_cell_122_16 (.BL(BL16),.BLN(BLN16),.WL(WL122));
sram_cell_6t_5 inst_cell_122_17 (.BL(BL17),.BLN(BLN17),.WL(WL122));
sram_cell_6t_5 inst_cell_122_18 (.BL(BL18),.BLN(BLN18),.WL(WL122));
sram_cell_6t_5 inst_cell_122_19 (.BL(BL19),.BLN(BLN19),.WL(WL122));
sram_cell_6t_5 inst_cell_122_20 (.BL(BL20),.BLN(BLN20),.WL(WL122));
sram_cell_6t_5 inst_cell_122_21 (.BL(BL21),.BLN(BLN21),.WL(WL122));
sram_cell_6t_5 inst_cell_122_22 (.BL(BL22),.BLN(BLN22),.WL(WL122));
sram_cell_6t_5 inst_cell_122_23 (.BL(BL23),.BLN(BLN23),.WL(WL122));
sram_cell_6t_5 inst_cell_122_24 (.BL(BL24),.BLN(BLN24),.WL(WL122));
sram_cell_6t_5 inst_cell_122_25 (.BL(BL25),.BLN(BLN25),.WL(WL122));
sram_cell_6t_5 inst_cell_122_26 (.BL(BL26),.BLN(BLN26),.WL(WL122));
sram_cell_6t_5 inst_cell_122_27 (.BL(BL27),.BLN(BLN27),.WL(WL122));
sram_cell_6t_5 inst_cell_122_28 (.BL(BL28),.BLN(BLN28),.WL(WL122));
sram_cell_6t_5 inst_cell_122_29 (.BL(BL29),.BLN(BLN29),.WL(WL122));
sram_cell_6t_5 inst_cell_122_30 (.BL(BL30),.BLN(BLN30),.WL(WL122));
sram_cell_6t_5 inst_cell_122_31 (.BL(BL31),.BLN(BLN31),.WL(WL122));
sram_cell_6t_5 inst_cell_122_32 (.BL(BL32),.BLN(BLN32),.WL(WL122));
sram_cell_6t_5 inst_cell_122_33 (.BL(BL33),.BLN(BLN33),.WL(WL122));
sram_cell_6t_5 inst_cell_122_34 (.BL(BL34),.BLN(BLN34),.WL(WL122));
sram_cell_6t_5 inst_cell_122_35 (.BL(BL35),.BLN(BLN35),.WL(WL122));
sram_cell_6t_5 inst_cell_122_36 (.BL(BL36),.BLN(BLN36),.WL(WL122));
sram_cell_6t_5 inst_cell_122_37 (.BL(BL37),.BLN(BLN37),.WL(WL122));
sram_cell_6t_5 inst_cell_122_38 (.BL(BL38),.BLN(BLN38),.WL(WL122));
sram_cell_6t_5 inst_cell_122_39 (.BL(BL39),.BLN(BLN39),.WL(WL122));
sram_cell_6t_5 inst_cell_122_40 (.BL(BL40),.BLN(BLN40),.WL(WL122));
sram_cell_6t_5 inst_cell_122_41 (.BL(BL41),.BLN(BLN41),.WL(WL122));
sram_cell_6t_5 inst_cell_122_42 (.BL(BL42),.BLN(BLN42),.WL(WL122));
sram_cell_6t_5 inst_cell_122_43 (.BL(BL43),.BLN(BLN43),.WL(WL122));
sram_cell_6t_5 inst_cell_122_44 (.BL(BL44),.BLN(BLN44),.WL(WL122));
sram_cell_6t_5 inst_cell_122_45 (.BL(BL45),.BLN(BLN45),.WL(WL122));
sram_cell_6t_5 inst_cell_122_46 (.BL(BL46),.BLN(BLN46),.WL(WL122));
sram_cell_6t_5 inst_cell_122_47 (.BL(BL47),.BLN(BLN47),.WL(WL122));
sram_cell_6t_5 inst_cell_122_48 (.BL(BL48),.BLN(BLN48),.WL(WL122));
sram_cell_6t_5 inst_cell_122_49 (.BL(BL49),.BLN(BLN49),.WL(WL122));
sram_cell_6t_5 inst_cell_122_50 (.BL(BL50),.BLN(BLN50),.WL(WL122));
sram_cell_6t_5 inst_cell_122_51 (.BL(BL51),.BLN(BLN51),.WL(WL122));
sram_cell_6t_5 inst_cell_122_52 (.BL(BL52),.BLN(BLN52),.WL(WL122));
sram_cell_6t_5 inst_cell_122_53 (.BL(BL53),.BLN(BLN53),.WL(WL122));
sram_cell_6t_5 inst_cell_122_54 (.BL(BL54),.BLN(BLN54),.WL(WL122));
sram_cell_6t_5 inst_cell_122_55 (.BL(BL55),.BLN(BLN55),.WL(WL122));
sram_cell_6t_5 inst_cell_122_56 (.BL(BL56),.BLN(BLN56),.WL(WL122));
sram_cell_6t_5 inst_cell_122_57 (.BL(BL57),.BLN(BLN57),.WL(WL122));
sram_cell_6t_5 inst_cell_122_58 (.BL(BL58),.BLN(BLN58),.WL(WL122));
sram_cell_6t_5 inst_cell_122_59 (.BL(BL59),.BLN(BLN59),.WL(WL122));
sram_cell_6t_5 inst_cell_122_60 (.BL(BL60),.BLN(BLN60),.WL(WL122));
sram_cell_6t_5 inst_cell_122_61 (.BL(BL61),.BLN(BLN61),.WL(WL122));
sram_cell_6t_5 inst_cell_122_62 (.BL(BL62),.BLN(BLN62),.WL(WL122));
sram_cell_6t_5 inst_cell_122_63 (.BL(BL63),.BLN(BLN63),.WL(WL122));
sram_cell_6t_5 inst_cell_122_64 (.BL(BL64),.BLN(BLN64),.WL(WL122));
sram_cell_6t_5 inst_cell_122_65 (.BL(BL65),.BLN(BLN65),.WL(WL122));
sram_cell_6t_5 inst_cell_122_66 (.BL(BL66),.BLN(BLN66),.WL(WL122));
sram_cell_6t_5 inst_cell_122_67 (.BL(BL67),.BLN(BLN67),.WL(WL122));
sram_cell_6t_5 inst_cell_122_68 (.BL(BL68),.BLN(BLN68),.WL(WL122));
sram_cell_6t_5 inst_cell_122_69 (.BL(BL69),.BLN(BLN69),.WL(WL122));
sram_cell_6t_5 inst_cell_122_70 (.BL(BL70),.BLN(BLN70),.WL(WL122));
sram_cell_6t_5 inst_cell_122_71 (.BL(BL71),.BLN(BLN71),.WL(WL122));
sram_cell_6t_5 inst_cell_122_72 (.BL(BL72),.BLN(BLN72),.WL(WL122));
sram_cell_6t_5 inst_cell_122_73 (.BL(BL73),.BLN(BLN73),.WL(WL122));
sram_cell_6t_5 inst_cell_122_74 (.BL(BL74),.BLN(BLN74),.WL(WL122));
sram_cell_6t_5 inst_cell_122_75 (.BL(BL75),.BLN(BLN75),.WL(WL122));
sram_cell_6t_5 inst_cell_122_76 (.BL(BL76),.BLN(BLN76),.WL(WL122));
sram_cell_6t_5 inst_cell_122_77 (.BL(BL77),.BLN(BLN77),.WL(WL122));
sram_cell_6t_5 inst_cell_122_78 (.BL(BL78),.BLN(BLN78),.WL(WL122));
sram_cell_6t_5 inst_cell_122_79 (.BL(BL79),.BLN(BLN79),.WL(WL122));
sram_cell_6t_5 inst_cell_122_80 (.BL(BL80),.BLN(BLN80),.WL(WL122));
sram_cell_6t_5 inst_cell_122_81 (.BL(BL81),.BLN(BLN81),.WL(WL122));
sram_cell_6t_5 inst_cell_122_82 (.BL(BL82),.BLN(BLN82),.WL(WL122));
sram_cell_6t_5 inst_cell_122_83 (.BL(BL83),.BLN(BLN83),.WL(WL122));
sram_cell_6t_5 inst_cell_122_84 (.BL(BL84),.BLN(BLN84),.WL(WL122));
sram_cell_6t_5 inst_cell_122_85 (.BL(BL85),.BLN(BLN85),.WL(WL122));
sram_cell_6t_5 inst_cell_122_86 (.BL(BL86),.BLN(BLN86),.WL(WL122));
sram_cell_6t_5 inst_cell_122_87 (.BL(BL87),.BLN(BLN87),.WL(WL122));
sram_cell_6t_5 inst_cell_122_88 (.BL(BL88),.BLN(BLN88),.WL(WL122));
sram_cell_6t_5 inst_cell_122_89 (.BL(BL89),.BLN(BLN89),.WL(WL122));
sram_cell_6t_5 inst_cell_122_90 (.BL(BL90),.BLN(BLN90),.WL(WL122));
sram_cell_6t_5 inst_cell_122_91 (.BL(BL91),.BLN(BLN91),.WL(WL122));
sram_cell_6t_5 inst_cell_122_92 (.BL(BL92),.BLN(BLN92),.WL(WL122));
sram_cell_6t_5 inst_cell_122_93 (.BL(BL93),.BLN(BLN93),.WL(WL122));
sram_cell_6t_5 inst_cell_122_94 (.BL(BL94),.BLN(BLN94),.WL(WL122));
sram_cell_6t_5 inst_cell_122_95 (.BL(BL95),.BLN(BLN95),.WL(WL122));
sram_cell_6t_5 inst_cell_122_96 (.BL(BL96),.BLN(BLN96),.WL(WL122));
sram_cell_6t_5 inst_cell_122_97 (.BL(BL97),.BLN(BLN97),.WL(WL122));
sram_cell_6t_5 inst_cell_122_98 (.BL(BL98),.BLN(BLN98),.WL(WL122));
sram_cell_6t_5 inst_cell_122_99 (.BL(BL99),.BLN(BLN99),.WL(WL122));
sram_cell_6t_5 inst_cell_122_100 (.BL(BL100),.BLN(BLN100),.WL(WL122));
sram_cell_6t_5 inst_cell_122_101 (.BL(BL101),.BLN(BLN101),.WL(WL122));
sram_cell_6t_5 inst_cell_122_102 (.BL(BL102),.BLN(BLN102),.WL(WL122));
sram_cell_6t_5 inst_cell_122_103 (.BL(BL103),.BLN(BLN103),.WL(WL122));
sram_cell_6t_5 inst_cell_122_104 (.BL(BL104),.BLN(BLN104),.WL(WL122));
sram_cell_6t_5 inst_cell_122_105 (.BL(BL105),.BLN(BLN105),.WL(WL122));
sram_cell_6t_5 inst_cell_122_106 (.BL(BL106),.BLN(BLN106),.WL(WL122));
sram_cell_6t_5 inst_cell_122_107 (.BL(BL107),.BLN(BLN107),.WL(WL122));
sram_cell_6t_5 inst_cell_122_108 (.BL(BL108),.BLN(BLN108),.WL(WL122));
sram_cell_6t_5 inst_cell_122_109 (.BL(BL109),.BLN(BLN109),.WL(WL122));
sram_cell_6t_5 inst_cell_122_110 (.BL(BL110),.BLN(BLN110),.WL(WL122));
sram_cell_6t_5 inst_cell_122_111 (.BL(BL111),.BLN(BLN111),.WL(WL122));
sram_cell_6t_5 inst_cell_122_112 (.BL(BL112),.BLN(BLN112),.WL(WL122));
sram_cell_6t_5 inst_cell_122_113 (.BL(BL113),.BLN(BLN113),.WL(WL122));
sram_cell_6t_5 inst_cell_122_114 (.BL(BL114),.BLN(BLN114),.WL(WL122));
sram_cell_6t_5 inst_cell_122_115 (.BL(BL115),.BLN(BLN115),.WL(WL122));
sram_cell_6t_5 inst_cell_122_116 (.BL(BL116),.BLN(BLN116),.WL(WL122));
sram_cell_6t_5 inst_cell_122_117 (.BL(BL117),.BLN(BLN117),.WL(WL122));
sram_cell_6t_5 inst_cell_122_118 (.BL(BL118),.BLN(BLN118),.WL(WL122));
sram_cell_6t_5 inst_cell_122_119 (.BL(BL119),.BLN(BLN119),.WL(WL122));
sram_cell_6t_5 inst_cell_122_120 (.BL(BL120),.BLN(BLN120),.WL(WL122));
sram_cell_6t_5 inst_cell_122_121 (.BL(BL121),.BLN(BLN121),.WL(WL122));
sram_cell_6t_5 inst_cell_122_122 (.BL(BL122),.BLN(BLN122),.WL(WL122));
sram_cell_6t_5 inst_cell_122_123 (.BL(BL123),.BLN(BLN123),.WL(WL122));
sram_cell_6t_5 inst_cell_122_124 (.BL(BL124),.BLN(BLN124),.WL(WL122));
sram_cell_6t_5 inst_cell_122_125 (.BL(BL125),.BLN(BLN125),.WL(WL122));
sram_cell_6t_5 inst_cell_122_126 (.BL(BL126),.BLN(BLN126),.WL(WL122));
sram_cell_6t_5 inst_cell_122_127 (.BL(BL127),.BLN(BLN127),.WL(WL122));
sram_cell_6t_5 inst_cell_123_0 (.BL(BL0),.BLN(BLN0),.WL(WL123));
sram_cell_6t_5 inst_cell_123_1 (.BL(BL1),.BLN(BLN1),.WL(WL123));
sram_cell_6t_5 inst_cell_123_2 (.BL(BL2),.BLN(BLN2),.WL(WL123));
sram_cell_6t_5 inst_cell_123_3 (.BL(BL3),.BLN(BLN3),.WL(WL123));
sram_cell_6t_5 inst_cell_123_4 (.BL(BL4),.BLN(BLN4),.WL(WL123));
sram_cell_6t_5 inst_cell_123_5 (.BL(BL5),.BLN(BLN5),.WL(WL123));
sram_cell_6t_5 inst_cell_123_6 (.BL(BL6),.BLN(BLN6),.WL(WL123));
sram_cell_6t_5 inst_cell_123_7 (.BL(BL7),.BLN(BLN7),.WL(WL123));
sram_cell_6t_5 inst_cell_123_8 (.BL(BL8),.BLN(BLN8),.WL(WL123));
sram_cell_6t_5 inst_cell_123_9 (.BL(BL9),.BLN(BLN9),.WL(WL123));
sram_cell_6t_5 inst_cell_123_10 (.BL(BL10),.BLN(BLN10),.WL(WL123));
sram_cell_6t_5 inst_cell_123_11 (.BL(BL11),.BLN(BLN11),.WL(WL123));
sram_cell_6t_5 inst_cell_123_12 (.BL(BL12),.BLN(BLN12),.WL(WL123));
sram_cell_6t_5 inst_cell_123_13 (.BL(BL13),.BLN(BLN13),.WL(WL123));
sram_cell_6t_5 inst_cell_123_14 (.BL(BL14),.BLN(BLN14),.WL(WL123));
sram_cell_6t_5 inst_cell_123_15 (.BL(BL15),.BLN(BLN15),.WL(WL123));
sram_cell_6t_5 inst_cell_123_16 (.BL(BL16),.BLN(BLN16),.WL(WL123));
sram_cell_6t_5 inst_cell_123_17 (.BL(BL17),.BLN(BLN17),.WL(WL123));
sram_cell_6t_5 inst_cell_123_18 (.BL(BL18),.BLN(BLN18),.WL(WL123));
sram_cell_6t_5 inst_cell_123_19 (.BL(BL19),.BLN(BLN19),.WL(WL123));
sram_cell_6t_5 inst_cell_123_20 (.BL(BL20),.BLN(BLN20),.WL(WL123));
sram_cell_6t_5 inst_cell_123_21 (.BL(BL21),.BLN(BLN21),.WL(WL123));
sram_cell_6t_5 inst_cell_123_22 (.BL(BL22),.BLN(BLN22),.WL(WL123));
sram_cell_6t_5 inst_cell_123_23 (.BL(BL23),.BLN(BLN23),.WL(WL123));
sram_cell_6t_5 inst_cell_123_24 (.BL(BL24),.BLN(BLN24),.WL(WL123));
sram_cell_6t_5 inst_cell_123_25 (.BL(BL25),.BLN(BLN25),.WL(WL123));
sram_cell_6t_5 inst_cell_123_26 (.BL(BL26),.BLN(BLN26),.WL(WL123));
sram_cell_6t_5 inst_cell_123_27 (.BL(BL27),.BLN(BLN27),.WL(WL123));
sram_cell_6t_5 inst_cell_123_28 (.BL(BL28),.BLN(BLN28),.WL(WL123));
sram_cell_6t_5 inst_cell_123_29 (.BL(BL29),.BLN(BLN29),.WL(WL123));
sram_cell_6t_5 inst_cell_123_30 (.BL(BL30),.BLN(BLN30),.WL(WL123));
sram_cell_6t_5 inst_cell_123_31 (.BL(BL31),.BLN(BLN31),.WL(WL123));
sram_cell_6t_5 inst_cell_123_32 (.BL(BL32),.BLN(BLN32),.WL(WL123));
sram_cell_6t_5 inst_cell_123_33 (.BL(BL33),.BLN(BLN33),.WL(WL123));
sram_cell_6t_5 inst_cell_123_34 (.BL(BL34),.BLN(BLN34),.WL(WL123));
sram_cell_6t_5 inst_cell_123_35 (.BL(BL35),.BLN(BLN35),.WL(WL123));
sram_cell_6t_5 inst_cell_123_36 (.BL(BL36),.BLN(BLN36),.WL(WL123));
sram_cell_6t_5 inst_cell_123_37 (.BL(BL37),.BLN(BLN37),.WL(WL123));
sram_cell_6t_5 inst_cell_123_38 (.BL(BL38),.BLN(BLN38),.WL(WL123));
sram_cell_6t_5 inst_cell_123_39 (.BL(BL39),.BLN(BLN39),.WL(WL123));
sram_cell_6t_5 inst_cell_123_40 (.BL(BL40),.BLN(BLN40),.WL(WL123));
sram_cell_6t_5 inst_cell_123_41 (.BL(BL41),.BLN(BLN41),.WL(WL123));
sram_cell_6t_5 inst_cell_123_42 (.BL(BL42),.BLN(BLN42),.WL(WL123));
sram_cell_6t_5 inst_cell_123_43 (.BL(BL43),.BLN(BLN43),.WL(WL123));
sram_cell_6t_5 inst_cell_123_44 (.BL(BL44),.BLN(BLN44),.WL(WL123));
sram_cell_6t_5 inst_cell_123_45 (.BL(BL45),.BLN(BLN45),.WL(WL123));
sram_cell_6t_5 inst_cell_123_46 (.BL(BL46),.BLN(BLN46),.WL(WL123));
sram_cell_6t_5 inst_cell_123_47 (.BL(BL47),.BLN(BLN47),.WL(WL123));
sram_cell_6t_5 inst_cell_123_48 (.BL(BL48),.BLN(BLN48),.WL(WL123));
sram_cell_6t_5 inst_cell_123_49 (.BL(BL49),.BLN(BLN49),.WL(WL123));
sram_cell_6t_5 inst_cell_123_50 (.BL(BL50),.BLN(BLN50),.WL(WL123));
sram_cell_6t_5 inst_cell_123_51 (.BL(BL51),.BLN(BLN51),.WL(WL123));
sram_cell_6t_5 inst_cell_123_52 (.BL(BL52),.BLN(BLN52),.WL(WL123));
sram_cell_6t_5 inst_cell_123_53 (.BL(BL53),.BLN(BLN53),.WL(WL123));
sram_cell_6t_5 inst_cell_123_54 (.BL(BL54),.BLN(BLN54),.WL(WL123));
sram_cell_6t_5 inst_cell_123_55 (.BL(BL55),.BLN(BLN55),.WL(WL123));
sram_cell_6t_5 inst_cell_123_56 (.BL(BL56),.BLN(BLN56),.WL(WL123));
sram_cell_6t_5 inst_cell_123_57 (.BL(BL57),.BLN(BLN57),.WL(WL123));
sram_cell_6t_5 inst_cell_123_58 (.BL(BL58),.BLN(BLN58),.WL(WL123));
sram_cell_6t_5 inst_cell_123_59 (.BL(BL59),.BLN(BLN59),.WL(WL123));
sram_cell_6t_5 inst_cell_123_60 (.BL(BL60),.BLN(BLN60),.WL(WL123));
sram_cell_6t_5 inst_cell_123_61 (.BL(BL61),.BLN(BLN61),.WL(WL123));
sram_cell_6t_5 inst_cell_123_62 (.BL(BL62),.BLN(BLN62),.WL(WL123));
sram_cell_6t_5 inst_cell_123_63 (.BL(BL63),.BLN(BLN63),.WL(WL123));
sram_cell_6t_5 inst_cell_123_64 (.BL(BL64),.BLN(BLN64),.WL(WL123));
sram_cell_6t_5 inst_cell_123_65 (.BL(BL65),.BLN(BLN65),.WL(WL123));
sram_cell_6t_5 inst_cell_123_66 (.BL(BL66),.BLN(BLN66),.WL(WL123));
sram_cell_6t_5 inst_cell_123_67 (.BL(BL67),.BLN(BLN67),.WL(WL123));
sram_cell_6t_5 inst_cell_123_68 (.BL(BL68),.BLN(BLN68),.WL(WL123));
sram_cell_6t_5 inst_cell_123_69 (.BL(BL69),.BLN(BLN69),.WL(WL123));
sram_cell_6t_5 inst_cell_123_70 (.BL(BL70),.BLN(BLN70),.WL(WL123));
sram_cell_6t_5 inst_cell_123_71 (.BL(BL71),.BLN(BLN71),.WL(WL123));
sram_cell_6t_5 inst_cell_123_72 (.BL(BL72),.BLN(BLN72),.WL(WL123));
sram_cell_6t_5 inst_cell_123_73 (.BL(BL73),.BLN(BLN73),.WL(WL123));
sram_cell_6t_5 inst_cell_123_74 (.BL(BL74),.BLN(BLN74),.WL(WL123));
sram_cell_6t_5 inst_cell_123_75 (.BL(BL75),.BLN(BLN75),.WL(WL123));
sram_cell_6t_5 inst_cell_123_76 (.BL(BL76),.BLN(BLN76),.WL(WL123));
sram_cell_6t_5 inst_cell_123_77 (.BL(BL77),.BLN(BLN77),.WL(WL123));
sram_cell_6t_5 inst_cell_123_78 (.BL(BL78),.BLN(BLN78),.WL(WL123));
sram_cell_6t_5 inst_cell_123_79 (.BL(BL79),.BLN(BLN79),.WL(WL123));
sram_cell_6t_5 inst_cell_123_80 (.BL(BL80),.BLN(BLN80),.WL(WL123));
sram_cell_6t_5 inst_cell_123_81 (.BL(BL81),.BLN(BLN81),.WL(WL123));
sram_cell_6t_5 inst_cell_123_82 (.BL(BL82),.BLN(BLN82),.WL(WL123));
sram_cell_6t_5 inst_cell_123_83 (.BL(BL83),.BLN(BLN83),.WL(WL123));
sram_cell_6t_5 inst_cell_123_84 (.BL(BL84),.BLN(BLN84),.WL(WL123));
sram_cell_6t_5 inst_cell_123_85 (.BL(BL85),.BLN(BLN85),.WL(WL123));
sram_cell_6t_5 inst_cell_123_86 (.BL(BL86),.BLN(BLN86),.WL(WL123));
sram_cell_6t_5 inst_cell_123_87 (.BL(BL87),.BLN(BLN87),.WL(WL123));
sram_cell_6t_5 inst_cell_123_88 (.BL(BL88),.BLN(BLN88),.WL(WL123));
sram_cell_6t_5 inst_cell_123_89 (.BL(BL89),.BLN(BLN89),.WL(WL123));
sram_cell_6t_5 inst_cell_123_90 (.BL(BL90),.BLN(BLN90),.WL(WL123));
sram_cell_6t_5 inst_cell_123_91 (.BL(BL91),.BLN(BLN91),.WL(WL123));
sram_cell_6t_5 inst_cell_123_92 (.BL(BL92),.BLN(BLN92),.WL(WL123));
sram_cell_6t_5 inst_cell_123_93 (.BL(BL93),.BLN(BLN93),.WL(WL123));
sram_cell_6t_5 inst_cell_123_94 (.BL(BL94),.BLN(BLN94),.WL(WL123));
sram_cell_6t_5 inst_cell_123_95 (.BL(BL95),.BLN(BLN95),.WL(WL123));
sram_cell_6t_5 inst_cell_123_96 (.BL(BL96),.BLN(BLN96),.WL(WL123));
sram_cell_6t_5 inst_cell_123_97 (.BL(BL97),.BLN(BLN97),.WL(WL123));
sram_cell_6t_5 inst_cell_123_98 (.BL(BL98),.BLN(BLN98),.WL(WL123));
sram_cell_6t_5 inst_cell_123_99 (.BL(BL99),.BLN(BLN99),.WL(WL123));
sram_cell_6t_5 inst_cell_123_100 (.BL(BL100),.BLN(BLN100),.WL(WL123));
sram_cell_6t_5 inst_cell_123_101 (.BL(BL101),.BLN(BLN101),.WL(WL123));
sram_cell_6t_5 inst_cell_123_102 (.BL(BL102),.BLN(BLN102),.WL(WL123));
sram_cell_6t_5 inst_cell_123_103 (.BL(BL103),.BLN(BLN103),.WL(WL123));
sram_cell_6t_5 inst_cell_123_104 (.BL(BL104),.BLN(BLN104),.WL(WL123));
sram_cell_6t_5 inst_cell_123_105 (.BL(BL105),.BLN(BLN105),.WL(WL123));
sram_cell_6t_5 inst_cell_123_106 (.BL(BL106),.BLN(BLN106),.WL(WL123));
sram_cell_6t_5 inst_cell_123_107 (.BL(BL107),.BLN(BLN107),.WL(WL123));
sram_cell_6t_5 inst_cell_123_108 (.BL(BL108),.BLN(BLN108),.WL(WL123));
sram_cell_6t_5 inst_cell_123_109 (.BL(BL109),.BLN(BLN109),.WL(WL123));
sram_cell_6t_5 inst_cell_123_110 (.BL(BL110),.BLN(BLN110),.WL(WL123));
sram_cell_6t_5 inst_cell_123_111 (.BL(BL111),.BLN(BLN111),.WL(WL123));
sram_cell_6t_5 inst_cell_123_112 (.BL(BL112),.BLN(BLN112),.WL(WL123));
sram_cell_6t_5 inst_cell_123_113 (.BL(BL113),.BLN(BLN113),.WL(WL123));
sram_cell_6t_5 inst_cell_123_114 (.BL(BL114),.BLN(BLN114),.WL(WL123));
sram_cell_6t_5 inst_cell_123_115 (.BL(BL115),.BLN(BLN115),.WL(WL123));
sram_cell_6t_5 inst_cell_123_116 (.BL(BL116),.BLN(BLN116),.WL(WL123));
sram_cell_6t_5 inst_cell_123_117 (.BL(BL117),.BLN(BLN117),.WL(WL123));
sram_cell_6t_5 inst_cell_123_118 (.BL(BL118),.BLN(BLN118),.WL(WL123));
sram_cell_6t_5 inst_cell_123_119 (.BL(BL119),.BLN(BLN119),.WL(WL123));
sram_cell_6t_5 inst_cell_123_120 (.BL(BL120),.BLN(BLN120),.WL(WL123));
sram_cell_6t_5 inst_cell_123_121 (.BL(BL121),.BLN(BLN121),.WL(WL123));
sram_cell_6t_5 inst_cell_123_122 (.BL(BL122),.BLN(BLN122),.WL(WL123));
sram_cell_6t_5 inst_cell_123_123 (.BL(BL123),.BLN(BLN123),.WL(WL123));
sram_cell_6t_5 inst_cell_123_124 (.BL(BL124),.BLN(BLN124),.WL(WL123));
sram_cell_6t_5 inst_cell_123_125 (.BL(BL125),.BLN(BLN125),.WL(WL123));
sram_cell_6t_5 inst_cell_123_126 (.BL(BL126),.BLN(BLN126),.WL(WL123));
sram_cell_6t_5 inst_cell_123_127 (.BL(BL127),.BLN(BLN127),.WL(WL123));
sram_cell_6t_5 inst_cell_124_0 (.BL(BL0),.BLN(BLN0),.WL(WL124));
sram_cell_6t_5 inst_cell_124_1 (.BL(BL1),.BLN(BLN1),.WL(WL124));
sram_cell_6t_5 inst_cell_124_2 (.BL(BL2),.BLN(BLN2),.WL(WL124));
sram_cell_6t_5 inst_cell_124_3 (.BL(BL3),.BLN(BLN3),.WL(WL124));
sram_cell_6t_5 inst_cell_124_4 (.BL(BL4),.BLN(BLN4),.WL(WL124));
sram_cell_6t_5 inst_cell_124_5 (.BL(BL5),.BLN(BLN5),.WL(WL124));
sram_cell_6t_5 inst_cell_124_6 (.BL(BL6),.BLN(BLN6),.WL(WL124));
sram_cell_6t_5 inst_cell_124_7 (.BL(BL7),.BLN(BLN7),.WL(WL124));
sram_cell_6t_5 inst_cell_124_8 (.BL(BL8),.BLN(BLN8),.WL(WL124));
sram_cell_6t_5 inst_cell_124_9 (.BL(BL9),.BLN(BLN9),.WL(WL124));
sram_cell_6t_5 inst_cell_124_10 (.BL(BL10),.BLN(BLN10),.WL(WL124));
sram_cell_6t_5 inst_cell_124_11 (.BL(BL11),.BLN(BLN11),.WL(WL124));
sram_cell_6t_5 inst_cell_124_12 (.BL(BL12),.BLN(BLN12),.WL(WL124));
sram_cell_6t_5 inst_cell_124_13 (.BL(BL13),.BLN(BLN13),.WL(WL124));
sram_cell_6t_5 inst_cell_124_14 (.BL(BL14),.BLN(BLN14),.WL(WL124));
sram_cell_6t_5 inst_cell_124_15 (.BL(BL15),.BLN(BLN15),.WL(WL124));
sram_cell_6t_5 inst_cell_124_16 (.BL(BL16),.BLN(BLN16),.WL(WL124));
sram_cell_6t_5 inst_cell_124_17 (.BL(BL17),.BLN(BLN17),.WL(WL124));
sram_cell_6t_5 inst_cell_124_18 (.BL(BL18),.BLN(BLN18),.WL(WL124));
sram_cell_6t_5 inst_cell_124_19 (.BL(BL19),.BLN(BLN19),.WL(WL124));
sram_cell_6t_5 inst_cell_124_20 (.BL(BL20),.BLN(BLN20),.WL(WL124));
sram_cell_6t_5 inst_cell_124_21 (.BL(BL21),.BLN(BLN21),.WL(WL124));
sram_cell_6t_5 inst_cell_124_22 (.BL(BL22),.BLN(BLN22),.WL(WL124));
sram_cell_6t_5 inst_cell_124_23 (.BL(BL23),.BLN(BLN23),.WL(WL124));
sram_cell_6t_5 inst_cell_124_24 (.BL(BL24),.BLN(BLN24),.WL(WL124));
sram_cell_6t_5 inst_cell_124_25 (.BL(BL25),.BLN(BLN25),.WL(WL124));
sram_cell_6t_5 inst_cell_124_26 (.BL(BL26),.BLN(BLN26),.WL(WL124));
sram_cell_6t_5 inst_cell_124_27 (.BL(BL27),.BLN(BLN27),.WL(WL124));
sram_cell_6t_5 inst_cell_124_28 (.BL(BL28),.BLN(BLN28),.WL(WL124));
sram_cell_6t_5 inst_cell_124_29 (.BL(BL29),.BLN(BLN29),.WL(WL124));
sram_cell_6t_5 inst_cell_124_30 (.BL(BL30),.BLN(BLN30),.WL(WL124));
sram_cell_6t_5 inst_cell_124_31 (.BL(BL31),.BLN(BLN31),.WL(WL124));
sram_cell_6t_5 inst_cell_124_32 (.BL(BL32),.BLN(BLN32),.WL(WL124));
sram_cell_6t_5 inst_cell_124_33 (.BL(BL33),.BLN(BLN33),.WL(WL124));
sram_cell_6t_5 inst_cell_124_34 (.BL(BL34),.BLN(BLN34),.WL(WL124));
sram_cell_6t_5 inst_cell_124_35 (.BL(BL35),.BLN(BLN35),.WL(WL124));
sram_cell_6t_5 inst_cell_124_36 (.BL(BL36),.BLN(BLN36),.WL(WL124));
sram_cell_6t_5 inst_cell_124_37 (.BL(BL37),.BLN(BLN37),.WL(WL124));
sram_cell_6t_5 inst_cell_124_38 (.BL(BL38),.BLN(BLN38),.WL(WL124));
sram_cell_6t_5 inst_cell_124_39 (.BL(BL39),.BLN(BLN39),.WL(WL124));
sram_cell_6t_5 inst_cell_124_40 (.BL(BL40),.BLN(BLN40),.WL(WL124));
sram_cell_6t_5 inst_cell_124_41 (.BL(BL41),.BLN(BLN41),.WL(WL124));
sram_cell_6t_5 inst_cell_124_42 (.BL(BL42),.BLN(BLN42),.WL(WL124));
sram_cell_6t_5 inst_cell_124_43 (.BL(BL43),.BLN(BLN43),.WL(WL124));
sram_cell_6t_5 inst_cell_124_44 (.BL(BL44),.BLN(BLN44),.WL(WL124));
sram_cell_6t_5 inst_cell_124_45 (.BL(BL45),.BLN(BLN45),.WL(WL124));
sram_cell_6t_5 inst_cell_124_46 (.BL(BL46),.BLN(BLN46),.WL(WL124));
sram_cell_6t_5 inst_cell_124_47 (.BL(BL47),.BLN(BLN47),.WL(WL124));
sram_cell_6t_5 inst_cell_124_48 (.BL(BL48),.BLN(BLN48),.WL(WL124));
sram_cell_6t_5 inst_cell_124_49 (.BL(BL49),.BLN(BLN49),.WL(WL124));
sram_cell_6t_5 inst_cell_124_50 (.BL(BL50),.BLN(BLN50),.WL(WL124));
sram_cell_6t_5 inst_cell_124_51 (.BL(BL51),.BLN(BLN51),.WL(WL124));
sram_cell_6t_5 inst_cell_124_52 (.BL(BL52),.BLN(BLN52),.WL(WL124));
sram_cell_6t_5 inst_cell_124_53 (.BL(BL53),.BLN(BLN53),.WL(WL124));
sram_cell_6t_5 inst_cell_124_54 (.BL(BL54),.BLN(BLN54),.WL(WL124));
sram_cell_6t_5 inst_cell_124_55 (.BL(BL55),.BLN(BLN55),.WL(WL124));
sram_cell_6t_5 inst_cell_124_56 (.BL(BL56),.BLN(BLN56),.WL(WL124));
sram_cell_6t_5 inst_cell_124_57 (.BL(BL57),.BLN(BLN57),.WL(WL124));
sram_cell_6t_5 inst_cell_124_58 (.BL(BL58),.BLN(BLN58),.WL(WL124));
sram_cell_6t_5 inst_cell_124_59 (.BL(BL59),.BLN(BLN59),.WL(WL124));
sram_cell_6t_5 inst_cell_124_60 (.BL(BL60),.BLN(BLN60),.WL(WL124));
sram_cell_6t_5 inst_cell_124_61 (.BL(BL61),.BLN(BLN61),.WL(WL124));
sram_cell_6t_5 inst_cell_124_62 (.BL(BL62),.BLN(BLN62),.WL(WL124));
sram_cell_6t_5 inst_cell_124_63 (.BL(BL63),.BLN(BLN63),.WL(WL124));
sram_cell_6t_5 inst_cell_124_64 (.BL(BL64),.BLN(BLN64),.WL(WL124));
sram_cell_6t_5 inst_cell_124_65 (.BL(BL65),.BLN(BLN65),.WL(WL124));
sram_cell_6t_5 inst_cell_124_66 (.BL(BL66),.BLN(BLN66),.WL(WL124));
sram_cell_6t_5 inst_cell_124_67 (.BL(BL67),.BLN(BLN67),.WL(WL124));
sram_cell_6t_5 inst_cell_124_68 (.BL(BL68),.BLN(BLN68),.WL(WL124));
sram_cell_6t_5 inst_cell_124_69 (.BL(BL69),.BLN(BLN69),.WL(WL124));
sram_cell_6t_5 inst_cell_124_70 (.BL(BL70),.BLN(BLN70),.WL(WL124));
sram_cell_6t_5 inst_cell_124_71 (.BL(BL71),.BLN(BLN71),.WL(WL124));
sram_cell_6t_5 inst_cell_124_72 (.BL(BL72),.BLN(BLN72),.WL(WL124));
sram_cell_6t_5 inst_cell_124_73 (.BL(BL73),.BLN(BLN73),.WL(WL124));
sram_cell_6t_5 inst_cell_124_74 (.BL(BL74),.BLN(BLN74),.WL(WL124));
sram_cell_6t_5 inst_cell_124_75 (.BL(BL75),.BLN(BLN75),.WL(WL124));
sram_cell_6t_5 inst_cell_124_76 (.BL(BL76),.BLN(BLN76),.WL(WL124));
sram_cell_6t_5 inst_cell_124_77 (.BL(BL77),.BLN(BLN77),.WL(WL124));
sram_cell_6t_5 inst_cell_124_78 (.BL(BL78),.BLN(BLN78),.WL(WL124));
sram_cell_6t_5 inst_cell_124_79 (.BL(BL79),.BLN(BLN79),.WL(WL124));
sram_cell_6t_5 inst_cell_124_80 (.BL(BL80),.BLN(BLN80),.WL(WL124));
sram_cell_6t_5 inst_cell_124_81 (.BL(BL81),.BLN(BLN81),.WL(WL124));
sram_cell_6t_5 inst_cell_124_82 (.BL(BL82),.BLN(BLN82),.WL(WL124));
sram_cell_6t_5 inst_cell_124_83 (.BL(BL83),.BLN(BLN83),.WL(WL124));
sram_cell_6t_5 inst_cell_124_84 (.BL(BL84),.BLN(BLN84),.WL(WL124));
sram_cell_6t_5 inst_cell_124_85 (.BL(BL85),.BLN(BLN85),.WL(WL124));
sram_cell_6t_5 inst_cell_124_86 (.BL(BL86),.BLN(BLN86),.WL(WL124));
sram_cell_6t_5 inst_cell_124_87 (.BL(BL87),.BLN(BLN87),.WL(WL124));
sram_cell_6t_5 inst_cell_124_88 (.BL(BL88),.BLN(BLN88),.WL(WL124));
sram_cell_6t_5 inst_cell_124_89 (.BL(BL89),.BLN(BLN89),.WL(WL124));
sram_cell_6t_5 inst_cell_124_90 (.BL(BL90),.BLN(BLN90),.WL(WL124));
sram_cell_6t_5 inst_cell_124_91 (.BL(BL91),.BLN(BLN91),.WL(WL124));
sram_cell_6t_5 inst_cell_124_92 (.BL(BL92),.BLN(BLN92),.WL(WL124));
sram_cell_6t_5 inst_cell_124_93 (.BL(BL93),.BLN(BLN93),.WL(WL124));
sram_cell_6t_5 inst_cell_124_94 (.BL(BL94),.BLN(BLN94),.WL(WL124));
sram_cell_6t_5 inst_cell_124_95 (.BL(BL95),.BLN(BLN95),.WL(WL124));
sram_cell_6t_5 inst_cell_124_96 (.BL(BL96),.BLN(BLN96),.WL(WL124));
sram_cell_6t_5 inst_cell_124_97 (.BL(BL97),.BLN(BLN97),.WL(WL124));
sram_cell_6t_5 inst_cell_124_98 (.BL(BL98),.BLN(BLN98),.WL(WL124));
sram_cell_6t_5 inst_cell_124_99 (.BL(BL99),.BLN(BLN99),.WL(WL124));
sram_cell_6t_5 inst_cell_124_100 (.BL(BL100),.BLN(BLN100),.WL(WL124));
sram_cell_6t_5 inst_cell_124_101 (.BL(BL101),.BLN(BLN101),.WL(WL124));
sram_cell_6t_5 inst_cell_124_102 (.BL(BL102),.BLN(BLN102),.WL(WL124));
sram_cell_6t_5 inst_cell_124_103 (.BL(BL103),.BLN(BLN103),.WL(WL124));
sram_cell_6t_5 inst_cell_124_104 (.BL(BL104),.BLN(BLN104),.WL(WL124));
sram_cell_6t_5 inst_cell_124_105 (.BL(BL105),.BLN(BLN105),.WL(WL124));
sram_cell_6t_5 inst_cell_124_106 (.BL(BL106),.BLN(BLN106),.WL(WL124));
sram_cell_6t_5 inst_cell_124_107 (.BL(BL107),.BLN(BLN107),.WL(WL124));
sram_cell_6t_5 inst_cell_124_108 (.BL(BL108),.BLN(BLN108),.WL(WL124));
sram_cell_6t_5 inst_cell_124_109 (.BL(BL109),.BLN(BLN109),.WL(WL124));
sram_cell_6t_5 inst_cell_124_110 (.BL(BL110),.BLN(BLN110),.WL(WL124));
sram_cell_6t_5 inst_cell_124_111 (.BL(BL111),.BLN(BLN111),.WL(WL124));
sram_cell_6t_5 inst_cell_124_112 (.BL(BL112),.BLN(BLN112),.WL(WL124));
sram_cell_6t_5 inst_cell_124_113 (.BL(BL113),.BLN(BLN113),.WL(WL124));
sram_cell_6t_5 inst_cell_124_114 (.BL(BL114),.BLN(BLN114),.WL(WL124));
sram_cell_6t_5 inst_cell_124_115 (.BL(BL115),.BLN(BLN115),.WL(WL124));
sram_cell_6t_5 inst_cell_124_116 (.BL(BL116),.BLN(BLN116),.WL(WL124));
sram_cell_6t_5 inst_cell_124_117 (.BL(BL117),.BLN(BLN117),.WL(WL124));
sram_cell_6t_5 inst_cell_124_118 (.BL(BL118),.BLN(BLN118),.WL(WL124));
sram_cell_6t_5 inst_cell_124_119 (.BL(BL119),.BLN(BLN119),.WL(WL124));
sram_cell_6t_5 inst_cell_124_120 (.BL(BL120),.BLN(BLN120),.WL(WL124));
sram_cell_6t_5 inst_cell_124_121 (.BL(BL121),.BLN(BLN121),.WL(WL124));
sram_cell_6t_5 inst_cell_124_122 (.BL(BL122),.BLN(BLN122),.WL(WL124));
sram_cell_6t_5 inst_cell_124_123 (.BL(BL123),.BLN(BLN123),.WL(WL124));
sram_cell_6t_5 inst_cell_124_124 (.BL(BL124),.BLN(BLN124),.WL(WL124));
sram_cell_6t_5 inst_cell_124_125 (.BL(BL125),.BLN(BLN125),.WL(WL124));
sram_cell_6t_5 inst_cell_124_126 (.BL(BL126),.BLN(BLN126),.WL(WL124));
sram_cell_6t_5 inst_cell_124_127 (.BL(BL127),.BLN(BLN127),.WL(WL124));
sram_cell_6t_5 inst_cell_125_0 (.BL(BL0),.BLN(BLN0),.WL(WL125));
sram_cell_6t_5 inst_cell_125_1 (.BL(BL1),.BLN(BLN1),.WL(WL125));
sram_cell_6t_5 inst_cell_125_2 (.BL(BL2),.BLN(BLN2),.WL(WL125));
sram_cell_6t_5 inst_cell_125_3 (.BL(BL3),.BLN(BLN3),.WL(WL125));
sram_cell_6t_5 inst_cell_125_4 (.BL(BL4),.BLN(BLN4),.WL(WL125));
sram_cell_6t_5 inst_cell_125_5 (.BL(BL5),.BLN(BLN5),.WL(WL125));
sram_cell_6t_5 inst_cell_125_6 (.BL(BL6),.BLN(BLN6),.WL(WL125));
sram_cell_6t_5 inst_cell_125_7 (.BL(BL7),.BLN(BLN7),.WL(WL125));
sram_cell_6t_5 inst_cell_125_8 (.BL(BL8),.BLN(BLN8),.WL(WL125));
sram_cell_6t_5 inst_cell_125_9 (.BL(BL9),.BLN(BLN9),.WL(WL125));
sram_cell_6t_5 inst_cell_125_10 (.BL(BL10),.BLN(BLN10),.WL(WL125));
sram_cell_6t_5 inst_cell_125_11 (.BL(BL11),.BLN(BLN11),.WL(WL125));
sram_cell_6t_5 inst_cell_125_12 (.BL(BL12),.BLN(BLN12),.WL(WL125));
sram_cell_6t_5 inst_cell_125_13 (.BL(BL13),.BLN(BLN13),.WL(WL125));
sram_cell_6t_5 inst_cell_125_14 (.BL(BL14),.BLN(BLN14),.WL(WL125));
sram_cell_6t_5 inst_cell_125_15 (.BL(BL15),.BLN(BLN15),.WL(WL125));
sram_cell_6t_5 inst_cell_125_16 (.BL(BL16),.BLN(BLN16),.WL(WL125));
sram_cell_6t_5 inst_cell_125_17 (.BL(BL17),.BLN(BLN17),.WL(WL125));
sram_cell_6t_5 inst_cell_125_18 (.BL(BL18),.BLN(BLN18),.WL(WL125));
sram_cell_6t_5 inst_cell_125_19 (.BL(BL19),.BLN(BLN19),.WL(WL125));
sram_cell_6t_5 inst_cell_125_20 (.BL(BL20),.BLN(BLN20),.WL(WL125));
sram_cell_6t_5 inst_cell_125_21 (.BL(BL21),.BLN(BLN21),.WL(WL125));
sram_cell_6t_5 inst_cell_125_22 (.BL(BL22),.BLN(BLN22),.WL(WL125));
sram_cell_6t_5 inst_cell_125_23 (.BL(BL23),.BLN(BLN23),.WL(WL125));
sram_cell_6t_5 inst_cell_125_24 (.BL(BL24),.BLN(BLN24),.WL(WL125));
sram_cell_6t_5 inst_cell_125_25 (.BL(BL25),.BLN(BLN25),.WL(WL125));
sram_cell_6t_5 inst_cell_125_26 (.BL(BL26),.BLN(BLN26),.WL(WL125));
sram_cell_6t_5 inst_cell_125_27 (.BL(BL27),.BLN(BLN27),.WL(WL125));
sram_cell_6t_5 inst_cell_125_28 (.BL(BL28),.BLN(BLN28),.WL(WL125));
sram_cell_6t_5 inst_cell_125_29 (.BL(BL29),.BLN(BLN29),.WL(WL125));
sram_cell_6t_5 inst_cell_125_30 (.BL(BL30),.BLN(BLN30),.WL(WL125));
sram_cell_6t_5 inst_cell_125_31 (.BL(BL31),.BLN(BLN31),.WL(WL125));
sram_cell_6t_5 inst_cell_125_32 (.BL(BL32),.BLN(BLN32),.WL(WL125));
sram_cell_6t_5 inst_cell_125_33 (.BL(BL33),.BLN(BLN33),.WL(WL125));
sram_cell_6t_5 inst_cell_125_34 (.BL(BL34),.BLN(BLN34),.WL(WL125));
sram_cell_6t_5 inst_cell_125_35 (.BL(BL35),.BLN(BLN35),.WL(WL125));
sram_cell_6t_5 inst_cell_125_36 (.BL(BL36),.BLN(BLN36),.WL(WL125));
sram_cell_6t_5 inst_cell_125_37 (.BL(BL37),.BLN(BLN37),.WL(WL125));
sram_cell_6t_5 inst_cell_125_38 (.BL(BL38),.BLN(BLN38),.WL(WL125));
sram_cell_6t_5 inst_cell_125_39 (.BL(BL39),.BLN(BLN39),.WL(WL125));
sram_cell_6t_5 inst_cell_125_40 (.BL(BL40),.BLN(BLN40),.WL(WL125));
sram_cell_6t_5 inst_cell_125_41 (.BL(BL41),.BLN(BLN41),.WL(WL125));
sram_cell_6t_5 inst_cell_125_42 (.BL(BL42),.BLN(BLN42),.WL(WL125));
sram_cell_6t_5 inst_cell_125_43 (.BL(BL43),.BLN(BLN43),.WL(WL125));
sram_cell_6t_5 inst_cell_125_44 (.BL(BL44),.BLN(BLN44),.WL(WL125));
sram_cell_6t_5 inst_cell_125_45 (.BL(BL45),.BLN(BLN45),.WL(WL125));
sram_cell_6t_5 inst_cell_125_46 (.BL(BL46),.BLN(BLN46),.WL(WL125));
sram_cell_6t_5 inst_cell_125_47 (.BL(BL47),.BLN(BLN47),.WL(WL125));
sram_cell_6t_5 inst_cell_125_48 (.BL(BL48),.BLN(BLN48),.WL(WL125));
sram_cell_6t_5 inst_cell_125_49 (.BL(BL49),.BLN(BLN49),.WL(WL125));
sram_cell_6t_5 inst_cell_125_50 (.BL(BL50),.BLN(BLN50),.WL(WL125));
sram_cell_6t_5 inst_cell_125_51 (.BL(BL51),.BLN(BLN51),.WL(WL125));
sram_cell_6t_5 inst_cell_125_52 (.BL(BL52),.BLN(BLN52),.WL(WL125));
sram_cell_6t_5 inst_cell_125_53 (.BL(BL53),.BLN(BLN53),.WL(WL125));
sram_cell_6t_5 inst_cell_125_54 (.BL(BL54),.BLN(BLN54),.WL(WL125));
sram_cell_6t_5 inst_cell_125_55 (.BL(BL55),.BLN(BLN55),.WL(WL125));
sram_cell_6t_5 inst_cell_125_56 (.BL(BL56),.BLN(BLN56),.WL(WL125));
sram_cell_6t_5 inst_cell_125_57 (.BL(BL57),.BLN(BLN57),.WL(WL125));
sram_cell_6t_5 inst_cell_125_58 (.BL(BL58),.BLN(BLN58),.WL(WL125));
sram_cell_6t_5 inst_cell_125_59 (.BL(BL59),.BLN(BLN59),.WL(WL125));
sram_cell_6t_5 inst_cell_125_60 (.BL(BL60),.BLN(BLN60),.WL(WL125));
sram_cell_6t_5 inst_cell_125_61 (.BL(BL61),.BLN(BLN61),.WL(WL125));
sram_cell_6t_5 inst_cell_125_62 (.BL(BL62),.BLN(BLN62),.WL(WL125));
sram_cell_6t_5 inst_cell_125_63 (.BL(BL63),.BLN(BLN63),.WL(WL125));
sram_cell_6t_5 inst_cell_125_64 (.BL(BL64),.BLN(BLN64),.WL(WL125));
sram_cell_6t_5 inst_cell_125_65 (.BL(BL65),.BLN(BLN65),.WL(WL125));
sram_cell_6t_5 inst_cell_125_66 (.BL(BL66),.BLN(BLN66),.WL(WL125));
sram_cell_6t_5 inst_cell_125_67 (.BL(BL67),.BLN(BLN67),.WL(WL125));
sram_cell_6t_5 inst_cell_125_68 (.BL(BL68),.BLN(BLN68),.WL(WL125));
sram_cell_6t_5 inst_cell_125_69 (.BL(BL69),.BLN(BLN69),.WL(WL125));
sram_cell_6t_5 inst_cell_125_70 (.BL(BL70),.BLN(BLN70),.WL(WL125));
sram_cell_6t_5 inst_cell_125_71 (.BL(BL71),.BLN(BLN71),.WL(WL125));
sram_cell_6t_5 inst_cell_125_72 (.BL(BL72),.BLN(BLN72),.WL(WL125));
sram_cell_6t_5 inst_cell_125_73 (.BL(BL73),.BLN(BLN73),.WL(WL125));
sram_cell_6t_5 inst_cell_125_74 (.BL(BL74),.BLN(BLN74),.WL(WL125));
sram_cell_6t_5 inst_cell_125_75 (.BL(BL75),.BLN(BLN75),.WL(WL125));
sram_cell_6t_5 inst_cell_125_76 (.BL(BL76),.BLN(BLN76),.WL(WL125));
sram_cell_6t_5 inst_cell_125_77 (.BL(BL77),.BLN(BLN77),.WL(WL125));
sram_cell_6t_5 inst_cell_125_78 (.BL(BL78),.BLN(BLN78),.WL(WL125));
sram_cell_6t_5 inst_cell_125_79 (.BL(BL79),.BLN(BLN79),.WL(WL125));
sram_cell_6t_5 inst_cell_125_80 (.BL(BL80),.BLN(BLN80),.WL(WL125));
sram_cell_6t_5 inst_cell_125_81 (.BL(BL81),.BLN(BLN81),.WL(WL125));
sram_cell_6t_5 inst_cell_125_82 (.BL(BL82),.BLN(BLN82),.WL(WL125));
sram_cell_6t_5 inst_cell_125_83 (.BL(BL83),.BLN(BLN83),.WL(WL125));
sram_cell_6t_5 inst_cell_125_84 (.BL(BL84),.BLN(BLN84),.WL(WL125));
sram_cell_6t_5 inst_cell_125_85 (.BL(BL85),.BLN(BLN85),.WL(WL125));
sram_cell_6t_5 inst_cell_125_86 (.BL(BL86),.BLN(BLN86),.WL(WL125));
sram_cell_6t_5 inst_cell_125_87 (.BL(BL87),.BLN(BLN87),.WL(WL125));
sram_cell_6t_5 inst_cell_125_88 (.BL(BL88),.BLN(BLN88),.WL(WL125));
sram_cell_6t_5 inst_cell_125_89 (.BL(BL89),.BLN(BLN89),.WL(WL125));
sram_cell_6t_5 inst_cell_125_90 (.BL(BL90),.BLN(BLN90),.WL(WL125));
sram_cell_6t_5 inst_cell_125_91 (.BL(BL91),.BLN(BLN91),.WL(WL125));
sram_cell_6t_5 inst_cell_125_92 (.BL(BL92),.BLN(BLN92),.WL(WL125));
sram_cell_6t_5 inst_cell_125_93 (.BL(BL93),.BLN(BLN93),.WL(WL125));
sram_cell_6t_5 inst_cell_125_94 (.BL(BL94),.BLN(BLN94),.WL(WL125));
sram_cell_6t_5 inst_cell_125_95 (.BL(BL95),.BLN(BLN95),.WL(WL125));
sram_cell_6t_5 inst_cell_125_96 (.BL(BL96),.BLN(BLN96),.WL(WL125));
sram_cell_6t_5 inst_cell_125_97 (.BL(BL97),.BLN(BLN97),.WL(WL125));
sram_cell_6t_5 inst_cell_125_98 (.BL(BL98),.BLN(BLN98),.WL(WL125));
sram_cell_6t_5 inst_cell_125_99 (.BL(BL99),.BLN(BLN99),.WL(WL125));
sram_cell_6t_5 inst_cell_125_100 (.BL(BL100),.BLN(BLN100),.WL(WL125));
sram_cell_6t_5 inst_cell_125_101 (.BL(BL101),.BLN(BLN101),.WL(WL125));
sram_cell_6t_5 inst_cell_125_102 (.BL(BL102),.BLN(BLN102),.WL(WL125));
sram_cell_6t_5 inst_cell_125_103 (.BL(BL103),.BLN(BLN103),.WL(WL125));
sram_cell_6t_5 inst_cell_125_104 (.BL(BL104),.BLN(BLN104),.WL(WL125));
sram_cell_6t_5 inst_cell_125_105 (.BL(BL105),.BLN(BLN105),.WL(WL125));
sram_cell_6t_5 inst_cell_125_106 (.BL(BL106),.BLN(BLN106),.WL(WL125));
sram_cell_6t_5 inst_cell_125_107 (.BL(BL107),.BLN(BLN107),.WL(WL125));
sram_cell_6t_5 inst_cell_125_108 (.BL(BL108),.BLN(BLN108),.WL(WL125));
sram_cell_6t_5 inst_cell_125_109 (.BL(BL109),.BLN(BLN109),.WL(WL125));
sram_cell_6t_5 inst_cell_125_110 (.BL(BL110),.BLN(BLN110),.WL(WL125));
sram_cell_6t_5 inst_cell_125_111 (.BL(BL111),.BLN(BLN111),.WL(WL125));
sram_cell_6t_5 inst_cell_125_112 (.BL(BL112),.BLN(BLN112),.WL(WL125));
sram_cell_6t_5 inst_cell_125_113 (.BL(BL113),.BLN(BLN113),.WL(WL125));
sram_cell_6t_5 inst_cell_125_114 (.BL(BL114),.BLN(BLN114),.WL(WL125));
sram_cell_6t_5 inst_cell_125_115 (.BL(BL115),.BLN(BLN115),.WL(WL125));
sram_cell_6t_5 inst_cell_125_116 (.BL(BL116),.BLN(BLN116),.WL(WL125));
sram_cell_6t_5 inst_cell_125_117 (.BL(BL117),.BLN(BLN117),.WL(WL125));
sram_cell_6t_5 inst_cell_125_118 (.BL(BL118),.BLN(BLN118),.WL(WL125));
sram_cell_6t_5 inst_cell_125_119 (.BL(BL119),.BLN(BLN119),.WL(WL125));
sram_cell_6t_5 inst_cell_125_120 (.BL(BL120),.BLN(BLN120),.WL(WL125));
sram_cell_6t_5 inst_cell_125_121 (.BL(BL121),.BLN(BLN121),.WL(WL125));
sram_cell_6t_5 inst_cell_125_122 (.BL(BL122),.BLN(BLN122),.WL(WL125));
sram_cell_6t_5 inst_cell_125_123 (.BL(BL123),.BLN(BLN123),.WL(WL125));
sram_cell_6t_5 inst_cell_125_124 (.BL(BL124),.BLN(BLN124),.WL(WL125));
sram_cell_6t_5 inst_cell_125_125 (.BL(BL125),.BLN(BLN125),.WL(WL125));
sram_cell_6t_5 inst_cell_125_126 (.BL(BL126),.BLN(BLN126),.WL(WL125));
sram_cell_6t_5 inst_cell_125_127 (.BL(BL127),.BLN(BLN127),.WL(WL125));
sram_cell_6t_5 inst_cell_126_0 (.BL(BL0),.BLN(BLN0),.WL(WL126));
sram_cell_6t_5 inst_cell_126_1 (.BL(BL1),.BLN(BLN1),.WL(WL126));
sram_cell_6t_5 inst_cell_126_2 (.BL(BL2),.BLN(BLN2),.WL(WL126));
sram_cell_6t_5 inst_cell_126_3 (.BL(BL3),.BLN(BLN3),.WL(WL126));
sram_cell_6t_5 inst_cell_126_4 (.BL(BL4),.BLN(BLN4),.WL(WL126));
sram_cell_6t_5 inst_cell_126_5 (.BL(BL5),.BLN(BLN5),.WL(WL126));
sram_cell_6t_5 inst_cell_126_6 (.BL(BL6),.BLN(BLN6),.WL(WL126));
sram_cell_6t_5 inst_cell_126_7 (.BL(BL7),.BLN(BLN7),.WL(WL126));
sram_cell_6t_5 inst_cell_126_8 (.BL(BL8),.BLN(BLN8),.WL(WL126));
sram_cell_6t_5 inst_cell_126_9 (.BL(BL9),.BLN(BLN9),.WL(WL126));
sram_cell_6t_5 inst_cell_126_10 (.BL(BL10),.BLN(BLN10),.WL(WL126));
sram_cell_6t_5 inst_cell_126_11 (.BL(BL11),.BLN(BLN11),.WL(WL126));
sram_cell_6t_5 inst_cell_126_12 (.BL(BL12),.BLN(BLN12),.WL(WL126));
sram_cell_6t_5 inst_cell_126_13 (.BL(BL13),.BLN(BLN13),.WL(WL126));
sram_cell_6t_5 inst_cell_126_14 (.BL(BL14),.BLN(BLN14),.WL(WL126));
sram_cell_6t_5 inst_cell_126_15 (.BL(BL15),.BLN(BLN15),.WL(WL126));
sram_cell_6t_5 inst_cell_126_16 (.BL(BL16),.BLN(BLN16),.WL(WL126));
sram_cell_6t_5 inst_cell_126_17 (.BL(BL17),.BLN(BLN17),.WL(WL126));
sram_cell_6t_5 inst_cell_126_18 (.BL(BL18),.BLN(BLN18),.WL(WL126));
sram_cell_6t_5 inst_cell_126_19 (.BL(BL19),.BLN(BLN19),.WL(WL126));
sram_cell_6t_5 inst_cell_126_20 (.BL(BL20),.BLN(BLN20),.WL(WL126));
sram_cell_6t_5 inst_cell_126_21 (.BL(BL21),.BLN(BLN21),.WL(WL126));
sram_cell_6t_5 inst_cell_126_22 (.BL(BL22),.BLN(BLN22),.WL(WL126));
sram_cell_6t_5 inst_cell_126_23 (.BL(BL23),.BLN(BLN23),.WL(WL126));
sram_cell_6t_5 inst_cell_126_24 (.BL(BL24),.BLN(BLN24),.WL(WL126));
sram_cell_6t_5 inst_cell_126_25 (.BL(BL25),.BLN(BLN25),.WL(WL126));
sram_cell_6t_5 inst_cell_126_26 (.BL(BL26),.BLN(BLN26),.WL(WL126));
sram_cell_6t_5 inst_cell_126_27 (.BL(BL27),.BLN(BLN27),.WL(WL126));
sram_cell_6t_5 inst_cell_126_28 (.BL(BL28),.BLN(BLN28),.WL(WL126));
sram_cell_6t_5 inst_cell_126_29 (.BL(BL29),.BLN(BLN29),.WL(WL126));
sram_cell_6t_5 inst_cell_126_30 (.BL(BL30),.BLN(BLN30),.WL(WL126));
sram_cell_6t_5 inst_cell_126_31 (.BL(BL31),.BLN(BLN31),.WL(WL126));
sram_cell_6t_5 inst_cell_126_32 (.BL(BL32),.BLN(BLN32),.WL(WL126));
sram_cell_6t_5 inst_cell_126_33 (.BL(BL33),.BLN(BLN33),.WL(WL126));
sram_cell_6t_5 inst_cell_126_34 (.BL(BL34),.BLN(BLN34),.WL(WL126));
sram_cell_6t_5 inst_cell_126_35 (.BL(BL35),.BLN(BLN35),.WL(WL126));
sram_cell_6t_5 inst_cell_126_36 (.BL(BL36),.BLN(BLN36),.WL(WL126));
sram_cell_6t_5 inst_cell_126_37 (.BL(BL37),.BLN(BLN37),.WL(WL126));
sram_cell_6t_5 inst_cell_126_38 (.BL(BL38),.BLN(BLN38),.WL(WL126));
sram_cell_6t_5 inst_cell_126_39 (.BL(BL39),.BLN(BLN39),.WL(WL126));
sram_cell_6t_5 inst_cell_126_40 (.BL(BL40),.BLN(BLN40),.WL(WL126));
sram_cell_6t_5 inst_cell_126_41 (.BL(BL41),.BLN(BLN41),.WL(WL126));
sram_cell_6t_5 inst_cell_126_42 (.BL(BL42),.BLN(BLN42),.WL(WL126));
sram_cell_6t_5 inst_cell_126_43 (.BL(BL43),.BLN(BLN43),.WL(WL126));
sram_cell_6t_5 inst_cell_126_44 (.BL(BL44),.BLN(BLN44),.WL(WL126));
sram_cell_6t_5 inst_cell_126_45 (.BL(BL45),.BLN(BLN45),.WL(WL126));
sram_cell_6t_5 inst_cell_126_46 (.BL(BL46),.BLN(BLN46),.WL(WL126));
sram_cell_6t_5 inst_cell_126_47 (.BL(BL47),.BLN(BLN47),.WL(WL126));
sram_cell_6t_5 inst_cell_126_48 (.BL(BL48),.BLN(BLN48),.WL(WL126));
sram_cell_6t_5 inst_cell_126_49 (.BL(BL49),.BLN(BLN49),.WL(WL126));
sram_cell_6t_5 inst_cell_126_50 (.BL(BL50),.BLN(BLN50),.WL(WL126));
sram_cell_6t_5 inst_cell_126_51 (.BL(BL51),.BLN(BLN51),.WL(WL126));
sram_cell_6t_5 inst_cell_126_52 (.BL(BL52),.BLN(BLN52),.WL(WL126));
sram_cell_6t_5 inst_cell_126_53 (.BL(BL53),.BLN(BLN53),.WL(WL126));
sram_cell_6t_5 inst_cell_126_54 (.BL(BL54),.BLN(BLN54),.WL(WL126));
sram_cell_6t_5 inst_cell_126_55 (.BL(BL55),.BLN(BLN55),.WL(WL126));
sram_cell_6t_5 inst_cell_126_56 (.BL(BL56),.BLN(BLN56),.WL(WL126));
sram_cell_6t_5 inst_cell_126_57 (.BL(BL57),.BLN(BLN57),.WL(WL126));
sram_cell_6t_5 inst_cell_126_58 (.BL(BL58),.BLN(BLN58),.WL(WL126));
sram_cell_6t_5 inst_cell_126_59 (.BL(BL59),.BLN(BLN59),.WL(WL126));
sram_cell_6t_5 inst_cell_126_60 (.BL(BL60),.BLN(BLN60),.WL(WL126));
sram_cell_6t_5 inst_cell_126_61 (.BL(BL61),.BLN(BLN61),.WL(WL126));
sram_cell_6t_5 inst_cell_126_62 (.BL(BL62),.BLN(BLN62),.WL(WL126));
sram_cell_6t_5 inst_cell_126_63 (.BL(BL63),.BLN(BLN63),.WL(WL126));
sram_cell_6t_5 inst_cell_126_64 (.BL(BL64),.BLN(BLN64),.WL(WL126));
sram_cell_6t_5 inst_cell_126_65 (.BL(BL65),.BLN(BLN65),.WL(WL126));
sram_cell_6t_5 inst_cell_126_66 (.BL(BL66),.BLN(BLN66),.WL(WL126));
sram_cell_6t_5 inst_cell_126_67 (.BL(BL67),.BLN(BLN67),.WL(WL126));
sram_cell_6t_5 inst_cell_126_68 (.BL(BL68),.BLN(BLN68),.WL(WL126));
sram_cell_6t_5 inst_cell_126_69 (.BL(BL69),.BLN(BLN69),.WL(WL126));
sram_cell_6t_5 inst_cell_126_70 (.BL(BL70),.BLN(BLN70),.WL(WL126));
sram_cell_6t_5 inst_cell_126_71 (.BL(BL71),.BLN(BLN71),.WL(WL126));
sram_cell_6t_5 inst_cell_126_72 (.BL(BL72),.BLN(BLN72),.WL(WL126));
sram_cell_6t_5 inst_cell_126_73 (.BL(BL73),.BLN(BLN73),.WL(WL126));
sram_cell_6t_5 inst_cell_126_74 (.BL(BL74),.BLN(BLN74),.WL(WL126));
sram_cell_6t_5 inst_cell_126_75 (.BL(BL75),.BLN(BLN75),.WL(WL126));
sram_cell_6t_5 inst_cell_126_76 (.BL(BL76),.BLN(BLN76),.WL(WL126));
sram_cell_6t_5 inst_cell_126_77 (.BL(BL77),.BLN(BLN77),.WL(WL126));
sram_cell_6t_5 inst_cell_126_78 (.BL(BL78),.BLN(BLN78),.WL(WL126));
sram_cell_6t_5 inst_cell_126_79 (.BL(BL79),.BLN(BLN79),.WL(WL126));
sram_cell_6t_5 inst_cell_126_80 (.BL(BL80),.BLN(BLN80),.WL(WL126));
sram_cell_6t_5 inst_cell_126_81 (.BL(BL81),.BLN(BLN81),.WL(WL126));
sram_cell_6t_5 inst_cell_126_82 (.BL(BL82),.BLN(BLN82),.WL(WL126));
sram_cell_6t_5 inst_cell_126_83 (.BL(BL83),.BLN(BLN83),.WL(WL126));
sram_cell_6t_5 inst_cell_126_84 (.BL(BL84),.BLN(BLN84),.WL(WL126));
sram_cell_6t_5 inst_cell_126_85 (.BL(BL85),.BLN(BLN85),.WL(WL126));
sram_cell_6t_5 inst_cell_126_86 (.BL(BL86),.BLN(BLN86),.WL(WL126));
sram_cell_6t_5 inst_cell_126_87 (.BL(BL87),.BLN(BLN87),.WL(WL126));
sram_cell_6t_5 inst_cell_126_88 (.BL(BL88),.BLN(BLN88),.WL(WL126));
sram_cell_6t_5 inst_cell_126_89 (.BL(BL89),.BLN(BLN89),.WL(WL126));
sram_cell_6t_5 inst_cell_126_90 (.BL(BL90),.BLN(BLN90),.WL(WL126));
sram_cell_6t_5 inst_cell_126_91 (.BL(BL91),.BLN(BLN91),.WL(WL126));
sram_cell_6t_5 inst_cell_126_92 (.BL(BL92),.BLN(BLN92),.WL(WL126));
sram_cell_6t_5 inst_cell_126_93 (.BL(BL93),.BLN(BLN93),.WL(WL126));
sram_cell_6t_5 inst_cell_126_94 (.BL(BL94),.BLN(BLN94),.WL(WL126));
sram_cell_6t_5 inst_cell_126_95 (.BL(BL95),.BLN(BLN95),.WL(WL126));
sram_cell_6t_5 inst_cell_126_96 (.BL(BL96),.BLN(BLN96),.WL(WL126));
sram_cell_6t_5 inst_cell_126_97 (.BL(BL97),.BLN(BLN97),.WL(WL126));
sram_cell_6t_5 inst_cell_126_98 (.BL(BL98),.BLN(BLN98),.WL(WL126));
sram_cell_6t_5 inst_cell_126_99 (.BL(BL99),.BLN(BLN99),.WL(WL126));
sram_cell_6t_5 inst_cell_126_100 (.BL(BL100),.BLN(BLN100),.WL(WL126));
sram_cell_6t_5 inst_cell_126_101 (.BL(BL101),.BLN(BLN101),.WL(WL126));
sram_cell_6t_5 inst_cell_126_102 (.BL(BL102),.BLN(BLN102),.WL(WL126));
sram_cell_6t_5 inst_cell_126_103 (.BL(BL103),.BLN(BLN103),.WL(WL126));
sram_cell_6t_5 inst_cell_126_104 (.BL(BL104),.BLN(BLN104),.WL(WL126));
sram_cell_6t_5 inst_cell_126_105 (.BL(BL105),.BLN(BLN105),.WL(WL126));
sram_cell_6t_5 inst_cell_126_106 (.BL(BL106),.BLN(BLN106),.WL(WL126));
sram_cell_6t_5 inst_cell_126_107 (.BL(BL107),.BLN(BLN107),.WL(WL126));
sram_cell_6t_5 inst_cell_126_108 (.BL(BL108),.BLN(BLN108),.WL(WL126));
sram_cell_6t_5 inst_cell_126_109 (.BL(BL109),.BLN(BLN109),.WL(WL126));
sram_cell_6t_5 inst_cell_126_110 (.BL(BL110),.BLN(BLN110),.WL(WL126));
sram_cell_6t_5 inst_cell_126_111 (.BL(BL111),.BLN(BLN111),.WL(WL126));
sram_cell_6t_5 inst_cell_126_112 (.BL(BL112),.BLN(BLN112),.WL(WL126));
sram_cell_6t_5 inst_cell_126_113 (.BL(BL113),.BLN(BLN113),.WL(WL126));
sram_cell_6t_5 inst_cell_126_114 (.BL(BL114),.BLN(BLN114),.WL(WL126));
sram_cell_6t_5 inst_cell_126_115 (.BL(BL115),.BLN(BLN115),.WL(WL126));
sram_cell_6t_5 inst_cell_126_116 (.BL(BL116),.BLN(BLN116),.WL(WL126));
sram_cell_6t_5 inst_cell_126_117 (.BL(BL117),.BLN(BLN117),.WL(WL126));
sram_cell_6t_5 inst_cell_126_118 (.BL(BL118),.BLN(BLN118),.WL(WL126));
sram_cell_6t_5 inst_cell_126_119 (.BL(BL119),.BLN(BLN119),.WL(WL126));
sram_cell_6t_5 inst_cell_126_120 (.BL(BL120),.BLN(BLN120),.WL(WL126));
sram_cell_6t_5 inst_cell_126_121 (.BL(BL121),.BLN(BLN121),.WL(WL126));
sram_cell_6t_5 inst_cell_126_122 (.BL(BL122),.BLN(BLN122),.WL(WL126));
sram_cell_6t_5 inst_cell_126_123 (.BL(BL123),.BLN(BLN123),.WL(WL126));
sram_cell_6t_5 inst_cell_126_124 (.BL(BL124),.BLN(BLN124),.WL(WL126));
sram_cell_6t_5 inst_cell_126_125 (.BL(BL125),.BLN(BLN125),.WL(WL126));
sram_cell_6t_5 inst_cell_126_126 (.BL(BL126),.BLN(BLN126),.WL(WL126));
sram_cell_6t_5 inst_cell_126_127 (.BL(BL127),.BLN(BLN127),.WL(WL126));
sram_cell_6t_5 inst_cell_127_0 (.BL(BL0),.BLN(BLN0),.WL(WL127));
sram_cell_6t_5 inst_cell_127_1 (.BL(BL1),.BLN(BLN1),.WL(WL127));
sram_cell_6t_5 inst_cell_127_2 (.BL(BL2),.BLN(BLN2),.WL(WL127));
sram_cell_6t_5 inst_cell_127_3 (.BL(BL3),.BLN(BLN3),.WL(WL127));
sram_cell_6t_5 inst_cell_127_4 (.BL(BL4),.BLN(BLN4),.WL(WL127));
sram_cell_6t_5 inst_cell_127_5 (.BL(BL5),.BLN(BLN5),.WL(WL127));
sram_cell_6t_5 inst_cell_127_6 (.BL(BL6),.BLN(BLN6),.WL(WL127));
sram_cell_6t_5 inst_cell_127_7 (.BL(BL7),.BLN(BLN7),.WL(WL127));
sram_cell_6t_5 inst_cell_127_8 (.BL(BL8),.BLN(BLN8),.WL(WL127));
sram_cell_6t_5 inst_cell_127_9 (.BL(BL9),.BLN(BLN9),.WL(WL127));
sram_cell_6t_5 inst_cell_127_10 (.BL(BL10),.BLN(BLN10),.WL(WL127));
sram_cell_6t_5 inst_cell_127_11 (.BL(BL11),.BLN(BLN11),.WL(WL127));
sram_cell_6t_5 inst_cell_127_12 (.BL(BL12),.BLN(BLN12),.WL(WL127));
sram_cell_6t_5 inst_cell_127_13 (.BL(BL13),.BLN(BLN13),.WL(WL127));
sram_cell_6t_5 inst_cell_127_14 (.BL(BL14),.BLN(BLN14),.WL(WL127));
sram_cell_6t_5 inst_cell_127_15 (.BL(BL15),.BLN(BLN15),.WL(WL127));
sram_cell_6t_5 inst_cell_127_16 (.BL(BL16),.BLN(BLN16),.WL(WL127));
sram_cell_6t_5 inst_cell_127_17 (.BL(BL17),.BLN(BLN17),.WL(WL127));
sram_cell_6t_5 inst_cell_127_18 (.BL(BL18),.BLN(BLN18),.WL(WL127));
sram_cell_6t_5 inst_cell_127_19 (.BL(BL19),.BLN(BLN19),.WL(WL127));
sram_cell_6t_5 inst_cell_127_20 (.BL(BL20),.BLN(BLN20),.WL(WL127));
sram_cell_6t_5 inst_cell_127_21 (.BL(BL21),.BLN(BLN21),.WL(WL127));
sram_cell_6t_5 inst_cell_127_22 (.BL(BL22),.BLN(BLN22),.WL(WL127));
sram_cell_6t_5 inst_cell_127_23 (.BL(BL23),.BLN(BLN23),.WL(WL127));
sram_cell_6t_5 inst_cell_127_24 (.BL(BL24),.BLN(BLN24),.WL(WL127));
sram_cell_6t_5 inst_cell_127_25 (.BL(BL25),.BLN(BLN25),.WL(WL127));
sram_cell_6t_5 inst_cell_127_26 (.BL(BL26),.BLN(BLN26),.WL(WL127));
sram_cell_6t_5 inst_cell_127_27 (.BL(BL27),.BLN(BLN27),.WL(WL127));
sram_cell_6t_5 inst_cell_127_28 (.BL(BL28),.BLN(BLN28),.WL(WL127));
sram_cell_6t_5 inst_cell_127_29 (.BL(BL29),.BLN(BLN29),.WL(WL127));
sram_cell_6t_5 inst_cell_127_30 (.BL(BL30),.BLN(BLN30),.WL(WL127));
sram_cell_6t_5 inst_cell_127_31 (.BL(BL31),.BLN(BLN31),.WL(WL127));
sram_cell_6t_5 inst_cell_127_32 (.BL(BL32),.BLN(BLN32),.WL(WL127));
sram_cell_6t_5 inst_cell_127_33 (.BL(BL33),.BLN(BLN33),.WL(WL127));
sram_cell_6t_5 inst_cell_127_34 (.BL(BL34),.BLN(BLN34),.WL(WL127));
sram_cell_6t_5 inst_cell_127_35 (.BL(BL35),.BLN(BLN35),.WL(WL127));
sram_cell_6t_5 inst_cell_127_36 (.BL(BL36),.BLN(BLN36),.WL(WL127));
sram_cell_6t_5 inst_cell_127_37 (.BL(BL37),.BLN(BLN37),.WL(WL127));
sram_cell_6t_5 inst_cell_127_38 (.BL(BL38),.BLN(BLN38),.WL(WL127));
sram_cell_6t_5 inst_cell_127_39 (.BL(BL39),.BLN(BLN39),.WL(WL127));
sram_cell_6t_5 inst_cell_127_40 (.BL(BL40),.BLN(BLN40),.WL(WL127));
sram_cell_6t_5 inst_cell_127_41 (.BL(BL41),.BLN(BLN41),.WL(WL127));
sram_cell_6t_5 inst_cell_127_42 (.BL(BL42),.BLN(BLN42),.WL(WL127));
sram_cell_6t_5 inst_cell_127_43 (.BL(BL43),.BLN(BLN43),.WL(WL127));
sram_cell_6t_5 inst_cell_127_44 (.BL(BL44),.BLN(BLN44),.WL(WL127));
sram_cell_6t_5 inst_cell_127_45 (.BL(BL45),.BLN(BLN45),.WL(WL127));
sram_cell_6t_5 inst_cell_127_46 (.BL(BL46),.BLN(BLN46),.WL(WL127));
sram_cell_6t_5 inst_cell_127_47 (.BL(BL47),.BLN(BLN47),.WL(WL127));
sram_cell_6t_5 inst_cell_127_48 (.BL(BL48),.BLN(BLN48),.WL(WL127));
sram_cell_6t_5 inst_cell_127_49 (.BL(BL49),.BLN(BLN49),.WL(WL127));
sram_cell_6t_5 inst_cell_127_50 (.BL(BL50),.BLN(BLN50),.WL(WL127));
sram_cell_6t_5 inst_cell_127_51 (.BL(BL51),.BLN(BLN51),.WL(WL127));
sram_cell_6t_5 inst_cell_127_52 (.BL(BL52),.BLN(BLN52),.WL(WL127));
sram_cell_6t_5 inst_cell_127_53 (.BL(BL53),.BLN(BLN53),.WL(WL127));
sram_cell_6t_5 inst_cell_127_54 (.BL(BL54),.BLN(BLN54),.WL(WL127));
sram_cell_6t_5 inst_cell_127_55 (.BL(BL55),.BLN(BLN55),.WL(WL127));
sram_cell_6t_5 inst_cell_127_56 (.BL(BL56),.BLN(BLN56),.WL(WL127));
sram_cell_6t_5 inst_cell_127_57 (.BL(BL57),.BLN(BLN57),.WL(WL127));
sram_cell_6t_5 inst_cell_127_58 (.BL(BL58),.BLN(BLN58),.WL(WL127));
sram_cell_6t_5 inst_cell_127_59 (.BL(BL59),.BLN(BLN59),.WL(WL127));
sram_cell_6t_5 inst_cell_127_60 (.BL(BL60),.BLN(BLN60),.WL(WL127));
sram_cell_6t_5 inst_cell_127_61 (.BL(BL61),.BLN(BLN61),.WL(WL127));
sram_cell_6t_5 inst_cell_127_62 (.BL(BL62),.BLN(BLN62),.WL(WL127));
sram_cell_6t_5 inst_cell_127_63 (.BL(BL63),.BLN(BLN63),.WL(WL127));
sram_cell_6t_5 inst_cell_127_64 (.BL(BL64),.BLN(BLN64),.WL(WL127));
sram_cell_6t_5 inst_cell_127_65 (.BL(BL65),.BLN(BLN65),.WL(WL127));
sram_cell_6t_5 inst_cell_127_66 (.BL(BL66),.BLN(BLN66),.WL(WL127));
sram_cell_6t_5 inst_cell_127_67 (.BL(BL67),.BLN(BLN67),.WL(WL127));
sram_cell_6t_5 inst_cell_127_68 (.BL(BL68),.BLN(BLN68),.WL(WL127));
sram_cell_6t_5 inst_cell_127_69 (.BL(BL69),.BLN(BLN69),.WL(WL127));
sram_cell_6t_5 inst_cell_127_70 (.BL(BL70),.BLN(BLN70),.WL(WL127));
sram_cell_6t_5 inst_cell_127_71 (.BL(BL71),.BLN(BLN71),.WL(WL127));
sram_cell_6t_5 inst_cell_127_72 (.BL(BL72),.BLN(BLN72),.WL(WL127));
sram_cell_6t_5 inst_cell_127_73 (.BL(BL73),.BLN(BLN73),.WL(WL127));
sram_cell_6t_5 inst_cell_127_74 (.BL(BL74),.BLN(BLN74),.WL(WL127));
sram_cell_6t_5 inst_cell_127_75 (.BL(BL75),.BLN(BLN75),.WL(WL127));
sram_cell_6t_5 inst_cell_127_76 (.BL(BL76),.BLN(BLN76),.WL(WL127));
sram_cell_6t_5 inst_cell_127_77 (.BL(BL77),.BLN(BLN77),.WL(WL127));
sram_cell_6t_5 inst_cell_127_78 (.BL(BL78),.BLN(BLN78),.WL(WL127));
sram_cell_6t_5 inst_cell_127_79 (.BL(BL79),.BLN(BLN79),.WL(WL127));
sram_cell_6t_5 inst_cell_127_80 (.BL(BL80),.BLN(BLN80),.WL(WL127));
sram_cell_6t_5 inst_cell_127_81 (.BL(BL81),.BLN(BLN81),.WL(WL127));
sram_cell_6t_5 inst_cell_127_82 (.BL(BL82),.BLN(BLN82),.WL(WL127));
sram_cell_6t_5 inst_cell_127_83 (.BL(BL83),.BLN(BLN83),.WL(WL127));
sram_cell_6t_5 inst_cell_127_84 (.BL(BL84),.BLN(BLN84),.WL(WL127));
sram_cell_6t_5 inst_cell_127_85 (.BL(BL85),.BLN(BLN85),.WL(WL127));
sram_cell_6t_5 inst_cell_127_86 (.BL(BL86),.BLN(BLN86),.WL(WL127));
sram_cell_6t_5 inst_cell_127_87 (.BL(BL87),.BLN(BLN87),.WL(WL127));
sram_cell_6t_5 inst_cell_127_88 (.BL(BL88),.BLN(BLN88),.WL(WL127));
sram_cell_6t_5 inst_cell_127_89 (.BL(BL89),.BLN(BLN89),.WL(WL127));
sram_cell_6t_5 inst_cell_127_90 (.BL(BL90),.BLN(BLN90),.WL(WL127));
sram_cell_6t_5 inst_cell_127_91 (.BL(BL91),.BLN(BLN91),.WL(WL127));
sram_cell_6t_5 inst_cell_127_92 (.BL(BL92),.BLN(BLN92),.WL(WL127));
sram_cell_6t_5 inst_cell_127_93 (.BL(BL93),.BLN(BLN93),.WL(WL127));
sram_cell_6t_5 inst_cell_127_94 (.BL(BL94),.BLN(BLN94),.WL(WL127));
sram_cell_6t_5 inst_cell_127_95 (.BL(BL95),.BLN(BLN95),.WL(WL127));
sram_cell_6t_5 inst_cell_127_96 (.BL(BL96),.BLN(BLN96),.WL(WL127));
sram_cell_6t_5 inst_cell_127_97 (.BL(BL97),.BLN(BLN97),.WL(WL127));
sram_cell_6t_5 inst_cell_127_98 (.BL(BL98),.BLN(BLN98),.WL(WL127));
sram_cell_6t_5 inst_cell_127_99 (.BL(BL99),.BLN(BLN99),.WL(WL127));
sram_cell_6t_5 inst_cell_127_100 (.BL(BL100),.BLN(BLN100),.WL(WL127));
sram_cell_6t_5 inst_cell_127_101 (.BL(BL101),.BLN(BLN101),.WL(WL127));
sram_cell_6t_5 inst_cell_127_102 (.BL(BL102),.BLN(BLN102),.WL(WL127));
sram_cell_6t_5 inst_cell_127_103 (.BL(BL103),.BLN(BLN103),.WL(WL127));
sram_cell_6t_5 inst_cell_127_104 (.BL(BL104),.BLN(BLN104),.WL(WL127));
sram_cell_6t_5 inst_cell_127_105 (.BL(BL105),.BLN(BLN105),.WL(WL127));
sram_cell_6t_5 inst_cell_127_106 (.BL(BL106),.BLN(BLN106),.WL(WL127));
sram_cell_6t_5 inst_cell_127_107 (.BL(BL107),.BLN(BLN107),.WL(WL127));
sram_cell_6t_5 inst_cell_127_108 (.BL(BL108),.BLN(BLN108),.WL(WL127));
sram_cell_6t_5 inst_cell_127_109 (.BL(BL109),.BLN(BLN109),.WL(WL127));
sram_cell_6t_5 inst_cell_127_110 (.BL(BL110),.BLN(BLN110),.WL(WL127));
sram_cell_6t_5 inst_cell_127_111 (.BL(BL111),.BLN(BLN111),.WL(WL127));
sram_cell_6t_5 inst_cell_127_112 (.BL(BL112),.BLN(BLN112),.WL(WL127));
sram_cell_6t_5 inst_cell_127_113 (.BL(BL113),.BLN(BLN113),.WL(WL127));
sram_cell_6t_5 inst_cell_127_114 (.BL(BL114),.BLN(BLN114),.WL(WL127));
sram_cell_6t_5 inst_cell_127_115 (.BL(BL115),.BLN(BLN115),.WL(WL127));
sram_cell_6t_5 inst_cell_127_116 (.BL(BL116),.BLN(BLN116),.WL(WL127));
sram_cell_6t_5 inst_cell_127_117 (.BL(BL117),.BLN(BLN117),.WL(WL127));
sram_cell_6t_5 inst_cell_127_118 (.BL(BL118),.BLN(BLN118),.WL(WL127));
sram_cell_6t_5 inst_cell_127_119 (.BL(BL119),.BLN(BLN119),.WL(WL127));
sram_cell_6t_5 inst_cell_127_120 (.BL(BL120),.BLN(BLN120),.WL(WL127));
sram_cell_6t_5 inst_cell_127_121 (.BL(BL121),.BLN(BLN121),.WL(WL127));
sram_cell_6t_5 inst_cell_127_122 (.BL(BL122),.BLN(BLN122),.WL(WL127));
sram_cell_6t_5 inst_cell_127_123 (.BL(BL123),.BLN(BLN123),.WL(WL127));
sram_cell_6t_5 inst_cell_127_124 (.BL(BL124),.BLN(BLN124),.WL(WL127));
sram_cell_6t_5 inst_cell_127_125 (.BL(BL125),.BLN(BLN125),.WL(WL127));
sram_cell_6t_5 inst_cell_127_126 (.BL(BL126),.BLN(BLN126),.WL(WL127));
sram_cell_6t_5 inst_cell_127_127 (.BL(BL127),.BLN(BLN127),.WL(WL127));
columnMux inst_colMux0 (BL0,BLN0,BL1,BLN1,BL2,BLN2,BL3,BLN3,SL0,SL1,SL2,SL3,DL0,DLN0);
write_driver_compiler inst_writeDriver0 (.clk(clk_bar),.data(din0),.write_en(write_en),.BL(DL0),.BLN(DLN0));
sense_amp_clocked_compiler inst_senAmp0 (.bit(DL0),.bit_bar(DLN0),.sense_en(sense_en),.sense(dout0));
columnMux inst_colMux1 (BL4,BLN4,BL5,BLN5,BL6,BLN6,BL7,BLN7,SL0,SL1,SL2,SL3,DL1,DLN1);
write_driver_compiler inst_writeDriver1 (.clk(clk_bar),.data(din1),.write_en(write_en),.BL(DL1),.BLN(DLN1));
sense_amp_clocked_compiler inst_senAmp1 (.bit(DL1),.bit_bar(DLN1),.sense_en(sense_en),.sense(dout1));
columnMux inst_colMux2 (BL8,BLN8,BL9,BLN9,BL10,BLN10,BL11,BLN11,SL0,SL1,SL2,SL3,DL2,DLN2);
write_driver_compiler inst_writeDriver2 (.clk(clk_bar),.data(din2),.write_en(write_en),.BL(DL2),.BLN(DLN2));
sense_amp_clocked_compiler inst_senAmp2 (.bit(DL2),.bit_bar(DLN2),.sense_en(sense_en),.sense(dout2));
columnMux inst_colMux3 (BL12,BLN12,BL13,BLN13,BL14,BLN14,BL15,BLN15,SL0,SL1,SL2,SL3,DL3,DLN3);
write_driver_compiler inst_writeDriver3 (.clk(clk_bar),.data(din3),.write_en(write_en),.BL(DL3),.BLN(DLN3));
sense_amp_clocked_compiler inst_senAmp3 (.bit(DL3),.bit_bar(DLN3),.sense_en(sense_en),.sense(dout3));
columnMux inst_colMux4 (BL16,BLN16,BL17,BLN17,BL18,BLN18,BL19,BLN19,SL0,SL1,SL2,SL3,DL4,DLN4);
write_driver_compiler inst_writeDriver4 (.clk(clk_bar),.data(din4),.write_en(write_en),.BL(DL4),.BLN(DLN4));
sense_amp_clocked_compiler inst_senAmp4 (.bit(DL4),.bit_bar(DLN4),.sense_en(sense_en),.sense(dout4));
columnMux inst_colMux5 (BL20,BLN20,BL21,BLN21,BL22,BLN22,BL23,BLN23,SL0,SL1,SL2,SL3,DL5,DLN5);
write_driver_compiler inst_writeDriver5 (.clk(clk_bar),.data(din5),.write_en(write_en),.BL(DL5),.BLN(DLN5));
sense_amp_clocked_compiler inst_senAmp5 (.bit(DL5),.bit_bar(DLN5),.sense_en(sense_en),.sense(dout5));
columnMux inst_colMux6 (BL24,BLN24,BL25,BLN25,BL26,BLN26,BL27,BLN27,SL0,SL1,SL2,SL3,DL6,DLN6);
write_driver_compiler inst_writeDriver6 (.clk(clk_bar),.data(din6),.write_en(write_en),.BL(DL6),.BLN(DLN6));
sense_amp_clocked_compiler inst_senAmp6 (.bit(DL6),.bit_bar(DLN6),.sense_en(sense_en),.sense(dout6));
columnMux inst_colMux7 (BL28,BLN28,BL29,BLN29,BL30,BLN30,BL31,BLN31,SL0,SL1,SL2,SL3,DL7,DLN7);
write_driver_compiler inst_writeDriver7 (.clk(clk_bar),.data(din7),.write_en(write_en),.BL(DL7),.BLN(DLN7));
sense_amp_clocked_compiler inst_senAmp7 (.bit(DL7),.bit_bar(DLN7),.sense_en(sense_en),.sense(dout7));
columnMux inst_colMux8 (BL32,BLN32,BL33,BLN33,BL34,BLN34,BL35,BLN35,SL0,SL1,SL2,SL3,DL8,DLN8);
write_driver_compiler inst_writeDriver8 (.clk(clk_bar),.data(din8),.write_en(write_en),.BL(DL8),.BLN(DLN8));
sense_amp_clocked_compiler inst_senAmp8 (.bit(DL8),.bit_bar(DLN8),.sense_en(sense_en),.sense(dout8));
columnMux inst_colMux9 (BL36,BLN36,BL37,BLN37,BL38,BLN38,BL39,BLN39,SL0,SL1,SL2,SL3,DL9,DLN9);
write_driver_compiler inst_writeDriver9 (.clk(clk_bar),.data(din9),.write_en(write_en),.BL(DL9),.BLN(DLN9));
sense_amp_clocked_compiler inst_senAmp9 (.bit(DL9),.bit_bar(DLN9),.sense_en(sense_en),.sense(dout9));
columnMux inst_colMux10 (BL40,BLN40,BL41,BLN41,BL42,BLN42,BL43,BLN43,SL0,SL1,SL2,SL3,DL10,DLN10);
write_driver_compiler inst_writeDriver10 (.clk(clk_bar),.data(din10),.write_en(write_en),.BL(DL10),.BLN(DLN10));
sense_amp_clocked_compiler inst_senAmp10 (.bit(DL10),.bit_bar(DLN10),.sense_en(sense_en),.sense(dout10));
columnMux inst_colMux11 (BL44,BLN44,BL45,BLN45,BL46,BLN46,BL47,BLN47,SL0,SL1,SL2,SL3,DL11,DLN11);
write_driver_compiler inst_writeDriver11 (.clk(clk_bar),.data(din11),.write_en(write_en),.BL(DL11),.BLN(DLN11));
sense_amp_clocked_compiler inst_senAmp11 (.bit(DL11),.bit_bar(DLN11),.sense_en(sense_en),.sense(dout11));
columnMux inst_colMux12 (BL48,BLN48,BL49,BLN49,BL50,BLN50,BL51,BLN51,SL0,SL1,SL2,SL3,DL12,DLN12);
write_driver_compiler inst_writeDriver12 (.clk(clk_bar),.data(din12),.write_en(write_en),.BL(DL12),.BLN(DLN12));
sense_amp_clocked_compiler inst_senAmp12 (.bit(DL12),.bit_bar(DLN12),.sense_en(sense_en),.sense(dout12));
columnMux inst_colMux13 (BL52,BLN52,BL53,BLN53,BL54,BLN54,BL55,BLN55,SL0,SL1,SL2,SL3,DL13,DLN13);
write_driver_compiler inst_writeDriver13 (.clk(clk_bar),.data(din13),.write_en(write_en),.BL(DL13),.BLN(DLN13));
sense_amp_clocked_compiler inst_senAmp13 (.bit(DL13),.bit_bar(DLN13),.sense_en(sense_en),.sense(dout13));
columnMux inst_colMux14 (BL56,BLN56,BL57,BLN57,BL58,BLN58,BL59,BLN59,SL0,SL1,SL2,SL3,DL14,DLN14);
write_driver_compiler inst_writeDriver14 (.clk(clk_bar),.data(din14),.write_en(write_en),.BL(DL14),.BLN(DLN14));
sense_amp_clocked_compiler inst_senAmp14 (.bit(DL14),.bit_bar(DLN14),.sense_en(sense_en),.sense(dout14));
columnMux inst_colMux15 (BL60,BLN60,BL61,BLN61,BL62,BLN62,BL63,BLN63,SL0,SL1,SL2,SL3,DL15,DLN15);
write_driver_compiler inst_writeDriver15 (.clk(clk_bar),.data(din15),.write_en(write_en),.BL(DL15),.BLN(DLN15));
sense_amp_clocked_compiler inst_senAmp15 (.bit(DL15),.bit_bar(DLN15),.sense_en(sense_en),.sense(dout15));
columnMux inst_colMux16 (BL64,BLN64,BL65,BLN65,BL66,BLN66,BL67,BLN67,SL0,SL1,SL2,SL3,DL16,DLN16);
write_driver_compiler inst_writeDriver16 (.clk(clk_bar),.data(din16),.write_en(write_en),.BL(DL16),.BLN(DLN16));
sense_amp_clocked_compiler inst_senAmp16 (.bit(DL16),.bit_bar(DLN16),.sense_en(sense_en),.sense(dout16));
columnMux inst_colMux17 (BL68,BLN68,BL69,BLN69,BL70,BLN70,BL71,BLN71,SL0,SL1,SL2,SL3,DL17,DLN17);
write_driver_compiler inst_writeDriver17 (.clk(clk_bar),.data(din17),.write_en(write_en),.BL(DL17),.BLN(DLN17));
sense_amp_clocked_compiler inst_senAmp17 (.bit(DL17),.bit_bar(DLN17),.sense_en(sense_en),.sense(dout17));
columnMux inst_colMux18 (BL72,BLN72,BL73,BLN73,BL74,BLN74,BL75,BLN75,SL0,SL1,SL2,SL3,DL18,DLN18);
write_driver_compiler inst_writeDriver18 (.clk(clk_bar),.data(din18),.write_en(write_en),.BL(DL18),.BLN(DLN18));
sense_amp_clocked_compiler inst_senAmp18 (.bit(DL18),.bit_bar(DLN18),.sense_en(sense_en),.sense(dout18));
columnMux inst_colMux19 (BL76,BLN76,BL77,BLN77,BL78,BLN78,BL79,BLN79,SL0,SL1,SL2,SL3,DL19,DLN19);
write_driver_compiler inst_writeDriver19 (.clk(clk_bar),.data(din19),.write_en(write_en),.BL(DL19),.BLN(DLN19));
sense_amp_clocked_compiler inst_senAmp19 (.bit(DL19),.bit_bar(DLN19),.sense_en(sense_en),.sense(dout19));
columnMux inst_colMux20 (BL80,BLN80,BL81,BLN81,BL82,BLN82,BL83,BLN83,SL0,SL1,SL2,SL3,DL20,DLN20);
write_driver_compiler inst_writeDriver20 (.clk(clk_bar),.data(din20),.write_en(write_en),.BL(DL20),.BLN(DLN20));
sense_amp_clocked_compiler inst_senAmp20 (.bit(DL20),.bit_bar(DLN20),.sense_en(sense_en),.sense(dout20));
columnMux inst_colMux21 (BL84,BLN84,BL85,BLN85,BL86,BLN86,BL87,BLN87,SL0,SL1,SL2,SL3,DL21,DLN21);
write_driver_compiler inst_writeDriver21 (.clk(clk_bar),.data(din21),.write_en(write_en),.BL(DL21),.BLN(DLN21));
sense_amp_clocked_compiler inst_senAmp21 (.bit(DL21),.bit_bar(DLN21),.sense_en(sense_en),.sense(dout21));
columnMux inst_colMux22 (BL88,BLN88,BL89,BLN89,BL90,BLN90,BL91,BLN91,SL0,SL1,SL2,SL3,DL22,DLN22);
write_driver_compiler inst_writeDriver22 (.clk(clk_bar),.data(din22),.write_en(write_en),.BL(DL22),.BLN(DLN22));
sense_amp_clocked_compiler inst_senAmp22 (.bit(DL22),.bit_bar(DLN22),.sense_en(sense_en),.sense(dout22));
columnMux inst_colMux23 (BL92,BLN92,BL93,BLN93,BL94,BLN94,BL95,BLN95,SL0,SL1,SL2,SL3,DL23,DLN23);
write_driver_compiler inst_writeDriver23 (.clk(clk_bar),.data(din23),.write_en(write_en),.BL(DL23),.BLN(DLN23));
sense_amp_clocked_compiler inst_senAmp23 (.bit(DL23),.bit_bar(DLN23),.sense_en(sense_en),.sense(dout23));
columnMux inst_colMux24 (BL96,BLN96,BL97,BLN97,BL98,BLN98,BL99,BLN99,SL0,SL1,SL2,SL3,DL24,DLN24);
write_driver_compiler inst_writeDriver24 (.clk(clk_bar),.data(din24),.write_en(write_en),.BL(DL24),.BLN(DLN24));
sense_amp_clocked_compiler inst_senAmp24 (.bit(DL24),.bit_bar(DLN24),.sense_en(sense_en),.sense(dout24));
columnMux inst_colMux25 (BL100,BLN100,BL101,BLN101,BL102,BLN102,BL103,BLN103,SL0,SL1,SL2,SL3,DL25,DLN25);
write_driver_compiler inst_writeDriver25 (.clk(clk_bar),.data(din25),.write_en(write_en),.BL(DL25),.BLN(DLN25));
sense_amp_clocked_compiler inst_senAmp25 (.bit(DL25),.bit_bar(DLN25),.sense_en(sense_en),.sense(dout25));
columnMux inst_colMux26 (BL104,BLN104,BL105,BLN105,BL106,BLN106,BL107,BLN107,SL0,SL1,SL2,SL3,DL26,DLN26);
write_driver_compiler inst_writeDriver26 (.clk(clk_bar),.data(din26),.write_en(write_en),.BL(DL26),.BLN(DLN26));
sense_amp_clocked_compiler inst_senAmp26 (.bit(DL26),.bit_bar(DLN26),.sense_en(sense_en),.sense(dout26));
columnMux inst_colMux27 (BL108,BLN108,BL109,BLN109,BL110,BLN110,BL111,BLN111,SL0,SL1,SL2,SL3,DL27,DLN27);
write_driver_compiler inst_writeDriver27 (.clk(clk_bar),.data(din27),.write_en(write_en),.BL(DL27),.BLN(DLN27));
sense_amp_clocked_compiler inst_senAmp27 (.bit(DL27),.bit_bar(DLN27),.sense_en(sense_en),.sense(dout27));
columnMux inst_colMux28 (BL112,BLN112,BL113,BLN113,BL114,BLN114,BL115,BLN115,SL0,SL1,SL2,SL3,DL28,DLN28);
write_driver_compiler inst_writeDriver28 (.clk(clk_bar),.data(din28),.write_en(write_en),.BL(DL28),.BLN(DLN28));
sense_amp_clocked_compiler inst_senAmp28 (.bit(DL28),.bit_bar(DLN28),.sense_en(sense_en),.sense(dout28));
columnMux inst_colMux29 (BL116,BLN116,BL117,BLN117,BL118,BLN118,BL119,BLN119,SL0,SL1,SL2,SL3,DL29,DLN29);
write_driver_compiler inst_writeDriver29 (.clk(clk_bar),.data(din29),.write_en(write_en),.BL(DL29),.BLN(DLN29));
sense_amp_clocked_compiler inst_senAmp29 (.bit(DL29),.bit_bar(DLN29),.sense_en(sense_en),.sense(dout29));
columnMux inst_colMux30 (BL120,BLN120,BL121,BLN121,BL122,BLN122,BL123,BLN123,SL0,SL1,SL2,SL3,DL30,DLN30);
write_driver_compiler inst_writeDriver30 (.clk(clk_bar),.data(din30),.write_en(write_en),.BL(DL30),.BLN(DLN30));
sense_amp_clocked_compiler inst_senAmp30 (.bit(DL30),.bit_bar(DLN30),.sense_en(sense_en),.sense(dout30));
columnMux inst_colMux31 (BL124,BLN124,BL125,BLN125,BL126,BLN126,BL127,BLN127,SL0,SL1,SL2,SL3,DL31,DLN31);
write_driver_compiler inst_writeDriver31 (.clk(clk_bar),.data(din31),.write_en(write_en),.BL(DL31),.BLN(DLN31));
sense_amp_clocked_compiler inst_senAmp31 (.bit(DL31),.bit_bar(DLN31),.sense_en(sense_en),.sense(dout31));
precharge_compiler inst_precharge0 (.clk(clk_bar),.B(BL0),.B_bar(BLN0));
precharge_compiler inst_precharge1 (.clk(clk_bar),.B(BL1),.B_bar(BLN1));
precharge_compiler inst_precharge2 (.clk(clk_bar),.B(BL2),.B_bar(BLN2));
precharge_compiler inst_precharge3 (.clk(clk_bar),.B(BL3),.B_bar(BLN3));
precharge_compiler inst_precharge4 (.clk(clk_bar),.B(BL4),.B_bar(BLN4));
precharge_compiler inst_precharge5 (.clk(clk_bar),.B(BL5),.B_bar(BLN5));
precharge_compiler inst_precharge6 (.clk(clk_bar),.B(BL6),.B_bar(BLN6));
precharge_compiler inst_precharge7 (.clk(clk_bar),.B(BL7),.B_bar(BLN7));
precharge_compiler inst_precharge8 (.clk(clk_bar),.B(BL8),.B_bar(BLN8));
precharge_compiler inst_precharge9 (.clk(clk_bar),.B(BL9),.B_bar(BLN9));
precharge_compiler inst_precharge10 (.clk(clk_bar),.B(BL10),.B_bar(BLN10));
precharge_compiler inst_precharge11 (.clk(clk_bar),.B(BL11),.B_bar(BLN11));
precharge_compiler inst_precharge12 (.clk(clk_bar),.B(BL12),.B_bar(BLN12));
precharge_compiler inst_precharge13 (.clk(clk_bar),.B(BL13),.B_bar(BLN13));
precharge_compiler inst_precharge14 (.clk(clk_bar),.B(BL14),.B_bar(BLN14));
precharge_compiler inst_precharge15 (.clk(clk_bar),.B(BL15),.B_bar(BLN15));
precharge_compiler inst_precharge16 (.clk(clk_bar),.B(BL16),.B_bar(BLN16));
precharge_compiler inst_precharge17 (.clk(clk_bar),.B(BL17),.B_bar(BLN17));
precharge_compiler inst_precharge18 (.clk(clk_bar),.B(BL18),.B_bar(BLN18));
precharge_compiler inst_precharge19 (.clk(clk_bar),.B(BL19),.B_bar(BLN19));
precharge_compiler inst_precharge20 (.clk(clk_bar),.B(BL20),.B_bar(BLN20));
precharge_compiler inst_precharge21 (.clk(clk_bar),.B(BL21),.B_bar(BLN21));
precharge_compiler inst_precharge22 (.clk(clk_bar),.B(BL22),.B_bar(BLN22));
precharge_compiler inst_precharge23 (.clk(clk_bar),.B(BL23),.B_bar(BLN23));
precharge_compiler inst_precharge24 (.clk(clk_bar),.B(BL24),.B_bar(BLN24));
precharge_compiler inst_precharge25 (.clk(clk_bar),.B(BL25),.B_bar(BLN25));
precharge_compiler inst_precharge26 (.clk(clk_bar),.B(BL26),.B_bar(BLN26));
precharge_compiler inst_precharge27 (.clk(clk_bar),.B(BL27),.B_bar(BLN27));
precharge_compiler inst_precharge28 (.clk(clk_bar),.B(BL28),.B_bar(BLN28));
precharge_compiler inst_precharge29 (.clk(clk_bar),.B(BL29),.B_bar(BLN29));
precharge_compiler inst_precharge30 (.clk(clk_bar),.B(BL30),.B_bar(BLN30));
precharge_compiler inst_precharge31 (.clk(clk_bar),.B(BL31),.B_bar(BLN31));
precharge_compiler inst_precharge32 (.clk(clk_bar),.B(BL32),.B_bar(BLN32));
precharge_compiler inst_precharge33 (.clk(clk_bar),.B(BL33),.B_bar(BLN33));
precharge_compiler inst_precharge34 (.clk(clk_bar),.B(BL34),.B_bar(BLN34));
precharge_compiler inst_precharge35 (.clk(clk_bar),.B(BL35),.B_bar(BLN35));
precharge_compiler inst_precharge36 (.clk(clk_bar),.B(BL36),.B_bar(BLN36));
precharge_compiler inst_precharge37 (.clk(clk_bar),.B(BL37),.B_bar(BLN37));
precharge_compiler inst_precharge38 (.clk(clk_bar),.B(BL38),.B_bar(BLN38));
precharge_compiler inst_precharge39 (.clk(clk_bar),.B(BL39),.B_bar(BLN39));
precharge_compiler inst_precharge40 (.clk(clk_bar),.B(BL40),.B_bar(BLN40));
precharge_compiler inst_precharge41 (.clk(clk_bar),.B(BL41),.B_bar(BLN41));
precharge_compiler inst_precharge42 (.clk(clk_bar),.B(BL42),.B_bar(BLN42));
precharge_compiler inst_precharge43 (.clk(clk_bar),.B(BL43),.B_bar(BLN43));
precharge_compiler inst_precharge44 (.clk(clk_bar),.B(BL44),.B_bar(BLN44));
precharge_compiler inst_precharge45 (.clk(clk_bar),.B(BL45),.B_bar(BLN45));
precharge_compiler inst_precharge46 (.clk(clk_bar),.B(BL46),.B_bar(BLN46));
precharge_compiler inst_precharge47 (.clk(clk_bar),.B(BL47),.B_bar(BLN47));
precharge_compiler inst_precharge48 (.clk(clk_bar),.B(BL48),.B_bar(BLN48));
precharge_compiler inst_precharge49 (.clk(clk_bar),.B(BL49),.B_bar(BLN49));
precharge_compiler inst_precharge50 (.clk(clk_bar),.B(BL50),.B_bar(BLN50));
precharge_compiler inst_precharge51 (.clk(clk_bar),.B(BL51),.B_bar(BLN51));
precharge_compiler inst_precharge52 (.clk(clk_bar),.B(BL52),.B_bar(BLN52));
precharge_compiler inst_precharge53 (.clk(clk_bar),.B(BL53),.B_bar(BLN53));
precharge_compiler inst_precharge54 (.clk(clk_bar),.B(BL54),.B_bar(BLN54));
precharge_compiler inst_precharge55 (.clk(clk_bar),.B(BL55),.B_bar(BLN55));
precharge_compiler inst_precharge56 (.clk(clk_bar),.B(BL56),.B_bar(BLN56));
precharge_compiler inst_precharge57 (.clk(clk_bar),.B(BL57),.B_bar(BLN57));
precharge_compiler inst_precharge58 (.clk(clk_bar),.B(BL58),.B_bar(BLN58));
precharge_compiler inst_precharge59 (.clk(clk_bar),.B(BL59),.B_bar(BLN59));
precharge_compiler inst_precharge60 (.clk(clk_bar),.B(BL60),.B_bar(BLN60));
precharge_compiler inst_precharge61 (.clk(clk_bar),.B(BL61),.B_bar(BLN61));
precharge_compiler inst_precharge62 (.clk(clk_bar),.B(BL62),.B_bar(BLN62));
precharge_compiler inst_precharge63 (.clk(clk_bar),.B(BL63),.B_bar(BLN63));
precharge_compiler inst_precharge64 (.clk(clk_bar),.B(BL64),.B_bar(BLN64));
precharge_compiler inst_precharge65 (.clk(clk_bar),.B(BL65),.B_bar(BLN65));
precharge_compiler inst_precharge66 (.clk(clk_bar),.B(BL66),.B_bar(BLN66));
precharge_compiler inst_precharge67 (.clk(clk_bar),.B(BL67),.B_bar(BLN67));
precharge_compiler inst_precharge68 (.clk(clk_bar),.B(BL68),.B_bar(BLN68));
precharge_compiler inst_precharge69 (.clk(clk_bar),.B(BL69),.B_bar(BLN69));
precharge_compiler inst_precharge70 (.clk(clk_bar),.B(BL70),.B_bar(BLN70));
precharge_compiler inst_precharge71 (.clk(clk_bar),.B(BL71),.B_bar(BLN71));
precharge_compiler inst_precharge72 (.clk(clk_bar),.B(BL72),.B_bar(BLN72));
precharge_compiler inst_precharge73 (.clk(clk_bar),.B(BL73),.B_bar(BLN73));
precharge_compiler inst_precharge74 (.clk(clk_bar),.B(BL74),.B_bar(BLN74));
precharge_compiler inst_precharge75 (.clk(clk_bar),.B(BL75),.B_bar(BLN75));
precharge_compiler inst_precharge76 (.clk(clk_bar),.B(BL76),.B_bar(BLN76));
precharge_compiler inst_precharge77 (.clk(clk_bar),.B(BL77),.B_bar(BLN77));
precharge_compiler inst_precharge78 (.clk(clk_bar),.B(BL78),.B_bar(BLN78));
precharge_compiler inst_precharge79 (.clk(clk_bar),.B(BL79),.B_bar(BLN79));
precharge_compiler inst_precharge80 (.clk(clk_bar),.B(BL80),.B_bar(BLN80));
precharge_compiler inst_precharge81 (.clk(clk_bar),.B(BL81),.B_bar(BLN81));
precharge_compiler inst_precharge82 (.clk(clk_bar),.B(BL82),.B_bar(BLN82));
precharge_compiler inst_precharge83 (.clk(clk_bar),.B(BL83),.B_bar(BLN83));
precharge_compiler inst_precharge84 (.clk(clk_bar),.B(BL84),.B_bar(BLN84));
precharge_compiler inst_precharge85 (.clk(clk_bar),.B(BL85),.B_bar(BLN85));
precharge_compiler inst_precharge86 (.clk(clk_bar),.B(BL86),.B_bar(BLN86));
precharge_compiler inst_precharge87 (.clk(clk_bar),.B(BL87),.B_bar(BLN87));
precharge_compiler inst_precharge88 (.clk(clk_bar),.B(BL88),.B_bar(BLN88));
precharge_compiler inst_precharge89 (.clk(clk_bar),.B(BL89),.B_bar(BLN89));
precharge_compiler inst_precharge90 (.clk(clk_bar),.B(BL90),.B_bar(BLN90));
precharge_compiler inst_precharge91 (.clk(clk_bar),.B(BL91),.B_bar(BLN91));
precharge_compiler inst_precharge92 (.clk(clk_bar),.B(BL92),.B_bar(BLN92));
precharge_compiler inst_precharge93 (.clk(clk_bar),.B(BL93),.B_bar(BLN93));
precharge_compiler inst_precharge94 (.clk(clk_bar),.B(BL94),.B_bar(BLN94));
precharge_compiler inst_precharge95 (.clk(clk_bar),.B(BL95),.B_bar(BLN95));
precharge_compiler inst_precharge96 (.clk(clk_bar),.B(BL96),.B_bar(BLN96));
precharge_compiler inst_precharge97 (.clk(clk_bar),.B(BL97),.B_bar(BLN97));
precharge_compiler inst_precharge98 (.clk(clk_bar),.B(BL98),.B_bar(BLN98));
precharge_compiler inst_precharge99 (.clk(clk_bar),.B(BL99),.B_bar(BLN99));
precharge_compiler inst_precharge100 (.clk(clk_bar),.B(BL100),.B_bar(BLN100));
precharge_compiler inst_precharge101 (.clk(clk_bar),.B(BL101),.B_bar(BLN101));
precharge_compiler inst_precharge102 (.clk(clk_bar),.B(BL102),.B_bar(BLN102));
precharge_compiler inst_precharge103 (.clk(clk_bar),.B(BL103),.B_bar(BLN103));
precharge_compiler inst_precharge104 (.clk(clk_bar),.B(BL104),.B_bar(BLN104));
precharge_compiler inst_precharge105 (.clk(clk_bar),.B(BL105),.B_bar(BLN105));
precharge_compiler inst_precharge106 (.clk(clk_bar),.B(BL106),.B_bar(BLN106));
precharge_compiler inst_precharge107 (.clk(clk_bar),.B(BL107),.B_bar(BLN107));
precharge_compiler inst_precharge108 (.clk(clk_bar),.B(BL108),.B_bar(BLN108));
precharge_compiler inst_precharge109 (.clk(clk_bar),.B(BL109),.B_bar(BLN109));
precharge_compiler inst_precharge110 (.clk(clk_bar),.B(BL110),.B_bar(BLN110));
precharge_compiler inst_precharge111 (.clk(clk_bar),.B(BL111),.B_bar(BLN111));
precharge_compiler inst_precharge112 (.clk(clk_bar),.B(BL112),.B_bar(BLN112));
precharge_compiler inst_precharge113 (.clk(clk_bar),.B(BL113),.B_bar(BLN113));
precharge_compiler inst_precharge114 (.clk(clk_bar),.B(BL114),.B_bar(BLN114));
precharge_compiler inst_precharge115 (.clk(clk_bar),.B(BL115),.B_bar(BLN115));
precharge_compiler inst_precharge116 (.clk(clk_bar),.B(BL116),.B_bar(BLN116));
precharge_compiler inst_precharge117 (.clk(clk_bar),.B(BL117),.B_bar(BLN117));
precharge_compiler inst_precharge118 (.clk(clk_bar),.B(BL118),.B_bar(BLN118));
precharge_compiler inst_precharge119 (.clk(clk_bar),.B(BL119),.B_bar(BLN119));
precharge_compiler inst_precharge120 (.clk(clk_bar),.B(BL120),.B_bar(BLN120));
precharge_compiler inst_precharge121 (.clk(clk_bar),.B(BL121),.B_bar(BLN121));
precharge_compiler inst_precharge122 (.clk(clk_bar),.B(BL122),.B_bar(BLN122));
precharge_compiler inst_precharge123 (.clk(clk_bar),.B(BL123),.B_bar(BLN123));
precharge_compiler inst_precharge124 (.clk(clk_bar),.B(BL124),.B_bar(BLN124));
precharge_compiler inst_precharge125 (.clk(clk_bar),.B(BL125),.B_bar(BLN125));
precharge_compiler inst_precharge126 (.clk(clk_bar),.B(BL126),.B_bar(BLN126));
precharge_compiler inst_precharge127 (.clk(clk_bar),.B(BL127),.B_bar(BLN127));
endmodule
