module invRow(A0,A1,A2,A3,A4,A5,A6,A7,Abar0,Abar1,Abar2,Abar3,Abar4,Abar5,Abar6,Abar7);
input A0;
input A1;
input A2;
input A3;
input A4;
input A5;
input A6;
input A7;
output Abar0;
output Abar1;
output Abar2;
output Abar3;
output Abar4;
output Abar5;
output Abar6;
output Abar7;
INVD wire0 (.A(A0),.Y(Abar0));
INVD wire1 (.A(A1),.Y(Abar1));
INVD wire2 (.A(A2),.Y(Abar2));
INVD wire3 (.A(A3),.Y(Abar3));
INVD wire4 (.A(A4),.Y(Abar4));
INVD wire5 (.A(A5),.Y(Abar5));
INVD wire6 (.A(A6),.Y(Abar6));
INVD wire7 (.A(A7),.Y(Abar7));
endmodule
module invCol(A0,A1,A2,A3,Abar0,Abar1,Abar2,Abar3);
input A0;
input A1;
input A2;
input A3;
output Abar0;
output Abar1;
output Abar2;
output Abar3;
INVD wire0 (.A(A0),.Y(Abar0));
INVD wire1 (.A(A1),.Y(Abar1));
INVD wire2 (.A(A2),.Y(Abar2));
INVD wire3 (.A(A3),.Y(Abar3));
endmodule
module rowDecoder(A0,A0_inv,A1,A1_inv,A2,A2_inv,A3,A3_inv,A4,A4_inv,A5,A5_inv,A6,A6_inv,A7,A7_inv,CLK,YF0,YF1,YF2,YF3,YF4,YF5,YF6,YF7,YF8,YF9,YF10,YF11,YF12,YF13,YF14,YF15,YF16,YF17,YF18,YF19,YF20,YF21,YF22,YF23,YF24,YF25,YF26,YF27,YF28,YF29,YF30,YF31,YF32,YF33,YF34,YF35,YF36,YF37,YF38,YF39,YF40,YF41,YF42,YF43,YF44,YF45,YF46,YF47,YF48,YF49,YF50,YF51,YF52,YF53,YF54,YF55,YF56,YF57,YF58,YF59,YF60,YF61,YF62,YF63,YF64,YF65,YF66,YF67,YF68,YF69,YF70,YF71,YF72,YF73,YF74,YF75,YF76,YF77,YF78,YF79,YF80,YF81,YF82,YF83,YF84,YF85,YF86,YF87,YF88,YF89,YF90,YF91,YF92,YF93,YF94,YF95,YF96,YF97,YF98,YF99,YF100,YF101,YF102,YF103,YF104,YF105,YF106,YF107,YF108,YF109,YF110,YF111,YF112,YF113,YF114,YF115,YF116,YF117,YF118,YF119,YF120,YF121,YF122,YF123,YF124,YF125,YF126,YF127,YF128,YF129,YF130,YF131,YF132,YF133,YF134,YF135,YF136,YF137,YF138,YF139,YF140,YF141,YF142,YF143,YF144,YF145,YF146,YF147,YF148,YF149,YF150,YF151,YF152,YF153,YF154,YF155,YF156,YF157,YF158,YF159,YF160,YF161,YF162,YF163,YF164,YF165,YF166,YF167,YF168,YF169,YF170,YF171,YF172,YF173,YF174,YF175,YF176,YF177,YF178,YF179,YF180,YF181,YF182,YF183,YF184,YF185,YF186,YF187,YF188,YF189,YF190,YF191,YF192,YF193,YF194,YF195,YF196,YF197,YF198,YF199,YF200,YF201,YF202,YF203,YF204,YF205,YF206,YF207,YF208,YF209,YF210,YF211,YF212,YF213,YF214,YF215,YF216,YF217,YF218,YF219,YF220,YF221,YF222,YF223,YF224,YF225,YF226,YF227,YF228,YF229,YF230,YF231,YF232,YF233,YF234,YF235,YF236,YF237,YF238,YF239,YF240,YF241,YF242,YF243,YF244,YF245,YF246,YF247,YF248,YF249,YF250,YF251,YF252,YF253,YF254,YF255);
input A0;
input A0_inv;
input A1;
input A1_inv;
input A2;
input A2_inv;
input A3;
input A3_inv;
input A4;
input A4_inv;
input A5;
input A5_inv;
input A6;
input A6_inv;
input A7;
input A7_inv;
input CLK;
output YF0;
output YF1;
output YF2;
output YF3;
output YF4;
output YF5;
output YF6;
output YF7;
output YF8;
output YF9;
output YF10;
output YF11;
output YF12;
output YF13;
output YF14;
output YF15;
output YF16;
output YF17;
output YF18;
output YF19;
output YF20;
output YF21;
output YF22;
output YF23;
output YF24;
output YF25;
output YF26;
output YF27;
output YF28;
output YF29;
output YF30;
output YF31;
output YF32;
output YF33;
output YF34;
output YF35;
output YF36;
output YF37;
output YF38;
output YF39;
output YF40;
output YF41;
output YF42;
output YF43;
output YF44;
output YF45;
output YF46;
output YF47;
output YF48;
output YF49;
output YF50;
output YF51;
output YF52;
output YF53;
output YF54;
output YF55;
output YF56;
output YF57;
output YF58;
output YF59;
output YF60;
output YF61;
output YF62;
output YF63;
output YF64;
output YF65;
output YF66;
output YF67;
output YF68;
output YF69;
output YF70;
output YF71;
output YF72;
output YF73;
output YF74;
output YF75;
output YF76;
output YF77;
output YF78;
output YF79;
output YF80;
output YF81;
output YF82;
output YF83;
output YF84;
output YF85;
output YF86;
output YF87;
output YF88;
output YF89;
output YF90;
output YF91;
output YF92;
output YF93;
output YF94;
output YF95;
output YF96;
output YF97;
output YF98;
output YF99;
output YF100;
output YF101;
output YF102;
output YF103;
output YF104;
output YF105;
output YF106;
output YF107;
output YF108;
output YF109;
output YF110;
output YF111;
output YF112;
output YF113;
output YF114;
output YF115;
output YF116;
output YF117;
output YF118;
output YF119;
output YF120;
output YF121;
output YF122;
output YF123;
output YF124;
output YF125;
output YF126;
output YF127;
output YF128;
output YF129;
output YF130;
output YF131;
output YF132;
output YF133;
output YF134;
output YF135;
output YF136;
output YF137;
output YF138;
output YF139;
output YF140;
output YF141;
output YF142;
output YF143;
output YF144;
output YF145;
output YF146;
output YF147;
output YF148;
output YF149;
output YF150;
output YF151;
output YF152;
output YF153;
output YF154;
output YF155;
output YF156;
output YF157;
output YF158;
output YF159;
output YF160;
output YF161;
output YF162;
output YF163;
output YF164;
output YF165;
output YF166;
output YF167;
output YF168;
output YF169;
output YF170;
output YF171;
output YF172;
output YF173;
output YF174;
output YF175;
output YF176;
output YF177;
output YF178;
output YF179;
output YF180;
output YF181;
output YF182;
output YF183;
output YF184;
output YF185;
output YF186;
output YF187;
output YF188;
output YF189;
output YF190;
output YF191;
output YF192;
output YF193;
output YF194;
output YF195;
output YF196;
output YF197;
output YF198;
output YF199;
output YF200;
output YF201;
output YF202;
output YF203;
output YF204;
output YF205;
output YF206;
output YF207;
output YF208;
output YF209;
output YF210;
output YF211;
output YF212;
output YF213;
output YF214;
output YF215;
output YF216;
output YF217;
output YF218;
output YF219;
output YF220;
output YF221;
output YF222;
output YF223;
output YF224;
output YF225;
output YF226;
output YF227;
output YF228;
output YF229;
output YF230;
output YF231;
output YF232;
output YF233;
output YF234;
output YF235;
output YF236;
output YF237;
output YF238;
output YF239;
output YF240;
output YF241;
output YF242;
output YF243;
output YF244;
output YF245;
output YF246;
output YF247;
output YF248;
output YF249;
output YF250;
output YF251;
output YF252;
output YF253;
output YF254;
output YF255;
NANDC2x1 inst_and_b0_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire0_0_0));
INVC inst_inv_b0_0_0 (.A(imd_wire0_0_0),.Y(wire0_0_0));
NANDC2x1 inst_and_b0_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire0_0_1));
INVC inst_inv_b0_0_1 (.A(imd_wire0_0_1),.Y(wire0_0_1));
NANDC2x1 inst_and_b0_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire0_0_2));
INVC inst_inv_b0_0_2 (.A(imd_wire0_0_2),.Y(wire0_0_2));
NANDC2x1 inst_and_b0_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire0_0_3));
INVC inst_inv_b0_0_3 (.A(imd_wire0_0_3),.Y(wire0_0_3));
NANDC2x1 inst_and_b0_1_0 (.A(wire0_0_0),.B(wire0_0_1),.Y(imd_wire0_1_0));
INVC inst_inv_b0_1_0 (.A(imd_wire0_1_0),.Y(wire0_1_0));
NANDC2x1 inst_and_b0_1_1 (.A(wire0_0_2),.B(wire0_0_3),.Y(imd_wire0_1_1));
INVC inst_inv_b0_1_1 (.A(imd_wire0_1_1),.Y(wire0_1_1));
NANDC2x1 inst_and_b0_2_0 (.A(wire0_1_0),.B(wire0_1_1),.Y(imd_Y0));
INVC inst_inv_b0_2_0 (.A(imd_Y0),.Y(Y0));
NANDC2x1 inst_clockedAND_b0_0 (.A(CLK),.B(Y0),.Y(imd_YF0));
INVC inst_clockedinv_b0_0 (.A(imd_YF0),.Y(YF0));


NANDC2x1 inst_and_b1_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire1_0_0));
INVC inst_inv_b1_0_0 (.A(imd_wire1_0_0),.Y(wire1_0_0));
NANDC2x1 inst_and_b1_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire1_0_1));
INVC inst_inv_b1_0_1 (.A(imd_wire1_0_1),.Y(wire1_0_1));
NANDC2x1 inst_and_b1_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire1_0_2));
INVC inst_inv_b1_0_2 (.A(imd_wire1_0_2),.Y(wire1_0_2));
NANDC2x1 inst_and_b1_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire1_0_3));
INVC inst_inv_b1_0_3 (.A(imd_wire1_0_3),.Y(wire1_0_3));
NANDC2x1 inst_and_b1_1_0 (.A(wire1_0_0),.B(wire1_0_1),.Y(imd_wire1_1_0));
INVC inst_inv_b1_1_0 (.A(imd_wire1_1_0),.Y(wire1_1_0));
NANDC2x1 inst_and_b1_1_1 (.A(wire1_0_2),.B(wire1_0_3),.Y(imd_wire1_1_1));
INVC inst_inv_b1_1_1 (.A(imd_wire1_1_1),.Y(wire1_1_1));
NANDC2x1 inst_and_b1_2_0 (.A(wire1_1_0),.B(wire1_1_1),.Y(imd_Y1));
INVC inst_inv_b1_2_0 (.A(imd_Y1),.Y(Y1));
NANDC2x1 inst_clockedAND_b1_1 (.A(CLK),.B(Y1),.Y(imd_YF1));
INVC inst_clockedinv_b1_1 (.A(imd_YF1),.Y(YF1));


NANDC2x1 inst_and_b2_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire2_0_0));
INVC inst_inv_b2_0_0 (.A(imd_wire2_0_0),.Y(wire2_0_0));
NANDC2x1 inst_and_b2_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire2_0_1));
INVC inst_inv_b2_0_1 (.A(imd_wire2_0_1),.Y(wire2_0_1));
NANDC2x1 inst_and_b2_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire2_0_2));
INVC inst_inv_b2_0_2 (.A(imd_wire2_0_2),.Y(wire2_0_2));
NANDC2x1 inst_and_b2_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire2_0_3));
INVC inst_inv_b2_0_3 (.A(imd_wire2_0_3),.Y(wire2_0_3));
NANDC2x1 inst_and_b2_1_0 (.A(wire2_0_0),.B(wire2_0_1),.Y(imd_wire2_1_0));
INVC inst_inv_b2_1_0 (.A(imd_wire2_1_0),.Y(wire2_1_0));
NANDC2x1 inst_and_b2_1_1 (.A(wire2_0_2),.B(wire2_0_3),.Y(imd_wire2_1_1));
INVC inst_inv_b2_1_1 (.A(imd_wire2_1_1),.Y(wire2_1_1));
NANDC2x1 inst_and_b2_2_0 (.A(wire2_1_0),.B(wire2_1_1),.Y(imd_Y2));
INVC inst_inv_b2_2_0 (.A(imd_Y2),.Y(Y2));
NANDC2x1 inst_clockedAND_b2_2 (.A(CLK),.B(Y2),.Y(imd_YF2));
INVC inst_clockedinv_b2_2 (.A(imd_YF2),.Y(YF2));


NANDC2x1 inst_and_b3_0_0 (.A(A0),.B(A1),.Y(imd_wire3_0_0));
INVC inst_inv_b3_0_0 (.A(imd_wire3_0_0),.Y(wire3_0_0));
NANDC2x1 inst_and_b3_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire3_0_1));
INVC inst_inv_b3_0_1 (.A(imd_wire3_0_1),.Y(wire3_0_1));
NANDC2x1 inst_and_b3_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire3_0_2));
INVC inst_inv_b3_0_2 (.A(imd_wire3_0_2),.Y(wire3_0_2));
NANDC2x1 inst_and_b3_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire3_0_3));
INVC inst_inv_b3_0_3 (.A(imd_wire3_0_3),.Y(wire3_0_3));
NANDC2x1 inst_and_b3_1_0 (.A(wire3_0_0),.B(wire3_0_1),.Y(imd_wire3_1_0));
INVC inst_inv_b3_1_0 (.A(imd_wire3_1_0),.Y(wire3_1_0));
NANDC2x1 inst_and_b3_1_1 (.A(wire3_0_2),.B(wire3_0_3),.Y(imd_wire3_1_1));
INVC inst_inv_b3_1_1 (.A(imd_wire3_1_1),.Y(wire3_1_1));
NANDC2x1 inst_and_b3_2_0 (.A(wire3_1_0),.B(wire3_1_1),.Y(imd_Y3));
INVC inst_inv_b3_2_0 (.A(imd_Y3),.Y(Y3));
NANDC2x1 inst_clockedAND_b3_3 (.A(CLK),.B(Y3),.Y(imd_YF3));
INVC inst_clockedinv_b3_3 (.A(imd_YF3),.Y(YF3));


NANDC2x1 inst_and_b4_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire4_0_0));
INVC inst_inv_b4_0_0 (.A(imd_wire4_0_0),.Y(wire4_0_0));
NANDC2x1 inst_and_b4_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire4_0_1));
INVC inst_inv_b4_0_1 (.A(imd_wire4_0_1),.Y(wire4_0_1));
NANDC2x1 inst_and_b4_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire4_0_2));
INVC inst_inv_b4_0_2 (.A(imd_wire4_0_2),.Y(wire4_0_2));
NANDC2x1 inst_and_b4_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire4_0_3));
INVC inst_inv_b4_0_3 (.A(imd_wire4_0_3),.Y(wire4_0_3));
NANDC2x1 inst_and_b4_1_0 (.A(wire4_0_0),.B(wire4_0_1),.Y(imd_wire4_1_0));
INVC inst_inv_b4_1_0 (.A(imd_wire4_1_0),.Y(wire4_1_0));
NANDC2x1 inst_and_b4_1_1 (.A(wire4_0_2),.B(wire4_0_3),.Y(imd_wire4_1_1));
INVC inst_inv_b4_1_1 (.A(imd_wire4_1_1),.Y(wire4_1_1));
NANDC2x1 inst_and_b4_2_0 (.A(wire4_1_0),.B(wire4_1_1),.Y(imd_Y4));
INVC inst_inv_b4_2_0 (.A(imd_Y4),.Y(Y4));
NANDC2x1 inst_clockedAND_b4_4 (.A(CLK),.B(Y4),.Y(imd_YF4));
INVC inst_clockedinv_b4_4 (.A(imd_YF4),.Y(YF4));


NANDC2x1 inst_and_b5_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire5_0_0));
INVC inst_inv_b5_0_0 (.A(imd_wire5_0_0),.Y(wire5_0_0));
NANDC2x1 inst_and_b5_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire5_0_1));
INVC inst_inv_b5_0_1 (.A(imd_wire5_0_1),.Y(wire5_0_1));
NANDC2x1 inst_and_b5_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire5_0_2));
INVC inst_inv_b5_0_2 (.A(imd_wire5_0_2),.Y(wire5_0_2));
NANDC2x1 inst_and_b5_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire5_0_3));
INVC inst_inv_b5_0_3 (.A(imd_wire5_0_3),.Y(wire5_0_3));
NANDC2x1 inst_and_b5_1_0 (.A(wire5_0_0),.B(wire5_0_1),.Y(imd_wire5_1_0));
INVC inst_inv_b5_1_0 (.A(imd_wire5_1_0),.Y(wire5_1_0));
NANDC2x1 inst_and_b5_1_1 (.A(wire5_0_2),.B(wire5_0_3),.Y(imd_wire5_1_1));
INVC inst_inv_b5_1_1 (.A(imd_wire5_1_1),.Y(wire5_1_1));
NANDC2x1 inst_and_b5_2_0 (.A(wire5_1_0),.B(wire5_1_1),.Y(imd_Y5));
INVC inst_inv_b5_2_0 (.A(imd_Y5),.Y(Y5));
NANDC2x1 inst_clockedAND_b5_5 (.A(CLK),.B(Y5),.Y(imd_YF5));
INVC inst_clockedinv_b5_5 (.A(imd_YF5),.Y(YF5));


NANDC2x1 inst_and_b6_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire6_0_0));
INVC inst_inv_b6_0_0 (.A(imd_wire6_0_0),.Y(wire6_0_0));
NANDC2x1 inst_and_b6_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire6_0_1));
INVC inst_inv_b6_0_1 (.A(imd_wire6_0_1),.Y(wire6_0_1));
NANDC2x1 inst_and_b6_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire6_0_2));
INVC inst_inv_b6_0_2 (.A(imd_wire6_0_2),.Y(wire6_0_2));
NANDC2x1 inst_and_b6_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire6_0_3));
INVC inst_inv_b6_0_3 (.A(imd_wire6_0_3),.Y(wire6_0_3));
NANDC2x1 inst_and_b6_1_0 (.A(wire6_0_0),.B(wire6_0_1),.Y(imd_wire6_1_0));
INVC inst_inv_b6_1_0 (.A(imd_wire6_1_0),.Y(wire6_1_0));
NANDC2x1 inst_and_b6_1_1 (.A(wire6_0_2),.B(wire6_0_3),.Y(imd_wire6_1_1));
INVC inst_inv_b6_1_1 (.A(imd_wire6_1_1),.Y(wire6_1_1));
NANDC2x1 inst_and_b6_2_0 (.A(wire6_1_0),.B(wire6_1_1),.Y(imd_Y6));
INVC inst_inv_b6_2_0 (.A(imd_Y6),.Y(Y6));
NANDC2x1 inst_clockedAND_b6_6 (.A(CLK),.B(Y6),.Y(imd_YF6));
INVC inst_clockedinv_b6_6 (.A(imd_YF6),.Y(YF6));


NANDC2x1 inst_and_b7_0_0 (.A(A0),.B(A1),.Y(imd_wire7_0_0));
INVC inst_inv_b7_0_0 (.A(imd_wire7_0_0),.Y(wire7_0_0));
NANDC2x1 inst_and_b7_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire7_0_1));
INVC inst_inv_b7_0_1 (.A(imd_wire7_0_1),.Y(wire7_0_1));
NANDC2x1 inst_and_b7_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire7_0_2));
INVC inst_inv_b7_0_2 (.A(imd_wire7_0_2),.Y(wire7_0_2));
NANDC2x1 inst_and_b7_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire7_0_3));
INVC inst_inv_b7_0_3 (.A(imd_wire7_0_3),.Y(wire7_0_3));
NANDC2x1 inst_and_b7_1_0 (.A(wire7_0_0),.B(wire7_0_1),.Y(imd_wire7_1_0));
INVC inst_inv_b7_1_0 (.A(imd_wire7_1_0),.Y(wire7_1_0));
NANDC2x1 inst_and_b7_1_1 (.A(wire7_0_2),.B(wire7_0_3),.Y(imd_wire7_1_1));
INVC inst_inv_b7_1_1 (.A(imd_wire7_1_1),.Y(wire7_1_1));
NANDC2x1 inst_and_b7_2_0 (.A(wire7_1_0),.B(wire7_1_1),.Y(imd_Y7));
INVC inst_inv_b7_2_0 (.A(imd_Y7),.Y(Y7));
NANDC2x1 inst_clockedAND_b7_7 (.A(CLK),.B(Y7),.Y(imd_YF7));
INVC inst_clockedinv_b7_7 (.A(imd_YF7),.Y(YF7));


NANDC2x1 inst_and_b8_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire8_0_0));
INVC inst_inv_b8_0_0 (.A(imd_wire8_0_0),.Y(wire8_0_0));
NANDC2x1 inst_and_b8_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire8_0_1));
INVC inst_inv_b8_0_1 (.A(imd_wire8_0_1),.Y(wire8_0_1));
NANDC2x1 inst_and_b8_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire8_0_2));
INVC inst_inv_b8_0_2 (.A(imd_wire8_0_2),.Y(wire8_0_2));
NANDC2x1 inst_and_b8_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire8_0_3));
INVC inst_inv_b8_0_3 (.A(imd_wire8_0_3),.Y(wire8_0_3));
NANDC2x1 inst_and_b8_1_0 (.A(wire8_0_0),.B(wire8_0_1),.Y(imd_wire8_1_0));
INVC inst_inv_b8_1_0 (.A(imd_wire8_1_0),.Y(wire8_1_0));
NANDC2x1 inst_and_b8_1_1 (.A(wire8_0_2),.B(wire8_0_3),.Y(imd_wire8_1_1));
INVC inst_inv_b8_1_1 (.A(imd_wire8_1_1),.Y(wire8_1_1));
NANDC2x1 inst_and_b8_2_0 (.A(wire8_1_0),.B(wire8_1_1),.Y(imd_Y8));
INVC inst_inv_b8_2_0 (.A(imd_Y8),.Y(Y8));
NANDC2x1 inst_clockedAND_b8_8 (.A(CLK),.B(Y8),.Y(imd_YF8));
INVC inst_clockedinv_b8_8 (.A(imd_YF8),.Y(YF8));


NANDC2x1 inst_and_b9_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire9_0_0));
INVC inst_inv_b9_0_0 (.A(imd_wire9_0_0),.Y(wire9_0_0));
NANDC2x1 inst_and_b9_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire9_0_1));
INVC inst_inv_b9_0_1 (.A(imd_wire9_0_1),.Y(wire9_0_1));
NANDC2x1 inst_and_b9_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire9_0_2));
INVC inst_inv_b9_0_2 (.A(imd_wire9_0_2),.Y(wire9_0_2));
NANDC2x1 inst_and_b9_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire9_0_3));
INVC inst_inv_b9_0_3 (.A(imd_wire9_0_3),.Y(wire9_0_3));
NANDC2x1 inst_and_b9_1_0 (.A(wire9_0_0),.B(wire9_0_1),.Y(imd_wire9_1_0));
INVC inst_inv_b9_1_0 (.A(imd_wire9_1_0),.Y(wire9_1_0));
NANDC2x1 inst_and_b9_1_1 (.A(wire9_0_2),.B(wire9_0_3),.Y(imd_wire9_1_1));
INVC inst_inv_b9_1_1 (.A(imd_wire9_1_1),.Y(wire9_1_1));
NANDC2x1 inst_and_b9_2_0 (.A(wire9_1_0),.B(wire9_1_1),.Y(imd_Y9));
INVC inst_inv_b9_2_0 (.A(imd_Y9),.Y(Y9));
NANDC2x1 inst_clockedAND_b9_9 (.A(CLK),.B(Y9),.Y(imd_YF9));
INVC inst_clockedinv_b9_9 (.A(imd_YF9),.Y(YF9));


NANDC2x1 inst_and_b10_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire10_0_0));
INVC inst_inv_b10_0_0 (.A(imd_wire10_0_0),.Y(wire10_0_0));
NANDC2x1 inst_and_b10_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire10_0_1));
INVC inst_inv_b10_0_1 (.A(imd_wire10_0_1),.Y(wire10_0_1));
NANDC2x1 inst_and_b10_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire10_0_2));
INVC inst_inv_b10_0_2 (.A(imd_wire10_0_2),.Y(wire10_0_2));
NANDC2x1 inst_and_b10_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire10_0_3));
INVC inst_inv_b10_0_3 (.A(imd_wire10_0_3),.Y(wire10_0_3));
NANDC2x1 inst_and_b10_1_0 (.A(wire10_0_0),.B(wire10_0_1),.Y(imd_wire10_1_0));
INVC inst_inv_b10_1_0 (.A(imd_wire10_1_0),.Y(wire10_1_0));
NANDC2x1 inst_and_b10_1_1 (.A(wire10_0_2),.B(wire10_0_3),.Y(imd_wire10_1_1));
INVC inst_inv_b10_1_1 (.A(imd_wire10_1_1),.Y(wire10_1_1));
NANDC2x1 inst_and_b10_2_0 (.A(wire10_1_0),.B(wire10_1_1),.Y(imd_Y10));
INVC inst_inv_b10_2_0 (.A(imd_Y10),.Y(Y10));
NANDC2x1 inst_clockedAND_b10_10 (.A(CLK),.B(Y10),.Y(imd_YF10));
INVC inst_clockedinv_b10_10 (.A(imd_YF10),.Y(YF10));


NANDC2x1 inst_and_b11_0_0 (.A(A0),.B(A1),.Y(imd_wire11_0_0));
INVC inst_inv_b11_0_0 (.A(imd_wire11_0_0),.Y(wire11_0_0));
NANDC2x1 inst_and_b11_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire11_0_1));
INVC inst_inv_b11_0_1 (.A(imd_wire11_0_1),.Y(wire11_0_1));
NANDC2x1 inst_and_b11_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire11_0_2));
INVC inst_inv_b11_0_2 (.A(imd_wire11_0_2),.Y(wire11_0_2));
NANDC2x1 inst_and_b11_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire11_0_3));
INVC inst_inv_b11_0_3 (.A(imd_wire11_0_3),.Y(wire11_0_3));
NANDC2x1 inst_and_b11_1_0 (.A(wire11_0_0),.B(wire11_0_1),.Y(imd_wire11_1_0));
INVC inst_inv_b11_1_0 (.A(imd_wire11_1_0),.Y(wire11_1_0));
NANDC2x1 inst_and_b11_1_1 (.A(wire11_0_2),.B(wire11_0_3),.Y(imd_wire11_1_1));
INVC inst_inv_b11_1_1 (.A(imd_wire11_1_1),.Y(wire11_1_1));
NANDC2x1 inst_and_b11_2_0 (.A(wire11_1_0),.B(wire11_1_1),.Y(imd_Y11));
INVC inst_inv_b11_2_0 (.A(imd_Y11),.Y(Y11));
NANDC2x1 inst_clockedAND_b11_11 (.A(CLK),.B(Y11),.Y(imd_YF11));
INVC inst_clockedinv_b11_11 (.A(imd_YF11),.Y(YF11));


NANDC2x1 inst_and_b12_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire12_0_0));
INVC inst_inv_b12_0_0 (.A(imd_wire12_0_0),.Y(wire12_0_0));
NANDC2x1 inst_and_b12_0_1 (.A(A2),.B(A3),.Y(imd_wire12_0_1));
INVC inst_inv_b12_0_1 (.A(imd_wire12_0_1),.Y(wire12_0_1));
NANDC2x1 inst_and_b12_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire12_0_2));
INVC inst_inv_b12_0_2 (.A(imd_wire12_0_2),.Y(wire12_0_2));
NANDC2x1 inst_and_b12_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire12_0_3));
INVC inst_inv_b12_0_3 (.A(imd_wire12_0_3),.Y(wire12_0_3));
NANDC2x1 inst_and_b12_1_0 (.A(wire12_0_0),.B(wire12_0_1),.Y(imd_wire12_1_0));
INVC inst_inv_b12_1_0 (.A(imd_wire12_1_0),.Y(wire12_1_0));
NANDC2x1 inst_and_b12_1_1 (.A(wire12_0_2),.B(wire12_0_3),.Y(imd_wire12_1_1));
INVC inst_inv_b12_1_1 (.A(imd_wire12_1_1),.Y(wire12_1_1));
NANDC2x1 inst_and_b12_2_0 (.A(wire12_1_0),.B(wire12_1_1),.Y(imd_Y12));
INVC inst_inv_b12_2_0 (.A(imd_Y12),.Y(Y12));
NANDC2x1 inst_clockedAND_b12_12 (.A(CLK),.B(Y12),.Y(imd_YF12));
INVC inst_clockedinv_b12_12 (.A(imd_YF12),.Y(YF12));


NANDC2x1 inst_and_b13_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire13_0_0));
INVC inst_inv_b13_0_0 (.A(imd_wire13_0_0),.Y(wire13_0_0));
NANDC2x1 inst_and_b13_0_1 (.A(A2),.B(A3),.Y(imd_wire13_0_1));
INVC inst_inv_b13_0_1 (.A(imd_wire13_0_1),.Y(wire13_0_1));
NANDC2x1 inst_and_b13_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire13_0_2));
INVC inst_inv_b13_0_2 (.A(imd_wire13_0_2),.Y(wire13_0_2));
NANDC2x1 inst_and_b13_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire13_0_3));
INVC inst_inv_b13_0_3 (.A(imd_wire13_0_3),.Y(wire13_0_3));
NANDC2x1 inst_and_b13_1_0 (.A(wire13_0_0),.B(wire13_0_1),.Y(imd_wire13_1_0));
INVC inst_inv_b13_1_0 (.A(imd_wire13_1_0),.Y(wire13_1_0));
NANDC2x1 inst_and_b13_1_1 (.A(wire13_0_2),.B(wire13_0_3),.Y(imd_wire13_1_1));
INVC inst_inv_b13_1_1 (.A(imd_wire13_1_1),.Y(wire13_1_1));
NANDC2x1 inst_and_b13_2_0 (.A(wire13_1_0),.B(wire13_1_1),.Y(imd_Y13));
INVC inst_inv_b13_2_0 (.A(imd_Y13),.Y(Y13));
NANDC2x1 inst_clockedAND_b13_13 (.A(CLK),.B(Y13),.Y(imd_YF13));
INVC inst_clockedinv_b13_13 (.A(imd_YF13),.Y(YF13));


NANDC2x1 inst_and_b14_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire14_0_0));
INVC inst_inv_b14_0_0 (.A(imd_wire14_0_0),.Y(wire14_0_0));
NANDC2x1 inst_and_b14_0_1 (.A(A2),.B(A3),.Y(imd_wire14_0_1));
INVC inst_inv_b14_0_1 (.A(imd_wire14_0_1),.Y(wire14_0_1));
NANDC2x1 inst_and_b14_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire14_0_2));
INVC inst_inv_b14_0_2 (.A(imd_wire14_0_2),.Y(wire14_0_2));
NANDC2x1 inst_and_b14_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire14_0_3));
INVC inst_inv_b14_0_3 (.A(imd_wire14_0_3),.Y(wire14_0_3));
NANDC2x1 inst_and_b14_1_0 (.A(wire14_0_0),.B(wire14_0_1),.Y(imd_wire14_1_0));
INVC inst_inv_b14_1_0 (.A(imd_wire14_1_0),.Y(wire14_1_0));
NANDC2x1 inst_and_b14_1_1 (.A(wire14_0_2),.B(wire14_0_3),.Y(imd_wire14_1_1));
INVC inst_inv_b14_1_1 (.A(imd_wire14_1_1),.Y(wire14_1_1));
NANDC2x1 inst_and_b14_2_0 (.A(wire14_1_0),.B(wire14_1_1),.Y(imd_Y14));
INVC inst_inv_b14_2_0 (.A(imd_Y14),.Y(Y14));
NANDC2x1 inst_clockedAND_b14_14 (.A(CLK),.B(Y14),.Y(imd_YF14));
INVC inst_clockedinv_b14_14 (.A(imd_YF14),.Y(YF14));


NANDC2x1 inst_and_b15_0_0 (.A(A0),.B(A1),.Y(imd_wire15_0_0));
INVC inst_inv_b15_0_0 (.A(imd_wire15_0_0),.Y(wire15_0_0));
NANDC2x1 inst_and_b15_0_1 (.A(A2),.B(A3),.Y(imd_wire15_0_1));
INVC inst_inv_b15_0_1 (.A(imd_wire15_0_1),.Y(wire15_0_1));
NANDC2x1 inst_and_b15_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire15_0_2));
INVC inst_inv_b15_0_2 (.A(imd_wire15_0_2),.Y(wire15_0_2));
NANDC2x1 inst_and_b15_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire15_0_3));
INVC inst_inv_b15_0_3 (.A(imd_wire15_0_3),.Y(wire15_0_3));
NANDC2x1 inst_and_b15_1_0 (.A(wire15_0_0),.B(wire15_0_1),.Y(imd_wire15_1_0));
INVC inst_inv_b15_1_0 (.A(imd_wire15_1_0),.Y(wire15_1_0));
NANDC2x1 inst_and_b15_1_1 (.A(wire15_0_2),.B(wire15_0_3),.Y(imd_wire15_1_1));
INVC inst_inv_b15_1_1 (.A(imd_wire15_1_1),.Y(wire15_1_1));
NANDC2x1 inst_and_b15_2_0 (.A(wire15_1_0),.B(wire15_1_1),.Y(imd_Y15));
INVC inst_inv_b15_2_0 (.A(imd_Y15),.Y(Y15));
NANDC2x1 inst_clockedAND_b15_15 (.A(CLK),.B(Y15),.Y(imd_YF15));
INVC inst_clockedinv_b15_15 (.A(imd_YF15),.Y(YF15));


NANDC2x1 inst_and_b16_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire16_0_0));
INVC inst_inv_b16_0_0 (.A(imd_wire16_0_0),.Y(wire16_0_0));
NANDC2x1 inst_and_b16_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire16_0_1));
INVC inst_inv_b16_0_1 (.A(imd_wire16_0_1),.Y(wire16_0_1));
NANDC2x1 inst_and_b16_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire16_0_2));
INVC inst_inv_b16_0_2 (.A(imd_wire16_0_2),.Y(wire16_0_2));
NANDC2x1 inst_and_b16_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire16_0_3));
INVC inst_inv_b16_0_3 (.A(imd_wire16_0_3),.Y(wire16_0_3));
NANDC2x1 inst_and_b16_1_0 (.A(wire16_0_0),.B(wire16_0_1),.Y(imd_wire16_1_0));
INVC inst_inv_b16_1_0 (.A(imd_wire16_1_0),.Y(wire16_1_0));
NANDC2x1 inst_and_b16_1_1 (.A(wire16_0_2),.B(wire16_0_3),.Y(imd_wire16_1_1));
INVC inst_inv_b16_1_1 (.A(imd_wire16_1_1),.Y(wire16_1_1));
NANDC2x1 inst_and_b16_2_0 (.A(wire16_1_0),.B(wire16_1_1),.Y(imd_Y16));
INVC inst_inv_b16_2_0 (.A(imd_Y16),.Y(Y16));
NANDC2x1 inst_clockedAND_b16_16 (.A(CLK),.B(Y16),.Y(imd_YF16));
INVC inst_clockedinv_b16_16 (.A(imd_YF16),.Y(YF16));


NANDC2x1 inst_and_b17_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire17_0_0));
INVC inst_inv_b17_0_0 (.A(imd_wire17_0_0),.Y(wire17_0_0));
NANDC2x1 inst_and_b17_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire17_0_1));
INVC inst_inv_b17_0_1 (.A(imd_wire17_0_1),.Y(wire17_0_1));
NANDC2x1 inst_and_b17_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire17_0_2));
INVC inst_inv_b17_0_2 (.A(imd_wire17_0_2),.Y(wire17_0_2));
NANDC2x1 inst_and_b17_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire17_0_3));
INVC inst_inv_b17_0_3 (.A(imd_wire17_0_3),.Y(wire17_0_3));
NANDC2x1 inst_and_b17_1_0 (.A(wire17_0_0),.B(wire17_0_1),.Y(imd_wire17_1_0));
INVC inst_inv_b17_1_0 (.A(imd_wire17_1_0),.Y(wire17_1_0));
NANDC2x1 inst_and_b17_1_1 (.A(wire17_0_2),.B(wire17_0_3),.Y(imd_wire17_1_1));
INVC inst_inv_b17_1_1 (.A(imd_wire17_1_1),.Y(wire17_1_1));
NANDC2x1 inst_and_b17_2_0 (.A(wire17_1_0),.B(wire17_1_1),.Y(imd_Y17));
INVC inst_inv_b17_2_0 (.A(imd_Y17),.Y(Y17));
NANDC2x1 inst_clockedAND_b17_17 (.A(CLK),.B(Y17),.Y(imd_YF17));
INVC inst_clockedinv_b17_17 (.A(imd_YF17),.Y(YF17));


NANDC2x1 inst_and_b18_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire18_0_0));
INVC inst_inv_b18_0_0 (.A(imd_wire18_0_0),.Y(wire18_0_0));
NANDC2x1 inst_and_b18_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire18_0_1));
INVC inst_inv_b18_0_1 (.A(imd_wire18_0_1),.Y(wire18_0_1));
NANDC2x1 inst_and_b18_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire18_0_2));
INVC inst_inv_b18_0_2 (.A(imd_wire18_0_2),.Y(wire18_0_2));
NANDC2x1 inst_and_b18_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire18_0_3));
INVC inst_inv_b18_0_3 (.A(imd_wire18_0_3),.Y(wire18_0_3));
NANDC2x1 inst_and_b18_1_0 (.A(wire18_0_0),.B(wire18_0_1),.Y(imd_wire18_1_0));
INVC inst_inv_b18_1_0 (.A(imd_wire18_1_0),.Y(wire18_1_0));
NANDC2x1 inst_and_b18_1_1 (.A(wire18_0_2),.B(wire18_0_3),.Y(imd_wire18_1_1));
INVC inst_inv_b18_1_1 (.A(imd_wire18_1_1),.Y(wire18_1_1));
NANDC2x1 inst_and_b18_2_0 (.A(wire18_1_0),.B(wire18_1_1),.Y(imd_Y18));
INVC inst_inv_b18_2_0 (.A(imd_Y18),.Y(Y18));
NANDC2x1 inst_clockedAND_b18_18 (.A(CLK),.B(Y18),.Y(imd_YF18));
INVC inst_clockedinv_b18_18 (.A(imd_YF18),.Y(YF18));


NANDC2x1 inst_and_b19_0_0 (.A(A0),.B(A1),.Y(imd_wire19_0_0));
INVC inst_inv_b19_0_0 (.A(imd_wire19_0_0),.Y(wire19_0_0));
NANDC2x1 inst_and_b19_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire19_0_1));
INVC inst_inv_b19_0_1 (.A(imd_wire19_0_1),.Y(wire19_0_1));
NANDC2x1 inst_and_b19_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire19_0_2));
INVC inst_inv_b19_0_2 (.A(imd_wire19_0_2),.Y(wire19_0_2));
NANDC2x1 inst_and_b19_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire19_0_3));
INVC inst_inv_b19_0_3 (.A(imd_wire19_0_3),.Y(wire19_0_3));
NANDC2x1 inst_and_b19_1_0 (.A(wire19_0_0),.B(wire19_0_1),.Y(imd_wire19_1_0));
INVC inst_inv_b19_1_0 (.A(imd_wire19_1_0),.Y(wire19_1_0));
NANDC2x1 inst_and_b19_1_1 (.A(wire19_0_2),.B(wire19_0_3),.Y(imd_wire19_1_1));
INVC inst_inv_b19_1_1 (.A(imd_wire19_1_1),.Y(wire19_1_1));
NANDC2x1 inst_and_b19_2_0 (.A(wire19_1_0),.B(wire19_1_1),.Y(imd_Y19));
INVC inst_inv_b19_2_0 (.A(imd_Y19),.Y(Y19));
NANDC2x1 inst_clockedAND_b19_19 (.A(CLK),.B(Y19),.Y(imd_YF19));
INVC inst_clockedinv_b19_19 (.A(imd_YF19),.Y(YF19));


NANDC2x1 inst_and_b20_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire20_0_0));
INVC inst_inv_b20_0_0 (.A(imd_wire20_0_0),.Y(wire20_0_0));
NANDC2x1 inst_and_b20_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire20_0_1));
INVC inst_inv_b20_0_1 (.A(imd_wire20_0_1),.Y(wire20_0_1));
NANDC2x1 inst_and_b20_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire20_0_2));
INVC inst_inv_b20_0_2 (.A(imd_wire20_0_2),.Y(wire20_0_2));
NANDC2x1 inst_and_b20_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire20_0_3));
INVC inst_inv_b20_0_3 (.A(imd_wire20_0_3),.Y(wire20_0_3));
NANDC2x1 inst_and_b20_1_0 (.A(wire20_0_0),.B(wire20_0_1),.Y(imd_wire20_1_0));
INVC inst_inv_b20_1_0 (.A(imd_wire20_1_0),.Y(wire20_1_0));
NANDC2x1 inst_and_b20_1_1 (.A(wire20_0_2),.B(wire20_0_3),.Y(imd_wire20_1_1));
INVC inst_inv_b20_1_1 (.A(imd_wire20_1_1),.Y(wire20_1_1));
NANDC2x1 inst_and_b20_2_0 (.A(wire20_1_0),.B(wire20_1_1),.Y(imd_Y20));
INVC inst_inv_b20_2_0 (.A(imd_Y20),.Y(Y20));
NANDC2x1 inst_clockedAND_b20_20 (.A(CLK),.B(Y20),.Y(imd_YF20));
INVC inst_clockedinv_b20_20 (.A(imd_YF20),.Y(YF20));


NANDC2x1 inst_and_b21_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire21_0_0));
INVC inst_inv_b21_0_0 (.A(imd_wire21_0_0),.Y(wire21_0_0));
NANDC2x1 inst_and_b21_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire21_0_1));
INVC inst_inv_b21_0_1 (.A(imd_wire21_0_1),.Y(wire21_0_1));
NANDC2x1 inst_and_b21_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire21_0_2));
INVC inst_inv_b21_0_2 (.A(imd_wire21_0_2),.Y(wire21_0_2));
NANDC2x1 inst_and_b21_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire21_0_3));
INVC inst_inv_b21_0_3 (.A(imd_wire21_0_3),.Y(wire21_0_3));
NANDC2x1 inst_and_b21_1_0 (.A(wire21_0_0),.B(wire21_0_1),.Y(imd_wire21_1_0));
INVC inst_inv_b21_1_0 (.A(imd_wire21_1_0),.Y(wire21_1_0));
NANDC2x1 inst_and_b21_1_1 (.A(wire21_0_2),.B(wire21_0_3),.Y(imd_wire21_1_1));
INVC inst_inv_b21_1_1 (.A(imd_wire21_1_1),.Y(wire21_1_1));
NANDC2x1 inst_and_b21_2_0 (.A(wire21_1_0),.B(wire21_1_1),.Y(imd_Y21));
INVC inst_inv_b21_2_0 (.A(imd_Y21),.Y(Y21));
NANDC2x1 inst_clockedAND_b21_21 (.A(CLK),.B(Y21),.Y(imd_YF21));
INVC inst_clockedinv_b21_21 (.A(imd_YF21),.Y(YF21));


NANDC2x1 inst_and_b22_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire22_0_0));
INVC inst_inv_b22_0_0 (.A(imd_wire22_0_0),.Y(wire22_0_0));
NANDC2x1 inst_and_b22_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire22_0_1));
INVC inst_inv_b22_0_1 (.A(imd_wire22_0_1),.Y(wire22_0_1));
NANDC2x1 inst_and_b22_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire22_0_2));
INVC inst_inv_b22_0_2 (.A(imd_wire22_0_2),.Y(wire22_0_2));
NANDC2x1 inst_and_b22_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire22_0_3));
INVC inst_inv_b22_0_3 (.A(imd_wire22_0_3),.Y(wire22_0_3));
NANDC2x1 inst_and_b22_1_0 (.A(wire22_0_0),.B(wire22_0_1),.Y(imd_wire22_1_0));
INVC inst_inv_b22_1_0 (.A(imd_wire22_1_0),.Y(wire22_1_0));
NANDC2x1 inst_and_b22_1_1 (.A(wire22_0_2),.B(wire22_0_3),.Y(imd_wire22_1_1));
INVC inst_inv_b22_1_1 (.A(imd_wire22_1_1),.Y(wire22_1_1));
NANDC2x1 inst_and_b22_2_0 (.A(wire22_1_0),.B(wire22_1_1),.Y(imd_Y22));
INVC inst_inv_b22_2_0 (.A(imd_Y22),.Y(Y22));
NANDC2x1 inst_clockedAND_b22_22 (.A(CLK),.B(Y22),.Y(imd_YF22));
INVC inst_clockedinv_b22_22 (.A(imd_YF22),.Y(YF22));


NANDC2x1 inst_and_b23_0_0 (.A(A0),.B(A1),.Y(imd_wire23_0_0));
INVC inst_inv_b23_0_0 (.A(imd_wire23_0_0),.Y(wire23_0_0));
NANDC2x1 inst_and_b23_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire23_0_1));
INVC inst_inv_b23_0_1 (.A(imd_wire23_0_1),.Y(wire23_0_1));
NANDC2x1 inst_and_b23_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire23_0_2));
INVC inst_inv_b23_0_2 (.A(imd_wire23_0_2),.Y(wire23_0_2));
NANDC2x1 inst_and_b23_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire23_0_3));
INVC inst_inv_b23_0_3 (.A(imd_wire23_0_3),.Y(wire23_0_3));
NANDC2x1 inst_and_b23_1_0 (.A(wire23_0_0),.B(wire23_0_1),.Y(imd_wire23_1_0));
INVC inst_inv_b23_1_0 (.A(imd_wire23_1_0),.Y(wire23_1_0));
NANDC2x1 inst_and_b23_1_1 (.A(wire23_0_2),.B(wire23_0_3),.Y(imd_wire23_1_1));
INVC inst_inv_b23_1_1 (.A(imd_wire23_1_1),.Y(wire23_1_1));
NANDC2x1 inst_and_b23_2_0 (.A(wire23_1_0),.B(wire23_1_1),.Y(imd_Y23));
INVC inst_inv_b23_2_0 (.A(imd_Y23),.Y(Y23));
NANDC2x1 inst_clockedAND_b23_23 (.A(CLK),.B(Y23),.Y(imd_YF23));
INVC inst_clockedinv_b23_23 (.A(imd_YF23),.Y(YF23));


NANDC2x1 inst_and_b24_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire24_0_0));
INVC inst_inv_b24_0_0 (.A(imd_wire24_0_0),.Y(wire24_0_0));
NANDC2x1 inst_and_b24_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire24_0_1));
INVC inst_inv_b24_0_1 (.A(imd_wire24_0_1),.Y(wire24_0_1));
NANDC2x1 inst_and_b24_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire24_0_2));
INVC inst_inv_b24_0_2 (.A(imd_wire24_0_2),.Y(wire24_0_2));
NANDC2x1 inst_and_b24_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire24_0_3));
INVC inst_inv_b24_0_3 (.A(imd_wire24_0_3),.Y(wire24_0_3));
NANDC2x1 inst_and_b24_1_0 (.A(wire24_0_0),.B(wire24_0_1),.Y(imd_wire24_1_0));
INVC inst_inv_b24_1_0 (.A(imd_wire24_1_0),.Y(wire24_1_0));
NANDC2x1 inst_and_b24_1_1 (.A(wire24_0_2),.B(wire24_0_3),.Y(imd_wire24_1_1));
INVC inst_inv_b24_1_1 (.A(imd_wire24_1_1),.Y(wire24_1_1));
NANDC2x1 inst_and_b24_2_0 (.A(wire24_1_0),.B(wire24_1_1),.Y(imd_Y24));
INVC inst_inv_b24_2_0 (.A(imd_Y24),.Y(Y24));
NANDC2x1 inst_clockedAND_b24_24 (.A(CLK),.B(Y24),.Y(imd_YF24));
INVC inst_clockedinv_b24_24 (.A(imd_YF24),.Y(YF24));


NANDC2x1 inst_and_b25_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire25_0_0));
INVC inst_inv_b25_0_0 (.A(imd_wire25_0_0),.Y(wire25_0_0));
NANDC2x1 inst_and_b25_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire25_0_1));
INVC inst_inv_b25_0_1 (.A(imd_wire25_0_1),.Y(wire25_0_1));
NANDC2x1 inst_and_b25_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire25_0_2));
INVC inst_inv_b25_0_2 (.A(imd_wire25_0_2),.Y(wire25_0_2));
NANDC2x1 inst_and_b25_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire25_0_3));
INVC inst_inv_b25_0_3 (.A(imd_wire25_0_3),.Y(wire25_0_3));
NANDC2x1 inst_and_b25_1_0 (.A(wire25_0_0),.B(wire25_0_1),.Y(imd_wire25_1_0));
INVC inst_inv_b25_1_0 (.A(imd_wire25_1_0),.Y(wire25_1_0));
NANDC2x1 inst_and_b25_1_1 (.A(wire25_0_2),.B(wire25_0_3),.Y(imd_wire25_1_1));
INVC inst_inv_b25_1_1 (.A(imd_wire25_1_1),.Y(wire25_1_1));
NANDC2x1 inst_and_b25_2_0 (.A(wire25_1_0),.B(wire25_1_1),.Y(imd_Y25));
INVC inst_inv_b25_2_0 (.A(imd_Y25),.Y(Y25));
NANDC2x1 inst_clockedAND_b25_25 (.A(CLK),.B(Y25),.Y(imd_YF25));
INVC inst_clockedinv_b25_25 (.A(imd_YF25),.Y(YF25));


NANDC2x1 inst_and_b26_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire26_0_0));
INVC inst_inv_b26_0_0 (.A(imd_wire26_0_0),.Y(wire26_0_0));
NANDC2x1 inst_and_b26_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire26_0_1));
INVC inst_inv_b26_0_1 (.A(imd_wire26_0_1),.Y(wire26_0_1));
NANDC2x1 inst_and_b26_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire26_0_2));
INVC inst_inv_b26_0_2 (.A(imd_wire26_0_2),.Y(wire26_0_2));
NANDC2x1 inst_and_b26_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire26_0_3));
INVC inst_inv_b26_0_3 (.A(imd_wire26_0_3),.Y(wire26_0_3));
NANDC2x1 inst_and_b26_1_0 (.A(wire26_0_0),.B(wire26_0_1),.Y(imd_wire26_1_0));
INVC inst_inv_b26_1_0 (.A(imd_wire26_1_0),.Y(wire26_1_0));
NANDC2x1 inst_and_b26_1_1 (.A(wire26_0_2),.B(wire26_0_3),.Y(imd_wire26_1_1));
INVC inst_inv_b26_1_1 (.A(imd_wire26_1_1),.Y(wire26_1_1));
NANDC2x1 inst_and_b26_2_0 (.A(wire26_1_0),.B(wire26_1_1),.Y(imd_Y26));
INVC inst_inv_b26_2_0 (.A(imd_Y26),.Y(Y26));
NANDC2x1 inst_clockedAND_b26_26 (.A(CLK),.B(Y26),.Y(imd_YF26));
INVC inst_clockedinv_b26_26 (.A(imd_YF26),.Y(YF26));


NANDC2x1 inst_and_b27_0_0 (.A(A0),.B(A1),.Y(imd_wire27_0_0));
INVC inst_inv_b27_0_0 (.A(imd_wire27_0_0),.Y(wire27_0_0));
NANDC2x1 inst_and_b27_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire27_0_1));
INVC inst_inv_b27_0_1 (.A(imd_wire27_0_1),.Y(wire27_0_1));
NANDC2x1 inst_and_b27_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire27_0_2));
INVC inst_inv_b27_0_2 (.A(imd_wire27_0_2),.Y(wire27_0_2));
NANDC2x1 inst_and_b27_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire27_0_3));
INVC inst_inv_b27_0_3 (.A(imd_wire27_0_3),.Y(wire27_0_3));
NANDC2x1 inst_and_b27_1_0 (.A(wire27_0_0),.B(wire27_0_1),.Y(imd_wire27_1_0));
INVC inst_inv_b27_1_0 (.A(imd_wire27_1_0),.Y(wire27_1_0));
NANDC2x1 inst_and_b27_1_1 (.A(wire27_0_2),.B(wire27_0_3),.Y(imd_wire27_1_1));
INVC inst_inv_b27_1_1 (.A(imd_wire27_1_1),.Y(wire27_1_1));
NANDC2x1 inst_and_b27_2_0 (.A(wire27_1_0),.B(wire27_1_1),.Y(imd_Y27));
INVC inst_inv_b27_2_0 (.A(imd_Y27),.Y(Y27));
NANDC2x1 inst_clockedAND_b27_27 (.A(CLK),.B(Y27),.Y(imd_YF27));
INVC inst_clockedinv_b27_27 (.A(imd_YF27),.Y(YF27));


NANDC2x1 inst_and_b28_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire28_0_0));
INVC inst_inv_b28_0_0 (.A(imd_wire28_0_0),.Y(wire28_0_0));
NANDC2x1 inst_and_b28_0_1 (.A(A2),.B(A3),.Y(imd_wire28_0_1));
INVC inst_inv_b28_0_1 (.A(imd_wire28_0_1),.Y(wire28_0_1));
NANDC2x1 inst_and_b28_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire28_0_2));
INVC inst_inv_b28_0_2 (.A(imd_wire28_0_2),.Y(wire28_0_2));
NANDC2x1 inst_and_b28_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire28_0_3));
INVC inst_inv_b28_0_3 (.A(imd_wire28_0_3),.Y(wire28_0_3));
NANDC2x1 inst_and_b28_1_0 (.A(wire28_0_0),.B(wire28_0_1),.Y(imd_wire28_1_0));
INVC inst_inv_b28_1_0 (.A(imd_wire28_1_0),.Y(wire28_1_0));
NANDC2x1 inst_and_b28_1_1 (.A(wire28_0_2),.B(wire28_0_3),.Y(imd_wire28_1_1));
INVC inst_inv_b28_1_1 (.A(imd_wire28_1_1),.Y(wire28_1_1));
NANDC2x1 inst_and_b28_2_0 (.A(wire28_1_0),.B(wire28_1_1),.Y(imd_Y28));
INVC inst_inv_b28_2_0 (.A(imd_Y28),.Y(Y28));
NANDC2x1 inst_clockedAND_b28_28 (.A(CLK),.B(Y28),.Y(imd_YF28));
INVC inst_clockedinv_b28_28 (.A(imd_YF28),.Y(YF28));


NANDC2x1 inst_and_b29_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire29_0_0));
INVC inst_inv_b29_0_0 (.A(imd_wire29_0_0),.Y(wire29_0_0));
NANDC2x1 inst_and_b29_0_1 (.A(A2),.B(A3),.Y(imd_wire29_0_1));
INVC inst_inv_b29_0_1 (.A(imd_wire29_0_1),.Y(wire29_0_1));
NANDC2x1 inst_and_b29_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire29_0_2));
INVC inst_inv_b29_0_2 (.A(imd_wire29_0_2),.Y(wire29_0_2));
NANDC2x1 inst_and_b29_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire29_0_3));
INVC inst_inv_b29_0_3 (.A(imd_wire29_0_3),.Y(wire29_0_3));
NANDC2x1 inst_and_b29_1_0 (.A(wire29_0_0),.B(wire29_0_1),.Y(imd_wire29_1_0));
INVC inst_inv_b29_1_0 (.A(imd_wire29_1_0),.Y(wire29_1_0));
NANDC2x1 inst_and_b29_1_1 (.A(wire29_0_2),.B(wire29_0_3),.Y(imd_wire29_1_1));
INVC inst_inv_b29_1_1 (.A(imd_wire29_1_1),.Y(wire29_1_1));
NANDC2x1 inst_and_b29_2_0 (.A(wire29_1_0),.B(wire29_1_1),.Y(imd_Y29));
INVC inst_inv_b29_2_0 (.A(imd_Y29),.Y(Y29));
NANDC2x1 inst_clockedAND_b29_29 (.A(CLK),.B(Y29),.Y(imd_YF29));
INVC inst_clockedinv_b29_29 (.A(imd_YF29),.Y(YF29));


NANDC2x1 inst_and_b30_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire30_0_0));
INVC inst_inv_b30_0_0 (.A(imd_wire30_0_0),.Y(wire30_0_0));
NANDC2x1 inst_and_b30_0_1 (.A(A2),.B(A3),.Y(imd_wire30_0_1));
INVC inst_inv_b30_0_1 (.A(imd_wire30_0_1),.Y(wire30_0_1));
NANDC2x1 inst_and_b30_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire30_0_2));
INVC inst_inv_b30_0_2 (.A(imd_wire30_0_2),.Y(wire30_0_2));
NANDC2x1 inst_and_b30_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire30_0_3));
INVC inst_inv_b30_0_3 (.A(imd_wire30_0_3),.Y(wire30_0_3));
NANDC2x1 inst_and_b30_1_0 (.A(wire30_0_0),.B(wire30_0_1),.Y(imd_wire30_1_0));
INVC inst_inv_b30_1_0 (.A(imd_wire30_1_0),.Y(wire30_1_0));
NANDC2x1 inst_and_b30_1_1 (.A(wire30_0_2),.B(wire30_0_3),.Y(imd_wire30_1_1));
INVC inst_inv_b30_1_1 (.A(imd_wire30_1_1),.Y(wire30_1_1));
NANDC2x1 inst_and_b30_2_0 (.A(wire30_1_0),.B(wire30_1_1),.Y(imd_Y30));
INVC inst_inv_b30_2_0 (.A(imd_Y30),.Y(Y30));
NANDC2x1 inst_clockedAND_b30_30 (.A(CLK),.B(Y30),.Y(imd_YF30));
INVC inst_clockedinv_b30_30 (.A(imd_YF30),.Y(YF30));


NANDC2x1 inst_and_b31_0_0 (.A(A0),.B(A1),.Y(imd_wire31_0_0));
INVC inst_inv_b31_0_0 (.A(imd_wire31_0_0),.Y(wire31_0_0));
NANDC2x1 inst_and_b31_0_1 (.A(A2),.B(A3),.Y(imd_wire31_0_1));
INVC inst_inv_b31_0_1 (.A(imd_wire31_0_1),.Y(wire31_0_1));
NANDC2x1 inst_and_b31_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire31_0_2));
INVC inst_inv_b31_0_2 (.A(imd_wire31_0_2),.Y(wire31_0_2));
NANDC2x1 inst_and_b31_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire31_0_3));
INVC inst_inv_b31_0_3 (.A(imd_wire31_0_3),.Y(wire31_0_3));
NANDC2x1 inst_and_b31_1_0 (.A(wire31_0_0),.B(wire31_0_1),.Y(imd_wire31_1_0));
INVC inst_inv_b31_1_0 (.A(imd_wire31_1_0),.Y(wire31_1_0));
NANDC2x1 inst_and_b31_1_1 (.A(wire31_0_2),.B(wire31_0_3),.Y(imd_wire31_1_1));
INVC inst_inv_b31_1_1 (.A(imd_wire31_1_1),.Y(wire31_1_1));
NANDC2x1 inst_and_b31_2_0 (.A(wire31_1_0),.B(wire31_1_1),.Y(imd_Y31));
INVC inst_inv_b31_2_0 (.A(imd_Y31),.Y(Y31));
NANDC2x1 inst_clockedAND_b31_31 (.A(CLK),.B(Y31),.Y(imd_YF31));
INVC inst_clockedinv_b31_31 (.A(imd_YF31),.Y(YF31));


NANDC2x1 inst_and_b32_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire32_0_0));
INVC inst_inv_b32_0_0 (.A(imd_wire32_0_0),.Y(wire32_0_0));
NANDC2x1 inst_and_b32_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire32_0_1));
INVC inst_inv_b32_0_1 (.A(imd_wire32_0_1),.Y(wire32_0_1));
NANDC2x1 inst_and_b32_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire32_0_2));
INVC inst_inv_b32_0_2 (.A(imd_wire32_0_2),.Y(wire32_0_2));
NANDC2x1 inst_and_b32_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire32_0_3));
INVC inst_inv_b32_0_3 (.A(imd_wire32_0_3),.Y(wire32_0_3));
NANDC2x1 inst_and_b32_1_0 (.A(wire32_0_0),.B(wire32_0_1),.Y(imd_wire32_1_0));
INVC inst_inv_b32_1_0 (.A(imd_wire32_1_0),.Y(wire32_1_0));
NANDC2x1 inst_and_b32_1_1 (.A(wire32_0_2),.B(wire32_0_3),.Y(imd_wire32_1_1));
INVC inst_inv_b32_1_1 (.A(imd_wire32_1_1),.Y(wire32_1_1));
NANDC2x1 inst_and_b32_2_0 (.A(wire32_1_0),.B(wire32_1_1),.Y(imd_Y32));
INVC inst_inv_b32_2_0 (.A(imd_Y32),.Y(Y32));
NANDC2x1 inst_clockedAND_b32_32 (.A(CLK),.B(Y32),.Y(imd_YF32));
INVC inst_clockedinv_b32_32 (.A(imd_YF32),.Y(YF32));


NANDC2x1 inst_and_b33_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire33_0_0));
INVC inst_inv_b33_0_0 (.A(imd_wire33_0_0),.Y(wire33_0_0));
NANDC2x1 inst_and_b33_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire33_0_1));
INVC inst_inv_b33_0_1 (.A(imd_wire33_0_1),.Y(wire33_0_1));
NANDC2x1 inst_and_b33_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire33_0_2));
INVC inst_inv_b33_0_2 (.A(imd_wire33_0_2),.Y(wire33_0_2));
NANDC2x1 inst_and_b33_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire33_0_3));
INVC inst_inv_b33_0_3 (.A(imd_wire33_0_3),.Y(wire33_0_3));
NANDC2x1 inst_and_b33_1_0 (.A(wire33_0_0),.B(wire33_0_1),.Y(imd_wire33_1_0));
INVC inst_inv_b33_1_0 (.A(imd_wire33_1_0),.Y(wire33_1_0));
NANDC2x1 inst_and_b33_1_1 (.A(wire33_0_2),.B(wire33_0_3),.Y(imd_wire33_1_1));
INVC inst_inv_b33_1_1 (.A(imd_wire33_1_1),.Y(wire33_1_1));
NANDC2x1 inst_and_b33_2_0 (.A(wire33_1_0),.B(wire33_1_1),.Y(imd_Y33));
INVC inst_inv_b33_2_0 (.A(imd_Y33),.Y(Y33));
NANDC2x1 inst_clockedAND_b33_33 (.A(CLK),.B(Y33),.Y(imd_YF33));
INVC inst_clockedinv_b33_33 (.A(imd_YF33),.Y(YF33));


NANDC2x1 inst_and_b34_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire34_0_0));
INVC inst_inv_b34_0_0 (.A(imd_wire34_0_0),.Y(wire34_0_0));
NANDC2x1 inst_and_b34_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire34_0_1));
INVC inst_inv_b34_0_1 (.A(imd_wire34_0_1),.Y(wire34_0_1));
NANDC2x1 inst_and_b34_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire34_0_2));
INVC inst_inv_b34_0_2 (.A(imd_wire34_0_2),.Y(wire34_0_2));
NANDC2x1 inst_and_b34_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire34_0_3));
INVC inst_inv_b34_0_3 (.A(imd_wire34_0_3),.Y(wire34_0_3));
NANDC2x1 inst_and_b34_1_0 (.A(wire34_0_0),.B(wire34_0_1),.Y(imd_wire34_1_0));
INVC inst_inv_b34_1_0 (.A(imd_wire34_1_0),.Y(wire34_1_0));
NANDC2x1 inst_and_b34_1_1 (.A(wire34_0_2),.B(wire34_0_3),.Y(imd_wire34_1_1));
INVC inst_inv_b34_1_1 (.A(imd_wire34_1_1),.Y(wire34_1_1));
NANDC2x1 inst_and_b34_2_0 (.A(wire34_1_0),.B(wire34_1_1),.Y(imd_Y34));
INVC inst_inv_b34_2_0 (.A(imd_Y34),.Y(Y34));
NANDC2x1 inst_clockedAND_b34_34 (.A(CLK),.B(Y34),.Y(imd_YF34));
INVC inst_clockedinv_b34_34 (.A(imd_YF34),.Y(YF34));


NANDC2x1 inst_and_b35_0_0 (.A(A0),.B(A1),.Y(imd_wire35_0_0));
INVC inst_inv_b35_0_0 (.A(imd_wire35_0_0),.Y(wire35_0_0));
NANDC2x1 inst_and_b35_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire35_0_1));
INVC inst_inv_b35_0_1 (.A(imd_wire35_0_1),.Y(wire35_0_1));
NANDC2x1 inst_and_b35_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire35_0_2));
INVC inst_inv_b35_0_2 (.A(imd_wire35_0_2),.Y(wire35_0_2));
NANDC2x1 inst_and_b35_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire35_0_3));
INVC inst_inv_b35_0_3 (.A(imd_wire35_0_3),.Y(wire35_0_3));
NANDC2x1 inst_and_b35_1_0 (.A(wire35_0_0),.B(wire35_0_1),.Y(imd_wire35_1_0));
INVC inst_inv_b35_1_0 (.A(imd_wire35_1_0),.Y(wire35_1_0));
NANDC2x1 inst_and_b35_1_1 (.A(wire35_0_2),.B(wire35_0_3),.Y(imd_wire35_1_1));
INVC inst_inv_b35_1_1 (.A(imd_wire35_1_1),.Y(wire35_1_1));
NANDC2x1 inst_and_b35_2_0 (.A(wire35_1_0),.B(wire35_1_1),.Y(imd_Y35));
INVC inst_inv_b35_2_0 (.A(imd_Y35),.Y(Y35));
NANDC2x1 inst_clockedAND_b35_35 (.A(CLK),.B(Y35),.Y(imd_YF35));
INVC inst_clockedinv_b35_35 (.A(imd_YF35),.Y(YF35));


NANDC2x1 inst_and_b36_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire36_0_0));
INVC inst_inv_b36_0_0 (.A(imd_wire36_0_0),.Y(wire36_0_0));
NANDC2x1 inst_and_b36_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire36_0_1));
INVC inst_inv_b36_0_1 (.A(imd_wire36_0_1),.Y(wire36_0_1));
NANDC2x1 inst_and_b36_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire36_0_2));
INVC inst_inv_b36_0_2 (.A(imd_wire36_0_2),.Y(wire36_0_2));
NANDC2x1 inst_and_b36_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire36_0_3));
INVC inst_inv_b36_0_3 (.A(imd_wire36_0_3),.Y(wire36_0_3));
NANDC2x1 inst_and_b36_1_0 (.A(wire36_0_0),.B(wire36_0_1),.Y(imd_wire36_1_0));
INVC inst_inv_b36_1_0 (.A(imd_wire36_1_0),.Y(wire36_1_0));
NANDC2x1 inst_and_b36_1_1 (.A(wire36_0_2),.B(wire36_0_3),.Y(imd_wire36_1_1));
INVC inst_inv_b36_1_1 (.A(imd_wire36_1_1),.Y(wire36_1_1));
NANDC2x1 inst_and_b36_2_0 (.A(wire36_1_0),.B(wire36_1_1),.Y(imd_Y36));
INVC inst_inv_b36_2_0 (.A(imd_Y36),.Y(Y36));
NANDC2x1 inst_clockedAND_b36_36 (.A(CLK),.B(Y36),.Y(imd_YF36));
INVC inst_clockedinv_b36_36 (.A(imd_YF36),.Y(YF36));


NANDC2x1 inst_and_b37_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire37_0_0));
INVC inst_inv_b37_0_0 (.A(imd_wire37_0_0),.Y(wire37_0_0));
NANDC2x1 inst_and_b37_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire37_0_1));
INVC inst_inv_b37_0_1 (.A(imd_wire37_0_1),.Y(wire37_0_1));
NANDC2x1 inst_and_b37_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire37_0_2));
INVC inst_inv_b37_0_2 (.A(imd_wire37_0_2),.Y(wire37_0_2));
NANDC2x1 inst_and_b37_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire37_0_3));
INVC inst_inv_b37_0_3 (.A(imd_wire37_0_3),.Y(wire37_0_3));
NANDC2x1 inst_and_b37_1_0 (.A(wire37_0_0),.B(wire37_0_1),.Y(imd_wire37_1_0));
INVC inst_inv_b37_1_0 (.A(imd_wire37_1_0),.Y(wire37_1_0));
NANDC2x1 inst_and_b37_1_1 (.A(wire37_0_2),.B(wire37_0_3),.Y(imd_wire37_1_1));
INVC inst_inv_b37_1_1 (.A(imd_wire37_1_1),.Y(wire37_1_1));
NANDC2x1 inst_and_b37_2_0 (.A(wire37_1_0),.B(wire37_1_1),.Y(imd_Y37));
INVC inst_inv_b37_2_0 (.A(imd_Y37),.Y(Y37));
NANDC2x1 inst_clockedAND_b37_37 (.A(CLK),.B(Y37),.Y(imd_YF37));
INVC inst_clockedinv_b37_37 (.A(imd_YF37),.Y(YF37));


NANDC2x1 inst_and_b38_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire38_0_0));
INVC inst_inv_b38_0_0 (.A(imd_wire38_0_0),.Y(wire38_0_0));
NANDC2x1 inst_and_b38_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire38_0_1));
INVC inst_inv_b38_0_1 (.A(imd_wire38_0_1),.Y(wire38_0_1));
NANDC2x1 inst_and_b38_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire38_0_2));
INVC inst_inv_b38_0_2 (.A(imd_wire38_0_2),.Y(wire38_0_2));
NANDC2x1 inst_and_b38_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire38_0_3));
INVC inst_inv_b38_0_3 (.A(imd_wire38_0_3),.Y(wire38_0_3));
NANDC2x1 inst_and_b38_1_0 (.A(wire38_0_0),.B(wire38_0_1),.Y(imd_wire38_1_0));
INVC inst_inv_b38_1_0 (.A(imd_wire38_1_0),.Y(wire38_1_0));
NANDC2x1 inst_and_b38_1_1 (.A(wire38_0_2),.B(wire38_0_3),.Y(imd_wire38_1_1));
INVC inst_inv_b38_1_1 (.A(imd_wire38_1_1),.Y(wire38_1_1));
NANDC2x1 inst_and_b38_2_0 (.A(wire38_1_0),.B(wire38_1_1),.Y(imd_Y38));
INVC inst_inv_b38_2_0 (.A(imd_Y38),.Y(Y38));
NANDC2x1 inst_clockedAND_b38_38 (.A(CLK),.B(Y38),.Y(imd_YF38));
INVC inst_clockedinv_b38_38 (.A(imd_YF38),.Y(YF38));


NANDC2x1 inst_and_b39_0_0 (.A(A0),.B(A1),.Y(imd_wire39_0_0));
INVC inst_inv_b39_0_0 (.A(imd_wire39_0_0),.Y(wire39_0_0));
NANDC2x1 inst_and_b39_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire39_0_1));
INVC inst_inv_b39_0_1 (.A(imd_wire39_0_1),.Y(wire39_0_1));
NANDC2x1 inst_and_b39_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire39_0_2));
INVC inst_inv_b39_0_2 (.A(imd_wire39_0_2),.Y(wire39_0_2));
NANDC2x1 inst_and_b39_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire39_0_3));
INVC inst_inv_b39_0_3 (.A(imd_wire39_0_3),.Y(wire39_0_3));
NANDC2x1 inst_and_b39_1_0 (.A(wire39_0_0),.B(wire39_0_1),.Y(imd_wire39_1_0));
INVC inst_inv_b39_1_0 (.A(imd_wire39_1_0),.Y(wire39_1_0));
NANDC2x1 inst_and_b39_1_1 (.A(wire39_0_2),.B(wire39_0_3),.Y(imd_wire39_1_1));
INVC inst_inv_b39_1_1 (.A(imd_wire39_1_1),.Y(wire39_1_1));
NANDC2x1 inst_and_b39_2_0 (.A(wire39_1_0),.B(wire39_1_1),.Y(imd_Y39));
INVC inst_inv_b39_2_0 (.A(imd_Y39),.Y(Y39));
NANDC2x1 inst_clockedAND_b39_39 (.A(CLK),.B(Y39),.Y(imd_YF39));
INVC inst_clockedinv_b39_39 (.A(imd_YF39),.Y(YF39));


NANDC2x1 inst_and_b40_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire40_0_0));
INVC inst_inv_b40_0_0 (.A(imd_wire40_0_0),.Y(wire40_0_0));
NANDC2x1 inst_and_b40_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire40_0_1));
INVC inst_inv_b40_0_1 (.A(imd_wire40_0_1),.Y(wire40_0_1));
NANDC2x1 inst_and_b40_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire40_0_2));
INVC inst_inv_b40_0_2 (.A(imd_wire40_0_2),.Y(wire40_0_2));
NANDC2x1 inst_and_b40_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire40_0_3));
INVC inst_inv_b40_0_3 (.A(imd_wire40_0_3),.Y(wire40_0_3));
NANDC2x1 inst_and_b40_1_0 (.A(wire40_0_0),.B(wire40_0_1),.Y(imd_wire40_1_0));
INVC inst_inv_b40_1_0 (.A(imd_wire40_1_0),.Y(wire40_1_0));
NANDC2x1 inst_and_b40_1_1 (.A(wire40_0_2),.B(wire40_0_3),.Y(imd_wire40_1_1));
INVC inst_inv_b40_1_1 (.A(imd_wire40_1_1),.Y(wire40_1_1));
NANDC2x1 inst_and_b40_2_0 (.A(wire40_1_0),.B(wire40_1_1),.Y(imd_Y40));
INVC inst_inv_b40_2_0 (.A(imd_Y40),.Y(Y40));
NANDC2x1 inst_clockedAND_b40_40 (.A(CLK),.B(Y40),.Y(imd_YF40));
INVC inst_clockedinv_b40_40 (.A(imd_YF40),.Y(YF40));


NANDC2x1 inst_and_b41_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire41_0_0));
INVC inst_inv_b41_0_0 (.A(imd_wire41_0_0),.Y(wire41_0_0));
NANDC2x1 inst_and_b41_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire41_0_1));
INVC inst_inv_b41_0_1 (.A(imd_wire41_0_1),.Y(wire41_0_1));
NANDC2x1 inst_and_b41_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire41_0_2));
INVC inst_inv_b41_0_2 (.A(imd_wire41_0_2),.Y(wire41_0_2));
NANDC2x1 inst_and_b41_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire41_0_3));
INVC inst_inv_b41_0_3 (.A(imd_wire41_0_3),.Y(wire41_0_3));
NANDC2x1 inst_and_b41_1_0 (.A(wire41_0_0),.B(wire41_0_1),.Y(imd_wire41_1_0));
INVC inst_inv_b41_1_0 (.A(imd_wire41_1_0),.Y(wire41_1_0));
NANDC2x1 inst_and_b41_1_1 (.A(wire41_0_2),.B(wire41_0_3),.Y(imd_wire41_1_1));
INVC inst_inv_b41_1_1 (.A(imd_wire41_1_1),.Y(wire41_1_1));
NANDC2x1 inst_and_b41_2_0 (.A(wire41_1_0),.B(wire41_1_1),.Y(imd_Y41));
INVC inst_inv_b41_2_0 (.A(imd_Y41),.Y(Y41));
NANDC2x1 inst_clockedAND_b41_41 (.A(CLK),.B(Y41),.Y(imd_YF41));
INVC inst_clockedinv_b41_41 (.A(imd_YF41),.Y(YF41));


NANDC2x1 inst_and_b42_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire42_0_0));
INVC inst_inv_b42_0_0 (.A(imd_wire42_0_0),.Y(wire42_0_0));
NANDC2x1 inst_and_b42_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire42_0_1));
INVC inst_inv_b42_0_1 (.A(imd_wire42_0_1),.Y(wire42_0_1));
NANDC2x1 inst_and_b42_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire42_0_2));
INVC inst_inv_b42_0_2 (.A(imd_wire42_0_2),.Y(wire42_0_2));
NANDC2x1 inst_and_b42_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire42_0_3));
INVC inst_inv_b42_0_3 (.A(imd_wire42_0_3),.Y(wire42_0_3));
NANDC2x1 inst_and_b42_1_0 (.A(wire42_0_0),.B(wire42_0_1),.Y(imd_wire42_1_0));
INVC inst_inv_b42_1_0 (.A(imd_wire42_1_0),.Y(wire42_1_0));
NANDC2x1 inst_and_b42_1_1 (.A(wire42_0_2),.B(wire42_0_3),.Y(imd_wire42_1_1));
INVC inst_inv_b42_1_1 (.A(imd_wire42_1_1),.Y(wire42_1_1));
NANDC2x1 inst_and_b42_2_0 (.A(wire42_1_0),.B(wire42_1_1),.Y(imd_Y42));
INVC inst_inv_b42_2_0 (.A(imd_Y42),.Y(Y42));
NANDC2x1 inst_clockedAND_b42_42 (.A(CLK),.B(Y42),.Y(imd_YF42));
INVC inst_clockedinv_b42_42 (.A(imd_YF42),.Y(YF42));


NANDC2x1 inst_and_b43_0_0 (.A(A0),.B(A1),.Y(imd_wire43_0_0));
INVC inst_inv_b43_0_0 (.A(imd_wire43_0_0),.Y(wire43_0_0));
NANDC2x1 inst_and_b43_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire43_0_1));
INVC inst_inv_b43_0_1 (.A(imd_wire43_0_1),.Y(wire43_0_1));
NANDC2x1 inst_and_b43_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire43_0_2));
INVC inst_inv_b43_0_2 (.A(imd_wire43_0_2),.Y(wire43_0_2));
NANDC2x1 inst_and_b43_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire43_0_3));
INVC inst_inv_b43_0_3 (.A(imd_wire43_0_3),.Y(wire43_0_3));
NANDC2x1 inst_and_b43_1_0 (.A(wire43_0_0),.B(wire43_0_1),.Y(imd_wire43_1_0));
INVC inst_inv_b43_1_0 (.A(imd_wire43_1_0),.Y(wire43_1_0));
NANDC2x1 inst_and_b43_1_1 (.A(wire43_0_2),.B(wire43_0_3),.Y(imd_wire43_1_1));
INVC inst_inv_b43_1_1 (.A(imd_wire43_1_1),.Y(wire43_1_1));
NANDC2x1 inst_and_b43_2_0 (.A(wire43_1_0),.B(wire43_1_1),.Y(imd_Y43));
INVC inst_inv_b43_2_0 (.A(imd_Y43),.Y(Y43));
NANDC2x1 inst_clockedAND_b43_43 (.A(CLK),.B(Y43),.Y(imd_YF43));
INVC inst_clockedinv_b43_43 (.A(imd_YF43),.Y(YF43));


NANDC2x1 inst_and_b44_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire44_0_0));
INVC inst_inv_b44_0_0 (.A(imd_wire44_0_0),.Y(wire44_0_0));
NANDC2x1 inst_and_b44_0_1 (.A(A2),.B(A3),.Y(imd_wire44_0_1));
INVC inst_inv_b44_0_1 (.A(imd_wire44_0_1),.Y(wire44_0_1));
NANDC2x1 inst_and_b44_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire44_0_2));
INVC inst_inv_b44_0_2 (.A(imd_wire44_0_2),.Y(wire44_0_2));
NANDC2x1 inst_and_b44_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire44_0_3));
INVC inst_inv_b44_0_3 (.A(imd_wire44_0_3),.Y(wire44_0_3));
NANDC2x1 inst_and_b44_1_0 (.A(wire44_0_0),.B(wire44_0_1),.Y(imd_wire44_1_0));
INVC inst_inv_b44_1_0 (.A(imd_wire44_1_0),.Y(wire44_1_0));
NANDC2x1 inst_and_b44_1_1 (.A(wire44_0_2),.B(wire44_0_3),.Y(imd_wire44_1_1));
INVC inst_inv_b44_1_1 (.A(imd_wire44_1_1),.Y(wire44_1_1));
NANDC2x1 inst_and_b44_2_0 (.A(wire44_1_0),.B(wire44_1_1),.Y(imd_Y44));
INVC inst_inv_b44_2_0 (.A(imd_Y44),.Y(Y44));
NANDC2x1 inst_clockedAND_b44_44 (.A(CLK),.B(Y44),.Y(imd_YF44));
INVC inst_clockedinv_b44_44 (.A(imd_YF44),.Y(YF44));


NANDC2x1 inst_and_b45_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire45_0_0));
INVC inst_inv_b45_0_0 (.A(imd_wire45_0_0),.Y(wire45_0_0));
NANDC2x1 inst_and_b45_0_1 (.A(A2),.B(A3),.Y(imd_wire45_0_1));
INVC inst_inv_b45_0_1 (.A(imd_wire45_0_1),.Y(wire45_0_1));
NANDC2x1 inst_and_b45_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire45_0_2));
INVC inst_inv_b45_0_2 (.A(imd_wire45_0_2),.Y(wire45_0_2));
NANDC2x1 inst_and_b45_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire45_0_3));
INVC inst_inv_b45_0_3 (.A(imd_wire45_0_3),.Y(wire45_0_3));
NANDC2x1 inst_and_b45_1_0 (.A(wire45_0_0),.B(wire45_0_1),.Y(imd_wire45_1_0));
INVC inst_inv_b45_1_0 (.A(imd_wire45_1_0),.Y(wire45_1_0));
NANDC2x1 inst_and_b45_1_1 (.A(wire45_0_2),.B(wire45_0_3),.Y(imd_wire45_1_1));
INVC inst_inv_b45_1_1 (.A(imd_wire45_1_1),.Y(wire45_1_1));
NANDC2x1 inst_and_b45_2_0 (.A(wire45_1_0),.B(wire45_1_1),.Y(imd_Y45));
INVC inst_inv_b45_2_0 (.A(imd_Y45),.Y(Y45));
NANDC2x1 inst_clockedAND_b45_45 (.A(CLK),.B(Y45),.Y(imd_YF45));
INVC inst_clockedinv_b45_45 (.A(imd_YF45),.Y(YF45));


NANDC2x1 inst_and_b46_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire46_0_0));
INVC inst_inv_b46_0_0 (.A(imd_wire46_0_0),.Y(wire46_0_0));
NANDC2x1 inst_and_b46_0_1 (.A(A2),.B(A3),.Y(imd_wire46_0_1));
INVC inst_inv_b46_0_1 (.A(imd_wire46_0_1),.Y(wire46_0_1));
NANDC2x1 inst_and_b46_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire46_0_2));
INVC inst_inv_b46_0_2 (.A(imd_wire46_0_2),.Y(wire46_0_2));
NANDC2x1 inst_and_b46_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire46_0_3));
INVC inst_inv_b46_0_3 (.A(imd_wire46_0_3),.Y(wire46_0_3));
NANDC2x1 inst_and_b46_1_0 (.A(wire46_0_0),.B(wire46_0_1),.Y(imd_wire46_1_0));
INVC inst_inv_b46_1_0 (.A(imd_wire46_1_0),.Y(wire46_1_0));
NANDC2x1 inst_and_b46_1_1 (.A(wire46_0_2),.B(wire46_0_3),.Y(imd_wire46_1_1));
INVC inst_inv_b46_1_1 (.A(imd_wire46_1_1),.Y(wire46_1_1));
NANDC2x1 inst_and_b46_2_0 (.A(wire46_1_0),.B(wire46_1_1),.Y(imd_Y46));
INVC inst_inv_b46_2_0 (.A(imd_Y46),.Y(Y46));
NANDC2x1 inst_clockedAND_b46_46 (.A(CLK),.B(Y46),.Y(imd_YF46));
INVC inst_clockedinv_b46_46 (.A(imd_YF46),.Y(YF46));


NANDC2x1 inst_and_b47_0_0 (.A(A0),.B(A1),.Y(imd_wire47_0_0));
INVC inst_inv_b47_0_0 (.A(imd_wire47_0_0),.Y(wire47_0_0));
NANDC2x1 inst_and_b47_0_1 (.A(A2),.B(A3),.Y(imd_wire47_0_1));
INVC inst_inv_b47_0_1 (.A(imd_wire47_0_1),.Y(wire47_0_1));
NANDC2x1 inst_and_b47_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire47_0_2));
INVC inst_inv_b47_0_2 (.A(imd_wire47_0_2),.Y(wire47_0_2));
NANDC2x1 inst_and_b47_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire47_0_3));
INVC inst_inv_b47_0_3 (.A(imd_wire47_0_3),.Y(wire47_0_3));
NANDC2x1 inst_and_b47_1_0 (.A(wire47_0_0),.B(wire47_0_1),.Y(imd_wire47_1_0));
INVC inst_inv_b47_1_0 (.A(imd_wire47_1_0),.Y(wire47_1_0));
NANDC2x1 inst_and_b47_1_1 (.A(wire47_0_2),.B(wire47_0_3),.Y(imd_wire47_1_1));
INVC inst_inv_b47_1_1 (.A(imd_wire47_1_1),.Y(wire47_1_1));
NANDC2x1 inst_and_b47_2_0 (.A(wire47_1_0),.B(wire47_1_1),.Y(imd_Y47));
INVC inst_inv_b47_2_0 (.A(imd_Y47),.Y(Y47));
NANDC2x1 inst_clockedAND_b47_47 (.A(CLK),.B(Y47),.Y(imd_YF47));
INVC inst_clockedinv_b47_47 (.A(imd_YF47),.Y(YF47));


NANDC2x1 inst_and_b48_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire48_0_0));
INVC inst_inv_b48_0_0 (.A(imd_wire48_0_0),.Y(wire48_0_0));
NANDC2x1 inst_and_b48_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire48_0_1));
INVC inst_inv_b48_0_1 (.A(imd_wire48_0_1),.Y(wire48_0_1));
NANDC2x1 inst_and_b48_0_2 (.A(A4),.B(A5),.Y(imd_wire48_0_2));
INVC inst_inv_b48_0_2 (.A(imd_wire48_0_2),.Y(wire48_0_2));
NANDC2x1 inst_and_b48_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire48_0_3));
INVC inst_inv_b48_0_3 (.A(imd_wire48_0_3),.Y(wire48_0_3));
NANDC2x1 inst_and_b48_1_0 (.A(wire48_0_0),.B(wire48_0_1),.Y(imd_wire48_1_0));
INVC inst_inv_b48_1_0 (.A(imd_wire48_1_0),.Y(wire48_1_0));
NANDC2x1 inst_and_b48_1_1 (.A(wire48_0_2),.B(wire48_0_3),.Y(imd_wire48_1_1));
INVC inst_inv_b48_1_1 (.A(imd_wire48_1_1),.Y(wire48_1_1));
NANDC2x1 inst_and_b48_2_0 (.A(wire48_1_0),.B(wire48_1_1),.Y(imd_Y48));
INVC inst_inv_b48_2_0 (.A(imd_Y48),.Y(Y48));
NANDC2x1 inst_clockedAND_b48_48 (.A(CLK),.B(Y48),.Y(imd_YF48));
INVC inst_clockedinv_b48_48 (.A(imd_YF48),.Y(YF48));


NANDC2x1 inst_and_b49_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire49_0_0));
INVC inst_inv_b49_0_0 (.A(imd_wire49_0_0),.Y(wire49_0_0));
NANDC2x1 inst_and_b49_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire49_0_1));
INVC inst_inv_b49_0_1 (.A(imd_wire49_0_1),.Y(wire49_0_1));
NANDC2x1 inst_and_b49_0_2 (.A(A4),.B(A5),.Y(imd_wire49_0_2));
INVC inst_inv_b49_0_2 (.A(imd_wire49_0_2),.Y(wire49_0_2));
NANDC2x1 inst_and_b49_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire49_0_3));
INVC inst_inv_b49_0_3 (.A(imd_wire49_0_3),.Y(wire49_0_3));
NANDC2x1 inst_and_b49_1_0 (.A(wire49_0_0),.B(wire49_0_1),.Y(imd_wire49_1_0));
INVC inst_inv_b49_1_0 (.A(imd_wire49_1_0),.Y(wire49_1_0));
NANDC2x1 inst_and_b49_1_1 (.A(wire49_0_2),.B(wire49_0_3),.Y(imd_wire49_1_1));
INVC inst_inv_b49_1_1 (.A(imd_wire49_1_1),.Y(wire49_1_1));
NANDC2x1 inst_and_b49_2_0 (.A(wire49_1_0),.B(wire49_1_1),.Y(imd_Y49));
INVC inst_inv_b49_2_0 (.A(imd_Y49),.Y(Y49));
NANDC2x1 inst_clockedAND_b49_49 (.A(CLK),.B(Y49),.Y(imd_YF49));
INVC inst_clockedinv_b49_49 (.A(imd_YF49),.Y(YF49));


NANDC2x1 inst_and_b50_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire50_0_0));
INVC inst_inv_b50_0_0 (.A(imd_wire50_0_0),.Y(wire50_0_0));
NANDC2x1 inst_and_b50_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire50_0_1));
INVC inst_inv_b50_0_1 (.A(imd_wire50_0_1),.Y(wire50_0_1));
NANDC2x1 inst_and_b50_0_2 (.A(A4),.B(A5),.Y(imd_wire50_0_2));
INVC inst_inv_b50_0_2 (.A(imd_wire50_0_2),.Y(wire50_0_2));
NANDC2x1 inst_and_b50_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire50_0_3));
INVC inst_inv_b50_0_3 (.A(imd_wire50_0_3),.Y(wire50_0_3));
NANDC2x1 inst_and_b50_1_0 (.A(wire50_0_0),.B(wire50_0_1),.Y(imd_wire50_1_0));
INVC inst_inv_b50_1_0 (.A(imd_wire50_1_0),.Y(wire50_1_0));
NANDC2x1 inst_and_b50_1_1 (.A(wire50_0_2),.B(wire50_0_3),.Y(imd_wire50_1_1));
INVC inst_inv_b50_1_1 (.A(imd_wire50_1_1),.Y(wire50_1_1));
NANDC2x1 inst_and_b50_2_0 (.A(wire50_1_0),.B(wire50_1_1),.Y(imd_Y50));
INVC inst_inv_b50_2_0 (.A(imd_Y50),.Y(Y50));
NANDC2x1 inst_clockedAND_b50_50 (.A(CLK),.B(Y50),.Y(imd_YF50));
INVC inst_clockedinv_b50_50 (.A(imd_YF50),.Y(YF50));


NANDC2x1 inst_and_b51_0_0 (.A(A0),.B(A1),.Y(imd_wire51_0_0));
INVC inst_inv_b51_0_0 (.A(imd_wire51_0_0),.Y(wire51_0_0));
NANDC2x1 inst_and_b51_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire51_0_1));
INVC inst_inv_b51_0_1 (.A(imd_wire51_0_1),.Y(wire51_0_1));
NANDC2x1 inst_and_b51_0_2 (.A(A4),.B(A5),.Y(imd_wire51_0_2));
INVC inst_inv_b51_0_2 (.A(imd_wire51_0_2),.Y(wire51_0_2));
NANDC2x1 inst_and_b51_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire51_0_3));
INVC inst_inv_b51_0_3 (.A(imd_wire51_0_3),.Y(wire51_0_3));
NANDC2x1 inst_and_b51_1_0 (.A(wire51_0_0),.B(wire51_0_1),.Y(imd_wire51_1_0));
INVC inst_inv_b51_1_0 (.A(imd_wire51_1_0),.Y(wire51_1_0));
NANDC2x1 inst_and_b51_1_1 (.A(wire51_0_2),.B(wire51_0_3),.Y(imd_wire51_1_1));
INVC inst_inv_b51_1_1 (.A(imd_wire51_1_1),.Y(wire51_1_1));
NANDC2x1 inst_and_b51_2_0 (.A(wire51_1_0),.B(wire51_1_1),.Y(imd_Y51));
INVC inst_inv_b51_2_0 (.A(imd_Y51),.Y(Y51));
NANDC2x1 inst_clockedAND_b51_51 (.A(CLK),.B(Y51),.Y(imd_YF51));
INVC inst_clockedinv_b51_51 (.A(imd_YF51),.Y(YF51));


NANDC2x1 inst_and_b52_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire52_0_0));
INVC inst_inv_b52_0_0 (.A(imd_wire52_0_0),.Y(wire52_0_0));
NANDC2x1 inst_and_b52_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire52_0_1));
INVC inst_inv_b52_0_1 (.A(imd_wire52_0_1),.Y(wire52_0_1));
NANDC2x1 inst_and_b52_0_2 (.A(A4),.B(A5),.Y(imd_wire52_0_2));
INVC inst_inv_b52_0_2 (.A(imd_wire52_0_2),.Y(wire52_0_2));
NANDC2x1 inst_and_b52_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire52_0_3));
INVC inst_inv_b52_0_3 (.A(imd_wire52_0_3),.Y(wire52_0_3));
NANDC2x1 inst_and_b52_1_0 (.A(wire52_0_0),.B(wire52_0_1),.Y(imd_wire52_1_0));
INVC inst_inv_b52_1_0 (.A(imd_wire52_1_0),.Y(wire52_1_0));
NANDC2x1 inst_and_b52_1_1 (.A(wire52_0_2),.B(wire52_0_3),.Y(imd_wire52_1_1));
INVC inst_inv_b52_1_1 (.A(imd_wire52_1_1),.Y(wire52_1_1));
NANDC2x1 inst_and_b52_2_0 (.A(wire52_1_0),.B(wire52_1_1),.Y(imd_Y52));
INVC inst_inv_b52_2_0 (.A(imd_Y52),.Y(Y52));
NANDC2x1 inst_clockedAND_b52_52 (.A(CLK),.B(Y52),.Y(imd_YF52));
INVC inst_clockedinv_b52_52 (.A(imd_YF52),.Y(YF52));


NANDC2x1 inst_and_b53_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire53_0_0));
INVC inst_inv_b53_0_0 (.A(imd_wire53_0_0),.Y(wire53_0_0));
NANDC2x1 inst_and_b53_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire53_0_1));
INVC inst_inv_b53_0_1 (.A(imd_wire53_0_1),.Y(wire53_0_1));
NANDC2x1 inst_and_b53_0_2 (.A(A4),.B(A5),.Y(imd_wire53_0_2));
INVC inst_inv_b53_0_2 (.A(imd_wire53_0_2),.Y(wire53_0_2));
NANDC2x1 inst_and_b53_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire53_0_3));
INVC inst_inv_b53_0_3 (.A(imd_wire53_0_3),.Y(wire53_0_3));
NANDC2x1 inst_and_b53_1_0 (.A(wire53_0_0),.B(wire53_0_1),.Y(imd_wire53_1_0));
INVC inst_inv_b53_1_0 (.A(imd_wire53_1_0),.Y(wire53_1_0));
NANDC2x1 inst_and_b53_1_1 (.A(wire53_0_2),.B(wire53_0_3),.Y(imd_wire53_1_1));
INVC inst_inv_b53_1_1 (.A(imd_wire53_1_1),.Y(wire53_1_1));
NANDC2x1 inst_and_b53_2_0 (.A(wire53_1_0),.B(wire53_1_1),.Y(imd_Y53));
INVC inst_inv_b53_2_0 (.A(imd_Y53),.Y(Y53));
NANDC2x1 inst_clockedAND_b53_53 (.A(CLK),.B(Y53),.Y(imd_YF53));
INVC inst_clockedinv_b53_53 (.A(imd_YF53),.Y(YF53));


NANDC2x1 inst_and_b54_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire54_0_0));
INVC inst_inv_b54_0_0 (.A(imd_wire54_0_0),.Y(wire54_0_0));
NANDC2x1 inst_and_b54_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire54_0_1));
INVC inst_inv_b54_0_1 (.A(imd_wire54_0_1),.Y(wire54_0_1));
NANDC2x1 inst_and_b54_0_2 (.A(A4),.B(A5),.Y(imd_wire54_0_2));
INVC inst_inv_b54_0_2 (.A(imd_wire54_0_2),.Y(wire54_0_2));
NANDC2x1 inst_and_b54_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire54_0_3));
INVC inst_inv_b54_0_3 (.A(imd_wire54_0_3),.Y(wire54_0_3));
NANDC2x1 inst_and_b54_1_0 (.A(wire54_0_0),.B(wire54_0_1),.Y(imd_wire54_1_0));
INVC inst_inv_b54_1_0 (.A(imd_wire54_1_0),.Y(wire54_1_0));
NANDC2x1 inst_and_b54_1_1 (.A(wire54_0_2),.B(wire54_0_3),.Y(imd_wire54_1_1));
INVC inst_inv_b54_1_1 (.A(imd_wire54_1_1),.Y(wire54_1_1));
NANDC2x1 inst_and_b54_2_0 (.A(wire54_1_0),.B(wire54_1_1),.Y(imd_Y54));
INVC inst_inv_b54_2_0 (.A(imd_Y54),.Y(Y54));
NANDC2x1 inst_clockedAND_b54_54 (.A(CLK),.B(Y54),.Y(imd_YF54));
INVC inst_clockedinv_b54_54 (.A(imd_YF54),.Y(YF54));


NANDC2x1 inst_and_b55_0_0 (.A(A0),.B(A1),.Y(imd_wire55_0_0));
INVC inst_inv_b55_0_0 (.A(imd_wire55_0_0),.Y(wire55_0_0));
NANDC2x1 inst_and_b55_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire55_0_1));
INVC inst_inv_b55_0_1 (.A(imd_wire55_0_1),.Y(wire55_0_1));
NANDC2x1 inst_and_b55_0_2 (.A(A4),.B(A5),.Y(imd_wire55_0_2));
INVC inst_inv_b55_0_2 (.A(imd_wire55_0_2),.Y(wire55_0_2));
NANDC2x1 inst_and_b55_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire55_0_3));
INVC inst_inv_b55_0_3 (.A(imd_wire55_0_3),.Y(wire55_0_3));
NANDC2x1 inst_and_b55_1_0 (.A(wire55_0_0),.B(wire55_0_1),.Y(imd_wire55_1_0));
INVC inst_inv_b55_1_0 (.A(imd_wire55_1_0),.Y(wire55_1_0));
NANDC2x1 inst_and_b55_1_1 (.A(wire55_0_2),.B(wire55_0_3),.Y(imd_wire55_1_1));
INVC inst_inv_b55_1_1 (.A(imd_wire55_1_1),.Y(wire55_1_1));
NANDC2x1 inst_and_b55_2_0 (.A(wire55_1_0),.B(wire55_1_1),.Y(imd_Y55));
INVC inst_inv_b55_2_0 (.A(imd_Y55),.Y(Y55));
NANDC2x1 inst_clockedAND_b55_55 (.A(CLK),.B(Y55),.Y(imd_YF55));
INVC inst_clockedinv_b55_55 (.A(imd_YF55),.Y(YF55));


NANDC2x1 inst_and_b56_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire56_0_0));
INVC inst_inv_b56_0_0 (.A(imd_wire56_0_0),.Y(wire56_0_0));
NANDC2x1 inst_and_b56_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire56_0_1));
INVC inst_inv_b56_0_1 (.A(imd_wire56_0_1),.Y(wire56_0_1));
NANDC2x1 inst_and_b56_0_2 (.A(A4),.B(A5),.Y(imd_wire56_0_2));
INVC inst_inv_b56_0_2 (.A(imd_wire56_0_2),.Y(wire56_0_2));
NANDC2x1 inst_and_b56_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire56_0_3));
INVC inst_inv_b56_0_3 (.A(imd_wire56_0_3),.Y(wire56_0_3));
NANDC2x1 inst_and_b56_1_0 (.A(wire56_0_0),.B(wire56_0_1),.Y(imd_wire56_1_0));
INVC inst_inv_b56_1_0 (.A(imd_wire56_1_0),.Y(wire56_1_0));
NANDC2x1 inst_and_b56_1_1 (.A(wire56_0_2),.B(wire56_0_3),.Y(imd_wire56_1_1));
INVC inst_inv_b56_1_1 (.A(imd_wire56_1_1),.Y(wire56_1_1));
NANDC2x1 inst_and_b56_2_0 (.A(wire56_1_0),.B(wire56_1_1),.Y(imd_Y56));
INVC inst_inv_b56_2_0 (.A(imd_Y56),.Y(Y56));
NANDC2x1 inst_clockedAND_b56_56 (.A(CLK),.B(Y56),.Y(imd_YF56));
INVC inst_clockedinv_b56_56 (.A(imd_YF56),.Y(YF56));


NANDC2x1 inst_and_b57_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire57_0_0));
INVC inst_inv_b57_0_0 (.A(imd_wire57_0_0),.Y(wire57_0_0));
NANDC2x1 inst_and_b57_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire57_0_1));
INVC inst_inv_b57_0_1 (.A(imd_wire57_0_1),.Y(wire57_0_1));
NANDC2x1 inst_and_b57_0_2 (.A(A4),.B(A5),.Y(imd_wire57_0_2));
INVC inst_inv_b57_0_2 (.A(imd_wire57_0_2),.Y(wire57_0_2));
NANDC2x1 inst_and_b57_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire57_0_3));
INVC inst_inv_b57_0_3 (.A(imd_wire57_0_3),.Y(wire57_0_3));
NANDC2x1 inst_and_b57_1_0 (.A(wire57_0_0),.B(wire57_0_1),.Y(imd_wire57_1_0));
INVC inst_inv_b57_1_0 (.A(imd_wire57_1_0),.Y(wire57_1_0));
NANDC2x1 inst_and_b57_1_1 (.A(wire57_0_2),.B(wire57_0_3),.Y(imd_wire57_1_1));
INVC inst_inv_b57_1_1 (.A(imd_wire57_1_1),.Y(wire57_1_1));
NANDC2x1 inst_and_b57_2_0 (.A(wire57_1_0),.B(wire57_1_1),.Y(imd_Y57));
INVC inst_inv_b57_2_0 (.A(imd_Y57),.Y(Y57));
NANDC2x1 inst_clockedAND_b57_57 (.A(CLK),.B(Y57),.Y(imd_YF57));
INVC inst_clockedinv_b57_57 (.A(imd_YF57),.Y(YF57));


NANDC2x1 inst_and_b58_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire58_0_0));
INVC inst_inv_b58_0_0 (.A(imd_wire58_0_0),.Y(wire58_0_0));
NANDC2x1 inst_and_b58_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire58_0_1));
INVC inst_inv_b58_0_1 (.A(imd_wire58_0_1),.Y(wire58_0_1));
NANDC2x1 inst_and_b58_0_2 (.A(A4),.B(A5),.Y(imd_wire58_0_2));
INVC inst_inv_b58_0_2 (.A(imd_wire58_0_2),.Y(wire58_0_2));
NANDC2x1 inst_and_b58_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire58_0_3));
INVC inst_inv_b58_0_3 (.A(imd_wire58_0_3),.Y(wire58_0_3));
NANDC2x1 inst_and_b58_1_0 (.A(wire58_0_0),.B(wire58_0_1),.Y(imd_wire58_1_0));
INVC inst_inv_b58_1_0 (.A(imd_wire58_1_0),.Y(wire58_1_0));
NANDC2x1 inst_and_b58_1_1 (.A(wire58_0_2),.B(wire58_0_3),.Y(imd_wire58_1_1));
INVC inst_inv_b58_1_1 (.A(imd_wire58_1_1),.Y(wire58_1_1));
NANDC2x1 inst_and_b58_2_0 (.A(wire58_1_0),.B(wire58_1_1),.Y(imd_Y58));
INVC inst_inv_b58_2_0 (.A(imd_Y58),.Y(Y58));
NANDC2x1 inst_clockedAND_b58_58 (.A(CLK),.B(Y58),.Y(imd_YF58));
INVC inst_clockedinv_b58_58 (.A(imd_YF58),.Y(YF58));


NANDC2x1 inst_and_b59_0_0 (.A(A0),.B(A1),.Y(imd_wire59_0_0));
INVC inst_inv_b59_0_0 (.A(imd_wire59_0_0),.Y(wire59_0_0));
NANDC2x1 inst_and_b59_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire59_0_1));
INVC inst_inv_b59_0_1 (.A(imd_wire59_0_1),.Y(wire59_0_1));
NANDC2x1 inst_and_b59_0_2 (.A(A4),.B(A5),.Y(imd_wire59_0_2));
INVC inst_inv_b59_0_2 (.A(imd_wire59_0_2),.Y(wire59_0_2));
NANDC2x1 inst_and_b59_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire59_0_3));
INVC inst_inv_b59_0_3 (.A(imd_wire59_0_3),.Y(wire59_0_3));
NANDC2x1 inst_and_b59_1_0 (.A(wire59_0_0),.B(wire59_0_1),.Y(imd_wire59_1_0));
INVC inst_inv_b59_1_0 (.A(imd_wire59_1_0),.Y(wire59_1_0));
NANDC2x1 inst_and_b59_1_1 (.A(wire59_0_2),.B(wire59_0_3),.Y(imd_wire59_1_1));
INVC inst_inv_b59_1_1 (.A(imd_wire59_1_1),.Y(wire59_1_1));
NANDC2x1 inst_and_b59_2_0 (.A(wire59_1_0),.B(wire59_1_1),.Y(imd_Y59));
INVC inst_inv_b59_2_0 (.A(imd_Y59),.Y(Y59));
NANDC2x1 inst_clockedAND_b59_59 (.A(CLK),.B(Y59),.Y(imd_YF59));
INVC inst_clockedinv_b59_59 (.A(imd_YF59),.Y(YF59));


NANDC2x1 inst_and_b60_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire60_0_0));
INVC inst_inv_b60_0_0 (.A(imd_wire60_0_0),.Y(wire60_0_0));
NANDC2x1 inst_and_b60_0_1 (.A(A2),.B(A3),.Y(imd_wire60_0_1));
INVC inst_inv_b60_0_1 (.A(imd_wire60_0_1),.Y(wire60_0_1));
NANDC2x1 inst_and_b60_0_2 (.A(A4),.B(A5),.Y(imd_wire60_0_2));
INVC inst_inv_b60_0_2 (.A(imd_wire60_0_2),.Y(wire60_0_2));
NANDC2x1 inst_and_b60_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire60_0_3));
INVC inst_inv_b60_0_3 (.A(imd_wire60_0_3),.Y(wire60_0_3));
NANDC2x1 inst_and_b60_1_0 (.A(wire60_0_0),.B(wire60_0_1),.Y(imd_wire60_1_0));
INVC inst_inv_b60_1_0 (.A(imd_wire60_1_0),.Y(wire60_1_0));
NANDC2x1 inst_and_b60_1_1 (.A(wire60_0_2),.B(wire60_0_3),.Y(imd_wire60_1_1));
INVC inst_inv_b60_1_1 (.A(imd_wire60_1_1),.Y(wire60_1_1));
NANDC2x1 inst_and_b60_2_0 (.A(wire60_1_0),.B(wire60_1_1),.Y(imd_Y60));
INVC inst_inv_b60_2_0 (.A(imd_Y60),.Y(Y60));
NANDC2x1 inst_clockedAND_b60_60 (.A(CLK),.B(Y60),.Y(imd_YF60));
INVC inst_clockedinv_b60_60 (.A(imd_YF60),.Y(YF60));


NANDC2x1 inst_and_b61_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire61_0_0));
INVC inst_inv_b61_0_0 (.A(imd_wire61_0_0),.Y(wire61_0_0));
NANDC2x1 inst_and_b61_0_1 (.A(A2),.B(A3),.Y(imd_wire61_0_1));
INVC inst_inv_b61_0_1 (.A(imd_wire61_0_1),.Y(wire61_0_1));
NANDC2x1 inst_and_b61_0_2 (.A(A4),.B(A5),.Y(imd_wire61_0_2));
INVC inst_inv_b61_0_2 (.A(imd_wire61_0_2),.Y(wire61_0_2));
NANDC2x1 inst_and_b61_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire61_0_3));
INVC inst_inv_b61_0_3 (.A(imd_wire61_0_3),.Y(wire61_0_3));
NANDC2x1 inst_and_b61_1_0 (.A(wire61_0_0),.B(wire61_0_1),.Y(imd_wire61_1_0));
INVC inst_inv_b61_1_0 (.A(imd_wire61_1_0),.Y(wire61_1_0));
NANDC2x1 inst_and_b61_1_1 (.A(wire61_0_2),.B(wire61_0_3),.Y(imd_wire61_1_1));
INVC inst_inv_b61_1_1 (.A(imd_wire61_1_1),.Y(wire61_1_1));
NANDC2x1 inst_and_b61_2_0 (.A(wire61_1_0),.B(wire61_1_1),.Y(imd_Y61));
INVC inst_inv_b61_2_0 (.A(imd_Y61),.Y(Y61));
NANDC2x1 inst_clockedAND_b61_61 (.A(CLK),.B(Y61),.Y(imd_YF61));
INVC inst_clockedinv_b61_61 (.A(imd_YF61),.Y(YF61));


NANDC2x1 inst_and_b62_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire62_0_0));
INVC inst_inv_b62_0_0 (.A(imd_wire62_0_0),.Y(wire62_0_0));
NANDC2x1 inst_and_b62_0_1 (.A(A2),.B(A3),.Y(imd_wire62_0_1));
INVC inst_inv_b62_0_1 (.A(imd_wire62_0_1),.Y(wire62_0_1));
NANDC2x1 inst_and_b62_0_2 (.A(A4),.B(A5),.Y(imd_wire62_0_2));
INVC inst_inv_b62_0_2 (.A(imd_wire62_0_2),.Y(wire62_0_2));
NANDC2x1 inst_and_b62_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire62_0_3));
INVC inst_inv_b62_0_3 (.A(imd_wire62_0_3),.Y(wire62_0_3));
NANDC2x1 inst_and_b62_1_0 (.A(wire62_0_0),.B(wire62_0_1),.Y(imd_wire62_1_0));
INVC inst_inv_b62_1_0 (.A(imd_wire62_1_0),.Y(wire62_1_0));
NANDC2x1 inst_and_b62_1_1 (.A(wire62_0_2),.B(wire62_0_3),.Y(imd_wire62_1_1));
INVC inst_inv_b62_1_1 (.A(imd_wire62_1_1),.Y(wire62_1_1));
NANDC2x1 inst_and_b62_2_0 (.A(wire62_1_0),.B(wire62_1_1),.Y(imd_Y62));
INVC inst_inv_b62_2_0 (.A(imd_Y62),.Y(Y62));
NANDC2x1 inst_clockedAND_b62_62 (.A(CLK),.B(Y62),.Y(imd_YF62));
INVC inst_clockedinv_b62_62 (.A(imd_YF62),.Y(YF62));


NANDC2x1 inst_and_b63_0_0 (.A(A0),.B(A1),.Y(imd_wire63_0_0));
INVC inst_inv_b63_0_0 (.A(imd_wire63_0_0),.Y(wire63_0_0));
NANDC2x1 inst_and_b63_0_1 (.A(A2),.B(A3),.Y(imd_wire63_0_1));
INVC inst_inv_b63_0_1 (.A(imd_wire63_0_1),.Y(wire63_0_1));
NANDC2x1 inst_and_b63_0_2 (.A(A4),.B(A5),.Y(imd_wire63_0_2));
INVC inst_inv_b63_0_2 (.A(imd_wire63_0_2),.Y(wire63_0_2));
NANDC2x1 inst_and_b63_0_3 (.A(A6_inv),.B(A7_inv),.Y(imd_wire63_0_3));
INVC inst_inv_b63_0_3 (.A(imd_wire63_0_3),.Y(wire63_0_3));
NANDC2x1 inst_and_b63_1_0 (.A(wire63_0_0),.B(wire63_0_1),.Y(imd_wire63_1_0));
INVC inst_inv_b63_1_0 (.A(imd_wire63_1_0),.Y(wire63_1_0));
NANDC2x1 inst_and_b63_1_1 (.A(wire63_0_2),.B(wire63_0_3),.Y(imd_wire63_1_1));
INVC inst_inv_b63_1_1 (.A(imd_wire63_1_1),.Y(wire63_1_1));
NANDC2x1 inst_and_b63_2_0 (.A(wire63_1_0),.B(wire63_1_1),.Y(imd_Y63));
INVC inst_inv_b63_2_0 (.A(imd_Y63),.Y(Y63));
NANDC2x1 inst_clockedAND_b63_63 (.A(CLK),.B(Y63),.Y(imd_YF63));
INVC inst_clockedinv_b63_63 (.A(imd_YF63),.Y(YF63));


NANDC2x1 inst_and_b64_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire64_0_0));
INVC inst_inv_b64_0_0 (.A(imd_wire64_0_0),.Y(wire64_0_0));
NANDC2x1 inst_and_b64_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire64_0_1));
INVC inst_inv_b64_0_1 (.A(imd_wire64_0_1),.Y(wire64_0_1));
NANDC2x1 inst_and_b64_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire64_0_2));
INVC inst_inv_b64_0_2 (.A(imd_wire64_0_2),.Y(wire64_0_2));
NANDC2x1 inst_and_b64_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire64_0_3));
INVC inst_inv_b64_0_3 (.A(imd_wire64_0_3),.Y(wire64_0_3));
NANDC2x1 inst_and_b64_1_0 (.A(wire64_0_0),.B(wire64_0_1),.Y(imd_wire64_1_0));
INVC inst_inv_b64_1_0 (.A(imd_wire64_1_0),.Y(wire64_1_0));
NANDC2x1 inst_and_b64_1_1 (.A(wire64_0_2),.B(wire64_0_3),.Y(imd_wire64_1_1));
INVC inst_inv_b64_1_1 (.A(imd_wire64_1_1),.Y(wire64_1_1));
NANDC2x1 inst_and_b64_2_0 (.A(wire64_1_0),.B(wire64_1_1),.Y(imd_Y64));
INVC inst_inv_b64_2_0 (.A(imd_Y64),.Y(Y64));
NANDC2x1 inst_clockedAND_b64_64 (.A(CLK),.B(Y64),.Y(imd_YF64));
INVC inst_clockedinv_b64_64 (.A(imd_YF64),.Y(YF64));


NANDC2x1 inst_and_b65_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire65_0_0));
INVC inst_inv_b65_0_0 (.A(imd_wire65_0_0),.Y(wire65_0_0));
NANDC2x1 inst_and_b65_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire65_0_1));
INVC inst_inv_b65_0_1 (.A(imd_wire65_0_1),.Y(wire65_0_1));
NANDC2x1 inst_and_b65_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire65_0_2));
INVC inst_inv_b65_0_2 (.A(imd_wire65_0_2),.Y(wire65_0_2));
NANDC2x1 inst_and_b65_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire65_0_3));
INVC inst_inv_b65_0_3 (.A(imd_wire65_0_3),.Y(wire65_0_3));
NANDC2x1 inst_and_b65_1_0 (.A(wire65_0_0),.B(wire65_0_1),.Y(imd_wire65_1_0));
INVC inst_inv_b65_1_0 (.A(imd_wire65_1_0),.Y(wire65_1_0));
NANDC2x1 inst_and_b65_1_1 (.A(wire65_0_2),.B(wire65_0_3),.Y(imd_wire65_1_1));
INVC inst_inv_b65_1_1 (.A(imd_wire65_1_1),.Y(wire65_1_1));
NANDC2x1 inst_and_b65_2_0 (.A(wire65_1_0),.B(wire65_1_1),.Y(imd_Y65));
INVC inst_inv_b65_2_0 (.A(imd_Y65),.Y(Y65));
NANDC2x1 inst_clockedAND_b65_65 (.A(CLK),.B(Y65),.Y(imd_YF65));
INVC inst_clockedinv_b65_65 (.A(imd_YF65),.Y(YF65));


NANDC2x1 inst_and_b66_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire66_0_0));
INVC inst_inv_b66_0_0 (.A(imd_wire66_0_0),.Y(wire66_0_0));
NANDC2x1 inst_and_b66_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire66_0_1));
INVC inst_inv_b66_0_1 (.A(imd_wire66_0_1),.Y(wire66_0_1));
NANDC2x1 inst_and_b66_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire66_0_2));
INVC inst_inv_b66_0_2 (.A(imd_wire66_0_2),.Y(wire66_0_2));
NANDC2x1 inst_and_b66_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire66_0_3));
INVC inst_inv_b66_0_3 (.A(imd_wire66_0_3),.Y(wire66_0_3));
NANDC2x1 inst_and_b66_1_0 (.A(wire66_0_0),.B(wire66_0_1),.Y(imd_wire66_1_0));
INVC inst_inv_b66_1_0 (.A(imd_wire66_1_0),.Y(wire66_1_0));
NANDC2x1 inst_and_b66_1_1 (.A(wire66_0_2),.B(wire66_0_3),.Y(imd_wire66_1_1));
INVC inst_inv_b66_1_1 (.A(imd_wire66_1_1),.Y(wire66_1_1));
NANDC2x1 inst_and_b66_2_0 (.A(wire66_1_0),.B(wire66_1_1),.Y(imd_Y66));
INVC inst_inv_b66_2_0 (.A(imd_Y66),.Y(Y66));
NANDC2x1 inst_clockedAND_b66_66 (.A(CLK),.B(Y66),.Y(imd_YF66));
INVC inst_clockedinv_b66_66 (.A(imd_YF66),.Y(YF66));


NANDC2x1 inst_and_b67_0_0 (.A(A0),.B(A1),.Y(imd_wire67_0_0));
INVC inst_inv_b67_0_0 (.A(imd_wire67_0_0),.Y(wire67_0_0));
NANDC2x1 inst_and_b67_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire67_0_1));
INVC inst_inv_b67_0_1 (.A(imd_wire67_0_1),.Y(wire67_0_1));
NANDC2x1 inst_and_b67_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire67_0_2));
INVC inst_inv_b67_0_2 (.A(imd_wire67_0_2),.Y(wire67_0_2));
NANDC2x1 inst_and_b67_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire67_0_3));
INVC inst_inv_b67_0_3 (.A(imd_wire67_0_3),.Y(wire67_0_3));
NANDC2x1 inst_and_b67_1_0 (.A(wire67_0_0),.B(wire67_0_1),.Y(imd_wire67_1_0));
INVC inst_inv_b67_1_0 (.A(imd_wire67_1_0),.Y(wire67_1_0));
NANDC2x1 inst_and_b67_1_1 (.A(wire67_0_2),.B(wire67_0_3),.Y(imd_wire67_1_1));
INVC inst_inv_b67_1_1 (.A(imd_wire67_1_1),.Y(wire67_1_1));
NANDC2x1 inst_and_b67_2_0 (.A(wire67_1_0),.B(wire67_1_1),.Y(imd_Y67));
INVC inst_inv_b67_2_0 (.A(imd_Y67),.Y(Y67));
NANDC2x1 inst_clockedAND_b67_67 (.A(CLK),.B(Y67),.Y(imd_YF67));
INVC inst_clockedinv_b67_67 (.A(imd_YF67),.Y(YF67));


NANDC2x1 inst_and_b68_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire68_0_0));
INVC inst_inv_b68_0_0 (.A(imd_wire68_0_0),.Y(wire68_0_0));
NANDC2x1 inst_and_b68_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire68_0_1));
INVC inst_inv_b68_0_1 (.A(imd_wire68_0_1),.Y(wire68_0_1));
NANDC2x1 inst_and_b68_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire68_0_2));
INVC inst_inv_b68_0_2 (.A(imd_wire68_0_2),.Y(wire68_0_2));
NANDC2x1 inst_and_b68_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire68_0_3));
INVC inst_inv_b68_0_3 (.A(imd_wire68_0_3),.Y(wire68_0_3));
NANDC2x1 inst_and_b68_1_0 (.A(wire68_0_0),.B(wire68_0_1),.Y(imd_wire68_1_0));
INVC inst_inv_b68_1_0 (.A(imd_wire68_1_0),.Y(wire68_1_0));
NANDC2x1 inst_and_b68_1_1 (.A(wire68_0_2),.B(wire68_0_3),.Y(imd_wire68_1_1));
INVC inst_inv_b68_1_1 (.A(imd_wire68_1_1),.Y(wire68_1_1));
NANDC2x1 inst_and_b68_2_0 (.A(wire68_1_0),.B(wire68_1_1),.Y(imd_Y68));
INVC inst_inv_b68_2_0 (.A(imd_Y68),.Y(Y68));
NANDC2x1 inst_clockedAND_b68_68 (.A(CLK),.B(Y68),.Y(imd_YF68));
INVC inst_clockedinv_b68_68 (.A(imd_YF68),.Y(YF68));


NANDC2x1 inst_and_b69_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire69_0_0));
INVC inst_inv_b69_0_0 (.A(imd_wire69_0_0),.Y(wire69_0_0));
NANDC2x1 inst_and_b69_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire69_0_1));
INVC inst_inv_b69_0_1 (.A(imd_wire69_0_1),.Y(wire69_0_1));
NANDC2x1 inst_and_b69_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire69_0_2));
INVC inst_inv_b69_0_2 (.A(imd_wire69_0_2),.Y(wire69_0_2));
NANDC2x1 inst_and_b69_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire69_0_3));
INVC inst_inv_b69_0_3 (.A(imd_wire69_0_3),.Y(wire69_0_3));
NANDC2x1 inst_and_b69_1_0 (.A(wire69_0_0),.B(wire69_0_1),.Y(imd_wire69_1_0));
INVC inst_inv_b69_1_0 (.A(imd_wire69_1_0),.Y(wire69_1_0));
NANDC2x1 inst_and_b69_1_1 (.A(wire69_0_2),.B(wire69_0_3),.Y(imd_wire69_1_1));
INVC inst_inv_b69_1_1 (.A(imd_wire69_1_1),.Y(wire69_1_1));
NANDC2x1 inst_and_b69_2_0 (.A(wire69_1_0),.B(wire69_1_1),.Y(imd_Y69));
INVC inst_inv_b69_2_0 (.A(imd_Y69),.Y(Y69));
NANDC2x1 inst_clockedAND_b69_69 (.A(CLK),.B(Y69),.Y(imd_YF69));
INVC inst_clockedinv_b69_69 (.A(imd_YF69),.Y(YF69));


NANDC2x1 inst_and_b70_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire70_0_0));
INVC inst_inv_b70_0_0 (.A(imd_wire70_0_0),.Y(wire70_0_0));
NANDC2x1 inst_and_b70_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire70_0_1));
INVC inst_inv_b70_0_1 (.A(imd_wire70_0_1),.Y(wire70_0_1));
NANDC2x1 inst_and_b70_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire70_0_2));
INVC inst_inv_b70_0_2 (.A(imd_wire70_0_2),.Y(wire70_0_2));
NANDC2x1 inst_and_b70_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire70_0_3));
INVC inst_inv_b70_0_3 (.A(imd_wire70_0_3),.Y(wire70_0_3));
NANDC2x1 inst_and_b70_1_0 (.A(wire70_0_0),.B(wire70_0_1),.Y(imd_wire70_1_0));
INVC inst_inv_b70_1_0 (.A(imd_wire70_1_0),.Y(wire70_1_0));
NANDC2x1 inst_and_b70_1_1 (.A(wire70_0_2),.B(wire70_0_3),.Y(imd_wire70_1_1));
INVC inst_inv_b70_1_1 (.A(imd_wire70_1_1),.Y(wire70_1_1));
NANDC2x1 inst_and_b70_2_0 (.A(wire70_1_0),.B(wire70_1_1),.Y(imd_Y70));
INVC inst_inv_b70_2_0 (.A(imd_Y70),.Y(Y70));
NANDC2x1 inst_clockedAND_b70_70 (.A(CLK),.B(Y70),.Y(imd_YF70));
INVC inst_clockedinv_b70_70 (.A(imd_YF70),.Y(YF70));


NANDC2x1 inst_and_b71_0_0 (.A(A0),.B(A1),.Y(imd_wire71_0_0));
INVC inst_inv_b71_0_0 (.A(imd_wire71_0_0),.Y(wire71_0_0));
NANDC2x1 inst_and_b71_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire71_0_1));
INVC inst_inv_b71_0_1 (.A(imd_wire71_0_1),.Y(wire71_0_1));
NANDC2x1 inst_and_b71_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire71_0_2));
INVC inst_inv_b71_0_2 (.A(imd_wire71_0_2),.Y(wire71_0_2));
NANDC2x1 inst_and_b71_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire71_0_3));
INVC inst_inv_b71_0_3 (.A(imd_wire71_0_3),.Y(wire71_0_3));
NANDC2x1 inst_and_b71_1_0 (.A(wire71_0_0),.B(wire71_0_1),.Y(imd_wire71_1_0));
INVC inst_inv_b71_1_0 (.A(imd_wire71_1_0),.Y(wire71_1_0));
NANDC2x1 inst_and_b71_1_1 (.A(wire71_0_2),.B(wire71_0_3),.Y(imd_wire71_1_1));
INVC inst_inv_b71_1_1 (.A(imd_wire71_1_1),.Y(wire71_1_1));
NANDC2x1 inst_and_b71_2_0 (.A(wire71_1_0),.B(wire71_1_1),.Y(imd_Y71));
INVC inst_inv_b71_2_0 (.A(imd_Y71),.Y(Y71));
NANDC2x1 inst_clockedAND_b71_71 (.A(CLK),.B(Y71),.Y(imd_YF71));
INVC inst_clockedinv_b71_71 (.A(imd_YF71),.Y(YF71));


NANDC2x1 inst_and_b72_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire72_0_0));
INVC inst_inv_b72_0_0 (.A(imd_wire72_0_0),.Y(wire72_0_0));
NANDC2x1 inst_and_b72_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire72_0_1));
INVC inst_inv_b72_0_1 (.A(imd_wire72_0_1),.Y(wire72_0_1));
NANDC2x1 inst_and_b72_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire72_0_2));
INVC inst_inv_b72_0_2 (.A(imd_wire72_0_2),.Y(wire72_0_2));
NANDC2x1 inst_and_b72_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire72_0_3));
INVC inst_inv_b72_0_3 (.A(imd_wire72_0_3),.Y(wire72_0_3));
NANDC2x1 inst_and_b72_1_0 (.A(wire72_0_0),.B(wire72_0_1),.Y(imd_wire72_1_0));
INVC inst_inv_b72_1_0 (.A(imd_wire72_1_0),.Y(wire72_1_0));
NANDC2x1 inst_and_b72_1_1 (.A(wire72_0_2),.B(wire72_0_3),.Y(imd_wire72_1_1));
INVC inst_inv_b72_1_1 (.A(imd_wire72_1_1),.Y(wire72_1_1));
NANDC2x1 inst_and_b72_2_0 (.A(wire72_1_0),.B(wire72_1_1),.Y(imd_Y72));
INVC inst_inv_b72_2_0 (.A(imd_Y72),.Y(Y72));
NANDC2x1 inst_clockedAND_b72_72 (.A(CLK),.B(Y72),.Y(imd_YF72));
INVC inst_clockedinv_b72_72 (.A(imd_YF72),.Y(YF72));


NANDC2x1 inst_and_b73_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire73_0_0));
INVC inst_inv_b73_0_0 (.A(imd_wire73_0_0),.Y(wire73_0_0));
NANDC2x1 inst_and_b73_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire73_0_1));
INVC inst_inv_b73_0_1 (.A(imd_wire73_0_1),.Y(wire73_0_1));
NANDC2x1 inst_and_b73_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire73_0_2));
INVC inst_inv_b73_0_2 (.A(imd_wire73_0_2),.Y(wire73_0_2));
NANDC2x1 inst_and_b73_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire73_0_3));
INVC inst_inv_b73_0_3 (.A(imd_wire73_0_3),.Y(wire73_0_3));
NANDC2x1 inst_and_b73_1_0 (.A(wire73_0_0),.B(wire73_0_1),.Y(imd_wire73_1_0));
INVC inst_inv_b73_1_0 (.A(imd_wire73_1_0),.Y(wire73_1_0));
NANDC2x1 inst_and_b73_1_1 (.A(wire73_0_2),.B(wire73_0_3),.Y(imd_wire73_1_1));
INVC inst_inv_b73_1_1 (.A(imd_wire73_1_1),.Y(wire73_1_1));
NANDC2x1 inst_and_b73_2_0 (.A(wire73_1_0),.B(wire73_1_1),.Y(imd_Y73));
INVC inst_inv_b73_2_0 (.A(imd_Y73),.Y(Y73));
NANDC2x1 inst_clockedAND_b73_73 (.A(CLK),.B(Y73),.Y(imd_YF73));
INVC inst_clockedinv_b73_73 (.A(imd_YF73),.Y(YF73));


NANDC2x1 inst_and_b74_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire74_0_0));
INVC inst_inv_b74_0_0 (.A(imd_wire74_0_0),.Y(wire74_0_0));
NANDC2x1 inst_and_b74_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire74_0_1));
INVC inst_inv_b74_0_1 (.A(imd_wire74_0_1),.Y(wire74_0_1));
NANDC2x1 inst_and_b74_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire74_0_2));
INVC inst_inv_b74_0_2 (.A(imd_wire74_0_2),.Y(wire74_0_2));
NANDC2x1 inst_and_b74_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire74_0_3));
INVC inst_inv_b74_0_3 (.A(imd_wire74_0_3),.Y(wire74_0_3));
NANDC2x1 inst_and_b74_1_0 (.A(wire74_0_0),.B(wire74_0_1),.Y(imd_wire74_1_0));
INVC inst_inv_b74_1_0 (.A(imd_wire74_1_0),.Y(wire74_1_0));
NANDC2x1 inst_and_b74_1_1 (.A(wire74_0_2),.B(wire74_0_3),.Y(imd_wire74_1_1));
INVC inst_inv_b74_1_1 (.A(imd_wire74_1_1),.Y(wire74_1_1));
NANDC2x1 inst_and_b74_2_0 (.A(wire74_1_0),.B(wire74_1_1),.Y(imd_Y74));
INVC inst_inv_b74_2_0 (.A(imd_Y74),.Y(Y74));
NANDC2x1 inst_clockedAND_b74_74 (.A(CLK),.B(Y74),.Y(imd_YF74));
INVC inst_clockedinv_b74_74 (.A(imd_YF74),.Y(YF74));


NANDC2x1 inst_and_b75_0_0 (.A(A0),.B(A1),.Y(imd_wire75_0_0));
INVC inst_inv_b75_0_0 (.A(imd_wire75_0_0),.Y(wire75_0_0));
NANDC2x1 inst_and_b75_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire75_0_1));
INVC inst_inv_b75_0_1 (.A(imd_wire75_0_1),.Y(wire75_0_1));
NANDC2x1 inst_and_b75_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire75_0_2));
INVC inst_inv_b75_0_2 (.A(imd_wire75_0_2),.Y(wire75_0_2));
NANDC2x1 inst_and_b75_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire75_0_3));
INVC inst_inv_b75_0_3 (.A(imd_wire75_0_3),.Y(wire75_0_3));
NANDC2x1 inst_and_b75_1_0 (.A(wire75_0_0),.B(wire75_0_1),.Y(imd_wire75_1_0));
INVC inst_inv_b75_1_0 (.A(imd_wire75_1_0),.Y(wire75_1_0));
NANDC2x1 inst_and_b75_1_1 (.A(wire75_0_2),.B(wire75_0_3),.Y(imd_wire75_1_1));
INVC inst_inv_b75_1_1 (.A(imd_wire75_1_1),.Y(wire75_1_1));
NANDC2x1 inst_and_b75_2_0 (.A(wire75_1_0),.B(wire75_1_1),.Y(imd_Y75));
INVC inst_inv_b75_2_0 (.A(imd_Y75),.Y(Y75));
NANDC2x1 inst_clockedAND_b75_75 (.A(CLK),.B(Y75),.Y(imd_YF75));
INVC inst_clockedinv_b75_75 (.A(imd_YF75),.Y(YF75));


NANDC2x1 inst_and_b76_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire76_0_0));
INVC inst_inv_b76_0_0 (.A(imd_wire76_0_0),.Y(wire76_0_0));
NANDC2x1 inst_and_b76_0_1 (.A(A2),.B(A3),.Y(imd_wire76_0_1));
INVC inst_inv_b76_0_1 (.A(imd_wire76_0_1),.Y(wire76_0_1));
NANDC2x1 inst_and_b76_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire76_0_2));
INVC inst_inv_b76_0_2 (.A(imd_wire76_0_2),.Y(wire76_0_2));
NANDC2x1 inst_and_b76_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire76_0_3));
INVC inst_inv_b76_0_3 (.A(imd_wire76_0_3),.Y(wire76_0_3));
NANDC2x1 inst_and_b76_1_0 (.A(wire76_0_0),.B(wire76_0_1),.Y(imd_wire76_1_0));
INVC inst_inv_b76_1_0 (.A(imd_wire76_1_0),.Y(wire76_1_0));
NANDC2x1 inst_and_b76_1_1 (.A(wire76_0_2),.B(wire76_0_3),.Y(imd_wire76_1_1));
INVC inst_inv_b76_1_1 (.A(imd_wire76_1_1),.Y(wire76_1_1));
NANDC2x1 inst_and_b76_2_0 (.A(wire76_1_0),.B(wire76_1_1),.Y(imd_Y76));
INVC inst_inv_b76_2_0 (.A(imd_Y76),.Y(Y76));
NANDC2x1 inst_clockedAND_b76_76 (.A(CLK),.B(Y76),.Y(imd_YF76));
INVC inst_clockedinv_b76_76 (.A(imd_YF76),.Y(YF76));


NANDC2x1 inst_and_b77_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire77_0_0));
INVC inst_inv_b77_0_0 (.A(imd_wire77_0_0),.Y(wire77_0_0));
NANDC2x1 inst_and_b77_0_1 (.A(A2),.B(A3),.Y(imd_wire77_0_1));
INVC inst_inv_b77_0_1 (.A(imd_wire77_0_1),.Y(wire77_0_1));
NANDC2x1 inst_and_b77_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire77_0_2));
INVC inst_inv_b77_0_2 (.A(imd_wire77_0_2),.Y(wire77_0_2));
NANDC2x1 inst_and_b77_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire77_0_3));
INVC inst_inv_b77_0_3 (.A(imd_wire77_0_3),.Y(wire77_0_3));
NANDC2x1 inst_and_b77_1_0 (.A(wire77_0_0),.B(wire77_0_1),.Y(imd_wire77_1_0));
INVC inst_inv_b77_1_0 (.A(imd_wire77_1_0),.Y(wire77_1_0));
NANDC2x1 inst_and_b77_1_1 (.A(wire77_0_2),.B(wire77_0_3),.Y(imd_wire77_1_1));
INVC inst_inv_b77_1_1 (.A(imd_wire77_1_1),.Y(wire77_1_1));
NANDC2x1 inst_and_b77_2_0 (.A(wire77_1_0),.B(wire77_1_1),.Y(imd_Y77));
INVC inst_inv_b77_2_0 (.A(imd_Y77),.Y(Y77));
NANDC2x1 inst_clockedAND_b77_77 (.A(CLK),.B(Y77),.Y(imd_YF77));
INVC inst_clockedinv_b77_77 (.A(imd_YF77),.Y(YF77));


NANDC2x1 inst_and_b78_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire78_0_0));
INVC inst_inv_b78_0_0 (.A(imd_wire78_0_0),.Y(wire78_0_0));
NANDC2x1 inst_and_b78_0_1 (.A(A2),.B(A3),.Y(imd_wire78_0_1));
INVC inst_inv_b78_0_1 (.A(imd_wire78_0_1),.Y(wire78_0_1));
NANDC2x1 inst_and_b78_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire78_0_2));
INVC inst_inv_b78_0_2 (.A(imd_wire78_0_2),.Y(wire78_0_2));
NANDC2x1 inst_and_b78_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire78_0_3));
INVC inst_inv_b78_0_3 (.A(imd_wire78_0_3),.Y(wire78_0_3));
NANDC2x1 inst_and_b78_1_0 (.A(wire78_0_0),.B(wire78_0_1),.Y(imd_wire78_1_0));
INVC inst_inv_b78_1_0 (.A(imd_wire78_1_0),.Y(wire78_1_0));
NANDC2x1 inst_and_b78_1_1 (.A(wire78_0_2),.B(wire78_0_3),.Y(imd_wire78_1_1));
INVC inst_inv_b78_1_1 (.A(imd_wire78_1_1),.Y(wire78_1_1));
NANDC2x1 inst_and_b78_2_0 (.A(wire78_1_0),.B(wire78_1_1),.Y(imd_Y78));
INVC inst_inv_b78_2_0 (.A(imd_Y78),.Y(Y78));
NANDC2x1 inst_clockedAND_b78_78 (.A(CLK),.B(Y78),.Y(imd_YF78));
INVC inst_clockedinv_b78_78 (.A(imd_YF78),.Y(YF78));


NANDC2x1 inst_and_b79_0_0 (.A(A0),.B(A1),.Y(imd_wire79_0_0));
INVC inst_inv_b79_0_0 (.A(imd_wire79_0_0),.Y(wire79_0_0));
NANDC2x1 inst_and_b79_0_1 (.A(A2),.B(A3),.Y(imd_wire79_0_1));
INVC inst_inv_b79_0_1 (.A(imd_wire79_0_1),.Y(wire79_0_1));
NANDC2x1 inst_and_b79_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire79_0_2));
INVC inst_inv_b79_0_2 (.A(imd_wire79_0_2),.Y(wire79_0_2));
NANDC2x1 inst_and_b79_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire79_0_3));
INVC inst_inv_b79_0_3 (.A(imd_wire79_0_3),.Y(wire79_0_3));
NANDC2x1 inst_and_b79_1_0 (.A(wire79_0_0),.B(wire79_0_1),.Y(imd_wire79_1_0));
INVC inst_inv_b79_1_0 (.A(imd_wire79_1_0),.Y(wire79_1_0));
NANDC2x1 inst_and_b79_1_1 (.A(wire79_0_2),.B(wire79_0_3),.Y(imd_wire79_1_1));
INVC inst_inv_b79_1_1 (.A(imd_wire79_1_1),.Y(wire79_1_1));
NANDC2x1 inst_and_b79_2_0 (.A(wire79_1_0),.B(wire79_1_1),.Y(imd_Y79));
INVC inst_inv_b79_2_0 (.A(imd_Y79),.Y(Y79));
NANDC2x1 inst_clockedAND_b79_79 (.A(CLK),.B(Y79),.Y(imd_YF79));
INVC inst_clockedinv_b79_79 (.A(imd_YF79),.Y(YF79));


NANDC2x1 inst_and_b80_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire80_0_0));
INVC inst_inv_b80_0_0 (.A(imd_wire80_0_0),.Y(wire80_0_0));
NANDC2x1 inst_and_b80_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire80_0_1));
INVC inst_inv_b80_0_1 (.A(imd_wire80_0_1),.Y(wire80_0_1));
NANDC2x1 inst_and_b80_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire80_0_2));
INVC inst_inv_b80_0_2 (.A(imd_wire80_0_2),.Y(wire80_0_2));
NANDC2x1 inst_and_b80_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire80_0_3));
INVC inst_inv_b80_0_3 (.A(imd_wire80_0_3),.Y(wire80_0_3));
NANDC2x1 inst_and_b80_1_0 (.A(wire80_0_0),.B(wire80_0_1),.Y(imd_wire80_1_0));
INVC inst_inv_b80_1_0 (.A(imd_wire80_1_0),.Y(wire80_1_0));
NANDC2x1 inst_and_b80_1_1 (.A(wire80_0_2),.B(wire80_0_3),.Y(imd_wire80_1_1));
INVC inst_inv_b80_1_1 (.A(imd_wire80_1_1),.Y(wire80_1_1));
NANDC2x1 inst_and_b80_2_0 (.A(wire80_1_0),.B(wire80_1_1),.Y(imd_Y80));
INVC inst_inv_b80_2_0 (.A(imd_Y80),.Y(Y80));
NANDC2x1 inst_clockedAND_b80_80 (.A(CLK),.B(Y80),.Y(imd_YF80));
INVC inst_clockedinv_b80_80 (.A(imd_YF80),.Y(YF80));


NANDC2x1 inst_and_b81_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire81_0_0));
INVC inst_inv_b81_0_0 (.A(imd_wire81_0_0),.Y(wire81_0_0));
NANDC2x1 inst_and_b81_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire81_0_1));
INVC inst_inv_b81_0_1 (.A(imd_wire81_0_1),.Y(wire81_0_1));
NANDC2x1 inst_and_b81_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire81_0_2));
INVC inst_inv_b81_0_2 (.A(imd_wire81_0_2),.Y(wire81_0_2));
NANDC2x1 inst_and_b81_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire81_0_3));
INVC inst_inv_b81_0_3 (.A(imd_wire81_0_3),.Y(wire81_0_3));
NANDC2x1 inst_and_b81_1_0 (.A(wire81_0_0),.B(wire81_0_1),.Y(imd_wire81_1_0));
INVC inst_inv_b81_1_0 (.A(imd_wire81_1_0),.Y(wire81_1_0));
NANDC2x1 inst_and_b81_1_1 (.A(wire81_0_2),.B(wire81_0_3),.Y(imd_wire81_1_1));
INVC inst_inv_b81_1_1 (.A(imd_wire81_1_1),.Y(wire81_1_1));
NANDC2x1 inst_and_b81_2_0 (.A(wire81_1_0),.B(wire81_1_1),.Y(imd_Y81));
INVC inst_inv_b81_2_0 (.A(imd_Y81),.Y(Y81));
NANDC2x1 inst_clockedAND_b81_81 (.A(CLK),.B(Y81),.Y(imd_YF81));
INVC inst_clockedinv_b81_81 (.A(imd_YF81),.Y(YF81));


NANDC2x1 inst_and_b82_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire82_0_0));
INVC inst_inv_b82_0_0 (.A(imd_wire82_0_0),.Y(wire82_0_0));
NANDC2x1 inst_and_b82_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire82_0_1));
INVC inst_inv_b82_0_1 (.A(imd_wire82_0_1),.Y(wire82_0_1));
NANDC2x1 inst_and_b82_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire82_0_2));
INVC inst_inv_b82_0_2 (.A(imd_wire82_0_2),.Y(wire82_0_2));
NANDC2x1 inst_and_b82_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire82_0_3));
INVC inst_inv_b82_0_3 (.A(imd_wire82_0_3),.Y(wire82_0_3));
NANDC2x1 inst_and_b82_1_0 (.A(wire82_0_0),.B(wire82_0_1),.Y(imd_wire82_1_0));
INVC inst_inv_b82_1_0 (.A(imd_wire82_1_0),.Y(wire82_1_0));
NANDC2x1 inst_and_b82_1_1 (.A(wire82_0_2),.B(wire82_0_3),.Y(imd_wire82_1_1));
INVC inst_inv_b82_1_1 (.A(imd_wire82_1_1),.Y(wire82_1_1));
NANDC2x1 inst_and_b82_2_0 (.A(wire82_1_0),.B(wire82_1_1),.Y(imd_Y82));
INVC inst_inv_b82_2_0 (.A(imd_Y82),.Y(Y82));
NANDC2x1 inst_clockedAND_b82_82 (.A(CLK),.B(Y82),.Y(imd_YF82));
INVC inst_clockedinv_b82_82 (.A(imd_YF82),.Y(YF82));


NANDC2x1 inst_and_b83_0_0 (.A(A0),.B(A1),.Y(imd_wire83_0_0));
INVC inst_inv_b83_0_0 (.A(imd_wire83_0_0),.Y(wire83_0_0));
NANDC2x1 inst_and_b83_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire83_0_1));
INVC inst_inv_b83_0_1 (.A(imd_wire83_0_1),.Y(wire83_0_1));
NANDC2x1 inst_and_b83_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire83_0_2));
INVC inst_inv_b83_0_2 (.A(imd_wire83_0_2),.Y(wire83_0_2));
NANDC2x1 inst_and_b83_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire83_0_3));
INVC inst_inv_b83_0_3 (.A(imd_wire83_0_3),.Y(wire83_0_3));
NANDC2x1 inst_and_b83_1_0 (.A(wire83_0_0),.B(wire83_0_1),.Y(imd_wire83_1_0));
INVC inst_inv_b83_1_0 (.A(imd_wire83_1_0),.Y(wire83_1_0));
NANDC2x1 inst_and_b83_1_1 (.A(wire83_0_2),.B(wire83_0_3),.Y(imd_wire83_1_1));
INVC inst_inv_b83_1_1 (.A(imd_wire83_1_1),.Y(wire83_1_1));
NANDC2x1 inst_and_b83_2_0 (.A(wire83_1_0),.B(wire83_1_1),.Y(imd_Y83));
INVC inst_inv_b83_2_0 (.A(imd_Y83),.Y(Y83));
NANDC2x1 inst_clockedAND_b83_83 (.A(CLK),.B(Y83),.Y(imd_YF83));
INVC inst_clockedinv_b83_83 (.A(imd_YF83),.Y(YF83));


NANDC2x1 inst_and_b84_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire84_0_0));
INVC inst_inv_b84_0_0 (.A(imd_wire84_0_0),.Y(wire84_0_0));
NANDC2x1 inst_and_b84_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire84_0_1));
INVC inst_inv_b84_0_1 (.A(imd_wire84_0_1),.Y(wire84_0_1));
NANDC2x1 inst_and_b84_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire84_0_2));
INVC inst_inv_b84_0_2 (.A(imd_wire84_0_2),.Y(wire84_0_2));
NANDC2x1 inst_and_b84_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire84_0_3));
INVC inst_inv_b84_0_3 (.A(imd_wire84_0_3),.Y(wire84_0_3));
NANDC2x1 inst_and_b84_1_0 (.A(wire84_0_0),.B(wire84_0_1),.Y(imd_wire84_1_0));
INVC inst_inv_b84_1_0 (.A(imd_wire84_1_0),.Y(wire84_1_0));
NANDC2x1 inst_and_b84_1_1 (.A(wire84_0_2),.B(wire84_0_3),.Y(imd_wire84_1_1));
INVC inst_inv_b84_1_1 (.A(imd_wire84_1_1),.Y(wire84_1_1));
NANDC2x1 inst_and_b84_2_0 (.A(wire84_1_0),.B(wire84_1_1),.Y(imd_Y84));
INVC inst_inv_b84_2_0 (.A(imd_Y84),.Y(Y84));
NANDC2x1 inst_clockedAND_b84_84 (.A(CLK),.B(Y84),.Y(imd_YF84));
INVC inst_clockedinv_b84_84 (.A(imd_YF84),.Y(YF84));


NANDC2x1 inst_and_b85_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire85_0_0));
INVC inst_inv_b85_0_0 (.A(imd_wire85_0_0),.Y(wire85_0_0));
NANDC2x1 inst_and_b85_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire85_0_1));
INVC inst_inv_b85_0_1 (.A(imd_wire85_0_1),.Y(wire85_0_1));
NANDC2x1 inst_and_b85_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire85_0_2));
INVC inst_inv_b85_0_2 (.A(imd_wire85_0_2),.Y(wire85_0_2));
NANDC2x1 inst_and_b85_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire85_0_3));
INVC inst_inv_b85_0_3 (.A(imd_wire85_0_3),.Y(wire85_0_3));
NANDC2x1 inst_and_b85_1_0 (.A(wire85_0_0),.B(wire85_0_1),.Y(imd_wire85_1_0));
INVC inst_inv_b85_1_0 (.A(imd_wire85_1_0),.Y(wire85_1_0));
NANDC2x1 inst_and_b85_1_1 (.A(wire85_0_2),.B(wire85_0_3),.Y(imd_wire85_1_1));
INVC inst_inv_b85_1_1 (.A(imd_wire85_1_1),.Y(wire85_1_1));
NANDC2x1 inst_and_b85_2_0 (.A(wire85_1_0),.B(wire85_1_1),.Y(imd_Y85));
INVC inst_inv_b85_2_0 (.A(imd_Y85),.Y(Y85));
NANDC2x1 inst_clockedAND_b85_85 (.A(CLK),.B(Y85),.Y(imd_YF85));
INVC inst_clockedinv_b85_85 (.A(imd_YF85),.Y(YF85));


NANDC2x1 inst_and_b86_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire86_0_0));
INVC inst_inv_b86_0_0 (.A(imd_wire86_0_0),.Y(wire86_0_0));
NANDC2x1 inst_and_b86_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire86_0_1));
INVC inst_inv_b86_0_1 (.A(imd_wire86_0_1),.Y(wire86_0_1));
NANDC2x1 inst_and_b86_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire86_0_2));
INVC inst_inv_b86_0_2 (.A(imd_wire86_0_2),.Y(wire86_0_2));
NANDC2x1 inst_and_b86_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire86_0_3));
INVC inst_inv_b86_0_3 (.A(imd_wire86_0_3),.Y(wire86_0_3));
NANDC2x1 inst_and_b86_1_0 (.A(wire86_0_0),.B(wire86_0_1),.Y(imd_wire86_1_0));
INVC inst_inv_b86_1_0 (.A(imd_wire86_1_0),.Y(wire86_1_0));
NANDC2x1 inst_and_b86_1_1 (.A(wire86_0_2),.B(wire86_0_3),.Y(imd_wire86_1_1));
INVC inst_inv_b86_1_1 (.A(imd_wire86_1_1),.Y(wire86_1_1));
NANDC2x1 inst_and_b86_2_0 (.A(wire86_1_0),.B(wire86_1_1),.Y(imd_Y86));
INVC inst_inv_b86_2_0 (.A(imd_Y86),.Y(Y86));
NANDC2x1 inst_clockedAND_b86_86 (.A(CLK),.B(Y86),.Y(imd_YF86));
INVC inst_clockedinv_b86_86 (.A(imd_YF86),.Y(YF86));


NANDC2x1 inst_and_b87_0_0 (.A(A0),.B(A1),.Y(imd_wire87_0_0));
INVC inst_inv_b87_0_0 (.A(imd_wire87_0_0),.Y(wire87_0_0));
NANDC2x1 inst_and_b87_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire87_0_1));
INVC inst_inv_b87_0_1 (.A(imd_wire87_0_1),.Y(wire87_0_1));
NANDC2x1 inst_and_b87_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire87_0_2));
INVC inst_inv_b87_0_2 (.A(imd_wire87_0_2),.Y(wire87_0_2));
NANDC2x1 inst_and_b87_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire87_0_3));
INVC inst_inv_b87_0_3 (.A(imd_wire87_0_3),.Y(wire87_0_3));
NANDC2x1 inst_and_b87_1_0 (.A(wire87_0_0),.B(wire87_0_1),.Y(imd_wire87_1_0));
INVC inst_inv_b87_1_0 (.A(imd_wire87_1_0),.Y(wire87_1_0));
NANDC2x1 inst_and_b87_1_1 (.A(wire87_0_2),.B(wire87_0_3),.Y(imd_wire87_1_1));
INVC inst_inv_b87_1_1 (.A(imd_wire87_1_1),.Y(wire87_1_1));
NANDC2x1 inst_and_b87_2_0 (.A(wire87_1_0),.B(wire87_1_1),.Y(imd_Y87));
INVC inst_inv_b87_2_0 (.A(imd_Y87),.Y(Y87));
NANDC2x1 inst_clockedAND_b87_87 (.A(CLK),.B(Y87),.Y(imd_YF87));
INVC inst_clockedinv_b87_87 (.A(imd_YF87),.Y(YF87));


NANDC2x1 inst_and_b88_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire88_0_0));
INVC inst_inv_b88_0_0 (.A(imd_wire88_0_0),.Y(wire88_0_0));
NANDC2x1 inst_and_b88_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire88_0_1));
INVC inst_inv_b88_0_1 (.A(imd_wire88_0_1),.Y(wire88_0_1));
NANDC2x1 inst_and_b88_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire88_0_2));
INVC inst_inv_b88_0_2 (.A(imd_wire88_0_2),.Y(wire88_0_2));
NANDC2x1 inst_and_b88_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire88_0_3));
INVC inst_inv_b88_0_3 (.A(imd_wire88_0_3),.Y(wire88_0_3));
NANDC2x1 inst_and_b88_1_0 (.A(wire88_0_0),.B(wire88_0_1),.Y(imd_wire88_1_0));
INVC inst_inv_b88_1_0 (.A(imd_wire88_1_0),.Y(wire88_1_0));
NANDC2x1 inst_and_b88_1_1 (.A(wire88_0_2),.B(wire88_0_3),.Y(imd_wire88_1_1));
INVC inst_inv_b88_1_1 (.A(imd_wire88_1_1),.Y(wire88_1_1));
NANDC2x1 inst_and_b88_2_0 (.A(wire88_1_0),.B(wire88_1_1),.Y(imd_Y88));
INVC inst_inv_b88_2_0 (.A(imd_Y88),.Y(Y88));
NANDC2x1 inst_clockedAND_b88_88 (.A(CLK),.B(Y88),.Y(imd_YF88));
INVC inst_clockedinv_b88_88 (.A(imd_YF88),.Y(YF88));


NANDC2x1 inst_and_b89_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire89_0_0));
INVC inst_inv_b89_0_0 (.A(imd_wire89_0_0),.Y(wire89_0_0));
NANDC2x1 inst_and_b89_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire89_0_1));
INVC inst_inv_b89_0_1 (.A(imd_wire89_0_1),.Y(wire89_0_1));
NANDC2x1 inst_and_b89_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire89_0_2));
INVC inst_inv_b89_0_2 (.A(imd_wire89_0_2),.Y(wire89_0_2));
NANDC2x1 inst_and_b89_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire89_0_3));
INVC inst_inv_b89_0_3 (.A(imd_wire89_0_3),.Y(wire89_0_3));
NANDC2x1 inst_and_b89_1_0 (.A(wire89_0_0),.B(wire89_0_1),.Y(imd_wire89_1_0));
INVC inst_inv_b89_1_0 (.A(imd_wire89_1_0),.Y(wire89_1_0));
NANDC2x1 inst_and_b89_1_1 (.A(wire89_0_2),.B(wire89_0_3),.Y(imd_wire89_1_1));
INVC inst_inv_b89_1_1 (.A(imd_wire89_1_1),.Y(wire89_1_1));
NANDC2x1 inst_and_b89_2_0 (.A(wire89_1_0),.B(wire89_1_1),.Y(imd_Y89));
INVC inst_inv_b89_2_0 (.A(imd_Y89),.Y(Y89));
NANDC2x1 inst_clockedAND_b89_89 (.A(CLK),.B(Y89),.Y(imd_YF89));
INVC inst_clockedinv_b89_89 (.A(imd_YF89),.Y(YF89));


NANDC2x1 inst_and_b90_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire90_0_0));
INVC inst_inv_b90_0_0 (.A(imd_wire90_0_0),.Y(wire90_0_0));
NANDC2x1 inst_and_b90_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire90_0_1));
INVC inst_inv_b90_0_1 (.A(imd_wire90_0_1),.Y(wire90_0_1));
NANDC2x1 inst_and_b90_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire90_0_2));
INVC inst_inv_b90_0_2 (.A(imd_wire90_0_2),.Y(wire90_0_2));
NANDC2x1 inst_and_b90_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire90_0_3));
INVC inst_inv_b90_0_3 (.A(imd_wire90_0_3),.Y(wire90_0_3));
NANDC2x1 inst_and_b90_1_0 (.A(wire90_0_0),.B(wire90_0_1),.Y(imd_wire90_1_0));
INVC inst_inv_b90_1_0 (.A(imd_wire90_1_0),.Y(wire90_1_0));
NANDC2x1 inst_and_b90_1_1 (.A(wire90_0_2),.B(wire90_0_3),.Y(imd_wire90_1_1));
INVC inst_inv_b90_1_1 (.A(imd_wire90_1_1),.Y(wire90_1_1));
NANDC2x1 inst_and_b90_2_0 (.A(wire90_1_0),.B(wire90_1_1),.Y(imd_Y90));
INVC inst_inv_b90_2_0 (.A(imd_Y90),.Y(Y90));
NANDC2x1 inst_clockedAND_b90_90 (.A(CLK),.B(Y90),.Y(imd_YF90));
INVC inst_clockedinv_b90_90 (.A(imd_YF90),.Y(YF90));


NANDC2x1 inst_and_b91_0_0 (.A(A0),.B(A1),.Y(imd_wire91_0_0));
INVC inst_inv_b91_0_0 (.A(imd_wire91_0_0),.Y(wire91_0_0));
NANDC2x1 inst_and_b91_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire91_0_1));
INVC inst_inv_b91_0_1 (.A(imd_wire91_0_1),.Y(wire91_0_1));
NANDC2x1 inst_and_b91_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire91_0_2));
INVC inst_inv_b91_0_2 (.A(imd_wire91_0_2),.Y(wire91_0_2));
NANDC2x1 inst_and_b91_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire91_0_3));
INVC inst_inv_b91_0_3 (.A(imd_wire91_0_3),.Y(wire91_0_3));
NANDC2x1 inst_and_b91_1_0 (.A(wire91_0_0),.B(wire91_0_1),.Y(imd_wire91_1_0));
INVC inst_inv_b91_1_0 (.A(imd_wire91_1_0),.Y(wire91_1_0));
NANDC2x1 inst_and_b91_1_1 (.A(wire91_0_2),.B(wire91_0_3),.Y(imd_wire91_1_1));
INVC inst_inv_b91_1_1 (.A(imd_wire91_1_1),.Y(wire91_1_1));
NANDC2x1 inst_and_b91_2_0 (.A(wire91_1_0),.B(wire91_1_1),.Y(imd_Y91));
INVC inst_inv_b91_2_0 (.A(imd_Y91),.Y(Y91));
NANDC2x1 inst_clockedAND_b91_91 (.A(CLK),.B(Y91),.Y(imd_YF91));
INVC inst_clockedinv_b91_91 (.A(imd_YF91),.Y(YF91));


NANDC2x1 inst_and_b92_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire92_0_0));
INVC inst_inv_b92_0_0 (.A(imd_wire92_0_0),.Y(wire92_0_0));
NANDC2x1 inst_and_b92_0_1 (.A(A2),.B(A3),.Y(imd_wire92_0_1));
INVC inst_inv_b92_0_1 (.A(imd_wire92_0_1),.Y(wire92_0_1));
NANDC2x1 inst_and_b92_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire92_0_2));
INVC inst_inv_b92_0_2 (.A(imd_wire92_0_2),.Y(wire92_0_2));
NANDC2x1 inst_and_b92_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire92_0_3));
INVC inst_inv_b92_0_3 (.A(imd_wire92_0_3),.Y(wire92_0_3));
NANDC2x1 inst_and_b92_1_0 (.A(wire92_0_0),.B(wire92_0_1),.Y(imd_wire92_1_0));
INVC inst_inv_b92_1_0 (.A(imd_wire92_1_0),.Y(wire92_1_0));
NANDC2x1 inst_and_b92_1_1 (.A(wire92_0_2),.B(wire92_0_3),.Y(imd_wire92_1_1));
INVC inst_inv_b92_1_1 (.A(imd_wire92_1_1),.Y(wire92_1_1));
NANDC2x1 inst_and_b92_2_0 (.A(wire92_1_0),.B(wire92_1_1),.Y(imd_Y92));
INVC inst_inv_b92_2_0 (.A(imd_Y92),.Y(Y92));
NANDC2x1 inst_clockedAND_b92_92 (.A(CLK),.B(Y92),.Y(imd_YF92));
INVC inst_clockedinv_b92_92 (.A(imd_YF92),.Y(YF92));


NANDC2x1 inst_and_b93_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire93_0_0));
INVC inst_inv_b93_0_0 (.A(imd_wire93_0_0),.Y(wire93_0_0));
NANDC2x1 inst_and_b93_0_1 (.A(A2),.B(A3),.Y(imd_wire93_0_1));
INVC inst_inv_b93_0_1 (.A(imd_wire93_0_1),.Y(wire93_0_1));
NANDC2x1 inst_and_b93_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire93_0_2));
INVC inst_inv_b93_0_2 (.A(imd_wire93_0_2),.Y(wire93_0_2));
NANDC2x1 inst_and_b93_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire93_0_3));
INVC inst_inv_b93_0_3 (.A(imd_wire93_0_3),.Y(wire93_0_3));
NANDC2x1 inst_and_b93_1_0 (.A(wire93_0_0),.B(wire93_0_1),.Y(imd_wire93_1_0));
INVC inst_inv_b93_1_0 (.A(imd_wire93_1_0),.Y(wire93_1_0));
NANDC2x1 inst_and_b93_1_1 (.A(wire93_0_2),.B(wire93_0_3),.Y(imd_wire93_1_1));
INVC inst_inv_b93_1_1 (.A(imd_wire93_1_1),.Y(wire93_1_1));
NANDC2x1 inst_and_b93_2_0 (.A(wire93_1_0),.B(wire93_1_1),.Y(imd_Y93));
INVC inst_inv_b93_2_0 (.A(imd_Y93),.Y(Y93));
NANDC2x1 inst_clockedAND_b93_93 (.A(CLK),.B(Y93),.Y(imd_YF93));
INVC inst_clockedinv_b93_93 (.A(imd_YF93),.Y(YF93));


NANDC2x1 inst_and_b94_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire94_0_0));
INVC inst_inv_b94_0_0 (.A(imd_wire94_0_0),.Y(wire94_0_0));
NANDC2x1 inst_and_b94_0_1 (.A(A2),.B(A3),.Y(imd_wire94_0_1));
INVC inst_inv_b94_0_1 (.A(imd_wire94_0_1),.Y(wire94_0_1));
NANDC2x1 inst_and_b94_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire94_0_2));
INVC inst_inv_b94_0_2 (.A(imd_wire94_0_2),.Y(wire94_0_2));
NANDC2x1 inst_and_b94_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire94_0_3));
INVC inst_inv_b94_0_3 (.A(imd_wire94_0_3),.Y(wire94_0_3));
NANDC2x1 inst_and_b94_1_0 (.A(wire94_0_0),.B(wire94_0_1),.Y(imd_wire94_1_0));
INVC inst_inv_b94_1_0 (.A(imd_wire94_1_0),.Y(wire94_1_0));
NANDC2x1 inst_and_b94_1_1 (.A(wire94_0_2),.B(wire94_0_3),.Y(imd_wire94_1_1));
INVC inst_inv_b94_1_1 (.A(imd_wire94_1_1),.Y(wire94_1_1));
NANDC2x1 inst_and_b94_2_0 (.A(wire94_1_0),.B(wire94_1_1),.Y(imd_Y94));
INVC inst_inv_b94_2_0 (.A(imd_Y94),.Y(Y94));
NANDC2x1 inst_clockedAND_b94_94 (.A(CLK),.B(Y94),.Y(imd_YF94));
INVC inst_clockedinv_b94_94 (.A(imd_YF94),.Y(YF94));


NANDC2x1 inst_and_b95_0_0 (.A(A0),.B(A1),.Y(imd_wire95_0_0));
INVC inst_inv_b95_0_0 (.A(imd_wire95_0_0),.Y(wire95_0_0));
NANDC2x1 inst_and_b95_0_1 (.A(A2),.B(A3),.Y(imd_wire95_0_1));
INVC inst_inv_b95_0_1 (.A(imd_wire95_0_1),.Y(wire95_0_1));
NANDC2x1 inst_and_b95_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire95_0_2));
INVC inst_inv_b95_0_2 (.A(imd_wire95_0_2),.Y(wire95_0_2));
NANDC2x1 inst_and_b95_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire95_0_3));
INVC inst_inv_b95_0_3 (.A(imd_wire95_0_3),.Y(wire95_0_3));
NANDC2x1 inst_and_b95_1_0 (.A(wire95_0_0),.B(wire95_0_1),.Y(imd_wire95_1_0));
INVC inst_inv_b95_1_0 (.A(imd_wire95_1_0),.Y(wire95_1_0));
NANDC2x1 inst_and_b95_1_1 (.A(wire95_0_2),.B(wire95_0_3),.Y(imd_wire95_1_1));
INVC inst_inv_b95_1_1 (.A(imd_wire95_1_1),.Y(wire95_1_1));
NANDC2x1 inst_and_b95_2_0 (.A(wire95_1_0),.B(wire95_1_1),.Y(imd_Y95));
INVC inst_inv_b95_2_0 (.A(imd_Y95),.Y(Y95));
NANDC2x1 inst_clockedAND_b95_95 (.A(CLK),.B(Y95),.Y(imd_YF95));
INVC inst_clockedinv_b95_95 (.A(imd_YF95),.Y(YF95));


NANDC2x1 inst_and_b96_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire96_0_0));
INVC inst_inv_b96_0_0 (.A(imd_wire96_0_0),.Y(wire96_0_0));
NANDC2x1 inst_and_b96_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire96_0_1));
INVC inst_inv_b96_0_1 (.A(imd_wire96_0_1),.Y(wire96_0_1));
NANDC2x1 inst_and_b96_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire96_0_2));
INVC inst_inv_b96_0_2 (.A(imd_wire96_0_2),.Y(wire96_0_2));
NANDC2x1 inst_and_b96_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire96_0_3));
INVC inst_inv_b96_0_3 (.A(imd_wire96_0_3),.Y(wire96_0_3));
NANDC2x1 inst_and_b96_1_0 (.A(wire96_0_0),.B(wire96_0_1),.Y(imd_wire96_1_0));
INVC inst_inv_b96_1_0 (.A(imd_wire96_1_0),.Y(wire96_1_0));
NANDC2x1 inst_and_b96_1_1 (.A(wire96_0_2),.B(wire96_0_3),.Y(imd_wire96_1_1));
INVC inst_inv_b96_1_1 (.A(imd_wire96_1_1),.Y(wire96_1_1));
NANDC2x1 inst_and_b96_2_0 (.A(wire96_1_0),.B(wire96_1_1),.Y(imd_Y96));
INVC inst_inv_b96_2_0 (.A(imd_Y96),.Y(Y96));
NANDC2x1 inst_clockedAND_b96_96 (.A(CLK),.B(Y96),.Y(imd_YF96));
INVC inst_clockedinv_b96_96 (.A(imd_YF96),.Y(YF96));


NANDC2x1 inst_and_b97_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire97_0_0));
INVC inst_inv_b97_0_0 (.A(imd_wire97_0_0),.Y(wire97_0_0));
NANDC2x1 inst_and_b97_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire97_0_1));
INVC inst_inv_b97_0_1 (.A(imd_wire97_0_1),.Y(wire97_0_1));
NANDC2x1 inst_and_b97_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire97_0_2));
INVC inst_inv_b97_0_2 (.A(imd_wire97_0_2),.Y(wire97_0_2));
NANDC2x1 inst_and_b97_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire97_0_3));
INVC inst_inv_b97_0_3 (.A(imd_wire97_0_3),.Y(wire97_0_3));
NANDC2x1 inst_and_b97_1_0 (.A(wire97_0_0),.B(wire97_0_1),.Y(imd_wire97_1_0));
INVC inst_inv_b97_1_0 (.A(imd_wire97_1_0),.Y(wire97_1_0));
NANDC2x1 inst_and_b97_1_1 (.A(wire97_0_2),.B(wire97_0_3),.Y(imd_wire97_1_1));
INVC inst_inv_b97_1_1 (.A(imd_wire97_1_1),.Y(wire97_1_1));
NANDC2x1 inst_and_b97_2_0 (.A(wire97_1_0),.B(wire97_1_1),.Y(imd_Y97));
INVC inst_inv_b97_2_0 (.A(imd_Y97),.Y(Y97));
NANDC2x1 inst_clockedAND_b97_97 (.A(CLK),.B(Y97),.Y(imd_YF97));
INVC inst_clockedinv_b97_97 (.A(imd_YF97),.Y(YF97));


NANDC2x1 inst_and_b98_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire98_0_0));
INVC inst_inv_b98_0_0 (.A(imd_wire98_0_0),.Y(wire98_0_0));
NANDC2x1 inst_and_b98_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire98_0_1));
INVC inst_inv_b98_0_1 (.A(imd_wire98_0_1),.Y(wire98_0_1));
NANDC2x1 inst_and_b98_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire98_0_2));
INVC inst_inv_b98_0_2 (.A(imd_wire98_0_2),.Y(wire98_0_2));
NANDC2x1 inst_and_b98_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire98_0_3));
INVC inst_inv_b98_0_3 (.A(imd_wire98_0_3),.Y(wire98_0_3));
NANDC2x1 inst_and_b98_1_0 (.A(wire98_0_0),.B(wire98_0_1),.Y(imd_wire98_1_0));
INVC inst_inv_b98_1_0 (.A(imd_wire98_1_0),.Y(wire98_1_0));
NANDC2x1 inst_and_b98_1_1 (.A(wire98_0_2),.B(wire98_0_3),.Y(imd_wire98_1_1));
INVC inst_inv_b98_1_1 (.A(imd_wire98_1_1),.Y(wire98_1_1));
NANDC2x1 inst_and_b98_2_0 (.A(wire98_1_0),.B(wire98_1_1),.Y(imd_Y98));
INVC inst_inv_b98_2_0 (.A(imd_Y98),.Y(Y98));
NANDC2x1 inst_clockedAND_b98_98 (.A(CLK),.B(Y98),.Y(imd_YF98));
INVC inst_clockedinv_b98_98 (.A(imd_YF98),.Y(YF98));


NANDC2x1 inst_and_b99_0_0 (.A(A0),.B(A1),.Y(imd_wire99_0_0));
INVC inst_inv_b99_0_0 (.A(imd_wire99_0_0),.Y(wire99_0_0));
NANDC2x1 inst_and_b99_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire99_0_1));
INVC inst_inv_b99_0_1 (.A(imd_wire99_0_1),.Y(wire99_0_1));
NANDC2x1 inst_and_b99_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire99_0_2));
INVC inst_inv_b99_0_2 (.A(imd_wire99_0_2),.Y(wire99_0_2));
NANDC2x1 inst_and_b99_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire99_0_3));
INVC inst_inv_b99_0_3 (.A(imd_wire99_0_3),.Y(wire99_0_3));
NANDC2x1 inst_and_b99_1_0 (.A(wire99_0_0),.B(wire99_0_1),.Y(imd_wire99_1_0));
INVC inst_inv_b99_1_0 (.A(imd_wire99_1_0),.Y(wire99_1_0));
NANDC2x1 inst_and_b99_1_1 (.A(wire99_0_2),.B(wire99_0_3),.Y(imd_wire99_1_1));
INVC inst_inv_b99_1_1 (.A(imd_wire99_1_1),.Y(wire99_1_1));
NANDC2x1 inst_and_b99_2_0 (.A(wire99_1_0),.B(wire99_1_1),.Y(imd_Y99));
INVC inst_inv_b99_2_0 (.A(imd_Y99),.Y(Y99));
NANDC2x1 inst_clockedAND_b99_99 (.A(CLK),.B(Y99),.Y(imd_YF99));
INVC inst_clockedinv_b99_99 (.A(imd_YF99),.Y(YF99));


NANDC2x1 inst_and_b100_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire100_0_0));
INVC inst_inv_b100_0_0 (.A(imd_wire100_0_0),.Y(wire100_0_0));
NANDC2x1 inst_and_b100_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire100_0_1));
INVC inst_inv_b100_0_1 (.A(imd_wire100_0_1),.Y(wire100_0_1));
NANDC2x1 inst_and_b100_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire100_0_2));
INVC inst_inv_b100_0_2 (.A(imd_wire100_0_2),.Y(wire100_0_2));
NANDC2x1 inst_and_b100_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire100_0_3));
INVC inst_inv_b100_0_3 (.A(imd_wire100_0_3),.Y(wire100_0_3));
NANDC2x1 inst_and_b100_1_0 (.A(wire100_0_0),.B(wire100_0_1),.Y(imd_wire100_1_0));
INVC inst_inv_b100_1_0 (.A(imd_wire100_1_0),.Y(wire100_1_0));
NANDC2x1 inst_and_b100_1_1 (.A(wire100_0_2),.B(wire100_0_3),.Y(imd_wire100_1_1));
INVC inst_inv_b100_1_1 (.A(imd_wire100_1_1),.Y(wire100_1_1));
NANDC2x1 inst_and_b100_2_0 (.A(wire100_1_0),.B(wire100_1_1),.Y(imd_Y100));
INVC inst_inv_b100_2_0 (.A(imd_Y100),.Y(Y100));
NANDC2x1 inst_clockedAND_b100_100 (.A(CLK),.B(Y100),.Y(imd_YF100));
INVC inst_clockedinv_b100_100 (.A(imd_YF100),.Y(YF100));


NANDC2x1 inst_and_b101_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire101_0_0));
INVC inst_inv_b101_0_0 (.A(imd_wire101_0_0),.Y(wire101_0_0));
NANDC2x1 inst_and_b101_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire101_0_1));
INVC inst_inv_b101_0_1 (.A(imd_wire101_0_1),.Y(wire101_0_1));
NANDC2x1 inst_and_b101_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire101_0_2));
INVC inst_inv_b101_0_2 (.A(imd_wire101_0_2),.Y(wire101_0_2));
NANDC2x1 inst_and_b101_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire101_0_3));
INVC inst_inv_b101_0_3 (.A(imd_wire101_0_3),.Y(wire101_0_3));
NANDC2x1 inst_and_b101_1_0 (.A(wire101_0_0),.B(wire101_0_1),.Y(imd_wire101_1_0));
INVC inst_inv_b101_1_0 (.A(imd_wire101_1_0),.Y(wire101_1_0));
NANDC2x1 inst_and_b101_1_1 (.A(wire101_0_2),.B(wire101_0_3),.Y(imd_wire101_1_1));
INVC inst_inv_b101_1_1 (.A(imd_wire101_1_1),.Y(wire101_1_1));
NANDC2x1 inst_and_b101_2_0 (.A(wire101_1_0),.B(wire101_1_1),.Y(imd_Y101));
INVC inst_inv_b101_2_0 (.A(imd_Y101),.Y(Y101));
NANDC2x1 inst_clockedAND_b101_101 (.A(CLK),.B(Y101),.Y(imd_YF101));
INVC inst_clockedinv_b101_101 (.A(imd_YF101),.Y(YF101));


NANDC2x1 inst_and_b102_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire102_0_0));
INVC inst_inv_b102_0_0 (.A(imd_wire102_0_0),.Y(wire102_0_0));
NANDC2x1 inst_and_b102_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire102_0_1));
INVC inst_inv_b102_0_1 (.A(imd_wire102_0_1),.Y(wire102_0_1));
NANDC2x1 inst_and_b102_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire102_0_2));
INVC inst_inv_b102_0_2 (.A(imd_wire102_0_2),.Y(wire102_0_2));
NANDC2x1 inst_and_b102_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire102_0_3));
INVC inst_inv_b102_0_3 (.A(imd_wire102_0_3),.Y(wire102_0_3));
NANDC2x1 inst_and_b102_1_0 (.A(wire102_0_0),.B(wire102_0_1),.Y(imd_wire102_1_0));
INVC inst_inv_b102_1_0 (.A(imd_wire102_1_0),.Y(wire102_1_0));
NANDC2x1 inst_and_b102_1_1 (.A(wire102_0_2),.B(wire102_0_3),.Y(imd_wire102_1_1));
INVC inst_inv_b102_1_1 (.A(imd_wire102_1_1),.Y(wire102_1_1));
NANDC2x1 inst_and_b102_2_0 (.A(wire102_1_0),.B(wire102_1_1),.Y(imd_Y102));
INVC inst_inv_b102_2_0 (.A(imd_Y102),.Y(Y102));
NANDC2x1 inst_clockedAND_b102_102 (.A(CLK),.B(Y102),.Y(imd_YF102));
INVC inst_clockedinv_b102_102 (.A(imd_YF102),.Y(YF102));


NANDC2x1 inst_and_b103_0_0 (.A(A0),.B(A1),.Y(imd_wire103_0_0));
INVC inst_inv_b103_0_0 (.A(imd_wire103_0_0),.Y(wire103_0_0));
NANDC2x1 inst_and_b103_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire103_0_1));
INVC inst_inv_b103_0_1 (.A(imd_wire103_0_1),.Y(wire103_0_1));
NANDC2x1 inst_and_b103_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire103_0_2));
INVC inst_inv_b103_0_2 (.A(imd_wire103_0_2),.Y(wire103_0_2));
NANDC2x1 inst_and_b103_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire103_0_3));
INVC inst_inv_b103_0_3 (.A(imd_wire103_0_3),.Y(wire103_0_3));
NANDC2x1 inst_and_b103_1_0 (.A(wire103_0_0),.B(wire103_0_1),.Y(imd_wire103_1_0));
INVC inst_inv_b103_1_0 (.A(imd_wire103_1_0),.Y(wire103_1_0));
NANDC2x1 inst_and_b103_1_1 (.A(wire103_0_2),.B(wire103_0_3),.Y(imd_wire103_1_1));
INVC inst_inv_b103_1_1 (.A(imd_wire103_1_1),.Y(wire103_1_1));
NANDC2x1 inst_and_b103_2_0 (.A(wire103_1_0),.B(wire103_1_1),.Y(imd_Y103));
INVC inst_inv_b103_2_0 (.A(imd_Y103),.Y(Y103));
NANDC2x1 inst_clockedAND_b103_103 (.A(CLK),.B(Y103),.Y(imd_YF103));
INVC inst_clockedinv_b103_103 (.A(imd_YF103),.Y(YF103));


NANDC2x1 inst_and_b104_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire104_0_0));
INVC inst_inv_b104_0_0 (.A(imd_wire104_0_0),.Y(wire104_0_0));
NANDC2x1 inst_and_b104_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire104_0_1));
INVC inst_inv_b104_0_1 (.A(imd_wire104_0_1),.Y(wire104_0_1));
NANDC2x1 inst_and_b104_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire104_0_2));
INVC inst_inv_b104_0_2 (.A(imd_wire104_0_2),.Y(wire104_0_2));
NANDC2x1 inst_and_b104_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire104_0_3));
INVC inst_inv_b104_0_3 (.A(imd_wire104_0_3),.Y(wire104_0_3));
NANDC2x1 inst_and_b104_1_0 (.A(wire104_0_0),.B(wire104_0_1),.Y(imd_wire104_1_0));
INVC inst_inv_b104_1_0 (.A(imd_wire104_1_0),.Y(wire104_1_0));
NANDC2x1 inst_and_b104_1_1 (.A(wire104_0_2),.B(wire104_0_3),.Y(imd_wire104_1_1));
INVC inst_inv_b104_1_1 (.A(imd_wire104_1_1),.Y(wire104_1_1));
NANDC2x1 inst_and_b104_2_0 (.A(wire104_1_0),.B(wire104_1_1),.Y(imd_Y104));
INVC inst_inv_b104_2_0 (.A(imd_Y104),.Y(Y104));
NANDC2x1 inst_clockedAND_b104_104 (.A(CLK),.B(Y104),.Y(imd_YF104));
INVC inst_clockedinv_b104_104 (.A(imd_YF104),.Y(YF104));


NANDC2x1 inst_and_b105_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire105_0_0));
INVC inst_inv_b105_0_0 (.A(imd_wire105_0_0),.Y(wire105_0_0));
NANDC2x1 inst_and_b105_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire105_0_1));
INVC inst_inv_b105_0_1 (.A(imd_wire105_0_1),.Y(wire105_0_1));
NANDC2x1 inst_and_b105_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire105_0_2));
INVC inst_inv_b105_0_2 (.A(imd_wire105_0_2),.Y(wire105_0_2));
NANDC2x1 inst_and_b105_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire105_0_3));
INVC inst_inv_b105_0_3 (.A(imd_wire105_0_3),.Y(wire105_0_3));
NANDC2x1 inst_and_b105_1_0 (.A(wire105_0_0),.B(wire105_0_1),.Y(imd_wire105_1_0));
INVC inst_inv_b105_1_0 (.A(imd_wire105_1_0),.Y(wire105_1_0));
NANDC2x1 inst_and_b105_1_1 (.A(wire105_0_2),.B(wire105_0_3),.Y(imd_wire105_1_1));
INVC inst_inv_b105_1_1 (.A(imd_wire105_1_1),.Y(wire105_1_1));
NANDC2x1 inst_and_b105_2_0 (.A(wire105_1_0),.B(wire105_1_1),.Y(imd_Y105));
INVC inst_inv_b105_2_0 (.A(imd_Y105),.Y(Y105));
NANDC2x1 inst_clockedAND_b105_105 (.A(CLK),.B(Y105),.Y(imd_YF105));
INVC inst_clockedinv_b105_105 (.A(imd_YF105),.Y(YF105));


NANDC2x1 inst_and_b106_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire106_0_0));
INVC inst_inv_b106_0_0 (.A(imd_wire106_0_0),.Y(wire106_0_0));
NANDC2x1 inst_and_b106_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire106_0_1));
INVC inst_inv_b106_0_1 (.A(imd_wire106_0_1),.Y(wire106_0_1));
NANDC2x1 inst_and_b106_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire106_0_2));
INVC inst_inv_b106_0_2 (.A(imd_wire106_0_2),.Y(wire106_0_2));
NANDC2x1 inst_and_b106_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire106_0_3));
INVC inst_inv_b106_0_3 (.A(imd_wire106_0_3),.Y(wire106_0_3));
NANDC2x1 inst_and_b106_1_0 (.A(wire106_0_0),.B(wire106_0_1),.Y(imd_wire106_1_0));
INVC inst_inv_b106_1_0 (.A(imd_wire106_1_0),.Y(wire106_1_0));
NANDC2x1 inst_and_b106_1_1 (.A(wire106_0_2),.B(wire106_0_3),.Y(imd_wire106_1_1));
INVC inst_inv_b106_1_1 (.A(imd_wire106_1_1),.Y(wire106_1_1));
NANDC2x1 inst_and_b106_2_0 (.A(wire106_1_0),.B(wire106_1_1),.Y(imd_Y106));
INVC inst_inv_b106_2_0 (.A(imd_Y106),.Y(Y106));
NANDC2x1 inst_clockedAND_b106_106 (.A(CLK),.B(Y106),.Y(imd_YF106));
INVC inst_clockedinv_b106_106 (.A(imd_YF106),.Y(YF106));


NANDC2x1 inst_and_b107_0_0 (.A(A0),.B(A1),.Y(imd_wire107_0_0));
INVC inst_inv_b107_0_0 (.A(imd_wire107_0_0),.Y(wire107_0_0));
NANDC2x1 inst_and_b107_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire107_0_1));
INVC inst_inv_b107_0_1 (.A(imd_wire107_0_1),.Y(wire107_0_1));
NANDC2x1 inst_and_b107_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire107_0_2));
INVC inst_inv_b107_0_2 (.A(imd_wire107_0_2),.Y(wire107_0_2));
NANDC2x1 inst_and_b107_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire107_0_3));
INVC inst_inv_b107_0_3 (.A(imd_wire107_0_3),.Y(wire107_0_3));
NANDC2x1 inst_and_b107_1_0 (.A(wire107_0_0),.B(wire107_0_1),.Y(imd_wire107_1_0));
INVC inst_inv_b107_1_0 (.A(imd_wire107_1_0),.Y(wire107_1_0));
NANDC2x1 inst_and_b107_1_1 (.A(wire107_0_2),.B(wire107_0_3),.Y(imd_wire107_1_1));
INVC inst_inv_b107_1_1 (.A(imd_wire107_1_1),.Y(wire107_1_1));
NANDC2x1 inst_and_b107_2_0 (.A(wire107_1_0),.B(wire107_1_1),.Y(imd_Y107));
INVC inst_inv_b107_2_0 (.A(imd_Y107),.Y(Y107));
NANDC2x1 inst_clockedAND_b107_107 (.A(CLK),.B(Y107),.Y(imd_YF107));
INVC inst_clockedinv_b107_107 (.A(imd_YF107),.Y(YF107));


NANDC2x1 inst_and_b108_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire108_0_0));
INVC inst_inv_b108_0_0 (.A(imd_wire108_0_0),.Y(wire108_0_0));
NANDC2x1 inst_and_b108_0_1 (.A(A2),.B(A3),.Y(imd_wire108_0_1));
INVC inst_inv_b108_0_1 (.A(imd_wire108_0_1),.Y(wire108_0_1));
NANDC2x1 inst_and_b108_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire108_0_2));
INVC inst_inv_b108_0_2 (.A(imd_wire108_0_2),.Y(wire108_0_2));
NANDC2x1 inst_and_b108_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire108_0_3));
INVC inst_inv_b108_0_3 (.A(imd_wire108_0_3),.Y(wire108_0_3));
NANDC2x1 inst_and_b108_1_0 (.A(wire108_0_0),.B(wire108_0_1),.Y(imd_wire108_1_0));
INVC inst_inv_b108_1_0 (.A(imd_wire108_1_0),.Y(wire108_1_0));
NANDC2x1 inst_and_b108_1_1 (.A(wire108_0_2),.B(wire108_0_3),.Y(imd_wire108_1_1));
INVC inst_inv_b108_1_1 (.A(imd_wire108_1_1),.Y(wire108_1_1));
NANDC2x1 inst_and_b108_2_0 (.A(wire108_1_0),.B(wire108_1_1),.Y(imd_Y108));
INVC inst_inv_b108_2_0 (.A(imd_Y108),.Y(Y108));
NANDC2x1 inst_clockedAND_b108_108 (.A(CLK),.B(Y108),.Y(imd_YF108));
INVC inst_clockedinv_b108_108 (.A(imd_YF108),.Y(YF108));


NANDC2x1 inst_and_b109_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire109_0_0));
INVC inst_inv_b109_0_0 (.A(imd_wire109_0_0),.Y(wire109_0_0));
NANDC2x1 inst_and_b109_0_1 (.A(A2),.B(A3),.Y(imd_wire109_0_1));
INVC inst_inv_b109_0_1 (.A(imd_wire109_0_1),.Y(wire109_0_1));
NANDC2x1 inst_and_b109_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire109_0_2));
INVC inst_inv_b109_0_2 (.A(imd_wire109_0_2),.Y(wire109_0_2));
NANDC2x1 inst_and_b109_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire109_0_3));
INVC inst_inv_b109_0_3 (.A(imd_wire109_0_3),.Y(wire109_0_3));
NANDC2x1 inst_and_b109_1_0 (.A(wire109_0_0),.B(wire109_0_1),.Y(imd_wire109_1_0));
INVC inst_inv_b109_1_0 (.A(imd_wire109_1_0),.Y(wire109_1_0));
NANDC2x1 inst_and_b109_1_1 (.A(wire109_0_2),.B(wire109_0_3),.Y(imd_wire109_1_1));
INVC inst_inv_b109_1_1 (.A(imd_wire109_1_1),.Y(wire109_1_1));
NANDC2x1 inst_and_b109_2_0 (.A(wire109_1_0),.B(wire109_1_1),.Y(imd_Y109));
INVC inst_inv_b109_2_0 (.A(imd_Y109),.Y(Y109));
NANDC2x1 inst_clockedAND_b109_109 (.A(CLK),.B(Y109),.Y(imd_YF109));
INVC inst_clockedinv_b109_109 (.A(imd_YF109),.Y(YF109));


NANDC2x1 inst_and_b110_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire110_0_0));
INVC inst_inv_b110_0_0 (.A(imd_wire110_0_0),.Y(wire110_0_0));
NANDC2x1 inst_and_b110_0_1 (.A(A2),.B(A3),.Y(imd_wire110_0_1));
INVC inst_inv_b110_0_1 (.A(imd_wire110_0_1),.Y(wire110_0_1));
NANDC2x1 inst_and_b110_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire110_0_2));
INVC inst_inv_b110_0_2 (.A(imd_wire110_0_2),.Y(wire110_0_2));
NANDC2x1 inst_and_b110_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire110_0_3));
INVC inst_inv_b110_0_3 (.A(imd_wire110_0_3),.Y(wire110_0_3));
NANDC2x1 inst_and_b110_1_0 (.A(wire110_0_0),.B(wire110_0_1),.Y(imd_wire110_1_0));
INVC inst_inv_b110_1_0 (.A(imd_wire110_1_0),.Y(wire110_1_0));
NANDC2x1 inst_and_b110_1_1 (.A(wire110_0_2),.B(wire110_0_3),.Y(imd_wire110_1_1));
INVC inst_inv_b110_1_1 (.A(imd_wire110_1_1),.Y(wire110_1_1));
NANDC2x1 inst_and_b110_2_0 (.A(wire110_1_0),.B(wire110_1_1),.Y(imd_Y110));
INVC inst_inv_b110_2_0 (.A(imd_Y110),.Y(Y110));
NANDC2x1 inst_clockedAND_b110_110 (.A(CLK),.B(Y110),.Y(imd_YF110));
INVC inst_clockedinv_b110_110 (.A(imd_YF110),.Y(YF110));


NANDC2x1 inst_and_b111_0_0 (.A(A0),.B(A1),.Y(imd_wire111_0_0));
INVC inst_inv_b111_0_0 (.A(imd_wire111_0_0),.Y(wire111_0_0));
NANDC2x1 inst_and_b111_0_1 (.A(A2),.B(A3),.Y(imd_wire111_0_1));
INVC inst_inv_b111_0_1 (.A(imd_wire111_0_1),.Y(wire111_0_1));
NANDC2x1 inst_and_b111_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire111_0_2));
INVC inst_inv_b111_0_2 (.A(imd_wire111_0_2),.Y(wire111_0_2));
NANDC2x1 inst_and_b111_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire111_0_3));
INVC inst_inv_b111_0_3 (.A(imd_wire111_0_3),.Y(wire111_0_3));
NANDC2x1 inst_and_b111_1_0 (.A(wire111_0_0),.B(wire111_0_1),.Y(imd_wire111_1_0));
INVC inst_inv_b111_1_0 (.A(imd_wire111_1_0),.Y(wire111_1_0));
NANDC2x1 inst_and_b111_1_1 (.A(wire111_0_2),.B(wire111_0_3),.Y(imd_wire111_1_1));
INVC inst_inv_b111_1_1 (.A(imd_wire111_1_1),.Y(wire111_1_1));
NANDC2x1 inst_and_b111_2_0 (.A(wire111_1_0),.B(wire111_1_1),.Y(imd_Y111));
INVC inst_inv_b111_2_0 (.A(imd_Y111),.Y(Y111));
NANDC2x1 inst_clockedAND_b111_111 (.A(CLK),.B(Y111),.Y(imd_YF111));
INVC inst_clockedinv_b111_111 (.A(imd_YF111),.Y(YF111));


NANDC2x1 inst_and_b112_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire112_0_0));
INVC inst_inv_b112_0_0 (.A(imd_wire112_0_0),.Y(wire112_0_0));
NANDC2x1 inst_and_b112_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire112_0_1));
INVC inst_inv_b112_0_1 (.A(imd_wire112_0_1),.Y(wire112_0_1));
NANDC2x1 inst_and_b112_0_2 (.A(A4),.B(A5),.Y(imd_wire112_0_2));
INVC inst_inv_b112_0_2 (.A(imd_wire112_0_2),.Y(wire112_0_2));
NANDC2x1 inst_and_b112_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire112_0_3));
INVC inst_inv_b112_0_3 (.A(imd_wire112_0_3),.Y(wire112_0_3));
NANDC2x1 inst_and_b112_1_0 (.A(wire112_0_0),.B(wire112_0_1),.Y(imd_wire112_1_0));
INVC inst_inv_b112_1_0 (.A(imd_wire112_1_0),.Y(wire112_1_0));
NANDC2x1 inst_and_b112_1_1 (.A(wire112_0_2),.B(wire112_0_3),.Y(imd_wire112_1_1));
INVC inst_inv_b112_1_1 (.A(imd_wire112_1_1),.Y(wire112_1_1));
NANDC2x1 inst_and_b112_2_0 (.A(wire112_1_0),.B(wire112_1_1),.Y(imd_Y112));
INVC inst_inv_b112_2_0 (.A(imd_Y112),.Y(Y112));
NANDC2x1 inst_clockedAND_b112_112 (.A(CLK),.B(Y112),.Y(imd_YF112));
INVC inst_clockedinv_b112_112 (.A(imd_YF112),.Y(YF112));


NANDC2x1 inst_and_b113_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire113_0_0));
INVC inst_inv_b113_0_0 (.A(imd_wire113_0_0),.Y(wire113_0_0));
NANDC2x1 inst_and_b113_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire113_0_1));
INVC inst_inv_b113_0_1 (.A(imd_wire113_0_1),.Y(wire113_0_1));
NANDC2x1 inst_and_b113_0_2 (.A(A4),.B(A5),.Y(imd_wire113_0_2));
INVC inst_inv_b113_0_2 (.A(imd_wire113_0_2),.Y(wire113_0_2));
NANDC2x1 inst_and_b113_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire113_0_3));
INVC inst_inv_b113_0_3 (.A(imd_wire113_0_3),.Y(wire113_0_3));
NANDC2x1 inst_and_b113_1_0 (.A(wire113_0_0),.B(wire113_0_1),.Y(imd_wire113_1_0));
INVC inst_inv_b113_1_0 (.A(imd_wire113_1_0),.Y(wire113_1_0));
NANDC2x1 inst_and_b113_1_1 (.A(wire113_0_2),.B(wire113_0_3),.Y(imd_wire113_1_1));
INVC inst_inv_b113_1_1 (.A(imd_wire113_1_1),.Y(wire113_1_1));
NANDC2x1 inst_and_b113_2_0 (.A(wire113_1_0),.B(wire113_1_1),.Y(imd_Y113));
INVC inst_inv_b113_2_0 (.A(imd_Y113),.Y(Y113));
NANDC2x1 inst_clockedAND_b113_113 (.A(CLK),.B(Y113),.Y(imd_YF113));
INVC inst_clockedinv_b113_113 (.A(imd_YF113),.Y(YF113));


NANDC2x1 inst_and_b114_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire114_0_0));
INVC inst_inv_b114_0_0 (.A(imd_wire114_0_0),.Y(wire114_0_0));
NANDC2x1 inst_and_b114_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire114_0_1));
INVC inst_inv_b114_0_1 (.A(imd_wire114_0_1),.Y(wire114_0_1));
NANDC2x1 inst_and_b114_0_2 (.A(A4),.B(A5),.Y(imd_wire114_0_2));
INVC inst_inv_b114_0_2 (.A(imd_wire114_0_2),.Y(wire114_0_2));
NANDC2x1 inst_and_b114_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire114_0_3));
INVC inst_inv_b114_0_3 (.A(imd_wire114_0_3),.Y(wire114_0_3));
NANDC2x1 inst_and_b114_1_0 (.A(wire114_0_0),.B(wire114_0_1),.Y(imd_wire114_1_0));
INVC inst_inv_b114_1_0 (.A(imd_wire114_1_0),.Y(wire114_1_0));
NANDC2x1 inst_and_b114_1_1 (.A(wire114_0_2),.B(wire114_0_3),.Y(imd_wire114_1_1));
INVC inst_inv_b114_1_1 (.A(imd_wire114_1_1),.Y(wire114_1_1));
NANDC2x1 inst_and_b114_2_0 (.A(wire114_1_0),.B(wire114_1_1),.Y(imd_Y114));
INVC inst_inv_b114_2_0 (.A(imd_Y114),.Y(Y114));
NANDC2x1 inst_clockedAND_b114_114 (.A(CLK),.B(Y114),.Y(imd_YF114));
INVC inst_clockedinv_b114_114 (.A(imd_YF114),.Y(YF114));


NANDC2x1 inst_and_b115_0_0 (.A(A0),.B(A1),.Y(imd_wire115_0_0));
INVC inst_inv_b115_0_0 (.A(imd_wire115_0_0),.Y(wire115_0_0));
NANDC2x1 inst_and_b115_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire115_0_1));
INVC inst_inv_b115_0_1 (.A(imd_wire115_0_1),.Y(wire115_0_1));
NANDC2x1 inst_and_b115_0_2 (.A(A4),.B(A5),.Y(imd_wire115_0_2));
INVC inst_inv_b115_0_2 (.A(imd_wire115_0_2),.Y(wire115_0_2));
NANDC2x1 inst_and_b115_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire115_0_3));
INVC inst_inv_b115_0_3 (.A(imd_wire115_0_3),.Y(wire115_0_3));
NANDC2x1 inst_and_b115_1_0 (.A(wire115_0_0),.B(wire115_0_1),.Y(imd_wire115_1_0));
INVC inst_inv_b115_1_0 (.A(imd_wire115_1_0),.Y(wire115_1_0));
NANDC2x1 inst_and_b115_1_1 (.A(wire115_0_2),.B(wire115_0_3),.Y(imd_wire115_1_1));
INVC inst_inv_b115_1_1 (.A(imd_wire115_1_1),.Y(wire115_1_1));
NANDC2x1 inst_and_b115_2_0 (.A(wire115_1_0),.B(wire115_1_1),.Y(imd_Y115));
INVC inst_inv_b115_2_0 (.A(imd_Y115),.Y(Y115));
NANDC2x1 inst_clockedAND_b115_115 (.A(CLK),.B(Y115),.Y(imd_YF115));
INVC inst_clockedinv_b115_115 (.A(imd_YF115),.Y(YF115));


NANDC2x1 inst_and_b116_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire116_0_0));
INVC inst_inv_b116_0_0 (.A(imd_wire116_0_0),.Y(wire116_0_0));
NANDC2x1 inst_and_b116_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire116_0_1));
INVC inst_inv_b116_0_1 (.A(imd_wire116_0_1),.Y(wire116_0_1));
NANDC2x1 inst_and_b116_0_2 (.A(A4),.B(A5),.Y(imd_wire116_0_2));
INVC inst_inv_b116_0_2 (.A(imd_wire116_0_2),.Y(wire116_0_2));
NANDC2x1 inst_and_b116_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire116_0_3));
INVC inst_inv_b116_0_3 (.A(imd_wire116_0_3),.Y(wire116_0_3));
NANDC2x1 inst_and_b116_1_0 (.A(wire116_0_0),.B(wire116_0_1),.Y(imd_wire116_1_0));
INVC inst_inv_b116_1_0 (.A(imd_wire116_1_0),.Y(wire116_1_0));
NANDC2x1 inst_and_b116_1_1 (.A(wire116_0_2),.B(wire116_0_3),.Y(imd_wire116_1_1));
INVC inst_inv_b116_1_1 (.A(imd_wire116_1_1),.Y(wire116_1_1));
NANDC2x1 inst_and_b116_2_0 (.A(wire116_1_0),.B(wire116_1_1),.Y(imd_Y116));
INVC inst_inv_b116_2_0 (.A(imd_Y116),.Y(Y116));
NANDC2x1 inst_clockedAND_b116_116 (.A(CLK),.B(Y116),.Y(imd_YF116));
INVC inst_clockedinv_b116_116 (.A(imd_YF116),.Y(YF116));


NANDC2x1 inst_and_b117_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire117_0_0));
INVC inst_inv_b117_0_0 (.A(imd_wire117_0_0),.Y(wire117_0_0));
NANDC2x1 inst_and_b117_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire117_0_1));
INVC inst_inv_b117_0_1 (.A(imd_wire117_0_1),.Y(wire117_0_1));
NANDC2x1 inst_and_b117_0_2 (.A(A4),.B(A5),.Y(imd_wire117_0_2));
INVC inst_inv_b117_0_2 (.A(imd_wire117_0_2),.Y(wire117_0_2));
NANDC2x1 inst_and_b117_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire117_0_3));
INVC inst_inv_b117_0_3 (.A(imd_wire117_0_3),.Y(wire117_0_3));
NANDC2x1 inst_and_b117_1_0 (.A(wire117_0_0),.B(wire117_0_1),.Y(imd_wire117_1_0));
INVC inst_inv_b117_1_0 (.A(imd_wire117_1_0),.Y(wire117_1_0));
NANDC2x1 inst_and_b117_1_1 (.A(wire117_0_2),.B(wire117_0_3),.Y(imd_wire117_1_1));
INVC inst_inv_b117_1_1 (.A(imd_wire117_1_1),.Y(wire117_1_1));
NANDC2x1 inst_and_b117_2_0 (.A(wire117_1_0),.B(wire117_1_1),.Y(imd_Y117));
INVC inst_inv_b117_2_0 (.A(imd_Y117),.Y(Y117));
NANDC2x1 inst_clockedAND_b117_117 (.A(CLK),.B(Y117),.Y(imd_YF117));
INVC inst_clockedinv_b117_117 (.A(imd_YF117),.Y(YF117));


NANDC2x1 inst_and_b118_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire118_0_0));
INVC inst_inv_b118_0_0 (.A(imd_wire118_0_0),.Y(wire118_0_0));
NANDC2x1 inst_and_b118_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire118_0_1));
INVC inst_inv_b118_0_1 (.A(imd_wire118_0_1),.Y(wire118_0_1));
NANDC2x1 inst_and_b118_0_2 (.A(A4),.B(A5),.Y(imd_wire118_0_2));
INVC inst_inv_b118_0_2 (.A(imd_wire118_0_2),.Y(wire118_0_2));
NANDC2x1 inst_and_b118_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire118_0_3));
INVC inst_inv_b118_0_3 (.A(imd_wire118_0_3),.Y(wire118_0_3));
NANDC2x1 inst_and_b118_1_0 (.A(wire118_0_0),.B(wire118_0_1),.Y(imd_wire118_1_0));
INVC inst_inv_b118_1_0 (.A(imd_wire118_1_0),.Y(wire118_1_0));
NANDC2x1 inst_and_b118_1_1 (.A(wire118_0_2),.B(wire118_0_3),.Y(imd_wire118_1_1));
INVC inst_inv_b118_1_1 (.A(imd_wire118_1_1),.Y(wire118_1_1));
NANDC2x1 inst_and_b118_2_0 (.A(wire118_1_0),.B(wire118_1_1),.Y(imd_Y118));
INVC inst_inv_b118_2_0 (.A(imd_Y118),.Y(Y118));
NANDC2x1 inst_clockedAND_b118_118 (.A(CLK),.B(Y118),.Y(imd_YF118));
INVC inst_clockedinv_b118_118 (.A(imd_YF118),.Y(YF118));


NANDC2x1 inst_and_b119_0_0 (.A(A0),.B(A1),.Y(imd_wire119_0_0));
INVC inst_inv_b119_0_0 (.A(imd_wire119_0_0),.Y(wire119_0_0));
NANDC2x1 inst_and_b119_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire119_0_1));
INVC inst_inv_b119_0_1 (.A(imd_wire119_0_1),.Y(wire119_0_1));
NANDC2x1 inst_and_b119_0_2 (.A(A4),.B(A5),.Y(imd_wire119_0_2));
INVC inst_inv_b119_0_2 (.A(imd_wire119_0_2),.Y(wire119_0_2));
NANDC2x1 inst_and_b119_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire119_0_3));
INVC inst_inv_b119_0_3 (.A(imd_wire119_0_3),.Y(wire119_0_3));
NANDC2x1 inst_and_b119_1_0 (.A(wire119_0_0),.B(wire119_0_1),.Y(imd_wire119_1_0));
INVC inst_inv_b119_1_0 (.A(imd_wire119_1_0),.Y(wire119_1_0));
NANDC2x1 inst_and_b119_1_1 (.A(wire119_0_2),.B(wire119_0_3),.Y(imd_wire119_1_1));
INVC inst_inv_b119_1_1 (.A(imd_wire119_1_1),.Y(wire119_1_1));
NANDC2x1 inst_and_b119_2_0 (.A(wire119_1_0),.B(wire119_1_1),.Y(imd_Y119));
INVC inst_inv_b119_2_0 (.A(imd_Y119),.Y(Y119));
NANDC2x1 inst_clockedAND_b119_119 (.A(CLK),.B(Y119),.Y(imd_YF119));
INVC inst_clockedinv_b119_119 (.A(imd_YF119),.Y(YF119));


NANDC2x1 inst_and_b120_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire120_0_0));
INVC inst_inv_b120_0_0 (.A(imd_wire120_0_0),.Y(wire120_0_0));
NANDC2x1 inst_and_b120_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire120_0_1));
INVC inst_inv_b120_0_1 (.A(imd_wire120_0_1),.Y(wire120_0_1));
NANDC2x1 inst_and_b120_0_2 (.A(A4),.B(A5),.Y(imd_wire120_0_2));
INVC inst_inv_b120_0_2 (.A(imd_wire120_0_2),.Y(wire120_0_2));
NANDC2x1 inst_and_b120_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire120_0_3));
INVC inst_inv_b120_0_3 (.A(imd_wire120_0_3),.Y(wire120_0_3));
NANDC2x1 inst_and_b120_1_0 (.A(wire120_0_0),.B(wire120_0_1),.Y(imd_wire120_1_0));
INVC inst_inv_b120_1_0 (.A(imd_wire120_1_0),.Y(wire120_1_0));
NANDC2x1 inst_and_b120_1_1 (.A(wire120_0_2),.B(wire120_0_3),.Y(imd_wire120_1_1));
INVC inst_inv_b120_1_1 (.A(imd_wire120_1_1),.Y(wire120_1_1));
NANDC2x1 inst_and_b120_2_0 (.A(wire120_1_0),.B(wire120_1_1),.Y(imd_Y120));
INVC inst_inv_b120_2_0 (.A(imd_Y120),.Y(Y120));
NANDC2x1 inst_clockedAND_b120_120 (.A(CLK),.B(Y120),.Y(imd_YF120));
INVC inst_clockedinv_b120_120 (.A(imd_YF120),.Y(YF120));


NANDC2x1 inst_and_b121_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire121_0_0));
INVC inst_inv_b121_0_0 (.A(imd_wire121_0_0),.Y(wire121_0_0));
NANDC2x1 inst_and_b121_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire121_0_1));
INVC inst_inv_b121_0_1 (.A(imd_wire121_0_1),.Y(wire121_0_1));
NANDC2x1 inst_and_b121_0_2 (.A(A4),.B(A5),.Y(imd_wire121_0_2));
INVC inst_inv_b121_0_2 (.A(imd_wire121_0_2),.Y(wire121_0_2));
NANDC2x1 inst_and_b121_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire121_0_3));
INVC inst_inv_b121_0_3 (.A(imd_wire121_0_3),.Y(wire121_0_3));
NANDC2x1 inst_and_b121_1_0 (.A(wire121_0_0),.B(wire121_0_1),.Y(imd_wire121_1_0));
INVC inst_inv_b121_1_0 (.A(imd_wire121_1_0),.Y(wire121_1_0));
NANDC2x1 inst_and_b121_1_1 (.A(wire121_0_2),.B(wire121_0_3),.Y(imd_wire121_1_1));
INVC inst_inv_b121_1_1 (.A(imd_wire121_1_1),.Y(wire121_1_1));
NANDC2x1 inst_and_b121_2_0 (.A(wire121_1_0),.B(wire121_1_1),.Y(imd_Y121));
INVC inst_inv_b121_2_0 (.A(imd_Y121),.Y(Y121));
NANDC2x1 inst_clockedAND_b121_121 (.A(CLK),.B(Y121),.Y(imd_YF121));
INVC inst_clockedinv_b121_121 (.A(imd_YF121),.Y(YF121));


NANDC2x1 inst_and_b122_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire122_0_0));
INVC inst_inv_b122_0_0 (.A(imd_wire122_0_0),.Y(wire122_0_0));
NANDC2x1 inst_and_b122_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire122_0_1));
INVC inst_inv_b122_0_1 (.A(imd_wire122_0_1),.Y(wire122_0_1));
NANDC2x1 inst_and_b122_0_2 (.A(A4),.B(A5),.Y(imd_wire122_0_2));
INVC inst_inv_b122_0_2 (.A(imd_wire122_0_2),.Y(wire122_0_2));
NANDC2x1 inst_and_b122_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire122_0_3));
INVC inst_inv_b122_0_3 (.A(imd_wire122_0_3),.Y(wire122_0_3));
NANDC2x1 inst_and_b122_1_0 (.A(wire122_0_0),.B(wire122_0_1),.Y(imd_wire122_1_0));
INVC inst_inv_b122_1_0 (.A(imd_wire122_1_0),.Y(wire122_1_0));
NANDC2x1 inst_and_b122_1_1 (.A(wire122_0_2),.B(wire122_0_3),.Y(imd_wire122_1_1));
INVC inst_inv_b122_1_1 (.A(imd_wire122_1_1),.Y(wire122_1_1));
NANDC2x1 inst_and_b122_2_0 (.A(wire122_1_0),.B(wire122_1_1),.Y(imd_Y122));
INVC inst_inv_b122_2_0 (.A(imd_Y122),.Y(Y122));
NANDC2x1 inst_clockedAND_b122_122 (.A(CLK),.B(Y122),.Y(imd_YF122));
INVC inst_clockedinv_b122_122 (.A(imd_YF122),.Y(YF122));


NANDC2x1 inst_and_b123_0_0 (.A(A0),.B(A1),.Y(imd_wire123_0_0));
INVC inst_inv_b123_0_0 (.A(imd_wire123_0_0),.Y(wire123_0_0));
NANDC2x1 inst_and_b123_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire123_0_1));
INVC inst_inv_b123_0_1 (.A(imd_wire123_0_1),.Y(wire123_0_1));
NANDC2x1 inst_and_b123_0_2 (.A(A4),.B(A5),.Y(imd_wire123_0_2));
INVC inst_inv_b123_0_2 (.A(imd_wire123_0_2),.Y(wire123_0_2));
NANDC2x1 inst_and_b123_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire123_0_3));
INVC inst_inv_b123_0_3 (.A(imd_wire123_0_3),.Y(wire123_0_3));
NANDC2x1 inst_and_b123_1_0 (.A(wire123_0_0),.B(wire123_0_1),.Y(imd_wire123_1_0));
INVC inst_inv_b123_1_0 (.A(imd_wire123_1_0),.Y(wire123_1_0));
NANDC2x1 inst_and_b123_1_1 (.A(wire123_0_2),.B(wire123_0_3),.Y(imd_wire123_1_1));
INVC inst_inv_b123_1_1 (.A(imd_wire123_1_1),.Y(wire123_1_1));
NANDC2x1 inst_and_b123_2_0 (.A(wire123_1_0),.B(wire123_1_1),.Y(imd_Y123));
INVC inst_inv_b123_2_0 (.A(imd_Y123),.Y(Y123));
NANDC2x1 inst_clockedAND_b123_123 (.A(CLK),.B(Y123),.Y(imd_YF123));
INVC inst_clockedinv_b123_123 (.A(imd_YF123),.Y(YF123));


NANDC2x1 inst_and_b124_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire124_0_0));
INVC inst_inv_b124_0_0 (.A(imd_wire124_0_0),.Y(wire124_0_0));
NANDC2x1 inst_and_b124_0_1 (.A(A2),.B(A3),.Y(imd_wire124_0_1));
INVC inst_inv_b124_0_1 (.A(imd_wire124_0_1),.Y(wire124_0_1));
NANDC2x1 inst_and_b124_0_2 (.A(A4),.B(A5),.Y(imd_wire124_0_2));
INVC inst_inv_b124_0_2 (.A(imd_wire124_0_2),.Y(wire124_0_2));
NANDC2x1 inst_and_b124_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire124_0_3));
INVC inst_inv_b124_0_3 (.A(imd_wire124_0_3),.Y(wire124_0_3));
NANDC2x1 inst_and_b124_1_0 (.A(wire124_0_0),.B(wire124_0_1),.Y(imd_wire124_1_0));
INVC inst_inv_b124_1_0 (.A(imd_wire124_1_0),.Y(wire124_1_0));
NANDC2x1 inst_and_b124_1_1 (.A(wire124_0_2),.B(wire124_0_3),.Y(imd_wire124_1_1));
INVC inst_inv_b124_1_1 (.A(imd_wire124_1_1),.Y(wire124_1_1));
NANDC2x1 inst_and_b124_2_0 (.A(wire124_1_0),.B(wire124_1_1),.Y(imd_Y124));
INVC inst_inv_b124_2_0 (.A(imd_Y124),.Y(Y124));
NANDC2x1 inst_clockedAND_b124_124 (.A(CLK),.B(Y124),.Y(imd_YF124));
INVC inst_clockedinv_b124_124 (.A(imd_YF124),.Y(YF124));


NANDC2x1 inst_and_b125_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire125_0_0));
INVC inst_inv_b125_0_0 (.A(imd_wire125_0_0),.Y(wire125_0_0));
NANDC2x1 inst_and_b125_0_1 (.A(A2),.B(A3),.Y(imd_wire125_0_1));
INVC inst_inv_b125_0_1 (.A(imd_wire125_0_1),.Y(wire125_0_1));
NANDC2x1 inst_and_b125_0_2 (.A(A4),.B(A5),.Y(imd_wire125_0_2));
INVC inst_inv_b125_0_2 (.A(imd_wire125_0_2),.Y(wire125_0_2));
NANDC2x1 inst_and_b125_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire125_0_3));
INVC inst_inv_b125_0_3 (.A(imd_wire125_0_3),.Y(wire125_0_3));
NANDC2x1 inst_and_b125_1_0 (.A(wire125_0_0),.B(wire125_0_1),.Y(imd_wire125_1_0));
INVC inst_inv_b125_1_0 (.A(imd_wire125_1_0),.Y(wire125_1_0));
NANDC2x1 inst_and_b125_1_1 (.A(wire125_0_2),.B(wire125_0_3),.Y(imd_wire125_1_1));
INVC inst_inv_b125_1_1 (.A(imd_wire125_1_1),.Y(wire125_1_1));
NANDC2x1 inst_and_b125_2_0 (.A(wire125_1_0),.B(wire125_1_1),.Y(imd_Y125));
INVC inst_inv_b125_2_0 (.A(imd_Y125),.Y(Y125));
NANDC2x1 inst_clockedAND_b125_125 (.A(CLK),.B(Y125),.Y(imd_YF125));
INVC inst_clockedinv_b125_125 (.A(imd_YF125),.Y(YF125));


NANDC2x1 inst_and_b126_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire126_0_0));
INVC inst_inv_b126_0_0 (.A(imd_wire126_0_0),.Y(wire126_0_0));
NANDC2x1 inst_and_b126_0_1 (.A(A2),.B(A3),.Y(imd_wire126_0_1));
INVC inst_inv_b126_0_1 (.A(imd_wire126_0_1),.Y(wire126_0_1));
NANDC2x1 inst_and_b126_0_2 (.A(A4),.B(A5),.Y(imd_wire126_0_2));
INVC inst_inv_b126_0_2 (.A(imd_wire126_0_2),.Y(wire126_0_2));
NANDC2x1 inst_and_b126_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire126_0_3));
INVC inst_inv_b126_0_3 (.A(imd_wire126_0_3),.Y(wire126_0_3));
NANDC2x1 inst_and_b126_1_0 (.A(wire126_0_0),.B(wire126_0_1),.Y(imd_wire126_1_0));
INVC inst_inv_b126_1_0 (.A(imd_wire126_1_0),.Y(wire126_1_0));
NANDC2x1 inst_and_b126_1_1 (.A(wire126_0_2),.B(wire126_0_3),.Y(imd_wire126_1_1));
INVC inst_inv_b126_1_1 (.A(imd_wire126_1_1),.Y(wire126_1_1));
NANDC2x1 inst_and_b126_2_0 (.A(wire126_1_0),.B(wire126_1_1),.Y(imd_Y126));
INVC inst_inv_b126_2_0 (.A(imd_Y126),.Y(Y126));
NANDC2x1 inst_clockedAND_b126_126 (.A(CLK),.B(Y126),.Y(imd_YF126));
INVC inst_clockedinv_b126_126 (.A(imd_YF126),.Y(YF126));


NANDC2x1 inst_and_b127_0_0 (.A(A0),.B(A1),.Y(imd_wire127_0_0));
INVC inst_inv_b127_0_0 (.A(imd_wire127_0_0),.Y(wire127_0_0));
NANDC2x1 inst_and_b127_0_1 (.A(A2),.B(A3),.Y(imd_wire127_0_1));
INVC inst_inv_b127_0_1 (.A(imd_wire127_0_1),.Y(wire127_0_1));
NANDC2x1 inst_and_b127_0_2 (.A(A4),.B(A5),.Y(imd_wire127_0_2));
INVC inst_inv_b127_0_2 (.A(imd_wire127_0_2),.Y(wire127_0_2));
NANDC2x1 inst_and_b127_0_3 (.A(A6),.B(A7_inv),.Y(imd_wire127_0_3));
INVC inst_inv_b127_0_3 (.A(imd_wire127_0_3),.Y(wire127_0_3));
NANDC2x1 inst_and_b127_1_0 (.A(wire127_0_0),.B(wire127_0_1),.Y(imd_wire127_1_0));
INVC inst_inv_b127_1_0 (.A(imd_wire127_1_0),.Y(wire127_1_0));
NANDC2x1 inst_and_b127_1_1 (.A(wire127_0_2),.B(wire127_0_3),.Y(imd_wire127_1_1));
INVC inst_inv_b127_1_1 (.A(imd_wire127_1_1),.Y(wire127_1_1));
NANDC2x1 inst_and_b127_2_0 (.A(wire127_1_0),.B(wire127_1_1),.Y(imd_Y127));
INVC inst_inv_b127_2_0 (.A(imd_Y127),.Y(Y127));
NANDC2x1 inst_clockedAND_b127_127 (.A(CLK),.B(Y127),.Y(imd_YF127));
INVC inst_clockedinv_b127_127 (.A(imd_YF127),.Y(YF127));


NANDC2x1 inst_and_b128_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire128_0_0));
INVC inst_inv_b128_0_0 (.A(imd_wire128_0_0),.Y(wire128_0_0));
NANDC2x1 inst_and_b128_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire128_0_1));
INVC inst_inv_b128_0_1 (.A(imd_wire128_0_1),.Y(wire128_0_1));
NANDC2x1 inst_and_b128_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire128_0_2));
INVC inst_inv_b128_0_2 (.A(imd_wire128_0_2),.Y(wire128_0_2));
NANDC2x1 inst_and_b128_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire128_0_3));
INVC inst_inv_b128_0_3 (.A(imd_wire128_0_3),.Y(wire128_0_3));
NANDC2x1 inst_and_b128_1_0 (.A(wire128_0_0),.B(wire128_0_1),.Y(imd_wire128_1_0));
INVC inst_inv_b128_1_0 (.A(imd_wire128_1_0),.Y(wire128_1_0));
NANDC2x1 inst_and_b128_1_1 (.A(wire128_0_2),.B(wire128_0_3),.Y(imd_wire128_1_1));
INVC inst_inv_b128_1_1 (.A(imd_wire128_1_1),.Y(wire128_1_1));
NANDC2x1 inst_and_b128_2_0 (.A(wire128_1_0),.B(wire128_1_1),.Y(imd_Y128));
INVC inst_inv_b128_2_0 (.A(imd_Y128),.Y(Y128));
NANDC2x1 inst_clockedAND_b128_128 (.A(CLK),.B(Y128),.Y(imd_YF128));
INVC inst_clockedinv_b128_128 (.A(imd_YF128),.Y(YF128));


NANDC2x1 inst_and_b129_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire129_0_0));
INVC inst_inv_b129_0_0 (.A(imd_wire129_0_0),.Y(wire129_0_0));
NANDC2x1 inst_and_b129_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire129_0_1));
INVC inst_inv_b129_0_1 (.A(imd_wire129_0_1),.Y(wire129_0_1));
NANDC2x1 inst_and_b129_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire129_0_2));
INVC inst_inv_b129_0_2 (.A(imd_wire129_0_2),.Y(wire129_0_2));
NANDC2x1 inst_and_b129_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire129_0_3));
INVC inst_inv_b129_0_3 (.A(imd_wire129_0_3),.Y(wire129_0_3));
NANDC2x1 inst_and_b129_1_0 (.A(wire129_0_0),.B(wire129_0_1),.Y(imd_wire129_1_0));
INVC inst_inv_b129_1_0 (.A(imd_wire129_1_0),.Y(wire129_1_0));
NANDC2x1 inst_and_b129_1_1 (.A(wire129_0_2),.B(wire129_0_3),.Y(imd_wire129_1_1));
INVC inst_inv_b129_1_1 (.A(imd_wire129_1_1),.Y(wire129_1_1));
NANDC2x1 inst_and_b129_2_0 (.A(wire129_1_0),.B(wire129_1_1),.Y(imd_Y129));
INVC inst_inv_b129_2_0 (.A(imd_Y129),.Y(Y129));
NANDC2x1 inst_clockedAND_b129_129 (.A(CLK),.B(Y129),.Y(imd_YF129));
INVC inst_clockedinv_b129_129 (.A(imd_YF129),.Y(YF129));


NANDC2x1 inst_and_b130_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire130_0_0));
INVC inst_inv_b130_0_0 (.A(imd_wire130_0_0),.Y(wire130_0_0));
NANDC2x1 inst_and_b130_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire130_0_1));
INVC inst_inv_b130_0_1 (.A(imd_wire130_0_1),.Y(wire130_0_1));
NANDC2x1 inst_and_b130_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire130_0_2));
INVC inst_inv_b130_0_2 (.A(imd_wire130_0_2),.Y(wire130_0_2));
NANDC2x1 inst_and_b130_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire130_0_3));
INVC inst_inv_b130_0_3 (.A(imd_wire130_0_3),.Y(wire130_0_3));
NANDC2x1 inst_and_b130_1_0 (.A(wire130_0_0),.B(wire130_0_1),.Y(imd_wire130_1_0));
INVC inst_inv_b130_1_0 (.A(imd_wire130_1_0),.Y(wire130_1_0));
NANDC2x1 inst_and_b130_1_1 (.A(wire130_0_2),.B(wire130_0_3),.Y(imd_wire130_1_1));
INVC inst_inv_b130_1_1 (.A(imd_wire130_1_1),.Y(wire130_1_1));
NANDC2x1 inst_and_b130_2_0 (.A(wire130_1_0),.B(wire130_1_1),.Y(imd_Y130));
INVC inst_inv_b130_2_0 (.A(imd_Y130),.Y(Y130));
NANDC2x1 inst_clockedAND_b130_130 (.A(CLK),.B(Y130),.Y(imd_YF130));
INVC inst_clockedinv_b130_130 (.A(imd_YF130),.Y(YF130));


NANDC2x1 inst_and_b131_0_0 (.A(A0),.B(A1),.Y(imd_wire131_0_0));
INVC inst_inv_b131_0_0 (.A(imd_wire131_0_0),.Y(wire131_0_0));
NANDC2x1 inst_and_b131_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire131_0_1));
INVC inst_inv_b131_0_1 (.A(imd_wire131_0_1),.Y(wire131_0_1));
NANDC2x1 inst_and_b131_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire131_0_2));
INVC inst_inv_b131_0_2 (.A(imd_wire131_0_2),.Y(wire131_0_2));
NANDC2x1 inst_and_b131_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire131_0_3));
INVC inst_inv_b131_0_3 (.A(imd_wire131_0_3),.Y(wire131_0_3));
NANDC2x1 inst_and_b131_1_0 (.A(wire131_0_0),.B(wire131_0_1),.Y(imd_wire131_1_0));
INVC inst_inv_b131_1_0 (.A(imd_wire131_1_0),.Y(wire131_1_0));
NANDC2x1 inst_and_b131_1_1 (.A(wire131_0_2),.B(wire131_0_3),.Y(imd_wire131_1_1));
INVC inst_inv_b131_1_1 (.A(imd_wire131_1_1),.Y(wire131_1_1));
NANDC2x1 inst_and_b131_2_0 (.A(wire131_1_0),.B(wire131_1_1),.Y(imd_Y131));
INVC inst_inv_b131_2_0 (.A(imd_Y131),.Y(Y131));
NANDC2x1 inst_clockedAND_b131_131 (.A(CLK),.B(Y131),.Y(imd_YF131));
INVC inst_clockedinv_b131_131 (.A(imd_YF131),.Y(YF131));


NANDC2x1 inst_and_b132_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire132_0_0));
INVC inst_inv_b132_0_0 (.A(imd_wire132_0_0),.Y(wire132_0_0));
NANDC2x1 inst_and_b132_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire132_0_1));
INVC inst_inv_b132_0_1 (.A(imd_wire132_0_1),.Y(wire132_0_1));
NANDC2x1 inst_and_b132_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire132_0_2));
INVC inst_inv_b132_0_2 (.A(imd_wire132_0_2),.Y(wire132_0_2));
NANDC2x1 inst_and_b132_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire132_0_3));
INVC inst_inv_b132_0_3 (.A(imd_wire132_0_3),.Y(wire132_0_3));
NANDC2x1 inst_and_b132_1_0 (.A(wire132_0_0),.B(wire132_0_1),.Y(imd_wire132_1_0));
INVC inst_inv_b132_1_0 (.A(imd_wire132_1_0),.Y(wire132_1_0));
NANDC2x1 inst_and_b132_1_1 (.A(wire132_0_2),.B(wire132_0_3),.Y(imd_wire132_1_1));
INVC inst_inv_b132_1_1 (.A(imd_wire132_1_1),.Y(wire132_1_1));
NANDC2x1 inst_and_b132_2_0 (.A(wire132_1_0),.B(wire132_1_1),.Y(imd_Y132));
INVC inst_inv_b132_2_0 (.A(imd_Y132),.Y(Y132));
NANDC2x1 inst_clockedAND_b132_132 (.A(CLK),.B(Y132),.Y(imd_YF132));
INVC inst_clockedinv_b132_132 (.A(imd_YF132),.Y(YF132));


NANDC2x1 inst_and_b133_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire133_0_0));
INVC inst_inv_b133_0_0 (.A(imd_wire133_0_0),.Y(wire133_0_0));
NANDC2x1 inst_and_b133_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire133_0_1));
INVC inst_inv_b133_0_1 (.A(imd_wire133_0_1),.Y(wire133_0_1));
NANDC2x1 inst_and_b133_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire133_0_2));
INVC inst_inv_b133_0_2 (.A(imd_wire133_0_2),.Y(wire133_0_2));
NANDC2x1 inst_and_b133_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire133_0_3));
INVC inst_inv_b133_0_3 (.A(imd_wire133_0_3),.Y(wire133_0_3));
NANDC2x1 inst_and_b133_1_0 (.A(wire133_0_0),.B(wire133_0_1),.Y(imd_wire133_1_0));
INVC inst_inv_b133_1_0 (.A(imd_wire133_1_0),.Y(wire133_1_0));
NANDC2x1 inst_and_b133_1_1 (.A(wire133_0_2),.B(wire133_0_3),.Y(imd_wire133_1_1));
INVC inst_inv_b133_1_1 (.A(imd_wire133_1_1),.Y(wire133_1_1));
NANDC2x1 inst_and_b133_2_0 (.A(wire133_1_0),.B(wire133_1_1),.Y(imd_Y133));
INVC inst_inv_b133_2_0 (.A(imd_Y133),.Y(Y133));
NANDC2x1 inst_clockedAND_b133_133 (.A(CLK),.B(Y133),.Y(imd_YF133));
INVC inst_clockedinv_b133_133 (.A(imd_YF133),.Y(YF133));


NANDC2x1 inst_and_b134_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire134_0_0));
INVC inst_inv_b134_0_0 (.A(imd_wire134_0_0),.Y(wire134_0_0));
NANDC2x1 inst_and_b134_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire134_0_1));
INVC inst_inv_b134_0_1 (.A(imd_wire134_0_1),.Y(wire134_0_1));
NANDC2x1 inst_and_b134_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire134_0_2));
INVC inst_inv_b134_0_2 (.A(imd_wire134_0_2),.Y(wire134_0_2));
NANDC2x1 inst_and_b134_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire134_0_3));
INVC inst_inv_b134_0_3 (.A(imd_wire134_0_3),.Y(wire134_0_3));
NANDC2x1 inst_and_b134_1_0 (.A(wire134_0_0),.B(wire134_0_1),.Y(imd_wire134_1_0));
INVC inst_inv_b134_1_0 (.A(imd_wire134_1_0),.Y(wire134_1_0));
NANDC2x1 inst_and_b134_1_1 (.A(wire134_0_2),.B(wire134_0_3),.Y(imd_wire134_1_1));
INVC inst_inv_b134_1_1 (.A(imd_wire134_1_1),.Y(wire134_1_1));
NANDC2x1 inst_and_b134_2_0 (.A(wire134_1_0),.B(wire134_1_1),.Y(imd_Y134));
INVC inst_inv_b134_2_0 (.A(imd_Y134),.Y(Y134));
NANDC2x1 inst_clockedAND_b134_134 (.A(CLK),.B(Y134),.Y(imd_YF134));
INVC inst_clockedinv_b134_134 (.A(imd_YF134),.Y(YF134));


NANDC2x1 inst_and_b135_0_0 (.A(A0),.B(A1),.Y(imd_wire135_0_0));
INVC inst_inv_b135_0_0 (.A(imd_wire135_0_0),.Y(wire135_0_0));
NANDC2x1 inst_and_b135_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire135_0_1));
INVC inst_inv_b135_0_1 (.A(imd_wire135_0_1),.Y(wire135_0_1));
NANDC2x1 inst_and_b135_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire135_0_2));
INVC inst_inv_b135_0_2 (.A(imd_wire135_0_2),.Y(wire135_0_2));
NANDC2x1 inst_and_b135_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire135_0_3));
INVC inst_inv_b135_0_3 (.A(imd_wire135_0_3),.Y(wire135_0_3));
NANDC2x1 inst_and_b135_1_0 (.A(wire135_0_0),.B(wire135_0_1),.Y(imd_wire135_1_0));
INVC inst_inv_b135_1_0 (.A(imd_wire135_1_0),.Y(wire135_1_0));
NANDC2x1 inst_and_b135_1_1 (.A(wire135_0_2),.B(wire135_0_3),.Y(imd_wire135_1_1));
INVC inst_inv_b135_1_1 (.A(imd_wire135_1_1),.Y(wire135_1_1));
NANDC2x1 inst_and_b135_2_0 (.A(wire135_1_0),.B(wire135_1_1),.Y(imd_Y135));
INVC inst_inv_b135_2_0 (.A(imd_Y135),.Y(Y135));
NANDC2x1 inst_clockedAND_b135_135 (.A(CLK),.B(Y135),.Y(imd_YF135));
INVC inst_clockedinv_b135_135 (.A(imd_YF135),.Y(YF135));


NANDC2x1 inst_and_b136_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire136_0_0));
INVC inst_inv_b136_0_0 (.A(imd_wire136_0_0),.Y(wire136_0_0));
NANDC2x1 inst_and_b136_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire136_0_1));
INVC inst_inv_b136_0_1 (.A(imd_wire136_0_1),.Y(wire136_0_1));
NANDC2x1 inst_and_b136_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire136_0_2));
INVC inst_inv_b136_0_2 (.A(imd_wire136_0_2),.Y(wire136_0_2));
NANDC2x1 inst_and_b136_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire136_0_3));
INVC inst_inv_b136_0_3 (.A(imd_wire136_0_3),.Y(wire136_0_3));
NANDC2x1 inst_and_b136_1_0 (.A(wire136_0_0),.B(wire136_0_1),.Y(imd_wire136_1_0));
INVC inst_inv_b136_1_0 (.A(imd_wire136_1_0),.Y(wire136_1_0));
NANDC2x1 inst_and_b136_1_1 (.A(wire136_0_2),.B(wire136_0_3),.Y(imd_wire136_1_1));
INVC inst_inv_b136_1_1 (.A(imd_wire136_1_1),.Y(wire136_1_1));
NANDC2x1 inst_and_b136_2_0 (.A(wire136_1_0),.B(wire136_1_1),.Y(imd_Y136));
INVC inst_inv_b136_2_0 (.A(imd_Y136),.Y(Y136));
NANDC2x1 inst_clockedAND_b136_136 (.A(CLK),.B(Y136),.Y(imd_YF136));
INVC inst_clockedinv_b136_136 (.A(imd_YF136),.Y(YF136));


NANDC2x1 inst_and_b137_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire137_0_0));
INVC inst_inv_b137_0_0 (.A(imd_wire137_0_0),.Y(wire137_0_0));
NANDC2x1 inst_and_b137_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire137_0_1));
INVC inst_inv_b137_0_1 (.A(imd_wire137_0_1),.Y(wire137_0_1));
NANDC2x1 inst_and_b137_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire137_0_2));
INVC inst_inv_b137_0_2 (.A(imd_wire137_0_2),.Y(wire137_0_2));
NANDC2x1 inst_and_b137_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire137_0_3));
INVC inst_inv_b137_0_3 (.A(imd_wire137_0_3),.Y(wire137_0_3));
NANDC2x1 inst_and_b137_1_0 (.A(wire137_0_0),.B(wire137_0_1),.Y(imd_wire137_1_0));
INVC inst_inv_b137_1_0 (.A(imd_wire137_1_0),.Y(wire137_1_0));
NANDC2x1 inst_and_b137_1_1 (.A(wire137_0_2),.B(wire137_0_3),.Y(imd_wire137_1_1));
INVC inst_inv_b137_1_1 (.A(imd_wire137_1_1),.Y(wire137_1_1));
NANDC2x1 inst_and_b137_2_0 (.A(wire137_1_0),.B(wire137_1_1),.Y(imd_Y137));
INVC inst_inv_b137_2_0 (.A(imd_Y137),.Y(Y137));
NANDC2x1 inst_clockedAND_b137_137 (.A(CLK),.B(Y137),.Y(imd_YF137));
INVC inst_clockedinv_b137_137 (.A(imd_YF137),.Y(YF137));


NANDC2x1 inst_and_b138_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire138_0_0));
INVC inst_inv_b138_0_0 (.A(imd_wire138_0_0),.Y(wire138_0_0));
NANDC2x1 inst_and_b138_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire138_0_1));
INVC inst_inv_b138_0_1 (.A(imd_wire138_0_1),.Y(wire138_0_1));
NANDC2x1 inst_and_b138_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire138_0_2));
INVC inst_inv_b138_0_2 (.A(imd_wire138_0_2),.Y(wire138_0_2));
NANDC2x1 inst_and_b138_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire138_0_3));
INVC inst_inv_b138_0_3 (.A(imd_wire138_0_3),.Y(wire138_0_3));
NANDC2x1 inst_and_b138_1_0 (.A(wire138_0_0),.B(wire138_0_1),.Y(imd_wire138_1_0));
INVC inst_inv_b138_1_0 (.A(imd_wire138_1_0),.Y(wire138_1_0));
NANDC2x1 inst_and_b138_1_1 (.A(wire138_0_2),.B(wire138_0_3),.Y(imd_wire138_1_1));
INVC inst_inv_b138_1_1 (.A(imd_wire138_1_1),.Y(wire138_1_1));
NANDC2x1 inst_and_b138_2_0 (.A(wire138_1_0),.B(wire138_1_1),.Y(imd_Y138));
INVC inst_inv_b138_2_0 (.A(imd_Y138),.Y(Y138));
NANDC2x1 inst_clockedAND_b138_138 (.A(CLK),.B(Y138),.Y(imd_YF138));
INVC inst_clockedinv_b138_138 (.A(imd_YF138),.Y(YF138));


NANDC2x1 inst_and_b139_0_0 (.A(A0),.B(A1),.Y(imd_wire139_0_0));
INVC inst_inv_b139_0_0 (.A(imd_wire139_0_0),.Y(wire139_0_0));
NANDC2x1 inst_and_b139_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire139_0_1));
INVC inst_inv_b139_0_1 (.A(imd_wire139_0_1),.Y(wire139_0_1));
NANDC2x1 inst_and_b139_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire139_0_2));
INVC inst_inv_b139_0_2 (.A(imd_wire139_0_2),.Y(wire139_0_2));
NANDC2x1 inst_and_b139_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire139_0_3));
INVC inst_inv_b139_0_3 (.A(imd_wire139_0_3),.Y(wire139_0_3));
NANDC2x1 inst_and_b139_1_0 (.A(wire139_0_0),.B(wire139_0_1),.Y(imd_wire139_1_0));
INVC inst_inv_b139_1_0 (.A(imd_wire139_1_0),.Y(wire139_1_0));
NANDC2x1 inst_and_b139_1_1 (.A(wire139_0_2),.B(wire139_0_3),.Y(imd_wire139_1_1));
INVC inst_inv_b139_1_1 (.A(imd_wire139_1_1),.Y(wire139_1_1));
NANDC2x1 inst_and_b139_2_0 (.A(wire139_1_0),.B(wire139_1_1),.Y(imd_Y139));
INVC inst_inv_b139_2_0 (.A(imd_Y139),.Y(Y139));
NANDC2x1 inst_clockedAND_b139_139 (.A(CLK),.B(Y139),.Y(imd_YF139));
INVC inst_clockedinv_b139_139 (.A(imd_YF139),.Y(YF139));


NANDC2x1 inst_and_b140_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire140_0_0));
INVC inst_inv_b140_0_0 (.A(imd_wire140_0_0),.Y(wire140_0_0));
NANDC2x1 inst_and_b140_0_1 (.A(A2),.B(A3),.Y(imd_wire140_0_1));
INVC inst_inv_b140_0_1 (.A(imd_wire140_0_1),.Y(wire140_0_1));
NANDC2x1 inst_and_b140_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire140_0_2));
INVC inst_inv_b140_0_2 (.A(imd_wire140_0_2),.Y(wire140_0_2));
NANDC2x1 inst_and_b140_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire140_0_3));
INVC inst_inv_b140_0_3 (.A(imd_wire140_0_3),.Y(wire140_0_3));
NANDC2x1 inst_and_b140_1_0 (.A(wire140_0_0),.B(wire140_0_1),.Y(imd_wire140_1_0));
INVC inst_inv_b140_1_0 (.A(imd_wire140_1_0),.Y(wire140_1_0));
NANDC2x1 inst_and_b140_1_1 (.A(wire140_0_2),.B(wire140_0_3),.Y(imd_wire140_1_1));
INVC inst_inv_b140_1_1 (.A(imd_wire140_1_1),.Y(wire140_1_1));
NANDC2x1 inst_and_b140_2_0 (.A(wire140_1_0),.B(wire140_1_1),.Y(imd_Y140));
INVC inst_inv_b140_2_0 (.A(imd_Y140),.Y(Y140));
NANDC2x1 inst_clockedAND_b140_140 (.A(CLK),.B(Y140),.Y(imd_YF140));
INVC inst_clockedinv_b140_140 (.A(imd_YF140),.Y(YF140));


NANDC2x1 inst_and_b141_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire141_0_0));
INVC inst_inv_b141_0_0 (.A(imd_wire141_0_0),.Y(wire141_0_0));
NANDC2x1 inst_and_b141_0_1 (.A(A2),.B(A3),.Y(imd_wire141_0_1));
INVC inst_inv_b141_0_1 (.A(imd_wire141_0_1),.Y(wire141_0_1));
NANDC2x1 inst_and_b141_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire141_0_2));
INVC inst_inv_b141_0_2 (.A(imd_wire141_0_2),.Y(wire141_0_2));
NANDC2x1 inst_and_b141_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire141_0_3));
INVC inst_inv_b141_0_3 (.A(imd_wire141_0_3),.Y(wire141_0_3));
NANDC2x1 inst_and_b141_1_0 (.A(wire141_0_0),.B(wire141_0_1),.Y(imd_wire141_1_0));
INVC inst_inv_b141_1_0 (.A(imd_wire141_1_0),.Y(wire141_1_0));
NANDC2x1 inst_and_b141_1_1 (.A(wire141_0_2),.B(wire141_0_3),.Y(imd_wire141_1_1));
INVC inst_inv_b141_1_1 (.A(imd_wire141_1_1),.Y(wire141_1_1));
NANDC2x1 inst_and_b141_2_0 (.A(wire141_1_0),.B(wire141_1_1),.Y(imd_Y141));
INVC inst_inv_b141_2_0 (.A(imd_Y141),.Y(Y141));
NANDC2x1 inst_clockedAND_b141_141 (.A(CLK),.B(Y141),.Y(imd_YF141));
INVC inst_clockedinv_b141_141 (.A(imd_YF141),.Y(YF141));


NANDC2x1 inst_and_b142_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire142_0_0));
INVC inst_inv_b142_0_0 (.A(imd_wire142_0_0),.Y(wire142_0_0));
NANDC2x1 inst_and_b142_0_1 (.A(A2),.B(A3),.Y(imd_wire142_0_1));
INVC inst_inv_b142_0_1 (.A(imd_wire142_0_1),.Y(wire142_0_1));
NANDC2x1 inst_and_b142_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire142_0_2));
INVC inst_inv_b142_0_2 (.A(imd_wire142_0_2),.Y(wire142_0_2));
NANDC2x1 inst_and_b142_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire142_0_3));
INVC inst_inv_b142_0_3 (.A(imd_wire142_0_3),.Y(wire142_0_3));
NANDC2x1 inst_and_b142_1_0 (.A(wire142_0_0),.B(wire142_0_1),.Y(imd_wire142_1_0));
INVC inst_inv_b142_1_0 (.A(imd_wire142_1_0),.Y(wire142_1_0));
NANDC2x1 inst_and_b142_1_1 (.A(wire142_0_2),.B(wire142_0_3),.Y(imd_wire142_1_1));
INVC inst_inv_b142_1_1 (.A(imd_wire142_1_1),.Y(wire142_1_1));
NANDC2x1 inst_and_b142_2_0 (.A(wire142_1_0),.B(wire142_1_1),.Y(imd_Y142));
INVC inst_inv_b142_2_0 (.A(imd_Y142),.Y(Y142));
NANDC2x1 inst_clockedAND_b142_142 (.A(CLK),.B(Y142),.Y(imd_YF142));
INVC inst_clockedinv_b142_142 (.A(imd_YF142),.Y(YF142));


NANDC2x1 inst_and_b143_0_0 (.A(A0),.B(A1),.Y(imd_wire143_0_0));
INVC inst_inv_b143_0_0 (.A(imd_wire143_0_0),.Y(wire143_0_0));
NANDC2x1 inst_and_b143_0_1 (.A(A2),.B(A3),.Y(imd_wire143_0_1));
INVC inst_inv_b143_0_1 (.A(imd_wire143_0_1),.Y(wire143_0_1));
NANDC2x1 inst_and_b143_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire143_0_2));
INVC inst_inv_b143_0_2 (.A(imd_wire143_0_2),.Y(wire143_0_2));
NANDC2x1 inst_and_b143_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire143_0_3));
INVC inst_inv_b143_0_3 (.A(imd_wire143_0_3),.Y(wire143_0_3));
NANDC2x1 inst_and_b143_1_0 (.A(wire143_0_0),.B(wire143_0_1),.Y(imd_wire143_1_0));
INVC inst_inv_b143_1_0 (.A(imd_wire143_1_0),.Y(wire143_1_0));
NANDC2x1 inst_and_b143_1_1 (.A(wire143_0_2),.B(wire143_0_3),.Y(imd_wire143_1_1));
INVC inst_inv_b143_1_1 (.A(imd_wire143_1_1),.Y(wire143_1_1));
NANDC2x1 inst_and_b143_2_0 (.A(wire143_1_0),.B(wire143_1_1),.Y(imd_Y143));
INVC inst_inv_b143_2_0 (.A(imd_Y143),.Y(Y143));
NANDC2x1 inst_clockedAND_b143_143 (.A(CLK),.B(Y143),.Y(imd_YF143));
INVC inst_clockedinv_b143_143 (.A(imd_YF143),.Y(YF143));


NANDC2x1 inst_and_b144_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire144_0_0));
INVC inst_inv_b144_0_0 (.A(imd_wire144_0_0),.Y(wire144_0_0));
NANDC2x1 inst_and_b144_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire144_0_1));
INVC inst_inv_b144_0_1 (.A(imd_wire144_0_1),.Y(wire144_0_1));
NANDC2x1 inst_and_b144_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire144_0_2));
INVC inst_inv_b144_0_2 (.A(imd_wire144_0_2),.Y(wire144_0_2));
NANDC2x1 inst_and_b144_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire144_0_3));
INVC inst_inv_b144_0_3 (.A(imd_wire144_0_3),.Y(wire144_0_3));
NANDC2x1 inst_and_b144_1_0 (.A(wire144_0_0),.B(wire144_0_1),.Y(imd_wire144_1_0));
INVC inst_inv_b144_1_0 (.A(imd_wire144_1_0),.Y(wire144_1_0));
NANDC2x1 inst_and_b144_1_1 (.A(wire144_0_2),.B(wire144_0_3),.Y(imd_wire144_1_1));
INVC inst_inv_b144_1_1 (.A(imd_wire144_1_1),.Y(wire144_1_1));
NANDC2x1 inst_and_b144_2_0 (.A(wire144_1_0),.B(wire144_1_1),.Y(imd_Y144));
INVC inst_inv_b144_2_0 (.A(imd_Y144),.Y(Y144));
NANDC2x1 inst_clockedAND_b144_144 (.A(CLK),.B(Y144),.Y(imd_YF144));
INVC inst_clockedinv_b144_144 (.A(imd_YF144),.Y(YF144));


NANDC2x1 inst_and_b145_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire145_0_0));
INVC inst_inv_b145_0_0 (.A(imd_wire145_0_0),.Y(wire145_0_0));
NANDC2x1 inst_and_b145_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire145_0_1));
INVC inst_inv_b145_0_1 (.A(imd_wire145_0_1),.Y(wire145_0_1));
NANDC2x1 inst_and_b145_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire145_0_2));
INVC inst_inv_b145_0_2 (.A(imd_wire145_0_2),.Y(wire145_0_2));
NANDC2x1 inst_and_b145_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire145_0_3));
INVC inst_inv_b145_0_3 (.A(imd_wire145_0_3),.Y(wire145_0_3));
NANDC2x1 inst_and_b145_1_0 (.A(wire145_0_0),.B(wire145_0_1),.Y(imd_wire145_1_0));
INVC inst_inv_b145_1_0 (.A(imd_wire145_1_0),.Y(wire145_1_0));
NANDC2x1 inst_and_b145_1_1 (.A(wire145_0_2),.B(wire145_0_3),.Y(imd_wire145_1_1));
INVC inst_inv_b145_1_1 (.A(imd_wire145_1_1),.Y(wire145_1_1));
NANDC2x1 inst_and_b145_2_0 (.A(wire145_1_0),.B(wire145_1_1),.Y(imd_Y145));
INVC inst_inv_b145_2_0 (.A(imd_Y145),.Y(Y145));
NANDC2x1 inst_clockedAND_b145_145 (.A(CLK),.B(Y145),.Y(imd_YF145));
INVC inst_clockedinv_b145_145 (.A(imd_YF145),.Y(YF145));


NANDC2x1 inst_and_b146_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire146_0_0));
INVC inst_inv_b146_0_0 (.A(imd_wire146_0_0),.Y(wire146_0_0));
NANDC2x1 inst_and_b146_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire146_0_1));
INVC inst_inv_b146_0_1 (.A(imd_wire146_0_1),.Y(wire146_0_1));
NANDC2x1 inst_and_b146_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire146_0_2));
INVC inst_inv_b146_0_2 (.A(imd_wire146_0_2),.Y(wire146_0_2));
NANDC2x1 inst_and_b146_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire146_0_3));
INVC inst_inv_b146_0_3 (.A(imd_wire146_0_3),.Y(wire146_0_3));
NANDC2x1 inst_and_b146_1_0 (.A(wire146_0_0),.B(wire146_0_1),.Y(imd_wire146_1_0));
INVC inst_inv_b146_1_0 (.A(imd_wire146_1_0),.Y(wire146_1_0));
NANDC2x1 inst_and_b146_1_1 (.A(wire146_0_2),.B(wire146_0_3),.Y(imd_wire146_1_1));
INVC inst_inv_b146_1_1 (.A(imd_wire146_1_1),.Y(wire146_1_1));
NANDC2x1 inst_and_b146_2_0 (.A(wire146_1_0),.B(wire146_1_1),.Y(imd_Y146));
INVC inst_inv_b146_2_0 (.A(imd_Y146),.Y(Y146));
NANDC2x1 inst_clockedAND_b146_146 (.A(CLK),.B(Y146),.Y(imd_YF146));
INVC inst_clockedinv_b146_146 (.A(imd_YF146),.Y(YF146));


NANDC2x1 inst_and_b147_0_0 (.A(A0),.B(A1),.Y(imd_wire147_0_0));
INVC inst_inv_b147_0_0 (.A(imd_wire147_0_0),.Y(wire147_0_0));
NANDC2x1 inst_and_b147_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire147_0_1));
INVC inst_inv_b147_0_1 (.A(imd_wire147_0_1),.Y(wire147_0_1));
NANDC2x1 inst_and_b147_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire147_0_2));
INVC inst_inv_b147_0_2 (.A(imd_wire147_0_2),.Y(wire147_0_2));
NANDC2x1 inst_and_b147_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire147_0_3));
INVC inst_inv_b147_0_3 (.A(imd_wire147_0_3),.Y(wire147_0_3));
NANDC2x1 inst_and_b147_1_0 (.A(wire147_0_0),.B(wire147_0_1),.Y(imd_wire147_1_0));
INVC inst_inv_b147_1_0 (.A(imd_wire147_1_0),.Y(wire147_1_0));
NANDC2x1 inst_and_b147_1_1 (.A(wire147_0_2),.B(wire147_0_3),.Y(imd_wire147_1_1));
INVC inst_inv_b147_1_1 (.A(imd_wire147_1_1),.Y(wire147_1_1));
NANDC2x1 inst_and_b147_2_0 (.A(wire147_1_0),.B(wire147_1_1),.Y(imd_Y147));
INVC inst_inv_b147_2_0 (.A(imd_Y147),.Y(Y147));
NANDC2x1 inst_clockedAND_b147_147 (.A(CLK),.B(Y147),.Y(imd_YF147));
INVC inst_clockedinv_b147_147 (.A(imd_YF147),.Y(YF147));


NANDC2x1 inst_and_b148_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire148_0_0));
INVC inst_inv_b148_0_0 (.A(imd_wire148_0_0),.Y(wire148_0_0));
NANDC2x1 inst_and_b148_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire148_0_1));
INVC inst_inv_b148_0_1 (.A(imd_wire148_0_1),.Y(wire148_0_1));
NANDC2x1 inst_and_b148_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire148_0_2));
INVC inst_inv_b148_0_2 (.A(imd_wire148_0_2),.Y(wire148_0_2));
NANDC2x1 inst_and_b148_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire148_0_3));
INVC inst_inv_b148_0_3 (.A(imd_wire148_0_3),.Y(wire148_0_3));
NANDC2x1 inst_and_b148_1_0 (.A(wire148_0_0),.B(wire148_0_1),.Y(imd_wire148_1_0));
INVC inst_inv_b148_1_0 (.A(imd_wire148_1_0),.Y(wire148_1_0));
NANDC2x1 inst_and_b148_1_1 (.A(wire148_0_2),.B(wire148_0_3),.Y(imd_wire148_1_1));
INVC inst_inv_b148_1_1 (.A(imd_wire148_1_1),.Y(wire148_1_1));
NANDC2x1 inst_and_b148_2_0 (.A(wire148_1_0),.B(wire148_1_1),.Y(imd_Y148));
INVC inst_inv_b148_2_0 (.A(imd_Y148),.Y(Y148));
NANDC2x1 inst_clockedAND_b148_148 (.A(CLK),.B(Y148),.Y(imd_YF148));
INVC inst_clockedinv_b148_148 (.A(imd_YF148),.Y(YF148));


NANDC2x1 inst_and_b149_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire149_0_0));
INVC inst_inv_b149_0_0 (.A(imd_wire149_0_0),.Y(wire149_0_0));
NANDC2x1 inst_and_b149_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire149_0_1));
INVC inst_inv_b149_0_1 (.A(imd_wire149_0_1),.Y(wire149_0_1));
NANDC2x1 inst_and_b149_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire149_0_2));
INVC inst_inv_b149_0_2 (.A(imd_wire149_0_2),.Y(wire149_0_2));
NANDC2x1 inst_and_b149_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire149_0_3));
INVC inst_inv_b149_0_3 (.A(imd_wire149_0_3),.Y(wire149_0_3));
NANDC2x1 inst_and_b149_1_0 (.A(wire149_0_0),.B(wire149_0_1),.Y(imd_wire149_1_0));
INVC inst_inv_b149_1_0 (.A(imd_wire149_1_0),.Y(wire149_1_0));
NANDC2x1 inst_and_b149_1_1 (.A(wire149_0_2),.B(wire149_0_3),.Y(imd_wire149_1_1));
INVC inst_inv_b149_1_1 (.A(imd_wire149_1_1),.Y(wire149_1_1));
NANDC2x1 inst_and_b149_2_0 (.A(wire149_1_0),.B(wire149_1_1),.Y(imd_Y149));
INVC inst_inv_b149_2_0 (.A(imd_Y149),.Y(Y149));
NANDC2x1 inst_clockedAND_b149_149 (.A(CLK),.B(Y149),.Y(imd_YF149));
INVC inst_clockedinv_b149_149 (.A(imd_YF149),.Y(YF149));


NANDC2x1 inst_and_b150_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire150_0_0));
INVC inst_inv_b150_0_0 (.A(imd_wire150_0_0),.Y(wire150_0_0));
NANDC2x1 inst_and_b150_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire150_0_1));
INVC inst_inv_b150_0_1 (.A(imd_wire150_0_1),.Y(wire150_0_1));
NANDC2x1 inst_and_b150_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire150_0_2));
INVC inst_inv_b150_0_2 (.A(imd_wire150_0_2),.Y(wire150_0_2));
NANDC2x1 inst_and_b150_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire150_0_3));
INVC inst_inv_b150_0_3 (.A(imd_wire150_0_3),.Y(wire150_0_3));
NANDC2x1 inst_and_b150_1_0 (.A(wire150_0_0),.B(wire150_0_1),.Y(imd_wire150_1_0));
INVC inst_inv_b150_1_0 (.A(imd_wire150_1_0),.Y(wire150_1_0));
NANDC2x1 inst_and_b150_1_1 (.A(wire150_0_2),.B(wire150_0_3),.Y(imd_wire150_1_1));
INVC inst_inv_b150_1_1 (.A(imd_wire150_1_1),.Y(wire150_1_1));
NANDC2x1 inst_and_b150_2_0 (.A(wire150_1_0),.B(wire150_1_1),.Y(imd_Y150));
INVC inst_inv_b150_2_0 (.A(imd_Y150),.Y(Y150));
NANDC2x1 inst_clockedAND_b150_150 (.A(CLK),.B(Y150),.Y(imd_YF150));
INVC inst_clockedinv_b150_150 (.A(imd_YF150),.Y(YF150));


NANDC2x1 inst_and_b151_0_0 (.A(A0),.B(A1),.Y(imd_wire151_0_0));
INVC inst_inv_b151_0_0 (.A(imd_wire151_0_0),.Y(wire151_0_0));
NANDC2x1 inst_and_b151_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire151_0_1));
INVC inst_inv_b151_0_1 (.A(imd_wire151_0_1),.Y(wire151_0_1));
NANDC2x1 inst_and_b151_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire151_0_2));
INVC inst_inv_b151_0_2 (.A(imd_wire151_0_2),.Y(wire151_0_2));
NANDC2x1 inst_and_b151_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire151_0_3));
INVC inst_inv_b151_0_3 (.A(imd_wire151_0_3),.Y(wire151_0_3));
NANDC2x1 inst_and_b151_1_0 (.A(wire151_0_0),.B(wire151_0_1),.Y(imd_wire151_1_0));
INVC inst_inv_b151_1_0 (.A(imd_wire151_1_0),.Y(wire151_1_0));
NANDC2x1 inst_and_b151_1_1 (.A(wire151_0_2),.B(wire151_0_3),.Y(imd_wire151_1_1));
INVC inst_inv_b151_1_1 (.A(imd_wire151_1_1),.Y(wire151_1_1));
NANDC2x1 inst_and_b151_2_0 (.A(wire151_1_0),.B(wire151_1_1),.Y(imd_Y151));
INVC inst_inv_b151_2_0 (.A(imd_Y151),.Y(Y151));
NANDC2x1 inst_clockedAND_b151_151 (.A(CLK),.B(Y151),.Y(imd_YF151));
INVC inst_clockedinv_b151_151 (.A(imd_YF151),.Y(YF151));


NANDC2x1 inst_and_b152_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire152_0_0));
INVC inst_inv_b152_0_0 (.A(imd_wire152_0_0),.Y(wire152_0_0));
NANDC2x1 inst_and_b152_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire152_0_1));
INVC inst_inv_b152_0_1 (.A(imd_wire152_0_1),.Y(wire152_0_1));
NANDC2x1 inst_and_b152_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire152_0_2));
INVC inst_inv_b152_0_2 (.A(imd_wire152_0_2),.Y(wire152_0_2));
NANDC2x1 inst_and_b152_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire152_0_3));
INVC inst_inv_b152_0_3 (.A(imd_wire152_0_3),.Y(wire152_0_3));
NANDC2x1 inst_and_b152_1_0 (.A(wire152_0_0),.B(wire152_0_1),.Y(imd_wire152_1_0));
INVC inst_inv_b152_1_0 (.A(imd_wire152_1_0),.Y(wire152_1_0));
NANDC2x1 inst_and_b152_1_1 (.A(wire152_0_2),.B(wire152_0_3),.Y(imd_wire152_1_1));
INVC inst_inv_b152_1_1 (.A(imd_wire152_1_1),.Y(wire152_1_1));
NANDC2x1 inst_and_b152_2_0 (.A(wire152_1_0),.B(wire152_1_1),.Y(imd_Y152));
INVC inst_inv_b152_2_0 (.A(imd_Y152),.Y(Y152));
NANDC2x1 inst_clockedAND_b152_152 (.A(CLK),.B(Y152),.Y(imd_YF152));
INVC inst_clockedinv_b152_152 (.A(imd_YF152),.Y(YF152));


NANDC2x1 inst_and_b153_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire153_0_0));
INVC inst_inv_b153_0_0 (.A(imd_wire153_0_0),.Y(wire153_0_0));
NANDC2x1 inst_and_b153_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire153_0_1));
INVC inst_inv_b153_0_1 (.A(imd_wire153_0_1),.Y(wire153_0_1));
NANDC2x1 inst_and_b153_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire153_0_2));
INVC inst_inv_b153_0_2 (.A(imd_wire153_0_2),.Y(wire153_0_2));
NANDC2x1 inst_and_b153_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire153_0_3));
INVC inst_inv_b153_0_3 (.A(imd_wire153_0_3),.Y(wire153_0_3));
NANDC2x1 inst_and_b153_1_0 (.A(wire153_0_0),.B(wire153_0_1),.Y(imd_wire153_1_0));
INVC inst_inv_b153_1_0 (.A(imd_wire153_1_0),.Y(wire153_1_0));
NANDC2x1 inst_and_b153_1_1 (.A(wire153_0_2),.B(wire153_0_3),.Y(imd_wire153_1_1));
INVC inst_inv_b153_1_1 (.A(imd_wire153_1_1),.Y(wire153_1_1));
NANDC2x1 inst_and_b153_2_0 (.A(wire153_1_0),.B(wire153_1_1),.Y(imd_Y153));
INVC inst_inv_b153_2_0 (.A(imd_Y153),.Y(Y153));
NANDC2x1 inst_clockedAND_b153_153 (.A(CLK),.B(Y153),.Y(imd_YF153));
INVC inst_clockedinv_b153_153 (.A(imd_YF153),.Y(YF153));


NANDC2x1 inst_and_b154_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire154_0_0));
INVC inst_inv_b154_0_0 (.A(imd_wire154_0_0),.Y(wire154_0_0));
NANDC2x1 inst_and_b154_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire154_0_1));
INVC inst_inv_b154_0_1 (.A(imd_wire154_0_1),.Y(wire154_0_1));
NANDC2x1 inst_and_b154_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire154_0_2));
INVC inst_inv_b154_0_2 (.A(imd_wire154_0_2),.Y(wire154_0_2));
NANDC2x1 inst_and_b154_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire154_0_3));
INVC inst_inv_b154_0_3 (.A(imd_wire154_0_3),.Y(wire154_0_3));
NANDC2x1 inst_and_b154_1_0 (.A(wire154_0_0),.B(wire154_0_1),.Y(imd_wire154_1_0));
INVC inst_inv_b154_1_0 (.A(imd_wire154_1_0),.Y(wire154_1_0));
NANDC2x1 inst_and_b154_1_1 (.A(wire154_0_2),.B(wire154_0_3),.Y(imd_wire154_1_1));
INVC inst_inv_b154_1_1 (.A(imd_wire154_1_1),.Y(wire154_1_1));
NANDC2x1 inst_and_b154_2_0 (.A(wire154_1_0),.B(wire154_1_1),.Y(imd_Y154));
INVC inst_inv_b154_2_0 (.A(imd_Y154),.Y(Y154));
NANDC2x1 inst_clockedAND_b154_154 (.A(CLK),.B(Y154),.Y(imd_YF154));
INVC inst_clockedinv_b154_154 (.A(imd_YF154),.Y(YF154));


NANDC2x1 inst_and_b155_0_0 (.A(A0),.B(A1),.Y(imd_wire155_0_0));
INVC inst_inv_b155_0_0 (.A(imd_wire155_0_0),.Y(wire155_0_0));
NANDC2x1 inst_and_b155_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire155_0_1));
INVC inst_inv_b155_0_1 (.A(imd_wire155_0_1),.Y(wire155_0_1));
NANDC2x1 inst_and_b155_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire155_0_2));
INVC inst_inv_b155_0_2 (.A(imd_wire155_0_2),.Y(wire155_0_2));
NANDC2x1 inst_and_b155_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire155_0_3));
INVC inst_inv_b155_0_3 (.A(imd_wire155_0_3),.Y(wire155_0_3));
NANDC2x1 inst_and_b155_1_0 (.A(wire155_0_0),.B(wire155_0_1),.Y(imd_wire155_1_0));
INVC inst_inv_b155_1_0 (.A(imd_wire155_1_0),.Y(wire155_1_0));
NANDC2x1 inst_and_b155_1_1 (.A(wire155_0_2),.B(wire155_0_3),.Y(imd_wire155_1_1));
INVC inst_inv_b155_1_1 (.A(imd_wire155_1_1),.Y(wire155_1_1));
NANDC2x1 inst_and_b155_2_0 (.A(wire155_1_0),.B(wire155_1_1),.Y(imd_Y155));
INVC inst_inv_b155_2_0 (.A(imd_Y155),.Y(Y155));
NANDC2x1 inst_clockedAND_b155_155 (.A(CLK),.B(Y155),.Y(imd_YF155));
INVC inst_clockedinv_b155_155 (.A(imd_YF155),.Y(YF155));


NANDC2x1 inst_and_b156_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire156_0_0));
INVC inst_inv_b156_0_0 (.A(imd_wire156_0_0),.Y(wire156_0_0));
NANDC2x1 inst_and_b156_0_1 (.A(A2),.B(A3),.Y(imd_wire156_0_1));
INVC inst_inv_b156_0_1 (.A(imd_wire156_0_1),.Y(wire156_0_1));
NANDC2x1 inst_and_b156_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire156_0_2));
INVC inst_inv_b156_0_2 (.A(imd_wire156_0_2),.Y(wire156_0_2));
NANDC2x1 inst_and_b156_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire156_0_3));
INVC inst_inv_b156_0_3 (.A(imd_wire156_0_3),.Y(wire156_0_3));
NANDC2x1 inst_and_b156_1_0 (.A(wire156_0_0),.B(wire156_0_1),.Y(imd_wire156_1_0));
INVC inst_inv_b156_1_0 (.A(imd_wire156_1_0),.Y(wire156_1_0));
NANDC2x1 inst_and_b156_1_1 (.A(wire156_0_2),.B(wire156_0_3),.Y(imd_wire156_1_1));
INVC inst_inv_b156_1_1 (.A(imd_wire156_1_1),.Y(wire156_1_1));
NANDC2x1 inst_and_b156_2_0 (.A(wire156_1_0),.B(wire156_1_1),.Y(imd_Y156));
INVC inst_inv_b156_2_0 (.A(imd_Y156),.Y(Y156));
NANDC2x1 inst_clockedAND_b156_156 (.A(CLK),.B(Y156),.Y(imd_YF156));
INVC inst_clockedinv_b156_156 (.A(imd_YF156),.Y(YF156));


NANDC2x1 inst_and_b157_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire157_0_0));
INVC inst_inv_b157_0_0 (.A(imd_wire157_0_0),.Y(wire157_0_0));
NANDC2x1 inst_and_b157_0_1 (.A(A2),.B(A3),.Y(imd_wire157_0_1));
INVC inst_inv_b157_0_1 (.A(imd_wire157_0_1),.Y(wire157_0_1));
NANDC2x1 inst_and_b157_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire157_0_2));
INVC inst_inv_b157_0_2 (.A(imd_wire157_0_2),.Y(wire157_0_2));
NANDC2x1 inst_and_b157_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire157_0_3));
INVC inst_inv_b157_0_3 (.A(imd_wire157_0_3),.Y(wire157_0_3));
NANDC2x1 inst_and_b157_1_0 (.A(wire157_0_0),.B(wire157_0_1),.Y(imd_wire157_1_0));
INVC inst_inv_b157_1_0 (.A(imd_wire157_1_0),.Y(wire157_1_0));
NANDC2x1 inst_and_b157_1_1 (.A(wire157_0_2),.B(wire157_0_3),.Y(imd_wire157_1_1));
INVC inst_inv_b157_1_1 (.A(imd_wire157_1_1),.Y(wire157_1_1));
NANDC2x1 inst_and_b157_2_0 (.A(wire157_1_0),.B(wire157_1_1),.Y(imd_Y157));
INVC inst_inv_b157_2_0 (.A(imd_Y157),.Y(Y157));
NANDC2x1 inst_clockedAND_b157_157 (.A(CLK),.B(Y157),.Y(imd_YF157));
INVC inst_clockedinv_b157_157 (.A(imd_YF157),.Y(YF157));


NANDC2x1 inst_and_b158_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire158_0_0));
INVC inst_inv_b158_0_0 (.A(imd_wire158_0_0),.Y(wire158_0_0));
NANDC2x1 inst_and_b158_0_1 (.A(A2),.B(A3),.Y(imd_wire158_0_1));
INVC inst_inv_b158_0_1 (.A(imd_wire158_0_1),.Y(wire158_0_1));
NANDC2x1 inst_and_b158_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire158_0_2));
INVC inst_inv_b158_0_2 (.A(imd_wire158_0_2),.Y(wire158_0_2));
NANDC2x1 inst_and_b158_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire158_0_3));
INVC inst_inv_b158_0_3 (.A(imd_wire158_0_3),.Y(wire158_0_3));
NANDC2x1 inst_and_b158_1_0 (.A(wire158_0_0),.B(wire158_0_1),.Y(imd_wire158_1_0));
INVC inst_inv_b158_1_0 (.A(imd_wire158_1_0),.Y(wire158_1_0));
NANDC2x1 inst_and_b158_1_1 (.A(wire158_0_2),.B(wire158_0_3),.Y(imd_wire158_1_1));
INVC inst_inv_b158_1_1 (.A(imd_wire158_1_1),.Y(wire158_1_1));
NANDC2x1 inst_and_b158_2_0 (.A(wire158_1_0),.B(wire158_1_1),.Y(imd_Y158));
INVC inst_inv_b158_2_0 (.A(imd_Y158),.Y(Y158));
NANDC2x1 inst_clockedAND_b158_158 (.A(CLK),.B(Y158),.Y(imd_YF158));
INVC inst_clockedinv_b158_158 (.A(imd_YF158),.Y(YF158));


NANDC2x1 inst_and_b159_0_0 (.A(A0),.B(A1),.Y(imd_wire159_0_0));
INVC inst_inv_b159_0_0 (.A(imd_wire159_0_0),.Y(wire159_0_0));
NANDC2x1 inst_and_b159_0_1 (.A(A2),.B(A3),.Y(imd_wire159_0_1));
INVC inst_inv_b159_0_1 (.A(imd_wire159_0_1),.Y(wire159_0_1));
NANDC2x1 inst_and_b159_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire159_0_2));
INVC inst_inv_b159_0_2 (.A(imd_wire159_0_2),.Y(wire159_0_2));
NANDC2x1 inst_and_b159_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire159_0_3));
INVC inst_inv_b159_0_3 (.A(imd_wire159_0_3),.Y(wire159_0_3));
NANDC2x1 inst_and_b159_1_0 (.A(wire159_0_0),.B(wire159_0_1),.Y(imd_wire159_1_0));
INVC inst_inv_b159_1_0 (.A(imd_wire159_1_0),.Y(wire159_1_0));
NANDC2x1 inst_and_b159_1_1 (.A(wire159_0_2),.B(wire159_0_3),.Y(imd_wire159_1_1));
INVC inst_inv_b159_1_1 (.A(imd_wire159_1_1),.Y(wire159_1_1));
NANDC2x1 inst_and_b159_2_0 (.A(wire159_1_0),.B(wire159_1_1),.Y(imd_Y159));
INVC inst_inv_b159_2_0 (.A(imd_Y159),.Y(Y159));
NANDC2x1 inst_clockedAND_b159_159 (.A(CLK),.B(Y159),.Y(imd_YF159));
INVC inst_clockedinv_b159_159 (.A(imd_YF159),.Y(YF159));


NANDC2x1 inst_and_b160_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire160_0_0));
INVC inst_inv_b160_0_0 (.A(imd_wire160_0_0),.Y(wire160_0_0));
NANDC2x1 inst_and_b160_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire160_0_1));
INVC inst_inv_b160_0_1 (.A(imd_wire160_0_1),.Y(wire160_0_1));
NANDC2x1 inst_and_b160_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire160_0_2));
INVC inst_inv_b160_0_2 (.A(imd_wire160_0_2),.Y(wire160_0_2));
NANDC2x1 inst_and_b160_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire160_0_3));
INVC inst_inv_b160_0_3 (.A(imd_wire160_0_3),.Y(wire160_0_3));
NANDC2x1 inst_and_b160_1_0 (.A(wire160_0_0),.B(wire160_0_1),.Y(imd_wire160_1_0));
INVC inst_inv_b160_1_0 (.A(imd_wire160_1_0),.Y(wire160_1_0));
NANDC2x1 inst_and_b160_1_1 (.A(wire160_0_2),.B(wire160_0_3),.Y(imd_wire160_1_1));
INVC inst_inv_b160_1_1 (.A(imd_wire160_1_1),.Y(wire160_1_1));
NANDC2x1 inst_and_b160_2_0 (.A(wire160_1_0),.B(wire160_1_1),.Y(imd_Y160));
INVC inst_inv_b160_2_0 (.A(imd_Y160),.Y(Y160));
NANDC2x1 inst_clockedAND_b160_160 (.A(CLK),.B(Y160),.Y(imd_YF160));
INVC inst_clockedinv_b160_160 (.A(imd_YF160),.Y(YF160));


NANDC2x1 inst_and_b161_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire161_0_0));
INVC inst_inv_b161_0_0 (.A(imd_wire161_0_0),.Y(wire161_0_0));
NANDC2x1 inst_and_b161_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire161_0_1));
INVC inst_inv_b161_0_1 (.A(imd_wire161_0_1),.Y(wire161_0_1));
NANDC2x1 inst_and_b161_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire161_0_2));
INVC inst_inv_b161_0_2 (.A(imd_wire161_0_2),.Y(wire161_0_2));
NANDC2x1 inst_and_b161_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire161_0_3));
INVC inst_inv_b161_0_3 (.A(imd_wire161_0_3),.Y(wire161_0_3));
NANDC2x1 inst_and_b161_1_0 (.A(wire161_0_0),.B(wire161_0_1),.Y(imd_wire161_1_0));
INVC inst_inv_b161_1_0 (.A(imd_wire161_1_0),.Y(wire161_1_0));
NANDC2x1 inst_and_b161_1_1 (.A(wire161_0_2),.B(wire161_0_3),.Y(imd_wire161_1_1));
INVC inst_inv_b161_1_1 (.A(imd_wire161_1_1),.Y(wire161_1_1));
NANDC2x1 inst_and_b161_2_0 (.A(wire161_1_0),.B(wire161_1_1),.Y(imd_Y161));
INVC inst_inv_b161_2_0 (.A(imd_Y161),.Y(Y161));
NANDC2x1 inst_clockedAND_b161_161 (.A(CLK),.B(Y161),.Y(imd_YF161));
INVC inst_clockedinv_b161_161 (.A(imd_YF161),.Y(YF161));


NANDC2x1 inst_and_b162_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire162_0_0));
INVC inst_inv_b162_0_0 (.A(imd_wire162_0_0),.Y(wire162_0_0));
NANDC2x1 inst_and_b162_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire162_0_1));
INVC inst_inv_b162_0_1 (.A(imd_wire162_0_1),.Y(wire162_0_1));
NANDC2x1 inst_and_b162_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire162_0_2));
INVC inst_inv_b162_0_2 (.A(imd_wire162_0_2),.Y(wire162_0_2));
NANDC2x1 inst_and_b162_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire162_0_3));
INVC inst_inv_b162_0_3 (.A(imd_wire162_0_3),.Y(wire162_0_3));
NANDC2x1 inst_and_b162_1_0 (.A(wire162_0_0),.B(wire162_0_1),.Y(imd_wire162_1_0));
INVC inst_inv_b162_1_0 (.A(imd_wire162_1_0),.Y(wire162_1_0));
NANDC2x1 inst_and_b162_1_1 (.A(wire162_0_2),.B(wire162_0_3),.Y(imd_wire162_1_1));
INVC inst_inv_b162_1_1 (.A(imd_wire162_1_1),.Y(wire162_1_1));
NANDC2x1 inst_and_b162_2_0 (.A(wire162_1_0),.B(wire162_1_1),.Y(imd_Y162));
INVC inst_inv_b162_2_0 (.A(imd_Y162),.Y(Y162));
NANDC2x1 inst_clockedAND_b162_162 (.A(CLK),.B(Y162),.Y(imd_YF162));
INVC inst_clockedinv_b162_162 (.A(imd_YF162),.Y(YF162));


NANDC2x1 inst_and_b163_0_0 (.A(A0),.B(A1),.Y(imd_wire163_0_0));
INVC inst_inv_b163_0_0 (.A(imd_wire163_0_0),.Y(wire163_0_0));
NANDC2x1 inst_and_b163_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire163_0_1));
INVC inst_inv_b163_0_1 (.A(imd_wire163_0_1),.Y(wire163_0_1));
NANDC2x1 inst_and_b163_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire163_0_2));
INVC inst_inv_b163_0_2 (.A(imd_wire163_0_2),.Y(wire163_0_2));
NANDC2x1 inst_and_b163_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire163_0_3));
INVC inst_inv_b163_0_3 (.A(imd_wire163_0_3),.Y(wire163_0_3));
NANDC2x1 inst_and_b163_1_0 (.A(wire163_0_0),.B(wire163_0_1),.Y(imd_wire163_1_0));
INVC inst_inv_b163_1_0 (.A(imd_wire163_1_0),.Y(wire163_1_0));
NANDC2x1 inst_and_b163_1_1 (.A(wire163_0_2),.B(wire163_0_3),.Y(imd_wire163_1_1));
INVC inst_inv_b163_1_1 (.A(imd_wire163_1_1),.Y(wire163_1_1));
NANDC2x1 inst_and_b163_2_0 (.A(wire163_1_0),.B(wire163_1_1),.Y(imd_Y163));
INVC inst_inv_b163_2_0 (.A(imd_Y163),.Y(Y163));
NANDC2x1 inst_clockedAND_b163_163 (.A(CLK),.B(Y163),.Y(imd_YF163));
INVC inst_clockedinv_b163_163 (.A(imd_YF163),.Y(YF163));


NANDC2x1 inst_and_b164_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire164_0_0));
INVC inst_inv_b164_0_0 (.A(imd_wire164_0_0),.Y(wire164_0_0));
NANDC2x1 inst_and_b164_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire164_0_1));
INVC inst_inv_b164_0_1 (.A(imd_wire164_0_1),.Y(wire164_0_1));
NANDC2x1 inst_and_b164_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire164_0_2));
INVC inst_inv_b164_0_2 (.A(imd_wire164_0_2),.Y(wire164_0_2));
NANDC2x1 inst_and_b164_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire164_0_3));
INVC inst_inv_b164_0_3 (.A(imd_wire164_0_3),.Y(wire164_0_3));
NANDC2x1 inst_and_b164_1_0 (.A(wire164_0_0),.B(wire164_0_1),.Y(imd_wire164_1_0));
INVC inst_inv_b164_1_0 (.A(imd_wire164_1_0),.Y(wire164_1_0));
NANDC2x1 inst_and_b164_1_1 (.A(wire164_0_2),.B(wire164_0_3),.Y(imd_wire164_1_1));
INVC inst_inv_b164_1_1 (.A(imd_wire164_1_1),.Y(wire164_1_1));
NANDC2x1 inst_and_b164_2_0 (.A(wire164_1_0),.B(wire164_1_1),.Y(imd_Y164));
INVC inst_inv_b164_2_0 (.A(imd_Y164),.Y(Y164));
NANDC2x1 inst_clockedAND_b164_164 (.A(CLK),.B(Y164),.Y(imd_YF164));
INVC inst_clockedinv_b164_164 (.A(imd_YF164),.Y(YF164));


NANDC2x1 inst_and_b165_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire165_0_0));
INVC inst_inv_b165_0_0 (.A(imd_wire165_0_0),.Y(wire165_0_0));
NANDC2x1 inst_and_b165_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire165_0_1));
INVC inst_inv_b165_0_1 (.A(imd_wire165_0_1),.Y(wire165_0_1));
NANDC2x1 inst_and_b165_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire165_0_2));
INVC inst_inv_b165_0_2 (.A(imd_wire165_0_2),.Y(wire165_0_2));
NANDC2x1 inst_and_b165_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire165_0_3));
INVC inst_inv_b165_0_3 (.A(imd_wire165_0_3),.Y(wire165_0_3));
NANDC2x1 inst_and_b165_1_0 (.A(wire165_0_0),.B(wire165_0_1),.Y(imd_wire165_1_0));
INVC inst_inv_b165_1_0 (.A(imd_wire165_1_0),.Y(wire165_1_0));
NANDC2x1 inst_and_b165_1_1 (.A(wire165_0_2),.B(wire165_0_3),.Y(imd_wire165_1_1));
INVC inst_inv_b165_1_1 (.A(imd_wire165_1_1),.Y(wire165_1_1));
NANDC2x1 inst_and_b165_2_0 (.A(wire165_1_0),.B(wire165_1_1),.Y(imd_Y165));
INVC inst_inv_b165_2_0 (.A(imd_Y165),.Y(Y165));
NANDC2x1 inst_clockedAND_b165_165 (.A(CLK),.B(Y165),.Y(imd_YF165));
INVC inst_clockedinv_b165_165 (.A(imd_YF165),.Y(YF165));


NANDC2x1 inst_and_b166_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire166_0_0));
INVC inst_inv_b166_0_0 (.A(imd_wire166_0_0),.Y(wire166_0_0));
NANDC2x1 inst_and_b166_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire166_0_1));
INVC inst_inv_b166_0_1 (.A(imd_wire166_0_1),.Y(wire166_0_1));
NANDC2x1 inst_and_b166_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire166_0_2));
INVC inst_inv_b166_0_2 (.A(imd_wire166_0_2),.Y(wire166_0_2));
NANDC2x1 inst_and_b166_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire166_0_3));
INVC inst_inv_b166_0_3 (.A(imd_wire166_0_3),.Y(wire166_0_3));
NANDC2x1 inst_and_b166_1_0 (.A(wire166_0_0),.B(wire166_0_1),.Y(imd_wire166_1_0));
INVC inst_inv_b166_1_0 (.A(imd_wire166_1_0),.Y(wire166_1_0));
NANDC2x1 inst_and_b166_1_1 (.A(wire166_0_2),.B(wire166_0_3),.Y(imd_wire166_1_1));
INVC inst_inv_b166_1_1 (.A(imd_wire166_1_1),.Y(wire166_1_1));
NANDC2x1 inst_and_b166_2_0 (.A(wire166_1_0),.B(wire166_1_1),.Y(imd_Y166));
INVC inst_inv_b166_2_0 (.A(imd_Y166),.Y(Y166));
NANDC2x1 inst_clockedAND_b166_166 (.A(CLK),.B(Y166),.Y(imd_YF166));
INVC inst_clockedinv_b166_166 (.A(imd_YF166),.Y(YF166));


NANDC2x1 inst_and_b167_0_0 (.A(A0),.B(A1),.Y(imd_wire167_0_0));
INVC inst_inv_b167_0_0 (.A(imd_wire167_0_0),.Y(wire167_0_0));
NANDC2x1 inst_and_b167_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire167_0_1));
INVC inst_inv_b167_0_1 (.A(imd_wire167_0_1),.Y(wire167_0_1));
NANDC2x1 inst_and_b167_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire167_0_2));
INVC inst_inv_b167_0_2 (.A(imd_wire167_0_2),.Y(wire167_0_2));
NANDC2x1 inst_and_b167_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire167_0_3));
INVC inst_inv_b167_0_3 (.A(imd_wire167_0_3),.Y(wire167_0_3));
NANDC2x1 inst_and_b167_1_0 (.A(wire167_0_0),.B(wire167_0_1),.Y(imd_wire167_1_0));
INVC inst_inv_b167_1_0 (.A(imd_wire167_1_0),.Y(wire167_1_0));
NANDC2x1 inst_and_b167_1_1 (.A(wire167_0_2),.B(wire167_0_3),.Y(imd_wire167_1_1));
INVC inst_inv_b167_1_1 (.A(imd_wire167_1_1),.Y(wire167_1_1));
NANDC2x1 inst_and_b167_2_0 (.A(wire167_1_0),.B(wire167_1_1),.Y(imd_Y167));
INVC inst_inv_b167_2_0 (.A(imd_Y167),.Y(Y167));
NANDC2x1 inst_clockedAND_b167_167 (.A(CLK),.B(Y167),.Y(imd_YF167));
INVC inst_clockedinv_b167_167 (.A(imd_YF167),.Y(YF167));


NANDC2x1 inst_and_b168_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire168_0_0));
INVC inst_inv_b168_0_0 (.A(imd_wire168_0_0),.Y(wire168_0_0));
NANDC2x1 inst_and_b168_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire168_0_1));
INVC inst_inv_b168_0_1 (.A(imd_wire168_0_1),.Y(wire168_0_1));
NANDC2x1 inst_and_b168_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire168_0_2));
INVC inst_inv_b168_0_2 (.A(imd_wire168_0_2),.Y(wire168_0_2));
NANDC2x1 inst_and_b168_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire168_0_3));
INVC inst_inv_b168_0_3 (.A(imd_wire168_0_3),.Y(wire168_0_3));
NANDC2x1 inst_and_b168_1_0 (.A(wire168_0_0),.B(wire168_0_1),.Y(imd_wire168_1_0));
INVC inst_inv_b168_1_0 (.A(imd_wire168_1_0),.Y(wire168_1_0));
NANDC2x1 inst_and_b168_1_1 (.A(wire168_0_2),.B(wire168_0_3),.Y(imd_wire168_1_1));
INVC inst_inv_b168_1_1 (.A(imd_wire168_1_1),.Y(wire168_1_1));
NANDC2x1 inst_and_b168_2_0 (.A(wire168_1_0),.B(wire168_1_1),.Y(imd_Y168));
INVC inst_inv_b168_2_0 (.A(imd_Y168),.Y(Y168));
NANDC2x1 inst_clockedAND_b168_168 (.A(CLK),.B(Y168),.Y(imd_YF168));
INVC inst_clockedinv_b168_168 (.A(imd_YF168),.Y(YF168));


NANDC2x1 inst_and_b169_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire169_0_0));
INVC inst_inv_b169_0_0 (.A(imd_wire169_0_0),.Y(wire169_0_0));
NANDC2x1 inst_and_b169_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire169_0_1));
INVC inst_inv_b169_0_1 (.A(imd_wire169_0_1),.Y(wire169_0_1));
NANDC2x1 inst_and_b169_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire169_0_2));
INVC inst_inv_b169_0_2 (.A(imd_wire169_0_2),.Y(wire169_0_2));
NANDC2x1 inst_and_b169_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire169_0_3));
INVC inst_inv_b169_0_3 (.A(imd_wire169_0_3),.Y(wire169_0_3));
NANDC2x1 inst_and_b169_1_0 (.A(wire169_0_0),.B(wire169_0_1),.Y(imd_wire169_1_0));
INVC inst_inv_b169_1_0 (.A(imd_wire169_1_0),.Y(wire169_1_0));
NANDC2x1 inst_and_b169_1_1 (.A(wire169_0_2),.B(wire169_0_3),.Y(imd_wire169_1_1));
INVC inst_inv_b169_1_1 (.A(imd_wire169_1_1),.Y(wire169_1_1));
NANDC2x1 inst_and_b169_2_0 (.A(wire169_1_0),.B(wire169_1_1),.Y(imd_Y169));
INVC inst_inv_b169_2_0 (.A(imd_Y169),.Y(Y169));
NANDC2x1 inst_clockedAND_b169_169 (.A(CLK),.B(Y169),.Y(imd_YF169));
INVC inst_clockedinv_b169_169 (.A(imd_YF169),.Y(YF169));


NANDC2x1 inst_and_b170_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire170_0_0));
INVC inst_inv_b170_0_0 (.A(imd_wire170_0_0),.Y(wire170_0_0));
NANDC2x1 inst_and_b170_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire170_0_1));
INVC inst_inv_b170_0_1 (.A(imd_wire170_0_1),.Y(wire170_0_1));
NANDC2x1 inst_and_b170_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire170_0_2));
INVC inst_inv_b170_0_2 (.A(imd_wire170_0_2),.Y(wire170_0_2));
NANDC2x1 inst_and_b170_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire170_0_3));
INVC inst_inv_b170_0_3 (.A(imd_wire170_0_3),.Y(wire170_0_3));
NANDC2x1 inst_and_b170_1_0 (.A(wire170_0_0),.B(wire170_0_1),.Y(imd_wire170_1_0));
INVC inst_inv_b170_1_0 (.A(imd_wire170_1_0),.Y(wire170_1_0));
NANDC2x1 inst_and_b170_1_1 (.A(wire170_0_2),.B(wire170_0_3),.Y(imd_wire170_1_1));
INVC inst_inv_b170_1_1 (.A(imd_wire170_1_1),.Y(wire170_1_1));
NANDC2x1 inst_and_b170_2_0 (.A(wire170_1_0),.B(wire170_1_1),.Y(imd_Y170));
INVC inst_inv_b170_2_0 (.A(imd_Y170),.Y(Y170));
NANDC2x1 inst_clockedAND_b170_170 (.A(CLK),.B(Y170),.Y(imd_YF170));
INVC inst_clockedinv_b170_170 (.A(imd_YF170),.Y(YF170));


NANDC2x1 inst_and_b171_0_0 (.A(A0),.B(A1),.Y(imd_wire171_0_0));
INVC inst_inv_b171_0_0 (.A(imd_wire171_0_0),.Y(wire171_0_0));
NANDC2x1 inst_and_b171_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire171_0_1));
INVC inst_inv_b171_0_1 (.A(imd_wire171_0_1),.Y(wire171_0_1));
NANDC2x1 inst_and_b171_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire171_0_2));
INVC inst_inv_b171_0_2 (.A(imd_wire171_0_2),.Y(wire171_0_2));
NANDC2x1 inst_and_b171_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire171_0_3));
INVC inst_inv_b171_0_3 (.A(imd_wire171_0_3),.Y(wire171_0_3));
NANDC2x1 inst_and_b171_1_0 (.A(wire171_0_0),.B(wire171_0_1),.Y(imd_wire171_1_0));
INVC inst_inv_b171_1_0 (.A(imd_wire171_1_0),.Y(wire171_1_0));
NANDC2x1 inst_and_b171_1_1 (.A(wire171_0_2),.B(wire171_0_3),.Y(imd_wire171_1_1));
INVC inst_inv_b171_1_1 (.A(imd_wire171_1_1),.Y(wire171_1_1));
NANDC2x1 inst_and_b171_2_0 (.A(wire171_1_0),.B(wire171_1_1),.Y(imd_Y171));
INVC inst_inv_b171_2_0 (.A(imd_Y171),.Y(Y171));
NANDC2x1 inst_clockedAND_b171_171 (.A(CLK),.B(Y171),.Y(imd_YF171));
INVC inst_clockedinv_b171_171 (.A(imd_YF171),.Y(YF171));


NANDC2x1 inst_and_b172_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire172_0_0));
INVC inst_inv_b172_0_0 (.A(imd_wire172_0_0),.Y(wire172_0_0));
NANDC2x1 inst_and_b172_0_1 (.A(A2),.B(A3),.Y(imd_wire172_0_1));
INVC inst_inv_b172_0_1 (.A(imd_wire172_0_1),.Y(wire172_0_1));
NANDC2x1 inst_and_b172_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire172_0_2));
INVC inst_inv_b172_0_2 (.A(imd_wire172_0_2),.Y(wire172_0_2));
NANDC2x1 inst_and_b172_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire172_0_3));
INVC inst_inv_b172_0_3 (.A(imd_wire172_0_3),.Y(wire172_0_3));
NANDC2x1 inst_and_b172_1_0 (.A(wire172_0_0),.B(wire172_0_1),.Y(imd_wire172_1_0));
INVC inst_inv_b172_1_0 (.A(imd_wire172_1_0),.Y(wire172_1_0));
NANDC2x1 inst_and_b172_1_1 (.A(wire172_0_2),.B(wire172_0_3),.Y(imd_wire172_1_1));
INVC inst_inv_b172_1_1 (.A(imd_wire172_1_1),.Y(wire172_1_1));
NANDC2x1 inst_and_b172_2_0 (.A(wire172_1_0),.B(wire172_1_1),.Y(imd_Y172));
INVC inst_inv_b172_2_0 (.A(imd_Y172),.Y(Y172));
NANDC2x1 inst_clockedAND_b172_172 (.A(CLK),.B(Y172),.Y(imd_YF172));
INVC inst_clockedinv_b172_172 (.A(imd_YF172),.Y(YF172));


NANDC2x1 inst_and_b173_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire173_0_0));
INVC inst_inv_b173_0_0 (.A(imd_wire173_0_0),.Y(wire173_0_0));
NANDC2x1 inst_and_b173_0_1 (.A(A2),.B(A3),.Y(imd_wire173_0_1));
INVC inst_inv_b173_0_1 (.A(imd_wire173_0_1),.Y(wire173_0_1));
NANDC2x1 inst_and_b173_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire173_0_2));
INVC inst_inv_b173_0_2 (.A(imd_wire173_0_2),.Y(wire173_0_2));
NANDC2x1 inst_and_b173_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire173_0_3));
INVC inst_inv_b173_0_3 (.A(imd_wire173_0_3),.Y(wire173_0_3));
NANDC2x1 inst_and_b173_1_0 (.A(wire173_0_0),.B(wire173_0_1),.Y(imd_wire173_1_0));
INVC inst_inv_b173_1_0 (.A(imd_wire173_1_0),.Y(wire173_1_0));
NANDC2x1 inst_and_b173_1_1 (.A(wire173_0_2),.B(wire173_0_3),.Y(imd_wire173_1_1));
INVC inst_inv_b173_1_1 (.A(imd_wire173_1_1),.Y(wire173_1_1));
NANDC2x1 inst_and_b173_2_0 (.A(wire173_1_0),.B(wire173_1_1),.Y(imd_Y173));
INVC inst_inv_b173_2_0 (.A(imd_Y173),.Y(Y173));
NANDC2x1 inst_clockedAND_b173_173 (.A(CLK),.B(Y173),.Y(imd_YF173));
INVC inst_clockedinv_b173_173 (.A(imd_YF173),.Y(YF173));


NANDC2x1 inst_and_b174_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire174_0_0));
INVC inst_inv_b174_0_0 (.A(imd_wire174_0_0),.Y(wire174_0_0));
NANDC2x1 inst_and_b174_0_1 (.A(A2),.B(A3),.Y(imd_wire174_0_1));
INVC inst_inv_b174_0_1 (.A(imd_wire174_0_1),.Y(wire174_0_1));
NANDC2x1 inst_and_b174_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire174_0_2));
INVC inst_inv_b174_0_2 (.A(imd_wire174_0_2),.Y(wire174_0_2));
NANDC2x1 inst_and_b174_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire174_0_3));
INVC inst_inv_b174_0_3 (.A(imd_wire174_0_3),.Y(wire174_0_3));
NANDC2x1 inst_and_b174_1_0 (.A(wire174_0_0),.B(wire174_0_1),.Y(imd_wire174_1_0));
INVC inst_inv_b174_1_0 (.A(imd_wire174_1_0),.Y(wire174_1_0));
NANDC2x1 inst_and_b174_1_1 (.A(wire174_0_2),.B(wire174_0_3),.Y(imd_wire174_1_1));
INVC inst_inv_b174_1_1 (.A(imd_wire174_1_1),.Y(wire174_1_1));
NANDC2x1 inst_and_b174_2_0 (.A(wire174_1_0),.B(wire174_1_1),.Y(imd_Y174));
INVC inst_inv_b174_2_0 (.A(imd_Y174),.Y(Y174));
NANDC2x1 inst_clockedAND_b174_174 (.A(CLK),.B(Y174),.Y(imd_YF174));
INVC inst_clockedinv_b174_174 (.A(imd_YF174),.Y(YF174));


NANDC2x1 inst_and_b175_0_0 (.A(A0),.B(A1),.Y(imd_wire175_0_0));
INVC inst_inv_b175_0_0 (.A(imd_wire175_0_0),.Y(wire175_0_0));
NANDC2x1 inst_and_b175_0_1 (.A(A2),.B(A3),.Y(imd_wire175_0_1));
INVC inst_inv_b175_0_1 (.A(imd_wire175_0_1),.Y(wire175_0_1));
NANDC2x1 inst_and_b175_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire175_0_2));
INVC inst_inv_b175_0_2 (.A(imd_wire175_0_2),.Y(wire175_0_2));
NANDC2x1 inst_and_b175_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire175_0_3));
INVC inst_inv_b175_0_3 (.A(imd_wire175_0_3),.Y(wire175_0_3));
NANDC2x1 inst_and_b175_1_0 (.A(wire175_0_0),.B(wire175_0_1),.Y(imd_wire175_1_0));
INVC inst_inv_b175_1_0 (.A(imd_wire175_1_0),.Y(wire175_1_0));
NANDC2x1 inst_and_b175_1_1 (.A(wire175_0_2),.B(wire175_0_3),.Y(imd_wire175_1_1));
INVC inst_inv_b175_1_1 (.A(imd_wire175_1_1),.Y(wire175_1_1));
NANDC2x1 inst_and_b175_2_0 (.A(wire175_1_0),.B(wire175_1_1),.Y(imd_Y175));
INVC inst_inv_b175_2_0 (.A(imd_Y175),.Y(Y175));
NANDC2x1 inst_clockedAND_b175_175 (.A(CLK),.B(Y175),.Y(imd_YF175));
INVC inst_clockedinv_b175_175 (.A(imd_YF175),.Y(YF175));


NANDC2x1 inst_and_b176_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire176_0_0));
INVC inst_inv_b176_0_0 (.A(imd_wire176_0_0),.Y(wire176_0_0));
NANDC2x1 inst_and_b176_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire176_0_1));
INVC inst_inv_b176_0_1 (.A(imd_wire176_0_1),.Y(wire176_0_1));
NANDC2x1 inst_and_b176_0_2 (.A(A4),.B(A5),.Y(imd_wire176_0_2));
INVC inst_inv_b176_0_2 (.A(imd_wire176_0_2),.Y(wire176_0_2));
NANDC2x1 inst_and_b176_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire176_0_3));
INVC inst_inv_b176_0_3 (.A(imd_wire176_0_3),.Y(wire176_0_3));
NANDC2x1 inst_and_b176_1_0 (.A(wire176_0_0),.B(wire176_0_1),.Y(imd_wire176_1_0));
INVC inst_inv_b176_1_0 (.A(imd_wire176_1_0),.Y(wire176_1_0));
NANDC2x1 inst_and_b176_1_1 (.A(wire176_0_2),.B(wire176_0_3),.Y(imd_wire176_1_1));
INVC inst_inv_b176_1_1 (.A(imd_wire176_1_1),.Y(wire176_1_1));
NANDC2x1 inst_and_b176_2_0 (.A(wire176_1_0),.B(wire176_1_1),.Y(imd_Y176));
INVC inst_inv_b176_2_0 (.A(imd_Y176),.Y(Y176));
NANDC2x1 inst_clockedAND_b176_176 (.A(CLK),.B(Y176),.Y(imd_YF176));
INVC inst_clockedinv_b176_176 (.A(imd_YF176),.Y(YF176));


NANDC2x1 inst_and_b177_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire177_0_0));
INVC inst_inv_b177_0_0 (.A(imd_wire177_0_0),.Y(wire177_0_0));
NANDC2x1 inst_and_b177_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire177_0_1));
INVC inst_inv_b177_0_1 (.A(imd_wire177_0_1),.Y(wire177_0_1));
NANDC2x1 inst_and_b177_0_2 (.A(A4),.B(A5),.Y(imd_wire177_0_2));
INVC inst_inv_b177_0_2 (.A(imd_wire177_0_2),.Y(wire177_0_2));
NANDC2x1 inst_and_b177_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire177_0_3));
INVC inst_inv_b177_0_3 (.A(imd_wire177_0_3),.Y(wire177_0_3));
NANDC2x1 inst_and_b177_1_0 (.A(wire177_0_0),.B(wire177_0_1),.Y(imd_wire177_1_0));
INVC inst_inv_b177_1_0 (.A(imd_wire177_1_0),.Y(wire177_1_0));
NANDC2x1 inst_and_b177_1_1 (.A(wire177_0_2),.B(wire177_0_3),.Y(imd_wire177_1_1));
INVC inst_inv_b177_1_1 (.A(imd_wire177_1_1),.Y(wire177_1_1));
NANDC2x1 inst_and_b177_2_0 (.A(wire177_1_0),.B(wire177_1_1),.Y(imd_Y177));
INVC inst_inv_b177_2_0 (.A(imd_Y177),.Y(Y177));
NANDC2x1 inst_clockedAND_b177_177 (.A(CLK),.B(Y177),.Y(imd_YF177));
INVC inst_clockedinv_b177_177 (.A(imd_YF177),.Y(YF177));


NANDC2x1 inst_and_b178_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire178_0_0));
INVC inst_inv_b178_0_0 (.A(imd_wire178_0_0),.Y(wire178_0_0));
NANDC2x1 inst_and_b178_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire178_0_1));
INVC inst_inv_b178_0_1 (.A(imd_wire178_0_1),.Y(wire178_0_1));
NANDC2x1 inst_and_b178_0_2 (.A(A4),.B(A5),.Y(imd_wire178_0_2));
INVC inst_inv_b178_0_2 (.A(imd_wire178_0_2),.Y(wire178_0_2));
NANDC2x1 inst_and_b178_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire178_0_3));
INVC inst_inv_b178_0_3 (.A(imd_wire178_0_3),.Y(wire178_0_3));
NANDC2x1 inst_and_b178_1_0 (.A(wire178_0_0),.B(wire178_0_1),.Y(imd_wire178_1_0));
INVC inst_inv_b178_1_0 (.A(imd_wire178_1_0),.Y(wire178_1_0));
NANDC2x1 inst_and_b178_1_1 (.A(wire178_0_2),.B(wire178_0_3),.Y(imd_wire178_1_1));
INVC inst_inv_b178_1_1 (.A(imd_wire178_1_1),.Y(wire178_1_1));
NANDC2x1 inst_and_b178_2_0 (.A(wire178_1_0),.B(wire178_1_1),.Y(imd_Y178));
INVC inst_inv_b178_2_0 (.A(imd_Y178),.Y(Y178));
NANDC2x1 inst_clockedAND_b178_178 (.A(CLK),.B(Y178),.Y(imd_YF178));
INVC inst_clockedinv_b178_178 (.A(imd_YF178),.Y(YF178));


NANDC2x1 inst_and_b179_0_0 (.A(A0),.B(A1),.Y(imd_wire179_0_0));
INVC inst_inv_b179_0_0 (.A(imd_wire179_0_0),.Y(wire179_0_0));
NANDC2x1 inst_and_b179_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire179_0_1));
INVC inst_inv_b179_0_1 (.A(imd_wire179_0_1),.Y(wire179_0_1));
NANDC2x1 inst_and_b179_0_2 (.A(A4),.B(A5),.Y(imd_wire179_0_2));
INVC inst_inv_b179_0_2 (.A(imd_wire179_0_2),.Y(wire179_0_2));
NANDC2x1 inst_and_b179_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire179_0_3));
INVC inst_inv_b179_0_3 (.A(imd_wire179_0_3),.Y(wire179_0_3));
NANDC2x1 inst_and_b179_1_0 (.A(wire179_0_0),.B(wire179_0_1),.Y(imd_wire179_1_0));
INVC inst_inv_b179_1_0 (.A(imd_wire179_1_0),.Y(wire179_1_0));
NANDC2x1 inst_and_b179_1_1 (.A(wire179_0_2),.B(wire179_0_3),.Y(imd_wire179_1_1));
INVC inst_inv_b179_1_1 (.A(imd_wire179_1_1),.Y(wire179_1_1));
NANDC2x1 inst_and_b179_2_0 (.A(wire179_1_0),.B(wire179_1_1),.Y(imd_Y179));
INVC inst_inv_b179_2_0 (.A(imd_Y179),.Y(Y179));
NANDC2x1 inst_clockedAND_b179_179 (.A(CLK),.B(Y179),.Y(imd_YF179));
INVC inst_clockedinv_b179_179 (.A(imd_YF179),.Y(YF179));


NANDC2x1 inst_and_b180_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire180_0_0));
INVC inst_inv_b180_0_0 (.A(imd_wire180_0_0),.Y(wire180_0_0));
NANDC2x1 inst_and_b180_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire180_0_1));
INVC inst_inv_b180_0_1 (.A(imd_wire180_0_1),.Y(wire180_0_1));
NANDC2x1 inst_and_b180_0_2 (.A(A4),.B(A5),.Y(imd_wire180_0_2));
INVC inst_inv_b180_0_2 (.A(imd_wire180_0_2),.Y(wire180_0_2));
NANDC2x1 inst_and_b180_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire180_0_3));
INVC inst_inv_b180_0_3 (.A(imd_wire180_0_3),.Y(wire180_0_3));
NANDC2x1 inst_and_b180_1_0 (.A(wire180_0_0),.B(wire180_0_1),.Y(imd_wire180_1_0));
INVC inst_inv_b180_1_0 (.A(imd_wire180_1_0),.Y(wire180_1_0));
NANDC2x1 inst_and_b180_1_1 (.A(wire180_0_2),.B(wire180_0_3),.Y(imd_wire180_1_1));
INVC inst_inv_b180_1_1 (.A(imd_wire180_1_1),.Y(wire180_1_1));
NANDC2x1 inst_and_b180_2_0 (.A(wire180_1_0),.B(wire180_1_1),.Y(imd_Y180));
INVC inst_inv_b180_2_0 (.A(imd_Y180),.Y(Y180));
NANDC2x1 inst_clockedAND_b180_180 (.A(CLK),.B(Y180),.Y(imd_YF180));
INVC inst_clockedinv_b180_180 (.A(imd_YF180),.Y(YF180));


NANDC2x1 inst_and_b181_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire181_0_0));
INVC inst_inv_b181_0_0 (.A(imd_wire181_0_0),.Y(wire181_0_0));
NANDC2x1 inst_and_b181_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire181_0_1));
INVC inst_inv_b181_0_1 (.A(imd_wire181_0_1),.Y(wire181_0_1));
NANDC2x1 inst_and_b181_0_2 (.A(A4),.B(A5),.Y(imd_wire181_0_2));
INVC inst_inv_b181_0_2 (.A(imd_wire181_0_2),.Y(wire181_0_2));
NANDC2x1 inst_and_b181_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire181_0_3));
INVC inst_inv_b181_0_3 (.A(imd_wire181_0_3),.Y(wire181_0_3));
NANDC2x1 inst_and_b181_1_0 (.A(wire181_0_0),.B(wire181_0_1),.Y(imd_wire181_1_0));
INVC inst_inv_b181_1_0 (.A(imd_wire181_1_0),.Y(wire181_1_0));
NANDC2x1 inst_and_b181_1_1 (.A(wire181_0_2),.B(wire181_0_3),.Y(imd_wire181_1_1));
INVC inst_inv_b181_1_1 (.A(imd_wire181_1_1),.Y(wire181_1_1));
NANDC2x1 inst_and_b181_2_0 (.A(wire181_1_0),.B(wire181_1_1),.Y(imd_Y181));
INVC inst_inv_b181_2_0 (.A(imd_Y181),.Y(Y181));
NANDC2x1 inst_clockedAND_b181_181 (.A(CLK),.B(Y181),.Y(imd_YF181));
INVC inst_clockedinv_b181_181 (.A(imd_YF181),.Y(YF181));


NANDC2x1 inst_and_b182_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire182_0_0));
INVC inst_inv_b182_0_0 (.A(imd_wire182_0_0),.Y(wire182_0_0));
NANDC2x1 inst_and_b182_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire182_0_1));
INVC inst_inv_b182_0_1 (.A(imd_wire182_0_1),.Y(wire182_0_1));
NANDC2x1 inst_and_b182_0_2 (.A(A4),.B(A5),.Y(imd_wire182_0_2));
INVC inst_inv_b182_0_2 (.A(imd_wire182_0_2),.Y(wire182_0_2));
NANDC2x1 inst_and_b182_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire182_0_3));
INVC inst_inv_b182_0_3 (.A(imd_wire182_0_3),.Y(wire182_0_3));
NANDC2x1 inst_and_b182_1_0 (.A(wire182_0_0),.B(wire182_0_1),.Y(imd_wire182_1_0));
INVC inst_inv_b182_1_0 (.A(imd_wire182_1_0),.Y(wire182_1_0));
NANDC2x1 inst_and_b182_1_1 (.A(wire182_0_2),.B(wire182_0_3),.Y(imd_wire182_1_1));
INVC inst_inv_b182_1_1 (.A(imd_wire182_1_1),.Y(wire182_1_1));
NANDC2x1 inst_and_b182_2_0 (.A(wire182_1_0),.B(wire182_1_1),.Y(imd_Y182));
INVC inst_inv_b182_2_0 (.A(imd_Y182),.Y(Y182));
NANDC2x1 inst_clockedAND_b182_182 (.A(CLK),.B(Y182),.Y(imd_YF182));
INVC inst_clockedinv_b182_182 (.A(imd_YF182),.Y(YF182));


NANDC2x1 inst_and_b183_0_0 (.A(A0),.B(A1),.Y(imd_wire183_0_0));
INVC inst_inv_b183_0_0 (.A(imd_wire183_0_0),.Y(wire183_0_0));
NANDC2x1 inst_and_b183_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire183_0_1));
INVC inst_inv_b183_0_1 (.A(imd_wire183_0_1),.Y(wire183_0_1));
NANDC2x1 inst_and_b183_0_2 (.A(A4),.B(A5),.Y(imd_wire183_0_2));
INVC inst_inv_b183_0_2 (.A(imd_wire183_0_2),.Y(wire183_0_2));
NANDC2x1 inst_and_b183_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire183_0_3));
INVC inst_inv_b183_0_3 (.A(imd_wire183_0_3),.Y(wire183_0_3));
NANDC2x1 inst_and_b183_1_0 (.A(wire183_0_0),.B(wire183_0_1),.Y(imd_wire183_1_0));
INVC inst_inv_b183_1_0 (.A(imd_wire183_1_0),.Y(wire183_1_0));
NANDC2x1 inst_and_b183_1_1 (.A(wire183_0_2),.B(wire183_0_3),.Y(imd_wire183_1_1));
INVC inst_inv_b183_1_1 (.A(imd_wire183_1_1),.Y(wire183_1_1));
NANDC2x1 inst_and_b183_2_0 (.A(wire183_1_0),.B(wire183_1_1),.Y(imd_Y183));
INVC inst_inv_b183_2_0 (.A(imd_Y183),.Y(Y183));
NANDC2x1 inst_clockedAND_b183_183 (.A(CLK),.B(Y183),.Y(imd_YF183));
INVC inst_clockedinv_b183_183 (.A(imd_YF183),.Y(YF183));


NANDC2x1 inst_and_b184_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire184_0_0));
INVC inst_inv_b184_0_0 (.A(imd_wire184_0_0),.Y(wire184_0_0));
NANDC2x1 inst_and_b184_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire184_0_1));
INVC inst_inv_b184_0_1 (.A(imd_wire184_0_1),.Y(wire184_0_1));
NANDC2x1 inst_and_b184_0_2 (.A(A4),.B(A5),.Y(imd_wire184_0_2));
INVC inst_inv_b184_0_2 (.A(imd_wire184_0_2),.Y(wire184_0_2));
NANDC2x1 inst_and_b184_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire184_0_3));
INVC inst_inv_b184_0_3 (.A(imd_wire184_0_3),.Y(wire184_0_3));
NANDC2x1 inst_and_b184_1_0 (.A(wire184_0_0),.B(wire184_0_1),.Y(imd_wire184_1_0));
INVC inst_inv_b184_1_0 (.A(imd_wire184_1_0),.Y(wire184_1_0));
NANDC2x1 inst_and_b184_1_1 (.A(wire184_0_2),.B(wire184_0_3),.Y(imd_wire184_1_1));
INVC inst_inv_b184_1_1 (.A(imd_wire184_1_1),.Y(wire184_1_1));
NANDC2x1 inst_and_b184_2_0 (.A(wire184_1_0),.B(wire184_1_1),.Y(imd_Y184));
INVC inst_inv_b184_2_0 (.A(imd_Y184),.Y(Y184));
NANDC2x1 inst_clockedAND_b184_184 (.A(CLK),.B(Y184),.Y(imd_YF184));
INVC inst_clockedinv_b184_184 (.A(imd_YF184),.Y(YF184));


NANDC2x1 inst_and_b185_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire185_0_0));
INVC inst_inv_b185_0_0 (.A(imd_wire185_0_0),.Y(wire185_0_0));
NANDC2x1 inst_and_b185_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire185_0_1));
INVC inst_inv_b185_0_1 (.A(imd_wire185_0_1),.Y(wire185_0_1));
NANDC2x1 inst_and_b185_0_2 (.A(A4),.B(A5),.Y(imd_wire185_0_2));
INVC inst_inv_b185_0_2 (.A(imd_wire185_0_2),.Y(wire185_0_2));
NANDC2x1 inst_and_b185_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire185_0_3));
INVC inst_inv_b185_0_3 (.A(imd_wire185_0_3),.Y(wire185_0_3));
NANDC2x1 inst_and_b185_1_0 (.A(wire185_0_0),.B(wire185_0_1),.Y(imd_wire185_1_0));
INVC inst_inv_b185_1_0 (.A(imd_wire185_1_0),.Y(wire185_1_0));
NANDC2x1 inst_and_b185_1_1 (.A(wire185_0_2),.B(wire185_0_3),.Y(imd_wire185_1_1));
INVC inst_inv_b185_1_1 (.A(imd_wire185_1_1),.Y(wire185_1_1));
NANDC2x1 inst_and_b185_2_0 (.A(wire185_1_0),.B(wire185_1_1),.Y(imd_Y185));
INVC inst_inv_b185_2_0 (.A(imd_Y185),.Y(Y185));
NANDC2x1 inst_clockedAND_b185_185 (.A(CLK),.B(Y185),.Y(imd_YF185));
INVC inst_clockedinv_b185_185 (.A(imd_YF185),.Y(YF185));


NANDC2x1 inst_and_b186_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire186_0_0));
INVC inst_inv_b186_0_0 (.A(imd_wire186_0_0),.Y(wire186_0_0));
NANDC2x1 inst_and_b186_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire186_0_1));
INVC inst_inv_b186_0_1 (.A(imd_wire186_0_1),.Y(wire186_0_1));
NANDC2x1 inst_and_b186_0_2 (.A(A4),.B(A5),.Y(imd_wire186_0_2));
INVC inst_inv_b186_0_2 (.A(imd_wire186_0_2),.Y(wire186_0_2));
NANDC2x1 inst_and_b186_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire186_0_3));
INVC inst_inv_b186_0_3 (.A(imd_wire186_0_3),.Y(wire186_0_3));
NANDC2x1 inst_and_b186_1_0 (.A(wire186_0_0),.B(wire186_0_1),.Y(imd_wire186_1_0));
INVC inst_inv_b186_1_0 (.A(imd_wire186_1_0),.Y(wire186_1_0));
NANDC2x1 inst_and_b186_1_1 (.A(wire186_0_2),.B(wire186_0_3),.Y(imd_wire186_1_1));
INVC inst_inv_b186_1_1 (.A(imd_wire186_1_1),.Y(wire186_1_1));
NANDC2x1 inst_and_b186_2_0 (.A(wire186_1_0),.B(wire186_1_1),.Y(imd_Y186));
INVC inst_inv_b186_2_0 (.A(imd_Y186),.Y(Y186));
NANDC2x1 inst_clockedAND_b186_186 (.A(CLK),.B(Y186),.Y(imd_YF186));
INVC inst_clockedinv_b186_186 (.A(imd_YF186),.Y(YF186));


NANDC2x1 inst_and_b187_0_0 (.A(A0),.B(A1),.Y(imd_wire187_0_0));
INVC inst_inv_b187_0_0 (.A(imd_wire187_0_0),.Y(wire187_0_0));
NANDC2x1 inst_and_b187_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire187_0_1));
INVC inst_inv_b187_0_1 (.A(imd_wire187_0_1),.Y(wire187_0_1));
NANDC2x1 inst_and_b187_0_2 (.A(A4),.B(A5),.Y(imd_wire187_0_2));
INVC inst_inv_b187_0_2 (.A(imd_wire187_0_2),.Y(wire187_0_2));
NANDC2x1 inst_and_b187_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire187_0_3));
INVC inst_inv_b187_0_3 (.A(imd_wire187_0_3),.Y(wire187_0_3));
NANDC2x1 inst_and_b187_1_0 (.A(wire187_0_0),.B(wire187_0_1),.Y(imd_wire187_1_0));
INVC inst_inv_b187_1_0 (.A(imd_wire187_1_0),.Y(wire187_1_0));
NANDC2x1 inst_and_b187_1_1 (.A(wire187_0_2),.B(wire187_0_3),.Y(imd_wire187_1_1));
INVC inst_inv_b187_1_1 (.A(imd_wire187_1_1),.Y(wire187_1_1));
NANDC2x1 inst_and_b187_2_0 (.A(wire187_1_0),.B(wire187_1_1),.Y(imd_Y187));
INVC inst_inv_b187_2_0 (.A(imd_Y187),.Y(Y187));
NANDC2x1 inst_clockedAND_b187_187 (.A(CLK),.B(Y187),.Y(imd_YF187));
INVC inst_clockedinv_b187_187 (.A(imd_YF187),.Y(YF187));


NANDC2x1 inst_and_b188_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire188_0_0));
INVC inst_inv_b188_0_0 (.A(imd_wire188_0_0),.Y(wire188_0_0));
NANDC2x1 inst_and_b188_0_1 (.A(A2),.B(A3),.Y(imd_wire188_0_1));
INVC inst_inv_b188_0_1 (.A(imd_wire188_0_1),.Y(wire188_0_1));
NANDC2x1 inst_and_b188_0_2 (.A(A4),.B(A5),.Y(imd_wire188_0_2));
INVC inst_inv_b188_0_2 (.A(imd_wire188_0_2),.Y(wire188_0_2));
NANDC2x1 inst_and_b188_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire188_0_3));
INVC inst_inv_b188_0_3 (.A(imd_wire188_0_3),.Y(wire188_0_3));
NANDC2x1 inst_and_b188_1_0 (.A(wire188_0_0),.B(wire188_0_1),.Y(imd_wire188_1_0));
INVC inst_inv_b188_1_0 (.A(imd_wire188_1_0),.Y(wire188_1_0));
NANDC2x1 inst_and_b188_1_1 (.A(wire188_0_2),.B(wire188_0_3),.Y(imd_wire188_1_1));
INVC inst_inv_b188_1_1 (.A(imd_wire188_1_1),.Y(wire188_1_1));
NANDC2x1 inst_and_b188_2_0 (.A(wire188_1_0),.B(wire188_1_1),.Y(imd_Y188));
INVC inst_inv_b188_2_0 (.A(imd_Y188),.Y(Y188));
NANDC2x1 inst_clockedAND_b188_188 (.A(CLK),.B(Y188),.Y(imd_YF188));
INVC inst_clockedinv_b188_188 (.A(imd_YF188),.Y(YF188));


NANDC2x1 inst_and_b189_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire189_0_0));
INVC inst_inv_b189_0_0 (.A(imd_wire189_0_0),.Y(wire189_0_0));
NANDC2x1 inst_and_b189_0_1 (.A(A2),.B(A3),.Y(imd_wire189_0_1));
INVC inst_inv_b189_0_1 (.A(imd_wire189_0_1),.Y(wire189_0_1));
NANDC2x1 inst_and_b189_0_2 (.A(A4),.B(A5),.Y(imd_wire189_0_2));
INVC inst_inv_b189_0_2 (.A(imd_wire189_0_2),.Y(wire189_0_2));
NANDC2x1 inst_and_b189_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire189_0_3));
INVC inst_inv_b189_0_3 (.A(imd_wire189_0_3),.Y(wire189_0_3));
NANDC2x1 inst_and_b189_1_0 (.A(wire189_0_0),.B(wire189_0_1),.Y(imd_wire189_1_0));
INVC inst_inv_b189_1_0 (.A(imd_wire189_1_0),.Y(wire189_1_0));
NANDC2x1 inst_and_b189_1_1 (.A(wire189_0_2),.B(wire189_0_3),.Y(imd_wire189_1_1));
INVC inst_inv_b189_1_1 (.A(imd_wire189_1_1),.Y(wire189_1_1));
NANDC2x1 inst_and_b189_2_0 (.A(wire189_1_0),.B(wire189_1_1),.Y(imd_Y189));
INVC inst_inv_b189_2_0 (.A(imd_Y189),.Y(Y189));
NANDC2x1 inst_clockedAND_b189_189 (.A(CLK),.B(Y189),.Y(imd_YF189));
INVC inst_clockedinv_b189_189 (.A(imd_YF189),.Y(YF189));


NANDC2x1 inst_and_b190_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire190_0_0));
INVC inst_inv_b190_0_0 (.A(imd_wire190_0_0),.Y(wire190_0_0));
NANDC2x1 inst_and_b190_0_1 (.A(A2),.B(A3),.Y(imd_wire190_0_1));
INVC inst_inv_b190_0_1 (.A(imd_wire190_0_1),.Y(wire190_0_1));
NANDC2x1 inst_and_b190_0_2 (.A(A4),.B(A5),.Y(imd_wire190_0_2));
INVC inst_inv_b190_0_2 (.A(imd_wire190_0_2),.Y(wire190_0_2));
NANDC2x1 inst_and_b190_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire190_0_3));
INVC inst_inv_b190_0_3 (.A(imd_wire190_0_3),.Y(wire190_0_3));
NANDC2x1 inst_and_b190_1_0 (.A(wire190_0_0),.B(wire190_0_1),.Y(imd_wire190_1_0));
INVC inst_inv_b190_1_0 (.A(imd_wire190_1_0),.Y(wire190_1_0));
NANDC2x1 inst_and_b190_1_1 (.A(wire190_0_2),.B(wire190_0_3),.Y(imd_wire190_1_1));
INVC inst_inv_b190_1_1 (.A(imd_wire190_1_1),.Y(wire190_1_1));
NANDC2x1 inst_and_b190_2_0 (.A(wire190_1_0),.B(wire190_1_1),.Y(imd_Y190));
INVC inst_inv_b190_2_0 (.A(imd_Y190),.Y(Y190));
NANDC2x1 inst_clockedAND_b190_190 (.A(CLK),.B(Y190),.Y(imd_YF190));
INVC inst_clockedinv_b190_190 (.A(imd_YF190),.Y(YF190));


NANDC2x1 inst_and_b191_0_0 (.A(A0),.B(A1),.Y(imd_wire191_0_0));
INVC inst_inv_b191_0_0 (.A(imd_wire191_0_0),.Y(wire191_0_0));
NANDC2x1 inst_and_b191_0_1 (.A(A2),.B(A3),.Y(imd_wire191_0_1));
INVC inst_inv_b191_0_1 (.A(imd_wire191_0_1),.Y(wire191_0_1));
NANDC2x1 inst_and_b191_0_2 (.A(A4),.B(A5),.Y(imd_wire191_0_2));
INVC inst_inv_b191_0_2 (.A(imd_wire191_0_2),.Y(wire191_0_2));
NANDC2x1 inst_and_b191_0_3 (.A(A6_inv),.B(A7),.Y(imd_wire191_0_3));
INVC inst_inv_b191_0_3 (.A(imd_wire191_0_3),.Y(wire191_0_3));
NANDC2x1 inst_and_b191_1_0 (.A(wire191_0_0),.B(wire191_0_1),.Y(imd_wire191_1_0));
INVC inst_inv_b191_1_0 (.A(imd_wire191_1_0),.Y(wire191_1_0));
NANDC2x1 inst_and_b191_1_1 (.A(wire191_0_2),.B(wire191_0_3),.Y(imd_wire191_1_1));
INVC inst_inv_b191_1_1 (.A(imd_wire191_1_1),.Y(wire191_1_1));
NANDC2x1 inst_and_b191_2_0 (.A(wire191_1_0),.B(wire191_1_1),.Y(imd_Y191));
INVC inst_inv_b191_2_0 (.A(imd_Y191),.Y(Y191));
NANDC2x1 inst_clockedAND_b191_191 (.A(CLK),.B(Y191),.Y(imd_YF191));
INVC inst_clockedinv_b191_191 (.A(imd_YF191),.Y(YF191));


NANDC2x1 inst_and_b192_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire192_0_0));
INVC inst_inv_b192_0_0 (.A(imd_wire192_0_0),.Y(wire192_0_0));
NANDC2x1 inst_and_b192_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire192_0_1));
INVC inst_inv_b192_0_1 (.A(imd_wire192_0_1),.Y(wire192_0_1));
NANDC2x1 inst_and_b192_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire192_0_2));
INVC inst_inv_b192_0_2 (.A(imd_wire192_0_2),.Y(wire192_0_2));
NANDC2x1 inst_and_b192_0_3 (.A(A6),.B(A7),.Y(imd_wire192_0_3));
INVC inst_inv_b192_0_3 (.A(imd_wire192_0_3),.Y(wire192_0_3));
NANDC2x1 inst_and_b192_1_0 (.A(wire192_0_0),.B(wire192_0_1),.Y(imd_wire192_1_0));
INVC inst_inv_b192_1_0 (.A(imd_wire192_1_0),.Y(wire192_1_0));
NANDC2x1 inst_and_b192_1_1 (.A(wire192_0_2),.B(wire192_0_3),.Y(imd_wire192_1_1));
INVC inst_inv_b192_1_1 (.A(imd_wire192_1_1),.Y(wire192_1_1));
NANDC2x1 inst_and_b192_2_0 (.A(wire192_1_0),.B(wire192_1_1),.Y(imd_Y192));
INVC inst_inv_b192_2_0 (.A(imd_Y192),.Y(Y192));
NANDC2x1 inst_clockedAND_b192_192 (.A(CLK),.B(Y192),.Y(imd_YF192));
INVC inst_clockedinv_b192_192 (.A(imd_YF192),.Y(YF192));


NANDC2x1 inst_and_b193_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire193_0_0));
INVC inst_inv_b193_0_0 (.A(imd_wire193_0_0),.Y(wire193_0_0));
NANDC2x1 inst_and_b193_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire193_0_1));
INVC inst_inv_b193_0_1 (.A(imd_wire193_0_1),.Y(wire193_0_1));
NANDC2x1 inst_and_b193_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire193_0_2));
INVC inst_inv_b193_0_2 (.A(imd_wire193_0_2),.Y(wire193_0_2));
NANDC2x1 inst_and_b193_0_3 (.A(A6),.B(A7),.Y(imd_wire193_0_3));
INVC inst_inv_b193_0_3 (.A(imd_wire193_0_3),.Y(wire193_0_3));
NANDC2x1 inst_and_b193_1_0 (.A(wire193_0_0),.B(wire193_0_1),.Y(imd_wire193_1_0));
INVC inst_inv_b193_1_0 (.A(imd_wire193_1_0),.Y(wire193_1_0));
NANDC2x1 inst_and_b193_1_1 (.A(wire193_0_2),.B(wire193_0_3),.Y(imd_wire193_1_1));
INVC inst_inv_b193_1_1 (.A(imd_wire193_1_1),.Y(wire193_1_1));
NANDC2x1 inst_and_b193_2_0 (.A(wire193_1_0),.B(wire193_1_1),.Y(imd_Y193));
INVC inst_inv_b193_2_0 (.A(imd_Y193),.Y(Y193));
NANDC2x1 inst_clockedAND_b193_193 (.A(CLK),.B(Y193),.Y(imd_YF193));
INVC inst_clockedinv_b193_193 (.A(imd_YF193),.Y(YF193));


NANDC2x1 inst_and_b194_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire194_0_0));
INVC inst_inv_b194_0_0 (.A(imd_wire194_0_0),.Y(wire194_0_0));
NANDC2x1 inst_and_b194_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire194_0_1));
INVC inst_inv_b194_0_1 (.A(imd_wire194_0_1),.Y(wire194_0_1));
NANDC2x1 inst_and_b194_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire194_0_2));
INVC inst_inv_b194_0_2 (.A(imd_wire194_0_2),.Y(wire194_0_2));
NANDC2x1 inst_and_b194_0_3 (.A(A6),.B(A7),.Y(imd_wire194_0_3));
INVC inst_inv_b194_0_3 (.A(imd_wire194_0_3),.Y(wire194_0_3));
NANDC2x1 inst_and_b194_1_0 (.A(wire194_0_0),.B(wire194_0_1),.Y(imd_wire194_1_0));
INVC inst_inv_b194_1_0 (.A(imd_wire194_1_0),.Y(wire194_1_0));
NANDC2x1 inst_and_b194_1_1 (.A(wire194_0_2),.B(wire194_0_3),.Y(imd_wire194_1_1));
INVC inst_inv_b194_1_1 (.A(imd_wire194_1_1),.Y(wire194_1_1));
NANDC2x1 inst_and_b194_2_0 (.A(wire194_1_0),.B(wire194_1_1),.Y(imd_Y194));
INVC inst_inv_b194_2_0 (.A(imd_Y194),.Y(Y194));
NANDC2x1 inst_clockedAND_b194_194 (.A(CLK),.B(Y194),.Y(imd_YF194));
INVC inst_clockedinv_b194_194 (.A(imd_YF194),.Y(YF194));


NANDC2x1 inst_and_b195_0_0 (.A(A0),.B(A1),.Y(imd_wire195_0_0));
INVC inst_inv_b195_0_0 (.A(imd_wire195_0_0),.Y(wire195_0_0));
NANDC2x1 inst_and_b195_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire195_0_1));
INVC inst_inv_b195_0_1 (.A(imd_wire195_0_1),.Y(wire195_0_1));
NANDC2x1 inst_and_b195_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire195_0_2));
INVC inst_inv_b195_0_2 (.A(imd_wire195_0_2),.Y(wire195_0_2));
NANDC2x1 inst_and_b195_0_3 (.A(A6),.B(A7),.Y(imd_wire195_0_3));
INVC inst_inv_b195_0_3 (.A(imd_wire195_0_3),.Y(wire195_0_3));
NANDC2x1 inst_and_b195_1_0 (.A(wire195_0_0),.B(wire195_0_1),.Y(imd_wire195_1_0));
INVC inst_inv_b195_1_0 (.A(imd_wire195_1_0),.Y(wire195_1_0));
NANDC2x1 inst_and_b195_1_1 (.A(wire195_0_2),.B(wire195_0_3),.Y(imd_wire195_1_1));
INVC inst_inv_b195_1_1 (.A(imd_wire195_1_1),.Y(wire195_1_1));
NANDC2x1 inst_and_b195_2_0 (.A(wire195_1_0),.B(wire195_1_1),.Y(imd_Y195));
INVC inst_inv_b195_2_0 (.A(imd_Y195),.Y(Y195));
NANDC2x1 inst_clockedAND_b195_195 (.A(CLK),.B(Y195),.Y(imd_YF195));
INVC inst_clockedinv_b195_195 (.A(imd_YF195),.Y(YF195));


NANDC2x1 inst_and_b196_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire196_0_0));
INVC inst_inv_b196_0_0 (.A(imd_wire196_0_0),.Y(wire196_0_0));
NANDC2x1 inst_and_b196_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire196_0_1));
INVC inst_inv_b196_0_1 (.A(imd_wire196_0_1),.Y(wire196_0_1));
NANDC2x1 inst_and_b196_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire196_0_2));
INVC inst_inv_b196_0_2 (.A(imd_wire196_0_2),.Y(wire196_0_2));
NANDC2x1 inst_and_b196_0_3 (.A(A6),.B(A7),.Y(imd_wire196_0_3));
INVC inst_inv_b196_0_3 (.A(imd_wire196_0_3),.Y(wire196_0_3));
NANDC2x1 inst_and_b196_1_0 (.A(wire196_0_0),.B(wire196_0_1),.Y(imd_wire196_1_0));
INVC inst_inv_b196_1_0 (.A(imd_wire196_1_0),.Y(wire196_1_0));
NANDC2x1 inst_and_b196_1_1 (.A(wire196_0_2),.B(wire196_0_3),.Y(imd_wire196_1_1));
INVC inst_inv_b196_1_1 (.A(imd_wire196_1_1),.Y(wire196_1_1));
NANDC2x1 inst_and_b196_2_0 (.A(wire196_1_0),.B(wire196_1_1),.Y(imd_Y196));
INVC inst_inv_b196_2_0 (.A(imd_Y196),.Y(Y196));
NANDC2x1 inst_clockedAND_b196_196 (.A(CLK),.B(Y196),.Y(imd_YF196));
INVC inst_clockedinv_b196_196 (.A(imd_YF196),.Y(YF196));


NANDC2x1 inst_and_b197_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire197_0_0));
INVC inst_inv_b197_0_0 (.A(imd_wire197_0_0),.Y(wire197_0_0));
NANDC2x1 inst_and_b197_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire197_0_1));
INVC inst_inv_b197_0_1 (.A(imd_wire197_0_1),.Y(wire197_0_1));
NANDC2x1 inst_and_b197_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire197_0_2));
INVC inst_inv_b197_0_2 (.A(imd_wire197_0_2),.Y(wire197_0_2));
NANDC2x1 inst_and_b197_0_3 (.A(A6),.B(A7),.Y(imd_wire197_0_3));
INVC inst_inv_b197_0_3 (.A(imd_wire197_0_3),.Y(wire197_0_3));
NANDC2x1 inst_and_b197_1_0 (.A(wire197_0_0),.B(wire197_0_1),.Y(imd_wire197_1_0));
INVC inst_inv_b197_1_0 (.A(imd_wire197_1_0),.Y(wire197_1_0));
NANDC2x1 inst_and_b197_1_1 (.A(wire197_0_2),.B(wire197_0_3),.Y(imd_wire197_1_1));
INVC inst_inv_b197_1_1 (.A(imd_wire197_1_1),.Y(wire197_1_1));
NANDC2x1 inst_and_b197_2_0 (.A(wire197_1_0),.B(wire197_1_1),.Y(imd_Y197));
INVC inst_inv_b197_2_0 (.A(imd_Y197),.Y(Y197));
NANDC2x1 inst_clockedAND_b197_197 (.A(CLK),.B(Y197),.Y(imd_YF197));
INVC inst_clockedinv_b197_197 (.A(imd_YF197),.Y(YF197));


NANDC2x1 inst_and_b198_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire198_0_0));
INVC inst_inv_b198_0_0 (.A(imd_wire198_0_0),.Y(wire198_0_0));
NANDC2x1 inst_and_b198_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire198_0_1));
INVC inst_inv_b198_0_1 (.A(imd_wire198_0_1),.Y(wire198_0_1));
NANDC2x1 inst_and_b198_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire198_0_2));
INVC inst_inv_b198_0_2 (.A(imd_wire198_0_2),.Y(wire198_0_2));
NANDC2x1 inst_and_b198_0_3 (.A(A6),.B(A7),.Y(imd_wire198_0_3));
INVC inst_inv_b198_0_3 (.A(imd_wire198_0_3),.Y(wire198_0_3));
NANDC2x1 inst_and_b198_1_0 (.A(wire198_0_0),.B(wire198_0_1),.Y(imd_wire198_1_0));
INVC inst_inv_b198_1_0 (.A(imd_wire198_1_0),.Y(wire198_1_0));
NANDC2x1 inst_and_b198_1_1 (.A(wire198_0_2),.B(wire198_0_3),.Y(imd_wire198_1_1));
INVC inst_inv_b198_1_1 (.A(imd_wire198_1_1),.Y(wire198_1_1));
NANDC2x1 inst_and_b198_2_0 (.A(wire198_1_0),.B(wire198_1_1),.Y(imd_Y198));
INVC inst_inv_b198_2_0 (.A(imd_Y198),.Y(Y198));
NANDC2x1 inst_clockedAND_b198_198 (.A(CLK),.B(Y198),.Y(imd_YF198));
INVC inst_clockedinv_b198_198 (.A(imd_YF198),.Y(YF198));


NANDC2x1 inst_and_b199_0_0 (.A(A0),.B(A1),.Y(imd_wire199_0_0));
INVC inst_inv_b199_0_0 (.A(imd_wire199_0_0),.Y(wire199_0_0));
NANDC2x1 inst_and_b199_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire199_0_1));
INVC inst_inv_b199_0_1 (.A(imd_wire199_0_1),.Y(wire199_0_1));
NANDC2x1 inst_and_b199_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire199_0_2));
INVC inst_inv_b199_0_2 (.A(imd_wire199_0_2),.Y(wire199_0_2));
NANDC2x1 inst_and_b199_0_3 (.A(A6),.B(A7),.Y(imd_wire199_0_3));
INVC inst_inv_b199_0_3 (.A(imd_wire199_0_3),.Y(wire199_0_3));
NANDC2x1 inst_and_b199_1_0 (.A(wire199_0_0),.B(wire199_0_1),.Y(imd_wire199_1_0));
INVC inst_inv_b199_1_0 (.A(imd_wire199_1_0),.Y(wire199_1_0));
NANDC2x1 inst_and_b199_1_1 (.A(wire199_0_2),.B(wire199_0_3),.Y(imd_wire199_1_1));
INVC inst_inv_b199_1_1 (.A(imd_wire199_1_1),.Y(wire199_1_1));
NANDC2x1 inst_and_b199_2_0 (.A(wire199_1_0),.B(wire199_1_1),.Y(imd_Y199));
INVC inst_inv_b199_2_0 (.A(imd_Y199),.Y(Y199));
NANDC2x1 inst_clockedAND_b199_199 (.A(CLK),.B(Y199),.Y(imd_YF199));
INVC inst_clockedinv_b199_199 (.A(imd_YF199),.Y(YF199));


NANDC2x1 inst_and_b200_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire200_0_0));
INVC inst_inv_b200_0_0 (.A(imd_wire200_0_0),.Y(wire200_0_0));
NANDC2x1 inst_and_b200_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire200_0_1));
INVC inst_inv_b200_0_1 (.A(imd_wire200_0_1),.Y(wire200_0_1));
NANDC2x1 inst_and_b200_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire200_0_2));
INVC inst_inv_b200_0_2 (.A(imd_wire200_0_2),.Y(wire200_0_2));
NANDC2x1 inst_and_b200_0_3 (.A(A6),.B(A7),.Y(imd_wire200_0_3));
INVC inst_inv_b200_0_3 (.A(imd_wire200_0_3),.Y(wire200_0_3));
NANDC2x1 inst_and_b200_1_0 (.A(wire200_0_0),.B(wire200_0_1),.Y(imd_wire200_1_0));
INVC inst_inv_b200_1_0 (.A(imd_wire200_1_0),.Y(wire200_1_0));
NANDC2x1 inst_and_b200_1_1 (.A(wire200_0_2),.B(wire200_0_3),.Y(imd_wire200_1_1));
INVC inst_inv_b200_1_1 (.A(imd_wire200_1_1),.Y(wire200_1_1));
NANDC2x1 inst_and_b200_2_0 (.A(wire200_1_0),.B(wire200_1_1),.Y(imd_Y200));
INVC inst_inv_b200_2_0 (.A(imd_Y200),.Y(Y200));
NANDC2x1 inst_clockedAND_b200_200 (.A(CLK),.B(Y200),.Y(imd_YF200));
INVC inst_clockedinv_b200_200 (.A(imd_YF200),.Y(YF200));


NANDC2x1 inst_and_b201_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire201_0_0));
INVC inst_inv_b201_0_0 (.A(imd_wire201_0_0),.Y(wire201_0_0));
NANDC2x1 inst_and_b201_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire201_0_1));
INVC inst_inv_b201_0_1 (.A(imd_wire201_0_1),.Y(wire201_0_1));
NANDC2x1 inst_and_b201_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire201_0_2));
INVC inst_inv_b201_0_2 (.A(imd_wire201_0_2),.Y(wire201_0_2));
NANDC2x1 inst_and_b201_0_3 (.A(A6),.B(A7),.Y(imd_wire201_0_3));
INVC inst_inv_b201_0_3 (.A(imd_wire201_0_3),.Y(wire201_0_3));
NANDC2x1 inst_and_b201_1_0 (.A(wire201_0_0),.B(wire201_0_1),.Y(imd_wire201_1_0));
INVC inst_inv_b201_1_0 (.A(imd_wire201_1_0),.Y(wire201_1_0));
NANDC2x1 inst_and_b201_1_1 (.A(wire201_0_2),.B(wire201_0_3),.Y(imd_wire201_1_1));
INVC inst_inv_b201_1_1 (.A(imd_wire201_1_1),.Y(wire201_1_1));
NANDC2x1 inst_and_b201_2_0 (.A(wire201_1_0),.B(wire201_1_1),.Y(imd_Y201));
INVC inst_inv_b201_2_0 (.A(imd_Y201),.Y(Y201));
NANDC2x1 inst_clockedAND_b201_201 (.A(CLK),.B(Y201),.Y(imd_YF201));
INVC inst_clockedinv_b201_201 (.A(imd_YF201),.Y(YF201));


NANDC2x1 inst_and_b202_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire202_0_0));
INVC inst_inv_b202_0_0 (.A(imd_wire202_0_0),.Y(wire202_0_0));
NANDC2x1 inst_and_b202_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire202_0_1));
INVC inst_inv_b202_0_1 (.A(imd_wire202_0_1),.Y(wire202_0_1));
NANDC2x1 inst_and_b202_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire202_0_2));
INVC inst_inv_b202_0_2 (.A(imd_wire202_0_2),.Y(wire202_0_2));
NANDC2x1 inst_and_b202_0_3 (.A(A6),.B(A7),.Y(imd_wire202_0_3));
INVC inst_inv_b202_0_3 (.A(imd_wire202_0_3),.Y(wire202_0_3));
NANDC2x1 inst_and_b202_1_0 (.A(wire202_0_0),.B(wire202_0_1),.Y(imd_wire202_1_0));
INVC inst_inv_b202_1_0 (.A(imd_wire202_1_0),.Y(wire202_1_0));
NANDC2x1 inst_and_b202_1_1 (.A(wire202_0_2),.B(wire202_0_3),.Y(imd_wire202_1_1));
INVC inst_inv_b202_1_1 (.A(imd_wire202_1_1),.Y(wire202_1_1));
NANDC2x1 inst_and_b202_2_0 (.A(wire202_1_0),.B(wire202_1_1),.Y(imd_Y202));
INVC inst_inv_b202_2_0 (.A(imd_Y202),.Y(Y202));
NANDC2x1 inst_clockedAND_b202_202 (.A(CLK),.B(Y202),.Y(imd_YF202));
INVC inst_clockedinv_b202_202 (.A(imd_YF202),.Y(YF202));


NANDC2x1 inst_and_b203_0_0 (.A(A0),.B(A1),.Y(imd_wire203_0_0));
INVC inst_inv_b203_0_0 (.A(imd_wire203_0_0),.Y(wire203_0_0));
NANDC2x1 inst_and_b203_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire203_0_1));
INVC inst_inv_b203_0_1 (.A(imd_wire203_0_1),.Y(wire203_0_1));
NANDC2x1 inst_and_b203_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire203_0_2));
INVC inst_inv_b203_0_2 (.A(imd_wire203_0_2),.Y(wire203_0_2));
NANDC2x1 inst_and_b203_0_3 (.A(A6),.B(A7),.Y(imd_wire203_0_3));
INVC inst_inv_b203_0_3 (.A(imd_wire203_0_3),.Y(wire203_0_3));
NANDC2x1 inst_and_b203_1_0 (.A(wire203_0_0),.B(wire203_0_1),.Y(imd_wire203_1_0));
INVC inst_inv_b203_1_0 (.A(imd_wire203_1_0),.Y(wire203_1_0));
NANDC2x1 inst_and_b203_1_1 (.A(wire203_0_2),.B(wire203_0_3),.Y(imd_wire203_1_1));
INVC inst_inv_b203_1_1 (.A(imd_wire203_1_1),.Y(wire203_1_1));
NANDC2x1 inst_and_b203_2_0 (.A(wire203_1_0),.B(wire203_1_1),.Y(imd_Y203));
INVC inst_inv_b203_2_0 (.A(imd_Y203),.Y(Y203));
NANDC2x1 inst_clockedAND_b203_203 (.A(CLK),.B(Y203),.Y(imd_YF203));
INVC inst_clockedinv_b203_203 (.A(imd_YF203),.Y(YF203));


NANDC2x1 inst_and_b204_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire204_0_0));
INVC inst_inv_b204_0_0 (.A(imd_wire204_0_0),.Y(wire204_0_0));
NANDC2x1 inst_and_b204_0_1 (.A(A2),.B(A3),.Y(imd_wire204_0_1));
INVC inst_inv_b204_0_1 (.A(imd_wire204_0_1),.Y(wire204_0_1));
NANDC2x1 inst_and_b204_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire204_0_2));
INVC inst_inv_b204_0_2 (.A(imd_wire204_0_2),.Y(wire204_0_2));
NANDC2x1 inst_and_b204_0_3 (.A(A6),.B(A7),.Y(imd_wire204_0_3));
INVC inst_inv_b204_0_3 (.A(imd_wire204_0_3),.Y(wire204_0_3));
NANDC2x1 inst_and_b204_1_0 (.A(wire204_0_0),.B(wire204_0_1),.Y(imd_wire204_1_0));
INVC inst_inv_b204_1_0 (.A(imd_wire204_1_0),.Y(wire204_1_0));
NANDC2x1 inst_and_b204_1_1 (.A(wire204_0_2),.B(wire204_0_3),.Y(imd_wire204_1_1));
INVC inst_inv_b204_1_1 (.A(imd_wire204_1_1),.Y(wire204_1_1));
NANDC2x1 inst_and_b204_2_0 (.A(wire204_1_0),.B(wire204_1_1),.Y(imd_Y204));
INVC inst_inv_b204_2_0 (.A(imd_Y204),.Y(Y204));
NANDC2x1 inst_clockedAND_b204_204 (.A(CLK),.B(Y204),.Y(imd_YF204));
INVC inst_clockedinv_b204_204 (.A(imd_YF204),.Y(YF204));


NANDC2x1 inst_and_b205_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire205_0_0));
INVC inst_inv_b205_0_0 (.A(imd_wire205_0_0),.Y(wire205_0_0));
NANDC2x1 inst_and_b205_0_1 (.A(A2),.B(A3),.Y(imd_wire205_0_1));
INVC inst_inv_b205_0_1 (.A(imd_wire205_0_1),.Y(wire205_0_1));
NANDC2x1 inst_and_b205_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire205_0_2));
INVC inst_inv_b205_0_2 (.A(imd_wire205_0_2),.Y(wire205_0_2));
NANDC2x1 inst_and_b205_0_3 (.A(A6),.B(A7),.Y(imd_wire205_0_3));
INVC inst_inv_b205_0_3 (.A(imd_wire205_0_3),.Y(wire205_0_3));
NANDC2x1 inst_and_b205_1_0 (.A(wire205_0_0),.B(wire205_0_1),.Y(imd_wire205_1_0));
INVC inst_inv_b205_1_0 (.A(imd_wire205_1_0),.Y(wire205_1_0));
NANDC2x1 inst_and_b205_1_1 (.A(wire205_0_2),.B(wire205_0_3),.Y(imd_wire205_1_1));
INVC inst_inv_b205_1_1 (.A(imd_wire205_1_1),.Y(wire205_1_1));
NANDC2x1 inst_and_b205_2_0 (.A(wire205_1_0),.B(wire205_1_1),.Y(imd_Y205));
INVC inst_inv_b205_2_0 (.A(imd_Y205),.Y(Y205));
NANDC2x1 inst_clockedAND_b205_205 (.A(CLK),.B(Y205),.Y(imd_YF205));
INVC inst_clockedinv_b205_205 (.A(imd_YF205),.Y(YF205));


NANDC2x1 inst_and_b206_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire206_0_0));
INVC inst_inv_b206_0_0 (.A(imd_wire206_0_0),.Y(wire206_0_0));
NANDC2x1 inst_and_b206_0_1 (.A(A2),.B(A3),.Y(imd_wire206_0_1));
INVC inst_inv_b206_0_1 (.A(imd_wire206_0_1),.Y(wire206_0_1));
NANDC2x1 inst_and_b206_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire206_0_2));
INVC inst_inv_b206_0_2 (.A(imd_wire206_0_2),.Y(wire206_0_2));
NANDC2x1 inst_and_b206_0_3 (.A(A6),.B(A7),.Y(imd_wire206_0_3));
INVC inst_inv_b206_0_3 (.A(imd_wire206_0_3),.Y(wire206_0_3));
NANDC2x1 inst_and_b206_1_0 (.A(wire206_0_0),.B(wire206_0_1),.Y(imd_wire206_1_0));
INVC inst_inv_b206_1_0 (.A(imd_wire206_1_0),.Y(wire206_1_0));
NANDC2x1 inst_and_b206_1_1 (.A(wire206_0_2),.B(wire206_0_3),.Y(imd_wire206_1_1));
INVC inst_inv_b206_1_1 (.A(imd_wire206_1_1),.Y(wire206_1_1));
NANDC2x1 inst_and_b206_2_0 (.A(wire206_1_0),.B(wire206_1_1),.Y(imd_Y206));
INVC inst_inv_b206_2_0 (.A(imd_Y206),.Y(Y206));
NANDC2x1 inst_clockedAND_b206_206 (.A(CLK),.B(Y206),.Y(imd_YF206));
INVC inst_clockedinv_b206_206 (.A(imd_YF206),.Y(YF206));


NANDC2x1 inst_and_b207_0_0 (.A(A0),.B(A1),.Y(imd_wire207_0_0));
INVC inst_inv_b207_0_0 (.A(imd_wire207_0_0),.Y(wire207_0_0));
NANDC2x1 inst_and_b207_0_1 (.A(A2),.B(A3),.Y(imd_wire207_0_1));
INVC inst_inv_b207_0_1 (.A(imd_wire207_0_1),.Y(wire207_0_1));
NANDC2x1 inst_and_b207_0_2 (.A(A4_inv),.B(A5_inv),.Y(imd_wire207_0_2));
INVC inst_inv_b207_0_2 (.A(imd_wire207_0_2),.Y(wire207_0_2));
NANDC2x1 inst_and_b207_0_3 (.A(A6),.B(A7),.Y(imd_wire207_0_3));
INVC inst_inv_b207_0_3 (.A(imd_wire207_0_3),.Y(wire207_0_3));
NANDC2x1 inst_and_b207_1_0 (.A(wire207_0_0),.B(wire207_0_1),.Y(imd_wire207_1_0));
INVC inst_inv_b207_1_0 (.A(imd_wire207_1_0),.Y(wire207_1_0));
NANDC2x1 inst_and_b207_1_1 (.A(wire207_0_2),.B(wire207_0_3),.Y(imd_wire207_1_1));
INVC inst_inv_b207_1_1 (.A(imd_wire207_1_1),.Y(wire207_1_1));
NANDC2x1 inst_and_b207_2_0 (.A(wire207_1_0),.B(wire207_1_1),.Y(imd_Y207));
INVC inst_inv_b207_2_0 (.A(imd_Y207),.Y(Y207));
NANDC2x1 inst_clockedAND_b207_207 (.A(CLK),.B(Y207),.Y(imd_YF207));
INVC inst_clockedinv_b207_207 (.A(imd_YF207),.Y(YF207));


NANDC2x1 inst_and_b208_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire208_0_0));
INVC inst_inv_b208_0_0 (.A(imd_wire208_0_0),.Y(wire208_0_0));
NANDC2x1 inst_and_b208_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire208_0_1));
INVC inst_inv_b208_0_1 (.A(imd_wire208_0_1),.Y(wire208_0_1));
NANDC2x1 inst_and_b208_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire208_0_2));
INVC inst_inv_b208_0_2 (.A(imd_wire208_0_2),.Y(wire208_0_2));
NANDC2x1 inst_and_b208_0_3 (.A(A6),.B(A7),.Y(imd_wire208_0_3));
INVC inst_inv_b208_0_3 (.A(imd_wire208_0_3),.Y(wire208_0_3));
NANDC2x1 inst_and_b208_1_0 (.A(wire208_0_0),.B(wire208_0_1),.Y(imd_wire208_1_0));
INVC inst_inv_b208_1_0 (.A(imd_wire208_1_0),.Y(wire208_1_0));
NANDC2x1 inst_and_b208_1_1 (.A(wire208_0_2),.B(wire208_0_3),.Y(imd_wire208_1_1));
INVC inst_inv_b208_1_1 (.A(imd_wire208_1_1),.Y(wire208_1_1));
NANDC2x1 inst_and_b208_2_0 (.A(wire208_1_0),.B(wire208_1_1),.Y(imd_Y208));
INVC inst_inv_b208_2_0 (.A(imd_Y208),.Y(Y208));
NANDC2x1 inst_clockedAND_b208_208 (.A(CLK),.B(Y208),.Y(imd_YF208));
INVC inst_clockedinv_b208_208 (.A(imd_YF208),.Y(YF208));


NANDC2x1 inst_and_b209_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire209_0_0));
INVC inst_inv_b209_0_0 (.A(imd_wire209_0_0),.Y(wire209_0_0));
NANDC2x1 inst_and_b209_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire209_0_1));
INVC inst_inv_b209_0_1 (.A(imd_wire209_0_1),.Y(wire209_0_1));
NANDC2x1 inst_and_b209_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire209_0_2));
INVC inst_inv_b209_0_2 (.A(imd_wire209_0_2),.Y(wire209_0_2));
NANDC2x1 inst_and_b209_0_3 (.A(A6),.B(A7),.Y(imd_wire209_0_3));
INVC inst_inv_b209_0_3 (.A(imd_wire209_0_3),.Y(wire209_0_3));
NANDC2x1 inst_and_b209_1_0 (.A(wire209_0_0),.B(wire209_0_1),.Y(imd_wire209_1_0));
INVC inst_inv_b209_1_0 (.A(imd_wire209_1_0),.Y(wire209_1_0));
NANDC2x1 inst_and_b209_1_1 (.A(wire209_0_2),.B(wire209_0_3),.Y(imd_wire209_1_1));
INVC inst_inv_b209_1_1 (.A(imd_wire209_1_1),.Y(wire209_1_1));
NANDC2x1 inst_and_b209_2_0 (.A(wire209_1_0),.B(wire209_1_1),.Y(imd_Y209));
INVC inst_inv_b209_2_0 (.A(imd_Y209),.Y(Y209));
NANDC2x1 inst_clockedAND_b209_209 (.A(CLK),.B(Y209),.Y(imd_YF209));
INVC inst_clockedinv_b209_209 (.A(imd_YF209),.Y(YF209));


NANDC2x1 inst_and_b210_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire210_0_0));
INVC inst_inv_b210_0_0 (.A(imd_wire210_0_0),.Y(wire210_0_0));
NANDC2x1 inst_and_b210_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire210_0_1));
INVC inst_inv_b210_0_1 (.A(imd_wire210_0_1),.Y(wire210_0_1));
NANDC2x1 inst_and_b210_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire210_0_2));
INVC inst_inv_b210_0_2 (.A(imd_wire210_0_2),.Y(wire210_0_2));
NANDC2x1 inst_and_b210_0_3 (.A(A6),.B(A7),.Y(imd_wire210_0_3));
INVC inst_inv_b210_0_3 (.A(imd_wire210_0_3),.Y(wire210_0_3));
NANDC2x1 inst_and_b210_1_0 (.A(wire210_0_0),.B(wire210_0_1),.Y(imd_wire210_1_0));
INVC inst_inv_b210_1_0 (.A(imd_wire210_1_0),.Y(wire210_1_0));
NANDC2x1 inst_and_b210_1_1 (.A(wire210_0_2),.B(wire210_0_3),.Y(imd_wire210_1_1));
INVC inst_inv_b210_1_1 (.A(imd_wire210_1_1),.Y(wire210_1_1));
NANDC2x1 inst_and_b210_2_0 (.A(wire210_1_0),.B(wire210_1_1),.Y(imd_Y210));
INVC inst_inv_b210_2_0 (.A(imd_Y210),.Y(Y210));
NANDC2x1 inst_clockedAND_b210_210 (.A(CLK),.B(Y210),.Y(imd_YF210));
INVC inst_clockedinv_b210_210 (.A(imd_YF210),.Y(YF210));


NANDC2x1 inst_and_b211_0_0 (.A(A0),.B(A1),.Y(imd_wire211_0_0));
INVC inst_inv_b211_0_0 (.A(imd_wire211_0_0),.Y(wire211_0_0));
NANDC2x1 inst_and_b211_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire211_0_1));
INVC inst_inv_b211_0_1 (.A(imd_wire211_0_1),.Y(wire211_0_1));
NANDC2x1 inst_and_b211_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire211_0_2));
INVC inst_inv_b211_0_2 (.A(imd_wire211_0_2),.Y(wire211_0_2));
NANDC2x1 inst_and_b211_0_3 (.A(A6),.B(A7),.Y(imd_wire211_0_3));
INVC inst_inv_b211_0_3 (.A(imd_wire211_0_3),.Y(wire211_0_3));
NANDC2x1 inst_and_b211_1_0 (.A(wire211_0_0),.B(wire211_0_1),.Y(imd_wire211_1_0));
INVC inst_inv_b211_1_0 (.A(imd_wire211_1_0),.Y(wire211_1_0));
NANDC2x1 inst_and_b211_1_1 (.A(wire211_0_2),.B(wire211_0_3),.Y(imd_wire211_1_1));
INVC inst_inv_b211_1_1 (.A(imd_wire211_1_1),.Y(wire211_1_1));
NANDC2x1 inst_and_b211_2_0 (.A(wire211_1_0),.B(wire211_1_1),.Y(imd_Y211));
INVC inst_inv_b211_2_0 (.A(imd_Y211),.Y(Y211));
NANDC2x1 inst_clockedAND_b211_211 (.A(CLK),.B(Y211),.Y(imd_YF211));
INVC inst_clockedinv_b211_211 (.A(imd_YF211),.Y(YF211));


NANDC2x1 inst_and_b212_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire212_0_0));
INVC inst_inv_b212_0_0 (.A(imd_wire212_0_0),.Y(wire212_0_0));
NANDC2x1 inst_and_b212_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire212_0_1));
INVC inst_inv_b212_0_1 (.A(imd_wire212_0_1),.Y(wire212_0_1));
NANDC2x1 inst_and_b212_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire212_0_2));
INVC inst_inv_b212_0_2 (.A(imd_wire212_0_2),.Y(wire212_0_2));
NANDC2x1 inst_and_b212_0_3 (.A(A6),.B(A7),.Y(imd_wire212_0_3));
INVC inst_inv_b212_0_3 (.A(imd_wire212_0_3),.Y(wire212_0_3));
NANDC2x1 inst_and_b212_1_0 (.A(wire212_0_0),.B(wire212_0_1),.Y(imd_wire212_1_0));
INVC inst_inv_b212_1_0 (.A(imd_wire212_1_0),.Y(wire212_1_0));
NANDC2x1 inst_and_b212_1_1 (.A(wire212_0_2),.B(wire212_0_3),.Y(imd_wire212_1_1));
INVC inst_inv_b212_1_1 (.A(imd_wire212_1_1),.Y(wire212_1_1));
NANDC2x1 inst_and_b212_2_0 (.A(wire212_1_0),.B(wire212_1_1),.Y(imd_Y212));
INVC inst_inv_b212_2_0 (.A(imd_Y212),.Y(Y212));
NANDC2x1 inst_clockedAND_b212_212 (.A(CLK),.B(Y212),.Y(imd_YF212));
INVC inst_clockedinv_b212_212 (.A(imd_YF212),.Y(YF212));


NANDC2x1 inst_and_b213_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire213_0_0));
INVC inst_inv_b213_0_0 (.A(imd_wire213_0_0),.Y(wire213_0_0));
NANDC2x1 inst_and_b213_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire213_0_1));
INVC inst_inv_b213_0_1 (.A(imd_wire213_0_1),.Y(wire213_0_1));
NANDC2x1 inst_and_b213_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire213_0_2));
INVC inst_inv_b213_0_2 (.A(imd_wire213_0_2),.Y(wire213_0_2));
NANDC2x1 inst_and_b213_0_3 (.A(A6),.B(A7),.Y(imd_wire213_0_3));
INVC inst_inv_b213_0_3 (.A(imd_wire213_0_3),.Y(wire213_0_3));
NANDC2x1 inst_and_b213_1_0 (.A(wire213_0_0),.B(wire213_0_1),.Y(imd_wire213_1_0));
INVC inst_inv_b213_1_0 (.A(imd_wire213_1_0),.Y(wire213_1_0));
NANDC2x1 inst_and_b213_1_1 (.A(wire213_0_2),.B(wire213_0_3),.Y(imd_wire213_1_1));
INVC inst_inv_b213_1_1 (.A(imd_wire213_1_1),.Y(wire213_1_1));
NANDC2x1 inst_and_b213_2_0 (.A(wire213_1_0),.B(wire213_1_1),.Y(imd_Y213));
INVC inst_inv_b213_2_0 (.A(imd_Y213),.Y(Y213));
NANDC2x1 inst_clockedAND_b213_213 (.A(CLK),.B(Y213),.Y(imd_YF213));
INVC inst_clockedinv_b213_213 (.A(imd_YF213),.Y(YF213));


NANDC2x1 inst_and_b214_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire214_0_0));
INVC inst_inv_b214_0_0 (.A(imd_wire214_0_0),.Y(wire214_0_0));
NANDC2x1 inst_and_b214_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire214_0_1));
INVC inst_inv_b214_0_1 (.A(imd_wire214_0_1),.Y(wire214_0_1));
NANDC2x1 inst_and_b214_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire214_0_2));
INVC inst_inv_b214_0_2 (.A(imd_wire214_0_2),.Y(wire214_0_2));
NANDC2x1 inst_and_b214_0_3 (.A(A6),.B(A7),.Y(imd_wire214_0_3));
INVC inst_inv_b214_0_3 (.A(imd_wire214_0_3),.Y(wire214_0_3));
NANDC2x1 inst_and_b214_1_0 (.A(wire214_0_0),.B(wire214_0_1),.Y(imd_wire214_1_0));
INVC inst_inv_b214_1_0 (.A(imd_wire214_1_0),.Y(wire214_1_0));
NANDC2x1 inst_and_b214_1_1 (.A(wire214_0_2),.B(wire214_0_3),.Y(imd_wire214_1_1));
INVC inst_inv_b214_1_1 (.A(imd_wire214_1_1),.Y(wire214_1_1));
NANDC2x1 inst_and_b214_2_0 (.A(wire214_1_0),.B(wire214_1_1),.Y(imd_Y214));
INVC inst_inv_b214_2_0 (.A(imd_Y214),.Y(Y214));
NANDC2x1 inst_clockedAND_b214_214 (.A(CLK),.B(Y214),.Y(imd_YF214));
INVC inst_clockedinv_b214_214 (.A(imd_YF214),.Y(YF214));


NANDC2x1 inst_and_b215_0_0 (.A(A0),.B(A1),.Y(imd_wire215_0_0));
INVC inst_inv_b215_0_0 (.A(imd_wire215_0_0),.Y(wire215_0_0));
NANDC2x1 inst_and_b215_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire215_0_1));
INVC inst_inv_b215_0_1 (.A(imd_wire215_0_1),.Y(wire215_0_1));
NANDC2x1 inst_and_b215_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire215_0_2));
INVC inst_inv_b215_0_2 (.A(imd_wire215_0_2),.Y(wire215_0_2));
NANDC2x1 inst_and_b215_0_3 (.A(A6),.B(A7),.Y(imd_wire215_0_3));
INVC inst_inv_b215_0_3 (.A(imd_wire215_0_3),.Y(wire215_0_3));
NANDC2x1 inst_and_b215_1_0 (.A(wire215_0_0),.B(wire215_0_1),.Y(imd_wire215_1_0));
INVC inst_inv_b215_1_0 (.A(imd_wire215_1_0),.Y(wire215_1_0));
NANDC2x1 inst_and_b215_1_1 (.A(wire215_0_2),.B(wire215_0_3),.Y(imd_wire215_1_1));
INVC inst_inv_b215_1_1 (.A(imd_wire215_1_1),.Y(wire215_1_1));
NANDC2x1 inst_and_b215_2_0 (.A(wire215_1_0),.B(wire215_1_1),.Y(imd_Y215));
INVC inst_inv_b215_2_0 (.A(imd_Y215),.Y(Y215));
NANDC2x1 inst_clockedAND_b215_215 (.A(CLK),.B(Y215),.Y(imd_YF215));
INVC inst_clockedinv_b215_215 (.A(imd_YF215),.Y(YF215));


NANDC2x1 inst_and_b216_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire216_0_0));
INVC inst_inv_b216_0_0 (.A(imd_wire216_0_0),.Y(wire216_0_0));
NANDC2x1 inst_and_b216_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire216_0_1));
INVC inst_inv_b216_0_1 (.A(imd_wire216_0_1),.Y(wire216_0_1));
NANDC2x1 inst_and_b216_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire216_0_2));
INVC inst_inv_b216_0_2 (.A(imd_wire216_0_2),.Y(wire216_0_2));
NANDC2x1 inst_and_b216_0_3 (.A(A6),.B(A7),.Y(imd_wire216_0_3));
INVC inst_inv_b216_0_3 (.A(imd_wire216_0_3),.Y(wire216_0_3));
NANDC2x1 inst_and_b216_1_0 (.A(wire216_0_0),.B(wire216_0_1),.Y(imd_wire216_1_0));
INVC inst_inv_b216_1_0 (.A(imd_wire216_1_0),.Y(wire216_1_0));
NANDC2x1 inst_and_b216_1_1 (.A(wire216_0_2),.B(wire216_0_3),.Y(imd_wire216_1_1));
INVC inst_inv_b216_1_1 (.A(imd_wire216_1_1),.Y(wire216_1_1));
NANDC2x1 inst_and_b216_2_0 (.A(wire216_1_0),.B(wire216_1_1),.Y(imd_Y216));
INVC inst_inv_b216_2_0 (.A(imd_Y216),.Y(Y216));
NANDC2x1 inst_clockedAND_b216_216 (.A(CLK),.B(Y216),.Y(imd_YF216));
INVC inst_clockedinv_b216_216 (.A(imd_YF216),.Y(YF216));


NANDC2x1 inst_and_b217_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire217_0_0));
INVC inst_inv_b217_0_0 (.A(imd_wire217_0_0),.Y(wire217_0_0));
NANDC2x1 inst_and_b217_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire217_0_1));
INVC inst_inv_b217_0_1 (.A(imd_wire217_0_1),.Y(wire217_0_1));
NANDC2x1 inst_and_b217_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire217_0_2));
INVC inst_inv_b217_0_2 (.A(imd_wire217_0_2),.Y(wire217_0_2));
NANDC2x1 inst_and_b217_0_3 (.A(A6),.B(A7),.Y(imd_wire217_0_3));
INVC inst_inv_b217_0_3 (.A(imd_wire217_0_3),.Y(wire217_0_3));
NANDC2x1 inst_and_b217_1_0 (.A(wire217_0_0),.B(wire217_0_1),.Y(imd_wire217_1_0));
INVC inst_inv_b217_1_0 (.A(imd_wire217_1_0),.Y(wire217_1_0));
NANDC2x1 inst_and_b217_1_1 (.A(wire217_0_2),.B(wire217_0_3),.Y(imd_wire217_1_1));
INVC inst_inv_b217_1_1 (.A(imd_wire217_1_1),.Y(wire217_1_1));
NANDC2x1 inst_and_b217_2_0 (.A(wire217_1_0),.B(wire217_1_1),.Y(imd_Y217));
INVC inst_inv_b217_2_0 (.A(imd_Y217),.Y(Y217));
NANDC2x1 inst_clockedAND_b217_217 (.A(CLK),.B(Y217),.Y(imd_YF217));
INVC inst_clockedinv_b217_217 (.A(imd_YF217),.Y(YF217));


NANDC2x1 inst_and_b218_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire218_0_0));
INVC inst_inv_b218_0_0 (.A(imd_wire218_0_0),.Y(wire218_0_0));
NANDC2x1 inst_and_b218_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire218_0_1));
INVC inst_inv_b218_0_1 (.A(imd_wire218_0_1),.Y(wire218_0_1));
NANDC2x1 inst_and_b218_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire218_0_2));
INVC inst_inv_b218_0_2 (.A(imd_wire218_0_2),.Y(wire218_0_2));
NANDC2x1 inst_and_b218_0_3 (.A(A6),.B(A7),.Y(imd_wire218_0_3));
INVC inst_inv_b218_0_3 (.A(imd_wire218_0_3),.Y(wire218_0_3));
NANDC2x1 inst_and_b218_1_0 (.A(wire218_0_0),.B(wire218_0_1),.Y(imd_wire218_1_0));
INVC inst_inv_b218_1_0 (.A(imd_wire218_1_0),.Y(wire218_1_0));
NANDC2x1 inst_and_b218_1_1 (.A(wire218_0_2),.B(wire218_0_3),.Y(imd_wire218_1_1));
INVC inst_inv_b218_1_1 (.A(imd_wire218_1_1),.Y(wire218_1_1));
NANDC2x1 inst_and_b218_2_0 (.A(wire218_1_0),.B(wire218_1_1),.Y(imd_Y218));
INVC inst_inv_b218_2_0 (.A(imd_Y218),.Y(Y218));
NANDC2x1 inst_clockedAND_b218_218 (.A(CLK),.B(Y218),.Y(imd_YF218));
INVC inst_clockedinv_b218_218 (.A(imd_YF218),.Y(YF218));


NANDC2x1 inst_and_b219_0_0 (.A(A0),.B(A1),.Y(imd_wire219_0_0));
INVC inst_inv_b219_0_0 (.A(imd_wire219_0_0),.Y(wire219_0_0));
NANDC2x1 inst_and_b219_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire219_0_1));
INVC inst_inv_b219_0_1 (.A(imd_wire219_0_1),.Y(wire219_0_1));
NANDC2x1 inst_and_b219_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire219_0_2));
INVC inst_inv_b219_0_2 (.A(imd_wire219_0_2),.Y(wire219_0_2));
NANDC2x1 inst_and_b219_0_3 (.A(A6),.B(A7),.Y(imd_wire219_0_3));
INVC inst_inv_b219_0_3 (.A(imd_wire219_0_3),.Y(wire219_0_3));
NANDC2x1 inst_and_b219_1_0 (.A(wire219_0_0),.B(wire219_0_1),.Y(imd_wire219_1_0));
INVC inst_inv_b219_1_0 (.A(imd_wire219_1_0),.Y(wire219_1_0));
NANDC2x1 inst_and_b219_1_1 (.A(wire219_0_2),.B(wire219_0_3),.Y(imd_wire219_1_1));
INVC inst_inv_b219_1_1 (.A(imd_wire219_1_1),.Y(wire219_1_1));
NANDC2x1 inst_and_b219_2_0 (.A(wire219_1_0),.B(wire219_1_1),.Y(imd_Y219));
INVC inst_inv_b219_2_0 (.A(imd_Y219),.Y(Y219));
NANDC2x1 inst_clockedAND_b219_219 (.A(CLK),.B(Y219),.Y(imd_YF219));
INVC inst_clockedinv_b219_219 (.A(imd_YF219),.Y(YF219));


NANDC2x1 inst_and_b220_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire220_0_0));
INVC inst_inv_b220_0_0 (.A(imd_wire220_0_0),.Y(wire220_0_0));
NANDC2x1 inst_and_b220_0_1 (.A(A2),.B(A3),.Y(imd_wire220_0_1));
INVC inst_inv_b220_0_1 (.A(imd_wire220_0_1),.Y(wire220_0_1));
NANDC2x1 inst_and_b220_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire220_0_2));
INVC inst_inv_b220_0_2 (.A(imd_wire220_0_2),.Y(wire220_0_2));
NANDC2x1 inst_and_b220_0_3 (.A(A6),.B(A7),.Y(imd_wire220_0_3));
INVC inst_inv_b220_0_3 (.A(imd_wire220_0_3),.Y(wire220_0_3));
NANDC2x1 inst_and_b220_1_0 (.A(wire220_0_0),.B(wire220_0_1),.Y(imd_wire220_1_0));
INVC inst_inv_b220_1_0 (.A(imd_wire220_1_0),.Y(wire220_1_0));
NANDC2x1 inst_and_b220_1_1 (.A(wire220_0_2),.B(wire220_0_3),.Y(imd_wire220_1_1));
INVC inst_inv_b220_1_1 (.A(imd_wire220_1_1),.Y(wire220_1_1));
NANDC2x1 inst_and_b220_2_0 (.A(wire220_1_0),.B(wire220_1_1),.Y(imd_Y220));
INVC inst_inv_b220_2_0 (.A(imd_Y220),.Y(Y220));
NANDC2x1 inst_clockedAND_b220_220 (.A(CLK),.B(Y220),.Y(imd_YF220));
INVC inst_clockedinv_b220_220 (.A(imd_YF220),.Y(YF220));


NANDC2x1 inst_and_b221_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire221_0_0));
INVC inst_inv_b221_0_0 (.A(imd_wire221_0_0),.Y(wire221_0_0));
NANDC2x1 inst_and_b221_0_1 (.A(A2),.B(A3),.Y(imd_wire221_0_1));
INVC inst_inv_b221_0_1 (.A(imd_wire221_0_1),.Y(wire221_0_1));
NANDC2x1 inst_and_b221_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire221_0_2));
INVC inst_inv_b221_0_2 (.A(imd_wire221_0_2),.Y(wire221_0_2));
NANDC2x1 inst_and_b221_0_3 (.A(A6),.B(A7),.Y(imd_wire221_0_3));
INVC inst_inv_b221_0_3 (.A(imd_wire221_0_3),.Y(wire221_0_3));
NANDC2x1 inst_and_b221_1_0 (.A(wire221_0_0),.B(wire221_0_1),.Y(imd_wire221_1_0));
INVC inst_inv_b221_1_0 (.A(imd_wire221_1_0),.Y(wire221_1_0));
NANDC2x1 inst_and_b221_1_1 (.A(wire221_0_2),.B(wire221_0_3),.Y(imd_wire221_1_1));
INVC inst_inv_b221_1_1 (.A(imd_wire221_1_1),.Y(wire221_1_1));
NANDC2x1 inst_and_b221_2_0 (.A(wire221_1_0),.B(wire221_1_1),.Y(imd_Y221));
INVC inst_inv_b221_2_0 (.A(imd_Y221),.Y(Y221));
NANDC2x1 inst_clockedAND_b221_221 (.A(CLK),.B(Y221),.Y(imd_YF221));
INVC inst_clockedinv_b221_221 (.A(imd_YF221),.Y(YF221));


NANDC2x1 inst_and_b222_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire222_0_0));
INVC inst_inv_b222_0_0 (.A(imd_wire222_0_0),.Y(wire222_0_0));
NANDC2x1 inst_and_b222_0_1 (.A(A2),.B(A3),.Y(imd_wire222_0_1));
INVC inst_inv_b222_0_1 (.A(imd_wire222_0_1),.Y(wire222_0_1));
NANDC2x1 inst_and_b222_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire222_0_2));
INVC inst_inv_b222_0_2 (.A(imd_wire222_0_2),.Y(wire222_0_2));
NANDC2x1 inst_and_b222_0_3 (.A(A6),.B(A7),.Y(imd_wire222_0_3));
INVC inst_inv_b222_0_3 (.A(imd_wire222_0_3),.Y(wire222_0_3));
NANDC2x1 inst_and_b222_1_0 (.A(wire222_0_0),.B(wire222_0_1),.Y(imd_wire222_1_0));
INVC inst_inv_b222_1_0 (.A(imd_wire222_1_0),.Y(wire222_1_0));
NANDC2x1 inst_and_b222_1_1 (.A(wire222_0_2),.B(wire222_0_3),.Y(imd_wire222_1_1));
INVC inst_inv_b222_1_1 (.A(imd_wire222_1_1),.Y(wire222_1_1));
NANDC2x1 inst_and_b222_2_0 (.A(wire222_1_0),.B(wire222_1_1),.Y(imd_Y222));
INVC inst_inv_b222_2_0 (.A(imd_Y222),.Y(Y222));
NANDC2x1 inst_clockedAND_b222_222 (.A(CLK),.B(Y222),.Y(imd_YF222));
INVC inst_clockedinv_b222_222 (.A(imd_YF222),.Y(YF222));


NANDC2x1 inst_and_b223_0_0 (.A(A0),.B(A1),.Y(imd_wire223_0_0));
INVC inst_inv_b223_0_0 (.A(imd_wire223_0_0),.Y(wire223_0_0));
NANDC2x1 inst_and_b223_0_1 (.A(A2),.B(A3),.Y(imd_wire223_0_1));
INVC inst_inv_b223_0_1 (.A(imd_wire223_0_1),.Y(wire223_0_1));
NANDC2x1 inst_and_b223_0_2 (.A(A4),.B(A5_inv),.Y(imd_wire223_0_2));
INVC inst_inv_b223_0_2 (.A(imd_wire223_0_2),.Y(wire223_0_2));
NANDC2x1 inst_and_b223_0_3 (.A(A6),.B(A7),.Y(imd_wire223_0_3));
INVC inst_inv_b223_0_3 (.A(imd_wire223_0_3),.Y(wire223_0_3));
NANDC2x1 inst_and_b223_1_0 (.A(wire223_0_0),.B(wire223_0_1),.Y(imd_wire223_1_0));
INVC inst_inv_b223_1_0 (.A(imd_wire223_1_0),.Y(wire223_1_0));
NANDC2x1 inst_and_b223_1_1 (.A(wire223_0_2),.B(wire223_0_3),.Y(imd_wire223_1_1));
INVC inst_inv_b223_1_1 (.A(imd_wire223_1_1),.Y(wire223_1_1));
NANDC2x1 inst_and_b223_2_0 (.A(wire223_1_0),.B(wire223_1_1),.Y(imd_Y223));
INVC inst_inv_b223_2_0 (.A(imd_Y223),.Y(Y223));
NANDC2x1 inst_clockedAND_b223_223 (.A(CLK),.B(Y223),.Y(imd_YF223));
INVC inst_clockedinv_b223_223 (.A(imd_YF223),.Y(YF223));


NANDC2x1 inst_and_b224_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire224_0_0));
INVC inst_inv_b224_0_0 (.A(imd_wire224_0_0),.Y(wire224_0_0));
NANDC2x1 inst_and_b224_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire224_0_1));
INVC inst_inv_b224_0_1 (.A(imd_wire224_0_1),.Y(wire224_0_1));
NANDC2x1 inst_and_b224_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire224_0_2));
INVC inst_inv_b224_0_2 (.A(imd_wire224_0_2),.Y(wire224_0_2));
NANDC2x1 inst_and_b224_0_3 (.A(A6),.B(A7),.Y(imd_wire224_0_3));
INVC inst_inv_b224_0_3 (.A(imd_wire224_0_3),.Y(wire224_0_3));
NANDC2x1 inst_and_b224_1_0 (.A(wire224_0_0),.B(wire224_0_1),.Y(imd_wire224_1_0));
INVC inst_inv_b224_1_0 (.A(imd_wire224_1_0),.Y(wire224_1_0));
NANDC2x1 inst_and_b224_1_1 (.A(wire224_0_2),.B(wire224_0_3),.Y(imd_wire224_1_1));
INVC inst_inv_b224_1_1 (.A(imd_wire224_1_1),.Y(wire224_1_1));
NANDC2x1 inst_and_b224_2_0 (.A(wire224_1_0),.B(wire224_1_1),.Y(imd_Y224));
INVC inst_inv_b224_2_0 (.A(imd_Y224),.Y(Y224));
NANDC2x1 inst_clockedAND_b224_224 (.A(CLK),.B(Y224),.Y(imd_YF224));
INVC inst_clockedinv_b224_224 (.A(imd_YF224),.Y(YF224));


NANDC2x1 inst_and_b225_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire225_0_0));
INVC inst_inv_b225_0_0 (.A(imd_wire225_0_0),.Y(wire225_0_0));
NANDC2x1 inst_and_b225_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire225_0_1));
INVC inst_inv_b225_0_1 (.A(imd_wire225_0_1),.Y(wire225_0_1));
NANDC2x1 inst_and_b225_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire225_0_2));
INVC inst_inv_b225_0_2 (.A(imd_wire225_0_2),.Y(wire225_0_2));
NANDC2x1 inst_and_b225_0_3 (.A(A6),.B(A7),.Y(imd_wire225_0_3));
INVC inst_inv_b225_0_3 (.A(imd_wire225_0_3),.Y(wire225_0_3));
NANDC2x1 inst_and_b225_1_0 (.A(wire225_0_0),.B(wire225_0_1),.Y(imd_wire225_1_0));
INVC inst_inv_b225_1_0 (.A(imd_wire225_1_0),.Y(wire225_1_0));
NANDC2x1 inst_and_b225_1_1 (.A(wire225_0_2),.B(wire225_0_3),.Y(imd_wire225_1_1));
INVC inst_inv_b225_1_1 (.A(imd_wire225_1_1),.Y(wire225_1_1));
NANDC2x1 inst_and_b225_2_0 (.A(wire225_1_0),.B(wire225_1_1),.Y(imd_Y225));
INVC inst_inv_b225_2_0 (.A(imd_Y225),.Y(Y225));
NANDC2x1 inst_clockedAND_b225_225 (.A(CLK),.B(Y225),.Y(imd_YF225));
INVC inst_clockedinv_b225_225 (.A(imd_YF225),.Y(YF225));


NANDC2x1 inst_and_b226_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire226_0_0));
INVC inst_inv_b226_0_0 (.A(imd_wire226_0_0),.Y(wire226_0_0));
NANDC2x1 inst_and_b226_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire226_0_1));
INVC inst_inv_b226_0_1 (.A(imd_wire226_0_1),.Y(wire226_0_1));
NANDC2x1 inst_and_b226_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire226_0_2));
INVC inst_inv_b226_0_2 (.A(imd_wire226_0_2),.Y(wire226_0_2));
NANDC2x1 inst_and_b226_0_3 (.A(A6),.B(A7),.Y(imd_wire226_0_3));
INVC inst_inv_b226_0_3 (.A(imd_wire226_0_3),.Y(wire226_0_3));
NANDC2x1 inst_and_b226_1_0 (.A(wire226_0_0),.B(wire226_0_1),.Y(imd_wire226_1_0));
INVC inst_inv_b226_1_0 (.A(imd_wire226_1_0),.Y(wire226_1_0));
NANDC2x1 inst_and_b226_1_1 (.A(wire226_0_2),.B(wire226_0_3),.Y(imd_wire226_1_1));
INVC inst_inv_b226_1_1 (.A(imd_wire226_1_1),.Y(wire226_1_1));
NANDC2x1 inst_and_b226_2_0 (.A(wire226_1_0),.B(wire226_1_1),.Y(imd_Y226));
INVC inst_inv_b226_2_0 (.A(imd_Y226),.Y(Y226));
NANDC2x1 inst_clockedAND_b226_226 (.A(CLK),.B(Y226),.Y(imd_YF226));
INVC inst_clockedinv_b226_226 (.A(imd_YF226),.Y(YF226));


NANDC2x1 inst_and_b227_0_0 (.A(A0),.B(A1),.Y(imd_wire227_0_0));
INVC inst_inv_b227_0_0 (.A(imd_wire227_0_0),.Y(wire227_0_0));
NANDC2x1 inst_and_b227_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire227_0_1));
INVC inst_inv_b227_0_1 (.A(imd_wire227_0_1),.Y(wire227_0_1));
NANDC2x1 inst_and_b227_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire227_0_2));
INVC inst_inv_b227_0_2 (.A(imd_wire227_0_2),.Y(wire227_0_2));
NANDC2x1 inst_and_b227_0_3 (.A(A6),.B(A7),.Y(imd_wire227_0_3));
INVC inst_inv_b227_0_3 (.A(imd_wire227_0_3),.Y(wire227_0_3));
NANDC2x1 inst_and_b227_1_0 (.A(wire227_0_0),.B(wire227_0_1),.Y(imd_wire227_1_0));
INVC inst_inv_b227_1_0 (.A(imd_wire227_1_0),.Y(wire227_1_0));
NANDC2x1 inst_and_b227_1_1 (.A(wire227_0_2),.B(wire227_0_3),.Y(imd_wire227_1_1));
INVC inst_inv_b227_1_1 (.A(imd_wire227_1_1),.Y(wire227_1_1));
NANDC2x1 inst_and_b227_2_0 (.A(wire227_1_0),.B(wire227_1_1),.Y(imd_Y227));
INVC inst_inv_b227_2_0 (.A(imd_Y227),.Y(Y227));
NANDC2x1 inst_clockedAND_b227_227 (.A(CLK),.B(Y227),.Y(imd_YF227));
INVC inst_clockedinv_b227_227 (.A(imd_YF227),.Y(YF227));


NANDC2x1 inst_and_b228_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire228_0_0));
INVC inst_inv_b228_0_0 (.A(imd_wire228_0_0),.Y(wire228_0_0));
NANDC2x1 inst_and_b228_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire228_0_1));
INVC inst_inv_b228_0_1 (.A(imd_wire228_0_1),.Y(wire228_0_1));
NANDC2x1 inst_and_b228_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire228_0_2));
INVC inst_inv_b228_0_2 (.A(imd_wire228_0_2),.Y(wire228_0_2));
NANDC2x1 inst_and_b228_0_3 (.A(A6),.B(A7),.Y(imd_wire228_0_3));
INVC inst_inv_b228_0_3 (.A(imd_wire228_0_3),.Y(wire228_0_3));
NANDC2x1 inst_and_b228_1_0 (.A(wire228_0_0),.B(wire228_0_1),.Y(imd_wire228_1_0));
INVC inst_inv_b228_1_0 (.A(imd_wire228_1_0),.Y(wire228_1_0));
NANDC2x1 inst_and_b228_1_1 (.A(wire228_0_2),.B(wire228_0_3),.Y(imd_wire228_1_1));
INVC inst_inv_b228_1_1 (.A(imd_wire228_1_1),.Y(wire228_1_1));
NANDC2x1 inst_and_b228_2_0 (.A(wire228_1_0),.B(wire228_1_1),.Y(imd_Y228));
INVC inst_inv_b228_2_0 (.A(imd_Y228),.Y(Y228));
NANDC2x1 inst_clockedAND_b228_228 (.A(CLK),.B(Y228),.Y(imd_YF228));
INVC inst_clockedinv_b228_228 (.A(imd_YF228),.Y(YF228));


NANDC2x1 inst_and_b229_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire229_0_0));
INVC inst_inv_b229_0_0 (.A(imd_wire229_0_0),.Y(wire229_0_0));
NANDC2x1 inst_and_b229_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire229_0_1));
INVC inst_inv_b229_0_1 (.A(imd_wire229_0_1),.Y(wire229_0_1));
NANDC2x1 inst_and_b229_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire229_0_2));
INVC inst_inv_b229_0_2 (.A(imd_wire229_0_2),.Y(wire229_0_2));
NANDC2x1 inst_and_b229_0_3 (.A(A6),.B(A7),.Y(imd_wire229_0_3));
INVC inst_inv_b229_0_3 (.A(imd_wire229_0_3),.Y(wire229_0_3));
NANDC2x1 inst_and_b229_1_0 (.A(wire229_0_0),.B(wire229_0_1),.Y(imd_wire229_1_0));
INVC inst_inv_b229_1_0 (.A(imd_wire229_1_0),.Y(wire229_1_0));
NANDC2x1 inst_and_b229_1_1 (.A(wire229_0_2),.B(wire229_0_3),.Y(imd_wire229_1_1));
INVC inst_inv_b229_1_1 (.A(imd_wire229_1_1),.Y(wire229_1_1));
NANDC2x1 inst_and_b229_2_0 (.A(wire229_1_0),.B(wire229_1_1),.Y(imd_Y229));
INVC inst_inv_b229_2_0 (.A(imd_Y229),.Y(Y229));
NANDC2x1 inst_clockedAND_b229_229 (.A(CLK),.B(Y229),.Y(imd_YF229));
INVC inst_clockedinv_b229_229 (.A(imd_YF229),.Y(YF229));


NANDC2x1 inst_and_b230_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire230_0_0));
INVC inst_inv_b230_0_0 (.A(imd_wire230_0_0),.Y(wire230_0_0));
NANDC2x1 inst_and_b230_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire230_0_1));
INVC inst_inv_b230_0_1 (.A(imd_wire230_0_1),.Y(wire230_0_1));
NANDC2x1 inst_and_b230_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire230_0_2));
INVC inst_inv_b230_0_2 (.A(imd_wire230_0_2),.Y(wire230_0_2));
NANDC2x1 inst_and_b230_0_3 (.A(A6),.B(A7),.Y(imd_wire230_0_3));
INVC inst_inv_b230_0_3 (.A(imd_wire230_0_3),.Y(wire230_0_3));
NANDC2x1 inst_and_b230_1_0 (.A(wire230_0_0),.B(wire230_0_1),.Y(imd_wire230_1_0));
INVC inst_inv_b230_1_0 (.A(imd_wire230_1_0),.Y(wire230_1_0));
NANDC2x1 inst_and_b230_1_1 (.A(wire230_0_2),.B(wire230_0_3),.Y(imd_wire230_1_1));
INVC inst_inv_b230_1_1 (.A(imd_wire230_1_1),.Y(wire230_1_1));
NANDC2x1 inst_and_b230_2_0 (.A(wire230_1_0),.B(wire230_1_1),.Y(imd_Y230));
INVC inst_inv_b230_2_0 (.A(imd_Y230),.Y(Y230));
NANDC2x1 inst_clockedAND_b230_230 (.A(CLK),.B(Y230),.Y(imd_YF230));
INVC inst_clockedinv_b230_230 (.A(imd_YF230),.Y(YF230));


NANDC2x1 inst_and_b231_0_0 (.A(A0),.B(A1),.Y(imd_wire231_0_0));
INVC inst_inv_b231_0_0 (.A(imd_wire231_0_0),.Y(wire231_0_0));
NANDC2x1 inst_and_b231_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire231_0_1));
INVC inst_inv_b231_0_1 (.A(imd_wire231_0_1),.Y(wire231_0_1));
NANDC2x1 inst_and_b231_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire231_0_2));
INVC inst_inv_b231_0_2 (.A(imd_wire231_0_2),.Y(wire231_0_2));
NANDC2x1 inst_and_b231_0_3 (.A(A6),.B(A7),.Y(imd_wire231_0_3));
INVC inst_inv_b231_0_3 (.A(imd_wire231_0_3),.Y(wire231_0_3));
NANDC2x1 inst_and_b231_1_0 (.A(wire231_0_0),.B(wire231_0_1),.Y(imd_wire231_1_0));
INVC inst_inv_b231_1_0 (.A(imd_wire231_1_0),.Y(wire231_1_0));
NANDC2x1 inst_and_b231_1_1 (.A(wire231_0_2),.B(wire231_0_3),.Y(imd_wire231_1_1));
INVC inst_inv_b231_1_1 (.A(imd_wire231_1_1),.Y(wire231_1_1));
NANDC2x1 inst_and_b231_2_0 (.A(wire231_1_0),.B(wire231_1_1),.Y(imd_Y231));
INVC inst_inv_b231_2_0 (.A(imd_Y231),.Y(Y231));
NANDC2x1 inst_clockedAND_b231_231 (.A(CLK),.B(Y231),.Y(imd_YF231));
INVC inst_clockedinv_b231_231 (.A(imd_YF231),.Y(YF231));


NANDC2x1 inst_and_b232_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire232_0_0));
INVC inst_inv_b232_0_0 (.A(imd_wire232_0_0),.Y(wire232_0_0));
NANDC2x1 inst_and_b232_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire232_0_1));
INVC inst_inv_b232_0_1 (.A(imd_wire232_0_1),.Y(wire232_0_1));
NANDC2x1 inst_and_b232_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire232_0_2));
INVC inst_inv_b232_0_2 (.A(imd_wire232_0_2),.Y(wire232_0_2));
NANDC2x1 inst_and_b232_0_3 (.A(A6),.B(A7),.Y(imd_wire232_0_3));
INVC inst_inv_b232_0_3 (.A(imd_wire232_0_3),.Y(wire232_0_3));
NANDC2x1 inst_and_b232_1_0 (.A(wire232_0_0),.B(wire232_0_1),.Y(imd_wire232_1_0));
INVC inst_inv_b232_1_0 (.A(imd_wire232_1_0),.Y(wire232_1_0));
NANDC2x1 inst_and_b232_1_1 (.A(wire232_0_2),.B(wire232_0_3),.Y(imd_wire232_1_1));
INVC inst_inv_b232_1_1 (.A(imd_wire232_1_1),.Y(wire232_1_1));
NANDC2x1 inst_and_b232_2_0 (.A(wire232_1_0),.B(wire232_1_1),.Y(imd_Y232));
INVC inst_inv_b232_2_0 (.A(imd_Y232),.Y(Y232));
NANDC2x1 inst_clockedAND_b232_232 (.A(CLK),.B(Y232),.Y(imd_YF232));
INVC inst_clockedinv_b232_232 (.A(imd_YF232),.Y(YF232));


NANDC2x1 inst_and_b233_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire233_0_0));
INVC inst_inv_b233_0_0 (.A(imd_wire233_0_0),.Y(wire233_0_0));
NANDC2x1 inst_and_b233_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire233_0_1));
INVC inst_inv_b233_0_1 (.A(imd_wire233_0_1),.Y(wire233_0_1));
NANDC2x1 inst_and_b233_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire233_0_2));
INVC inst_inv_b233_0_2 (.A(imd_wire233_0_2),.Y(wire233_0_2));
NANDC2x1 inst_and_b233_0_3 (.A(A6),.B(A7),.Y(imd_wire233_0_3));
INVC inst_inv_b233_0_3 (.A(imd_wire233_0_3),.Y(wire233_0_3));
NANDC2x1 inst_and_b233_1_0 (.A(wire233_0_0),.B(wire233_0_1),.Y(imd_wire233_1_0));
INVC inst_inv_b233_1_0 (.A(imd_wire233_1_0),.Y(wire233_1_0));
NANDC2x1 inst_and_b233_1_1 (.A(wire233_0_2),.B(wire233_0_3),.Y(imd_wire233_1_1));
INVC inst_inv_b233_1_1 (.A(imd_wire233_1_1),.Y(wire233_1_1));
NANDC2x1 inst_and_b233_2_0 (.A(wire233_1_0),.B(wire233_1_1),.Y(imd_Y233));
INVC inst_inv_b233_2_0 (.A(imd_Y233),.Y(Y233));
NANDC2x1 inst_clockedAND_b233_233 (.A(CLK),.B(Y233),.Y(imd_YF233));
INVC inst_clockedinv_b233_233 (.A(imd_YF233),.Y(YF233));


NANDC2x1 inst_and_b234_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire234_0_0));
INVC inst_inv_b234_0_0 (.A(imd_wire234_0_0),.Y(wire234_0_0));
NANDC2x1 inst_and_b234_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire234_0_1));
INVC inst_inv_b234_0_1 (.A(imd_wire234_0_1),.Y(wire234_0_1));
NANDC2x1 inst_and_b234_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire234_0_2));
INVC inst_inv_b234_0_2 (.A(imd_wire234_0_2),.Y(wire234_0_2));
NANDC2x1 inst_and_b234_0_3 (.A(A6),.B(A7),.Y(imd_wire234_0_3));
INVC inst_inv_b234_0_3 (.A(imd_wire234_0_3),.Y(wire234_0_3));
NANDC2x1 inst_and_b234_1_0 (.A(wire234_0_0),.B(wire234_0_1),.Y(imd_wire234_1_0));
INVC inst_inv_b234_1_0 (.A(imd_wire234_1_0),.Y(wire234_1_0));
NANDC2x1 inst_and_b234_1_1 (.A(wire234_0_2),.B(wire234_0_3),.Y(imd_wire234_1_1));
INVC inst_inv_b234_1_1 (.A(imd_wire234_1_1),.Y(wire234_1_1));
NANDC2x1 inst_and_b234_2_0 (.A(wire234_1_0),.B(wire234_1_1),.Y(imd_Y234));
INVC inst_inv_b234_2_0 (.A(imd_Y234),.Y(Y234));
NANDC2x1 inst_clockedAND_b234_234 (.A(CLK),.B(Y234),.Y(imd_YF234));
INVC inst_clockedinv_b234_234 (.A(imd_YF234),.Y(YF234));


NANDC2x1 inst_and_b235_0_0 (.A(A0),.B(A1),.Y(imd_wire235_0_0));
INVC inst_inv_b235_0_0 (.A(imd_wire235_0_0),.Y(wire235_0_0));
NANDC2x1 inst_and_b235_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire235_0_1));
INVC inst_inv_b235_0_1 (.A(imd_wire235_0_1),.Y(wire235_0_1));
NANDC2x1 inst_and_b235_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire235_0_2));
INVC inst_inv_b235_0_2 (.A(imd_wire235_0_2),.Y(wire235_0_2));
NANDC2x1 inst_and_b235_0_3 (.A(A6),.B(A7),.Y(imd_wire235_0_3));
INVC inst_inv_b235_0_3 (.A(imd_wire235_0_3),.Y(wire235_0_3));
NANDC2x1 inst_and_b235_1_0 (.A(wire235_0_0),.B(wire235_0_1),.Y(imd_wire235_1_0));
INVC inst_inv_b235_1_0 (.A(imd_wire235_1_0),.Y(wire235_1_0));
NANDC2x1 inst_and_b235_1_1 (.A(wire235_0_2),.B(wire235_0_3),.Y(imd_wire235_1_1));
INVC inst_inv_b235_1_1 (.A(imd_wire235_1_1),.Y(wire235_1_1));
NANDC2x1 inst_and_b235_2_0 (.A(wire235_1_0),.B(wire235_1_1),.Y(imd_Y235));
INVC inst_inv_b235_2_0 (.A(imd_Y235),.Y(Y235));
NANDC2x1 inst_clockedAND_b235_235 (.A(CLK),.B(Y235),.Y(imd_YF235));
INVC inst_clockedinv_b235_235 (.A(imd_YF235),.Y(YF235));


NANDC2x1 inst_and_b236_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire236_0_0));
INVC inst_inv_b236_0_0 (.A(imd_wire236_0_0),.Y(wire236_0_0));
NANDC2x1 inst_and_b236_0_1 (.A(A2),.B(A3),.Y(imd_wire236_0_1));
INVC inst_inv_b236_0_1 (.A(imd_wire236_0_1),.Y(wire236_0_1));
NANDC2x1 inst_and_b236_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire236_0_2));
INVC inst_inv_b236_0_2 (.A(imd_wire236_0_2),.Y(wire236_0_2));
NANDC2x1 inst_and_b236_0_3 (.A(A6),.B(A7),.Y(imd_wire236_0_3));
INVC inst_inv_b236_0_3 (.A(imd_wire236_0_3),.Y(wire236_0_3));
NANDC2x1 inst_and_b236_1_0 (.A(wire236_0_0),.B(wire236_0_1),.Y(imd_wire236_1_0));
INVC inst_inv_b236_1_0 (.A(imd_wire236_1_0),.Y(wire236_1_0));
NANDC2x1 inst_and_b236_1_1 (.A(wire236_0_2),.B(wire236_0_3),.Y(imd_wire236_1_1));
INVC inst_inv_b236_1_1 (.A(imd_wire236_1_1),.Y(wire236_1_1));
NANDC2x1 inst_and_b236_2_0 (.A(wire236_1_0),.B(wire236_1_1),.Y(imd_Y236));
INVC inst_inv_b236_2_0 (.A(imd_Y236),.Y(Y236));
NANDC2x1 inst_clockedAND_b236_236 (.A(CLK),.B(Y236),.Y(imd_YF236));
INVC inst_clockedinv_b236_236 (.A(imd_YF236),.Y(YF236));


NANDC2x1 inst_and_b237_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire237_0_0));
INVC inst_inv_b237_0_0 (.A(imd_wire237_0_0),.Y(wire237_0_0));
NANDC2x1 inst_and_b237_0_1 (.A(A2),.B(A3),.Y(imd_wire237_0_1));
INVC inst_inv_b237_0_1 (.A(imd_wire237_0_1),.Y(wire237_0_1));
NANDC2x1 inst_and_b237_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire237_0_2));
INVC inst_inv_b237_0_2 (.A(imd_wire237_0_2),.Y(wire237_0_2));
NANDC2x1 inst_and_b237_0_3 (.A(A6),.B(A7),.Y(imd_wire237_0_3));
INVC inst_inv_b237_0_3 (.A(imd_wire237_0_3),.Y(wire237_0_3));
NANDC2x1 inst_and_b237_1_0 (.A(wire237_0_0),.B(wire237_0_1),.Y(imd_wire237_1_0));
INVC inst_inv_b237_1_0 (.A(imd_wire237_1_0),.Y(wire237_1_0));
NANDC2x1 inst_and_b237_1_1 (.A(wire237_0_2),.B(wire237_0_3),.Y(imd_wire237_1_1));
INVC inst_inv_b237_1_1 (.A(imd_wire237_1_1),.Y(wire237_1_1));
NANDC2x1 inst_and_b237_2_0 (.A(wire237_1_0),.B(wire237_1_1),.Y(imd_Y237));
INVC inst_inv_b237_2_0 (.A(imd_Y237),.Y(Y237));
NANDC2x1 inst_clockedAND_b237_237 (.A(CLK),.B(Y237),.Y(imd_YF237));
INVC inst_clockedinv_b237_237 (.A(imd_YF237),.Y(YF237));


NANDC2x1 inst_and_b238_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire238_0_0));
INVC inst_inv_b238_0_0 (.A(imd_wire238_0_0),.Y(wire238_0_0));
NANDC2x1 inst_and_b238_0_1 (.A(A2),.B(A3),.Y(imd_wire238_0_1));
INVC inst_inv_b238_0_1 (.A(imd_wire238_0_1),.Y(wire238_0_1));
NANDC2x1 inst_and_b238_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire238_0_2));
INVC inst_inv_b238_0_2 (.A(imd_wire238_0_2),.Y(wire238_0_2));
NANDC2x1 inst_and_b238_0_3 (.A(A6),.B(A7),.Y(imd_wire238_0_3));
INVC inst_inv_b238_0_3 (.A(imd_wire238_0_3),.Y(wire238_0_3));
NANDC2x1 inst_and_b238_1_0 (.A(wire238_0_0),.B(wire238_0_1),.Y(imd_wire238_1_0));
INVC inst_inv_b238_1_0 (.A(imd_wire238_1_0),.Y(wire238_1_0));
NANDC2x1 inst_and_b238_1_1 (.A(wire238_0_2),.B(wire238_0_3),.Y(imd_wire238_1_1));
INVC inst_inv_b238_1_1 (.A(imd_wire238_1_1),.Y(wire238_1_1));
NANDC2x1 inst_and_b238_2_0 (.A(wire238_1_0),.B(wire238_1_1),.Y(imd_Y238));
INVC inst_inv_b238_2_0 (.A(imd_Y238),.Y(Y238));
NANDC2x1 inst_clockedAND_b238_238 (.A(CLK),.B(Y238),.Y(imd_YF238));
INVC inst_clockedinv_b238_238 (.A(imd_YF238),.Y(YF238));


NANDC2x1 inst_and_b239_0_0 (.A(A0),.B(A1),.Y(imd_wire239_0_0));
INVC inst_inv_b239_0_0 (.A(imd_wire239_0_0),.Y(wire239_0_0));
NANDC2x1 inst_and_b239_0_1 (.A(A2),.B(A3),.Y(imd_wire239_0_1));
INVC inst_inv_b239_0_1 (.A(imd_wire239_0_1),.Y(wire239_0_1));
NANDC2x1 inst_and_b239_0_2 (.A(A4_inv),.B(A5),.Y(imd_wire239_0_2));
INVC inst_inv_b239_0_2 (.A(imd_wire239_0_2),.Y(wire239_0_2));
NANDC2x1 inst_and_b239_0_3 (.A(A6),.B(A7),.Y(imd_wire239_0_3));
INVC inst_inv_b239_0_3 (.A(imd_wire239_0_3),.Y(wire239_0_3));
NANDC2x1 inst_and_b239_1_0 (.A(wire239_0_0),.B(wire239_0_1),.Y(imd_wire239_1_0));
INVC inst_inv_b239_1_0 (.A(imd_wire239_1_0),.Y(wire239_1_0));
NANDC2x1 inst_and_b239_1_1 (.A(wire239_0_2),.B(wire239_0_3),.Y(imd_wire239_1_1));
INVC inst_inv_b239_1_1 (.A(imd_wire239_1_1),.Y(wire239_1_1));
NANDC2x1 inst_and_b239_2_0 (.A(wire239_1_0),.B(wire239_1_1),.Y(imd_Y239));
INVC inst_inv_b239_2_0 (.A(imd_Y239),.Y(Y239));
NANDC2x1 inst_clockedAND_b239_239 (.A(CLK),.B(Y239),.Y(imd_YF239));
INVC inst_clockedinv_b239_239 (.A(imd_YF239),.Y(YF239));


NANDC2x1 inst_and_b240_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire240_0_0));
INVC inst_inv_b240_0_0 (.A(imd_wire240_0_0),.Y(wire240_0_0));
NANDC2x1 inst_and_b240_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire240_0_1));
INVC inst_inv_b240_0_1 (.A(imd_wire240_0_1),.Y(wire240_0_1));
NANDC2x1 inst_and_b240_0_2 (.A(A4),.B(A5),.Y(imd_wire240_0_2));
INVC inst_inv_b240_0_2 (.A(imd_wire240_0_2),.Y(wire240_0_2));
NANDC2x1 inst_and_b240_0_3 (.A(A6),.B(A7),.Y(imd_wire240_0_3));
INVC inst_inv_b240_0_3 (.A(imd_wire240_0_3),.Y(wire240_0_3));
NANDC2x1 inst_and_b240_1_0 (.A(wire240_0_0),.B(wire240_0_1),.Y(imd_wire240_1_0));
INVC inst_inv_b240_1_0 (.A(imd_wire240_1_0),.Y(wire240_1_0));
NANDC2x1 inst_and_b240_1_1 (.A(wire240_0_2),.B(wire240_0_3),.Y(imd_wire240_1_1));
INVC inst_inv_b240_1_1 (.A(imd_wire240_1_1),.Y(wire240_1_1));
NANDC2x1 inst_and_b240_2_0 (.A(wire240_1_0),.B(wire240_1_1),.Y(imd_Y240));
INVC inst_inv_b240_2_0 (.A(imd_Y240),.Y(Y240));
NANDC2x1 inst_clockedAND_b240_240 (.A(CLK),.B(Y240),.Y(imd_YF240));
INVC inst_clockedinv_b240_240 (.A(imd_YF240),.Y(YF240));


NANDC2x1 inst_and_b241_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire241_0_0));
INVC inst_inv_b241_0_0 (.A(imd_wire241_0_0),.Y(wire241_0_0));
NANDC2x1 inst_and_b241_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire241_0_1));
INVC inst_inv_b241_0_1 (.A(imd_wire241_0_1),.Y(wire241_0_1));
NANDC2x1 inst_and_b241_0_2 (.A(A4),.B(A5),.Y(imd_wire241_0_2));
INVC inst_inv_b241_0_2 (.A(imd_wire241_0_2),.Y(wire241_0_2));
NANDC2x1 inst_and_b241_0_3 (.A(A6),.B(A7),.Y(imd_wire241_0_3));
INVC inst_inv_b241_0_3 (.A(imd_wire241_0_3),.Y(wire241_0_3));
NANDC2x1 inst_and_b241_1_0 (.A(wire241_0_0),.B(wire241_0_1),.Y(imd_wire241_1_0));
INVC inst_inv_b241_1_0 (.A(imd_wire241_1_0),.Y(wire241_1_0));
NANDC2x1 inst_and_b241_1_1 (.A(wire241_0_2),.B(wire241_0_3),.Y(imd_wire241_1_1));
INVC inst_inv_b241_1_1 (.A(imd_wire241_1_1),.Y(wire241_1_1));
NANDC2x1 inst_and_b241_2_0 (.A(wire241_1_0),.B(wire241_1_1),.Y(imd_Y241));
INVC inst_inv_b241_2_0 (.A(imd_Y241),.Y(Y241));
NANDC2x1 inst_clockedAND_b241_241 (.A(CLK),.B(Y241),.Y(imd_YF241));
INVC inst_clockedinv_b241_241 (.A(imd_YF241),.Y(YF241));


NANDC2x1 inst_and_b242_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire242_0_0));
INVC inst_inv_b242_0_0 (.A(imd_wire242_0_0),.Y(wire242_0_0));
NANDC2x1 inst_and_b242_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire242_0_1));
INVC inst_inv_b242_0_1 (.A(imd_wire242_0_1),.Y(wire242_0_1));
NANDC2x1 inst_and_b242_0_2 (.A(A4),.B(A5),.Y(imd_wire242_0_2));
INVC inst_inv_b242_0_2 (.A(imd_wire242_0_2),.Y(wire242_0_2));
NANDC2x1 inst_and_b242_0_3 (.A(A6),.B(A7),.Y(imd_wire242_0_3));
INVC inst_inv_b242_0_3 (.A(imd_wire242_0_3),.Y(wire242_0_3));
NANDC2x1 inst_and_b242_1_0 (.A(wire242_0_0),.B(wire242_0_1),.Y(imd_wire242_1_0));
INVC inst_inv_b242_1_0 (.A(imd_wire242_1_0),.Y(wire242_1_0));
NANDC2x1 inst_and_b242_1_1 (.A(wire242_0_2),.B(wire242_0_3),.Y(imd_wire242_1_1));
INVC inst_inv_b242_1_1 (.A(imd_wire242_1_1),.Y(wire242_1_1));
NANDC2x1 inst_and_b242_2_0 (.A(wire242_1_0),.B(wire242_1_1),.Y(imd_Y242));
INVC inst_inv_b242_2_0 (.A(imd_Y242),.Y(Y242));
NANDC2x1 inst_clockedAND_b242_242 (.A(CLK),.B(Y242),.Y(imd_YF242));
INVC inst_clockedinv_b242_242 (.A(imd_YF242),.Y(YF242));


NANDC2x1 inst_and_b243_0_0 (.A(A0),.B(A1),.Y(imd_wire243_0_0));
INVC inst_inv_b243_0_0 (.A(imd_wire243_0_0),.Y(wire243_0_0));
NANDC2x1 inst_and_b243_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire243_0_1));
INVC inst_inv_b243_0_1 (.A(imd_wire243_0_1),.Y(wire243_0_1));
NANDC2x1 inst_and_b243_0_2 (.A(A4),.B(A5),.Y(imd_wire243_0_2));
INVC inst_inv_b243_0_2 (.A(imd_wire243_0_2),.Y(wire243_0_2));
NANDC2x1 inst_and_b243_0_3 (.A(A6),.B(A7),.Y(imd_wire243_0_3));
INVC inst_inv_b243_0_3 (.A(imd_wire243_0_3),.Y(wire243_0_3));
NANDC2x1 inst_and_b243_1_0 (.A(wire243_0_0),.B(wire243_0_1),.Y(imd_wire243_1_0));
INVC inst_inv_b243_1_0 (.A(imd_wire243_1_0),.Y(wire243_1_0));
NANDC2x1 inst_and_b243_1_1 (.A(wire243_0_2),.B(wire243_0_3),.Y(imd_wire243_1_1));
INVC inst_inv_b243_1_1 (.A(imd_wire243_1_1),.Y(wire243_1_1));
NANDC2x1 inst_and_b243_2_0 (.A(wire243_1_0),.B(wire243_1_1),.Y(imd_Y243));
INVC inst_inv_b243_2_0 (.A(imd_Y243),.Y(Y243));
NANDC2x1 inst_clockedAND_b243_243 (.A(CLK),.B(Y243),.Y(imd_YF243));
INVC inst_clockedinv_b243_243 (.A(imd_YF243),.Y(YF243));


NANDC2x1 inst_and_b244_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire244_0_0));
INVC inst_inv_b244_0_0 (.A(imd_wire244_0_0),.Y(wire244_0_0));
NANDC2x1 inst_and_b244_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire244_0_1));
INVC inst_inv_b244_0_1 (.A(imd_wire244_0_1),.Y(wire244_0_1));
NANDC2x1 inst_and_b244_0_2 (.A(A4),.B(A5),.Y(imd_wire244_0_2));
INVC inst_inv_b244_0_2 (.A(imd_wire244_0_2),.Y(wire244_0_2));
NANDC2x1 inst_and_b244_0_3 (.A(A6),.B(A7),.Y(imd_wire244_0_3));
INVC inst_inv_b244_0_3 (.A(imd_wire244_0_3),.Y(wire244_0_3));
NANDC2x1 inst_and_b244_1_0 (.A(wire244_0_0),.B(wire244_0_1),.Y(imd_wire244_1_0));
INVC inst_inv_b244_1_0 (.A(imd_wire244_1_0),.Y(wire244_1_0));
NANDC2x1 inst_and_b244_1_1 (.A(wire244_0_2),.B(wire244_0_3),.Y(imd_wire244_1_1));
INVC inst_inv_b244_1_1 (.A(imd_wire244_1_1),.Y(wire244_1_1));
NANDC2x1 inst_and_b244_2_0 (.A(wire244_1_0),.B(wire244_1_1),.Y(imd_Y244));
INVC inst_inv_b244_2_0 (.A(imd_Y244),.Y(Y244));
NANDC2x1 inst_clockedAND_b244_244 (.A(CLK),.B(Y244),.Y(imd_YF244));
INVC inst_clockedinv_b244_244 (.A(imd_YF244),.Y(YF244));


NANDC2x1 inst_and_b245_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire245_0_0));
INVC inst_inv_b245_0_0 (.A(imd_wire245_0_0),.Y(wire245_0_0));
NANDC2x1 inst_and_b245_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire245_0_1));
INVC inst_inv_b245_0_1 (.A(imd_wire245_0_1),.Y(wire245_0_1));
NANDC2x1 inst_and_b245_0_2 (.A(A4),.B(A5),.Y(imd_wire245_0_2));
INVC inst_inv_b245_0_2 (.A(imd_wire245_0_2),.Y(wire245_0_2));
NANDC2x1 inst_and_b245_0_3 (.A(A6),.B(A7),.Y(imd_wire245_0_3));
INVC inst_inv_b245_0_3 (.A(imd_wire245_0_3),.Y(wire245_0_3));
NANDC2x1 inst_and_b245_1_0 (.A(wire245_0_0),.B(wire245_0_1),.Y(imd_wire245_1_0));
INVC inst_inv_b245_1_0 (.A(imd_wire245_1_0),.Y(wire245_1_0));
NANDC2x1 inst_and_b245_1_1 (.A(wire245_0_2),.B(wire245_0_3),.Y(imd_wire245_1_1));
INVC inst_inv_b245_1_1 (.A(imd_wire245_1_1),.Y(wire245_1_1));
NANDC2x1 inst_and_b245_2_0 (.A(wire245_1_0),.B(wire245_1_1),.Y(imd_Y245));
INVC inst_inv_b245_2_0 (.A(imd_Y245),.Y(Y245));
NANDC2x1 inst_clockedAND_b245_245 (.A(CLK),.B(Y245),.Y(imd_YF245));
INVC inst_clockedinv_b245_245 (.A(imd_YF245),.Y(YF245));


NANDC2x1 inst_and_b246_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire246_0_0));
INVC inst_inv_b246_0_0 (.A(imd_wire246_0_0),.Y(wire246_0_0));
NANDC2x1 inst_and_b246_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire246_0_1));
INVC inst_inv_b246_0_1 (.A(imd_wire246_0_1),.Y(wire246_0_1));
NANDC2x1 inst_and_b246_0_2 (.A(A4),.B(A5),.Y(imd_wire246_0_2));
INVC inst_inv_b246_0_2 (.A(imd_wire246_0_2),.Y(wire246_0_2));
NANDC2x1 inst_and_b246_0_3 (.A(A6),.B(A7),.Y(imd_wire246_0_3));
INVC inst_inv_b246_0_3 (.A(imd_wire246_0_3),.Y(wire246_0_3));
NANDC2x1 inst_and_b246_1_0 (.A(wire246_0_0),.B(wire246_0_1),.Y(imd_wire246_1_0));
INVC inst_inv_b246_1_0 (.A(imd_wire246_1_0),.Y(wire246_1_0));
NANDC2x1 inst_and_b246_1_1 (.A(wire246_0_2),.B(wire246_0_3),.Y(imd_wire246_1_1));
INVC inst_inv_b246_1_1 (.A(imd_wire246_1_1),.Y(wire246_1_1));
NANDC2x1 inst_and_b246_2_0 (.A(wire246_1_0),.B(wire246_1_1),.Y(imd_Y246));
INVC inst_inv_b246_2_0 (.A(imd_Y246),.Y(Y246));
NANDC2x1 inst_clockedAND_b246_246 (.A(CLK),.B(Y246),.Y(imd_YF246));
INVC inst_clockedinv_b246_246 (.A(imd_YF246),.Y(YF246));


NANDC2x1 inst_and_b247_0_0 (.A(A0),.B(A1),.Y(imd_wire247_0_0));
INVC inst_inv_b247_0_0 (.A(imd_wire247_0_0),.Y(wire247_0_0));
NANDC2x1 inst_and_b247_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire247_0_1));
INVC inst_inv_b247_0_1 (.A(imd_wire247_0_1),.Y(wire247_0_1));
NANDC2x1 inst_and_b247_0_2 (.A(A4),.B(A5),.Y(imd_wire247_0_2));
INVC inst_inv_b247_0_2 (.A(imd_wire247_0_2),.Y(wire247_0_2));
NANDC2x1 inst_and_b247_0_3 (.A(A6),.B(A7),.Y(imd_wire247_0_3));
INVC inst_inv_b247_0_3 (.A(imd_wire247_0_3),.Y(wire247_0_3));
NANDC2x1 inst_and_b247_1_0 (.A(wire247_0_0),.B(wire247_0_1),.Y(imd_wire247_1_0));
INVC inst_inv_b247_1_0 (.A(imd_wire247_1_0),.Y(wire247_1_0));
NANDC2x1 inst_and_b247_1_1 (.A(wire247_0_2),.B(wire247_0_3),.Y(imd_wire247_1_1));
INVC inst_inv_b247_1_1 (.A(imd_wire247_1_1),.Y(wire247_1_1));
NANDC2x1 inst_and_b247_2_0 (.A(wire247_1_0),.B(wire247_1_1),.Y(imd_Y247));
INVC inst_inv_b247_2_0 (.A(imd_Y247),.Y(Y247));
NANDC2x1 inst_clockedAND_b247_247 (.A(CLK),.B(Y247),.Y(imd_YF247));
INVC inst_clockedinv_b247_247 (.A(imd_YF247),.Y(YF247));


NANDC2x1 inst_and_b248_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire248_0_0));
INVC inst_inv_b248_0_0 (.A(imd_wire248_0_0),.Y(wire248_0_0));
NANDC2x1 inst_and_b248_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire248_0_1));
INVC inst_inv_b248_0_1 (.A(imd_wire248_0_1),.Y(wire248_0_1));
NANDC2x1 inst_and_b248_0_2 (.A(A4),.B(A5),.Y(imd_wire248_0_2));
INVC inst_inv_b248_0_2 (.A(imd_wire248_0_2),.Y(wire248_0_2));
NANDC2x1 inst_and_b248_0_3 (.A(A6),.B(A7),.Y(imd_wire248_0_3));
INVC inst_inv_b248_0_3 (.A(imd_wire248_0_3),.Y(wire248_0_3));
NANDC2x1 inst_and_b248_1_0 (.A(wire248_0_0),.B(wire248_0_1),.Y(imd_wire248_1_0));
INVC inst_inv_b248_1_0 (.A(imd_wire248_1_0),.Y(wire248_1_0));
NANDC2x1 inst_and_b248_1_1 (.A(wire248_0_2),.B(wire248_0_3),.Y(imd_wire248_1_1));
INVC inst_inv_b248_1_1 (.A(imd_wire248_1_1),.Y(wire248_1_1));
NANDC2x1 inst_and_b248_2_0 (.A(wire248_1_0),.B(wire248_1_1),.Y(imd_Y248));
INVC inst_inv_b248_2_0 (.A(imd_Y248),.Y(Y248));
NANDC2x1 inst_clockedAND_b248_248 (.A(CLK),.B(Y248),.Y(imd_YF248));
INVC inst_clockedinv_b248_248 (.A(imd_YF248),.Y(YF248));


NANDC2x1 inst_and_b249_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire249_0_0));
INVC inst_inv_b249_0_0 (.A(imd_wire249_0_0),.Y(wire249_0_0));
NANDC2x1 inst_and_b249_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire249_0_1));
INVC inst_inv_b249_0_1 (.A(imd_wire249_0_1),.Y(wire249_0_1));
NANDC2x1 inst_and_b249_0_2 (.A(A4),.B(A5),.Y(imd_wire249_0_2));
INVC inst_inv_b249_0_2 (.A(imd_wire249_0_2),.Y(wire249_0_2));
NANDC2x1 inst_and_b249_0_3 (.A(A6),.B(A7),.Y(imd_wire249_0_3));
INVC inst_inv_b249_0_3 (.A(imd_wire249_0_3),.Y(wire249_0_3));
NANDC2x1 inst_and_b249_1_0 (.A(wire249_0_0),.B(wire249_0_1),.Y(imd_wire249_1_0));
INVC inst_inv_b249_1_0 (.A(imd_wire249_1_0),.Y(wire249_1_0));
NANDC2x1 inst_and_b249_1_1 (.A(wire249_0_2),.B(wire249_0_3),.Y(imd_wire249_1_1));
INVC inst_inv_b249_1_1 (.A(imd_wire249_1_1),.Y(wire249_1_1));
NANDC2x1 inst_and_b249_2_0 (.A(wire249_1_0),.B(wire249_1_1),.Y(imd_Y249));
INVC inst_inv_b249_2_0 (.A(imd_Y249),.Y(Y249));
NANDC2x1 inst_clockedAND_b249_249 (.A(CLK),.B(Y249),.Y(imd_YF249));
INVC inst_clockedinv_b249_249 (.A(imd_YF249),.Y(YF249));


NANDC2x1 inst_and_b250_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire250_0_0));
INVC inst_inv_b250_0_0 (.A(imd_wire250_0_0),.Y(wire250_0_0));
NANDC2x1 inst_and_b250_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire250_0_1));
INVC inst_inv_b250_0_1 (.A(imd_wire250_0_1),.Y(wire250_0_1));
NANDC2x1 inst_and_b250_0_2 (.A(A4),.B(A5),.Y(imd_wire250_0_2));
INVC inst_inv_b250_0_2 (.A(imd_wire250_0_2),.Y(wire250_0_2));
NANDC2x1 inst_and_b250_0_3 (.A(A6),.B(A7),.Y(imd_wire250_0_3));
INVC inst_inv_b250_0_3 (.A(imd_wire250_0_3),.Y(wire250_0_3));
NANDC2x1 inst_and_b250_1_0 (.A(wire250_0_0),.B(wire250_0_1),.Y(imd_wire250_1_0));
INVC inst_inv_b250_1_0 (.A(imd_wire250_1_0),.Y(wire250_1_0));
NANDC2x1 inst_and_b250_1_1 (.A(wire250_0_2),.B(wire250_0_3),.Y(imd_wire250_1_1));
INVC inst_inv_b250_1_1 (.A(imd_wire250_1_1),.Y(wire250_1_1));
NANDC2x1 inst_and_b250_2_0 (.A(wire250_1_0),.B(wire250_1_1),.Y(imd_Y250));
INVC inst_inv_b250_2_0 (.A(imd_Y250),.Y(Y250));
NANDC2x1 inst_clockedAND_b250_250 (.A(CLK),.B(Y250),.Y(imd_YF250));
INVC inst_clockedinv_b250_250 (.A(imd_YF250),.Y(YF250));


NANDC2x1 inst_and_b251_0_0 (.A(A0),.B(A1),.Y(imd_wire251_0_0));
INVC inst_inv_b251_0_0 (.A(imd_wire251_0_0),.Y(wire251_0_0));
NANDC2x1 inst_and_b251_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire251_0_1));
INVC inst_inv_b251_0_1 (.A(imd_wire251_0_1),.Y(wire251_0_1));
NANDC2x1 inst_and_b251_0_2 (.A(A4),.B(A5),.Y(imd_wire251_0_2));
INVC inst_inv_b251_0_2 (.A(imd_wire251_0_2),.Y(wire251_0_2));
NANDC2x1 inst_and_b251_0_3 (.A(A6),.B(A7),.Y(imd_wire251_0_3));
INVC inst_inv_b251_0_3 (.A(imd_wire251_0_3),.Y(wire251_0_3));
NANDC2x1 inst_and_b251_1_0 (.A(wire251_0_0),.B(wire251_0_1),.Y(imd_wire251_1_0));
INVC inst_inv_b251_1_0 (.A(imd_wire251_1_0),.Y(wire251_1_0));
NANDC2x1 inst_and_b251_1_1 (.A(wire251_0_2),.B(wire251_0_3),.Y(imd_wire251_1_1));
INVC inst_inv_b251_1_1 (.A(imd_wire251_1_1),.Y(wire251_1_1));
NANDC2x1 inst_and_b251_2_0 (.A(wire251_1_0),.B(wire251_1_1),.Y(imd_Y251));
INVC inst_inv_b251_2_0 (.A(imd_Y251),.Y(Y251));
NANDC2x1 inst_clockedAND_b251_251 (.A(CLK),.B(Y251),.Y(imd_YF251));
INVC inst_clockedinv_b251_251 (.A(imd_YF251),.Y(YF251));


NANDC2x1 inst_and_b252_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire252_0_0));
INVC inst_inv_b252_0_0 (.A(imd_wire252_0_0),.Y(wire252_0_0));
NANDC2x1 inst_and_b252_0_1 (.A(A2),.B(A3),.Y(imd_wire252_0_1));
INVC inst_inv_b252_0_1 (.A(imd_wire252_0_1),.Y(wire252_0_1));
NANDC2x1 inst_and_b252_0_2 (.A(A4),.B(A5),.Y(imd_wire252_0_2));
INVC inst_inv_b252_0_2 (.A(imd_wire252_0_2),.Y(wire252_0_2));
NANDC2x1 inst_and_b252_0_3 (.A(A6),.B(A7),.Y(imd_wire252_0_3));
INVC inst_inv_b252_0_3 (.A(imd_wire252_0_3),.Y(wire252_0_3));
NANDC2x1 inst_and_b252_1_0 (.A(wire252_0_0),.B(wire252_0_1),.Y(imd_wire252_1_0));
INVC inst_inv_b252_1_0 (.A(imd_wire252_1_0),.Y(wire252_1_0));
NANDC2x1 inst_and_b252_1_1 (.A(wire252_0_2),.B(wire252_0_3),.Y(imd_wire252_1_1));
INVC inst_inv_b252_1_1 (.A(imd_wire252_1_1),.Y(wire252_1_1));
NANDC2x1 inst_and_b252_2_0 (.A(wire252_1_0),.B(wire252_1_1),.Y(imd_Y252));
INVC inst_inv_b252_2_0 (.A(imd_Y252),.Y(Y252));
NANDC2x1 inst_clockedAND_b252_252 (.A(CLK),.B(Y252),.Y(imd_YF252));
INVC inst_clockedinv_b252_252 (.A(imd_YF252),.Y(YF252));


NANDC2x1 inst_and_b253_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire253_0_0));
INVC inst_inv_b253_0_0 (.A(imd_wire253_0_0),.Y(wire253_0_0));
NANDC2x1 inst_and_b253_0_1 (.A(A2),.B(A3),.Y(imd_wire253_0_1));
INVC inst_inv_b253_0_1 (.A(imd_wire253_0_1),.Y(wire253_0_1));
NANDC2x1 inst_and_b253_0_2 (.A(A4),.B(A5),.Y(imd_wire253_0_2));
INVC inst_inv_b253_0_2 (.A(imd_wire253_0_2),.Y(wire253_0_2));
NANDC2x1 inst_and_b253_0_3 (.A(A6),.B(A7),.Y(imd_wire253_0_3));
INVC inst_inv_b253_0_3 (.A(imd_wire253_0_3),.Y(wire253_0_3));
NANDC2x1 inst_and_b253_1_0 (.A(wire253_0_0),.B(wire253_0_1),.Y(imd_wire253_1_0));
INVC inst_inv_b253_1_0 (.A(imd_wire253_1_0),.Y(wire253_1_0));
NANDC2x1 inst_and_b253_1_1 (.A(wire253_0_2),.B(wire253_0_3),.Y(imd_wire253_1_1));
INVC inst_inv_b253_1_1 (.A(imd_wire253_1_1),.Y(wire253_1_1));
NANDC2x1 inst_and_b253_2_0 (.A(wire253_1_0),.B(wire253_1_1),.Y(imd_Y253));
INVC inst_inv_b253_2_0 (.A(imd_Y253),.Y(Y253));
NANDC2x1 inst_clockedAND_b253_253 (.A(CLK),.B(Y253),.Y(imd_YF253));
INVC inst_clockedinv_b253_253 (.A(imd_YF253),.Y(YF253));


NANDC2x1 inst_and_b254_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire254_0_0));
INVC inst_inv_b254_0_0 (.A(imd_wire254_0_0),.Y(wire254_0_0));
NANDC2x1 inst_and_b254_0_1 (.A(A2),.B(A3),.Y(imd_wire254_0_1));
INVC inst_inv_b254_0_1 (.A(imd_wire254_0_1),.Y(wire254_0_1));
NANDC2x1 inst_and_b254_0_2 (.A(A4),.B(A5),.Y(imd_wire254_0_2));
INVC inst_inv_b254_0_2 (.A(imd_wire254_0_2),.Y(wire254_0_2));
NANDC2x1 inst_and_b254_0_3 (.A(A6),.B(A7),.Y(imd_wire254_0_3));
INVC inst_inv_b254_0_3 (.A(imd_wire254_0_3),.Y(wire254_0_3));
NANDC2x1 inst_and_b254_1_0 (.A(wire254_0_0),.B(wire254_0_1),.Y(imd_wire254_1_0));
INVC inst_inv_b254_1_0 (.A(imd_wire254_1_0),.Y(wire254_1_0));
NANDC2x1 inst_and_b254_1_1 (.A(wire254_0_2),.B(wire254_0_3),.Y(imd_wire254_1_1));
INVC inst_inv_b254_1_1 (.A(imd_wire254_1_1),.Y(wire254_1_1));
NANDC2x1 inst_and_b254_2_0 (.A(wire254_1_0),.B(wire254_1_1),.Y(imd_Y254));
INVC inst_inv_b254_2_0 (.A(imd_Y254),.Y(Y254));
NANDC2x1 inst_clockedAND_b254_254 (.A(CLK),.B(Y254),.Y(imd_YF254));
INVC inst_clockedinv_b254_254 (.A(imd_YF254),.Y(YF254));


NANDC2x1 inst_and_b255_0_0 (.A(A0),.B(A1),.Y(imd_wire255_0_0));
INVC inst_inv_b255_0_0 (.A(imd_wire255_0_0),.Y(wire255_0_0));
NANDC2x1 inst_and_b255_0_1 (.A(A2),.B(A3),.Y(imd_wire255_0_1));
INVC inst_inv_b255_0_1 (.A(imd_wire255_0_1),.Y(wire255_0_1));
NANDC2x1 inst_and_b255_0_2 (.A(A4),.B(A5),.Y(imd_wire255_0_2));
INVC inst_inv_b255_0_2 (.A(imd_wire255_0_2),.Y(wire255_0_2));
NANDC2x1 inst_and_b255_0_3 (.A(A6),.B(A7),.Y(imd_wire255_0_3));
INVC inst_inv_b255_0_3 (.A(imd_wire255_0_3),.Y(wire255_0_3));
NANDC2x1 inst_and_b255_1_0 (.A(wire255_0_0),.B(wire255_0_1),.Y(imd_wire255_1_0));
INVC inst_inv_b255_1_0 (.A(imd_wire255_1_0),.Y(wire255_1_0));
NANDC2x1 inst_and_b255_1_1 (.A(wire255_0_2),.B(wire255_0_3),.Y(imd_wire255_1_1));
INVC inst_inv_b255_1_1 (.A(imd_wire255_1_1),.Y(wire255_1_1));
NANDC2x1 inst_and_b255_2_0 (.A(wire255_1_0),.B(wire255_1_1),.Y(imd_Y255));
INVC inst_inv_b255_2_0 (.A(imd_Y255),.Y(Y255));
NANDC2x1 inst_clockedAND_b255_255 (.A(CLK),.B(Y255),.Y(imd_YF255));
INVC inst_clockedinv_b255_255 (.A(imd_YF255),.Y(YF255));


endmodule
module colDecoder(A0,A0_inv,A1,A1_inv,A2,A2_inv,A3,A3_inv,CLK,YF0,YF1,YF2,YF3,YF4,YF5,YF6,YF7,YF8,YF9,YF10,YF11,YF12,YF13,YF14,YF15);
input A0;
input A0_inv;
input A1;
input A1_inv;
input A2;
input A2_inv;
input A3;
input A3_inv;
input CLK;
output YF0;
output YF1;
output YF2;
output YF3;
output YF4;
output YF5;
output YF6;
output YF7;
output YF8;
output YF9;
output YF10;
output YF11;
output YF12;
output YF13;
output YF14;
output YF15;
NANDC2x1 inst_and_b0_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire0_0_0));
INVC inst_inv_b0_0_0 (.A(imd_wire0_0_0),.Y(wire0_0_0));
NANDC2x1 inst_and_b0_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire0_0_1));
INVC inst_inv_b0_0_1 (.A(imd_wire0_0_1),.Y(wire0_0_1));
NANDC2x1 inst_and_b0_1_0 (.A(wire0_0_0),.B(wire0_0_1),.Y(imd_Y0));
INVC inst_inv_b0_1_0 (.A(imd_Y0),.Y(Y0));
NANDC2x1 inst_clockedAND_b0_0 (.A(CLK),.B(Y0),.Y(imd_YF0));
INVC inst_clockedinv_b0_0 (.A(imd_YF0),.Y(YF0));


NANDC2x1 inst_and_b1_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire1_0_0));
INVC inst_inv_b1_0_0 (.A(imd_wire1_0_0),.Y(wire1_0_0));
NANDC2x1 inst_and_b1_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire1_0_1));
INVC inst_inv_b1_0_1 (.A(imd_wire1_0_1),.Y(wire1_0_1));
NANDC2x1 inst_and_b1_1_0 (.A(wire1_0_0),.B(wire1_0_1),.Y(imd_Y1));
INVC inst_inv_b1_1_0 (.A(imd_Y1),.Y(Y1));
NANDC2x1 inst_clockedAND_b1_1 (.A(CLK),.B(Y1),.Y(imd_YF1));
INVC inst_clockedinv_b1_1 (.A(imd_YF1),.Y(YF1));


NANDC2x1 inst_and_b2_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire2_0_0));
INVC inst_inv_b2_0_0 (.A(imd_wire2_0_0),.Y(wire2_0_0));
NANDC2x1 inst_and_b2_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire2_0_1));
INVC inst_inv_b2_0_1 (.A(imd_wire2_0_1),.Y(wire2_0_1));
NANDC2x1 inst_and_b2_1_0 (.A(wire2_0_0),.B(wire2_0_1),.Y(imd_Y2));
INVC inst_inv_b2_1_0 (.A(imd_Y2),.Y(Y2));
NANDC2x1 inst_clockedAND_b2_2 (.A(CLK),.B(Y2),.Y(imd_YF2));
INVC inst_clockedinv_b2_2 (.A(imd_YF2),.Y(YF2));


NANDC2x1 inst_and_b3_0_0 (.A(A0),.B(A1),.Y(imd_wire3_0_0));
INVC inst_inv_b3_0_0 (.A(imd_wire3_0_0),.Y(wire3_0_0));
NANDC2x1 inst_and_b3_0_1 (.A(A2_inv),.B(A3_inv),.Y(imd_wire3_0_1));
INVC inst_inv_b3_0_1 (.A(imd_wire3_0_1),.Y(wire3_0_1));
NANDC2x1 inst_and_b3_1_0 (.A(wire3_0_0),.B(wire3_0_1),.Y(imd_Y3));
INVC inst_inv_b3_1_0 (.A(imd_Y3),.Y(Y3));
NANDC2x1 inst_clockedAND_b3_3 (.A(CLK),.B(Y3),.Y(imd_YF3));
INVC inst_clockedinv_b3_3 (.A(imd_YF3),.Y(YF3));


NANDC2x1 inst_and_b4_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire4_0_0));
INVC inst_inv_b4_0_0 (.A(imd_wire4_0_0),.Y(wire4_0_0));
NANDC2x1 inst_and_b4_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire4_0_1));
INVC inst_inv_b4_0_1 (.A(imd_wire4_0_1),.Y(wire4_0_1));
NANDC2x1 inst_and_b4_1_0 (.A(wire4_0_0),.B(wire4_0_1),.Y(imd_Y4));
INVC inst_inv_b4_1_0 (.A(imd_Y4),.Y(Y4));
NANDC2x1 inst_clockedAND_b4_4 (.A(CLK),.B(Y4),.Y(imd_YF4));
INVC inst_clockedinv_b4_4 (.A(imd_YF4),.Y(YF4));


NANDC2x1 inst_and_b5_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire5_0_0));
INVC inst_inv_b5_0_0 (.A(imd_wire5_0_0),.Y(wire5_0_0));
NANDC2x1 inst_and_b5_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire5_0_1));
INVC inst_inv_b5_0_1 (.A(imd_wire5_0_1),.Y(wire5_0_1));
NANDC2x1 inst_and_b5_1_0 (.A(wire5_0_0),.B(wire5_0_1),.Y(imd_Y5));
INVC inst_inv_b5_1_0 (.A(imd_Y5),.Y(Y5));
NANDC2x1 inst_clockedAND_b5_5 (.A(CLK),.B(Y5),.Y(imd_YF5));
INVC inst_clockedinv_b5_5 (.A(imd_YF5),.Y(YF5));


NANDC2x1 inst_and_b6_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire6_0_0));
INVC inst_inv_b6_0_0 (.A(imd_wire6_0_0),.Y(wire6_0_0));
NANDC2x1 inst_and_b6_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire6_0_1));
INVC inst_inv_b6_0_1 (.A(imd_wire6_0_1),.Y(wire6_0_1));
NANDC2x1 inst_and_b6_1_0 (.A(wire6_0_0),.B(wire6_0_1),.Y(imd_Y6));
INVC inst_inv_b6_1_0 (.A(imd_Y6),.Y(Y6));
NANDC2x1 inst_clockedAND_b6_6 (.A(CLK),.B(Y6),.Y(imd_YF6));
INVC inst_clockedinv_b6_6 (.A(imd_YF6),.Y(YF6));


NANDC2x1 inst_and_b7_0_0 (.A(A0),.B(A1),.Y(imd_wire7_0_0));
INVC inst_inv_b7_0_0 (.A(imd_wire7_0_0),.Y(wire7_0_0));
NANDC2x1 inst_and_b7_0_1 (.A(A2),.B(A3_inv),.Y(imd_wire7_0_1));
INVC inst_inv_b7_0_1 (.A(imd_wire7_0_1),.Y(wire7_0_1));
NANDC2x1 inst_and_b7_1_0 (.A(wire7_0_0),.B(wire7_0_1),.Y(imd_Y7));
INVC inst_inv_b7_1_0 (.A(imd_Y7),.Y(Y7));
NANDC2x1 inst_clockedAND_b7_7 (.A(CLK),.B(Y7),.Y(imd_YF7));
INVC inst_clockedinv_b7_7 (.A(imd_YF7),.Y(YF7));


NANDC2x1 inst_and_b8_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire8_0_0));
INVC inst_inv_b8_0_0 (.A(imd_wire8_0_0),.Y(wire8_0_0));
NANDC2x1 inst_and_b8_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire8_0_1));
INVC inst_inv_b8_0_1 (.A(imd_wire8_0_1),.Y(wire8_0_1));
NANDC2x1 inst_and_b8_1_0 (.A(wire8_0_0),.B(wire8_0_1),.Y(imd_Y8));
INVC inst_inv_b8_1_0 (.A(imd_Y8),.Y(Y8));
NANDC2x1 inst_clockedAND_b8_8 (.A(CLK),.B(Y8),.Y(imd_YF8));
INVC inst_clockedinv_b8_8 (.A(imd_YF8),.Y(YF8));


NANDC2x1 inst_and_b9_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire9_0_0));
INVC inst_inv_b9_0_0 (.A(imd_wire9_0_0),.Y(wire9_0_0));
NANDC2x1 inst_and_b9_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire9_0_1));
INVC inst_inv_b9_0_1 (.A(imd_wire9_0_1),.Y(wire9_0_1));
NANDC2x1 inst_and_b9_1_0 (.A(wire9_0_0),.B(wire9_0_1),.Y(imd_Y9));
INVC inst_inv_b9_1_0 (.A(imd_Y9),.Y(Y9));
NANDC2x1 inst_clockedAND_b9_9 (.A(CLK),.B(Y9),.Y(imd_YF9));
INVC inst_clockedinv_b9_9 (.A(imd_YF9),.Y(YF9));


NANDC2x1 inst_and_b10_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire10_0_0));
INVC inst_inv_b10_0_0 (.A(imd_wire10_0_0),.Y(wire10_0_0));
NANDC2x1 inst_and_b10_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire10_0_1));
INVC inst_inv_b10_0_1 (.A(imd_wire10_0_1),.Y(wire10_0_1));
NANDC2x1 inst_and_b10_1_0 (.A(wire10_0_0),.B(wire10_0_1),.Y(imd_Y10));
INVC inst_inv_b10_1_0 (.A(imd_Y10),.Y(Y10));
NANDC2x1 inst_clockedAND_b10_10 (.A(CLK),.B(Y10),.Y(imd_YF10));
INVC inst_clockedinv_b10_10 (.A(imd_YF10),.Y(YF10));


NANDC2x1 inst_and_b11_0_0 (.A(A0),.B(A1),.Y(imd_wire11_0_0));
INVC inst_inv_b11_0_0 (.A(imd_wire11_0_0),.Y(wire11_0_0));
NANDC2x1 inst_and_b11_0_1 (.A(A2_inv),.B(A3),.Y(imd_wire11_0_1));
INVC inst_inv_b11_0_1 (.A(imd_wire11_0_1),.Y(wire11_0_1));
NANDC2x1 inst_and_b11_1_0 (.A(wire11_0_0),.B(wire11_0_1),.Y(imd_Y11));
INVC inst_inv_b11_1_0 (.A(imd_Y11),.Y(Y11));
NANDC2x1 inst_clockedAND_b11_11 (.A(CLK),.B(Y11),.Y(imd_YF11));
INVC inst_clockedinv_b11_11 (.A(imd_YF11),.Y(YF11));


NANDC2x1 inst_and_b12_0_0 (.A(A0_inv),.B(A1_inv),.Y(imd_wire12_0_0));
INVC inst_inv_b12_0_0 (.A(imd_wire12_0_0),.Y(wire12_0_0));
NANDC2x1 inst_and_b12_0_1 (.A(A2),.B(A3),.Y(imd_wire12_0_1));
INVC inst_inv_b12_0_1 (.A(imd_wire12_0_1),.Y(wire12_0_1));
NANDC2x1 inst_and_b12_1_0 (.A(wire12_0_0),.B(wire12_0_1),.Y(imd_Y12));
INVC inst_inv_b12_1_0 (.A(imd_Y12),.Y(Y12));
NANDC2x1 inst_clockedAND_b12_12 (.A(CLK),.B(Y12),.Y(imd_YF12));
INVC inst_clockedinv_b12_12 (.A(imd_YF12),.Y(YF12));


NANDC2x1 inst_and_b13_0_0 (.A(A0),.B(A1_inv),.Y(imd_wire13_0_0));
INVC inst_inv_b13_0_0 (.A(imd_wire13_0_0),.Y(wire13_0_0));
NANDC2x1 inst_and_b13_0_1 (.A(A2),.B(A3),.Y(imd_wire13_0_1));
INVC inst_inv_b13_0_1 (.A(imd_wire13_0_1),.Y(wire13_0_1));
NANDC2x1 inst_and_b13_1_0 (.A(wire13_0_0),.B(wire13_0_1),.Y(imd_Y13));
INVC inst_inv_b13_1_0 (.A(imd_Y13),.Y(Y13));
NANDC2x1 inst_clockedAND_b13_13 (.A(CLK),.B(Y13),.Y(imd_YF13));
INVC inst_clockedinv_b13_13 (.A(imd_YF13),.Y(YF13));


NANDC2x1 inst_and_b14_0_0 (.A(A0_inv),.B(A1),.Y(imd_wire14_0_0));
INVC inst_inv_b14_0_0 (.A(imd_wire14_0_0),.Y(wire14_0_0));
NANDC2x1 inst_and_b14_0_1 (.A(A2),.B(A3),.Y(imd_wire14_0_1));
INVC inst_inv_b14_0_1 (.A(imd_wire14_0_1),.Y(wire14_0_1));
NANDC2x1 inst_and_b14_1_0 (.A(wire14_0_0),.B(wire14_0_1),.Y(imd_Y14));
INVC inst_inv_b14_1_0 (.A(imd_Y14),.Y(Y14));
NANDC2x1 inst_clockedAND_b14_14 (.A(CLK),.B(Y14),.Y(imd_YF14));
INVC inst_clockedinv_b14_14 (.A(imd_YF14),.Y(YF14));


NANDC2x1 inst_and_b15_0_0 (.A(A0),.B(A1),.Y(imd_wire15_0_0));
INVC inst_inv_b15_0_0 (.A(imd_wire15_0_0),.Y(wire15_0_0));
NANDC2x1 inst_and_b15_0_1 (.A(A2),.B(A3),.Y(imd_wire15_0_1));
INVC inst_inv_b15_0_1 (.A(imd_wire15_0_1),.Y(wire15_0_1));
NANDC2x1 inst_and_b15_1_0 (.A(wire15_0_0),.B(wire15_0_1),.Y(imd_Y15));
INVC inst_inv_b15_1_0 (.A(imd_Y15),.Y(Y15));
NANDC2x1 inst_clockedAND_b15_15 (.A(CLK),.B(Y15),.Y(imd_YF15));
INVC inst_clockedinv_b15_15 (.A(imd_YF15),.Y(YF15));


endmodule
module columnMux(A0,Abar0,A1,Abar1,A2,Abar2,A3,Abar3,A4,Abar4,A5,Abar5,A6,Abar6,A7,Abar7,A8,Abar8,A9,Abar9,A10,Abar10,A11,Abar11,A12,Abar12,A13,Abar13,A14,Abar14,A15,Abar15,sel0,sel1,sel2,sel3,sel4,sel5,sel6,sel7,sel8,sel9,sel10,sel11,sel12,sel13,sel14,sel15,Y,Ybar);
input A0;
input Abar0;
input A1;
input Abar1;
input A2;
input Abar2;
input A3;
input Abar3;
input A4;
input Abar4;
input A5;
input Abar5;
input A6;
input Abar6;
input A7;
input Abar7;
input A8;
input Abar8;
input A9;
input Abar9;
input A10;
input Abar10;
input A11;
input Abar11;
input A12;
input Abar12;
input A13;
input Abar13;
input A14;
input Abar14;
input A15;
input Abar15;
input sel0;
input sel1;
input sel2;
input sel3;
input sel4;
input sel5;
input sel6;
input sel7;
input sel8;
input sel9;
input sel10;
input sel11;
input sel12;
input sel13;
input sel14;
input sel15;
output Y;
output Ybar;
muxTrans wire0 (.A(A0),.S(sel0),.Y(Y));
muxTrans wire1 (.A(Abar0),.S(sel0),.Y(Ybar));
muxTrans wire2 (.A(A1),.S(sel1),.Y(Y));
muxTrans wire3 (.A(Abar1),.S(sel1),.Y(Ybar));
muxTrans wire4 (.A(A2),.S(sel2),.Y(Y));
muxTrans wire5 (.A(Abar2),.S(sel2),.Y(Ybar));
muxTrans wire6 (.A(A3),.S(sel3),.Y(Y));
muxTrans wire7 (.A(Abar3),.S(sel3),.Y(Ybar));
muxTrans wire8 (.A(A4),.S(sel4),.Y(Y));
muxTrans wire9 (.A(Abar4),.S(sel4),.Y(Ybar));
muxTrans wire10 (.A(A5),.S(sel5),.Y(Y));
muxTrans wire11 (.A(Abar5),.S(sel5),.Y(Ybar));
muxTrans wire12 (.A(A6),.S(sel6),.Y(Y));
muxTrans wire13 (.A(Abar6),.S(sel6),.Y(Ybar));
muxTrans wire14 (.A(A7),.S(sel7),.Y(Y));
muxTrans wire15 (.A(Abar7),.S(sel7),.Y(Ybar));
muxTrans wire16 (.A(A8),.S(sel8),.Y(Y));
muxTrans wire17 (.A(Abar8),.S(sel8),.Y(Ybar));
muxTrans wire18 (.A(A9),.S(sel9),.Y(Y));
muxTrans wire19 (.A(Abar9),.S(sel9),.Y(Ybar));
muxTrans wire20 (.A(A10),.S(sel10),.Y(Y));
muxTrans wire21 (.A(Abar10),.S(sel10),.Y(Ybar));
muxTrans wire22 (.A(A11),.S(sel11),.Y(Y));
muxTrans wire23 (.A(Abar11),.S(sel11),.Y(Ybar));
muxTrans wire24 (.A(A12),.S(sel12),.Y(Y));
muxTrans wire25 (.A(Abar12),.S(sel12),.Y(Ybar));
muxTrans wire26 (.A(A13),.S(sel13),.Y(Y));
muxTrans wire27 (.A(Abar13),.S(sel13),.Y(Ybar));
muxTrans wire28 (.A(A14),.S(sel14),.Y(Y));
muxTrans wire29 (.A(Abar14),.S(sel14),.Y(Ybar));
muxTrans wire30 (.A(A15),.S(sel15),.Y(Y));
muxTrans wire31 (.A(Abar15),.S(sel15),.Y(Ybar));
endmodule
module sram_4kb_256x128x8(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,addr8,addr9,addr10,addr11,din0,din1,din2,din3,din4,din5,din6,din7,dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7,clk,write_en,sense_en);
input addr0;
input addr1;
input addr2;
input addr3;
input addr4;
input addr5;
input addr6;
input addr7;
input addr8;
input addr9;
input addr10;
input addr11;
input din0;
input din1;
input din2;
input din3;
input din4;
input din5;
input din6;
input din7;
output dout0;
output dout1;
output dout2;
output dout3;
output dout4;
output dout5;
output dout6;
output dout7;
input clk;
input write_en;
input sense_en;

specify
    (sense_en  => dout0  ) = 8.6;   
    (sense_en  => dout1  ) = 3.6;   
    (sense_en  => dout2  ) = 2.6;   
    (sense_en  => dout3  ) = 4.6;   
    (sense_en  => dout4  ) = 6.6;   
    (sense_en  => dout5  ) = 8.6;   
    (sense_en  => dout6  ) = 8.6;   
    (sense_en  => dout7  ) = 1.6;   
endspecify

inverter_compiler inst_invComp (.A0(clk),.A0_bar(clk_bar));
invRow inst_invRow(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,inv_addr0,inv_addr1,inv_addr2,inv_addr3,inv_addr4,inv_addr5,inv_addr6,inv_addr7);
invCol inst_invCol(addr8,addr9,addr10,addr11,inv_addr8,inv_addr9,inv_addr10,inv_addr11);
rowDecoder inst_rowDec (addr0,inv_addr0,addr1,inv_addr1,addr2,inv_addr2,addr3,inv_addr3,addr4,inv_addr4,addr5,inv_addr5,addr6,inv_addr6,addr7,inv_addr7,clk_bar,WL0,WL1,WL2,WL3,WL4,WL5,WL6,WL7,WL8,WL9,WL10,WL11,WL12,WL13,WL14,WL15,WL16,WL17,WL18,WL19,WL20,WL21,WL22,WL23,WL24,WL25,WL26,WL27,WL28,WL29,WL30,WL31,WL32,WL33,WL34,WL35,WL36,WL37,WL38,WL39,WL40,WL41,WL42,WL43,WL44,WL45,WL46,WL47,WL48,WL49,WL50,WL51,WL52,WL53,WL54,WL55,WL56,WL57,WL58,WL59,WL60,WL61,WL62,WL63,WL64,WL65,WL66,WL67,WL68,WL69,WL70,WL71,WL72,WL73,WL74,WL75,WL76,WL77,WL78,WL79,WL80,WL81,WL82,WL83,WL84,WL85,WL86,WL87,WL88,WL89,WL90,WL91,WL92,WL93,WL94,WL95,WL96,WL97,WL98,WL99,WL100,WL101,WL102,WL103,WL104,WL105,WL106,WL107,WL108,WL109,WL110,WL111,WL112,WL113,WL114,WL115,WL116,WL117,WL118,WL119,WL120,WL121,WL122,WL123,WL124,WL125,WL126,WL127,WL128,WL129,WL130,WL131,WL132,WL133,WL134,WL135,WL136,WL137,WL138,WL139,WL140,WL141,WL142,WL143,WL144,WL145,WL146,WL147,WL148,WL149,WL150,WL151,WL152,WL153,WL154,WL155,WL156,WL157,WL158,WL159,WL160,WL161,WL162,WL163,WL164,WL165,WL166,WL167,WL168,WL169,WL170,WL171,WL172,WL173,WL174,WL175,WL176,WL177,WL178,WL179,WL180,WL181,WL182,WL183,WL184,WL185,WL186,WL187,WL188,WL189,WL190,WL191,WL192,WL193,WL194,WL195,WL196,WL197,WL198,WL199,WL200,WL201,WL202,WL203,WL204,WL205,WL206,WL207,WL208,WL209,WL210,WL211,WL212,WL213,WL214,WL215,WL216,WL217,WL218,WL219,WL220,WL221,WL222,WL223,WL224,WL225,WL226,WL227,WL228,WL229,WL230,WL231,WL232,WL233,WL234,WL235,WL236,WL237,WL238,WL239,WL240,WL241,WL242,WL243,WL244,WL245,WL246,WL247,WL248,WL249,WL250,WL251,WL252,WL253,WL254,WL255);
colDecoder inst_colDec (addr8,inv_addr8,addr9,inv_addr9,addr10,inv_addr10,addr11,inv_addr11,clk_bar,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15);
sram_cell_6t_5 inst_cell_0_0 (.BL(BL0),.BLN(BLN0),.WL(WL0));
sram_cell_6t_5 inst_cell_0_1 (.BL(BL1),.BLN(BLN1),.WL(WL0));
sram_cell_6t_5 inst_cell_0_2 (.BL(BL2),.BLN(BLN2),.WL(WL0));
sram_cell_6t_5 inst_cell_0_3 (.BL(BL3),.BLN(BLN3),.WL(WL0));
sram_cell_6t_5 inst_cell_0_4 (.BL(BL4),.BLN(BLN4),.WL(WL0));
sram_cell_6t_5 inst_cell_0_5 (.BL(BL5),.BLN(BLN5),.WL(WL0));
sram_cell_6t_5 inst_cell_0_6 (.BL(BL6),.BLN(BLN6),.WL(WL0));
sram_cell_6t_5 inst_cell_0_7 (.BL(BL7),.BLN(BLN7),.WL(WL0));
sram_cell_6t_5 inst_cell_0_8 (.BL(BL8),.BLN(BLN8),.WL(WL0));
sram_cell_6t_5 inst_cell_0_9 (.BL(BL9),.BLN(BLN9),.WL(WL0));
sram_cell_6t_5 inst_cell_0_10 (.BL(BL10),.BLN(BLN10),.WL(WL0));
sram_cell_6t_5 inst_cell_0_11 (.BL(BL11),.BLN(BLN11),.WL(WL0));
sram_cell_6t_5 inst_cell_0_12 (.BL(BL12),.BLN(BLN12),.WL(WL0));
sram_cell_6t_5 inst_cell_0_13 (.BL(BL13),.BLN(BLN13),.WL(WL0));
sram_cell_6t_5 inst_cell_0_14 (.BL(BL14),.BLN(BLN14),.WL(WL0));
sram_cell_6t_5 inst_cell_0_15 (.BL(BL15),.BLN(BLN15),.WL(WL0));
sram_cell_6t_5 inst_cell_0_16 (.BL(BL16),.BLN(BLN16),.WL(WL0));
sram_cell_6t_5 inst_cell_0_17 (.BL(BL17),.BLN(BLN17),.WL(WL0));
sram_cell_6t_5 inst_cell_0_18 (.BL(BL18),.BLN(BLN18),.WL(WL0));
sram_cell_6t_5 inst_cell_0_19 (.BL(BL19),.BLN(BLN19),.WL(WL0));
sram_cell_6t_5 inst_cell_0_20 (.BL(BL20),.BLN(BLN20),.WL(WL0));
sram_cell_6t_5 inst_cell_0_21 (.BL(BL21),.BLN(BLN21),.WL(WL0));
sram_cell_6t_5 inst_cell_0_22 (.BL(BL22),.BLN(BLN22),.WL(WL0));
sram_cell_6t_5 inst_cell_0_23 (.BL(BL23),.BLN(BLN23),.WL(WL0));
sram_cell_6t_5 inst_cell_0_24 (.BL(BL24),.BLN(BLN24),.WL(WL0));
sram_cell_6t_5 inst_cell_0_25 (.BL(BL25),.BLN(BLN25),.WL(WL0));
sram_cell_6t_5 inst_cell_0_26 (.BL(BL26),.BLN(BLN26),.WL(WL0));
sram_cell_6t_5 inst_cell_0_27 (.BL(BL27),.BLN(BLN27),.WL(WL0));
sram_cell_6t_5 inst_cell_0_28 (.BL(BL28),.BLN(BLN28),.WL(WL0));
sram_cell_6t_5 inst_cell_0_29 (.BL(BL29),.BLN(BLN29),.WL(WL0));
sram_cell_6t_5 inst_cell_0_30 (.BL(BL30),.BLN(BLN30),.WL(WL0));
sram_cell_6t_5 inst_cell_0_31 (.BL(BL31),.BLN(BLN31),.WL(WL0));
sram_cell_6t_5 inst_cell_0_32 (.BL(BL32),.BLN(BLN32),.WL(WL0));
sram_cell_6t_5 inst_cell_0_33 (.BL(BL33),.BLN(BLN33),.WL(WL0));
sram_cell_6t_5 inst_cell_0_34 (.BL(BL34),.BLN(BLN34),.WL(WL0));
sram_cell_6t_5 inst_cell_0_35 (.BL(BL35),.BLN(BLN35),.WL(WL0));
sram_cell_6t_5 inst_cell_0_36 (.BL(BL36),.BLN(BLN36),.WL(WL0));
sram_cell_6t_5 inst_cell_0_37 (.BL(BL37),.BLN(BLN37),.WL(WL0));
sram_cell_6t_5 inst_cell_0_38 (.BL(BL38),.BLN(BLN38),.WL(WL0));
sram_cell_6t_5 inst_cell_0_39 (.BL(BL39),.BLN(BLN39),.WL(WL0));
sram_cell_6t_5 inst_cell_0_40 (.BL(BL40),.BLN(BLN40),.WL(WL0));
sram_cell_6t_5 inst_cell_0_41 (.BL(BL41),.BLN(BLN41),.WL(WL0));
sram_cell_6t_5 inst_cell_0_42 (.BL(BL42),.BLN(BLN42),.WL(WL0));
sram_cell_6t_5 inst_cell_0_43 (.BL(BL43),.BLN(BLN43),.WL(WL0));
sram_cell_6t_5 inst_cell_0_44 (.BL(BL44),.BLN(BLN44),.WL(WL0));
sram_cell_6t_5 inst_cell_0_45 (.BL(BL45),.BLN(BLN45),.WL(WL0));
sram_cell_6t_5 inst_cell_0_46 (.BL(BL46),.BLN(BLN46),.WL(WL0));
sram_cell_6t_5 inst_cell_0_47 (.BL(BL47),.BLN(BLN47),.WL(WL0));
sram_cell_6t_5 inst_cell_0_48 (.BL(BL48),.BLN(BLN48),.WL(WL0));
sram_cell_6t_5 inst_cell_0_49 (.BL(BL49),.BLN(BLN49),.WL(WL0));
sram_cell_6t_5 inst_cell_0_50 (.BL(BL50),.BLN(BLN50),.WL(WL0));
sram_cell_6t_5 inst_cell_0_51 (.BL(BL51),.BLN(BLN51),.WL(WL0));
sram_cell_6t_5 inst_cell_0_52 (.BL(BL52),.BLN(BLN52),.WL(WL0));
sram_cell_6t_5 inst_cell_0_53 (.BL(BL53),.BLN(BLN53),.WL(WL0));
sram_cell_6t_5 inst_cell_0_54 (.BL(BL54),.BLN(BLN54),.WL(WL0));
sram_cell_6t_5 inst_cell_0_55 (.BL(BL55),.BLN(BLN55),.WL(WL0));
sram_cell_6t_5 inst_cell_0_56 (.BL(BL56),.BLN(BLN56),.WL(WL0));
sram_cell_6t_5 inst_cell_0_57 (.BL(BL57),.BLN(BLN57),.WL(WL0));
sram_cell_6t_5 inst_cell_0_58 (.BL(BL58),.BLN(BLN58),.WL(WL0));
sram_cell_6t_5 inst_cell_0_59 (.BL(BL59),.BLN(BLN59),.WL(WL0));
sram_cell_6t_5 inst_cell_0_60 (.BL(BL60),.BLN(BLN60),.WL(WL0));
sram_cell_6t_5 inst_cell_0_61 (.BL(BL61),.BLN(BLN61),.WL(WL0));
sram_cell_6t_5 inst_cell_0_62 (.BL(BL62),.BLN(BLN62),.WL(WL0));
sram_cell_6t_5 inst_cell_0_63 (.BL(BL63),.BLN(BLN63),.WL(WL0));
sram_cell_6t_5 inst_cell_0_64 (.BL(BL64),.BLN(BLN64),.WL(WL0));
sram_cell_6t_5 inst_cell_0_65 (.BL(BL65),.BLN(BLN65),.WL(WL0));
sram_cell_6t_5 inst_cell_0_66 (.BL(BL66),.BLN(BLN66),.WL(WL0));
sram_cell_6t_5 inst_cell_0_67 (.BL(BL67),.BLN(BLN67),.WL(WL0));
sram_cell_6t_5 inst_cell_0_68 (.BL(BL68),.BLN(BLN68),.WL(WL0));
sram_cell_6t_5 inst_cell_0_69 (.BL(BL69),.BLN(BLN69),.WL(WL0));
sram_cell_6t_5 inst_cell_0_70 (.BL(BL70),.BLN(BLN70),.WL(WL0));
sram_cell_6t_5 inst_cell_0_71 (.BL(BL71),.BLN(BLN71),.WL(WL0));
sram_cell_6t_5 inst_cell_0_72 (.BL(BL72),.BLN(BLN72),.WL(WL0));
sram_cell_6t_5 inst_cell_0_73 (.BL(BL73),.BLN(BLN73),.WL(WL0));
sram_cell_6t_5 inst_cell_0_74 (.BL(BL74),.BLN(BLN74),.WL(WL0));
sram_cell_6t_5 inst_cell_0_75 (.BL(BL75),.BLN(BLN75),.WL(WL0));
sram_cell_6t_5 inst_cell_0_76 (.BL(BL76),.BLN(BLN76),.WL(WL0));
sram_cell_6t_5 inst_cell_0_77 (.BL(BL77),.BLN(BLN77),.WL(WL0));
sram_cell_6t_5 inst_cell_0_78 (.BL(BL78),.BLN(BLN78),.WL(WL0));
sram_cell_6t_5 inst_cell_0_79 (.BL(BL79),.BLN(BLN79),.WL(WL0));
sram_cell_6t_5 inst_cell_0_80 (.BL(BL80),.BLN(BLN80),.WL(WL0));
sram_cell_6t_5 inst_cell_0_81 (.BL(BL81),.BLN(BLN81),.WL(WL0));
sram_cell_6t_5 inst_cell_0_82 (.BL(BL82),.BLN(BLN82),.WL(WL0));
sram_cell_6t_5 inst_cell_0_83 (.BL(BL83),.BLN(BLN83),.WL(WL0));
sram_cell_6t_5 inst_cell_0_84 (.BL(BL84),.BLN(BLN84),.WL(WL0));
sram_cell_6t_5 inst_cell_0_85 (.BL(BL85),.BLN(BLN85),.WL(WL0));
sram_cell_6t_5 inst_cell_0_86 (.BL(BL86),.BLN(BLN86),.WL(WL0));
sram_cell_6t_5 inst_cell_0_87 (.BL(BL87),.BLN(BLN87),.WL(WL0));
sram_cell_6t_5 inst_cell_0_88 (.BL(BL88),.BLN(BLN88),.WL(WL0));
sram_cell_6t_5 inst_cell_0_89 (.BL(BL89),.BLN(BLN89),.WL(WL0));
sram_cell_6t_5 inst_cell_0_90 (.BL(BL90),.BLN(BLN90),.WL(WL0));
sram_cell_6t_5 inst_cell_0_91 (.BL(BL91),.BLN(BLN91),.WL(WL0));
sram_cell_6t_5 inst_cell_0_92 (.BL(BL92),.BLN(BLN92),.WL(WL0));
sram_cell_6t_5 inst_cell_0_93 (.BL(BL93),.BLN(BLN93),.WL(WL0));
sram_cell_6t_5 inst_cell_0_94 (.BL(BL94),.BLN(BLN94),.WL(WL0));
sram_cell_6t_5 inst_cell_0_95 (.BL(BL95),.BLN(BLN95),.WL(WL0));
sram_cell_6t_5 inst_cell_0_96 (.BL(BL96),.BLN(BLN96),.WL(WL0));
sram_cell_6t_5 inst_cell_0_97 (.BL(BL97),.BLN(BLN97),.WL(WL0));
sram_cell_6t_5 inst_cell_0_98 (.BL(BL98),.BLN(BLN98),.WL(WL0));
sram_cell_6t_5 inst_cell_0_99 (.BL(BL99),.BLN(BLN99),.WL(WL0));
sram_cell_6t_5 inst_cell_0_100 (.BL(BL100),.BLN(BLN100),.WL(WL0));
sram_cell_6t_5 inst_cell_0_101 (.BL(BL101),.BLN(BLN101),.WL(WL0));
sram_cell_6t_5 inst_cell_0_102 (.BL(BL102),.BLN(BLN102),.WL(WL0));
sram_cell_6t_5 inst_cell_0_103 (.BL(BL103),.BLN(BLN103),.WL(WL0));
sram_cell_6t_5 inst_cell_0_104 (.BL(BL104),.BLN(BLN104),.WL(WL0));
sram_cell_6t_5 inst_cell_0_105 (.BL(BL105),.BLN(BLN105),.WL(WL0));
sram_cell_6t_5 inst_cell_0_106 (.BL(BL106),.BLN(BLN106),.WL(WL0));
sram_cell_6t_5 inst_cell_0_107 (.BL(BL107),.BLN(BLN107),.WL(WL0));
sram_cell_6t_5 inst_cell_0_108 (.BL(BL108),.BLN(BLN108),.WL(WL0));
sram_cell_6t_5 inst_cell_0_109 (.BL(BL109),.BLN(BLN109),.WL(WL0));
sram_cell_6t_5 inst_cell_0_110 (.BL(BL110),.BLN(BLN110),.WL(WL0));
sram_cell_6t_5 inst_cell_0_111 (.BL(BL111),.BLN(BLN111),.WL(WL0));
sram_cell_6t_5 inst_cell_0_112 (.BL(BL112),.BLN(BLN112),.WL(WL0));
sram_cell_6t_5 inst_cell_0_113 (.BL(BL113),.BLN(BLN113),.WL(WL0));
sram_cell_6t_5 inst_cell_0_114 (.BL(BL114),.BLN(BLN114),.WL(WL0));
sram_cell_6t_5 inst_cell_0_115 (.BL(BL115),.BLN(BLN115),.WL(WL0));
sram_cell_6t_5 inst_cell_0_116 (.BL(BL116),.BLN(BLN116),.WL(WL0));
sram_cell_6t_5 inst_cell_0_117 (.BL(BL117),.BLN(BLN117),.WL(WL0));
sram_cell_6t_5 inst_cell_0_118 (.BL(BL118),.BLN(BLN118),.WL(WL0));
sram_cell_6t_5 inst_cell_0_119 (.BL(BL119),.BLN(BLN119),.WL(WL0));
sram_cell_6t_5 inst_cell_0_120 (.BL(BL120),.BLN(BLN120),.WL(WL0));
sram_cell_6t_5 inst_cell_0_121 (.BL(BL121),.BLN(BLN121),.WL(WL0));
sram_cell_6t_5 inst_cell_0_122 (.BL(BL122),.BLN(BLN122),.WL(WL0));
sram_cell_6t_5 inst_cell_0_123 (.BL(BL123),.BLN(BLN123),.WL(WL0));
sram_cell_6t_5 inst_cell_0_124 (.BL(BL124),.BLN(BLN124),.WL(WL0));
sram_cell_6t_5 inst_cell_0_125 (.BL(BL125),.BLN(BLN125),.WL(WL0));
sram_cell_6t_5 inst_cell_0_126 (.BL(BL126),.BLN(BLN126),.WL(WL0));
sram_cell_6t_5 inst_cell_0_127 (.BL(BL127),.BLN(BLN127),.WL(WL0));
sram_cell_6t_5 inst_cell_1_0 (.BL(BL0),.BLN(BLN0),.WL(WL1));
sram_cell_6t_5 inst_cell_1_1 (.BL(BL1),.BLN(BLN1),.WL(WL1));
sram_cell_6t_5 inst_cell_1_2 (.BL(BL2),.BLN(BLN2),.WL(WL1));
sram_cell_6t_5 inst_cell_1_3 (.BL(BL3),.BLN(BLN3),.WL(WL1));
sram_cell_6t_5 inst_cell_1_4 (.BL(BL4),.BLN(BLN4),.WL(WL1));
sram_cell_6t_5 inst_cell_1_5 (.BL(BL5),.BLN(BLN5),.WL(WL1));
sram_cell_6t_5 inst_cell_1_6 (.BL(BL6),.BLN(BLN6),.WL(WL1));
sram_cell_6t_5 inst_cell_1_7 (.BL(BL7),.BLN(BLN7),.WL(WL1));
sram_cell_6t_5 inst_cell_1_8 (.BL(BL8),.BLN(BLN8),.WL(WL1));
sram_cell_6t_5 inst_cell_1_9 (.BL(BL9),.BLN(BLN9),.WL(WL1));
sram_cell_6t_5 inst_cell_1_10 (.BL(BL10),.BLN(BLN10),.WL(WL1));
sram_cell_6t_5 inst_cell_1_11 (.BL(BL11),.BLN(BLN11),.WL(WL1));
sram_cell_6t_5 inst_cell_1_12 (.BL(BL12),.BLN(BLN12),.WL(WL1));
sram_cell_6t_5 inst_cell_1_13 (.BL(BL13),.BLN(BLN13),.WL(WL1));
sram_cell_6t_5 inst_cell_1_14 (.BL(BL14),.BLN(BLN14),.WL(WL1));
sram_cell_6t_5 inst_cell_1_15 (.BL(BL15),.BLN(BLN15),.WL(WL1));
sram_cell_6t_5 inst_cell_1_16 (.BL(BL16),.BLN(BLN16),.WL(WL1));
sram_cell_6t_5 inst_cell_1_17 (.BL(BL17),.BLN(BLN17),.WL(WL1));
sram_cell_6t_5 inst_cell_1_18 (.BL(BL18),.BLN(BLN18),.WL(WL1));
sram_cell_6t_5 inst_cell_1_19 (.BL(BL19),.BLN(BLN19),.WL(WL1));
sram_cell_6t_5 inst_cell_1_20 (.BL(BL20),.BLN(BLN20),.WL(WL1));
sram_cell_6t_5 inst_cell_1_21 (.BL(BL21),.BLN(BLN21),.WL(WL1));
sram_cell_6t_5 inst_cell_1_22 (.BL(BL22),.BLN(BLN22),.WL(WL1));
sram_cell_6t_5 inst_cell_1_23 (.BL(BL23),.BLN(BLN23),.WL(WL1));
sram_cell_6t_5 inst_cell_1_24 (.BL(BL24),.BLN(BLN24),.WL(WL1));
sram_cell_6t_5 inst_cell_1_25 (.BL(BL25),.BLN(BLN25),.WL(WL1));
sram_cell_6t_5 inst_cell_1_26 (.BL(BL26),.BLN(BLN26),.WL(WL1));
sram_cell_6t_5 inst_cell_1_27 (.BL(BL27),.BLN(BLN27),.WL(WL1));
sram_cell_6t_5 inst_cell_1_28 (.BL(BL28),.BLN(BLN28),.WL(WL1));
sram_cell_6t_5 inst_cell_1_29 (.BL(BL29),.BLN(BLN29),.WL(WL1));
sram_cell_6t_5 inst_cell_1_30 (.BL(BL30),.BLN(BLN30),.WL(WL1));
sram_cell_6t_5 inst_cell_1_31 (.BL(BL31),.BLN(BLN31),.WL(WL1));
sram_cell_6t_5 inst_cell_1_32 (.BL(BL32),.BLN(BLN32),.WL(WL1));
sram_cell_6t_5 inst_cell_1_33 (.BL(BL33),.BLN(BLN33),.WL(WL1));
sram_cell_6t_5 inst_cell_1_34 (.BL(BL34),.BLN(BLN34),.WL(WL1));
sram_cell_6t_5 inst_cell_1_35 (.BL(BL35),.BLN(BLN35),.WL(WL1));
sram_cell_6t_5 inst_cell_1_36 (.BL(BL36),.BLN(BLN36),.WL(WL1));
sram_cell_6t_5 inst_cell_1_37 (.BL(BL37),.BLN(BLN37),.WL(WL1));
sram_cell_6t_5 inst_cell_1_38 (.BL(BL38),.BLN(BLN38),.WL(WL1));
sram_cell_6t_5 inst_cell_1_39 (.BL(BL39),.BLN(BLN39),.WL(WL1));
sram_cell_6t_5 inst_cell_1_40 (.BL(BL40),.BLN(BLN40),.WL(WL1));
sram_cell_6t_5 inst_cell_1_41 (.BL(BL41),.BLN(BLN41),.WL(WL1));
sram_cell_6t_5 inst_cell_1_42 (.BL(BL42),.BLN(BLN42),.WL(WL1));
sram_cell_6t_5 inst_cell_1_43 (.BL(BL43),.BLN(BLN43),.WL(WL1));
sram_cell_6t_5 inst_cell_1_44 (.BL(BL44),.BLN(BLN44),.WL(WL1));
sram_cell_6t_5 inst_cell_1_45 (.BL(BL45),.BLN(BLN45),.WL(WL1));
sram_cell_6t_5 inst_cell_1_46 (.BL(BL46),.BLN(BLN46),.WL(WL1));
sram_cell_6t_5 inst_cell_1_47 (.BL(BL47),.BLN(BLN47),.WL(WL1));
sram_cell_6t_5 inst_cell_1_48 (.BL(BL48),.BLN(BLN48),.WL(WL1));
sram_cell_6t_5 inst_cell_1_49 (.BL(BL49),.BLN(BLN49),.WL(WL1));
sram_cell_6t_5 inst_cell_1_50 (.BL(BL50),.BLN(BLN50),.WL(WL1));
sram_cell_6t_5 inst_cell_1_51 (.BL(BL51),.BLN(BLN51),.WL(WL1));
sram_cell_6t_5 inst_cell_1_52 (.BL(BL52),.BLN(BLN52),.WL(WL1));
sram_cell_6t_5 inst_cell_1_53 (.BL(BL53),.BLN(BLN53),.WL(WL1));
sram_cell_6t_5 inst_cell_1_54 (.BL(BL54),.BLN(BLN54),.WL(WL1));
sram_cell_6t_5 inst_cell_1_55 (.BL(BL55),.BLN(BLN55),.WL(WL1));
sram_cell_6t_5 inst_cell_1_56 (.BL(BL56),.BLN(BLN56),.WL(WL1));
sram_cell_6t_5 inst_cell_1_57 (.BL(BL57),.BLN(BLN57),.WL(WL1));
sram_cell_6t_5 inst_cell_1_58 (.BL(BL58),.BLN(BLN58),.WL(WL1));
sram_cell_6t_5 inst_cell_1_59 (.BL(BL59),.BLN(BLN59),.WL(WL1));
sram_cell_6t_5 inst_cell_1_60 (.BL(BL60),.BLN(BLN60),.WL(WL1));
sram_cell_6t_5 inst_cell_1_61 (.BL(BL61),.BLN(BLN61),.WL(WL1));
sram_cell_6t_5 inst_cell_1_62 (.BL(BL62),.BLN(BLN62),.WL(WL1));
sram_cell_6t_5 inst_cell_1_63 (.BL(BL63),.BLN(BLN63),.WL(WL1));
sram_cell_6t_5 inst_cell_1_64 (.BL(BL64),.BLN(BLN64),.WL(WL1));
sram_cell_6t_5 inst_cell_1_65 (.BL(BL65),.BLN(BLN65),.WL(WL1));
sram_cell_6t_5 inst_cell_1_66 (.BL(BL66),.BLN(BLN66),.WL(WL1));
sram_cell_6t_5 inst_cell_1_67 (.BL(BL67),.BLN(BLN67),.WL(WL1));
sram_cell_6t_5 inst_cell_1_68 (.BL(BL68),.BLN(BLN68),.WL(WL1));
sram_cell_6t_5 inst_cell_1_69 (.BL(BL69),.BLN(BLN69),.WL(WL1));
sram_cell_6t_5 inst_cell_1_70 (.BL(BL70),.BLN(BLN70),.WL(WL1));
sram_cell_6t_5 inst_cell_1_71 (.BL(BL71),.BLN(BLN71),.WL(WL1));
sram_cell_6t_5 inst_cell_1_72 (.BL(BL72),.BLN(BLN72),.WL(WL1));
sram_cell_6t_5 inst_cell_1_73 (.BL(BL73),.BLN(BLN73),.WL(WL1));
sram_cell_6t_5 inst_cell_1_74 (.BL(BL74),.BLN(BLN74),.WL(WL1));
sram_cell_6t_5 inst_cell_1_75 (.BL(BL75),.BLN(BLN75),.WL(WL1));
sram_cell_6t_5 inst_cell_1_76 (.BL(BL76),.BLN(BLN76),.WL(WL1));
sram_cell_6t_5 inst_cell_1_77 (.BL(BL77),.BLN(BLN77),.WL(WL1));
sram_cell_6t_5 inst_cell_1_78 (.BL(BL78),.BLN(BLN78),.WL(WL1));
sram_cell_6t_5 inst_cell_1_79 (.BL(BL79),.BLN(BLN79),.WL(WL1));
sram_cell_6t_5 inst_cell_1_80 (.BL(BL80),.BLN(BLN80),.WL(WL1));
sram_cell_6t_5 inst_cell_1_81 (.BL(BL81),.BLN(BLN81),.WL(WL1));
sram_cell_6t_5 inst_cell_1_82 (.BL(BL82),.BLN(BLN82),.WL(WL1));
sram_cell_6t_5 inst_cell_1_83 (.BL(BL83),.BLN(BLN83),.WL(WL1));
sram_cell_6t_5 inst_cell_1_84 (.BL(BL84),.BLN(BLN84),.WL(WL1));
sram_cell_6t_5 inst_cell_1_85 (.BL(BL85),.BLN(BLN85),.WL(WL1));
sram_cell_6t_5 inst_cell_1_86 (.BL(BL86),.BLN(BLN86),.WL(WL1));
sram_cell_6t_5 inst_cell_1_87 (.BL(BL87),.BLN(BLN87),.WL(WL1));
sram_cell_6t_5 inst_cell_1_88 (.BL(BL88),.BLN(BLN88),.WL(WL1));
sram_cell_6t_5 inst_cell_1_89 (.BL(BL89),.BLN(BLN89),.WL(WL1));
sram_cell_6t_5 inst_cell_1_90 (.BL(BL90),.BLN(BLN90),.WL(WL1));
sram_cell_6t_5 inst_cell_1_91 (.BL(BL91),.BLN(BLN91),.WL(WL1));
sram_cell_6t_5 inst_cell_1_92 (.BL(BL92),.BLN(BLN92),.WL(WL1));
sram_cell_6t_5 inst_cell_1_93 (.BL(BL93),.BLN(BLN93),.WL(WL1));
sram_cell_6t_5 inst_cell_1_94 (.BL(BL94),.BLN(BLN94),.WL(WL1));
sram_cell_6t_5 inst_cell_1_95 (.BL(BL95),.BLN(BLN95),.WL(WL1));
sram_cell_6t_5 inst_cell_1_96 (.BL(BL96),.BLN(BLN96),.WL(WL1));
sram_cell_6t_5 inst_cell_1_97 (.BL(BL97),.BLN(BLN97),.WL(WL1));
sram_cell_6t_5 inst_cell_1_98 (.BL(BL98),.BLN(BLN98),.WL(WL1));
sram_cell_6t_5 inst_cell_1_99 (.BL(BL99),.BLN(BLN99),.WL(WL1));
sram_cell_6t_5 inst_cell_1_100 (.BL(BL100),.BLN(BLN100),.WL(WL1));
sram_cell_6t_5 inst_cell_1_101 (.BL(BL101),.BLN(BLN101),.WL(WL1));
sram_cell_6t_5 inst_cell_1_102 (.BL(BL102),.BLN(BLN102),.WL(WL1));
sram_cell_6t_5 inst_cell_1_103 (.BL(BL103),.BLN(BLN103),.WL(WL1));
sram_cell_6t_5 inst_cell_1_104 (.BL(BL104),.BLN(BLN104),.WL(WL1));
sram_cell_6t_5 inst_cell_1_105 (.BL(BL105),.BLN(BLN105),.WL(WL1));
sram_cell_6t_5 inst_cell_1_106 (.BL(BL106),.BLN(BLN106),.WL(WL1));
sram_cell_6t_5 inst_cell_1_107 (.BL(BL107),.BLN(BLN107),.WL(WL1));
sram_cell_6t_5 inst_cell_1_108 (.BL(BL108),.BLN(BLN108),.WL(WL1));
sram_cell_6t_5 inst_cell_1_109 (.BL(BL109),.BLN(BLN109),.WL(WL1));
sram_cell_6t_5 inst_cell_1_110 (.BL(BL110),.BLN(BLN110),.WL(WL1));
sram_cell_6t_5 inst_cell_1_111 (.BL(BL111),.BLN(BLN111),.WL(WL1));
sram_cell_6t_5 inst_cell_1_112 (.BL(BL112),.BLN(BLN112),.WL(WL1));
sram_cell_6t_5 inst_cell_1_113 (.BL(BL113),.BLN(BLN113),.WL(WL1));
sram_cell_6t_5 inst_cell_1_114 (.BL(BL114),.BLN(BLN114),.WL(WL1));
sram_cell_6t_5 inst_cell_1_115 (.BL(BL115),.BLN(BLN115),.WL(WL1));
sram_cell_6t_5 inst_cell_1_116 (.BL(BL116),.BLN(BLN116),.WL(WL1));
sram_cell_6t_5 inst_cell_1_117 (.BL(BL117),.BLN(BLN117),.WL(WL1));
sram_cell_6t_5 inst_cell_1_118 (.BL(BL118),.BLN(BLN118),.WL(WL1));
sram_cell_6t_5 inst_cell_1_119 (.BL(BL119),.BLN(BLN119),.WL(WL1));
sram_cell_6t_5 inst_cell_1_120 (.BL(BL120),.BLN(BLN120),.WL(WL1));
sram_cell_6t_5 inst_cell_1_121 (.BL(BL121),.BLN(BLN121),.WL(WL1));
sram_cell_6t_5 inst_cell_1_122 (.BL(BL122),.BLN(BLN122),.WL(WL1));
sram_cell_6t_5 inst_cell_1_123 (.BL(BL123),.BLN(BLN123),.WL(WL1));
sram_cell_6t_5 inst_cell_1_124 (.BL(BL124),.BLN(BLN124),.WL(WL1));
sram_cell_6t_5 inst_cell_1_125 (.BL(BL125),.BLN(BLN125),.WL(WL1));
sram_cell_6t_5 inst_cell_1_126 (.BL(BL126),.BLN(BLN126),.WL(WL1));
sram_cell_6t_5 inst_cell_1_127 (.BL(BL127),.BLN(BLN127),.WL(WL1));
sram_cell_6t_5 inst_cell_2_0 (.BL(BL0),.BLN(BLN0),.WL(WL2));
sram_cell_6t_5 inst_cell_2_1 (.BL(BL1),.BLN(BLN1),.WL(WL2));
sram_cell_6t_5 inst_cell_2_2 (.BL(BL2),.BLN(BLN2),.WL(WL2));
sram_cell_6t_5 inst_cell_2_3 (.BL(BL3),.BLN(BLN3),.WL(WL2));
sram_cell_6t_5 inst_cell_2_4 (.BL(BL4),.BLN(BLN4),.WL(WL2));
sram_cell_6t_5 inst_cell_2_5 (.BL(BL5),.BLN(BLN5),.WL(WL2));
sram_cell_6t_5 inst_cell_2_6 (.BL(BL6),.BLN(BLN6),.WL(WL2));
sram_cell_6t_5 inst_cell_2_7 (.BL(BL7),.BLN(BLN7),.WL(WL2));
sram_cell_6t_5 inst_cell_2_8 (.BL(BL8),.BLN(BLN8),.WL(WL2));
sram_cell_6t_5 inst_cell_2_9 (.BL(BL9),.BLN(BLN9),.WL(WL2));
sram_cell_6t_5 inst_cell_2_10 (.BL(BL10),.BLN(BLN10),.WL(WL2));
sram_cell_6t_5 inst_cell_2_11 (.BL(BL11),.BLN(BLN11),.WL(WL2));
sram_cell_6t_5 inst_cell_2_12 (.BL(BL12),.BLN(BLN12),.WL(WL2));
sram_cell_6t_5 inst_cell_2_13 (.BL(BL13),.BLN(BLN13),.WL(WL2));
sram_cell_6t_5 inst_cell_2_14 (.BL(BL14),.BLN(BLN14),.WL(WL2));
sram_cell_6t_5 inst_cell_2_15 (.BL(BL15),.BLN(BLN15),.WL(WL2));
sram_cell_6t_5 inst_cell_2_16 (.BL(BL16),.BLN(BLN16),.WL(WL2));
sram_cell_6t_5 inst_cell_2_17 (.BL(BL17),.BLN(BLN17),.WL(WL2));
sram_cell_6t_5 inst_cell_2_18 (.BL(BL18),.BLN(BLN18),.WL(WL2));
sram_cell_6t_5 inst_cell_2_19 (.BL(BL19),.BLN(BLN19),.WL(WL2));
sram_cell_6t_5 inst_cell_2_20 (.BL(BL20),.BLN(BLN20),.WL(WL2));
sram_cell_6t_5 inst_cell_2_21 (.BL(BL21),.BLN(BLN21),.WL(WL2));
sram_cell_6t_5 inst_cell_2_22 (.BL(BL22),.BLN(BLN22),.WL(WL2));
sram_cell_6t_5 inst_cell_2_23 (.BL(BL23),.BLN(BLN23),.WL(WL2));
sram_cell_6t_5 inst_cell_2_24 (.BL(BL24),.BLN(BLN24),.WL(WL2));
sram_cell_6t_5 inst_cell_2_25 (.BL(BL25),.BLN(BLN25),.WL(WL2));
sram_cell_6t_5 inst_cell_2_26 (.BL(BL26),.BLN(BLN26),.WL(WL2));
sram_cell_6t_5 inst_cell_2_27 (.BL(BL27),.BLN(BLN27),.WL(WL2));
sram_cell_6t_5 inst_cell_2_28 (.BL(BL28),.BLN(BLN28),.WL(WL2));
sram_cell_6t_5 inst_cell_2_29 (.BL(BL29),.BLN(BLN29),.WL(WL2));
sram_cell_6t_5 inst_cell_2_30 (.BL(BL30),.BLN(BLN30),.WL(WL2));
sram_cell_6t_5 inst_cell_2_31 (.BL(BL31),.BLN(BLN31),.WL(WL2));
sram_cell_6t_5 inst_cell_2_32 (.BL(BL32),.BLN(BLN32),.WL(WL2));
sram_cell_6t_5 inst_cell_2_33 (.BL(BL33),.BLN(BLN33),.WL(WL2));
sram_cell_6t_5 inst_cell_2_34 (.BL(BL34),.BLN(BLN34),.WL(WL2));
sram_cell_6t_5 inst_cell_2_35 (.BL(BL35),.BLN(BLN35),.WL(WL2));
sram_cell_6t_5 inst_cell_2_36 (.BL(BL36),.BLN(BLN36),.WL(WL2));
sram_cell_6t_5 inst_cell_2_37 (.BL(BL37),.BLN(BLN37),.WL(WL2));
sram_cell_6t_5 inst_cell_2_38 (.BL(BL38),.BLN(BLN38),.WL(WL2));
sram_cell_6t_5 inst_cell_2_39 (.BL(BL39),.BLN(BLN39),.WL(WL2));
sram_cell_6t_5 inst_cell_2_40 (.BL(BL40),.BLN(BLN40),.WL(WL2));
sram_cell_6t_5 inst_cell_2_41 (.BL(BL41),.BLN(BLN41),.WL(WL2));
sram_cell_6t_5 inst_cell_2_42 (.BL(BL42),.BLN(BLN42),.WL(WL2));
sram_cell_6t_5 inst_cell_2_43 (.BL(BL43),.BLN(BLN43),.WL(WL2));
sram_cell_6t_5 inst_cell_2_44 (.BL(BL44),.BLN(BLN44),.WL(WL2));
sram_cell_6t_5 inst_cell_2_45 (.BL(BL45),.BLN(BLN45),.WL(WL2));
sram_cell_6t_5 inst_cell_2_46 (.BL(BL46),.BLN(BLN46),.WL(WL2));
sram_cell_6t_5 inst_cell_2_47 (.BL(BL47),.BLN(BLN47),.WL(WL2));
sram_cell_6t_5 inst_cell_2_48 (.BL(BL48),.BLN(BLN48),.WL(WL2));
sram_cell_6t_5 inst_cell_2_49 (.BL(BL49),.BLN(BLN49),.WL(WL2));
sram_cell_6t_5 inst_cell_2_50 (.BL(BL50),.BLN(BLN50),.WL(WL2));
sram_cell_6t_5 inst_cell_2_51 (.BL(BL51),.BLN(BLN51),.WL(WL2));
sram_cell_6t_5 inst_cell_2_52 (.BL(BL52),.BLN(BLN52),.WL(WL2));
sram_cell_6t_5 inst_cell_2_53 (.BL(BL53),.BLN(BLN53),.WL(WL2));
sram_cell_6t_5 inst_cell_2_54 (.BL(BL54),.BLN(BLN54),.WL(WL2));
sram_cell_6t_5 inst_cell_2_55 (.BL(BL55),.BLN(BLN55),.WL(WL2));
sram_cell_6t_5 inst_cell_2_56 (.BL(BL56),.BLN(BLN56),.WL(WL2));
sram_cell_6t_5 inst_cell_2_57 (.BL(BL57),.BLN(BLN57),.WL(WL2));
sram_cell_6t_5 inst_cell_2_58 (.BL(BL58),.BLN(BLN58),.WL(WL2));
sram_cell_6t_5 inst_cell_2_59 (.BL(BL59),.BLN(BLN59),.WL(WL2));
sram_cell_6t_5 inst_cell_2_60 (.BL(BL60),.BLN(BLN60),.WL(WL2));
sram_cell_6t_5 inst_cell_2_61 (.BL(BL61),.BLN(BLN61),.WL(WL2));
sram_cell_6t_5 inst_cell_2_62 (.BL(BL62),.BLN(BLN62),.WL(WL2));
sram_cell_6t_5 inst_cell_2_63 (.BL(BL63),.BLN(BLN63),.WL(WL2));
sram_cell_6t_5 inst_cell_2_64 (.BL(BL64),.BLN(BLN64),.WL(WL2));
sram_cell_6t_5 inst_cell_2_65 (.BL(BL65),.BLN(BLN65),.WL(WL2));
sram_cell_6t_5 inst_cell_2_66 (.BL(BL66),.BLN(BLN66),.WL(WL2));
sram_cell_6t_5 inst_cell_2_67 (.BL(BL67),.BLN(BLN67),.WL(WL2));
sram_cell_6t_5 inst_cell_2_68 (.BL(BL68),.BLN(BLN68),.WL(WL2));
sram_cell_6t_5 inst_cell_2_69 (.BL(BL69),.BLN(BLN69),.WL(WL2));
sram_cell_6t_5 inst_cell_2_70 (.BL(BL70),.BLN(BLN70),.WL(WL2));
sram_cell_6t_5 inst_cell_2_71 (.BL(BL71),.BLN(BLN71),.WL(WL2));
sram_cell_6t_5 inst_cell_2_72 (.BL(BL72),.BLN(BLN72),.WL(WL2));
sram_cell_6t_5 inst_cell_2_73 (.BL(BL73),.BLN(BLN73),.WL(WL2));
sram_cell_6t_5 inst_cell_2_74 (.BL(BL74),.BLN(BLN74),.WL(WL2));
sram_cell_6t_5 inst_cell_2_75 (.BL(BL75),.BLN(BLN75),.WL(WL2));
sram_cell_6t_5 inst_cell_2_76 (.BL(BL76),.BLN(BLN76),.WL(WL2));
sram_cell_6t_5 inst_cell_2_77 (.BL(BL77),.BLN(BLN77),.WL(WL2));
sram_cell_6t_5 inst_cell_2_78 (.BL(BL78),.BLN(BLN78),.WL(WL2));
sram_cell_6t_5 inst_cell_2_79 (.BL(BL79),.BLN(BLN79),.WL(WL2));
sram_cell_6t_5 inst_cell_2_80 (.BL(BL80),.BLN(BLN80),.WL(WL2));
sram_cell_6t_5 inst_cell_2_81 (.BL(BL81),.BLN(BLN81),.WL(WL2));
sram_cell_6t_5 inst_cell_2_82 (.BL(BL82),.BLN(BLN82),.WL(WL2));
sram_cell_6t_5 inst_cell_2_83 (.BL(BL83),.BLN(BLN83),.WL(WL2));
sram_cell_6t_5 inst_cell_2_84 (.BL(BL84),.BLN(BLN84),.WL(WL2));
sram_cell_6t_5 inst_cell_2_85 (.BL(BL85),.BLN(BLN85),.WL(WL2));
sram_cell_6t_5 inst_cell_2_86 (.BL(BL86),.BLN(BLN86),.WL(WL2));
sram_cell_6t_5 inst_cell_2_87 (.BL(BL87),.BLN(BLN87),.WL(WL2));
sram_cell_6t_5 inst_cell_2_88 (.BL(BL88),.BLN(BLN88),.WL(WL2));
sram_cell_6t_5 inst_cell_2_89 (.BL(BL89),.BLN(BLN89),.WL(WL2));
sram_cell_6t_5 inst_cell_2_90 (.BL(BL90),.BLN(BLN90),.WL(WL2));
sram_cell_6t_5 inst_cell_2_91 (.BL(BL91),.BLN(BLN91),.WL(WL2));
sram_cell_6t_5 inst_cell_2_92 (.BL(BL92),.BLN(BLN92),.WL(WL2));
sram_cell_6t_5 inst_cell_2_93 (.BL(BL93),.BLN(BLN93),.WL(WL2));
sram_cell_6t_5 inst_cell_2_94 (.BL(BL94),.BLN(BLN94),.WL(WL2));
sram_cell_6t_5 inst_cell_2_95 (.BL(BL95),.BLN(BLN95),.WL(WL2));
sram_cell_6t_5 inst_cell_2_96 (.BL(BL96),.BLN(BLN96),.WL(WL2));
sram_cell_6t_5 inst_cell_2_97 (.BL(BL97),.BLN(BLN97),.WL(WL2));
sram_cell_6t_5 inst_cell_2_98 (.BL(BL98),.BLN(BLN98),.WL(WL2));
sram_cell_6t_5 inst_cell_2_99 (.BL(BL99),.BLN(BLN99),.WL(WL2));
sram_cell_6t_5 inst_cell_2_100 (.BL(BL100),.BLN(BLN100),.WL(WL2));
sram_cell_6t_5 inst_cell_2_101 (.BL(BL101),.BLN(BLN101),.WL(WL2));
sram_cell_6t_5 inst_cell_2_102 (.BL(BL102),.BLN(BLN102),.WL(WL2));
sram_cell_6t_5 inst_cell_2_103 (.BL(BL103),.BLN(BLN103),.WL(WL2));
sram_cell_6t_5 inst_cell_2_104 (.BL(BL104),.BLN(BLN104),.WL(WL2));
sram_cell_6t_5 inst_cell_2_105 (.BL(BL105),.BLN(BLN105),.WL(WL2));
sram_cell_6t_5 inst_cell_2_106 (.BL(BL106),.BLN(BLN106),.WL(WL2));
sram_cell_6t_5 inst_cell_2_107 (.BL(BL107),.BLN(BLN107),.WL(WL2));
sram_cell_6t_5 inst_cell_2_108 (.BL(BL108),.BLN(BLN108),.WL(WL2));
sram_cell_6t_5 inst_cell_2_109 (.BL(BL109),.BLN(BLN109),.WL(WL2));
sram_cell_6t_5 inst_cell_2_110 (.BL(BL110),.BLN(BLN110),.WL(WL2));
sram_cell_6t_5 inst_cell_2_111 (.BL(BL111),.BLN(BLN111),.WL(WL2));
sram_cell_6t_5 inst_cell_2_112 (.BL(BL112),.BLN(BLN112),.WL(WL2));
sram_cell_6t_5 inst_cell_2_113 (.BL(BL113),.BLN(BLN113),.WL(WL2));
sram_cell_6t_5 inst_cell_2_114 (.BL(BL114),.BLN(BLN114),.WL(WL2));
sram_cell_6t_5 inst_cell_2_115 (.BL(BL115),.BLN(BLN115),.WL(WL2));
sram_cell_6t_5 inst_cell_2_116 (.BL(BL116),.BLN(BLN116),.WL(WL2));
sram_cell_6t_5 inst_cell_2_117 (.BL(BL117),.BLN(BLN117),.WL(WL2));
sram_cell_6t_5 inst_cell_2_118 (.BL(BL118),.BLN(BLN118),.WL(WL2));
sram_cell_6t_5 inst_cell_2_119 (.BL(BL119),.BLN(BLN119),.WL(WL2));
sram_cell_6t_5 inst_cell_2_120 (.BL(BL120),.BLN(BLN120),.WL(WL2));
sram_cell_6t_5 inst_cell_2_121 (.BL(BL121),.BLN(BLN121),.WL(WL2));
sram_cell_6t_5 inst_cell_2_122 (.BL(BL122),.BLN(BLN122),.WL(WL2));
sram_cell_6t_5 inst_cell_2_123 (.BL(BL123),.BLN(BLN123),.WL(WL2));
sram_cell_6t_5 inst_cell_2_124 (.BL(BL124),.BLN(BLN124),.WL(WL2));
sram_cell_6t_5 inst_cell_2_125 (.BL(BL125),.BLN(BLN125),.WL(WL2));
sram_cell_6t_5 inst_cell_2_126 (.BL(BL126),.BLN(BLN126),.WL(WL2));
sram_cell_6t_5 inst_cell_2_127 (.BL(BL127),.BLN(BLN127),.WL(WL2));
sram_cell_6t_5 inst_cell_3_0 (.BL(BL0),.BLN(BLN0),.WL(WL3));
sram_cell_6t_5 inst_cell_3_1 (.BL(BL1),.BLN(BLN1),.WL(WL3));
sram_cell_6t_5 inst_cell_3_2 (.BL(BL2),.BLN(BLN2),.WL(WL3));
sram_cell_6t_5 inst_cell_3_3 (.BL(BL3),.BLN(BLN3),.WL(WL3));
sram_cell_6t_5 inst_cell_3_4 (.BL(BL4),.BLN(BLN4),.WL(WL3));
sram_cell_6t_5 inst_cell_3_5 (.BL(BL5),.BLN(BLN5),.WL(WL3));
sram_cell_6t_5 inst_cell_3_6 (.BL(BL6),.BLN(BLN6),.WL(WL3));
sram_cell_6t_5 inst_cell_3_7 (.BL(BL7),.BLN(BLN7),.WL(WL3));
sram_cell_6t_5 inst_cell_3_8 (.BL(BL8),.BLN(BLN8),.WL(WL3));
sram_cell_6t_5 inst_cell_3_9 (.BL(BL9),.BLN(BLN9),.WL(WL3));
sram_cell_6t_5 inst_cell_3_10 (.BL(BL10),.BLN(BLN10),.WL(WL3));
sram_cell_6t_5 inst_cell_3_11 (.BL(BL11),.BLN(BLN11),.WL(WL3));
sram_cell_6t_5 inst_cell_3_12 (.BL(BL12),.BLN(BLN12),.WL(WL3));
sram_cell_6t_5 inst_cell_3_13 (.BL(BL13),.BLN(BLN13),.WL(WL3));
sram_cell_6t_5 inst_cell_3_14 (.BL(BL14),.BLN(BLN14),.WL(WL3));
sram_cell_6t_5 inst_cell_3_15 (.BL(BL15),.BLN(BLN15),.WL(WL3));
sram_cell_6t_5 inst_cell_3_16 (.BL(BL16),.BLN(BLN16),.WL(WL3));
sram_cell_6t_5 inst_cell_3_17 (.BL(BL17),.BLN(BLN17),.WL(WL3));
sram_cell_6t_5 inst_cell_3_18 (.BL(BL18),.BLN(BLN18),.WL(WL3));
sram_cell_6t_5 inst_cell_3_19 (.BL(BL19),.BLN(BLN19),.WL(WL3));
sram_cell_6t_5 inst_cell_3_20 (.BL(BL20),.BLN(BLN20),.WL(WL3));
sram_cell_6t_5 inst_cell_3_21 (.BL(BL21),.BLN(BLN21),.WL(WL3));
sram_cell_6t_5 inst_cell_3_22 (.BL(BL22),.BLN(BLN22),.WL(WL3));
sram_cell_6t_5 inst_cell_3_23 (.BL(BL23),.BLN(BLN23),.WL(WL3));
sram_cell_6t_5 inst_cell_3_24 (.BL(BL24),.BLN(BLN24),.WL(WL3));
sram_cell_6t_5 inst_cell_3_25 (.BL(BL25),.BLN(BLN25),.WL(WL3));
sram_cell_6t_5 inst_cell_3_26 (.BL(BL26),.BLN(BLN26),.WL(WL3));
sram_cell_6t_5 inst_cell_3_27 (.BL(BL27),.BLN(BLN27),.WL(WL3));
sram_cell_6t_5 inst_cell_3_28 (.BL(BL28),.BLN(BLN28),.WL(WL3));
sram_cell_6t_5 inst_cell_3_29 (.BL(BL29),.BLN(BLN29),.WL(WL3));
sram_cell_6t_5 inst_cell_3_30 (.BL(BL30),.BLN(BLN30),.WL(WL3));
sram_cell_6t_5 inst_cell_3_31 (.BL(BL31),.BLN(BLN31),.WL(WL3));
sram_cell_6t_5 inst_cell_3_32 (.BL(BL32),.BLN(BLN32),.WL(WL3));
sram_cell_6t_5 inst_cell_3_33 (.BL(BL33),.BLN(BLN33),.WL(WL3));
sram_cell_6t_5 inst_cell_3_34 (.BL(BL34),.BLN(BLN34),.WL(WL3));
sram_cell_6t_5 inst_cell_3_35 (.BL(BL35),.BLN(BLN35),.WL(WL3));
sram_cell_6t_5 inst_cell_3_36 (.BL(BL36),.BLN(BLN36),.WL(WL3));
sram_cell_6t_5 inst_cell_3_37 (.BL(BL37),.BLN(BLN37),.WL(WL3));
sram_cell_6t_5 inst_cell_3_38 (.BL(BL38),.BLN(BLN38),.WL(WL3));
sram_cell_6t_5 inst_cell_3_39 (.BL(BL39),.BLN(BLN39),.WL(WL3));
sram_cell_6t_5 inst_cell_3_40 (.BL(BL40),.BLN(BLN40),.WL(WL3));
sram_cell_6t_5 inst_cell_3_41 (.BL(BL41),.BLN(BLN41),.WL(WL3));
sram_cell_6t_5 inst_cell_3_42 (.BL(BL42),.BLN(BLN42),.WL(WL3));
sram_cell_6t_5 inst_cell_3_43 (.BL(BL43),.BLN(BLN43),.WL(WL3));
sram_cell_6t_5 inst_cell_3_44 (.BL(BL44),.BLN(BLN44),.WL(WL3));
sram_cell_6t_5 inst_cell_3_45 (.BL(BL45),.BLN(BLN45),.WL(WL3));
sram_cell_6t_5 inst_cell_3_46 (.BL(BL46),.BLN(BLN46),.WL(WL3));
sram_cell_6t_5 inst_cell_3_47 (.BL(BL47),.BLN(BLN47),.WL(WL3));
sram_cell_6t_5 inst_cell_3_48 (.BL(BL48),.BLN(BLN48),.WL(WL3));
sram_cell_6t_5 inst_cell_3_49 (.BL(BL49),.BLN(BLN49),.WL(WL3));
sram_cell_6t_5 inst_cell_3_50 (.BL(BL50),.BLN(BLN50),.WL(WL3));
sram_cell_6t_5 inst_cell_3_51 (.BL(BL51),.BLN(BLN51),.WL(WL3));
sram_cell_6t_5 inst_cell_3_52 (.BL(BL52),.BLN(BLN52),.WL(WL3));
sram_cell_6t_5 inst_cell_3_53 (.BL(BL53),.BLN(BLN53),.WL(WL3));
sram_cell_6t_5 inst_cell_3_54 (.BL(BL54),.BLN(BLN54),.WL(WL3));
sram_cell_6t_5 inst_cell_3_55 (.BL(BL55),.BLN(BLN55),.WL(WL3));
sram_cell_6t_5 inst_cell_3_56 (.BL(BL56),.BLN(BLN56),.WL(WL3));
sram_cell_6t_5 inst_cell_3_57 (.BL(BL57),.BLN(BLN57),.WL(WL3));
sram_cell_6t_5 inst_cell_3_58 (.BL(BL58),.BLN(BLN58),.WL(WL3));
sram_cell_6t_5 inst_cell_3_59 (.BL(BL59),.BLN(BLN59),.WL(WL3));
sram_cell_6t_5 inst_cell_3_60 (.BL(BL60),.BLN(BLN60),.WL(WL3));
sram_cell_6t_5 inst_cell_3_61 (.BL(BL61),.BLN(BLN61),.WL(WL3));
sram_cell_6t_5 inst_cell_3_62 (.BL(BL62),.BLN(BLN62),.WL(WL3));
sram_cell_6t_5 inst_cell_3_63 (.BL(BL63),.BLN(BLN63),.WL(WL3));
sram_cell_6t_5 inst_cell_3_64 (.BL(BL64),.BLN(BLN64),.WL(WL3));
sram_cell_6t_5 inst_cell_3_65 (.BL(BL65),.BLN(BLN65),.WL(WL3));
sram_cell_6t_5 inst_cell_3_66 (.BL(BL66),.BLN(BLN66),.WL(WL3));
sram_cell_6t_5 inst_cell_3_67 (.BL(BL67),.BLN(BLN67),.WL(WL3));
sram_cell_6t_5 inst_cell_3_68 (.BL(BL68),.BLN(BLN68),.WL(WL3));
sram_cell_6t_5 inst_cell_3_69 (.BL(BL69),.BLN(BLN69),.WL(WL3));
sram_cell_6t_5 inst_cell_3_70 (.BL(BL70),.BLN(BLN70),.WL(WL3));
sram_cell_6t_5 inst_cell_3_71 (.BL(BL71),.BLN(BLN71),.WL(WL3));
sram_cell_6t_5 inst_cell_3_72 (.BL(BL72),.BLN(BLN72),.WL(WL3));
sram_cell_6t_5 inst_cell_3_73 (.BL(BL73),.BLN(BLN73),.WL(WL3));
sram_cell_6t_5 inst_cell_3_74 (.BL(BL74),.BLN(BLN74),.WL(WL3));
sram_cell_6t_5 inst_cell_3_75 (.BL(BL75),.BLN(BLN75),.WL(WL3));
sram_cell_6t_5 inst_cell_3_76 (.BL(BL76),.BLN(BLN76),.WL(WL3));
sram_cell_6t_5 inst_cell_3_77 (.BL(BL77),.BLN(BLN77),.WL(WL3));
sram_cell_6t_5 inst_cell_3_78 (.BL(BL78),.BLN(BLN78),.WL(WL3));
sram_cell_6t_5 inst_cell_3_79 (.BL(BL79),.BLN(BLN79),.WL(WL3));
sram_cell_6t_5 inst_cell_3_80 (.BL(BL80),.BLN(BLN80),.WL(WL3));
sram_cell_6t_5 inst_cell_3_81 (.BL(BL81),.BLN(BLN81),.WL(WL3));
sram_cell_6t_5 inst_cell_3_82 (.BL(BL82),.BLN(BLN82),.WL(WL3));
sram_cell_6t_5 inst_cell_3_83 (.BL(BL83),.BLN(BLN83),.WL(WL3));
sram_cell_6t_5 inst_cell_3_84 (.BL(BL84),.BLN(BLN84),.WL(WL3));
sram_cell_6t_5 inst_cell_3_85 (.BL(BL85),.BLN(BLN85),.WL(WL3));
sram_cell_6t_5 inst_cell_3_86 (.BL(BL86),.BLN(BLN86),.WL(WL3));
sram_cell_6t_5 inst_cell_3_87 (.BL(BL87),.BLN(BLN87),.WL(WL3));
sram_cell_6t_5 inst_cell_3_88 (.BL(BL88),.BLN(BLN88),.WL(WL3));
sram_cell_6t_5 inst_cell_3_89 (.BL(BL89),.BLN(BLN89),.WL(WL3));
sram_cell_6t_5 inst_cell_3_90 (.BL(BL90),.BLN(BLN90),.WL(WL3));
sram_cell_6t_5 inst_cell_3_91 (.BL(BL91),.BLN(BLN91),.WL(WL3));
sram_cell_6t_5 inst_cell_3_92 (.BL(BL92),.BLN(BLN92),.WL(WL3));
sram_cell_6t_5 inst_cell_3_93 (.BL(BL93),.BLN(BLN93),.WL(WL3));
sram_cell_6t_5 inst_cell_3_94 (.BL(BL94),.BLN(BLN94),.WL(WL3));
sram_cell_6t_5 inst_cell_3_95 (.BL(BL95),.BLN(BLN95),.WL(WL3));
sram_cell_6t_5 inst_cell_3_96 (.BL(BL96),.BLN(BLN96),.WL(WL3));
sram_cell_6t_5 inst_cell_3_97 (.BL(BL97),.BLN(BLN97),.WL(WL3));
sram_cell_6t_5 inst_cell_3_98 (.BL(BL98),.BLN(BLN98),.WL(WL3));
sram_cell_6t_5 inst_cell_3_99 (.BL(BL99),.BLN(BLN99),.WL(WL3));
sram_cell_6t_5 inst_cell_3_100 (.BL(BL100),.BLN(BLN100),.WL(WL3));
sram_cell_6t_5 inst_cell_3_101 (.BL(BL101),.BLN(BLN101),.WL(WL3));
sram_cell_6t_5 inst_cell_3_102 (.BL(BL102),.BLN(BLN102),.WL(WL3));
sram_cell_6t_5 inst_cell_3_103 (.BL(BL103),.BLN(BLN103),.WL(WL3));
sram_cell_6t_5 inst_cell_3_104 (.BL(BL104),.BLN(BLN104),.WL(WL3));
sram_cell_6t_5 inst_cell_3_105 (.BL(BL105),.BLN(BLN105),.WL(WL3));
sram_cell_6t_5 inst_cell_3_106 (.BL(BL106),.BLN(BLN106),.WL(WL3));
sram_cell_6t_5 inst_cell_3_107 (.BL(BL107),.BLN(BLN107),.WL(WL3));
sram_cell_6t_5 inst_cell_3_108 (.BL(BL108),.BLN(BLN108),.WL(WL3));
sram_cell_6t_5 inst_cell_3_109 (.BL(BL109),.BLN(BLN109),.WL(WL3));
sram_cell_6t_5 inst_cell_3_110 (.BL(BL110),.BLN(BLN110),.WL(WL3));
sram_cell_6t_5 inst_cell_3_111 (.BL(BL111),.BLN(BLN111),.WL(WL3));
sram_cell_6t_5 inst_cell_3_112 (.BL(BL112),.BLN(BLN112),.WL(WL3));
sram_cell_6t_5 inst_cell_3_113 (.BL(BL113),.BLN(BLN113),.WL(WL3));
sram_cell_6t_5 inst_cell_3_114 (.BL(BL114),.BLN(BLN114),.WL(WL3));
sram_cell_6t_5 inst_cell_3_115 (.BL(BL115),.BLN(BLN115),.WL(WL3));
sram_cell_6t_5 inst_cell_3_116 (.BL(BL116),.BLN(BLN116),.WL(WL3));
sram_cell_6t_5 inst_cell_3_117 (.BL(BL117),.BLN(BLN117),.WL(WL3));
sram_cell_6t_5 inst_cell_3_118 (.BL(BL118),.BLN(BLN118),.WL(WL3));
sram_cell_6t_5 inst_cell_3_119 (.BL(BL119),.BLN(BLN119),.WL(WL3));
sram_cell_6t_5 inst_cell_3_120 (.BL(BL120),.BLN(BLN120),.WL(WL3));
sram_cell_6t_5 inst_cell_3_121 (.BL(BL121),.BLN(BLN121),.WL(WL3));
sram_cell_6t_5 inst_cell_3_122 (.BL(BL122),.BLN(BLN122),.WL(WL3));
sram_cell_6t_5 inst_cell_3_123 (.BL(BL123),.BLN(BLN123),.WL(WL3));
sram_cell_6t_5 inst_cell_3_124 (.BL(BL124),.BLN(BLN124),.WL(WL3));
sram_cell_6t_5 inst_cell_3_125 (.BL(BL125),.BLN(BLN125),.WL(WL3));
sram_cell_6t_5 inst_cell_3_126 (.BL(BL126),.BLN(BLN126),.WL(WL3));
sram_cell_6t_5 inst_cell_3_127 (.BL(BL127),.BLN(BLN127),.WL(WL3));
sram_cell_6t_5 inst_cell_4_0 (.BL(BL0),.BLN(BLN0),.WL(WL4));
sram_cell_6t_5 inst_cell_4_1 (.BL(BL1),.BLN(BLN1),.WL(WL4));
sram_cell_6t_5 inst_cell_4_2 (.BL(BL2),.BLN(BLN2),.WL(WL4));
sram_cell_6t_5 inst_cell_4_3 (.BL(BL3),.BLN(BLN3),.WL(WL4));
sram_cell_6t_5 inst_cell_4_4 (.BL(BL4),.BLN(BLN4),.WL(WL4));
sram_cell_6t_5 inst_cell_4_5 (.BL(BL5),.BLN(BLN5),.WL(WL4));
sram_cell_6t_5 inst_cell_4_6 (.BL(BL6),.BLN(BLN6),.WL(WL4));
sram_cell_6t_5 inst_cell_4_7 (.BL(BL7),.BLN(BLN7),.WL(WL4));
sram_cell_6t_5 inst_cell_4_8 (.BL(BL8),.BLN(BLN8),.WL(WL4));
sram_cell_6t_5 inst_cell_4_9 (.BL(BL9),.BLN(BLN9),.WL(WL4));
sram_cell_6t_5 inst_cell_4_10 (.BL(BL10),.BLN(BLN10),.WL(WL4));
sram_cell_6t_5 inst_cell_4_11 (.BL(BL11),.BLN(BLN11),.WL(WL4));
sram_cell_6t_5 inst_cell_4_12 (.BL(BL12),.BLN(BLN12),.WL(WL4));
sram_cell_6t_5 inst_cell_4_13 (.BL(BL13),.BLN(BLN13),.WL(WL4));
sram_cell_6t_5 inst_cell_4_14 (.BL(BL14),.BLN(BLN14),.WL(WL4));
sram_cell_6t_5 inst_cell_4_15 (.BL(BL15),.BLN(BLN15),.WL(WL4));
sram_cell_6t_5 inst_cell_4_16 (.BL(BL16),.BLN(BLN16),.WL(WL4));
sram_cell_6t_5 inst_cell_4_17 (.BL(BL17),.BLN(BLN17),.WL(WL4));
sram_cell_6t_5 inst_cell_4_18 (.BL(BL18),.BLN(BLN18),.WL(WL4));
sram_cell_6t_5 inst_cell_4_19 (.BL(BL19),.BLN(BLN19),.WL(WL4));
sram_cell_6t_5 inst_cell_4_20 (.BL(BL20),.BLN(BLN20),.WL(WL4));
sram_cell_6t_5 inst_cell_4_21 (.BL(BL21),.BLN(BLN21),.WL(WL4));
sram_cell_6t_5 inst_cell_4_22 (.BL(BL22),.BLN(BLN22),.WL(WL4));
sram_cell_6t_5 inst_cell_4_23 (.BL(BL23),.BLN(BLN23),.WL(WL4));
sram_cell_6t_5 inst_cell_4_24 (.BL(BL24),.BLN(BLN24),.WL(WL4));
sram_cell_6t_5 inst_cell_4_25 (.BL(BL25),.BLN(BLN25),.WL(WL4));
sram_cell_6t_5 inst_cell_4_26 (.BL(BL26),.BLN(BLN26),.WL(WL4));
sram_cell_6t_5 inst_cell_4_27 (.BL(BL27),.BLN(BLN27),.WL(WL4));
sram_cell_6t_5 inst_cell_4_28 (.BL(BL28),.BLN(BLN28),.WL(WL4));
sram_cell_6t_5 inst_cell_4_29 (.BL(BL29),.BLN(BLN29),.WL(WL4));
sram_cell_6t_5 inst_cell_4_30 (.BL(BL30),.BLN(BLN30),.WL(WL4));
sram_cell_6t_5 inst_cell_4_31 (.BL(BL31),.BLN(BLN31),.WL(WL4));
sram_cell_6t_5 inst_cell_4_32 (.BL(BL32),.BLN(BLN32),.WL(WL4));
sram_cell_6t_5 inst_cell_4_33 (.BL(BL33),.BLN(BLN33),.WL(WL4));
sram_cell_6t_5 inst_cell_4_34 (.BL(BL34),.BLN(BLN34),.WL(WL4));
sram_cell_6t_5 inst_cell_4_35 (.BL(BL35),.BLN(BLN35),.WL(WL4));
sram_cell_6t_5 inst_cell_4_36 (.BL(BL36),.BLN(BLN36),.WL(WL4));
sram_cell_6t_5 inst_cell_4_37 (.BL(BL37),.BLN(BLN37),.WL(WL4));
sram_cell_6t_5 inst_cell_4_38 (.BL(BL38),.BLN(BLN38),.WL(WL4));
sram_cell_6t_5 inst_cell_4_39 (.BL(BL39),.BLN(BLN39),.WL(WL4));
sram_cell_6t_5 inst_cell_4_40 (.BL(BL40),.BLN(BLN40),.WL(WL4));
sram_cell_6t_5 inst_cell_4_41 (.BL(BL41),.BLN(BLN41),.WL(WL4));
sram_cell_6t_5 inst_cell_4_42 (.BL(BL42),.BLN(BLN42),.WL(WL4));
sram_cell_6t_5 inst_cell_4_43 (.BL(BL43),.BLN(BLN43),.WL(WL4));
sram_cell_6t_5 inst_cell_4_44 (.BL(BL44),.BLN(BLN44),.WL(WL4));
sram_cell_6t_5 inst_cell_4_45 (.BL(BL45),.BLN(BLN45),.WL(WL4));
sram_cell_6t_5 inst_cell_4_46 (.BL(BL46),.BLN(BLN46),.WL(WL4));
sram_cell_6t_5 inst_cell_4_47 (.BL(BL47),.BLN(BLN47),.WL(WL4));
sram_cell_6t_5 inst_cell_4_48 (.BL(BL48),.BLN(BLN48),.WL(WL4));
sram_cell_6t_5 inst_cell_4_49 (.BL(BL49),.BLN(BLN49),.WL(WL4));
sram_cell_6t_5 inst_cell_4_50 (.BL(BL50),.BLN(BLN50),.WL(WL4));
sram_cell_6t_5 inst_cell_4_51 (.BL(BL51),.BLN(BLN51),.WL(WL4));
sram_cell_6t_5 inst_cell_4_52 (.BL(BL52),.BLN(BLN52),.WL(WL4));
sram_cell_6t_5 inst_cell_4_53 (.BL(BL53),.BLN(BLN53),.WL(WL4));
sram_cell_6t_5 inst_cell_4_54 (.BL(BL54),.BLN(BLN54),.WL(WL4));
sram_cell_6t_5 inst_cell_4_55 (.BL(BL55),.BLN(BLN55),.WL(WL4));
sram_cell_6t_5 inst_cell_4_56 (.BL(BL56),.BLN(BLN56),.WL(WL4));
sram_cell_6t_5 inst_cell_4_57 (.BL(BL57),.BLN(BLN57),.WL(WL4));
sram_cell_6t_5 inst_cell_4_58 (.BL(BL58),.BLN(BLN58),.WL(WL4));
sram_cell_6t_5 inst_cell_4_59 (.BL(BL59),.BLN(BLN59),.WL(WL4));
sram_cell_6t_5 inst_cell_4_60 (.BL(BL60),.BLN(BLN60),.WL(WL4));
sram_cell_6t_5 inst_cell_4_61 (.BL(BL61),.BLN(BLN61),.WL(WL4));
sram_cell_6t_5 inst_cell_4_62 (.BL(BL62),.BLN(BLN62),.WL(WL4));
sram_cell_6t_5 inst_cell_4_63 (.BL(BL63),.BLN(BLN63),.WL(WL4));
sram_cell_6t_5 inst_cell_4_64 (.BL(BL64),.BLN(BLN64),.WL(WL4));
sram_cell_6t_5 inst_cell_4_65 (.BL(BL65),.BLN(BLN65),.WL(WL4));
sram_cell_6t_5 inst_cell_4_66 (.BL(BL66),.BLN(BLN66),.WL(WL4));
sram_cell_6t_5 inst_cell_4_67 (.BL(BL67),.BLN(BLN67),.WL(WL4));
sram_cell_6t_5 inst_cell_4_68 (.BL(BL68),.BLN(BLN68),.WL(WL4));
sram_cell_6t_5 inst_cell_4_69 (.BL(BL69),.BLN(BLN69),.WL(WL4));
sram_cell_6t_5 inst_cell_4_70 (.BL(BL70),.BLN(BLN70),.WL(WL4));
sram_cell_6t_5 inst_cell_4_71 (.BL(BL71),.BLN(BLN71),.WL(WL4));
sram_cell_6t_5 inst_cell_4_72 (.BL(BL72),.BLN(BLN72),.WL(WL4));
sram_cell_6t_5 inst_cell_4_73 (.BL(BL73),.BLN(BLN73),.WL(WL4));
sram_cell_6t_5 inst_cell_4_74 (.BL(BL74),.BLN(BLN74),.WL(WL4));
sram_cell_6t_5 inst_cell_4_75 (.BL(BL75),.BLN(BLN75),.WL(WL4));
sram_cell_6t_5 inst_cell_4_76 (.BL(BL76),.BLN(BLN76),.WL(WL4));
sram_cell_6t_5 inst_cell_4_77 (.BL(BL77),.BLN(BLN77),.WL(WL4));
sram_cell_6t_5 inst_cell_4_78 (.BL(BL78),.BLN(BLN78),.WL(WL4));
sram_cell_6t_5 inst_cell_4_79 (.BL(BL79),.BLN(BLN79),.WL(WL4));
sram_cell_6t_5 inst_cell_4_80 (.BL(BL80),.BLN(BLN80),.WL(WL4));
sram_cell_6t_5 inst_cell_4_81 (.BL(BL81),.BLN(BLN81),.WL(WL4));
sram_cell_6t_5 inst_cell_4_82 (.BL(BL82),.BLN(BLN82),.WL(WL4));
sram_cell_6t_5 inst_cell_4_83 (.BL(BL83),.BLN(BLN83),.WL(WL4));
sram_cell_6t_5 inst_cell_4_84 (.BL(BL84),.BLN(BLN84),.WL(WL4));
sram_cell_6t_5 inst_cell_4_85 (.BL(BL85),.BLN(BLN85),.WL(WL4));
sram_cell_6t_5 inst_cell_4_86 (.BL(BL86),.BLN(BLN86),.WL(WL4));
sram_cell_6t_5 inst_cell_4_87 (.BL(BL87),.BLN(BLN87),.WL(WL4));
sram_cell_6t_5 inst_cell_4_88 (.BL(BL88),.BLN(BLN88),.WL(WL4));
sram_cell_6t_5 inst_cell_4_89 (.BL(BL89),.BLN(BLN89),.WL(WL4));
sram_cell_6t_5 inst_cell_4_90 (.BL(BL90),.BLN(BLN90),.WL(WL4));
sram_cell_6t_5 inst_cell_4_91 (.BL(BL91),.BLN(BLN91),.WL(WL4));
sram_cell_6t_5 inst_cell_4_92 (.BL(BL92),.BLN(BLN92),.WL(WL4));
sram_cell_6t_5 inst_cell_4_93 (.BL(BL93),.BLN(BLN93),.WL(WL4));
sram_cell_6t_5 inst_cell_4_94 (.BL(BL94),.BLN(BLN94),.WL(WL4));
sram_cell_6t_5 inst_cell_4_95 (.BL(BL95),.BLN(BLN95),.WL(WL4));
sram_cell_6t_5 inst_cell_4_96 (.BL(BL96),.BLN(BLN96),.WL(WL4));
sram_cell_6t_5 inst_cell_4_97 (.BL(BL97),.BLN(BLN97),.WL(WL4));
sram_cell_6t_5 inst_cell_4_98 (.BL(BL98),.BLN(BLN98),.WL(WL4));
sram_cell_6t_5 inst_cell_4_99 (.BL(BL99),.BLN(BLN99),.WL(WL4));
sram_cell_6t_5 inst_cell_4_100 (.BL(BL100),.BLN(BLN100),.WL(WL4));
sram_cell_6t_5 inst_cell_4_101 (.BL(BL101),.BLN(BLN101),.WL(WL4));
sram_cell_6t_5 inst_cell_4_102 (.BL(BL102),.BLN(BLN102),.WL(WL4));
sram_cell_6t_5 inst_cell_4_103 (.BL(BL103),.BLN(BLN103),.WL(WL4));
sram_cell_6t_5 inst_cell_4_104 (.BL(BL104),.BLN(BLN104),.WL(WL4));
sram_cell_6t_5 inst_cell_4_105 (.BL(BL105),.BLN(BLN105),.WL(WL4));
sram_cell_6t_5 inst_cell_4_106 (.BL(BL106),.BLN(BLN106),.WL(WL4));
sram_cell_6t_5 inst_cell_4_107 (.BL(BL107),.BLN(BLN107),.WL(WL4));
sram_cell_6t_5 inst_cell_4_108 (.BL(BL108),.BLN(BLN108),.WL(WL4));
sram_cell_6t_5 inst_cell_4_109 (.BL(BL109),.BLN(BLN109),.WL(WL4));
sram_cell_6t_5 inst_cell_4_110 (.BL(BL110),.BLN(BLN110),.WL(WL4));
sram_cell_6t_5 inst_cell_4_111 (.BL(BL111),.BLN(BLN111),.WL(WL4));
sram_cell_6t_5 inst_cell_4_112 (.BL(BL112),.BLN(BLN112),.WL(WL4));
sram_cell_6t_5 inst_cell_4_113 (.BL(BL113),.BLN(BLN113),.WL(WL4));
sram_cell_6t_5 inst_cell_4_114 (.BL(BL114),.BLN(BLN114),.WL(WL4));
sram_cell_6t_5 inst_cell_4_115 (.BL(BL115),.BLN(BLN115),.WL(WL4));
sram_cell_6t_5 inst_cell_4_116 (.BL(BL116),.BLN(BLN116),.WL(WL4));
sram_cell_6t_5 inst_cell_4_117 (.BL(BL117),.BLN(BLN117),.WL(WL4));
sram_cell_6t_5 inst_cell_4_118 (.BL(BL118),.BLN(BLN118),.WL(WL4));
sram_cell_6t_5 inst_cell_4_119 (.BL(BL119),.BLN(BLN119),.WL(WL4));
sram_cell_6t_5 inst_cell_4_120 (.BL(BL120),.BLN(BLN120),.WL(WL4));
sram_cell_6t_5 inst_cell_4_121 (.BL(BL121),.BLN(BLN121),.WL(WL4));
sram_cell_6t_5 inst_cell_4_122 (.BL(BL122),.BLN(BLN122),.WL(WL4));
sram_cell_6t_5 inst_cell_4_123 (.BL(BL123),.BLN(BLN123),.WL(WL4));
sram_cell_6t_5 inst_cell_4_124 (.BL(BL124),.BLN(BLN124),.WL(WL4));
sram_cell_6t_5 inst_cell_4_125 (.BL(BL125),.BLN(BLN125),.WL(WL4));
sram_cell_6t_5 inst_cell_4_126 (.BL(BL126),.BLN(BLN126),.WL(WL4));
sram_cell_6t_5 inst_cell_4_127 (.BL(BL127),.BLN(BLN127),.WL(WL4));
sram_cell_6t_5 inst_cell_5_0 (.BL(BL0),.BLN(BLN0),.WL(WL5));
sram_cell_6t_5 inst_cell_5_1 (.BL(BL1),.BLN(BLN1),.WL(WL5));
sram_cell_6t_5 inst_cell_5_2 (.BL(BL2),.BLN(BLN2),.WL(WL5));
sram_cell_6t_5 inst_cell_5_3 (.BL(BL3),.BLN(BLN3),.WL(WL5));
sram_cell_6t_5 inst_cell_5_4 (.BL(BL4),.BLN(BLN4),.WL(WL5));
sram_cell_6t_5 inst_cell_5_5 (.BL(BL5),.BLN(BLN5),.WL(WL5));
sram_cell_6t_5 inst_cell_5_6 (.BL(BL6),.BLN(BLN6),.WL(WL5));
sram_cell_6t_5 inst_cell_5_7 (.BL(BL7),.BLN(BLN7),.WL(WL5));
sram_cell_6t_5 inst_cell_5_8 (.BL(BL8),.BLN(BLN8),.WL(WL5));
sram_cell_6t_5 inst_cell_5_9 (.BL(BL9),.BLN(BLN9),.WL(WL5));
sram_cell_6t_5 inst_cell_5_10 (.BL(BL10),.BLN(BLN10),.WL(WL5));
sram_cell_6t_5 inst_cell_5_11 (.BL(BL11),.BLN(BLN11),.WL(WL5));
sram_cell_6t_5 inst_cell_5_12 (.BL(BL12),.BLN(BLN12),.WL(WL5));
sram_cell_6t_5 inst_cell_5_13 (.BL(BL13),.BLN(BLN13),.WL(WL5));
sram_cell_6t_5 inst_cell_5_14 (.BL(BL14),.BLN(BLN14),.WL(WL5));
sram_cell_6t_5 inst_cell_5_15 (.BL(BL15),.BLN(BLN15),.WL(WL5));
sram_cell_6t_5 inst_cell_5_16 (.BL(BL16),.BLN(BLN16),.WL(WL5));
sram_cell_6t_5 inst_cell_5_17 (.BL(BL17),.BLN(BLN17),.WL(WL5));
sram_cell_6t_5 inst_cell_5_18 (.BL(BL18),.BLN(BLN18),.WL(WL5));
sram_cell_6t_5 inst_cell_5_19 (.BL(BL19),.BLN(BLN19),.WL(WL5));
sram_cell_6t_5 inst_cell_5_20 (.BL(BL20),.BLN(BLN20),.WL(WL5));
sram_cell_6t_5 inst_cell_5_21 (.BL(BL21),.BLN(BLN21),.WL(WL5));
sram_cell_6t_5 inst_cell_5_22 (.BL(BL22),.BLN(BLN22),.WL(WL5));
sram_cell_6t_5 inst_cell_5_23 (.BL(BL23),.BLN(BLN23),.WL(WL5));
sram_cell_6t_5 inst_cell_5_24 (.BL(BL24),.BLN(BLN24),.WL(WL5));
sram_cell_6t_5 inst_cell_5_25 (.BL(BL25),.BLN(BLN25),.WL(WL5));
sram_cell_6t_5 inst_cell_5_26 (.BL(BL26),.BLN(BLN26),.WL(WL5));
sram_cell_6t_5 inst_cell_5_27 (.BL(BL27),.BLN(BLN27),.WL(WL5));
sram_cell_6t_5 inst_cell_5_28 (.BL(BL28),.BLN(BLN28),.WL(WL5));
sram_cell_6t_5 inst_cell_5_29 (.BL(BL29),.BLN(BLN29),.WL(WL5));
sram_cell_6t_5 inst_cell_5_30 (.BL(BL30),.BLN(BLN30),.WL(WL5));
sram_cell_6t_5 inst_cell_5_31 (.BL(BL31),.BLN(BLN31),.WL(WL5));
sram_cell_6t_5 inst_cell_5_32 (.BL(BL32),.BLN(BLN32),.WL(WL5));
sram_cell_6t_5 inst_cell_5_33 (.BL(BL33),.BLN(BLN33),.WL(WL5));
sram_cell_6t_5 inst_cell_5_34 (.BL(BL34),.BLN(BLN34),.WL(WL5));
sram_cell_6t_5 inst_cell_5_35 (.BL(BL35),.BLN(BLN35),.WL(WL5));
sram_cell_6t_5 inst_cell_5_36 (.BL(BL36),.BLN(BLN36),.WL(WL5));
sram_cell_6t_5 inst_cell_5_37 (.BL(BL37),.BLN(BLN37),.WL(WL5));
sram_cell_6t_5 inst_cell_5_38 (.BL(BL38),.BLN(BLN38),.WL(WL5));
sram_cell_6t_5 inst_cell_5_39 (.BL(BL39),.BLN(BLN39),.WL(WL5));
sram_cell_6t_5 inst_cell_5_40 (.BL(BL40),.BLN(BLN40),.WL(WL5));
sram_cell_6t_5 inst_cell_5_41 (.BL(BL41),.BLN(BLN41),.WL(WL5));
sram_cell_6t_5 inst_cell_5_42 (.BL(BL42),.BLN(BLN42),.WL(WL5));
sram_cell_6t_5 inst_cell_5_43 (.BL(BL43),.BLN(BLN43),.WL(WL5));
sram_cell_6t_5 inst_cell_5_44 (.BL(BL44),.BLN(BLN44),.WL(WL5));
sram_cell_6t_5 inst_cell_5_45 (.BL(BL45),.BLN(BLN45),.WL(WL5));
sram_cell_6t_5 inst_cell_5_46 (.BL(BL46),.BLN(BLN46),.WL(WL5));
sram_cell_6t_5 inst_cell_5_47 (.BL(BL47),.BLN(BLN47),.WL(WL5));
sram_cell_6t_5 inst_cell_5_48 (.BL(BL48),.BLN(BLN48),.WL(WL5));
sram_cell_6t_5 inst_cell_5_49 (.BL(BL49),.BLN(BLN49),.WL(WL5));
sram_cell_6t_5 inst_cell_5_50 (.BL(BL50),.BLN(BLN50),.WL(WL5));
sram_cell_6t_5 inst_cell_5_51 (.BL(BL51),.BLN(BLN51),.WL(WL5));
sram_cell_6t_5 inst_cell_5_52 (.BL(BL52),.BLN(BLN52),.WL(WL5));
sram_cell_6t_5 inst_cell_5_53 (.BL(BL53),.BLN(BLN53),.WL(WL5));
sram_cell_6t_5 inst_cell_5_54 (.BL(BL54),.BLN(BLN54),.WL(WL5));
sram_cell_6t_5 inst_cell_5_55 (.BL(BL55),.BLN(BLN55),.WL(WL5));
sram_cell_6t_5 inst_cell_5_56 (.BL(BL56),.BLN(BLN56),.WL(WL5));
sram_cell_6t_5 inst_cell_5_57 (.BL(BL57),.BLN(BLN57),.WL(WL5));
sram_cell_6t_5 inst_cell_5_58 (.BL(BL58),.BLN(BLN58),.WL(WL5));
sram_cell_6t_5 inst_cell_5_59 (.BL(BL59),.BLN(BLN59),.WL(WL5));
sram_cell_6t_5 inst_cell_5_60 (.BL(BL60),.BLN(BLN60),.WL(WL5));
sram_cell_6t_5 inst_cell_5_61 (.BL(BL61),.BLN(BLN61),.WL(WL5));
sram_cell_6t_5 inst_cell_5_62 (.BL(BL62),.BLN(BLN62),.WL(WL5));
sram_cell_6t_5 inst_cell_5_63 (.BL(BL63),.BLN(BLN63),.WL(WL5));
sram_cell_6t_5 inst_cell_5_64 (.BL(BL64),.BLN(BLN64),.WL(WL5));
sram_cell_6t_5 inst_cell_5_65 (.BL(BL65),.BLN(BLN65),.WL(WL5));
sram_cell_6t_5 inst_cell_5_66 (.BL(BL66),.BLN(BLN66),.WL(WL5));
sram_cell_6t_5 inst_cell_5_67 (.BL(BL67),.BLN(BLN67),.WL(WL5));
sram_cell_6t_5 inst_cell_5_68 (.BL(BL68),.BLN(BLN68),.WL(WL5));
sram_cell_6t_5 inst_cell_5_69 (.BL(BL69),.BLN(BLN69),.WL(WL5));
sram_cell_6t_5 inst_cell_5_70 (.BL(BL70),.BLN(BLN70),.WL(WL5));
sram_cell_6t_5 inst_cell_5_71 (.BL(BL71),.BLN(BLN71),.WL(WL5));
sram_cell_6t_5 inst_cell_5_72 (.BL(BL72),.BLN(BLN72),.WL(WL5));
sram_cell_6t_5 inst_cell_5_73 (.BL(BL73),.BLN(BLN73),.WL(WL5));
sram_cell_6t_5 inst_cell_5_74 (.BL(BL74),.BLN(BLN74),.WL(WL5));
sram_cell_6t_5 inst_cell_5_75 (.BL(BL75),.BLN(BLN75),.WL(WL5));
sram_cell_6t_5 inst_cell_5_76 (.BL(BL76),.BLN(BLN76),.WL(WL5));
sram_cell_6t_5 inst_cell_5_77 (.BL(BL77),.BLN(BLN77),.WL(WL5));
sram_cell_6t_5 inst_cell_5_78 (.BL(BL78),.BLN(BLN78),.WL(WL5));
sram_cell_6t_5 inst_cell_5_79 (.BL(BL79),.BLN(BLN79),.WL(WL5));
sram_cell_6t_5 inst_cell_5_80 (.BL(BL80),.BLN(BLN80),.WL(WL5));
sram_cell_6t_5 inst_cell_5_81 (.BL(BL81),.BLN(BLN81),.WL(WL5));
sram_cell_6t_5 inst_cell_5_82 (.BL(BL82),.BLN(BLN82),.WL(WL5));
sram_cell_6t_5 inst_cell_5_83 (.BL(BL83),.BLN(BLN83),.WL(WL5));
sram_cell_6t_5 inst_cell_5_84 (.BL(BL84),.BLN(BLN84),.WL(WL5));
sram_cell_6t_5 inst_cell_5_85 (.BL(BL85),.BLN(BLN85),.WL(WL5));
sram_cell_6t_5 inst_cell_5_86 (.BL(BL86),.BLN(BLN86),.WL(WL5));
sram_cell_6t_5 inst_cell_5_87 (.BL(BL87),.BLN(BLN87),.WL(WL5));
sram_cell_6t_5 inst_cell_5_88 (.BL(BL88),.BLN(BLN88),.WL(WL5));
sram_cell_6t_5 inst_cell_5_89 (.BL(BL89),.BLN(BLN89),.WL(WL5));
sram_cell_6t_5 inst_cell_5_90 (.BL(BL90),.BLN(BLN90),.WL(WL5));
sram_cell_6t_5 inst_cell_5_91 (.BL(BL91),.BLN(BLN91),.WL(WL5));
sram_cell_6t_5 inst_cell_5_92 (.BL(BL92),.BLN(BLN92),.WL(WL5));
sram_cell_6t_5 inst_cell_5_93 (.BL(BL93),.BLN(BLN93),.WL(WL5));
sram_cell_6t_5 inst_cell_5_94 (.BL(BL94),.BLN(BLN94),.WL(WL5));
sram_cell_6t_5 inst_cell_5_95 (.BL(BL95),.BLN(BLN95),.WL(WL5));
sram_cell_6t_5 inst_cell_5_96 (.BL(BL96),.BLN(BLN96),.WL(WL5));
sram_cell_6t_5 inst_cell_5_97 (.BL(BL97),.BLN(BLN97),.WL(WL5));
sram_cell_6t_5 inst_cell_5_98 (.BL(BL98),.BLN(BLN98),.WL(WL5));
sram_cell_6t_5 inst_cell_5_99 (.BL(BL99),.BLN(BLN99),.WL(WL5));
sram_cell_6t_5 inst_cell_5_100 (.BL(BL100),.BLN(BLN100),.WL(WL5));
sram_cell_6t_5 inst_cell_5_101 (.BL(BL101),.BLN(BLN101),.WL(WL5));
sram_cell_6t_5 inst_cell_5_102 (.BL(BL102),.BLN(BLN102),.WL(WL5));
sram_cell_6t_5 inst_cell_5_103 (.BL(BL103),.BLN(BLN103),.WL(WL5));
sram_cell_6t_5 inst_cell_5_104 (.BL(BL104),.BLN(BLN104),.WL(WL5));
sram_cell_6t_5 inst_cell_5_105 (.BL(BL105),.BLN(BLN105),.WL(WL5));
sram_cell_6t_5 inst_cell_5_106 (.BL(BL106),.BLN(BLN106),.WL(WL5));
sram_cell_6t_5 inst_cell_5_107 (.BL(BL107),.BLN(BLN107),.WL(WL5));
sram_cell_6t_5 inst_cell_5_108 (.BL(BL108),.BLN(BLN108),.WL(WL5));
sram_cell_6t_5 inst_cell_5_109 (.BL(BL109),.BLN(BLN109),.WL(WL5));
sram_cell_6t_5 inst_cell_5_110 (.BL(BL110),.BLN(BLN110),.WL(WL5));
sram_cell_6t_5 inst_cell_5_111 (.BL(BL111),.BLN(BLN111),.WL(WL5));
sram_cell_6t_5 inst_cell_5_112 (.BL(BL112),.BLN(BLN112),.WL(WL5));
sram_cell_6t_5 inst_cell_5_113 (.BL(BL113),.BLN(BLN113),.WL(WL5));
sram_cell_6t_5 inst_cell_5_114 (.BL(BL114),.BLN(BLN114),.WL(WL5));
sram_cell_6t_5 inst_cell_5_115 (.BL(BL115),.BLN(BLN115),.WL(WL5));
sram_cell_6t_5 inst_cell_5_116 (.BL(BL116),.BLN(BLN116),.WL(WL5));
sram_cell_6t_5 inst_cell_5_117 (.BL(BL117),.BLN(BLN117),.WL(WL5));
sram_cell_6t_5 inst_cell_5_118 (.BL(BL118),.BLN(BLN118),.WL(WL5));
sram_cell_6t_5 inst_cell_5_119 (.BL(BL119),.BLN(BLN119),.WL(WL5));
sram_cell_6t_5 inst_cell_5_120 (.BL(BL120),.BLN(BLN120),.WL(WL5));
sram_cell_6t_5 inst_cell_5_121 (.BL(BL121),.BLN(BLN121),.WL(WL5));
sram_cell_6t_5 inst_cell_5_122 (.BL(BL122),.BLN(BLN122),.WL(WL5));
sram_cell_6t_5 inst_cell_5_123 (.BL(BL123),.BLN(BLN123),.WL(WL5));
sram_cell_6t_5 inst_cell_5_124 (.BL(BL124),.BLN(BLN124),.WL(WL5));
sram_cell_6t_5 inst_cell_5_125 (.BL(BL125),.BLN(BLN125),.WL(WL5));
sram_cell_6t_5 inst_cell_5_126 (.BL(BL126),.BLN(BLN126),.WL(WL5));
sram_cell_6t_5 inst_cell_5_127 (.BL(BL127),.BLN(BLN127),.WL(WL5));
sram_cell_6t_5 inst_cell_6_0 (.BL(BL0),.BLN(BLN0),.WL(WL6));
sram_cell_6t_5 inst_cell_6_1 (.BL(BL1),.BLN(BLN1),.WL(WL6));
sram_cell_6t_5 inst_cell_6_2 (.BL(BL2),.BLN(BLN2),.WL(WL6));
sram_cell_6t_5 inst_cell_6_3 (.BL(BL3),.BLN(BLN3),.WL(WL6));
sram_cell_6t_5 inst_cell_6_4 (.BL(BL4),.BLN(BLN4),.WL(WL6));
sram_cell_6t_5 inst_cell_6_5 (.BL(BL5),.BLN(BLN5),.WL(WL6));
sram_cell_6t_5 inst_cell_6_6 (.BL(BL6),.BLN(BLN6),.WL(WL6));
sram_cell_6t_5 inst_cell_6_7 (.BL(BL7),.BLN(BLN7),.WL(WL6));
sram_cell_6t_5 inst_cell_6_8 (.BL(BL8),.BLN(BLN8),.WL(WL6));
sram_cell_6t_5 inst_cell_6_9 (.BL(BL9),.BLN(BLN9),.WL(WL6));
sram_cell_6t_5 inst_cell_6_10 (.BL(BL10),.BLN(BLN10),.WL(WL6));
sram_cell_6t_5 inst_cell_6_11 (.BL(BL11),.BLN(BLN11),.WL(WL6));
sram_cell_6t_5 inst_cell_6_12 (.BL(BL12),.BLN(BLN12),.WL(WL6));
sram_cell_6t_5 inst_cell_6_13 (.BL(BL13),.BLN(BLN13),.WL(WL6));
sram_cell_6t_5 inst_cell_6_14 (.BL(BL14),.BLN(BLN14),.WL(WL6));
sram_cell_6t_5 inst_cell_6_15 (.BL(BL15),.BLN(BLN15),.WL(WL6));
sram_cell_6t_5 inst_cell_6_16 (.BL(BL16),.BLN(BLN16),.WL(WL6));
sram_cell_6t_5 inst_cell_6_17 (.BL(BL17),.BLN(BLN17),.WL(WL6));
sram_cell_6t_5 inst_cell_6_18 (.BL(BL18),.BLN(BLN18),.WL(WL6));
sram_cell_6t_5 inst_cell_6_19 (.BL(BL19),.BLN(BLN19),.WL(WL6));
sram_cell_6t_5 inst_cell_6_20 (.BL(BL20),.BLN(BLN20),.WL(WL6));
sram_cell_6t_5 inst_cell_6_21 (.BL(BL21),.BLN(BLN21),.WL(WL6));
sram_cell_6t_5 inst_cell_6_22 (.BL(BL22),.BLN(BLN22),.WL(WL6));
sram_cell_6t_5 inst_cell_6_23 (.BL(BL23),.BLN(BLN23),.WL(WL6));
sram_cell_6t_5 inst_cell_6_24 (.BL(BL24),.BLN(BLN24),.WL(WL6));
sram_cell_6t_5 inst_cell_6_25 (.BL(BL25),.BLN(BLN25),.WL(WL6));
sram_cell_6t_5 inst_cell_6_26 (.BL(BL26),.BLN(BLN26),.WL(WL6));
sram_cell_6t_5 inst_cell_6_27 (.BL(BL27),.BLN(BLN27),.WL(WL6));
sram_cell_6t_5 inst_cell_6_28 (.BL(BL28),.BLN(BLN28),.WL(WL6));
sram_cell_6t_5 inst_cell_6_29 (.BL(BL29),.BLN(BLN29),.WL(WL6));
sram_cell_6t_5 inst_cell_6_30 (.BL(BL30),.BLN(BLN30),.WL(WL6));
sram_cell_6t_5 inst_cell_6_31 (.BL(BL31),.BLN(BLN31),.WL(WL6));
sram_cell_6t_5 inst_cell_6_32 (.BL(BL32),.BLN(BLN32),.WL(WL6));
sram_cell_6t_5 inst_cell_6_33 (.BL(BL33),.BLN(BLN33),.WL(WL6));
sram_cell_6t_5 inst_cell_6_34 (.BL(BL34),.BLN(BLN34),.WL(WL6));
sram_cell_6t_5 inst_cell_6_35 (.BL(BL35),.BLN(BLN35),.WL(WL6));
sram_cell_6t_5 inst_cell_6_36 (.BL(BL36),.BLN(BLN36),.WL(WL6));
sram_cell_6t_5 inst_cell_6_37 (.BL(BL37),.BLN(BLN37),.WL(WL6));
sram_cell_6t_5 inst_cell_6_38 (.BL(BL38),.BLN(BLN38),.WL(WL6));
sram_cell_6t_5 inst_cell_6_39 (.BL(BL39),.BLN(BLN39),.WL(WL6));
sram_cell_6t_5 inst_cell_6_40 (.BL(BL40),.BLN(BLN40),.WL(WL6));
sram_cell_6t_5 inst_cell_6_41 (.BL(BL41),.BLN(BLN41),.WL(WL6));
sram_cell_6t_5 inst_cell_6_42 (.BL(BL42),.BLN(BLN42),.WL(WL6));
sram_cell_6t_5 inst_cell_6_43 (.BL(BL43),.BLN(BLN43),.WL(WL6));
sram_cell_6t_5 inst_cell_6_44 (.BL(BL44),.BLN(BLN44),.WL(WL6));
sram_cell_6t_5 inst_cell_6_45 (.BL(BL45),.BLN(BLN45),.WL(WL6));
sram_cell_6t_5 inst_cell_6_46 (.BL(BL46),.BLN(BLN46),.WL(WL6));
sram_cell_6t_5 inst_cell_6_47 (.BL(BL47),.BLN(BLN47),.WL(WL6));
sram_cell_6t_5 inst_cell_6_48 (.BL(BL48),.BLN(BLN48),.WL(WL6));
sram_cell_6t_5 inst_cell_6_49 (.BL(BL49),.BLN(BLN49),.WL(WL6));
sram_cell_6t_5 inst_cell_6_50 (.BL(BL50),.BLN(BLN50),.WL(WL6));
sram_cell_6t_5 inst_cell_6_51 (.BL(BL51),.BLN(BLN51),.WL(WL6));
sram_cell_6t_5 inst_cell_6_52 (.BL(BL52),.BLN(BLN52),.WL(WL6));
sram_cell_6t_5 inst_cell_6_53 (.BL(BL53),.BLN(BLN53),.WL(WL6));
sram_cell_6t_5 inst_cell_6_54 (.BL(BL54),.BLN(BLN54),.WL(WL6));
sram_cell_6t_5 inst_cell_6_55 (.BL(BL55),.BLN(BLN55),.WL(WL6));
sram_cell_6t_5 inst_cell_6_56 (.BL(BL56),.BLN(BLN56),.WL(WL6));
sram_cell_6t_5 inst_cell_6_57 (.BL(BL57),.BLN(BLN57),.WL(WL6));
sram_cell_6t_5 inst_cell_6_58 (.BL(BL58),.BLN(BLN58),.WL(WL6));
sram_cell_6t_5 inst_cell_6_59 (.BL(BL59),.BLN(BLN59),.WL(WL6));
sram_cell_6t_5 inst_cell_6_60 (.BL(BL60),.BLN(BLN60),.WL(WL6));
sram_cell_6t_5 inst_cell_6_61 (.BL(BL61),.BLN(BLN61),.WL(WL6));
sram_cell_6t_5 inst_cell_6_62 (.BL(BL62),.BLN(BLN62),.WL(WL6));
sram_cell_6t_5 inst_cell_6_63 (.BL(BL63),.BLN(BLN63),.WL(WL6));
sram_cell_6t_5 inst_cell_6_64 (.BL(BL64),.BLN(BLN64),.WL(WL6));
sram_cell_6t_5 inst_cell_6_65 (.BL(BL65),.BLN(BLN65),.WL(WL6));
sram_cell_6t_5 inst_cell_6_66 (.BL(BL66),.BLN(BLN66),.WL(WL6));
sram_cell_6t_5 inst_cell_6_67 (.BL(BL67),.BLN(BLN67),.WL(WL6));
sram_cell_6t_5 inst_cell_6_68 (.BL(BL68),.BLN(BLN68),.WL(WL6));
sram_cell_6t_5 inst_cell_6_69 (.BL(BL69),.BLN(BLN69),.WL(WL6));
sram_cell_6t_5 inst_cell_6_70 (.BL(BL70),.BLN(BLN70),.WL(WL6));
sram_cell_6t_5 inst_cell_6_71 (.BL(BL71),.BLN(BLN71),.WL(WL6));
sram_cell_6t_5 inst_cell_6_72 (.BL(BL72),.BLN(BLN72),.WL(WL6));
sram_cell_6t_5 inst_cell_6_73 (.BL(BL73),.BLN(BLN73),.WL(WL6));
sram_cell_6t_5 inst_cell_6_74 (.BL(BL74),.BLN(BLN74),.WL(WL6));
sram_cell_6t_5 inst_cell_6_75 (.BL(BL75),.BLN(BLN75),.WL(WL6));
sram_cell_6t_5 inst_cell_6_76 (.BL(BL76),.BLN(BLN76),.WL(WL6));
sram_cell_6t_5 inst_cell_6_77 (.BL(BL77),.BLN(BLN77),.WL(WL6));
sram_cell_6t_5 inst_cell_6_78 (.BL(BL78),.BLN(BLN78),.WL(WL6));
sram_cell_6t_5 inst_cell_6_79 (.BL(BL79),.BLN(BLN79),.WL(WL6));
sram_cell_6t_5 inst_cell_6_80 (.BL(BL80),.BLN(BLN80),.WL(WL6));
sram_cell_6t_5 inst_cell_6_81 (.BL(BL81),.BLN(BLN81),.WL(WL6));
sram_cell_6t_5 inst_cell_6_82 (.BL(BL82),.BLN(BLN82),.WL(WL6));
sram_cell_6t_5 inst_cell_6_83 (.BL(BL83),.BLN(BLN83),.WL(WL6));
sram_cell_6t_5 inst_cell_6_84 (.BL(BL84),.BLN(BLN84),.WL(WL6));
sram_cell_6t_5 inst_cell_6_85 (.BL(BL85),.BLN(BLN85),.WL(WL6));
sram_cell_6t_5 inst_cell_6_86 (.BL(BL86),.BLN(BLN86),.WL(WL6));
sram_cell_6t_5 inst_cell_6_87 (.BL(BL87),.BLN(BLN87),.WL(WL6));
sram_cell_6t_5 inst_cell_6_88 (.BL(BL88),.BLN(BLN88),.WL(WL6));
sram_cell_6t_5 inst_cell_6_89 (.BL(BL89),.BLN(BLN89),.WL(WL6));
sram_cell_6t_5 inst_cell_6_90 (.BL(BL90),.BLN(BLN90),.WL(WL6));
sram_cell_6t_5 inst_cell_6_91 (.BL(BL91),.BLN(BLN91),.WL(WL6));
sram_cell_6t_5 inst_cell_6_92 (.BL(BL92),.BLN(BLN92),.WL(WL6));
sram_cell_6t_5 inst_cell_6_93 (.BL(BL93),.BLN(BLN93),.WL(WL6));
sram_cell_6t_5 inst_cell_6_94 (.BL(BL94),.BLN(BLN94),.WL(WL6));
sram_cell_6t_5 inst_cell_6_95 (.BL(BL95),.BLN(BLN95),.WL(WL6));
sram_cell_6t_5 inst_cell_6_96 (.BL(BL96),.BLN(BLN96),.WL(WL6));
sram_cell_6t_5 inst_cell_6_97 (.BL(BL97),.BLN(BLN97),.WL(WL6));
sram_cell_6t_5 inst_cell_6_98 (.BL(BL98),.BLN(BLN98),.WL(WL6));
sram_cell_6t_5 inst_cell_6_99 (.BL(BL99),.BLN(BLN99),.WL(WL6));
sram_cell_6t_5 inst_cell_6_100 (.BL(BL100),.BLN(BLN100),.WL(WL6));
sram_cell_6t_5 inst_cell_6_101 (.BL(BL101),.BLN(BLN101),.WL(WL6));
sram_cell_6t_5 inst_cell_6_102 (.BL(BL102),.BLN(BLN102),.WL(WL6));
sram_cell_6t_5 inst_cell_6_103 (.BL(BL103),.BLN(BLN103),.WL(WL6));
sram_cell_6t_5 inst_cell_6_104 (.BL(BL104),.BLN(BLN104),.WL(WL6));
sram_cell_6t_5 inst_cell_6_105 (.BL(BL105),.BLN(BLN105),.WL(WL6));
sram_cell_6t_5 inst_cell_6_106 (.BL(BL106),.BLN(BLN106),.WL(WL6));
sram_cell_6t_5 inst_cell_6_107 (.BL(BL107),.BLN(BLN107),.WL(WL6));
sram_cell_6t_5 inst_cell_6_108 (.BL(BL108),.BLN(BLN108),.WL(WL6));
sram_cell_6t_5 inst_cell_6_109 (.BL(BL109),.BLN(BLN109),.WL(WL6));
sram_cell_6t_5 inst_cell_6_110 (.BL(BL110),.BLN(BLN110),.WL(WL6));
sram_cell_6t_5 inst_cell_6_111 (.BL(BL111),.BLN(BLN111),.WL(WL6));
sram_cell_6t_5 inst_cell_6_112 (.BL(BL112),.BLN(BLN112),.WL(WL6));
sram_cell_6t_5 inst_cell_6_113 (.BL(BL113),.BLN(BLN113),.WL(WL6));
sram_cell_6t_5 inst_cell_6_114 (.BL(BL114),.BLN(BLN114),.WL(WL6));
sram_cell_6t_5 inst_cell_6_115 (.BL(BL115),.BLN(BLN115),.WL(WL6));
sram_cell_6t_5 inst_cell_6_116 (.BL(BL116),.BLN(BLN116),.WL(WL6));
sram_cell_6t_5 inst_cell_6_117 (.BL(BL117),.BLN(BLN117),.WL(WL6));
sram_cell_6t_5 inst_cell_6_118 (.BL(BL118),.BLN(BLN118),.WL(WL6));
sram_cell_6t_5 inst_cell_6_119 (.BL(BL119),.BLN(BLN119),.WL(WL6));
sram_cell_6t_5 inst_cell_6_120 (.BL(BL120),.BLN(BLN120),.WL(WL6));
sram_cell_6t_5 inst_cell_6_121 (.BL(BL121),.BLN(BLN121),.WL(WL6));
sram_cell_6t_5 inst_cell_6_122 (.BL(BL122),.BLN(BLN122),.WL(WL6));
sram_cell_6t_5 inst_cell_6_123 (.BL(BL123),.BLN(BLN123),.WL(WL6));
sram_cell_6t_5 inst_cell_6_124 (.BL(BL124),.BLN(BLN124),.WL(WL6));
sram_cell_6t_5 inst_cell_6_125 (.BL(BL125),.BLN(BLN125),.WL(WL6));
sram_cell_6t_5 inst_cell_6_126 (.BL(BL126),.BLN(BLN126),.WL(WL6));
sram_cell_6t_5 inst_cell_6_127 (.BL(BL127),.BLN(BLN127),.WL(WL6));
sram_cell_6t_5 inst_cell_7_0 (.BL(BL0),.BLN(BLN0),.WL(WL7));
sram_cell_6t_5 inst_cell_7_1 (.BL(BL1),.BLN(BLN1),.WL(WL7));
sram_cell_6t_5 inst_cell_7_2 (.BL(BL2),.BLN(BLN2),.WL(WL7));
sram_cell_6t_5 inst_cell_7_3 (.BL(BL3),.BLN(BLN3),.WL(WL7));
sram_cell_6t_5 inst_cell_7_4 (.BL(BL4),.BLN(BLN4),.WL(WL7));
sram_cell_6t_5 inst_cell_7_5 (.BL(BL5),.BLN(BLN5),.WL(WL7));
sram_cell_6t_5 inst_cell_7_6 (.BL(BL6),.BLN(BLN6),.WL(WL7));
sram_cell_6t_5 inst_cell_7_7 (.BL(BL7),.BLN(BLN7),.WL(WL7));
sram_cell_6t_5 inst_cell_7_8 (.BL(BL8),.BLN(BLN8),.WL(WL7));
sram_cell_6t_5 inst_cell_7_9 (.BL(BL9),.BLN(BLN9),.WL(WL7));
sram_cell_6t_5 inst_cell_7_10 (.BL(BL10),.BLN(BLN10),.WL(WL7));
sram_cell_6t_5 inst_cell_7_11 (.BL(BL11),.BLN(BLN11),.WL(WL7));
sram_cell_6t_5 inst_cell_7_12 (.BL(BL12),.BLN(BLN12),.WL(WL7));
sram_cell_6t_5 inst_cell_7_13 (.BL(BL13),.BLN(BLN13),.WL(WL7));
sram_cell_6t_5 inst_cell_7_14 (.BL(BL14),.BLN(BLN14),.WL(WL7));
sram_cell_6t_5 inst_cell_7_15 (.BL(BL15),.BLN(BLN15),.WL(WL7));
sram_cell_6t_5 inst_cell_7_16 (.BL(BL16),.BLN(BLN16),.WL(WL7));
sram_cell_6t_5 inst_cell_7_17 (.BL(BL17),.BLN(BLN17),.WL(WL7));
sram_cell_6t_5 inst_cell_7_18 (.BL(BL18),.BLN(BLN18),.WL(WL7));
sram_cell_6t_5 inst_cell_7_19 (.BL(BL19),.BLN(BLN19),.WL(WL7));
sram_cell_6t_5 inst_cell_7_20 (.BL(BL20),.BLN(BLN20),.WL(WL7));
sram_cell_6t_5 inst_cell_7_21 (.BL(BL21),.BLN(BLN21),.WL(WL7));
sram_cell_6t_5 inst_cell_7_22 (.BL(BL22),.BLN(BLN22),.WL(WL7));
sram_cell_6t_5 inst_cell_7_23 (.BL(BL23),.BLN(BLN23),.WL(WL7));
sram_cell_6t_5 inst_cell_7_24 (.BL(BL24),.BLN(BLN24),.WL(WL7));
sram_cell_6t_5 inst_cell_7_25 (.BL(BL25),.BLN(BLN25),.WL(WL7));
sram_cell_6t_5 inst_cell_7_26 (.BL(BL26),.BLN(BLN26),.WL(WL7));
sram_cell_6t_5 inst_cell_7_27 (.BL(BL27),.BLN(BLN27),.WL(WL7));
sram_cell_6t_5 inst_cell_7_28 (.BL(BL28),.BLN(BLN28),.WL(WL7));
sram_cell_6t_5 inst_cell_7_29 (.BL(BL29),.BLN(BLN29),.WL(WL7));
sram_cell_6t_5 inst_cell_7_30 (.BL(BL30),.BLN(BLN30),.WL(WL7));
sram_cell_6t_5 inst_cell_7_31 (.BL(BL31),.BLN(BLN31),.WL(WL7));
sram_cell_6t_5 inst_cell_7_32 (.BL(BL32),.BLN(BLN32),.WL(WL7));
sram_cell_6t_5 inst_cell_7_33 (.BL(BL33),.BLN(BLN33),.WL(WL7));
sram_cell_6t_5 inst_cell_7_34 (.BL(BL34),.BLN(BLN34),.WL(WL7));
sram_cell_6t_5 inst_cell_7_35 (.BL(BL35),.BLN(BLN35),.WL(WL7));
sram_cell_6t_5 inst_cell_7_36 (.BL(BL36),.BLN(BLN36),.WL(WL7));
sram_cell_6t_5 inst_cell_7_37 (.BL(BL37),.BLN(BLN37),.WL(WL7));
sram_cell_6t_5 inst_cell_7_38 (.BL(BL38),.BLN(BLN38),.WL(WL7));
sram_cell_6t_5 inst_cell_7_39 (.BL(BL39),.BLN(BLN39),.WL(WL7));
sram_cell_6t_5 inst_cell_7_40 (.BL(BL40),.BLN(BLN40),.WL(WL7));
sram_cell_6t_5 inst_cell_7_41 (.BL(BL41),.BLN(BLN41),.WL(WL7));
sram_cell_6t_5 inst_cell_7_42 (.BL(BL42),.BLN(BLN42),.WL(WL7));
sram_cell_6t_5 inst_cell_7_43 (.BL(BL43),.BLN(BLN43),.WL(WL7));
sram_cell_6t_5 inst_cell_7_44 (.BL(BL44),.BLN(BLN44),.WL(WL7));
sram_cell_6t_5 inst_cell_7_45 (.BL(BL45),.BLN(BLN45),.WL(WL7));
sram_cell_6t_5 inst_cell_7_46 (.BL(BL46),.BLN(BLN46),.WL(WL7));
sram_cell_6t_5 inst_cell_7_47 (.BL(BL47),.BLN(BLN47),.WL(WL7));
sram_cell_6t_5 inst_cell_7_48 (.BL(BL48),.BLN(BLN48),.WL(WL7));
sram_cell_6t_5 inst_cell_7_49 (.BL(BL49),.BLN(BLN49),.WL(WL7));
sram_cell_6t_5 inst_cell_7_50 (.BL(BL50),.BLN(BLN50),.WL(WL7));
sram_cell_6t_5 inst_cell_7_51 (.BL(BL51),.BLN(BLN51),.WL(WL7));
sram_cell_6t_5 inst_cell_7_52 (.BL(BL52),.BLN(BLN52),.WL(WL7));
sram_cell_6t_5 inst_cell_7_53 (.BL(BL53),.BLN(BLN53),.WL(WL7));
sram_cell_6t_5 inst_cell_7_54 (.BL(BL54),.BLN(BLN54),.WL(WL7));
sram_cell_6t_5 inst_cell_7_55 (.BL(BL55),.BLN(BLN55),.WL(WL7));
sram_cell_6t_5 inst_cell_7_56 (.BL(BL56),.BLN(BLN56),.WL(WL7));
sram_cell_6t_5 inst_cell_7_57 (.BL(BL57),.BLN(BLN57),.WL(WL7));
sram_cell_6t_5 inst_cell_7_58 (.BL(BL58),.BLN(BLN58),.WL(WL7));
sram_cell_6t_5 inst_cell_7_59 (.BL(BL59),.BLN(BLN59),.WL(WL7));
sram_cell_6t_5 inst_cell_7_60 (.BL(BL60),.BLN(BLN60),.WL(WL7));
sram_cell_6t_5 inst_cell_7_61 (.BL(BL61),.BLN(BLN61),.WL(WL7));
sram_cell_6t_5 inst_cell_7_62 (.BL(BL62),.BLN(BLN62),.WL(WL7));
sram_cell_6t_5 inst_cell_7_63 (.BL(BL63),.BLN(BLN63),.WL(WL7));
sram_cell_6t_5 inst_cell_7_64 (.BL(BL64),.BLN(BLN64),.WL(WL7));
sram_cell_6t_5 inst_cell_7_65 (.BL(BL65),.BLN(BLN65),.WL(WL7));
sram_cell_6t_5 inst_cell_7_66 (.BL(BL66),.BLN(BLN66),.WL(WL7));
sram_cell_6t_5 inst_cell_7_67 (.BL(BL67),.BLN(BLN67),.WL(WL7));
sram_cell_6t_5 inst_cell_7_68 (.BL(BL68),.BLN(BLN68),.WL(WL7));
sram_cell_6t_5 inst_cell_7_69 (.BL(BL69),.BLN(BLN69),.WL(WL7));
sram_cell_6t_5 inst_cell_7_70 (.BL(BL70),.BLN(BLN70),.WL(WL7));
sram_cell_6t_5 inst_cell_7_71 (.BL(BL71),.BLN(BLN71),.WL(WL7));
sram_cell_6t_5 inst_cell_7_72 (.BL(BL72),.BLN(BLN72),.WL(WL7));
sram_cell_6t_5 inst_cell_7_73 (.BL(BL73),.BLN(BLN73),.WL(WL7));
sram_cell_6t_5 inst_cell_7_74 (.BL(BL74),.BLN(BLN74),.WL(WL7));
sram_cell_6t_5 inst_cell_7_75 (.BL(BL75),.BLN(BLN75),.WL(WL7));
sram_cell_6t_5 inst_cell_7_76 (.BL(BL76),.BLN(BLN76),.WL(WL7));
sram_cell_6t_5 inst_cell_7_77 (.BL(BL77),.BLN(BLN77),.WL(WL7));
sram_cell_6t_5 inst_cell_7_78 (.BL(BL78),.BLN(BLN78),.WL(WL7));
sram_cell_6t_5 inst_cell_7_79 (.BL(BL79),.BLN(BLN79),.WL(WL7));
sram_cell_6t_5 inst_cell_7_80 (.BL(BL80),.BLN(BLN80),.WL(WL7));
sram_cell_6t_5 inst_cell_7_81 (.BL(BL81),.BLN(BLN81),.WL(WL7));
sram_cell_6t_5 inst_cell_7_82 (.BL(BL82),.BLN(BLN82),.WL(WL7));
sram_cell_6t_5 inst_cell_7_83 (.BL(BL83),.BLN(BLN83),.WL(WL7));
sram_cell_6t_5 inst_cell_7_84 (.BL(BL84),.BLN(BLN84),.WL(WL7));
sram_cell_6t_5 inst_cell_7_85 (.BL(BL85),.BLN(BLN85),.WL(WL7));
sram_cell_6t_5 inst_cell_7_86 (.BL(BL86),.BLN(BLN86),.WL(WL7));
sram_cell_6t_5 inst_cell_7_87 (.BL(BL87),.BLN(BLN87),.WL(WL7));
sram_cell_6t_5 inst_cell_7_88 (.BL(BL88),.BLN(BLN88),.WL(WL7));
sram_cell_6t_5 inst_cell_7_89 (.BL(BL89),.BLN(BLN89),.WL(WL7));
sram_cell_6t_5 inst_cell_7_90 (.BL(BL90),.BLN(BLN90),.WL(WL7));
sram_cell_6t_5 inst_cell_7_91 (.BL(BL91),.BLN(BLN91),.WL(WL7));
sram_cell_6t_5 inst_cell_7_92 (.BL(BL92),.BLN(BLN92),.WL(WL7));
sram_cell_6t_5 inst_cell_7_93 (.BL(BL93),.BLN(BLN93),.WL(WL7));
sram_cell_6t_5 inst_cell_7_94 (.BL(BL94),.BLN(BLN94),.WL(WL7));
sram_cell_6t_5 inst_cell_7_95 (.BL(BL95),.BLN(BLN95),.WL(WL7));
sram_cell_6t_5 inst_cell_7_96 (.BL(BL96),.BLN(BLN96),.WL(WL7));
sram_cell_6t_5 inst_cell_7_97 (.BL(BL97),.BLN(BLN97),.WL(WL7));
sram_cell_6t_5 inst_cell_7_98 (.BL(BL98),.BLN(BLN98),.WL(WL7));
sram_cell_6t_5 inst_cell_7_99 (.BL(BL99),.BLN(BLN99),.WL(WL7));
sram_cell_6t_5 inst_cell_7_100 (.BL(BL100),.BLN(BLN100),.WL(WL7));
sram_cell_6t_5 inst_cell_7_101 (.BL(BL101),.BLN(BLN101),.WL(WL7));
sram_cell_6t_5 inst_cell_7_102 (.BL(BL102),.BLN(BLN102),.WL(WL7));
sram_cell_6t_5 inst_cell_7_103 (.BL(BL103),.BLN(BLN103),.WL(WL7));
sram_cell_6t_5 inst_cell_7_104 (.BL(BL104),.BLN(BLN104),.WL(WL7));
sram_cell_6t_5 inst_cell_7_105 (.BL(BL105),.BLN(BLN105),.WL(WL7));
sram_cell_6t_5 inst_cell_7_106 (.BL(BL106),.BLN(BLN106),.WL(WL7));
sram_cell_6t_5 inst_cell_7_107 (.BL(BL107),.BLN(BLN107),.WL(WL7));
sram_cell_6t_5 inst_cell_7_108 (.BL(BL108),.BLN(BLN108),.WL(WL7));
sram_cell_6t_5 inst_cell_7_109 (.BL(BL109),.BLN(BLN109),.WL(WL7));
sram_cell_6t_5 inst_cell_7_110 (.BL(BL110),.BLN(BLN110),.WL(WL7));
sram_cell_6t_5 inst_cell_7_111 (.BL(BL111),.BLN(BLN111),.WL(WL7));
sram_cell_6t_5 inst_cell_7_112 (.BL(BL112),.BLN(BLN112),.WL(WL7));
sram_cell_6t_5 inst_cell_7_113 (.BL(BL113),.BLN(BLN113),.WL(WL7));
sram_cell_6t_5 inst_cell_7_114 (.BL(BL114),.BLN(BLN114),.WL(WL7));
sram_cell_6t_5 inst_cell_7_115 (.BL(BL115),.BLN(BLN115),.WL(WL7));
sram_cell_6t_5 inst_cell_7_116 (.BL(BL116),.BLN(BLN116),.WL(WL7));
sram_cell_6t_5 inst_cell_7_117 (.BL(BL117),.BLN(BLN117),.WL(WL7));
sram_cell_6t_5 inst_cell_7_118 (.BL(BL118),.BLN(BLN118),.WL(WL7));
sram_cell_6t_5 inst_cell_7_119 (.BL(BL119),.BLN(BLN119),.WL(WL7));
sram_cell_6t_5 inst_cell_7_120 (.BL(BL120),.BLN(BLN120),.WL(WL7));
sram_cell_6t_5 inst_cell_7_121 (.BL(BL121),.BLN(BLN121),.WL(WL7));
sram_cell_6t_5 inst_cell_7_122 (.BL(BL122),.BLN(BLN122),.WL(WL7));
sram_cell_6t_5 inst_cell_7_123 (.BL(BL123),.BLN(BLN123),.WL(WL7));
sram_cell_6t_5 inst_cell_7_124 (.BL(BL124),.BLN(BLN124),.WL(WL7));
sram_cell_6t_5 inst_cell_7_125 (.BL(BL125),.BLN(BLN125),.WL(WL7));
sram_cell_6t_5 inst_cell_7_126 (.BL(BL126),.BLN(BLN126),.WL(WL7));
sram_cell_6t_5 inst_cell_7_127 (.BL(BL127),.BLN(BLN127),.WL(WL7));
sram_cell_6t_5 inst_cell_8_0 (.BL(BL0),.BLN(BLN0),.WL(WL8));
sram_cell_6t_5 inst_cell_8_1 (.BL(BL1),.BLN(BLN1),.WL(WL8));
sram_cell_6t_5 inst_cell_8_2 (.BL(BL2),.BLN(BLN2),.WL(WL8));
sram_cell_6t_5 inst_cell_8_3 (.BL(BL3),.BLN(BLN3),.WL(WL8));
sram_cell_6t_5 inst_cell_8_4 (.BL(BL4),.BLN(BLN4),.WL(WL8));
sram_cell_6t_5 inst_cell_8_5 (.BL(BL5),.BLN(BLN5),.WL(WL8));
sram_cell_6t_5 inst_cell_8_6 (.BL(BL6),.BLN(BLN6),.WL(WL8));
sram_cell_6t_5 inst_cell_8_7 (.BL(BL7),.BLN(BLN7),.WL(WL8));
sram_cell_6t_5 inst_cell_8_8 (.BL(BL8),.BLN(BLN8),.WL(WL8));
sram_cell_6t_5 inst_cell_8_9 (.BL(BL9),.BLN(BLN9),.WL(WL8));
sram_cell_6t_5 inst_cell_8_10 (.BL(BL10),.BLN(BLN10),.WL(WL8));
sram_cell_6t_5 inst_cell_8_11 (.BL(BL11),.BLN(BLN11),.WL(WL8));
sram_cell_6t_5 inst_cell_8_12 (.BL(BL12),.BLN(BLN12),.WL(WL8));
sram_cell_6t_5 inst_cell_8_13 (.BL(BL13),.BLN(BLN13),.WL(WL8));
sram_cell_6t_5 inst_cell_8_14 (.BL(BL14),.BLN(BLN14),.WL(WL8));
sram_cell_6t_5 inst_cell_8_15 (.BL(BL15),.BLN(BLN15),.WL(WL8));
sram_cell_6t_5 inst_cell_8_16 (.BL(BL16),.BLN(BLN16),.WL(WL8));
sram_cell_6t_5 inst_cell_8_17 (.BL(BL17),.BLN(BLN17),.WL(WL8));
sram_cell_6t_5 inst_cell_8_18 (.BL(BL18),.BLN(BLN18),.WL(WL8));
sram_cell_6t_5 inst_cell_8_19 (.BL(BL19),.BLN(BLN19),.WL(WL8));
sram_cell_6t_5 inst_cell_8_20 (.BL(BL20),.BLN(BLN20),.WL(WL8));
sram_cell_6t_5 inst_cell_8_21 (.BL(BL21),.BLN(BLN21),.WL(WL8));
sram_cell_6t_5 inst_cell_8_22 (.BL(BL22),.BLN(BLN22),.WL(WL8));
sram_cell_6t_5 inst_cell_8_23 (.BL(BL23),.BLN(BLN23),.WL(WL8));
sram_cell_6t_5 inst_cell_8_24 (.BL(BL24),.BLN(BLN24),.WL(WL8));
sram_cell_6t_5 inst_cell_8_25 (.BL(BL25),.BLN(BLN25),.WL(WL8));
sram_cell_6t_5 inst_cell_8_26 (.BL(BL26),.BLN(BLN26),.WL(WL8));
sram_cell_6t_5 inst_cell_8_27 (.BL(BL27),.BLN(BLN27),.WL(WL8));
sram_cell_6t_5 inst_cell_8_28 (.BL(BL28),.BLN(BLN28),.WL(WL8));
sram_cell_6t_5 inst_cell_8_29 (.BL(BL29),.BLN(BLN29),.WL(WL8));
sram_cell_6t_5 inst_cell_8_30 (.BL(BL30),.BLN(BLN30),.WL(WL8));
sram_cell_6t_5 inst_cell_8_31 (.BL(BL31),.BLN(BLN31),.WL(WL8));
sram_cell_6t_5 inst_cell_8_32 (.BL(BL32),.BLN(BLN32),.WL(WL8));
sram_cell_6t_5 inst_cell_8_33 (.BL(BL33),.BLN(BLN33),.WL(WL8));
sram_cell_6t_5 inst_cell_8_34 (.BL(BL34),.BLN(BLN34),.WL(WL8));
sram_cell_6t_5 inst_cell_8_35 (.BL(BL35),.BLN(BLN35),.WL(WL8));
sram_cell_6t_5 inst_cell_8_36 (.BL(BL36),.BLN(BLN36),.WL(WL8));
sram_cell_6t_5 inst_cell_8_37 (.BL(BL37),.BLN(BLN37),.WL(WL8));
sram_cell_6t_5 inst_cell_8_38 (.BL(BL38),.BLN(BLN38),.WL(WL8));
sram_cell_6t_5 inst_cell_8_39 (.BL(BL39),.BLN(BLN39),.WL(WL8));
sram_cell_6t_5 inst_cell_8_40 (.BL(BL40),.BLN(BLN40),.WL(WL8));
sram_cell_6t_5 inst_cell_8_41 (.BL(BL41),.BLN(BLN41),.WL(WL8));
sram_cell_6t_5 inst_cell_8_42 (.BL(BL42),.BLN(BLN42),.WL(WL8));
sram_cell_6t_5 inst_cell_8_43 (.BL(BL43),.BLN(BLN43),.WL(WL8));
sram_cell_6t_5 inst_cell_8_44 (.BL(BL44),.BLN(BLN44),.WL(WL8));
sram_cell_6t_5 inst_cell_8_45 (.BL(BL45),.BLN(BLN45),.WL(WL8));
sram_cell_6t_5 inst_cell_8_46 (.BL(BL46),.BLN(BLN46),.WL(WL8));
sram_cell_6t_5 inst_cell_8_47 (.BL(BL47),.BLN(BLN47),.WL(WL8));
sram_cell_6t_5 inst_cell_8_48 (.BL(BL48),.BLN(BLN48),.WL(WL8));
sram_cell_6t_5 inst_cell_8_49 (.BL(BL49),.BLN(BLN49),.WL(WL8));
sram_cell_6t_5 inst_cell_8_50 (.BL(BL50),.BLN(BLN50),.WL(WL8));
sram_cell_6t_5 inst_cell_8_51 (.BL(BL51),.BLN(BLN51),.WL(WL8));
sram_cell_6t_5 inst_cell_8_52 (.BL(BL52),.BLN(BLN52),.WL(WL8));
sram_cell_6t_5 inst_cell_8_53 (.BL(BL53),.BLN(BLN53),.WL(WL8));
sram_cell_6t_5 inst_cell_8_54 (.BL(BL54),.BLN(BLN54),.WL(WL8));
sram_cell_6t_5 inst_cell_8_55 (.BL(BL55),.BLN(BLN55),.WL(WL8));
sram_cell_6t_5 inst_cell_8_56 (.BL(BL56),.BLN(BLN56),.WL(WL8));
sram_cell_6t_5 inst_cell_8_57 (.BL(BL57),.BLN(BLN57),.WL(WL8));
sram_cell_6t_5 inst_cell_8_58 (.BL(BL58),.BLN(BLN58),.WL(WL8));
sram_cell_6t_5 inst_cell_8_59 (.BL(BL59),.BLN(BLN59),.WL(WL8));
sram_cell_6t_5 inst_cell_8_60 (.BL(BL60),.BLN(BLN60),.WL(WL8));
sram_cell_6t_5 inst_cell_8_61 (.BL(BL61),.BLN(BLN61),.WL(WL8));
sram_cell_6t_5 inst_cell_8_62 (.BL(BL62),.BLN(BLN62),.WL(WL8));
sram_cell_6t_5 inst_cell_8_63 (.BL(BL63),.BLN(BLN63),.WL(WL8));
sram_cell_6t_5 inst_cell_8_64 (.BL(BL64),.BLN(BLN64),.WL(WL8));
sram_cell_6t_5 inst_cell_8_65 (.BL(BL65),.BLN(BLN65),.WL(WL8));
sram_cell_6t_5 inst_cell_8_66 (.BL(BL66),.BLN(BLN66),.WL(WL8));
sram_cell_6t_5 inst_cell_8_67 (.BL(BL67),.BLN(BLN67),.WL(WL8));
sram_cell_6t_5 inst_cell_8_68 (.BL(BL68),.BLN(BLN68),.WL(WL8));
sram_cell_6t_5 inst_cell_8_69 (.BL(BL69),.BLN(BLN69),.WL(WL8));
sram_cell_6t_5 inst_cell_8_70 (.BL(BL70),.BLN(BLN70),.WL(WL8));
sram_cell_6t_5 inst_cell_8_71 (.BL(BL71),.BLN(BLN71),.WL(WL8));
sram_cell_6t_5 inst_cell_8_72 (.BL(BL72),.BLN(BLN72),.WL(WL8));
sram_cell_6t_5 inst_cell_8_73 (.BL(BL73),.BLN(BLN73),.WL(WL8));
sram_cell_6t_5 inst_cell_8_74 (.BL(BL74),.BLN(BLN74),.WL(WL8));
sram_cell_6t_5 inst_cell_8_75 (.BL(BL75),.BLN(BLN75),.WL(WL8));
sram_cell_6t_5 inst_cell_8_76 (.BL(BL76),.BLN(BLN76),.WL(WL8));
sram_cell_6t_5 inst_cell_8_77 (.BL(BL77),.BLN(BLN77),.WL(WL8));
sram_cell_6t_5 inst_cell_8_78 (.BL(BL78),.BLN(BLN78),.WL(WL8));
sram_cell_6t_5 inst_cell_8_79 (.BL(BL79),.BLN(BLN79),.WL(WL8));
sram_cell_6t_5 inst_cell_8_80 (.BL(BL80),.BLN(BLN80),.WL(WL8));
sram_cell_6t_5 inst_cell_8_81 (.BL(BL81),.BLN(BLN81),.WL(WL8));
sram_cell_6t_5 inst_cell_8_82 (.BL(BL82),.BLN(BLN82),.WL(WL8));
sram_cell_6t_5 inst_cell_8_83 (.BL(BL83),.BLN(BLN83),.WL(WL8));
sram_cell_6t_5 inst_cell_8_84 (.BL(BL84),.BLN(BLN84),.WL(WL8));
sram_cell_6t_5 inst_cell_8_85 (.BL(BL85),.BLN(BLN85),.WL(WL8));
sram_cell_6t_5 inst_cell_8_86 (.BL(BL86),.BLN(BLN86),.WL(WL8));
sram_cell_6t_5 inst_cell_8_87 (.BL(BL87),.BLN(BLN87),.WL(WL8));
sram_cell_6t_5 inst_cell_8_88 (.BL(BL88),.BLN(BLN88),.WL(WL8));
sram_cell_6t_5 inst_cell_8_89 (.BL(BL89),.BLN(BLN89),.WL(WL8));
sram_cell_6t_5 inst_cell_8_90 (.BL(BL90),.BLN(BLN90),.WL(WL8));
sram_cell_6t_5 inst_cell_8_91 (.BL(BL91),.BLN(BLN91),.WL(WL8));
sram_cell_6t_5 inst_cell_8_92 (.BL(BL92),.BLN(BLN92),.WL(WL8));
sram_cell_6t_5 inst_cell_8_93 (.BL(BL93),.BLN(BLN93),.WL(WL8));
sram_cell_6t_5 inst_cell_8_94 (.BL(BL94),.BLN(BLN94),.WL(WL8));
sram_cell_6t_5 inst_cell_8_95 (.BL(BL95),.BLN(BLN95),.WL(WL8));
sram_cell_6t_5 inst_cell_8_96 (.BL(BL96),.BLN(BLN96),.WL(WL8));
sram_cell_6t_5 inst_cell_8_97 (.BL(BL97),.BLN(BLN97),.WL(WL8));
sram_cell_6t_5 inst_cell_8_98 (.BL(BL98),.BLN(BLN98),.WL(WL8));
sram_cell_6t_5 inst_cell_8_99 (.BL(BL99),.BLN(BLN99),.WL(WL8));
sram_cell_6t_5 inst_cell_8_100 (.BL(BL100),.BLN(BLN100),.WL(WL8));
sram_cell_6t_5 inst_cell_8_101 (.BL(BL101),.BLN(BLN101),.WL(WL8));
sram_cell_6t_5 inst_cell_8_102 (.BL(BL102),.BLN(BLN102),.WL(WL8));
sram_cell_6t_5 inst_cell_8_103 (.BL(BL103),.BLN(BLN103),.WL(WL8));
sram_cell_6t_5 inst_cell_8_104 (.BL(BL104),.BLN(BLN104),.WL(WL8));
sram_cell_6t_5 inst_cell_8_105 (.BL(BL105),.BLN(BLN105),.WL(WL8));
sram_cell_6t_5 inst_cell_8_106 (.BL(BL106),.BLN(BLN106),.WL(WL8));
sram_cell_6t_5 inst_cell_8_107 (.BL(BL107),.BLN(BLN107),.WL(WL8));
sram_cell_6t_5 inst_cell_8_108 (.BL(BL108),.BLN(BLN108),.WL(WL8));
sram_cell_6t_5 inst_cell_8_109 (.BL(BL109),.BLN(BLN109),.WL(WL8));
sram_cell_6t_5 inst_cell_8_110 (.BL(BL110),.BLN(BLN110),.WL(WL8));
sram_cell_6t_5 inst_cell_8_111 (.BL(BL111),.BLN(BLN111),.WL(WL8));
sram_cell_6t_5 inst_cell_8_112 (.BL(BL112),.BLN(BLN112),.WL(WL8));
sram_cell_6t_5 inst_cell_8_113 (.BL(BL113),.BLN(BLN113),.WL(WL8));
sram_cell_6t_5 inst_cell_8_114 (.BL(BL114),.BLN(BLN114),.WL(WL8));
sram_cell_6t_5 inst_cell_8_115 (.BL(BL115),.BLN(BLN115),.WL(WL8));
sram_cell_6t_5 inst_cell_8_116 (.BL(BL116),.BLN(BLN116),.WL(WL8));
sram_cell_6t_5 inst_cell_8_117 (.BL(BL117),.BLN(BLN117),.WL(WL8));
sram_cell_6t_5 inst_cell_8_118 (.BL(BL118),.BLN(BLN118),.WL(WL8));
sram_cell_6t_5 inst_cell_8_119 (.BL(BL119),.BLN(BLN119),.WL(WL8));
sram_cell_6t_5 inst_cell_8_120 (.BL(BL120),.BLN(BLN120),.WL(WL8));
sram_cell_6t_5 inst_cell_8_121 (.BL(BL121),.BLN(BLN121),.WL(WL8));
sram_cell_6t_5 inst_cell_8_122 (.BL(BL122),.BLN(BLN122),.WL(WL8));
sram_cell_6t_5 inst_cell_8_123 (.BL(BL123),.BLN(BLN123),.WL(WL8));
sram_cell_6t_5 inst_cell_8_124 (.BL(BL124),.BLN(BLN124),.WL(WL8));
sram_cell_6t_5 inst_cell_8_125 (.BL(BL125),.BLN(BLN125),.WL(WL8));
sram_cell_6t_5 inst_cell_8_126 (.BL(BL126),.BLN(BLN126),.WL(WL8));
sram_cell_6t_5 inst_cell_8_127 (.BL(BL127),.BLN(BLN127),.WL(WL8));
sram_cell_6t_5 inst_cell_9_0 (.BL(BL0),.BLN(BLN0),.WL(WL9));
sram_cell_6t_5 inst_cell_9_1 (.BL(BL1),.BLN(BLN1),.WL(WL9));
sram_cell_6t_5 inst_cell_9_2 (.BL(BL2),.BLN(BLN2),.WL(WL9));
sram_cell_6t_5 inst_cell_9_3 (.BL(BL3),.BLN(BLN3),.WL(WL9));
sram_cell_6t_5 inst_cell_9_4 (.BL(BL4),.BLN(BLN4),.WL(WL9));
sram_cell_6t_5 inst_cell_9_5 (.BL(BL5),.BLN(BLN5),.WL(WL9));
sram_cell_6t_5 inst_cell_9_6 (.BL(BL6),.BLN(BLN6),.WL(WL9));
sram_cell_6t_5 inst_cell_9_7 (.BL(BL7),.BLN(BLN7),.WL(WL9));
sram_cell_6t_5 inst_cell_9_8 (.BL(BL8),.BLN(BLN8),.WL(WL9));
sram_cell_6t_5 inst_cell_9_9 (.BL(BL9),.BLN(BLN9),.WL(WL9));
sram_cell_6t_5 inst_cell_9_10 (.BL(BL10),.BLN(BLN10),.WL(WL9));
sram_cell_6t_5 inst_cell_9_11 (.BL(BL11),.BLN(BLN11),.WL(WL9));
sram_cell_6t_5 inst_cell_9_12 (.BL(BL12),.BLN(BLN12),.WL(WL9));
sram_cell_6t_5 inst_cell_9_13 (.BL(BL13),.BLN(BLN13),.WL(WL9));
sram_cell_6t_5 inst_cell_9_14 (.BL(BL14),.BLN(BLN14),.WL(WL9));
sram_cell_6t_5 inst_cell_9_15 (.BL(BL15),.BLN(BLN15),.WL(WL9));
sram_cell_6t_5 inst_cell_9_16 (.BL(BL16),.BLN(BLN16),.WL(WL9));
sram_cell_6t_5 inst_cell_9_17 (.BL(BL17),.BLN(BLN17),.WL(WL9));
sram_cell_6t_5 inst_cell_9_18 (.BL(BL18),.BLN(BLN18),.WL(WL9));
sram_cell_6t_5 inst_cell_9_19 (.BL(BL19),.BLN(BLN19),.WL(WL9));
sram_cell_6t_5 inst_cell_9_20 (.BL(BL20),.BLN(BLN20),.WL(WL9));
sram_cell_6t_5 inst_cell_9_21 (.BL(BL21),.BLN(BLN21),.WL(WL9));
sram_cell_6t_5 inst_cell_9_22 (.BL(BL22),.BLN(BLN22),.WL(WL9));
sram_cell_6t_5 inst_cell_9_23 (.BL(BL23),.BLN(BLN23),.WL(WL9));
sram_cell_6t_5 inst_cell_9_24 (.BL(BL24),.BLN(BLN24),.WL(WL9));
sram_cell_6t_5 inst_cell_9_25 (.BL(BL25),.BLN(BLN25),.WL(WL9));
sram_cell_6t_5 inst_cell_9_26 (.BL(BL26),.BLN(BLN26),.WL(WL9));
sram_cell_6t_5 inst_cell_9_27 (.BL(BL27),.BLN(BLN27),.WL(WL9));
sram_cell_6t_5 inst_cell_9_28 (.BL(BL28),.BLN(BLN28),.WL(WL9));
sram_cell_6t_5 inst_cell_9_29 (.BL(BL29),.BLN(BLN29),.WL(WL9));
sram_cell_6t_5 inst_cell_9_30 (.BL(BL30),.BLN(BLN30),.WL(WL9));
sram_cell_6t_5 inst_cell_9_31 (.BL(BL31),.BLN(BLN31),.WL(WL9));
sram_cell_6t_5 inst_cell_9_32 (.BL(BL32),.BLN(BLN32),.WL(WL9));
sram_cell_6t_5 inst_cell_9_33 (.BL(BL33),.BLN(BLN33),.WL(WL9));
sram_cell_6t_5 inst_cell_9_34 (.BL(BL34),.BLN(BLN34),.WL(WL9));
sram_cell_6t_5 inst_cell_9_35 (.BL(BL35),.BLN(BLN35),.WL(WL9));
sram_cell_6t_5 inst_cell_9_36 (.BL(BL36),.BLN(BLN36),.WL(WL9));
sram_cell_6t_5 inst_cell_9_37 (.BL(BL37),.BLN(BLN37),.WL(WL9));
sram_cell_6t_5 inst_cell_9_38 (.BL(BL38),.BLN(BLN38),.WL(WL9));
sram_cell_6t_5 inst_cell_9_39 (.BL(BL39),.BLN(BLN39),.WL(WL9));
sram_cell_6t_5 inst_cell_9_40 (.BL(BL40),.BLN(BLN40),.WL(WL9));
sram_cell_6t_5 inst_cell_9_41 (.BL(BL41),.BLN(BLN41),.WL(WL9));
sram_cell_6t_5 inst_cell_9_42 (.BL(BL42),.BLN(BLN42),.WL(WL9));
sram_cell_6t_5 inst_cell_9_43 (.BL(BL43),.BLN(BLN43),.WL(WL9));
sram_cell_6t_5 inst_cell_9_44 (.BL(BL44),.BLN(BLN44),.WL(WL9));
sram_cell_6t_5 inst_cell_9_45 (.BL(BL45),.BLN(BLN45),.WL(WL9));
sram_cell_6t_5 inst_cell_9_46 (.BL(BL46),.BLN(BLN46),.WL(WL9));
sram_cell_6t_5 inst_cell_9_47 (.BL(BL47),.BLN(BLN47),.WL(WL9));
sram_cell_6t_5 inst_cell_9_48 (.BL(BL48),.BLN(BLN48),.WL(WL9));
sram_cell_6t_5 inst_cell_9_49 (.BL(BL49),.BLN(BLN49),.WL(WL9));
sram_cell_6t_5 inst_cell_9_50 (.BL(BL50),.BLN(BLN50),.WL(WL9));
sram_cell_6t_5 inst_cell_9_51 (.BL(BL51),.BLN(BLN51),.WL(WL9));
sram_cell_6t_5 inst_cell_9_52 (.BL(BL52),.BLN(BLN52),.WL(WL9));
sram_cell_6t_5 inst_cell_9_53 (.BL(BL53),.BLN(BLN53),.WL(WL9));
sram_cell_6t_5 inst_cell_9_54 (.BL(BL54),.BLN(BLN54),.WL(WL9));
sram_cell_6t_5 inst_cell_9_55 (.BL(BL55),.BLN(BLN55),.WL(WL9));
sram_cell_6t_5 inst_cell_9_56 (.BL(BL56),.BLN(BLN56),.WL(WL9));
sram_cell_6t_5 inst_cell_9_57 (.BL(BL57),.BLN(BLN57),.WL(WL9));
sram_cell_6t_5 inst_cell_9_58 (.BL(BL58),.BLN(BLN58),.WL(WL9));
sram_cell_6t_5 inst_cell_9_59 (.BL(BL59),.BLN(BLN59),.WL(WL9));
sram_cell_6t_5 inst_cell_9_60 (.BL(BL60),.BLN(BLN60),.WL(WL9));
sram_cell_6t_5 inst_cell_9_61 (.BL(BL61),.BLN(BLN61),.WL(WL9));
sram_cell_6t_5 inst_cell_9_62 (.BL(BL62),.BLN(BLN62),.WL(WL9));
sram_cell_6t_5 inst_cell_9_63 (.BL(BL63),.BLN(BLN63),.WL(WL9));
sram_cell_6t_5 inst_cell_9_64 (.BL(BL64),.BLN(BLN64),.WL(WL9));
sram_cell_6t_5 inst_cell_9_65 (.BL(BL65),.BLN(BLN65),.WL(WL9));
sram_cell_6t_5 inst_cell_9_66 (.BL(BL66),.BLN(BLN66),.WL(WL9));
sram_cell_6t_5 inst_cell_9_67 (.BL(BL67),.BLN(BLN67),.WL(WL9));
sram_cell_6t_5 inst_cell_9_68 (.BL(BL68),.BLN(BLN68),.WL(WL9));
sram_cell_6t_5 inst_cell_9_69 (.BL(BL69),.BLN(BLN69),.WL(WL9));
sram_cell_6t_5 inst_cell_9_70 (.BL(BL70),.BLN(BLN70),.WL(WL9));
sram_cell_6t_5 inst_cell_9_71 (.BL(BL71),.BLN(BLN71),.WL(WL9));
sram_cell_6t_5 inst_cell_9_72 (.BL(BL72),.BLN(BLN72),.WL(WL9));
sram_cell_6t_5 inst_cell_9_73 (.BL(BL73),.BLN(BLN73),.WL(WL9));
sram_cell_6t_5 inst_cell_9_74 (.BL(BL74),.BLN(BLN74),.WL(WL9));
sram_cell_6t_5 inst_cell_9_75 (.BL(BL75),.BLN(BLN75),.WL(WL9));
sram_cell_6t_5 inst_cell_9_76 (.BL(BL76),.BLN(BLN76),.WL(WL9));
sram_cell_6t_5 inst_cell_9_77 (.BL(BL77),.BLN(BLN77),.WL(WL9));
sram_cell_6t_5 inst_cell_9_78 (.BL(BL78),.BLN(BLN78),.WL(WL9));
sram_cell_6t_5 inst_cell_9_79 (.BL(BL79),.BLN(BLN79),.WL(WL9));
sram_cell_6t_5 inst_cell_9_80 (.BL(BL80),.BLN(BLN80),.WL(WL9));
sram_cell_6t_5 inst_cell_9_81 (.BL(BL81),.BLN(BLN81),.WL(WL9));
sram_cell_6t_5 inst_cell_9_82 (.BL(BL82),.BLN(BLN82),.WL(WL9));
sram_cell_6t_5 inst_cell_9_83 (.BL(BL83),.BLN(BLN83),.WL(WL9));
sram_cell_6t_5 inst_cell_9_84 (.BL(BL84),.BLN(BLN84),.WL(WL9));
sram_cell_6t_5 inst_cell_9_85 (.BL(BL85),.BLN(BLN85),.WL(WL9));
sram_cell_6t_5 inst_cell_9_86 (.BL(BL86),.BLN(BLN86),.WL(WL9));
sram_cell_6t_5 inst_cell_9_87 (.BL(BL87),.BLN(BLN87),.WL(WL9));
sram_cell_6t_5 inst_cell_9_88 (.BL(BL88),.BLN(BLN88),.WL(WL9));
sram_cell_6t_5 inst_cell_9_89 (.BL(BL89),.BLN(BLN89),.WL(WL9));
sram_cell_6t_5 inst_cell_9_90 (.BL(BL90),.BLN(BLN90),.WL(WL9));
sram_cell_6t_5 inst_cell_9_91 (.BL(BL91),.BLN(BLN91),.WL(WL9));
sram_cell_6t_5 inst_cell_9_92 (.BL(BL92),.BLN(BLN92),.WL(WL9));
sram_cell_6t_5 inst_cell_9_93 (.BL(BL93),.BLN(BLN93),.WL(WL9));
sram_cell_6t_5 inst_cell_9_94 (.BL(BL94),.BLN(BLN94),.WL(WL9));
sram_cell_6t_5 inst_cell_9_95 (.BL(BL95),.BLN(BLN95),.WL(WL9));
sram_cell_6t_5 inst_cell_9_96 (.BL(BL96),.BLN(BLN96),.WL(WL9));
sram_cell_6t_5 inst_cell_9_97 (.BL(BL97),.BLN(BLN97),.WL(WL9));
sram_cell_6t_5 inst_cell_9_98 (.BL(BL98),.BLN(BLN98),.WL(WL9));
sram_cell_6t_5 inst_cell_9_99 (.BL(BL99),.BLN(BLN99),.WL(WL9));
sram_cell_6t_5 inst_cell_9_100 (.BL(BL100),.BLN(BLN100),.WL(WL9));
sram_cell_6t_5 inst_cell_9_101 (.BL(BL101),.BLN(BLN101),.WL(WL9));
sram_cell_6t_5 inst_cell_9_102 (.BL(BL102),.BLN(BLN102),.WL(WL9));
sram_cell_6t_5 inst_cell_9_103 (.BL(BL103),.BLN(BLN103),.WL(WL9));
sram_cell_6t_5 inst_cell_9_104 (.BL(BL104),.BLN(BLN104),.WL(WL9));
sram_cell_6t_5 inst_cell_9_105 (.BL(BL105),.BLN(BLN105),.WL(WL9));
sram_cell_6t_5 inst_cell_9_106 (.BL(BL106),.BLN(BLN106),.WL(WL9));
sram_cell_6t_5 inst_cell_9_107 (.BL(BL107),.BLN(BLN107),.WL(WL9));
sram_cell_6t_5 inst_cell_9_108 (.BL(BL108),.BLN(BLN108),.WL(WL9));
sram_cell_6t_5 inst_cell_9_109 (.BL(BL109),.BLN(BLN109),.WL(WL9));
sram_cell_6t_5 inst_cell_9_110 (.BL(BL110),.BLN(BLN110),.WL(WL9));
sram_cell_6t_5 inst_cell_9_111 (.BL(BL111),.BLN(BLN111),.WL(WL9));
sram_cell_6t_5 inst_cell_9_112 (.BL(BL112),.BLN(BLN112),.WL(WL9));
sram_cell_6t_5 inst_cell_9_113 (.BL(BL113),.BLN(BLN113),.WL(WL9));
sram_cell_6t_5 inst_cell_9_114 (.BL(BL114),.BLN(BLN114),.WL(WL9));
sram_cell_6t_5 inst_cell_9_115 (.BL(BL115),.BLN(BLN115),.WL(WL9));
sram_cell_6t_5 inst_cell_9_116 (.BL(BL116),.BLN(BLN116),.WL(WL9));
sram_cell_6t_5 inst_cell_9_117 (.BL(BL117),.BLN(BLN117),.WL(WL9));
sram_cell_6t_5 inst_cell_9_118 (.BL(BL118),.BLN(BLN118),.WL(WL9));
sram_cell_6t_5 inst_cell_9_119 (.BL(BL119),.BLN(BLN119),.WL(WL9));
sram_cell_6t_5 inst_cell_9_120 (.BL(BL120),.BLN(BLN120),.WL(WL9));
sram_cell_6t_5 inst_cell_9_121 (.BL(BL121),.BLN(BLN121),.WL(WL9));
sram_cell_6t_5 inst_cell_9_122 (.BL(BL122),.BLN(BLN122),.WL(WL9));
sram_cell_6t_5 inst_cell_9_123 (.BL(BL123),.BLN(BLN123),.WL(WL9));
sram_cell_6t_5 inst_cell_9_124 (.BL(BL124),.BLN(BLN124),.WL(WL9));
sram_cell_6t_5 inst_cell_9_125 (.BL(BL125),.BLN(BLN125),.WL(WL9));
sram_cell_6t_5 inst_cell_9_126 (.BL(BL126),.BLN(BLN126),.WL(WL9));
sram_cell_6t_5 inst_cell_9_127 (.BL(BL127),.BLN(BLN127),.WL(WL9));
sram_cell_6t_5 inst_cell_10_0 (.BL(BL0),.BLN(BLN0),.WL(WL10));
sram_cell_6t_5 inst_cell_10_1 (.BL(BL1),.BLN(BLN1),.WL(WL10));
sram_cell_6t_5 inst_cell_10_2 (.BL(BL2),.BLN(BLN2),.WL(WL10));
sram_cell_6t_5 inst_cell_10_3 (.BL(BL3),.BLN(BLN3),.WL(WL10));
sram_cell_6t_5 inst_cell_10_4 (.BL(BL4),.BLN(BLN4),.WL(WL10));
sram_cell_6t_5 inst_cell_10_5 (.BL(BL5),.BLN(BLN5),.WL(WL10));
sram_cell_6t_5 inst_cell_10_6 (.BL(BL6),.BLN(BLN6),.WL(WL10));
sram_cell_6t_5 inst_cell_10_7 (.BL(BL7),.BLN(BLN7),.WL(WL10));
sram_cell_6t_5 inst_cell_10_8 (.BL(BL8),.BLN(BLN8),.WL(WL10));
sram_cell_6t_5 inst_cell_10_9 (.BL(BL9),.BLN(BLN9),.WL(WL10));
sram_cell_6t_5 inst_cell_10_10 (.BL(BL10),.BLN(BLN10),.WL(WL10));
sram_cell_6t_5 inst_cell_10_11 (.BL(BL11),.BLN(BLN11),.WL(WL10));
sram_cell_6t_5 inst_cell_10_12 (.BL(BL12),.BLN(BLN12),.WL(WL10));
sram_cell_6t_5 inst_cell_10_13 (.BL(BL13),.BLN(BLN13),.WL(WL10));
sram_cell_6t_5 inst_cell_10_14 (.BL(BL14),.BLN(BLN14),.WL(WL10));
sram_cell_6t_5 inst_cell_10_15 (.BL(BL15),.BLN(BLN15),.WL(WL10));
sram_cell_6t_5 inst_cell_10_16 (.BL(BL16),.BLN(BLN16),.WL(WL10));
sram_cell_6t_5 inst_cell_10_17 (.BL(BL17),.BLN(BLN17),.WL(WL10));
sram_cell_6t_5 inst_cell_10_18 (.BL(BL18),.BLN(BLN18),.WL(WL10));
sram_cell_6t_5 inst_cell_10_19 (.BL(BL19),.BLN(BLN19),.WL(WL10));
sram_cell_6t_5 inst_cell_10_20 (.BL(BL20),.BLN(BLN20),.WL(WL10));
sram_cell_6t_5 inst_cell_10_21 (.BL(BL21),.BLN(BLN21),.WL(WL10));
sram_cell_6t_5 inst_cell_10_22 (.BL(BL22),.BLN(BLN22),.WL(WL10));
sram_cell_6t_5 inst_cell_10_23 (.BL(BL23),.BLN(BLN23),.WL(WL10));
sram_cell_6t_5 inst_cell_10_24 (.BL(BL24),.BLN(BLN24),.WL(WL10));
sram_cell_6t_5 inst_cell_10_25 (.BL(BL25),.BLN(BLN25),.WL(WL10));
sram_cell_6t_5 inst_cell_10_26 (.BL(BL26),.BLN(BLN26),.WL(WL10));
sram_cell_6t_5 inst_cell_10_27 (.BL(BL27),.BLN(BLN27),.WL(WL10));
sram_cell_6t_5 inst_cell_10_28 (.BL(BL28),.BLN(BLN28),.WL(WL10));
sram_cell_6t_5 inst_cell_10_29 (.BL(BL29),.BLN(BLN29),.WL(WL10));
sram_cell_6t_5 inst_cell_10_30 (.BL(BL30),.BLN(BLN30),.WL(WL10));
sram_cell_6t_5 inst_cell_10_31 (.BL(BL31),.BLN(BLN31),.WL(WL10));
sram_cell_6t_5 inst_cell_10_32 (.BL(BL32),.BLN(BLN32),.WL(WL10));
sram_cell_6t_5 inst_cell_10_33 (.BL(BL33),.BLN(BLN33),.WL(WL10));
sram_cell_6t_5 inst_cell_10_34 (.BL(BL34),.BLN(BLN34),.WL(WL10));
sram_cell_6t_5 inst_cell_10_35 (.BL(BL35),.BLN(BLN35),.WL(WL10));
sram_cell_6t_5 inst_cell_10_36 (.BL(BL36),.BLN(BLN36),.WL(WL10));
sram_cell_6t_5 inst_cell_10_37 (.BL(BL37),.BLN(BLN37),.WL(WL10));
sram_cell_6t_5 inst_cell_10_38 (.BL(BL38),.BLN(BLN38),.WL(WL10));
sram_cell_6t_5 inst_cell_10_39 (.BL(BL39),.BLN(BLN39),.WL(WL10));
sram_cell_6t_5 inst_cell_10_40 (.BL(BL40),.BLN(BLN40),.WL(WL10));
sram_cell_6t_5 inst_cell_10_41 (.BL(BL41),.BLN(BLN41),.WL(WL10));
sram_cell_6t_5 inst_cell_10_42 (.BL(BL42),.BLN(BLN42),.WL(WL10));
sram_cell_6t_5 inst_cell_10_43 (.BL(BL43),.BLN(BLN43),.WL(WL10));
sram_cell_6t_5 inst_cell_10_44 (.BL(BL44),.BLN(BLN44),.WL(WL10));
sram_cell_6t_5 inst_cell_10_45 (.BL(BL45),.BLN(BLN45),.WL(WL10));
sram_cell_6t_5 inst_cell_10_46 (.BL(BL46),.BLN(BLN46),.WL(WL10));
sram_cell_6t_5 inst_cell_10_47 (.BL(BL47),.BLN(BLN47),.WL(WL10));
sram_cell_6t_5 inst_cell_10_48 (.BL(BL48),.BLN(BLN48),.WL(WL10));
sram_cell_6t_5 inst_cell_10_49 (.BL(BL49),.BLN(BLN49),.WL(WL10));
sram_cell_6t_5 inst_cell_10_50 (.BL(BL50),.BLN(BLN50),.WL(WL10));
sram_cell_6t_5 inst_cell_10_51 (.BL(BL51),.BLN(BLN51),.WL(WL10));
sram_cell_6t_5 inst_cell_10_52 (.BL(BL52),.BLN(BLN52),.WL(WL10));
sram_cell_6t_5 inst_cell_10_53 (.BL(BL53),.BLN(BLN53),.WL(WL10));
sram_cell_6t_5 inst_cell_10_54 (.BL(BL54),.BLN(BLN54),.WL(WL10));
sram_cell_6t_5 inst_cell_10_55 (.BL(BL55),.BLN(BLN55),.WL(WL10));
sram_cell_6t_5 inst_cell_10_56 (.BL(BL56),.BLN(BLN56),.WL(WL10));
sram_cell_6t_5 inst_cell_10_57 (.BL(BL57),.BLN(BLN57),.WL(WL10));
sram_cell_6t_5 inst_cell_10_58 (.BL(BL58),.BLN(BLN58),.WL(WL10));
sram_cell_6t_5 inst_cell_10_59 (.BL(BL59),.BLN(BLN59),.WL(WL10));
sram_cell_6t_5 inst_cell_10_60 (.BL(BL60),.BLN(BLN60),.WL(WL10));
sram_cell_6t_5 inst_cell_10_61 (.BL(BL61),.BLN(BLN61),.WL(WL10));
sram_cell_6t_5 inst_cell_10_62 (.BL(BL62),.BLN(BLN62),.WL(WL10));
sram_cell_6t_5 inst_cell_10_63 (.BL(BL63),.BLN(BLN63),.WL(WL10));
sram_cell_6t_5 inst_cell_10_64 (.BL(BL64),.BLN(BLN64),.WL(WL10));
sram_cell_6t_5 inst_cell_10_65 (.BL(BL65),.BLN(BLN65),.WL(WL10));
sram_cell_6t_5 inst_cell_10_66 (.BL(BL66),.BLN(BLN66),.WL(WL10));
sram_cell_6t_5 inst_cell_10_67 (.BL(BL67),.BLN(BLN67),.WL(WL10));
sram_cell_6t_5 inst_cell_10_68 (.BL(BL68),.BLN(BLN68),.WL(WL10));
sram_cell_6t_5 inst_cell_10_69 (.BL(BL69),.BLN(BLN69),.WL(WL10));
sram_cell_6t_5 inst_cell_10_70 (.BL(BL70),.BLN(BLN70),.WL(WL10));
sram_cell_6t_5 inst_cell_10_71 (.BL(BL71),.BLN(BLN71),.WL(WL10));
sram_cell_6t_5 inst_cell_10_72 (.BL(BL72),.BLN(BLN72),.WL(WL10));
sram_cell_6t_5 inst_cell_10_73 (.BL(BL73),.BLN(BLN73),.WL(WL10));
sram_cell_6t_5 inst_cell_10_74 (.BL(BL74),.BLN(BLN74),.WL(WL10));
sram_cell_6t_5 inst_cell_10_75 (.BL(BL75),.BLN(BLN75),.WL(WL10));
sram_cell_6t_5 inst_cell_10_76 (.BL(BL76),.BLN(BLN76),.WL(WL10));
sram_cell_6t_5 inst_cell_10_77 (.BL(BL77),.BLN(BLN77),.WL(WL10));
sram_cell_6t_5 inst_cell_10_78 (.BL(BL78),.BLN(BLN78),.WL(WL10));
sram_cell_6t_5 inst_cell_10_79 (.BL(BL79),.BLN(BLN79),.WL(WL10));
sram_cell_6t_5 inst_cell_10_80 (.BL(BL80),.BLN(BLN80),.WL(WL10));
sram_cell_6t_5 inst_cell_10_81 (.BL(BL81),.BLN(BLN81),.WL(WL10));
sram_cell_6t_5 inst_cell_10_82 (.BL(BL82),.BLN(BLN82),.WL(WL10));
sram_cell_6t_5 inst_cell_10_83 (.BL(BL83),.BLN(BLN83),.WL(WL10));
sram_cell_6t_5 inst_cell_10_84 (.BL(BL84),.BLN(BLN84),.WL(WL10));
sram_cell_6t_5 inst_cell_10_85 (.BL(BL85),.BLN(BLN85),.WL(WL10));
sram_cell_6t_5 inst_cell_10_86 (.BL(BL86),.BLN(BLN86),.WL(WL10));
sram_cell_6t_5 inst_cell_10_87 (.BL(BL87),.BLN(BLN87),.WL(WL10));
sram_cell_6t_5 inst_cell_10_88 (.BL(BL88),.BLN(BLN88),.WL(WL10));
sram_cell_6t_5 inst_cell_10_89 (.BL(BL89),.BLN(BLN89),.WL(WL10));
sram_cell_6t_5 inst_cell_10_90 (.BL(BL90),.BLN(BLN90),.WL(WL10));
sram_cell_6t_5 inst_cell_10_91 (.BL(BL91),.BLN(BLN91),.WL(WL10));
sram_cell_6t_5 inst_cell_10_92 (.BL(BL92),.BLN(BLN92),.WL(WL10));
sram_cell_6t_5 inst_cell_10_93 (.BL(BL93),.BLN(BLN93),.WL(WL10));
sram_cell_6t_5 inst_cell_10_94 (.BL(BL94),.BLN(BLN94),.WL(WL10));
sram_cell_6t_5 inst_cell_10_95 (.BL(BL95),.BLN(BLN95),.WL(WL10));
sram_cell_6t_5 inst_cell_10_96 (.BL(BL96),.BLN(BLN96),.WL(WL10));
sram_cell_6t_5 inst_cell_10_97 (.BL(BL97),.BLN(BLN97),.WL(WL10));
sram_cell_6t_5 inst_cell_10_98 (.BL(BL98),.BLN(BLN98),.WL(WL10));
sram_cell_6t_5 inst_cell_10_99 (.BL(BL99),.BLN(BLN99),.WL(WL10));
sram_cell_6t_5 inst_cell_10_100 (.BL(BL100),.BLN(BLN100),.WL(WL10));
sram_cell_6t_5 inst_cell_10_101 (.BL(BL101),.BLN(BLN101),.WL(WL10));
sram_cell_6t_5 inst_cell_10_102 (.BL(BL102),.BLN(BLN102),.WL(WL10));
sram_cell_6t_5 inst_cell_10_103 (.BL(BL103),.BLN(BLN103),.WL(WL10));
sram_cell_6t_5 inst_cell_10_104 (.BL(BL104),.BLN(BLN104),.WL(WL10));
sram_cell_6t_5 inst_cell_10_105 (.BL(BL105),.BLN(BLN105),.WL(WL10));
sram_cell_6t_5 inst_cell_10_106 (.BL(BL106),.BLN(BLN106),.WL(WL10));
sram_cell_6t_5 inst_cell_10_107 (.BL(BL107),.BLN(BLN107),.WL(WL10));
sram_cell_6t_5 inst_cell_10_108 (.BL(BL108),.BLN(BLN108),.WL(WL10));
sram_cell_6t_5 inst_cell_10_109 (.BL(BL109),.BLN(BLN109),.WL(WL10));
sram_cell_6t_5 inst_cell_10_110 (.BL(BL110),.BLN(BLN110),.WL(WL10));
sram_cell_6t_5 inst_cell_10_111 (.BL(BL111),.BLN(BLN111),.WL(WL10));
sram_cell_6t_5 inst_cell_10_112 (.BL(BL112),.BLN(BLN112),.WL(WL10));
sram_cell_6t_5 inst_cell_10_113 (.BL(BL113),.BLN(BLN113),.WL(WL10));
sram_cell_6t_5 inst_cell_10_114 (.BL(BL114),.BLN(BLN114),.WL(WL10));
sram_cell_6t_5 inst_cell_10_115 (.BL(BL115),.BLN(BLN115),.WL(WL10));
sram_cell_6t_5 inst_cell_10_116 (.BL(BL116),.BLN(BLN116),.WL(WL10));
sram_cell_6t_5 inst_cell_10_117 (.BL(BL117),.BLN(BLN117),.WL(WL10));
sram_cell_6t_5 inst_cell_10_118 (.BL(BL118),.BLN(BLN118),.WL(WL10));
sram_cell_6t_5 inst_cell_10_119 (.BL(BL119),.BLN(BLN119),.WL(WL10));
sram_cell_6t_5 inst_cell_10_120 (.BL(BL120),.BLN(BLN120),.WL(WL10));
sram_cell_6t_5 inst_cell_10_121 (.BL(BL121),.BLN(BLN121),.WL(WL10));
sram_cell_6t_5 inst_cell_10_122 (.BL(BL122),.BLN(BLN122),.WL(WL10));
sram_cell_6t_5 inst_cell_10_123 (.BL(BL123),.BLN(BLN123),.WL(WL10));
sram_cell_6t_5 inst_cell_10_124 (.BL(BL124),.BLN(BLN124),.WL(WL10));
sram_cell_6t_5 inst_cell_10_125 (.BL(BL125),.BLN(BLN125),.WL(WL10));
sram_cell_6t_5 inst_cell_10_126 (.BL(BL126),.BLN(BLN126),.WL(WL10));
sram_cell_6t_5 inst_cell_10_127 (.BL(BL127),.BLN(BLN127),.WL(WL10));
sram_cell_6t_5 inst_cell_11_0 (.BL(BL0),.BLN(BLN0),.WL(WL11));
sram_cell_6t_5 inst_cell_11_1 (.BL(BL1),.BLN(BLN1),.WL(WL11));
sram_cell_6t_5 inst_cell_11_2 (.BL(BL2),.BLN(BLN2),.WL(WL11));
sram_cell_6t_5 inst_cell_11_3 (.BL(BL3),.BLN(BLN3),.WL(WL11));
sram_cell_6t_5 inst_cell_11_4 (.BL(BL4),.BLN(BLN4),.WL(WL11));
sram_cell_6t_5 inst_cell_11_5 (.BL(BL5),.BLN(BLN5),.WL(WL11));
sram_cell_6t_5 inst_cell_11_6 (.BL(BL6),.BLN(BLN6),.WL(WL11));
sram_cell_6t_5 inst_cell_11_7 (.BL(BL7),.BLN(BLN7),.WL(WL11));
sram_cell_6t_5 inst_cell_11_8 (.BL(BL8),.BLN(BLN8),.WL(WL11));
sram_cell_6t_5 inst_cell_11_9 (.BL(BL9),.BLN(BLN9),.WL(WL11));
sram_cell_6t_5 inst_cell_11_10 (.BL(BL10),.BLN(BLN10),.WL(WL11));
sram_cell_6t_5 inst_cell_11_11 (.BL(BL11),.BLN(BLN11),.WL(WL11));
sram_cell_6t_5 inst_cell_11_12 (.BL(BL12),.BLN(BLN12),.WL(WL11));
sram_cell_6t_5 inst_cell_11_13 (.BL(BL13),.BLN(BLN13),.WL(WL11));
sram_cell_6t_5 inst_cell_11_14 (.BL(BL14),.BLN(BLN14),.WL(WL11));
sram_cell_6t_5 inst_cell_11_15 (.BL(BL15),.BLN(BLN15),.WL(WL11));
sram_cell_6t_5 inst_cell_11_16 (.BL(BL16),.BLN(BLN16),.WL(WL11));
sram_cell_6t_5 inst_cell_11_17 (.BL(BL17),.BLN(BLN17),.WL(WL11));
sram_cell_6t_5 inst_cell_11_18 (.BL(BL18),.BLN(BLN18),.WL(WL11));
sram_cell_6t_5 inst_cell_11_19 (.BL(BL19),.BLN(BLN19),.WL(WL11));
sram_cell_6t_5 inst_cell_11_20 (.BL(BL20),.BLN(BLN20),.WL(WL11));
sram_cell_6t_5 inst_cell_11_21 (.BL(BL21),.BLN(BLN21),.WL(WL11));
sram_cell_6t_5 inst_cell_11_22 (.BL(BL22),.BLN(BLN22),.WL(WL11));
sram_cell_6t_5 inst_cell_11_23 (.BL(BL23),.BLN(BLN23),.WL(WL11));
sram_cell_6t_5 inst_cell_11_24 (.BL(BL24),.BLN(BLN24),.WL(WL11));
sram_cell_6t_5 inst_cell_11_25 (.BL(BL25),.BLN(BLN25),.WL(WL11));
sram_cell_6t_5 inst_cell_11_26 (.BL(BL26),.BLN(BLN26),.WL(WL11));
sram_cell_6t_5 inst_cell_11_27 (.BL(BL27),.BLN(BLN27),.WL(WL11));
sram_cell_6t_5 inst_cell_11_28 (.BL(BL28),.BLN(BLN28),.WL(WL11));
sram_cell_6t_5 inst_cell_11_29 (.BL(BL29),.BLN(BLN29),.WL(WL11));
sram_cell_6t_5 inst_cell_11_30 (.BL(BL30),.BLN(BLN30),.WL(WL11));
sram_cell_6t_5 inst_cell_11_31 (.BL(BL31),.BLN(BLN31),.WL(WL11));
sram_cell_6t_5 inst_cell_11_32 (.BL(BL32),.BLN(BLN32),.WL(WL11));
sram_cell_6t_5 inst_cell_11_33 (.BL(BL33),.BLN(BLN33),.WL(WL11));
sram_cell_6t_5 inst_cell_11_34 (.BL(BL34),.BLN(BLN34),.WL(WL11));
sram_cell_6t_5 inst_cell_11_35 (.BL(BL35),.BLN(BLN35),.WL(WL11));
sram_cell_6t_5 inst_cell_11_36 (.BL(BL36),.BLN(BLN36),.WL(WL11));
sram_cell_6t_5 inst_cell_11_37 (.BL(BL37),.BLN(BLN37),.WL(WL11));
sram_cell_6t_5 inst_cell_11_38 (.BL(BL38),.BLN(BLN38),.WL(WL11));
sram_cell_6t_5 inst_cell_11_39 (.BL(BL39),.BLN(BLN39),.WL(WL11));
sram_cell_6t_5 inst_cell_11_40 (.BL(BL40),.BLN(BLN40),.WL(WL11));
sram_cell_6t_5 inst_cell_11_41 (.BL(BL41),.BLN(BLN41),.WL(WL11));
sram_cell_6t_5 inst_cell_11_42 (.BL(BL42),.BLN(BLN42),.WL(WL11));
sram_cell_6t_5 inst_cell_11_43 (.BL(BL43),.BLN(BLN43),.WL(WL11));
sram_cell_6t_5 inst_cell_11_44 (.BL(BL44),.BLN(BLN44),.WL(WL11));
sram_cell_6t_5 inst_cell_11_45 (.BL(BL45),.BLN(BLN45),.WL(WL11));
sram_cell_6t_5 inst_cell_11_46 (.BL(BL46),.BLN(BLN46),.WL(WL11));
sram_cell_6t_5 inst_cell_11_47 (.BL(BL47),.BLN(BLN47),.WL(WL11));
sram_cell_6t_5 inst_cell_11_48 (.BL(BL48),.BLN(BLN48),.WL(WL11));
sram_cell_6t_5 inst_cell_11_49 (.BL(BL49),.BLN(BLN49),.WL(WL11));
sram_cell_6t_5 inst_cell_11_50 (.BL(BL50),.BLN(BLN50),.WL(WL11));
sram_cell_6t_5 inst_cell_11_51 (.BL(BL51),.BLN(BLN51),.WL(WL11));
sram_cell_6t_5 inst_cell_11_52 (.BL(BL52),.BLN(BLN52),.WL(WL11));
sram_cell_6t_5 inst_cell_11_53 (.BL(BL53),.BLN(BLN53),.WL(WL11));
sram_cell_6t_5 inst_cell_11_54 (.BL(BL54),.BLN(BLN54),.WL(WL11));
sram_cell_6t_5 inst_cell_11_55 (.BL(BL55),.BLN(BLN55),.WL(WL11));
sram_cell_6t_5 inst_cell_11_56 (.BL(BL56),.BLN(BLN56),.WL(WL11));
sram_cell_6t_5 inst_cell_11_57 (.BL(BL57),.BLN(BLN57),.WL(WL11));
sram_cell_6t_5 inst_cell_11_58 (.BL(BL58),.BLN(BLN58),.WL(WL11));
sram_cell_6t_5 inst_cell_11_59 (.BL(BL59),.BLN(BLN59),.WL(WL11));
sram_cell_6t_5 inst_cell_11_60 (.BL(BL60),.BLN(BLN60),.WL(WL11));
sram_cell_6t_5 inst_cell_11_61 (.BL(BL61),.BLN(BLN61),.WL(WL11));
sram_cell_6t_5 inst_cell_11_62 (.BL(BL62),.BLN(BLN62),.WL(WL11));
sram_cell_6t_5 inst_cell_11_63 (.BL(BL63),.BLN(BLN63),.WL(WL11));
sram_cell_6t_5 inst_cell_11_64 (.BL(BL64),.BLN(BLN64),.WL(WL11));
sram_cell_6t_5 inst_cell_11_65 (.BL(BL65),.BLN(BLN65),.WL(WL11));
sram_cell_6t_5 inst_cell_11_66 (.BL(BL66),.BLN(BLN66),.WL(WL11));
sram_cell_6t_5 inst_cell_11_67 (.BL(BL67),.BLN(BLN67),.WL(WL11));
sram_cell_6t_5 inst_cell_11_68 (.BL(BL68),.BLN(BLN68),.WL(WL11));
sram_cell_6t_5 inst_cell_11_69 (.BL(BL69),.BLN(BLN69),.WL(WL11));
sram_cell_6t_5 inst_cell_11_70 (.BL(BL70),.BLN(BLN70),.WL(WL11));
sram_cell_6t_5 inst_cell_11_71 (.BL(BL71),.BLN(BLN71),.WL(WL11));
sram_cell_6t_5 inst_cell_11_72 (.BL(BL72),.BLN(BLN72),.WL(WL11));
sram_cell_6t_5 inst_cell_11_73 (.BL(BL73),.BLN(BLN73),.WL(WL11));
sram_cell_6t_5 inst_cell_11_74 (.BL(BL74),.BLN(BLN74),.WL(WL11));
sram_cell_6t_5 inst_cell_11_75 (.BL(BL75),.BLN(BLN75),.WL(WL11));
sram_cell_6t_5 inst_cell_11_76 (.BL(BL76),.BLN(BLN76),.WL(WL11));
sram_cell_6t_5 inst_cell_11_77 (.BL(BL77),.BLN(BLN77),.WL(WL11));
sram_cell_6t_5 inst_cell_11_78 (.BL(BL78),.BLN(BLN78),.WL(WL11));
sram_cell_6t_5 inst_cell_11_79 (.BL(BL79),.BLN(BLN79),.WL(WL11));
sram_cell_6t_5 inst_cell_11_80 (.BL(BL80),.BLN(BLN80),.WL(WL11));
sram_cell_6t_5 inst_cell_11_81 (.BL(BL81),.BLN(BLN81),.WL(WL11));
sram_cell_6t_5 inst_cell_11_82 (.BL(BL82),.BLN(BLN82),.WL(WL11));
sram_cell_6t_5 inst_cell_11_83 (.BL(BL83),.BLN(BLN83),.WL(WL11));
sram_cell_6t_5 inst_cell_11_84 (.BL(BL84),.BLN(BLN84),.WL(WL11));
sram_cell_6t_5 inst_cell_11_85 (.BL(BL85),.BLN(BLN85),.WL(WL11));
sram_cell_6t_5 inst_cell_11_86 (.BL(BL86),.BLN(BLN86),.WL(WL11));
sram_cell_6t_5 inst_cell_11_87 (.BL(BL87),.BLN(BLN87),.WL(WL11));
sram_cell_6t_5 inst_cell_11_88 (.BL(BL88),.BLN(BLN88),.WL(WL11));
sram_cell_6t_5 inst_cell_11_89 (.BL(BL89),.BLN(BLN89),.WL(WL11));
sram_cell_6t_5 inst_cell_11_90 (.BL(BL90),.BLN(BLN90),.WL(WL11));
sram_cell_6t_5 inst_cell_11_91 (.BL(BL91),.BLN(BLN91),.WL(WL11));
sram_cell_6t_5 inst_cell_11_92 (.BL(BL92),.BLN(BLN92),.WL(WL11));
sram_cell_6t_5 inst_cell_11_93 (.BL(BL93),.BLN(BLN93),.WL(WL11));
sram_cell_6t_5 inst_cell_11_94 (.BL(BL94),.BLN(BLN94),.WL(WL11));
sram_cell_6t_5 inst_cell_11_95 (.BL(BL95),.BLN(BLN95),.WL(WL11));
sram_cell_6t_5 inst_cell_11_96 (.BL(BL96),.BLN(BLN96),.WL(WL11));
sram_cell_6t_5 inst_cell_11_97 (.BL(BL97),.BLN(BLN97),.WL(WL11));
sram_cell_6t_5 inst_cell_11_98 (.BL(BL98),.BLN(BLN98),.WL(WL11));
sram_cell_6t_5 inst_cell_11_99 (.BL(BL99),.BLN(BLN99),.WL(WL11));
sram_cell_6t_5 inst_cell_11_100 (.BL(BL100),.BLN(BLN100),.WL(WL11));
sram_cell_6t_5 inst_cell_11_101 (.BL(BL101),.BLN(BLN101),.WL(WL11));
sram_cell_6t_5 inst_cell_11_102 (.BL(BL102),.BLN(BLN102),.WL(WL11));
sram_cell_6t_5 inst_cell_11_103 (.BL(BL103),.BLN(BLN103),.WL(WL11));
sram_cell_6t_5 inst_cell_11_104 (.BL(BL104),.BLN(BLN104),.WL(WL11));
sram_cell_6t_5 inst_cell_11_105 (.BL(BL105),.BLN(BLN105),.WL(WL11));
sram_cell_6t_5 inst_cell_11_106 (.BL(BL106),.BLN(BLN106),.WL(WL11));
sram_cell_6t_5 inst_cell_11_107 (.BL(BL107),.BLN(BLN107),.WL(WL11));
sram_cell_6t_5 inst_cell_11_108 (.BL(BL108),.BLN(BLN108),.WL(WL11));
sram_cell_6t_5 inst_cell_11_109 (.BL(BL109),.BLN(BLN109),.WL(WL11));
sram_cell_6t_5 inst_cell_11_110 (.BL(BL110),.BLN(BLN110),.WL(WL11));
sram_cell_6t_5 inst_cell_11_111 (.BL(BL111),.BLN(BLN111),.WL(WL11));
sram_cell_6t_5 inst_cell_11_112 (.BL(BL112),.BLN(BLN112),.WL(WL11));
sram_cell_6t_5 inst_cell_11_113 (.BL(BL113),.BLN(BLN113),.WL(WL11));
sram_cell_6t_5 inst_cell_11_114 (.BL(BL114),.BLN(BLN114),.WL(WL11));
sram_cell_6t_5 inst_cell_11_115 (.BL(BL115),.BLN(BLN115),.WL(WL11));
sram_cell_6t_5 inst_cell_11_116 (.BL(BL116),.BLN(BLN116),.WL(WL11));
sram_cell_6t_5 inst_cell_11_117 (.BL(BL117),.BLN(BLN117),.WL(WL11));
sram_cell_6t_5 inst_cell_11_118 (.BL(BL118),.BLN(BLN118),.WL(WL11));
sram_cell_6t_5 inst_cell_11_119 (.BL(BL119),.BLN(BLN119),.WL(WL11));
sram_cell_6t_5 inst_cell_11_120 (.BL(BL120),.BLN(BLN120),.WL(WL11));
sram_cell_6t_5 inst_cell_11_121 (.BL(BL121),.BLN(BLN121),.WL(WL11));
sram_cell_6t_5 inst_cell_11_122 (.BL(BL122),.BLN(BLN122),.WL(WL11));
sram_cell_6t_5 inst_cell_11_123 (.BL(BL123),.BLN(BLN123),.WL(WL11));
sram_cell_6t_5 inst_cell_11_124 (.BL(BL124),.BLN(BLN124),.WL(WL11));
sram_cell_6t_5 inst_cell_11_125 (.BL(BL125),.BLN(BLN125),.WL(WL11));
sram_cell_6t_5 inst_cell_11_126 (.BL(BL126),.BLN(BLN126),.WL(WL11));
sram_cell_6t_5 inst_cell_11_127 (.BL(BL127),.BLN(BLN127),.WL(WL11));
sram_cell_6t_5 inst_cell_12_0 (.BL(BL0),.BLN(BLN0),.WL(WL12));
sram_cell_6t_5 inst_cell_12_1 (.BL(BL1),.BLN(BLN1),.WL(WL12));
sram_cell_6t_5 inst_cell_12_2 (.BL(BL2),.BLN(BLN2),.WL(WL12));
sram_cell_6t_5 inst_cell_12_3 (.BL(BL3),.BLN(BLN3),.WL(WL12));
sram_cell_6t_5 inst_cell_12_4 (.BL(BL4),.BLN(BLN4),.WL(WL12));
sram_cell_6t_5 inst_cell_12_5 (.BL(BL5),.BLN(BLN5),.WL(WL12));
sram_cell_6t_5 inst_cell_12_6 (.BL(BL6),.BLN(BLN6),.WL(WL12));
sram_cell_6t_5 inst_cell_12_7 (.BL(BL7),.BLN(BLN7),.WL(WL12));
sram_cell_6t_5 inst_cell_12_8 (.BL(BL8),.BLN(BLN8),.WL(WL12));
sram_cell_6t_5 inst_cell_12_9 (.BL(BL9),.BLN(BLN9),.WL(WL12));
sram_cell_6t_5 inst_cell_12_10 (.BL(BL10),.BLN(BLN10),.WL(WL12));
sram_cell_6t_5 inst_cell_12_11 (.BL(BL11),.BLN(BLN11),.WL(WL12));
sram_cell_6t_5 inst_cell_12_12 (.BL(BL12),.BLN(BLN12),.WL(WL12));
sram_cell_6t_5 inst_cell_12_13 (.BL(BL13),.BLN(BLN13),.WL(WL12));
sram_cell_6t_5 inst_cell_12_14 (.BL(BL14),.BLN(BLN14),.WL(WL12));
sram_cell_6t_5 inst_cell_12_15 (.BL(BL15),.BLN(BLN15),.WL(WL12));
sram_cell_6t_5 inst_cell_12_16 (.BL(BL16),.BLN(BLN16),.WL(WL12));
sram_cell_6t_5 inst_cell_12_17 (.BL(BL17),.BLN(BLN17),.WL(WL12));
sram_cell_6t_5 inst_cell_12_18 (.BL(BL18),.BLN(BLN18),.WL(WL12));
sram_cell_6t_5 inst_cell_12_19 (.BL(BL19),.BLN(BLN19),.WL(WL12));
sram_cell_6t_5 inst_cell_12_20 (.BL(BL20),.BLN(BLN20),.WL(WL12));
sram_cell_6t_5 inst_cell_12_21 (.BL(BL21),.BLN(BLN21),.WL(WL12));
sram_cell_6t_5 inst_cell_12_22 (.BL(BL22),.BLN(BLN22),.WL(WL12));
sram_cell_6t_5 inst_cell_12_23 (.BL(BL23),.BLN(BLN23),.WL(WL12));
sram_cell_6t_5 inst_cell_12_24 (.BL(BL24),.BLN(BLN24),.WL(WL12));
sram_cell_6t_5 inst_cell_12_25 (.BL(BL25),.BLN(BLN25),.WL(WL12));
sram_cell_6t_5 inst_cell_12_26 (.BL(BL26),.BLN(BLN26),.WL(WL12));
sram_cell_6t_5 inst_cell_12_27 (.BL(BL27),.BLN(BLN27),.WL(WL12));
sram_cell_6t_5 inst_cell_12_28 (.BL(BL28),.BLN(BLN28),.WL(WL12));
sram_cell_6t_5 inst_cell_12_29 (.BL(BL29),.BLN(BLN29),.WL(WL12));
sram_cell_6t_5 inst_cell_12_30 (.BL(BL30),.BLN(BLN30),.WL(WL12));
sram_cell_6t_5 inst_cell_12_31 (.BL(BL31),.BLN(BLN31),.WL(WL12));
sram_cell_6t_5 inst_cell_12_32 (.BL(BL32),.BLN(BLN32),.WL(WL12));
sram_cell_6t_5 inst_cell_12_33 (.BL(BL33),.BLN(BLN33),.WL(WL12));
sram_cell_6t_5 inst_cell_12_34 (.BL(BL34),.BLN(BLN34),.WL(WL12));
sram_cell_6t_5 inst_cell_12_35 (.BL(BL35),.BLN(BLN35),.WL(WL12));
sram_cell_6t_5 inst_cell_12_36 (.BL(BL36),.BLN(BLN36),.WL(WL12));
sram_cell_6t_5 inst_cell_12_37 (.BL(BL37),.BLN(BLN37),.WL(WL12));
sram_cell_6t_5 inst_cell_12_38 (.BL(BL38),.BLN(BLN38),.WL(WL12));
sram_cell_6t_5 inst_cell_12_39 (.BL(BL39),.BLN(BLN39),.WL(WL12));
sram_cell_6t_5 inst_cell_12_40 (.BL(BL40),.BLN(BLN40),.WL(WL12));
sram_cell_6t_5 inst_cell_12_41 (.BL(BL41),.BLN(BLN41),.WL(WL12));
sram_cell_6t_5 inst_cell_12_42 (.BL(BL42),.BLN(BLN42),.WL(WL12));
sram_cell_6t_5 inst_cell_12_43 (.BL(BL43),.BLN(BLN43),.WL(WL12));
sram_cell_6t_5 inst_cell_12_44 (.BL(BL44),.BLN(BLN44),.WL(WL12));
sram_cell_6t_5 inst_cell_12_45 (.BL(BL45),.BLN(BLN45),.WL(WL12));
sram_cell_6t_5 inst_cell_12_46 (.BL(BL46),.BLN(BLN46),.WL(WL12));
sram_cell_6t_5 inst_cell_12_47 (.BL(BL47),.BLN(BLN47),.WL(WL12));
sram_cell_6t_5 inst_cell_12_48 (.BL(BL48),.BLN(BLN48),.WL(WL12));
sram_cell_6t_5 inst_cell_12_49 (.BL(BL49),.BLN(BLN49),.WL(WL12));
sram_cell_6t_5 inst_cell_12_50 (.BL(BL50),.BLN(BLN50),.WL(WL12));
sram_cell_6t_5 inst_cell_12_51 (.BL(BL51),.BLN(BLN51),.WL(WL12));
sram_cell_6t_5 inst_cell_12_52 (.BL(BL52),.BLN(BLN52),.WL(WL12));
sram_cell_6t_5 inst_cell_12_53 (.BL(BL53),.BLN(BLN53),.WL(WL12));
sram_cell_6t_5 inst_cell_12_54 (.BL(BL54),.BLN(BLN54),.WL(WL12));
sram_cell_6t_5 inst_cell_12_55 (.BL(BL55),.BLN(BLN55),.WL(WL12));
sram_cell_6t_5 inst_cell_12_56 (.BL(BL56),.BLN(BLN56),.WL(WL12));
sram_cell_6t_5 inst_cell_12_57 (.BL(BL57),.BLN(BLN57),.WL(WL12));
sram_cell_6t_5 inst_cell_12_58 (.BL(BL58),.BLN(BLN58),.WL(WL12));
sram_cell_6t_5 inst_cell_12_59 (.BL(BL59),.BLN(BLN59),.WL(WL12));
sram_cell_6t_5 inst_cell_12_60 (.BL(BL60),.BLN(BLN60),.WL(WL12));
sram_cell_6t_5 inst_cell_12_61 (.BL(BL61),.BLN(BLN61),.WL(WL12));
sram_cell_6t_5 inst_cell_12_62 (.BL(BL62),.BLN(BLN62),.WL(WL12));
sram_cell_6t_5 inst_cell_12_63 (.BL(BL63),.BLN(BLN63),.WL(WL12));
sram_cell_6t_5 inst_cell_12_64 (.BL(BL64),.BLN(BLN64),.WL(WL12));
sram_cell_6t_5 inst_cell_12_65 (.BL(BL65),.BLN(BLN65),.WL(WL12));
sram_cell_6t_5 inst_cell_12_66 (.BL(BL66),.BLN(BLN66),.WL(WL12));
sram_cell_6t_5 inst_cell_12_67 (.BL(BL67),.BLN(BLN67),.WL(WL12));
sram_cell_6t_5 inst_cell_12_68 (.BL(BL68),.BLN(BLN68),.WL(WL12));
sram_cell_6t_5 inst_cell_12_69 (.BL(BL69),.BLN(BLN69),.WL(WL12));
sram_cell_6t_5 inst_cell_12_70 (.BL(BL70),.BLN(BLN70),.WL(WL12));
sram_cell_6t_5 inst_cell_12_71 (.BL(BL71),.BLN(BLN71),.WL(WL12));
sram_cell_6t_5 inst_cell_12_72 (.BL(BL72),.BLN(BLN72),.WL(WL12));
sram_cell_6t_5 inst_cell_12_73 (.BL(BL73),.BLN(BLN73),.WL(WL12));
sram_cell_6t_5 inst_cell_12_74 (.BL(BL74),.BLN(BLN74),.WL(WL12));
sram_cell_6t_5 inst_cell_12_75 (.BL(BL75),.BLN(BLN75),.WL(WL12));
sram_cell_6t_5 inst_cell_12_76 (.BL(BL76),.BLN(BLN76),.WL(WL12));
sram_cell_6t_5 inst_cell_12_77 (.BL(BL77),.BLN(BLN77),.WL(WL12));
sram_cell_6t_5 inst_cell_12_78 (.BL(BL78),.BLN(BLN78),.WL(WL12));
sram_cell_6t_5 inst_cell_12_79 (.BL(BL79),.BLN(BLN79),.WL(WL12));
sram_cell_6t_5 inst_cell_12_80 (.BL(BL80),.BLN(BLN80),.WL(WL12));
sram_cell_6t_5 inst_cell_12_81 (.BL(BL81),.BLN(BLN81),.WL(WL12));
sram_cell_6t_5 inst_cell_12_82 (.BL(BL82),.BLN(BLN82),.WL(WL12));
sram_cell_6t_5 inst_cell_12_83 (.BL(BL83),.BLN(BLN83),.WL(WL12));
sram_cell_6t_5 inst_cell_12_84 (.BL(BL84),.BLN(BLN84),.WL(WL12));
sram_cell_6t_5 inst_cell_12_85 (.BL(BL85),.BLN(BLN85),.WL(WL12));
sram_cell_6t_5 inst_cell_12_86 (.BL(BL86),.BLN(BLN86),.WL(WL12));
sram_cell_6t_5 inst_cell_12_87 (.BL(BL87),.BLN(BLN87),.WL(WL12));
sram_cell_6t_5 inst_cell_12_88 (.BL(BL88),.BLN(BLN88),.WL(WL12));
sram_cell_6t_5 inst_cell_12_89 (.BL(BL89),.BLN(BLN89),.WL(WL12));
sram_cell_6t_5 inst_cell_12_90 (.BL(BL90),.BLN(BLN90),.WL(WL12));
sram_cell_6t_5 inst_cell_12_91 (.BL(BL91),.BLN(BLN91),.WL(WL12));
sram_cell_6t_5 inst_cell_12_92 (.BL(BL92),.BLN(BLN92),.WL(WL12));
sram_cell_6t_5 inst_cell_12_93 (.BL(BL93),.BLN(BLN93),.WL(WL12));
sram_cell_6t_5 inst_cell_12_94 (.BL(BL94),.BLN(BLN94),.WL(WL12));
sram_cell_6t_5 inst_cell_12_95 (.BL(BL95),.BLN(BLN95),.WL(WL12));
sram_cell_6t_5 inst_cell_12_96 (.BL(BL96),.BLN(BLN96),.WL(WL12));
sram_cell_6t_5 inst_cell_12_97 (.BL(BL97),.BLN(BLN97),.WL(WL12));
sram_cell_6t_5 inst_cell_12_98 (.BL(BL98),.BLN(BLN98),.WL(WL12));
sram_cell_6t_5 inst_cell_12_99 (.BL(BL99),.BLN(BLN99),.WL(WL12));
sram_cell_6t_5 inst_cell_12_100 (.BL(BL100),.BLN(BLN100),.WL(WL12));
sram_cell_6t_5 inst_cell_12_101 (.BL(BL101),.BLN(BLN101),.WL(WL12));
sram_cell_6t_5 inst_cell_12_102 (.BL(BL102),.BLN(BLN102),.WL(WL12));
sram_cell_6t_5 inst_cell_12_103 (.BL(BL103),.BLN(BLN103),.WL(WL12));
sram_cell_6t_5 inst_cell_12_104 (.BL(BL104),.BLN(BLN104),.WL(WL12));
sram_cell_6t_5 inst_cell_12_105 (.BL(BL105),.BLN(BLN105),.WL(WL12));
sram_cell_6t_5 inst_cell_12_106 (.BL(BL106),.BLN(BLN106),.WL(WL12));
sram_cell_6t_5 inst_cell_12_107 (.BL(BL107),.BLN(BLN107),.WL(WL12));
sram_cell_6t_5 inst_cell_12_108 (.BL(BL108),.BLN(BLN108),.WL(WL12));
sram_cell_6t_5 inst_cell_12_109 (.BL(BL109),.BLN(BLN109),.WL(WL12));
sram_cell_6t_5 inst_cell_12_110 (.BL(BL110),.BLN(BLN110),.WL(WL12));
sram_cell_6t_5 inst_cell_12_111 (.BL(BL111),.BLN(BLN111),.WL(WL12));
sram_cell_6t_5 inst_cell_12_112 (.BL(BL112),.BLN(BLN112),.WL(WL12));
sram_cell_6t_5 inst_cell_12_113 (.BL(BL113),.BLN(BLN113),.WL(WL12));
sram_cell_6t_5 inst_cell_12_114 (.BL(BL114),.BLN(BLN114),.WL(WL12));
sram_cell_6t_5 inst_cell_12_115 (.BL(BL115),.BLN(BLN115),.WL(WL12));
sram_cell_6t_5 inst_cell_12_116 (.BL(BL116),.BLN(BLN116),.WL(WL12));
sram_cell_6t_5 inst_cell_12_117 (.BL(BL117),.BLN(BLN117),.WL(WL12));
sram_cell_6t_5 inst_cell_12_118 (.BL(BL118),.BLN(BLN118),.WL(WL12));
sram_cell_6t_5 inst_cell_12_119 (.BL(BL119),.BLN(BLN119),.WL(WL12));
sram_cell_6t_5 inst_cell_12_120 (.BL(BL120),.BLN(BLN120),.WL(WL12));
sram_cell_6t_5 inst_cell_12_121 (.BL(BL121),.BLN(BLN121),.WL(WL12));
sram_cell_6t_5 inst_cell_12_122 (.BL(BL122),.BLN(BLN122),.WL(WL12));
sram_cell_6t_5 inst_cell_12_123 (.BL(BL123),.BLN(BLN123),.WL(WL12));
sram_cell_6t_5 inst_cell_12_124 (.BL(BL124),.BLN(BLN124),.WL(WL12));
sram_cell_6t_5 inst_cell_12_125 (.BL(BL125),.BLN(BLN125),.WL(WL12));
sram_cell_6t_5 inst_cell_12_126 (.BL(BL126),.BLN(BLN126),.WL(WL12));
sram_cell_6t_5 inst_cell_12_127 (.BL(BL127),.BLN(BLN127),.WL(WL12));
sram_cell_6t_5 inst_cell_13_0 (.BL(BL0),.BLN(BLN0),.WL(WL13));
sram_cell_6t_5 inst_cell_13_1 (.BL(BL1),.BLN(BLN1),.WL(WL13));
sram_cell_6t_5 inst_cell_13_2 (.BL(BL2),.BLN(BLN2),.WL(WL13));
sram_cell_6t_5 inst_cell_13_3 (.BL(BL3),.BLN(BLN3),.WL(WL13));
sram_cell_6t_5 inst_cell_13_4 (.BL(BL4),.BLN(BLN4),.WL(WL13));
sram_cell_6t_5 inst_cell_13_5 (.BL(BL5),.BLN(BLN5),.WL(WL13));
sram_cell_6t_5 inst_cell_13_6 (.BL(BL6),.BLN(BLN6),.WL(WL13));
sram_cell_6t_5 inst_cell_13_7 (.BL(BL7),.BLN(BLN7),.WL(WL13));
sram_cell_6t_5 inst_cell_13_8 (.BL(BL8),.BLN(BLN8),.WL(WL13));
sram_cell_6t_5 inst_cell_13_9 (.BL(BL9),.BLN(BLN9),.WL(WL13));
sram_cell_6t_5 inst_cell_13_10 (.BL(BL10),.BLN(BLN10),.WL(WL13));
sram_cell_6t_5 inst_cell_13_11 (.BL(BL11),.BLN(BLN11),.WL(WL13));
sram_cell_6t_5 inst_cell_13_12 (.BL(BL12),.BLN(BLN12),.WL(WL13));
sram_cell_6t_5 inst_cell_13_13 (.BL(BL13),.BLN(BLN13),.WL(WL13));
sram_cell_6t_5 inst_cell_13_14 (.BL(BL14),.BLN(BLN14),.WL(WL13));
sram_cell_6t_5 inst_cell_13_15 (.BL(BL15),.BLN(BLN15),.WL(WL13));
sram_cell_6t_5 inst_cell_13_16 (.BL(BL16),.BLN(BLN16),.WL(WL13));
sram_cell_6t_5 inst_cell_13_17 (.BL(BL17),.BLN(BLN17),.WL(WL13));
sram_cell_6t_5 inst_cell_13_18 (.BL(BL18),.BLN(BLN18),.WL(WL13));
sram_cell_6t_5 inst_cell_13_19 (.BL(BL19),.BLN(BLN19),.WL(WL13));
sram_cell_6t_5 inst_cell_13_20 (.BL(BL20),.BLN(BLN20),.WL(WL13));
sram_cell_6t_5 inst_cell_13_21 (.BL(BL21),.BLN(BLN21),.WL(WL13));
sram_cell_6t_5 inst_cell_13_22 (.BL(BL22),.BLN(BLN22),.WL(WL13));
sram_cell_6t_5 inst_cell_13_23 (.BL(BL23),.BLN(BLN23),.WL(WL13));
sram_cell_6t_5 inst_cell_13_24 (.BL(BL24),.BLN(BLN24),.WL(WL13));
sram_cell_6t_5 inst_cell_13_25 (.BL(BL25),.BLN(BLN25),.WL(WL13));
sram_cell_6t_5 inst_cell_13_26 (.BL(BL26),.BLN(BLN26),.WL(WL13));
sram_cell_6t_5 inst_cell_13_27 (.BL(BL27),.BLN(BLN27),.WL(WL13));
sram_cell_6t_5 inst_cell_13_28 (.BL(BL28),.BLN(BLN28),.WL(WL13));
sram_cell_6t_5 inst_cell_13_29 (.BL(BL29),.BLN(BLN29),.WL(WL13));
sram_cell_6t_5 inst_cell_13_30 (.BL(BL30),.BLN(BLN30),.WL(WL13));
sram_cell_6t_5 inst_cell_13_31 (.BL(BL31),.BLN(BLN31),.WL(WL13));
sram_cell_6t_5 inst_cell_13_32 (.BL(BL32),.BLN(BLN32),.WL(WL13));
sram_cell_6t_5 inst_cell_13_33 (.BL(BL33),.BLN(BLN33),.WL(WL13));
sram_cell_6t_5 inst_cell_13_34 (.BL(BL34),.BLN(BLN34),.WL(WL13));
sram_cell_6t_5 inst_cell_13_35 (.BL(BL35),.BLN(BLN35),.WL(WL13));
sram_cell_6t_5 inst_cell_13_36 (.BL(BL36),.BLN(BLN36),.WL(WL13));
sram_cell_6t_5 inst_cell_13_37 (.BL(BL37),.BLN(BLN37),.WL(WL13));
sram_cell_6t_5 inst_cell_13_38 (.BL(BL38),.BLN(BLN38),.WL(WL13));
sram_cell_6t_5 inst_cell_13_39 (.BL(BL39),.BLN(BLN39),.WL(WL13));
sram_cell_6t_5 inst_cell_13_40 (.BL(BL40),.BLN(BLN40),.WL(WL13));
sram_cell_6t_5 inst_cell_13_41 (.BL(BL41),.BLN(BLN41),.WL(WL13));
sram_cell_6t_5 inst_cell_13_42 (.BL(BL42),.BLN(BLN42),.WL(WL13));
sram_cell_6t_5 inst_cell_13_43 (.BL(BL43),.BLN(BLN43),.WL(WL13));
sram_cell_6t_5 inst_cell_13_44 (.BL(BL44),.BLN(BLN44),.WL(WL13));
sram_cell_6t_5 inst_cell_13_45 (.BL(BL45),.BLN(BLN45),.WL(WL13));
sram_cell_6t_5 inst_cell_13_46 (.BL(BL46),.BLN(BLN46),.WL(WL13));
sram_cell_6t_5 inst_cell_13_47 (.BL(BL47),.BLN(BLN47),.WL(WL13));
sram_cell_6t_5 inst_cell_13_48 (.BL(BL48),.BLN(BLN48),.WL(WL13));
sram_cell_6t_5 inst_cell_13_49 (.BL(BL49),.BLN(BLN49),.WL(WL13));
sram_cell_6t_5 inst_cell_13_50 (.BL(BL50),.BLN(BLN50),.WL(WL13));
sram_cell_6t_5 inst_cell_13_51 (.BL(BL51),.BLN(BLN51),.WL(WL13));
sram_cell_6t_5 inst_cell_13_52 (.BL(BL52),.BLN(BLN52),.WL(WL13));
sram_cell_6t_5 inst_cell_13_53 (.BL(BL53),.BLN(BLN53),.WL(WL13));
sram_cell_6t_5 inst_cell_13_54 (.BL(BL54),.BLN(BLN54),.WL(WL13));
sram_cell_6t_5 inst_cell_13_55 (.BL(BL55),.BLN(BLN55),.WL(WL13));
sram_cell_6t_5 inst_cell_13_56 (.BL(BL56),.BLN(BLN56),.WL(WL13));
sram_cell_6t_5 inst_cell_13_57 (.BL(BL57),.BLN(BLN57),.WL(WL13));
sram_cell_6t_5 inst_cell_13_58 (.BL(BL58),.BLN(BLN58),.WL(WL13));
sram_cell_6t_5 inst_cell_13_59 (.BL(BL59),.BLN(BLN59),.WL(WL13));
sram_cell_6t_5 inst_cell_13_60 (.BL(BL60),.BLN(BLN60),.WL(WL13));
sram_cell_6t_5 inst_cell_13_61 (.BL(BL61),.BLN(BLN61),.WL(WL13));
sram_cell_6t_5 inst_cell_13_62 (.BL(BL62),.BLN(BLN62),.WL(WL13));
sram_cell_6t_5 inst_cell_13_63 (.BL(BL63),.BLN(BLN63),.WL(WL13));
sram_cell_6t_5 inst_cell_13_64 (.BL(BL64),.BLN(BLN64),.WL(WL13));
sram_cell_6t_5 inst_cell_13_65 (.BL(BL65),.BLN(BLN65),.WL(WL13));
sram_cell_6t_5 inst_cell_13_66 (.BL(BL66),.BLN(BLN66),.WL(WL13));
sram_cell_6t_5 inst_cell_13_67 (.BL(BL67),.BLN(BLN67),.WL(WL13));
sram_cell_6t_5 inst_cell_13_68 (.BL(BL68),.BLN(BLN68),.WL(WL13));
sram_cell_6t_5 inst_cell_13_69 (.BL(BL69),.BLN(BLN69),.WL(WL13));
sram_cell_6t_5 inst_cell_13_70 (.BL(BL70),.BLN(BLN70),.WL(WL13));
sram_cell_6t_5 inst_cell_13_71 (.BL(BL71),.BLN(BLN71),.WL(WL13));
sram_cell_6t_5 inst_cell_13_72 (.BL(BL72),.BLN(BLN72),.WL(WL13));
sram_cell_6t_5 inst_cell_13_73 (.BL(BL73),.BLN(BLN73),.WL(WL13));
sram_cell_6t_5 inst_cell_13_74 (.BL(BL74),.BLN(BLN74),.WL(WL13));
sram_cell_6t_5 inst_cell_13_75 (.BL(BL75),.BLN(BLN75),.WL(WL13));
sram_cell_6t_5 inst_cell_13_76 (.BL(BL76),.BLN(BLN76),.WL(WL13));
sram_cell_6t_5 inst_cell_13_77 (.BL(BL77),.BLN(BLN77),.WL(WL13));
sram_cell_6t_5 inst_cell_13_78 (.BL(BL78),.BLN(BLN78),.WL(WL13));
sram_cell_6t_5 inst_cell_13_79 (.BL(BL79),.BLN(BLN79),.WL(WL13));
sram_cell_6t_5 inst_cell_13_80 (.BL(BL80),.BLN(BLN80),.WL(WL13));
sram_cell_6t_5 inst_cell_13_81 (.BL(BL81),.BLN(BLN81),.WL(WL13));
sram_cell_6t_5 inst_cell_13_82 (.BL(BL82),.BLN(BLN82),.WL(WL13));
sram_cell_6t_5 inst_cell_13_83 (.BL(BL83),.BLN(BLN83),.WL(WL13));
sram_cell_6t_5 inst_cell_13_84 (.BL(BL84),.BLN(BLN84),.WL(WL13));
sram_cell_6t_5 inst_cell_13_85 (.BL(BL85),.BLN(BLN85),.WL(WL13));
sram_cell_6t_5 inst_cell_13_86 (.BL(BL86),.BLN(BLN86),.WL(WL13));
sram_cell_6t_5 inst_cell_13_87 (.BL(BL87),.BLN(BLN87),.WL(WL13));
sram_cell_6t_5 inst_cell_13_88 (.BL(BL88),.BLN(BLN88),.WL(WL13));
sram_cell_6t_5 inst_cell_13_89 (.BL(BL89),.BLN(BLN89),.WL(WL13));
sram_cell_6t_5 inst_cell_13_90 (.BL(BL90),.BLN(BLN90),.WL(WL13));
sram_cell_6t_5 inst_cell_13_91 (.BL(BL91),.BLN(BLN91),.WL(WL13));
sram_cell_6t_5 inst_cell_13_92 (.BL(BL92),.BLN(BLN92),.WL(WL13));
sram_cell_6t_5 inst_cell_13_93 (.BL(BL93),.BLN(BLN93),.WL(WL13));
sram_cell_6t_5 inst_cell_13_94 (.BL(BL94),.BLN(BLN94),.WL(WL13));
sram_cell_6t_5 inst_cell_13_95 (.BL(BL95),.BLN(BLN95),.WL(WL13));
sram_cell_6t_5 inst_cell_13_96 (.BL(BL96),.BLN(BLN96),.WL(WL13));
sram_cell_6t_5 inst_cell_13_97 (.BL(BL97),.BLN(BLN97),.WL(WL13));
sram_cell_6t_5 inst_cell_13_98 (.BL(BL98),.BLN(BLN98),.WL(WL13));
sram_cell_6t_5 inst_cell_13_99 (.BL(BL99),.BLN(BLN99),.WL(WL13));
sram_cell_6t_5 inst_cell_13_100 (.BL(BL100),.BLN(BLN100),.WL(WL13));
sram_cell_6t_5 inst_cell_13_101 (.BL(BL101),.BLN(BLN101),.WL(WL13));
sram_cell_6t_5 inst_cell_13_102 (.BL(BL102),.BLN(BLN102),.WL(WL13));
sram_cell_6t_5 inst_cell_13_103 (.BL(BL103),.BLN(BLN103),.WL(WL13));
sram_cell_6t_5 inst_cell_13_104 (.BL(BL104),.BLN(BLN104),.WL(WL13));
sram_cell_6t_5 inst_cell_13_105 (.BL(BL105),.BLN(BLN105),.WL(WL13));
sram_cell_6t_5 inst_cell_13_106 (.BL(BL106),.BLN(BLN106),.WL(WL13));
sram_cell_6t_5 inst_cell_13_107 (.BL(BL107),.BLN(BLN107),.WL(WL13));
sram_cell_6t_5 inst_cell_13_108 (.BL(BL108),.BLN(BLN108),.WL(WL13));
sram_cell_6t_5 inst_cell_13_109 (.BL(BL109),.BLN(BLN109),.WL(WL13));
sram_cell_6t_5 inst_cell_13_110 (.BL(BL110),.BLN(BLN110),.WL(WL13));
sram_cell_6t_5 inst_cell_13_111 (.BL(BL111),.BLN(BLN111),.WL(WL13));
sram_cell_6t_5 inst_cell_13_112 (.BL(BL112),.BLN(BLN112),.WL(WL13));
sram_cell_6t_5 inst_cell_13_113 (.BL(BL113),.BLN(BLN113),.WL(WL13));
sram_cell_6t_5 inst_cell_13_114 (.BL(BL114),.BLN(BLN114),.WL(WL13));
sram_cell_6t_5 inst_cell_13_115 (.BL(BL115),.BLN(BLN115),.WL(WL13));
sram_cell_6t_5 inst_cell_13_116 (.BL(BL116),.BLN(BLN116),.WL(WL13));
sram_cell_6t_5 inst_cell_13_117 (.BL(BL117),.BLN(BLN117),.WL(WL13));
sram_cell_6t_5 inst_cell_13_118 (.BL(BL118),.BLN(BLN118),.WL(WL13));
sram_cell_6t_5 inst_cell_13_119 (.BL(BL119),.BLN(BLN119),.WL(WL13));
sram_cell_6t_5 inst_cell_13_120 (.BL(BL120),.BLN(BLN120),.WL(WL13));
sram_cell_6t_5 inst_cell_13_121 (.BL(BL121),.BLN(BLN121),.WL(WL13));
sram_cell_6t_5 inst_cell_13_122 (.BL(BL122),.BLN(BLN122),.WL(WL13));
sram_cell_6t_5 inst_cell_13_123 (.BL(BL123),.BLN(BLN123),.WL(WL13));
sram_cell_6t_5 inst_cell_13_124 (.BL(BL124),.BLN(BLN124),.WL(WL13));
sram_cell_6t_5 inst_cell_13_125 (.BL(BL125),.BLN(BLN125),.WL(WL13));
sram_cell_6t_5 inst_cell_13_126 (.BL(BL126),.BLN(BLN126),.WL(WL13));
sram_cell_6t_5 inst_cell_13_127 (.BL(BL127),.BLN(BLN127),.WL(WL13));
sram_cell_6t_5 inst_cell_14_0 (.BL(BL0),.BLN(BLN0),.WL(WL14));
sram_cell_6t_5 inst_cell_14_1 (.BL(BL1),.BLN(BLN1),.WL(WL14));
sram_cell_6t_5 inst_cell_14_2 (.BL(BL2),.BLN(BLN2),.WL(WL14));
sram_cell_6t_5 inst_cell_14_3 (.BL(BL3),.BLN(BLN3),.WL(WL14));
sram_cell_6t_5 inst_cell_14_4 (.BL(BL4),.BLN(BLN4),.WL(WL14));
sram_cell_6t_5 inst_cell_14_5 (.BL(BL5),.BLN(BLN5),.WL(WL14));
sram_cell_6t_5 inst_cell_14_6 (.BL(BL6),.BLN(BLN6),.WL(WL14));
sram_cell_6t_5 inst_cell_14_7 (.BL(BL7),.BLN(BLN7),.WL(WL14));
sram_cell_6t_5 inst_cell_14_8 (.BL(BL8),.BLN(BLN8),.WL(WL14));
sram_cell_6t_5 inst_cell_14_9 (.BL(BL9),.BLN(BLN9),.WL(WL14));
sram_cell_6t_5 inst_cell_14_10 (.BL(BL10),.BLN(BLN10),.WL(WL14));
sram_cell_6t_5 inst_cell_14_11 (.BL(BL11),.BLN(BLN11),.WL(WL14));
sram_cell_6t_5 inst_cell_14_12 (.BL(BL12),.BLN(BLN12),.WL(WL14));
sram_cell_6t_5 inst_cell_14_13 (.BL(BL13),.BLN(BLN13),.WL(WL14));
sram_cell_6t_5 inst_cell_14_14 (.BL(BL14),.BLN(BLN14),.WL(WL14));
sram_cell_6t_5 inst_cell_14_15 (.BL(BL15),.BLN(BLN15),.WL(WL14));
sram_cell_6t_5 inst_cell_14_16 (.BL(BL16),.BLN(BLN16),.WL(WL14));
sram_cell_6t_5 inst_cell_14_17 (.BL(BL17),.BLN(BLN17),.WL(WL14));
sram_cell_6t_5 inst_cell_14_18 (.BL(BL18),.BLN(BLN18),.WL(WL14));
sram_cell_6t_5 inst_cell_14_19 (.BL(BL19),.BLN(BLN19),.WL(WL14));
sram_cell_6t_5 inst_cell_14_20 (.BL(BL20),.BLN(BLN20),.WL(WL14));
sram_cell_6t_5 inst_cell_14_21 (.BL(BL21),.BLN(BLN21),.WL(WL14));
sram_cell_6t_5 inst_cell_14_22 (.BL(BL22),.BLN(BLN22),.WL(WL14));
sram_cell_6t_5 inst_cell_14_23 (.BL(BL23),.BLN(BLN23),.WL(WL14));
sram_cell_6t_5 inst_cell_14_24 (.BL(BL24),.BLN(BLN24),.WL(WL14));
sram_cell_6t_5 inst_cell_14_25 (.BL(BL25),.BLN(BLN25),.WL(WL14));
sram_cell_6t_5 inst_cell_14_26 (.BL(BL26),.BLN(BLN26),.WL(WL14));
sram_cell_6t_5 inst_cell_14_27 (.BL(BL27),.BLN(BLN27),.WL(WL14));
sram_cell_6t_5 inst_cell_14_28 (.BL(BL28),.BLN(BLN28),.WL(WL14));
sram_cell_6t_5 inst_cell_14_29 (.BL(BL29),.BLN(BLN29),.WL(WL14));
sram_cell_6t_5 inst_cell_14_30 (.BL(BL30),.BLN(BLN30),.WL(WL14));
sram_cell_6t_5 inst_cell_14_31 (.BL(BL31),.BLN(BLN31),.WL(WL14));
sram_cell_6t_5 inst_cell_14_32 (.BL(BL32),.BLN(BLN32),.WL(WL14));
sram_cell_6t_5 inst_cell_14_33 (.BL(BL33),.BLN(BLN33),.WL(WL14));
sram_cell_6t_5 inst_cell_14_34 (.BL(BL34),.BLN(BLN34),.WL(WL14));
sram_cell_6t_5 inst_cell_14_35 (.BL(BL35),.BLN(BLN35),.WL(WL14));
sram_cell_6t_5 inst_cell_14_36 (.BL(BL36),.BLN(BLN36),.WL(WL14));
sram_cell_6t_5 inst_cell_14_37 (.BL(BL37),.BLN(BLN37),.WL(WL14));
sram_cell_6t_5 inst_cell_14_38 (.BL(BL38),.BLN(BLN38),.WL(WL14));
sram_cell_6t_5 inst_cell_14_39 (.BL(BL39),.BLN(BLN39),.WL(WL14));
sram_cell_6t_5 inst_cell_14_40 (.BL(BL40),.BLN(BLN40),.WL(WL14));
sram_cell_6t_5 inst_cell_14_41 (.BL(BL41),.BLN(BLN41),.WL(WL14));
sram_cell_6t_5 inst_cell_14_42 (.BL(BL42),.BLN(BLN42),.WL(WL14));
sram_cell_6t_5 inst_cell_14_43 (.BL(BL43),.BLN(BLN43),.WL(WL14));
sram_cell_6t_5 inst_cell_14_44 (.BL(BL44),.BLN(BLN44),.WL(WL14));
sram_cell_6t_5 inst_cell_14_45 (.BL(BL45),.BLN(BLN45),.WL(WL14));
sram_cell_6t_5 inst_cell_14_46 (.BL(BL46),.BLN(BLN46),.WL(WL14));
sram_cell_6t_5 inst_cell_14_47 (.BL(BL47),.BLN(BLN47),.WL(WL14));
sram_cell_6t_5 inst_cell_14_48 (.BL(BL48),.BLN(BLN48),.WL(WL14));
sram_cell_6t_5 inst_cell_14_49 (.BL(BL49),.BLN(BLN49),.WL(WL14));
sram_cell_6t_5 inst_cell_14_50 (.BL(BL50),.BLN(BLN50),.WL(WL14));
sram_cell_6t_5 inst_cell_14_51 (.BL(BL51),.BLN(BLN51),.WL(WL14));
sram_cell_6t_5 inst_cell_14_52 (.BL(BL52),.BLN(BLN52),.WL(WL14));
sram_cell_6t_5 inst_cell_14_53 (.BL(BL53),.BLN(BLN53),.WL(WL14));
sram_cell_6t_5 inst_cell_14_54 (.BL(BL54),.BLN(BLN54),.WL(WL14));
sram_cell_6t_5 inst_cell_14_55 (.BL(BL55),.BLN(BLN55),.WL(WL14));
sram_cell_6t_5 inst_cell_14_56 (.BL(BL56),.BLN(BLN56),.WL(WL14));
sram_cell_6t_5 inst_cell_14_57 (.BL(BL57),.BLN(BLN57),.WL(WL14));
sram_cell_6t_5 inst_cell_14_58 (.BL(BL58),.BLN(BLN58),.WL(WL14));
sram_cell_6t_5 inst_cell_14_59 (.BL(BL59),.BLN(BLN59),.WL(WL14));
sram_cell_6t_5 inst_cell_14_60 (.BL(BL60),.BLN(BLN60),.WL(WL14));
sram_cell_6t_5 inst_cell_14_61 (.BL(BL61),.BLN(BLN61),.WL(WL14));
sram_cell_6t_5 inst_cell_14_62 (.BL(BL62),.BLN(BLN62),.WL(WL14));
sram_cell_6t_5 inst_cell_14_63 (.BL(BL63),.BLN(BLN63),.WL(WL14));
sram_cell_6t_5 inst_cell_14_64 (.BL(BL64),.BLN(BLN64),.WL(WL14));
sram_cell_6t_5 inst_cell_14_65 (.BL(BL65),.BLN(BLN65),.WL(WL14));
sram_cell_6t_5 inst_cell_14_66 (.BL(BL66),.BLN(BLN66),.WL(WL14));
sram_cell_6t_5 inst_cell_14_67 (.BL(BL67),.BLN(BLN67),.WL(WL14));
sram_cell_6t_5 inst_cell_14_68 (.BL(BL68),.BLN(BLN68),.WL(WL14));
sram_cell_6t_5 inst_cell_14_69 (.BL(BL69),.BLN(BLN69),.WL(WL14));
sram_cell_6t_5 inst_cell_14_70 (.BL(BL70),.BLN(BLN70),.WL(WL14));
sram_cell_6t_5 inst_cell_14_71 (.BL(BL71),.BLN(BLN71),.WL(WL14));
sram_cell_6t_5 inst_cell_14_72 (.BL(BL72),.BLN(BLN72),.WL(WL14));
sram_cell_6t_5 inst_cell_14_73 (.BL(BL73),.BLN(BLN73),.WL(WL14));
sram_cell_6t_5 inst_cell_14_74 (.BL(BL74),.BLN(BLN74),.WL(WL14));
sram_cell_6t_5 inst_cell_14_75 (.BL(BL75),.BLN(BLN75),.WL(WL14));
sram_cell_6t_5 inst_cell_14_76 (.BL(BL76),.BLN(BLN76),.WL(WL14));
sram_cell_6t_5 inst_cell_14_77 (.BL(BL77),.BLN(BLN77),.WL(WL14));
sram_cell_6t_5 inst_cell_14_78 (.BL(BL78),.BLN(BLN78),.WL(WL14));
sram_cell_6t_5 inst_cell_14_79 (.BL(BL79),.BLN(BLN79),.WL(WL14));
sram_cell_6t_5 inst_cell_14_80 (.BL(BL80),.BLN(BLN80),.WL(WL14));
sram_cell_6t_5 inst_cell_14_81 (.BL(BL81),.BLN(BLN81),.WL(WL14));
sram_cell_6t_5 inst_cell_14_82 (.BL(BL82),.BLN(BLN82),.WL(WL14));
sram_cell_6t_5 inst_cell_14_83 (.BL(BL83),.BLN(BLN83),.WL(WL14));
sram_cell_6t_5 inst_cell_14_84 (.BL(BL84),.BLN(BLN84),.WL(WL14));
sram_cell_6t_5 inst_cell_14_85 (.BL(BL85),.BLN(BLN85),.WL(WL14));
sram_cell_6t_5 inst_cell_14_86 (.BL(BL86),.BLN(BLN86),.WL(WL14));
sram_cell_6t_5 inst_cell_14_87 (.BL(BL87),.BLN(BLN87),.WL(WL14));
sram_cell_6t_5 inst_cell_14_88 (.BL(BL88),.BLN(BLN88),.WL(WL14));
sram_cell_6t_5 inst_cell_14_89 (.BL(BL89),.BLN(BLN89),.WL(WL14));
sram_cell_6t_5 inst_cell_14_90 (.BL(BL90),.BLN(BLN90),.WL(WL14));
sram_cell_6t_5 inst_cell_14_91 (.BL(BL91),.BLN(BLN91),.WL(WL14));
sram_cell_6t_5 inst_cell_14_92 (.BL(BL92),.BLN(BLN92),.WL(WL14));
sram_cell_6t_5 inst_cell_14_93 (.BL(BL93),.BLN(BLN93),.WL(WL14));
sram_cell_6t_5 inst_cell_14_94 (.BL(BL94),.BLN(BLN94),.WL(WL14));
sram_cell_6t_5 inst_cell_14_95 (.BL(BL95),.BLN(BLN95),.WL(WL14));
sram_cell_6t_5 inst_cell_14_96 (.BL(BL96),.BLN(BLN96),.WL(WL14));
sram_cell_6t_5 inst_cell_14_97 (.BL(BL97),.BLN(BLN97),.WL(WL14));
sram_cell_6t_5 inst_cell_14_98 (.BL(BL98),.BLN(BLN98),.WL(WL14));
sram_cell_6t_5 inst_cell_14_99 (.BL(BL99),.BLN(BLN99),.WL(WL14));
sram_cell_6t_5 inst_cell_14_100 (.BL(BL100),.BLN(BLN100),.WL(WL14));
sram_cell_6t_5 inst_cell_14_101 (.BL(BL101),.BLN(BLN101),.WL(WL14));
sram_cell_6t_5 inst_cell_14_102 (.BL(BL102),.BLN(BLN102),.WL(WL14));
sram_cell_6t_5 inst_cell_14_103 (.BL(BL103),.BLN(BLN103),.WL(WL14));
sram_cell_6t_5 inst_cell_14_104 (.BL(BL104),.BLN(BLN104),.WL(WL14));
sram_cell_6t_5 inst_cell_14_105 (.BL(BL105),.BLN(BLN105),.WL(WL14));
sram_cell_6t_5 inst_cell_14_106 (.BL(BL106),.BLN(BLN106),.WL(WL14));
sram_cell_6t_5 inst_cell_14_107 (.BL(BL107),.BLN(BLN107),.WL(WL14));
sram_cell_6t_5 inst_cell_14_108 (.BL(BL108),.BLN(BLN108),.WL(WL14));
sram_cell_6t_5 inst_cell_14_109 (.BL(BL109),.BLN(BLN109),.WL(WL14));
sram_cell_6t_5 inst_cell_14_110 (.BL(BL110),.BLN(BLN110),.WL(WL14));
sram_cell_6t_5 inst_cell_14_111 (.BL(BL111),.BLN(BLN111),.WL(WL14));
sram_cell_6t_5 inst_cell_14_112 (.BL(BL112),.BLN(BLN112),.WL(WL14));
sram_cell_6t_5 inst_cell_14_113 (.BL(BL113),.BLN(BLN113),.WL(WL14));
sram_cell_6t_5 inst_cell_14_114 (.BL(BL114),.BLN(BLN114),.WL(WL14));
sram_cell_6t_5 inst_cell_14_115 (.BL(BL115),.BLN(BLN115),.WL(WL14));
sram_cell_6t_5 inst_cell_14_116 (.BL(BL116),.BLN(BLN116),.WL(WL14));
sram_cell_6t_5 inst_cell_14_117 (.BL(BL117),.BLN(BLN117),.WL(WL14));
sram_cell_6t_5 inst_cell_14_118 (.BL(BL118),.BLN(BLN118),.WL(WL14));
sram_cell_6t_5 inst_cell_14_119 (.BL(BL119),.BLN(BLN119),.WL(WL14));
sram_cell_6t_5 inst_cell_14_120 (.BL(BL120),.BLN(BLN120),.WL(WL14));
sram_cell_6t_5 inst_cell_14_121 (.BL(BL121),.BLN(BLN121),.WL(WL14));
sram_cell_6t_5 inst_cell_14_122 (.BL(BL122),.BLN(BLN122),.WL(WL14));
sram_cell_6t_5 inst_cell_14_123 (.BL(BL123),.BLN(BLN123),.WL(WL14));
sram_cell_6t_5 inst_cell_14_124 (.BL(BL124),.BLN(BLN124),.WL(WL14));
sram_cell_6t_5 inst_cell_14_125 (.BL(BL125),.BLN(BLN125),.WL(WL14));
sram_cell_6t_5 inst_cell_14_126 (.BL(BL126),.BLN(BLN126),.WL(WL14));
sram_cell_6t_5 inst_cell_14_127 (.BL(BL127),.BLN(BLN127),.WL(WL14));
sram_cell_6t_5 inst_cell_15_0 (.BL(BL0),.BLN(BLN0),.WL(WL15));
sram_cell_6t_5 inst_cell_15_1 (.BL(BL1),.BLN(BLN1),.WL(WL15));
sram_cell_6t_5 inst_cell_15_2 (.BL(BL2),.BLN(BLN2),.WL(WL15));
sram_cell_6t_5 inst_cell_15_3 (.BL(BL3),.BLN(BLN3),.WL(WL15));
sram_cell_6t_5 inst_cell_15_4 (.BL(BL4),.BLN(BLN4),.WL(WL15));
sram_cell_6t_5 inst_cell_15_5 (.BL(BL5),.BLN(BLN5),.WL(WL15));
sram_cell_6t_5 inst_cell_15_6 (.BL(BL6),.BLN(BLN6),.WL(WL15));
sram_cell_6t_5 inst_cell_15_7 (.BL(BL7),.BLN(BLN7),.WL(WL15));
sram_cell_6t_5 inst_cell_15_8 (.BL(BL8),.BLN(BLN8),.WL(WL15));
sram_cell_6t_5 inst_cell_15_9 (.BL(BL9),.BLN(BLN9),.WL(WL15));
sram_cell_6t_5 inst_cell_15_10 (.BL(BL10),.BLN(BLN10),.WL(WL15));
sram_cell_6t_5 inst_cell_15_11 (.BL(BL11),.BLN(BLN11),.WL(WL15));
sram_cell_6t_5 inst_cell_15_12 (.BL(BL12),.BLN(BLN12),.WL(WL15));
sram_cell_6t_5 inst_cell_15_13 (.BL(BL13),.BLN(BLN13),.WL(WL15));
sram_cell_6t_5 inst_cell_15_14 (.BL(BL14),.BLN(BLN14),.WL(WL15));
sram_cell_6t_5 inst_cell_15_15 (.BL(BL15),.BLN(BLN15),.WL(WL15));
sram_cell_6t_5 inst_cell_15_16 (.BL(BL16),.BLN(BLN16),.WL(WL15));
sram_cell_6t_5 inst_cell_15_17 (.BL(BL17),.BLN(BLN17),.WL(WL15));
sram_cell_6t_5 inst_cell_15_18 (.BL(BL18),.BLN(BLN18),.WL(WL15));
sram_cell_6t_5 inst_cell_15_19 (.BL(BL19),.BLN(BLN19),.WL(WL15));
sram_cell_6t_5 inst_cell_15_20 (.BL(BL20),.BLN(BLN20),.WL(WL15));
sram_cell_6t_5 inst_cell_15_21 (.BL(BL21),.BLN(BLN21),.WL(WL15));
sram_cell_6t_5 inst_cell_15_22 (.BL(BL22),.BLN(BLN22),.WL(WL15));
sram_cell_6t_5 inst_cell_15_23 (.BL(BL23),.BLN(BLN23),.WL(WL15));
sram_cell_6t_5 inst_cell_15_24 (.BL(BL24),.BLN(BLN24),.WL(WL15));
sram_cell_6t_5 inst_cell_15_25 (.BL(BL25),.BLN(BLN25),.WL(WL15));
sram_cell_6t_5 inst_cell_15_26 (.BL(BL26),.BLN(BLN26),.WL(WL15));
sram_cell_6t_5 inst_cell_15_27 (.BL(BL27),.BLN(BLN27),.WL(WL15));
sram_cell_6t_5 inst_cell_15_28 (.BL(BL28),.BLN(BLN28),.WL(WL15));
sram_cell_6t_5 inst_cell_15_29 (.BL(BL29),.BLN(BLN29),.WL(WL15));
sram_cell_6t_5 inst_cell_15_30 (.BL(BL30),.BLN(BLN30),.WL(WL15));
sram_cell_6t_5 inst_cell_15_31 (.BL(BL31),.BLN(BLN31),.WL(WL15));
sram_cell_6t_5 inst_cell_15_32 (.BL(BL32),.BLN(BLN32),.WL(WL15));
sram_cell_6t_5 inst_cell_15_33 (.BL(BL33),.BLN(BLN33),.WL(WL15));
sram_cell_6t_5 inst_cell_15_34 (.BL(BL34),.BLN(BLN34),.WL(WL15));
sram_cell_6t_5 inst_cell_15_35 (.BL(BL35),.BLN(BLN35),.WL(WL15));
sram_cell_6t_5 inst_cell_15_36 (.BL(BL36),.BLN(BLN36),.WL(WL15));
sram_cell_6t_5 inst_cell_15_37 (.BL(BL37),.BLN(BLN37),.WL(WL15));
sram_cell_6t_5 inst_cell_15_38 (.BL(BL38),.BLN(BLN38),.WL(WL15));
sram_cell_6t_5 inst_cell_15_39 (.BL(BL39),.BLN(BLN39),.WL(WL15));
sram_cell_6t_5 inst_cell_15_40 (.BL(BL40),.BLN(BLN40),.WL(WL15));
sram_cell_6t_5 inst_cell_15_41 (.BL(BL41),.BLN(BLN41),.WL(WL15));
sram_cell_6t_5 inst_cell_15_42 (.BL(BL42),.BLN(BLN42),.WL(WL15));
sram_cell_6t_5 inst_cell_15_43 (.BL(BL43),.BLN(BLN43),.WL(WL15));
sram_cell_6t_5 inst_cell_15_44 (.BL(BL44),.BLN(BLN44),.WL(WL15));
sram_cell_6t_5 inst_cell_15_45 (.BL(BL45),.BLN(BLN45),.WL(WL15));
sram_cell_6t_5 inst_cell_15_46 (.BL(BL46),.BLN(BLN46),.WL(WL15));
sram_cell_6t_5 inst_cell_15_47 (.BL(BL47),.BLN(BLN47),.WL(WL15));
sram_cell_6t_5 inst_cell_15_48 (.BL(BL48),.BLN(BLN48),.WL(WL15));
sram_cell_6t_5 inst_cell_15_49 (.BL(BL49),.BLN(BLN49),.WL(WL15));
sram_cell_6t_5 inst_cell_15_50 (.BL(BL50),.BLN(BLN50),.WL(WL15));
sram_cell_6t_5 inst_cell_15_51 (.BL(BL51),.BLN(BLN51),.WL(WL15));
sram_cell_6t_5 inst_cell_15_52 (.BL(BL52),.BLN(BLN52),.WL(WL15));
sram_cell_6t_5 inst_cell_15_53 (.BL(BL53),.BLN(BLN53),.WL(WL15));
sram_cell_6t_5 inst_cell_15_54 (.BL(BL54),.BLN(BLN54),.WL(WL15));
sram_cell_6t_5 inst_cell_15_55 (.BL(BL55),.BLN(BLN55),.WL(WL15));
sram_cell_6t_5 inst_cell_15_56 (.BL(BL56),.BLN(BLN56),.WL(WL15));
sram_cell_6t_5 inst_cell_15_57 (.BL(BL57),.BLN(BLN57),.WL(WL15));
sram_cell_6t_5 inst_cell_15_58 (.BL(BL58),.BLN(BLN58),.WL(WL15));
sram_cell_6t_5 inst_cell_15_59 (.BL(BL59),.BLN(BLN59),.WL(WL15));
sram_cell_6t_5 inst_cell_15_60 (.BL(BL60),.BLN(BLN60),.WL(WL15));
sram_cell_6t_5 inst_cell_15_61 (.BL(BL61),.BLN(BLN61),.WL(WL15));
sram_cell_6t_5 inst_cell_15_62 (.BL(BL62),.BLN(BLN62),.WL(WL15));
sram_cell_6t_5 inst_cell_15_63 (.BL(BL63),.BLN(BLN63),.WL(WL15));
sram_cell_6t_5 inst_cell_15_64 (.BL(BL64),.BLN(BLN64),.WL(WL15));
sram_cell_6t_5 inst_cell_15_65 (.BL(BL65),.BLN(BLN65),.WL(WL15));
sram_cell_6t_5 inst_cell_15_66 (.BL(BL66),.BLN(BLN66),.WL(WL15));
sram_cell_6t_5 inst_cell_15_67 (.BL(BL67),.BLN(BLN67),.WL(WL15));
sram_cell_6t_5 inst_cell_15_68 (.BL(BL68),.BLN(BLN68),.WL(WL15));
sram_cell_6t_5 inst_cell_15_69 (.BL(BL69),.BLN(BLN69),.WL(WL15));
sram_cell_6t_5 inst_cell_15_70 (.BL(BL70),.BLN(BLN70),.WL(WL15));
sram_cell_6t_5 inst_cell_15_71 (.BL(BL71),.BLN(BLN71),.WL(WL15));
sram_cell_6t_5 inst_cell_15_72 (.BL(BL72),.BLN(BLN72),.WL(WL15));
sram_cell_6t_5 inst_cell_15_73 (.BL(BL73),.BLN(BLN73),.WL(WL15));
sram_cell_6t_5 inst_cell_15_74 (.BL(BL74),.BLN(BLN74),.WL(WL15));
sram_cell_6t_5 inst_cell_15_75 (.BL(BL75),.BLN(BLN75),.WL(WL15));
sram_cell_6t_5 inst_cell_15_76 (.BL(BL76),.BLN(BLN76),.WL(WL15));
sram_cell_6t_5 inst_cell_15_77 (.BL(BL77),.BLN(BLN77),.WL(WL15));
sram_cell_6t_5 inst_cell_15_78 (.BL(BL78),.BLN(BLN78),.WL(WL15));
sram_cell_6t_5 inst_cell_15_79 (.BL(BL79),.BLN(BLN79),.WL(WL15));
sram_cell_6t_5 inst_cell_15_80 (.BL(BL80),.BLN(BLN80),.WL(WL15));
sram_cell_6t_5 inst_cell_15_81 (.BL(BL81),.BLN(BLN81),.WL(WL15));
sram_cell_6t_5 inst_cell_15_82 (.BL(BL82),.BLN(BLN82),.WL(WL15));
sram_cell_6t_5 inst_cell_15_83 (.BL(BL83),.BLN(BLN83),.WL(WL15));
sram_cell_6t_5 inst_cell_15_84 (.BL(BL84),.BLN(BLN84),.WL(WL15));
sram_cell_6t_5 inst_cell_15_85 (.BL(BL85),.BLN(BLN85),.WL(WL15));
sram_cell_6t_5 inst_cell_15_86 (.BL(BL86),.BLN(BLN86),.WL(WL15));
sram_cell_6t_5 inst_cell_15_87 (.BL(BL87),.BLN(BLN87),.WL(WL15));
sram_cell_6t_5 inst_cell_15_88 (.BL(BL88),.BLN(BLN88),.WL(WL15));
sram_cell_6t_5 inst_cell_15_89 (.BL(BL89),.BLN(BLN89),.WL(WL15));
sram_cell_6t_5 inst_cell_15_90 (.BL(BL90),.BLN(BLN90),.WL(WL15));
sram_cell_6t_5 inst_cell_15_91 (.BL(BL91),.BLN(BLN91),.WL(WL15));
sram_cell_6t_5 inst_cell_15_92 (.BL(BL92),.BLN(BLN92),.WL(WL15));
sram_cell_6t_5 inst_cell_15_93 (.BL(BL93),.BLN(BLN93),.WL(WL15));
sram_cell_6t_5 inst_cell_15_94 (.BL(BL94),.BLN(BLN94),.WL(WL15));
sram_cell_6t_5 inst_cell_15_95 (.BL(BL95),.BLN(BLN95),.WL(WL15));
sram_cell_6t_5 inst_cell_15_96 (.BL(BL96),.BLN(BLN96),.WL(WL15));
sram_cell_6t_5 inst_cell_15_97 (.BL(BL97),.BLN(BLN97),.WL(WL15));
sram_cell_6t_5 inst_cell_15_98 (.BL(BL98),.BLN(BLN98),.WL(WL15));
sram_cell_6t_5 inst_cell_15_99 (.BL(BL99),.BLN(BLN99),.WL(WL15));
sram_cell_6t_5 inst_cell_15_100 (.BL(BL100),.BLN(BLN100),.WL(WL15));
sram_cell_6t_5 inst_cell_15_101 (.BL(BL101),.BLN(BLN101),.WL(WL15));
sram_cell_6t_5 inst_cell_15_102 (.BL(BL102),.BLN(BLN102),.WL(WL15));
sram_cell_6t_5 inst_cell_15_103 (.BL(BL103),.BLN(BLN103),.WL(WL15));
sram_cell_6t_5 inst_cell_15_104 (.BL(BL104),.BLN(BLN104),.WL(WL15));
sram_cell_6t_5 inst_cell_15_105 (.BL(BL105),.BLN(BLN105),.WL(WL15));
sram_cell_6t_5 inst_cell_15_106 (.BL(BL106),.BLN(BLN106),.WL(WL15));
sram_cell_6t_5 inst_cell_15_107 (.BL(BL107),.BLN(BLN107),.WL(WL15));
sram_cell_6t_5 inst_cell_15_108 (.BL(BL108),.BLN(BLN108),.WL(WL15));
sram_cell_6t_5 inst_cell_15_109 (.BL(BL109),.BLN(BLN109),.WL(WL15));
sram_cell_6t_5 inst_cell_15_110 (.BL(BL110),.BLN(BLN110),.WL(WL15));
sram_cell_6t_5 inst_cell_15_111 (.BL(BL111),.BLN(BLN111),.WL(WL15));
sram_cell_6t_5 inst_cell_15_112 (.BL(BL112),.BLN(BLN112),.WL(WL15));
sram_cell_6t_5 inst_cell_15_113 (.BL(BL113),.BLN(BLN113),.WL(WL15));
sram_cell_6t_5 inst_cell_15_114 (.BL(BL114),.BLN(BLN114),.WL(WL15));
sram_cell_6t_5 inst_cell_15_115 (.BL(BL115),.BLN(BLN115),.WL(WL15));
sram_cell_6t_5 inst_cell_15_116 (.BL(BL116),.BLN(BLN116),.WL(WL15));
sram_cell_6t_5 inst_cell_15_117 (.BL(BL117),.BLN(BLN117),.WL(WL15));
sram_cell_6t_5 inst_cell_15_118 (.BL(BL118),.BLN(BLN118),.WL(WL15));
sram_cell_6t_5 inst_cell_15_119 (.BL(BL119),.BLN(BLN119),.WL(WL15));
sram_cell_6t_5 inst_cell_15_120 (.BL(BL120),.BLN(BLN120),.WL(WL15));
sram_cell_6t_5 inst_cell_15_121 (.BL(BL121),.BLN(BLN121),.WL(WL15));
sram_cell_6t_5 inst_cell_15_122 (.BL(BL122),.BLN(BLN122),.WL(WL15));
sram_cell_6t_5 inst_cell_15_123 (.BL(BL123),.BLN(BLN123),.WL(WL15));
sram_cell_6t_5 inst_cell_15_124 (.BL(BL124),.BLN(BLN124),.WL(WL15));
sram_cell_6t_5 inst_cell_15_125 (.BL(BL125),.BLN(BLN125),.WL(WL15));
sram_cell_6t_5 inst_cell_15_126 (.BL(BL126),.BLN(BLN126),.WL(WL15));
sram_cell_6t_5 inst_cell_15_127 (.BL(BL127),.BLN(BLN127),.WL(WL15));
sram_cell_6t_5 inst_cell_16_0 (.BL(BL0),.BLN(BLN0),.WL(WL16));
sram_cell_6t_5 inst_cell_16_1 (.BL(BL1),.BLN(BLN1),.WL(WL16));
sram_cell_6t_5 inst_cell_16_2 (.BL(BL2),.BLN(BLN2),.WL(WL16));
sram_cell_6t_5 inst_cell_16_3 (.BL(BL3),.BLN(BLN3),.WL(WL16));
sram_cell_6t_5 inst_cell_16_4 (.BL(BL4),.BLN(BLN4),.WL(WL16));
sram_cell_6t_5 inst_cell_16_5 (.BL(BL5),.BLN(BLN5),.WL(WL16));
sram_cell_6t_5 inst_cell_16_6 (.BL(BL6),.BLN(BLN6),.WL(WL16));
sram_cell_6t_5 inst_cell_16_7 (.BL(BL7),.BLN(BLN7),.WL(WL16));
sram_cell_6t_5 inst_cell_16_8 (.BL(BL8),.BLN(BLN8),.WL(WL16));
sram_cell_6t_5 inst_cell_16_9 (.BL(BL9),.BLN(BLN9),.WL(WL16));
sram_cell_6t_5 inst_cell_16_10 (.BL(BL10),.BLN(BLN10),.WL(WL16));
sram_cell_6t_5 inst_cell_16_11 (.BL(BL11),.BLN(BLN11),.WL(WL16));
sram_cell_6t_5 inst_cell_16_12 (.BL(BL12),.BLN(BLN12),.WL(WL16));
sram_cell_6t_5 inst_cell_16_13 (.BL(BL13),.BLN(BLN13),.WL(WL16));
sram_cell_6t_5 inst_cell_16_14 (.BL(BL14),.BLN(BLN14),.WL(WL16));
sram_cell_6t_5 inst_cell_16_15 (.BL(BL15),.BLN(BLN15),.WL(WL16));
sram_cell_6t_5 inst_cell_16_16 (.BL(BL16),.BLN(BLN16),.WL(WL16));
sram_cell_6t_5 inst_cell_16_17 (.BL(BL17),.BLN(BLN17),.WL(WL16));
sram_cell_6t_5 inst_cell_16_18 (.BL(BL18),.BLN(BLN18),.WL(WL16));
sram_cell_6t_5 inst_cell_16_19 (.BL(BL19),.BLN(BLN19),.WL(WL16));
sram_cell_6t_5 inst_cell_16_20 (.BL(BL20),.BLN(BLN20),.WL(WL16));
sram_cell_6t_5 inst_cell_16_21 (.BL(BL21),.BLN(BLN21),.WL(WL16));
sram_cell_6t_5 inst_cell_16_22 (.BL(BL22),.BLN(BLN22),.WL(WL16));
sram_cell_6t_5 inst_cell_16_23 (.BL(BL23),.BLN(BLN23),.WL(WL16));
sram_cell_6t_5 inst_cell_16_24 (.BL(BL24),.BLN(BLN24),.WL(WL16));
sram_cell_6t_5 inst_cell_16_25 (.BL(BL25),.BLN(BLN25),.WL(WL16));
sram_cell_6t_5 inst_cell_16_26 (.BL(BL26),.BLN(BLN26),.WL(WL16));
sram_cell_6t_5 inst_cell_16_27 (.BL(BL27),.BLN(BLN27),.WL(WL16));
sram_cell_6t_5 inst_cell_16_28 (.BL(BL28),.BLN(BLN28),.WL(WL16));
sram_cell_6t_5 inst_cell_16_29 (.BL(BL29),.BLN(BLN29),.WL(WL16));
sram_cell_6t_5 inst_cell_16_30 (.BL(BL30),.BLN(BLN30),.WL(WL16));
sram_cell_6t_5 inst_cell_16_31 (.BL(BL31),.BLN(BLN31),.WL(WL16));
sram_cell_6t_5 inst_cell_16_32 (.BL(BL32),.BLN(BLN32),.WL(WL16));
sram_cell_6t_5 inst_cell_16_33 (.BL(BL33),.BLN(BLN33),.WL(WL16));
sram_cell_6t_5 inst_cell_16_34 (.BL(BL34),.BLN(BLN34),.WL(WL16));
sram_cell_6t_5 inst_cell_16_35 (.BL(BL35),.BLN(BLN35),.WL(WL16));
sram_cell_6t_5 inst_cell_16_36 (.BL(BL36),.BLN(BLN36),.WL(WL16));
sram_cell_6t_5 inst_cell_16_37 (.BL(BL37),.BLN(BLN37),.WL(WL16));
sram_cell_6t_5 inst_cell_16_38 (.BL(BL38),.BLN(BLN38),.WL(WL16));
sram_cell_6t_5 inst_cell_16_39 (.BL(BL39),.BLN(BLN39),.WL(WL16));
sram_cell_6t_5 inst_cell_16_40 (.BL(BL40),.BLN(BLN40),.WL(WL16));
sram_cell_6t_5 inst_cell_16_41 (.BL(BL41),.BLN(BLN41),.WL(WL16));
sram_cell_6t_5 inst_cell_16_42 (.BL(BL42),.BLN(BLN42),.WL(WL16));
sram_cell_6t_5 inst_cell_16_43 (.BL(BL43),.BLN(BLN43),.WL(WL16));
sram_cell_6t_5 inst_cell_16_44 (.BL(BL44),.BLN(BLN44),.WL(WL16));
sram_cell_6t_5 inst_cell_16_45 (.BL(BL45),.BLN(BLN45),.WL(WL16));
sram_cell_6t_5 inst_cell_16_46 (.BL(BL46),.BLN(BLN46),.WL(WL16));
sram_cell_6t_5 inst_cell_16_47 (.BL(BL47),.BLN(BLN47),.WL(WL16));
sram_cell_6t_5 inst_cell_16_48 (.BL(BL48),.BLN(BLN48),.WL(WL16));
sram_cell_6t_5 inst_cell_16_49 (.BL(BL49),.BLN(BLN49),.WL(WL16));
sram_cell_6t_5 inst_cell_16_50 (.BL(BL50),.BLN(BLN50),.WL(WL16));
sram_cell_6t_5 inst_cell_16_51 (.BL(BL51),.BLN(BLN51),.WL(WL16));
sram_cell_6t_5 inst_cell_16_52 (.BL(BL52),.BLN(BLN52),.WL(WL16));
sram_cell_6t_5 inst_cell_16_53 (.BL(BL53),.BLN(BLN53),.WL(WL16));
sram_cell_6t_5 inst_cell_16_54 (.BL(BL54),.BLN(BLN54),.WL(WL16));
sram_cell_6t_5 inst_cell_16_55 (.BL(BL55),.BLN(BLN55),.WL(WL16));
sram_cell_6t_5 inst_cell_16_56 (.BL(BL56),.BLN(BLN56),.WL(WL16));
sram_cell_6t_5 inst_cell_16_57 (.BL(BL57),.BLN(BLN57),.WL(WL16));
sram_cell_6t_5 inst_cell_16_58 (.BL(BL58),.BLN(BLN58),.WL(WL16));
sram_cell_6t_5 inst_cell_16_59 (.BL(BL59),.BLN(BLN59),.WL(WL16));
sram_cell_6t_5 inst_cell_16_60 (.BL(BL60),.BLN(BLN60),.WL(WL16));
sram_cell_6t_5 inst_cell_16_61 (.BL(BL61),.BLN(BLN61),.WL(WL16));
sram_cell_6t_5 inst_cell_16_62 (.BL(BL62),.BLN(BLN62),.WL(WL16));
sram_cell_6t_5 inst_cell_16_63 (.BL(BL63),.BLN(BLN63),.WL(WL16));
sram_cell_6t_5 inst_cell_16_64 (.BL(BL64),.BLN(BLN64),.WL(WL16));
sram_cell_6t_5 inst_cell_16_65 (.BL(BL65),.BLN(BLN65),.WL(WL16));
sram_cell_6t_5 inst_cell_16_66 (.BL(BL66),.BLN(BLN66),.WL(WL16));
sram_cell_6t_5 inst_cell_16_67 (.BL(BL67),.BLN(BLN67),.WL(WL16));
sram_cell_6t_5 inst_cell_16_68 (.BL(BL68),.BLN(BLN68),.WL(WL16));
sram_cell_6t_5 inst_cell_16_69 (.BL(BL69),.BLN(BLN69),.WL(WL16));
sram_cell_6t_5 inst_cell_16_70 (.BL(BL70),.BLN(BLN70),.WL(WL16));
sram_cell_6t_5 inst_cell_16_71 (.BL(BL71),.BLN(BLN71),.WL(WL16));
sram_cell_6t_5 inst_cell_16_72 (.BL(BL72),.BLN(BLN72),.WL(WL16));
sram_cell_6t_5 inst_cell_16_73 (.BL(BL73),.BLN(BLN73),.WL(WL16));
sram_cell_6t_5 inst_cell_16_74 (.BL(BL74),.BLN(BLN74),.WL(WL16));
sram_cell_6t_5 inst_cell_16_75 (.BL(BL75),.BLN(BLN75),.WL(WL16));
sram_cell_6t_5 inst_cell_16_76 (.BL(BL76),.BLN(BLN76),.WL(WL16));
sram_cell_6t_5 inst_cell_16_77 (.BL(BL77),.BLN(BLN77),.WL(WL16));
sram_cell_6t_5 inst_cell_16_78 (.BL(BL78),.BLN(BLN78),.WL(WL16));
sram_cell_6t_5 inst_cell_16_79 (.BL(BL79),.BLN(BLN79),.WL(WL16));
sram_cell_6t_5 inst_cell_16_80 (.BL(BL80),.BLN(BLN80),.WL(WL16));
sram_cell_6t_5 inst_cell_16_81 (.BL(BL81),.BLN(BLN81),.WL(WL16));
sram_cell_6t_5 inst_cell_16_82 (.BL(BL82),.BLN(BLN82),.WL(WL16));
sram_cell_6t_5 inst_cell_16_83 (.BL(BL83),.BLN(BLN83),.WL(WL16));
sram_cell_6t_5 inst_cell_16_84 (.BL(BL84),.BLN(BLN84),.WL(WL16));
sram_cell_6t_5 inst_cell_16_85 (.BL(BL85),.BLN(BLN85),.WL(WL16));
sram_cell_6t_5 inst_cell_16_86 (.BL(BL86),.BLN(BLN86),.WL(WL16));
sram_cell_6t_5 inst_cell_16_87 (.BL(BL87),.BLN(BLN87),.WL(WL16));
sram_cell_6t_5 inst_cell_16_88 (.BL(BL88),.BLN(BLN88),.WL(WL16));
sram_cell_6t_5 inst_cell_16_89 (.BL(BL89),.BLN(BLN89),.WL(WL16));
sram_cell_6t_5 inst_cell_16_90 (.BL(BL90),.BLN(BLN90),.WL(WL16));
sram_cell_6t_5 inst_cell_16_91 (.BL(BL91),.BLN(BLN91),.WL(WL16));
sram_cell_6t_5 inst_cell_16_92 (.BL(BL92),.BLN(BLN92),.WL(WL16));
sram_cell_6t_5 inst_cell_16_93 (.BL(BL93),.BLN(BLN93),.WL(WL16));
sram_cell_6t_5 inst_cell_16_94 (.BL(BL94),.BLN(BLN94),.WL(WL16));
sram_cell_6t_5 inst_cell_16_95 (.BL(BL95),.BLN(BLN95),.WL(WL16));
sram_cell_6t_5 inst_cell_16_96 (.BL(BL96),.BLN(BLN96),.WL(WL16));
sram_cell_6t_5 inst_cell_16_97 (.BL(BL97),.BLN(BLN97),.WL(WL16));
sram_cell_6t_5 inst_cell_16_98 (.BL(BL98),.BLN(BLN98),.WL(WL16));
sram_cell_6t_5 inst_cell_16_99 (.BL(BL99),.BLN(BLN99),.WL(WL16));
sram_cell_6t_5 inst_cell_16_100 (.BL(BL100),.BLN(BLN100),.WL(WL16));
sram_cell_6t_5 inst_cell_16_101 (.BL(BL101),.BLN(BLN101),.WL(WL16));
sram_cell_6t_5 inst_cell_16_102 (.BL(BL102),.BLN(BLN102),.WL(WL16));
sram_cell_6t_5 inst_cell_16_103 (.BL(BL103),.BLN(BLN103),.WL(WL16));
sram_cell_6t_5 inst_cell_16_104 (.BL(BL104),.BLN(BLN104),.WL(WL16));
sram_cell_6t_5 inst_cell_16_105 (.BL(BL105),.BLN(BLN105),.WL(WL16));
sram_cell_6t_5 inst_cell_16_106 (.BL(BL106),.BLN(BLN106),.WL(WL16));
sram_cell_6t_5 inst_cell_16_107 (.BL(BL107),.BLN(BLN107),.WL(WL16));
sram_cell_6t_5 inst_cell_16_108 (.BL(BL108),.BLN(BLN108),.WL(WL16));
sram_cell_6t_5 inst_cell_16_109 (.BL(BL109),.BLN(BLN109),.WL(WL16));
sram_cell_6t_5 inst_cell_16_110 (.BL(BL110),.BLN(BLN110),.WL(WL16));
sram_cell_6t_5 inst_cell_16_111 (.BL(BL111),.BLN(BLN111),.WL(WL16));
sram_cell_6t_5 inst_cell_16_112 (.BL(BL112),.BLN(BLN112),.WL(WL16));
sram_cell_6t_5 inst_cell_16_113 (.BL(BL113),.BLN(BLN113),.WL(WL16));
sram_cell_6t_5 inst_cell_16_114 (.BL(BL114),.BLN(BLN114),.WL(WL16));
sram_cell_6t_5 inst_cell_16_115 (.BL(BL115),.BLN(BLN115),.WL(WL16));
sram_cell_6t_5 inst_cell_16_116 (.BL(BL116),.BLN(BLN116),.WL(WL16));
sram_cell_6t_5 inst_cell_16_117 (.BL(BL117),.BLN(BLN117),.WL(WL16));
sram_cell_6t_5 inst_cell_16_118 (.BL(BL118),.BLN(BLN118),.WL(WL16));
sram_cell_6t_5 inst_cell_16_119 (.BL(BL119),.BLN(BLN119),.WL(WL16));
sram_cell_6t_5 inst_cell_16_120 (.BL(BL120),.BLN(BLN120),.WL(WL16));
sram_cell_6t_5 inst_cell_16_121 (.BL(BL121),.BLN(BLN121),.WL(WL16));
sram_cell_6t_5 inst_cell_16_122 (.BL(BL122),.BLN(BLN122),.WL(WL16));
sram_cell_6t_5 inst_cell_16_123 (.BL(BL123),.BLN(BLN123),.WL(WL16));
sram_cell_6t_5 inst_cell_16_124 (.BL(BL124),.BLN(BLN124),.WL(WL16));
sram_cell_6t_5 inst_cell_16_125 (.BL(BL125),.BLN(BLN125),.WL(WL16));
sram_cell_6t_5 inst_cell_16_126 (.BL(BL126),.BLN(BLN126),.WL(WL16));
sram_cell_6t_5 inst_cell_16_127 (.BL(BL127),.BLN(BLN127),.WL(WL16));
sram_cell_6t_5 inst_cell_17_0 (.BL(BL0),.BLN(BLN0),.WL(WL17));
sram_cell_6t_5 inst_cell_17_1 (.BL(BL1),.BLN(BLN1),.WL(WL17));
sram_cell_6t_5 inst_cell_17_2 (.BL(BL2),.BLN(BLN2),.WL(WL17));
sram_cell_6t_5 inst_cell_17_3 (.BL(BL3),.BLN(BLN3),.WL(WL17));
sram_cell_6t_5 inst_cell_17_4 (.BL(BL4),.BLN(BLN4),.WL(WL17));
sram_cell_6t_5 inst_cell_17_5 (.BL(BL5),.BLN(BLN5),.WL(WL17));
sram_cell_6t_5 inst_cell_17_6 (.BL(BL6),.BLN(BLN6),.WL(WL17));
sram_cell_6t_5 inst_cell_17_7 (.BL(BL7),.BLN(BLN7),.WL(WL17));
sram_cell_6t_5 inst_cell_17_8 (.BL(BL8),.BLN(BLN8),.WL(WL17));
sram_cell_6t_5 inst_cell_17_9 (.BL(BL9),.BLN(BLN9),.WL(WL17));
sram_cell_6t_5 inst_cell_17_10 (.BL(BL10),.BLN(BLN10),.WL(WL17));
sram_cell_6t_5 inst_cell_17_11 (.BL(BL11),.BLN(BLN11),.WL(WL17));
sram_cell_6t_5 inst_cell_17_12 (.BL(BL12),.BLN(BLN12),.WL(WL17));
sram_cell_6t_5 inst_cell_17_13 (.BL(BL13),.BLN(BLN13),.WL(WL17));
sram_cell_6t_5 inst_cell_17_14 (.BL(BL14),.BLN(BLN14),.WL(WL17));
sram_cell_6t_5 inst_cell_17_15 (.BL(BL15),.BLN(BLN15),.WL(WL17));
sram_cell_6t_5 inst_cell_17_16 (.BL(BL16),.BLN(BLN16),.WL(WL17));
sram_cell_6t_5 inst_cell_17_17 (.BL(BL17),.BLN(BLN17),.WL(WL17));
sram_cell_6t_5 inst_cell_17_18 (.BL(BL18),.BLN(BLN18),.WL(WL17));
sram_cell_6t_5 inst_cell_17_19 (.BL(BL19),.BLN(BLN19),.WL(WL17));
sram_cell_6t_5 inst_cell_17_20 (.BL(BL20),.BLN(BLN20),.WL(WL17));
sram_cell_6t_5 inst_cell_17_21 (.BL(BL21),.BLN(BLN21),.WL(WL17));
sram_cell_6t_5 inst_cell_17_22 (.BL(BL22),.BLN(BLN22),.WL(WL17));
sram_cell_6t_5 inst_cell_17_23 (.BL(BL23),.BLN(BLN23),.WL(WL17));
sram_cell_6t_5 inst_cell_17_24 (.BL(BL24),.BLN(BLN24),.WL(WL17));
sram_cell_6t_5 inst_cell_17_25 (.BL(BL25),.BLN(BLN25),.WL(WL17));
sram_cell_6t_5 inst_cell_17_26 (.BL(BL26),.BLN(BLN26),.WL(WL17));
sram_cell_6t_5 inst_cell_17_27 (.BL(BL27),.BLN(BLN27),.WL(WL17));
sram_cell_6t_5 inst_cell_17_28 (.BL(BL28),.BLN(BLN28),.WL(WL17));
sram_cell_6t_5 inst_cell_17_29 (.BL(BL29),.BLN(BLN29),.WL(WL17));
sram_cell_6t_5 inst_cell_17_30 (.BL(BL30),.BLN(BLN30),.WL(WL17));
sram_cell_6t_5 inst_cell_17_31 (.BL(BL31),.BLN(BLN31),.WL(WL17));
sram_cell_6t_5 inst_cell_17_32 (.BL(BL32),.BLN(BLN32),.WL(WL17));
sram_cell_6t_5 inst_cell_17_33 (.BL(BL33),.BLN(BLN33),.WL(WL17));
sram_cell_6t_5 inst_cell_17_34 (.BL(BL34),.BLN(BLN34),.WL(WL17));
sram_cell_6t_5 inst_cell_17_35 (.BL(BL35),.BLN(BLN35),.WL(WL17));
sram_cell_6t_5 inst_cell_17_36 (.BL(BL36),.BLN(BLN36),.WL(WL17));
sram_cell_6t_5 inst_cell_17_37 (.BL(BL37),.BLN(BLN37),.WL(WL17));
sram_cell_6t_5 inst_cell_17_38 (.BL(BL38),.BLN(BLN38),.WL(WL17));
sram_cell_6t_5 inst_cell_17_39 (.BL(BL39),.BLN(BLN39),.WL(WL17));
sram_cell_6t_5 inst_cell_17_40 (.BL(BL40),.BLN(BLN40),.WL(WL17));
sram_cell_6t_5 inst_cell_17_41 (.BL(BL41),.BLN(BLN41),.WL(WL17));
sram_cell_6t_5 inst_cell_17_42 (.BL(BL42),.BLN(BLN42),.WL(WL17));
sram_cell_6t_5 inst_cell_17_43 (.BL(BL43),.BLN(BLN43),.WL(WL17));
sram_cell_6t_5 inst_cell_17_44 (.BL(BL44),.BLN(BLN44),.WL(WL17));
sram_cell_6t_5 inst_cell_17_45 (.BL(BL45),.BLN(BLN45),.WL(WL17));
sram_cell_6t_5 inst_cell_17_46 (.BL(BL46),.BLN(BLN46),.WL(WL17));
sram_cell_6t_5 inst_cell_17_47 (.BL(BL47),.BLN(BLN47),.WL(WL17));
sram_cell_6t_5 inst_cell_17_48 (.BL(BL48),.BLN(BLN48),.WL(WL17));
sram_cell_6t_5 inst_cell_17_49 (.BL(BL49),.BLN(BLN49),.WL(WL17));
sram_cell_6t_5 inst_cell_17_50 (.BL(BL50),.BLN(BLN50),.WL(WL17));
sram_cell_6t_5 inst_cell_17_51 (.BL(BL51),.BLN(BLN51),.WL(WL17));
sram_cell_6t_5 inst_cell_17_52 (.BL(BL52),.BLN(BLN52),.WL(WL17));
sram_cell_6t_5 inst_cell_17_53 (.BL(BL53),.BLN(BLN53),.WL(WL17));
sram_cell_6t_5 inst_cell_17_54 (.BL(BL54),.BLN(BLN54),.WL(WL17));
sram_cell_6t_5 inst_cell_17_55 (.BL(BL55),.BLN(BLN55),.WL(WL17));
sram_cell_6t_5 inst_cell_17_56 (.BL(BL56),.BLN(BLN56),.WL(WL17));
sram_cell_6t_5 inst_cell_17_57 (.BL(BL57),.BLN(BLN57),.WL(WL17));
sram_cell_6t_5 inst_cell_17_58 (.BL(BL58),.BLN(BLN58),.WL(WL17));
sram_cell_6t_5 inst_cell_17_59 (.BL(BL59),.BLN(BLN59),.WL(WL17));
sram_cell_6t_5 inst_cell_17_60 (.BL(BL60),.BLN(BLN60),.WL(WL17));
sram_cell_6t_5 inst_cell_17_61 (.BL(BL61),.BLN(BLN61),.WL(WL17));
sram_cell_6t_5 inst_cell_17_62 (.BL(BL62),.BLN(BLN62),.WL(WL17));
sram_cell_6t_5 inst_cell_17_63 (.BL(BL63),.BLN(BLN63),.WL(WL17));
sram_cell_6t_5 inst_cell_17_64 (.BL(BL64),.BLN(BLN64),.WL(WL17));
sram_cell_6t_5 inst_cell_17_65 (.BL(BL65),.BLN(BLN65),.WL(WL17));
sram_cell_6t_5 inst_cell_17_66 (.BL(BL66),.BLN(BLN66),.WL(WL17));
sram_cell_6t_5 inst_cell_17_67 (.BL(BL67),.BLN(BLN67),.WL(WL17));
sram_cell_6t_5 inst_cell_17_68 (.BL(BL68),.BLN(BLN68),.WL(WL17));
sram_cell_6t_5 inst_cell_17_69 (.BL(BL69),.BLN(BLN69),.WL(WL17));
sram_cell_6t_5 inst_cell_17_70 (.BL(BL70),.BLN(BLN70),.WL(WL17));
sram_cell_6t_5 inst_cell_17_71 (.BL(BL71),.BLN(BLN71),.WL(WL17));
sram_cell_6t_5 inst_cell_17_72 (.BL(BL72),.BLN(BLN72),.WL(WL17));
sram_cell_6t_5 inst_cell_17_73 (.BL(BL73),.BLN(BLN73),.WL(WL17));
sram_cell_6t_5 inst_cell_17_74 (.BL(BL74),.BLN(BLN74),.WL(WL17));
sram_cell_6t_5 inst_cell_17_75 (.BL(BL75),.BLN(BLN75),.WL(WL17));
sram_cell_6t_5 inst_cell_17_76 (.BL(BL76),.BLN(BLN76),.WL(WL17));
sram_cell_6t_5 inst_cell_17_77 (.BL(BL77),.BLN(BLN77),.WL(WL17));
sram_cell_6t_5 inst_cell_17_78 (.BL(BL78),.BLN(BLN78),.WL(WL17));
sram_cell_6t_5 inst_cell_17_79 (.BL(BL79),.BLN(BLN79),.WL(WL17));
sram_cell_6t_5 inst_cell_17_80 (.BL(BL80),.BLN(BLN80),.WL(WL17));
sram_cell_6t_5 inst_cell_17_81 (.BL(BL81),.BLN(BLN81),.WL(WL17));
sram_cell_6t_5 inst_cell_17_82 (.BL(BL82),.BLN(BLN82),.WL(WL17));
sram_cell_6t_5 inst_cell_17_83 (.BL(BL83),.BLN(BLN83),.WL(WL17));
sram_cell_6t_5 inst_cell_17_84 (.BL(BL84),.BLN(BLN84),.WL(WL17));
sram_cell_6t_5 inst_cell_17_85 (.BL(BL85),.BLN(BLN85),.WL(WL17));
sram_cell_6t_5 inst_cell_17_86 (.BL(BL86),.BLN(BLN86),.WL(WL17));
sram_cell_6t_5 inst_cell_17_87 (.BL(BL87),.BLN(BLN87),.WL(WL17));
sram_cell_6t_5 inst_cell_17_88 (.BL(BL88),.BLN(BLN88),.WL(WL17));
sram_cell_6t_5 inst_cell_17_89 (.BL(BL89),.BLN(BLN89),.WL(WL17));
sram_cell_6t_5 inst_cell_17_90 (.BL(BL90),.BLN(BLN90),.WL(WL17));
sram_cell_6t_5 inst_cell_17_91 (.BL(BL91),.BLN(BLN91),.WL(WL17));
sram_cell_6t_5 inst_cell_17_92 (.BL(BL92),.BLN(BLN92),.WL(WL17));
sram_cell_6t_5 inst_cell_17_93 (.BL(BL93),.BLN(BLN93),.WL(WL17));
sram_cell_6t_5 inst_cell_17_94 (.BL(BL94),.BLN(BLN94),.WL(WL17));
sram_cell_6t_5 inst_cell_17_95 (.BL(BL95),.BLN(BLN95),.WL(WL17));
sram_cell_6t_5 inst_cell_17_96 (.BL(BL96),.BLN(BLN96),.WL(WL17));
sram_cell_6t_5 inst_cell_17_97 (.BL(BL97),.BLN(BLN97),.WL(WL17));
sram_cell_6t_5 inst_cell_17_98 (.BL(BL98),.BLN(BLN98),.WL(WL17));
sram_cell_6t_5 inst_cell_17_99 (.BL(BL99),.BLN(BLN99),.WL(WL17));
sram_cell_6t_5 inst_cell_17_100 (.BL(BL100),.BLN(BLN100),.WL(WL17));
sram_cell_6t_5 inst_cell_17_101 (.BL(BL101),.BLN(BLN101),.WL(WL17));
sram_cell_6t_5 inst_cell_17_102 (.BL(BL102),.BLN(BLN102),.WL(WL17));
sram_cell_6t_5 inst_cell_17_103 (.BL(BL103),.BLN(BLN103),.WL(WL17));
sram_cell_6t_5 inst_cell_17_104 (.BL(BL104),.BLN(BLN104),.WL(WL17));
sram_cell_6t_5 inst_cell_17_105 (.BL(BL105),.BLN(BLN105),.WL(WL17));
sram_cell_6t_5 inst_cell_17_106 (.BL(BL106),.BLN(BLN106),.WL(WL17));
sram_cell_6t_5 inst_cell_17_107 (.BL(BL107),.BLN(BLN107),.WL(WL17));
sram_cell_6t_5 inst_cell_17_108 (.BL(BL108),.BLN(BLN108),.WL(WL17));
sram_cell_6t_5 inst_cell_17_109 (.BL(BL109),.BLN(BLN109),.WL(WL17));
sram_cell_6t_5 inst_cell_17_110 (.BL(BL110),.BLN(BLN110),.WL(WL17));
sram_cell_6t_5 inst_cell_17_111 (.BL(BL111),.BLN(BLN111),.WL(WL17));
sram_cell_6t_5 inst_cell_17_112 (.BL(BL112),.BLN(BLN112),.WL(WL17));
sram_cell_6t_5 inst_cell_17_113 (.BL(BL113),.BLN(BLN113),.WL(WL17));
sram_cell_6t_5 inst_cell_17_114 (.BL(BL114),.BLN(BLN114),.WL(WL17));
sram_cell_6t_5 inst_cell_17_115 (.BL(BL115),.BLN(BLN115),.WL(WL17));
sram_cell_6t_5 inst_cell_17_116 (.BL(BL116),.BLN(BLN116),.WL(WL17));
sram_cell_6t_5 inst_cell_17_117 (.BL(BL117),.BLN(BLN117),.WL(WL17));
sram_cell_6t_5 inst_cell_17_118 (.BL(BL118),.BLN(BLN118),.WL(WL17));
sram_cell_6t_5 inst_cell_17_119 (.BL(BL119),.BLN(BLN119),.WL(WL17));
sram_cell_6t_5 inst_cell_17_120 (.BL(BL120),.BLN(BLN120),.WL(WL17));
sram_cell_6t_5 inst_cell_17_121 (.BL(BL121),.BLN(BLN121),.WL(WL17));
sram_cell_6t_5 inst_cell_17_122 (.BL(BL122),.BLN(BLN122),.WL(WL17));
sram_cell_6t_5 inst_cell_17_123 (.BL(BL123),.BLN(BLN123),.WL(WL17));
sram_cell_6t_5 inst_cell_17_124 (.BL(BL124),.BLN(BLN124),.WL(WL17));
sram_cell_6t_5 inst_cell_17_125 (.BL(BL125),.BLN(BLN125),.WL(WL17));
sram_cell_6t_5 inst_cell_17_126 (.BL(BL126),.BLN(BLN126),.WL(WL17));
sram_cell_6t_5 inst_cell_17_127 (.BL(BL127),.BLN(BLN127),.WL(WL17));
sram_cell_6t_5 inst_cell_18_0 (.BL(BL0),.BLN(BLN0),.WL(WL18));
sram_cell_6t_5 inst_cell_18_1 (.BL(BL1),.BLN(BLN1),.WL(WL18));
sram_cell_6t_5 inst_cell_18_2 (.BL(BL2),.BLN(BLN2),.WL(WL18));
sram_cell_6t_5 inst_cell_18_3 (.BL(BL3),.BLN(BLN3),.WL(WL18));
sram_cell_6t_5 inst_cell_18_4 (.BL(BL4),.BLN(BLN4),.WL(WL18));
sram_cell_6t_5 inst_cell_18_5 (.BL(BL5),.BLN(BLN5),.WL(WL18));
sram_cell_6t_5 inst_cell_18_6 (.BL(BL6),.BLN(BLN6),.WL(WL18));
sram_cell_6t_5 inst_cell_18_7 (.BL(BL7),.BLN(BLN7),.WL(WL18));
sram_cell_6t_5 inst_cell_18_8 (.BL(BL8),.BLN(BLN8),.WL(WL18));
sram_cell_6t_5 inst_cell_18_9 (.BL(BL9),.BLN(BLN9),.WL(WL18));
sram_cell_6t_5 inst_cell_18_10 (.BL(BL10),.BLN(BLN10),.WL(WL18));
sram_cell_6t_5 inst_cell_18_11 (.BL(BL11),.BLN(BLN11),.WL(WL18));
sram_cell_6t_5 inst_cell_18_12 (.BL(BL12),.BLN(BLN12),.WL(WL18));
sram_cell_6t_5 inst_cell_18_13 (.BL(BL13),.BLN(BLN13),.WL(WL18));
sram_cell_6t_5 inst_cell_18_14 (.BL(BL14),.BLN(BLN14),.WL(WL18));
sram_cell_6t_5 inst_cell_18_15 (.BL(BL15),.BLN(BLN15),.WL(WL18));
sram_cell_6t_5 inst_cell_18_16 (.BL(BL16),.BLN(BLN16),.WL(WL18));
sram_cell_6t_5 inst_cell_18_17 (.BL(BL17),.BLN(BLN17),.WL(WL18));
sram_cell_6t_5 inst_cell_18_18 (.BL(BL18),.BLN(BLN18),.WL(WL18));
sram_cell_6t_5 inst_cell_18_19 (.BL(BL19),.BLN(BLN19),.WL(WL18));
sram_cell_6t_5 inst_cell_18_20 (.BL(BL20),.BLN(BLN20),.WL(WL18));
sram_cell_6t_5 inst_cell_18_21 (.BL(BL21),.BLN(BLN21),.WL(WL18));
sram_cell_6t_5 inst_cell_18_22 (.BL(BL22),.BLN(BLN22),.WL(WL18));
sram_cell_6t_5 inst_cell_18_23 (.BL(BL23),.BLN(BLN23),.WL(WL18));
sram_cell_6t_5 inst_cell_18_24 (.BL(BL24),.BLN(BLN24),.WL(WL18));
sram_cell_6t_5 inst_cell_18_25 (.BL(BL25),.BLN(BLN25),.WL(WL18));
sram_cell_6t_5 inst_cell_18_26 (.BL(BL26),.BLN(BLN26),.WL(WL18));
sram_cell_6t_5 inst_cell_18_27 (.BL(BL27),.BLN(BLN27),.WL(WL18));
sram_cell_6t_5 inst_cell_18_28 (.BL(BL28),.BLN(BLN28),.WL(WL18));
sram_cell_6t_5 inst_cell_18_29 (.BL(BL29),.BLN(BLN29),.WL(WL18));
sram_cell_6t_5 inst_cell_18_30 (.BL(BL30),.BLN(BLN30),.WL(WL18));
sram_cell_6t_5 inst_cell_18_31 (.BL(BL31),.BLN(BLN31),.WL(WL18));
sram_cell_6t_5 inst_cell_18_32 (.BL(BL32),.BLN(BLN32),.WL(WL18));
sram_cell_6t_5 inst_cell_18_33 (.BL(BL33),.BLN(BLN33),.WL(WL18));
sram_cell_6t_5 inst_cell_18_34 (.BL(BL34),.BLN(BLN34),.WL(WL18));
sram_cell_6t_5 inst_cell_18_35 (.BL(BL35),.BLN(BLN35),.WL(WL18));
sram_cell_6t_5 inst_cell_18_36 (.BL(BL36),.BLN(BLN36),.WL(WL18));
sram_cell_6t_5 inst_cell_18_37 (.BL(BL37),.BLN(BLN37),.WL(WL18));
sram_cell_6t_5 inst_cell_18_38 (.BL(BL38),.BLN(BLN38),.WL(WL18));
sram_cell_6t_5 inst_cell_18_39 (.BL(BL39),.BLN(BLN39),.WL(WL18));
sram_cell_6t_5 inst_cell_18_40 (.BL(BL40),.BLN(BLN40),.WL(WL18));
sram_cell_6t_5 inst_cell_18_41 (.BL(BL41),.BLN(BLN41),.WL(WL18));
sram_cell_6t_5 inst_cell_18_42 (.BL(BL42),.BLN(BLN42),.WL(WL18));
sram_cell_6t_5 inst_cell_18_43 (.BL(BL43),.BLN(BLN43),.WL(WL18));
sram_cell_6t_5 inst_cell_18_44 (.BL(BL44),.BLN(BLN44),.WL(WL18));
sram_cell_6t_5 inst_cell_18_45 (.BL(BL45),.BLN(BLN45),.WL(WL18));
sram_cell_6t_5 inst_cell_18_46 (.BL(BL46),.BLN(BLN46),.WL(WL18));
sram_cell_6t_5 inst_cell_18_47 (.BL(BL47),.BLN(BLN47),.WL(WL18));
sram_cell_6t_5 inst_cell_18_48 (.BL(BL48),.BLN(BLN48),.WL(WL18));
sram_cell_6t_5 inst_cell_18_49 (.BL(BL49),.BLN(BLN49),.WL(WL18));
sram_cell_6t_5 inst_cell_18_50 (.BL(BL50),.BLN(BLN50),.WL(WL18));
sram_cell_6t_5 inst_cell_18_51 (.BL(BL51),.BLN(BLN51),.WL(WL18));
sram_cell_6t_5 inst_cell_18_52 (.BL(BL52),.BLN(BLN52),.WL(WL18));
sram_cell_6t_5 inst_cell_18_53 (.BL(BL53),.BLN(BLN53),.WL(WL18));
sram_cell_6t_5 inst_cell_18_54 (.BL(BL54),.BLN(BLN54),.WL(WL18));
sram_cell_6t_5 inst_cell_18_55 (.BL(BL55),.BLN(BLN55),.WL(WL18));
sram_cell_6t_5 inst_cell_18_56 (.BL(BL56),.BLN(BLN56),.WL(WL18));
sram_cell_6t_5 inst_cell_18_57 (.BL(BL57),.BLN(BLN57),.WL(WL18));
sram_cell_6t_5 inst_cell_18_58 (.BL(BL58),.BLN(BLN58),.WL(WL18));
sram_cell_6t_5 inst_cell_18_59 (.BL(BL59),.BLN(BLN59),.WL(WL18));
sram_cell_6t_5 inst_cell_18_60 (.BL(BL60),.BLN(BLN60),.WL(WL18));
sram_cell_6t_5 inst_cell_18_61 (.BL(BL61),.BLN(BLN61),.WL(WL18));
sram_cell_6t_5 inst_cell_18_62 (.BL(BL62),.BLN(BLN62),.WL(WL18));
sram_cell_6t_5 inst_cell_18_63 (.BL(BL63),.BLN(BLN63),.WL(WL18));
sram_cell_6t_5 inst_cell_18_64 (.BL(BL64),.BLN(BLN64),.WL(WL18));
sram_cell_6t_5 inst_cell_18_65 (.BL(BL65),.BLN(BLN65),.WL(WL18));
sram_cell_6t_5 inst_cell_18_66 (.BL(BL66),.BLN(BLN66),.WL(WL18));
sram_cell_6t_5 inst_cell_18_67 (.BL(BL67),.BLN(BLN67),.WL(WL18));
sram_cell_6t_5 inst_cell_18_68 (.BL(BL68),.BLN(BLN68),.WL(WL18));
sram_cell_6t_5 inst_cell_18_69 (.BL(BL69),.BLN(BLN69),.WL(WL18));
sram_cell_6t_5 inst_cell_18_70 (.BL(BL70),.BLN(BLN70),.WL(WL18));
sram_cell_6t_5 inst_cell_18_71 (.BL(BL71),.BLN(BLN71),.WL(WL18));
sram_cell_6t_5 inst_cell_18_72 (.BL(BL72),.BLN(BLN72),.WL(WL18));
sram_cell_6t_5 inst_cell_18_73 (.BL(BL73),.BLN(BLN73),.WL(WL18));
sram_cell_6t_5 inst_cell_18_74 (.BL(BL74),.BLN(BLN74),.WL(WL18));
sram_cell_6t_5 inst_cell_18_75 (.BL(BL75),.BLN(BLN75),.WL(WL18));
sram_cell_6t_5 inst_cell_18_76 (.BL(BL76),.BLN(BLN76),.WL(WL18));
sram_cell_6t_5 inst_cell_18_77 (.BL(BL77),.BLN(BLN77),.WL(WL18));
sram_cell_6t_5 inst_cell_18_78 (.BL(BL78),.BLN(BLN78),.WL(WL18));
sram_cell_6t_5 inst_cell_18_79 (.BL(BL79),.BLN(BLN79),.WL(WL18));
sram_cell_6t_5 inst_cell_18_80 (.BL(BL80),.BLN(BLN80),.WL(WL18));
sram_cell_6t_5 inst_cell_18_81 (.BL(BL81),.BLN(BLN81),.WL(WL18));
sram_cell_6t_5 inst_cell_18_82 (.BL(BL82),.BLN(BLN82),.WL(WL18));
sram_cell_6t_5 inst_cell_18_83 (.BL(BL83),.BLN(BLN83),.WL(WL18));
sram_cell_6t_5 inst_cell_18_84 (.BL(BL84),.BLN(BLN84),.WL(WL18));
sram_cell_6t_5 inst_cell_18_85 (.BL(BL85),.BLN(BLN85),.WL(WL18));
sram_cell_6t_5 inst_cell_18_86 (.BL(BL86),.BLN(BLN86),.WL(WL18));
sram_cell_6t_5 inst_cell_18_87 (.BL(BL87),.BLN(BLN87),.WL(WL18));
sram_cell_6t_5 inst_cell_18_88 (.BL(BL88),.BLN(BLN88),.WL(WL18));
sram_cell_6t_5 inst_cell_18_89 (.BL(BL89),.BLN(BLN89),.WL(WL18));
sram_cell_6t_5 inst_cell_18_90 (.BL(BL90),.BLN(BLN90),.WL(WL18));
sram_cell_6t_5 inst_cell_18_91 (.BL(BL91),.BLN(BLN91),.WL(WL18));
sram_cell_6t_5 inst_cell_18_92 (.BL(BL92),.BLN(BLN92),.WL(WL18));
sram_cell_6t_5 inst_cell_18_93 (.BL(BL93),.BLN(BLN93),.WL(WL18));
sram_cell_6t_5 inst_cell_18_94 (.BL(BL94),.BLN(BLN94),.WL(WL18));
sram_cell_6t_5 inst_cell_18_95 (.BL(BL95),.BLN(BLN95),.WL(WL18));
sram_cell_6t_5 inst_cell_18_96 (.BL(BL96),.BLN(BLN96),.WL(WL18));
sram_cell_6t_5 inst_cell_18_97 (.BL(BL97),.BLN(BLN97),.WL(WL18));
sram_cell_6t_5 inst_cell_18_98 (.BL(BL98),.BLN(BLN98),.WL(WL18));
sram_cell_6t_5 inst_cell_18_99 (.BL(BL99),.BLN(BLN99),.WL(WL18));
sram_cell_6t_5 inst_cell_18_100 (.BL(BL100),.BLN(BLN100),.WL(WL18));
sram_cell_6t_5 inst_cell_18_101 (.BL(BL101),.BLN(BLN101),.WL(WL18));
sram_cell_6t_5 inst_cell_18_102 (.BL(BL102),.BLN(BLN102),.WL(WL18));
sram_cell_6t_5 inst_cell_18_103 (.BL(BL103),.BLN(BLN103),.WL(WL18));
sram_cell_6t_5 inst_cell_18_104 (.BL(BL104),.BLN(BLN104),.WL(WL18));
sram_cell_6t_5 inst_cell_18_105 (.BL(BL105),.BLN(BLN105),.WL(WL18));
sram_cell_6t_5 inst_cell_18_106 (.BL(BL106),.BLN(BLN106),.WL(WL18));
sram_cell_6t_5 inst_cell_18_107 (.BL(BL107),.BLN(BLN107),.WL(WL18));
sram_cell_6t_5 inst_cell_18_108 (.BL(BL108),.BLN(BLN108),.WL(WL18));
sram_cell_6t_5 inst_cell_18_109 (.BL(BL109),.BLN(BLN109),.WL(WL18));
sram_cell_6t_5 inst_cell_18_110 (.BL(BL110),.BLN(BLN110),.WL(WL18));
sram_cell_6t_5 inst_cell_18_111 (.BL(BL111),.BLN(BLN111),.WL(WL18));
sram_cell_6t_5 inst_cell_18_112 (.BL(BL112),.BLN(BLN112),.WL(WL18));
sram_cell_6t_5 inst_cell_18_113 (.BL(BL113),.BLN(BLN113),.WL(WL18));
sram_cell_6t_5 inst_cell_18_114 (.BL(BL114),.BLN(BLN114),.WL(WL18));
sram_cell_6t_5 inst_cell_18_115 (.BL(BL115),.BLN(BLN115),.WL(WL18));
sram_cell_6t_5 inst_cell_18_116 (.BL(BL116),.BLN(BLN116),.WL(WL18));
sram_cell_6t_5 inst_cell_18_117 (.BL(BL117),.BLN(BLN117),.WL(WL18));
sram_cell_6t_5 inst_cell_18_118 (.BL(BL118),.BLN(BLN118),.WL(WL18));
sram_cell_6t_5 inst_cell_18_119 (.BL(BL119),.BLN(BLN119),.WL(WL18));
sram_cell_6t_5 inst_cell_18_120 (.BL(BL120),.BLN(BLN120),.WL(WL18));
sram_cell_6t_5 inst_cell_18_121 (.BL(BL121),.BLN(BLN121),.WL(WL18));
sram_cell_6t_5 inst_cell_18_122 (.BL(BL122),.BLN(BLN122),.WL(WL18));
sram_cell_6t_5 inst_cell_18_123 (.BL(BL123),.BLN(BLN123),.WL(WL18));
sram_cell_6t_5 inst_cell_18_124 (.BL(BL124),.BLN(BLN124),.WL(WL18));
sram_cell_6t_5 inst_cell_18_125 (.BL(BL125),.BLN(BLN125),.WL(WL18));
sram_cell_6t_5 inst_cell_18_126 (.BL(BL126),.BLN(BLN126),.WL(WL18));
sram_cell_6t_5 inst_cell_18_127 (.BL(BL127),.BLN(BLN127),.WL(WL18));
sram_cell_6t_5 inst_cell_19_0 (.BL(BL0),.BLN(BLN0),.WL(WL19));
sram_cell_6t_5 inst_cell_19_1 (.BL(BL1),.BLN(BLN1),.WL(WL19));
sram_cell_6t_5 inst_cell_19_2 (.BL(BL2),.BLN(BLN2),.WL(WL19));
sram_cell_6t_5 inst_cell_19_3 (.BL(BL3),.BLN(BLN3),.WL(WL19));
sram_cell_6t_5 inst_cell_19_4 (.BL(BL4),.BLN(BLN4),.WL(WL19));
sram_cell_6t_5 inst_cell_19_5 (.BL(BL5),.BLN(BLN5),.WL(WL19));
sram_cell_6t_5 inst_cell_19_6 (.BL(BL6),.BLN(BLN6),.WL(WL19));
sram_cell_6t_5 inst_cell_19_7 (.BL(BL7),.BLN(BLN7),.WL(WL19));
sram_cell_6t_5 inst_cell_19_8 (.BL(BL8),.BLN(BLN8),.WL(WL19));
sram_cell_6t_5 inst_cell_19_9 (.BL(BL9),.BLN(BLN9),.WL(WL19));
sram_cell_6t_5 inst_cell_19_10 (.BL(BL10),.BLN(BLN10),.WL(WL19));
sram_cell_6t_5 inst_cell_19_11 (.BL(BL11),.BLN(BLN11),.WL(WL19));
sram_cell_6t_5 inst_cell_19_12 (.BL(BL12),.BLN(BLN12),.WL(WL19));
sram_cell_6t_5 inst_cell_19_13 (.BL(BL13),.BLN(BLN13),.WL(WL19));
sram_cell_6t_5 inst_cell_19_14 (.BL(BL14),.BLN(BLN14),.WL(WL19));
sram_cell_6t_5 inst_cell_19_15 (.BL(BL15),.BLN(BLN15),.WL(WL19));
sram_cell_6t_5 inst_cell_19_16 (.BL(BL16),.BLN(BLN16),.WL(WL19));
sram_cell_6t_5 inst_cell_19_17 (.BL(BL17),.BLN(BLN17),.WL(WL19));
sram_cell_6t_5 inst_cell_19_18 (.BL(BL18),.BLN(BLN18),.WL(WL19));
sram_cell_6t_5 inst_cell_19_19 (.BL(BL19),.BLN(BLN19),.WL(WL19));
sram_cell_6t_5 inst_cell_19_20 (.BL(BL20),.BLN(BLN20),.WL(WL19));
sram_cell_6t_5 inst_cell_19_21 (.BL(BL21),.BLN(BLN21),.WL(WL19));
sram_cell_6t_5 inst_cell_19_22 (.BL(BL22),.BLN(BLN22),.WL(WL19));
sram_cell_6t_5 inst_cell_19_23 (.BL(BL23),.BLN(BLN23),.WL(WL19));
sram_cell_6t_5 inst_cell_19_24 (.BL(BL24),.BLN(BLN24),.WL(WL19));
sram_cell_6t_5 inst_cell_19_25 (.BL(BL25),.BLN(BLN25),.WL(WL19));
sram_cell_6t_5 inst_cell_19_26 (.BL(BL26),.BLN(BLN26),.WL(WL19));
sram_cell_6t_5 inst_cell_19_27 (.BL(BL27),.BLN(BLN27),.WL(WL19));
sram_cell_6t_5 inst_cell_19_28 (.BL(BL28),.BLN(BLN28),.WL(WL19));
sram_cell_6t_5 inst_cell_19_29 (.BL(BL29),.BLN(BLN29),.WL(WL19));
sram_cell_6t_5 inst_cell_19_30 (.BL(BL30),.BLN(BLN30),.WL(WL19));
sram_cell_6t_5 inst_cell_19_31 (.BL(BL31),.BLN(BLN31),.WL(WL19));
sram_cell_6t_5 inst_cell_19_32 (.BL(BL32),.BLN(BLN32),.WL(WL19));
sram_cell_6t_5 inst_cell_19_33 (.BL(BL33),.BLN(BLN33),.WL(WL19));
sram_cell_6t_5 inst_cell_19_34 (.BL(BL34),.BLN(BLN34),.WL(WL19));
sram_cell_6t_5 inst_cell_19_35 (.BL(BL35),.BLN(BLN35),.WL(WL19));
sram_cell_6t_5 inst_cell_19_36 (.BL(BL36),.BLN(BLN36),.WL(WL19));
sram_cell_6t_5 inst_cell_19_37 (.BL(BL37),.BLN(BLN37),.WL(WL19));
sram_cell_6t_5 inst_cell_19_38 (.BL(BL38),.BLN(BLN38),.WL(WL19));
sram_cell_6t_5 inst_cell_19_39 (.BL(BL39),.BLN(BLN39),.WL(WL19));
sram_cell_6t_5 inst_cell_19_40 (.BL(BL40),.BLN(BLN40),.WL(WL19));
sram_cell_6t_5 inst_cell_19_41 (.BL(BL41),.BLN(BLN41),.WL(WL19));
sram_cell_6t_5 inst_cell_19_42 (.BL(BL42),.BLN(BLN42),.WL(WL19));
sram_cell_6t_5 inst_cell_19_43 (.BL(BL43),.BLN(BLN43),.WL(WL19));
sram_cell_6t_5 inst_cell_19_44 (.BL(BL44),.BLN(BLN44),.WL(WL19));
sram_cell_6t_5 inst_cell_19_45 (.BL(BL45),.BLN(BLN45),.WL(WL19));
sram_cell_6t_5 inst_cell_19_46 (.BL(BL46),.BLN(BLN46),.WL(WL19));
sram_cell_6t_5 inst_cell_19_47 (.BL(BL47),.BLN(BLN47),.WL(WL19));
sram_cell_6t_5 inst_cell_19_48 (.BL(BL48),.BLN(BLN48),.WL(WL19));
sram_cell_6t_5 inst_cell_19_49 (.BL(BL49),.BLN(BLN49),.WL(WL19));
sram_cell_6t_5 inst_cell_19_50 (.BL(BL50),.BLN(BLN50),.WL(WL19));
sram_cell_6t_5 inst_cell_19_51 (.BL(BL51),.BLN(BLN51),.WL(WL19));
sram_cell_6t_5 inst_cell_19_52 (.BL(BL52),.BLN(BLN52),.WL(WL19));
sram_cell_6t_5 inst_cell_19_53 (.BL(BL53),.BLN(BLN53),.WL(WL19));
sram_cell_6t_5 inst_cell_19_54 (.BL(BL54),.BLN(BLN54),.WL(WL19));
sram_cell_6t_5 inst_cell_19_55 (.BL(BL55),.BLN(BLN55),.WL(WL19));
sram_cell_6t_5 inst_cell_19_56 (.BL(BL56),.BLN(BLN56),.WL(WL19));
sram_cell_6t_5 inst_cell_19_57 (.BL(BL57),.BLN(BLN57),.WL(WL19));
sram_cell_6t_5 inst_cell_19_58 (.BL(BL58),.BLN(BLN58),.WL(WL19));
sram_cell_6t_5 inst_cell_19_59 (.BL(BL59),.BLN(BLN59),.WL(WL19));
sram_cell_6t_5 inst_cell_19_60 (.BL(BL60),.BLN(BLN60),.WL(WL19));
sram_cell_6t_5 inst_cell_19_61 (.BL(BL61),.BLN(BLN61),.WL(WL19));
sram_cell_6t_5 inst_cell_19_62 (.BL(BL62),.BLN(BLN62),.WL(WL19));
sram_cell_6t_5 inst_cell_19_63 (.BL(BL63),.BLN(BLN63),.WL(WL19));
sram_cell_6t_5 inst_cell_19_64 (.BL(BL64),.BLN(BLN64),.WL(WL19));
sram_cell_6t_5 inst_cell_19_65 (.BL(BL65),.BLN(BLN65),.WL(WL19));
sram_cell_6t_5 inst_cell_19_66 (.BL(BL66),.BLN(BLN66),.WL(WL19));
sram_cell_6t_5 inst_cell_19_67 (.BL(BL67),.BLN(BLN67),.WL(WL19));
sram_cell_6t_5 inst_cell_19_68 (.BL(BL68),.BLN(BLN68),.WL(WL19));
sram_cell_6t_5 inst_cell_19_69 (.BL(BL69),.BLN(BLN69),.WL(WL19));
sram_cell_6t_5 inst_cell_19_70 (.BL(BL70),.BLN(BLN70),.WL(WL19));
sram_cell_6t_5 inst_cell_19_71 (.BL(BL71),.BLN(BLN71),.WL(WL19));
sram_cell_6t_5 inst_cell_19_72 (.BL(BL72),.BLN(BLN72),.WL(WL19));
sram_cell_6t_5 inst_cell_19_73 (.BL(BL73),.BLN(BLN73),.WL(WL19));
sram_cell_6t_5 inst_cell_19_74 (.BL(BL74),.BLN(BLN74),.WL(WL19));
sram_cell_6t_5 inst_cell_19_75 (.BL(BL75),.BLN(BLN75),.WL(WL19));
sram_cell_6t_5 inst_cell_19_76 (.BL(BL76),.BLN(BLN76),.WL(WL19));
sram_cell_6t_5 inst_cell_19_77 (.BL(BL77),.BLN(BLN77),.WL(WL19));
sram_cell_6t_5 inst_cell_19_78 (.BL(BL78),.BLN(BLN78),.WL(WL19));
sram_cell_6t_5 inst_cell_19_79 (.BL(BL79),.BLN(BLN79),.WL(WL19));
sram_cell_6t_5 inst_cell_19_80 (.BL(BL80),.BLN(BLN80),.WL(WL19));
sram_cell_6t_5 inst_cell_19_81 (.BL(BL81),.BLN(BLN81),.WL(WL19));
sram_cell_6t_5 inst_cell_19_82 (.BL(BL82),.BLN(BLN82),.WL(WL19));
sram_cell_6t_5 inst_cell_19_83 (.BL(BL83),.BLN(BLN83),.WL(WL19));
sram_cell_6t_5 inst_cell_19_84 (.BL(BL84),.BLN(BLN84),.WL(WL19));
sram_cell_6t_5 inst_cell_19_85 (.BL(BL85),.BLN(BLN85),.WL(WL19));
sram_cell_6t_5 inst_cell_19_86 (.BL(BL86),.BLN(BLN86),.WL(WL19));
sram_cell_6t_5 inst_cell_19_87 (.BL(BL87),.BLN(BLN87),.WL(WL19));
sram_cell_6t_5 inst_cell_19_88 (.BL(BL88),.BLN(BLN88),.WL(WL19));
sram_cell_6t_5 inst_cell_19_89 (.BL(BL89),.BLN(BLN89),.WL(WL19));
sram_cell_6t_5 inst_cell_19_90 (.BL(BL90),.BLN(BLN90),.WL(WL19));
sram_cell_6t_5 inst_cell_19_91 (.BL(BL91),.BLN(BLN91),.WL(WL19));
sram_cell_6t_5 inst_cell_19_92 (.BL(BL92),.BLN(BLN92),.WL(WL19));
sram_cell_6t_5 inst_cell_19_93 (.BL(BL93),.BLN(BLN93),.WL(WL19));
sram_cell_6t_5 inst_cell_19_94 (.BL(BL94),.BLN(BLN94),.WL(WL19));
sram_cell_6t_5 inst_cell_19_95 (.BL(BL95),.BLN(BLN95),.WL(WL19));
sram_cell_6t_5 inst_cell_19_96 (.BL(BL96),.BLN(BLN96),.WL(WL19));
sram_cell_6t_5 inst_cell_19_97 (.BL(BL97),.BLN(BLN97),.WL(WL19));
sram_cell_6t_5 inst_cell_19_98 (.BL(BL98),.BLN(BLN98),.WL(WL19));
sram_cell_6t_5 inst_cell_19_99 (.BL(BL99),.BLN(BLN99),.WL(WL19));
sram_cell_6t_5 inst_cell_19_100 (.BL(BL100),.BLN(BLN100),.WL(WL19));
sram_cell_6t_5 inst_cell_19_101 (.BL(BL101),.BLN(BLN101),.WL(WL19));
sram_cell_6t_5 inst_cell_19_102 (.BL(BL102),.BLN(BLN102),.WL(WL19));
sram_cell_6t_5 inst_cell_19_103 (.BL(BL103),.BLN(BLN103),.WL(WL19));
sram_cell_6t_5 inst_cell_19_104 (.BL(BL104),.BLN(BLN104),.WL(WL19));
sram_cell_6t_5 inst_cell_19_105 (.BL(BL105),.BLN(BLN105),.WL(WL19));
sram_cell_6t_5 inst_cell_19_106 (.BL(BL106),.BLN(BLN106),.WL(WL19));
sram_cell_6t_5 inst_cell_19_107 (.BL(BL107),.BLN(BLN107),.WL(WL19));
sram_cell_6t_5 inst_cell_19_108 (.BL(BL108),.BLN(BLN108),.WL(WL19));
sram_cell_6t_5 inst_cell_19_109 (.BL(BL109),.BLN(BLN109),.WL(WL19));
sram_cell_6t_5 inst_cell_19_110 (.BL(BL110),.BLN(BLN110),.WL(WL19));
sram_cell_6t_5 inst_cell_19_111 (.BL(BL111),.BLN(BLN111),.WL(WL19));
sram_cell_6t_5 inst_cell_19_112 (.BL(BL112),.BLN(BLN112),.WL(WL19));
sram_cell_6t_5 inst_cell_19_113 (.BL(BL113),.BLN(BLN113),.WL(WL19));
sram_cell_6t_5 inst_cell_19_114 (.BL(BL114),.BLN(BLN114),.WL(WL19));
sram_cell_6t_5 inst_cell_19_115 (.BL(BL115),.BLN(BLN115),.WL(WL19));
sram_cell_6t_5 inst_cell_19_116 (.BL(BL116),.BLN(BLN116),.WL(WL19));
sram_cell_6t_5 inst_cell_19_117 (.BL(BL117),.BLN(BLN117),.WL(WL19));
sram_cell_6t_5 inst_cell_19_118 (.BL(BL118),.BLN(BLN118),.WL(WL19));
sram_cell_6t_5 inst_cell_19_119 (.BL(BL119),.BLN(BLN119),.WL(WL19));
sram_cell_6t_5 inst_cell_19_120 (.BL(BL120),.BLN(BLN120),.WL(WL19));
sram_cell_6t_5 inst_cell_19_121 (.BL(BL121),.BLN(BLN121),.WL(WL19));
sram_cell_6t_5 inst_cell_19_122 (.BL(BL122),.BLN(BLN122),.WL(WL19));
sram_cell_6t_5 inst_cell_19_123 (.BL(BL123),.BLN(BLN123),.WL(WL19));
sram_cell_6t_5 inst_cell_19_124 (.BL(BL124),.BLN(BLN124),.WL(WL19));
sram_cell_6t_5 inst_cell_19_125 (.BL(BL125),.BLN(BLN125),.WL(WL19));
sram_cell_6t_5 inst_cell_19_126 (.BL(BL126),.BLN(BLN126),.WL(WL19));
sram_cell_6t_5 inst_cell_19_127 (.BL(BL127),.BLN(BLN127),.WL(WL19));
sram_cell_6t_5 inst_cell_20_0 (.BL(BL0),.BLN(BLN0),.WL(WL20));
sram_cell_6t_5 inst_cell_20_1 (.BL(BL1),.BLN(BLN1),.WL(WL20));
sram_cell_6t_5 inst_cell_20_2 (.BL(BL2),.BLN(BLN2),.WL(WL20));
sram_cell_6t_5 inst_cell_20_3 (.BL(BL3),.BLN(BLN3),.WL(WL20));
sram_cell_6t_5 inst_cell_20_4 (.BL(BL4),.BLN(BLN4),.WL(WL20));
sram_cell_6t_5 inst_cell_20_5 (.BL(BL5),.BLN(BLN5),.WL(WL20));
sram_cell_6t_5 inst_cell_20_6 (.BL(BL6),.BLN(BLN6),.WL(WL20));
sram_cell_6t_5 inst_cell_20_7 (.BL(BL7),.BLN(BLN7),.WL(WL20));
sram_cell_6t_5 inst_cell_20_8 (.BL(BL8),.BLN(BLN8),.WL(WL20));
sram_cell_6t_5 inst_cell_20_9 (.BL(BL9),.BLN(BLN9),.WL(WL20));
sram_cell_6t_5 inst_cell_20_10 (.BL(BL10),.BLN(BLN10),.WL(WL20));
sram_cell_6t_5 inst_cell_20_11 (.BL(BL11),.BLN(BLN11),.WL(WL20));
sram_cell_6t_5 inst_cell_20_12 (.BL(BL12),.BLN(BLN12),.WL(WL20));
sram_cell_6t_5 inst_cell_20_13 (.BL(BL13),.BLN(BLN13),.WL(WL20));
sram_cell_6t_5 inst_cell_20_14 (.BL(BL14),.BLN(BLN14),.WL(WL20));
sram_cell_6t_5 inst_cell_20_15 (.BL(BL15),.BLN(BLN15),.WL(WL20));
sram_cell_6t_5 inst_cell_20_16 (.BL(BL16),.BLN(BLN16),.WL(WL20));
sram_cell_6t_5 inst_cell_20_17 (.BL(BL17),.BLN(BLN17),.WL(WL20));
sram_cell_6t_5 inst_cell_20_18 (.BL(BL18),.BLN(BLN18),.WL(WL20));
sram_cell_6t_5 inst_cell_20_19 (.BL(BL19),.BLN(BLN19),.WL(WL20));
sram_cell_6t_5 inst_cell_20_20 (.BL(BL20),.BLN(BLN20),.WL(WL20));
sram_cell_6t_5 inst_cell_20_21 (.BL(BL21),.BLN(BLN21),.WL(WL20));
sram_cell_6t_5 inst_cell_20_22 (.BL(BL22),.BLN(BLN22),.WL(WL20));
sram_cell_6t_5 inst_cell_20_23 (.BL(BL23),.BLN(BLN23),.WL(WL20));
sram_cell_6t_5 inst_cell_20_24 (.BL(BL24),.BLN(BLN24),.WL(WL20));
sram_cell_6t_5 inst_cell_20_25 (.BL(BL25),.BLN(BLN25),.WL(WL20));
sram_cell_6t_5 inst_cell_20_26 (.BL(BL26),.BLN(BLN26),.WL(WL20));
sram_cell_6t_5 inst_cell_20_27 (.BL(BL27),.BLN(BLN27),.WL(WL20));
sram_cell_6t_5 inst_cell_20_28 (.BL(BL28),.BLN(BLN28),.WL(WL20));
sram_cell_6t_5 inst_cell_20_29 (.BL(BL29),.BLN(BLN29),.WL(WL20));
sram_cell_6t_5 inst_cell_20_30 (.BL(BL30),.BLN(BLN30),.WL(WL20));
sram_cell_6t_5 inst_cell_20_31 (.BL(BL31),.BLN(BLN31),.WL(WL20));
sram_cell_6t_5 inst_cell_20_32 (.BL(BL32),.BLN(BLN32),.WL(WL20));
sram_cell_6t_5 inst_cell_20_33 (.BL(BL33),.BLN(BLN33),.WL(WL20));
sram_cell_6t_5 inst_cell_20_34 (.BL(BL34),.BLN(BLN34),.WL(WL20));
sram_cell_6t_5 inst_cell_20_35 (.BL(BL35),.BLN(BLN35),.WL(WL20));
sram_cell_6t_5 inst_cell_20_36 (.BL(BL36),.BLN(BLN36),.WL(WL20));
sram_cell_6t_5 inst_cell_20_37 (.BL(BL37),.BLN(BLN37),.WL(WL20));
sram_cell_6t_5 inst_cell_20_38 (.BL(BL38),.BLN(BLN38),.WL(WL20));
sram_cell_6t_5 inst_cell_20_39 (.BL(BL39),.BLN(BLN39),.WL(WL20));
sram_cell_6t_5 inst_cell_20_40 (.BL(BL40),.BLN(BLN40),.WL(WL20));
sram_cell_6t_5 inst_cell_20_41 (.BL(BL41),.BLN(BLN41),.WL(WL20));
sram_cell_6t_5 inst_cell_20_42 (.BL(BL42),.BLN(BLN42),.WL(WL20));
sram_cell_6t_5 inst_cell_20_43 (.BL(BL43),.BLN(BLN43),.WL(WL20));
sram_cell_6t_5 inst_cell_20_44 (.BL(BL44),.BLN(BLN44),.WL(WL20));
sram_cell_6t_5 inst_cell_20_45 (.BL(BL45),.BLN(BLN45),.WL(WL20));
sram_cell_6t_5 inst_cell_20_46 (.BL(BL46),.BLN(BLN46),.WL(WL20));
sram_cell_6t_5 inst_cell_20_47 (.BL(BL47),.BLN(BLN47),.WL(WL20));
sram_cell_6t_5 inst_cell_20_48 (.BL(BL48),.BLN(BLN48),.WL(WL20));
sram_cell_6t_5 inst_cell_20_49 (.BL(BL49),.BLN(BLN49),.WL(WL20));
sram_cell_6t_5 inst_cell_20_50 (.BL(BL50),.BLN(BLN50),.WL(WL20));
sram_cell_6t_5 inst_cell_20_51 (.BL(BL51),.BLN(BLN51),.WL(WL20));
sram_cell_6t_5 inst_cell_20_52 (.BL(BL52),.BLN(BLN52),.WL(WL20));
sram_cell_6t_5 inst_cell_20_53 (.BL(BL53),.BLN(BLN53),.WL(WL20));
sram_cell_6t_5 inst_cell_20_54 (.BL(BL54),.BLN(BLN54),.WL(WL20));
sram_cell_6t_5 inst_cell_20_55 (.BL(BL55),.BLN(BLN55),.WL(WL20));
sram_cell_6t_5 inst_cell_20_56 (.BL(BL56),.BLN(BLN56),.WL(WL20));
sram_cell_6t_5 inst_cell_20_57 (.BL(BL57),.BLN(BLN57),.WL(WL20));
sram_cell_6t_5 inst_cell_20_58 (.BL(BL58),.BLN(BLN58),.WL(WL20));
sram_cell_6t_5 inst_cell_20_59 (.BL(BL59),.BLN(BLN59),.WL(WL20));
sram_cell_6t_5 inst_cell_20_60 (.BL(BL60),.BLN(BLN60),.WL(WL20));
sram_cell_6t_5 inst_cell_20_61 (.BL(BL61),.BLN(BLN61),.WL(WL20));
sram_cell_6t_5 inst_cell_20_62 (.BL(BL62),.BLN(BLN62),.WL(WL20));
sram_cell_6t_5 inst_cell_20_63 (.BL(BL63),.BLN(BLN63),.WL(WL20));
sram_cell_6t_5 inst_cell_20_64 (.BL(BL64),.BLN(BLN64),.WL(WL20));
sram_cell_6t_5 inst_cell_20_65 (.BL(BL65),.BLN(BLN65),.WL(WL20));
sram_cell_6t_5 inst_cell_20_66 (.BL(BL66),.BLN(BLN66),.WL(WL20));
sram_cell_6t_5 inst_cell_20_67 (.BL(BL67),.BLN(BLN67),.WL(WL20));
sram_cell_6t_5 inst_cell_20_68 (.BL(BL68),.BLN(BLN68),.WL(WL20));
sram_cell_6t_5 inst_cell_20_69 (.BL(BL69),.BLN(BLN69),.WL(WL20));
sram_cell_6t_5 inst_cell_20_70 (.BL(BL70),.BLN(BLN70),.WL(WL20));
sram_cell_6t_5 inst_cell_20_71 (.BL(BL71),.BLN(BLN71),.WL(WL20));
sram_cell_6t_5 inst_cell_20_72 (.BL(BL72),.BLN(BLN72),.WL(WL20));
sram_cell_6t_5 inst_cell_20_73 (.BL(BL73),.BLN(BLN73),.WL(WL20));
sram_cell_6t_5 inst_cell_20_74 (.BL(BL74),.BLN(BLN74),.WL(WL20));
sram_cell_6t_5 inst_cell_20_75 (.BL(BL75),.BLN(BLN75),.WL(WL20));
sram_cell_6t_5 inst_cell_20_76 (.BL(BL76),.BLN(BLN76),.WL(WL20));
sram_cell_6t_5 inst_cell_20_77 (.BL(BL77),.BLN(BLN77),.WL(WL20));
sram_cell_6t_5 inst_cell_20_78 (.BL(BL78),.BLN(BLN78),.WL(WL20));
sram_cell_6t_5 inst_cell_20_79 (.BL(BL79),.BLN(BLN79),.WL(WL20));
sram_cell_6t_5 inst_cell_20_80 (.BL(BL80),.BLN(BLN80),.WL(WL20));
sram_cell_6t_5 inst_cell_20_81 (.BL(BL81),.BLN(BLN81),.WL(WL20));
sram_cell_6t_5 inst_cell_20_82 (.BL(BL82),.BLN(BLN82),.WL(WL20));
sram_cell_6t_5 inst_cell_20_83 (.BL(BL83),.BLN(BLN83),.WL(WL20));
sram_cell_6t_5 inst_cell_20_84 (.BL(BL84),.BLN(BLN84),.WL(WL20));
sram_cell_6t_5 inst_cell_20_85 (.BL(BL85),.BLN(BLN85),.WL(WL20));
sram_cell_6t_5 inst_cell_20_86 (.BL(BL86),.BLN(BLN86),.WL(WL20));
sram_cell_6t_5 inst_cell_20_87 (.BL(BL87),.BLN(BLN87),.WL(WL20));
sram_cell_6t_5 inst_cell_20_88 (.BL(BL88),.BLN(BLN88),.WL(WL20));
sram_cell_6t_5 inst_cell_20_89 (.BL(BL89),.BLN(BLN89),.WL(WL20));
sram_cell_6t_5 inst_cell_20_90 (.BL(BL90),.BLN(BLN90),.WL(WL20));
sram_cell_6t_5 inst_cell_20_91 (.BL(BL91),.BLN(BLN91),.WL(WL20));
sram_cell_6t_5 inst_cell_20_92 (.BL(BL92),.BLN(BLN92),.WL(WL20));
sram_cell_6t_5 inst_cell_20_93 (.BL(BL93),.BLN(BLN93),.WL(WL20));
sram_cell_6t_5 inst_cell_20_94 (.BL(BL94),.BLN(BLN94),.WL(WL20));
sram_cell_6t_5 inst_cell_20_95 (.BL(BL95),.BLN(BLN95),.WL(WL20));
sram_cell_6t_5 inst_cell_20_96 (.BL(BL96),.BLN(BLN96),.WL(WL20));
sram_cell_6t_5 inst_cell_20_97 (.BL(BL97),.BLN(BLN97),.WL(WL20));
sram_cell_6t_5 inst_cell_20_98 (.BL(BL98),.BLN(BLN98),.WL(WL20));
sram_cell_6t_5 inst_cell_20_99 (.BL(BL99),.BLN(BLN99),.WL(WL20));
sram_cell_6t_5 inst_cell_20_100 (.BL(BL100),.BLN(BLN100),.WL(WL20));
sram_cell_6t_5 inst_cell_20_101 (.BL(BL101),.BLN(BLN101),.WL(WL20));
sram_cell_6t_5 inst_cell_20_102 (.BL(BL102),.BLN(BLN102),.WL(WL20));
sram_cell_6t_5 inst_cell_20_103 (.BL(BL103),.BLN(BLN103),.WL(WL20));
sram_cell_6t_5 inst_cell_20_104 (.BL(BL104),.BLN(BLN104),.WL(WL20));
sram_cell_6t_5 inst_cell_20_105 (.BL(BL105),.BLN(BLN105),.WL(WL20));
sram_cell_6t_5 inst_cell_20_106 (.BL(BL106),.BLN(BLN106),.WL(WL20));
sram_cell_6t_5 inst_cell_20_107 (.BL(BL107),.BLN(BLN107),.WL(WL20));
sram_cell_6t_5 inst_cell_20_108 (.BL(BL108),.BLN(BLN108),.WL(WL20));
sram_cell_6t_5 inst_cell_20_109 (.BL(BL109),.BLN(BLN109),.WL(WL20));
sram_cell_6t_5 inst_cell_20_110 (.BL(BL110),.BLN(BLN110),.WL(WL20));
sram_cell_6t_5 inst_cell_20_111 (.BL(BL111),.BLN(BLN111),.WL(WL20));
sram_cell_6t_5 inst_cell_20_112 (.BL(BL112),.BLN(BLN112),.WL(WL20));
sram_cell_6t_5 inst_cell_20_113 (.BL(BL113),.BLN(BLN113),.WL(WL20));
sram_cell_6t_5 inst_cell_20_114 (.BL(BL114),.BLN(BLN114),.WL(WL20));
sram_cell_6t_5 inst_cell_20_115 (.BL(BL115),.BLN(BLN115),.WL(WL20));
sram_cell_6t_5 inst_cell_20_116 (.BL(BL116),.BLN(BLN116),.WL(WL20));
sram_cell_6t_5 inst_cell_20_117 (.BL(BL117),.BLN(BLN117),.WL(WL20));
sram_cell_6t_5 inst_cell_20_118 (.BL(BL118),.BLN(BLN118),.WL(WL20));
sram_cell_6t_5 inst_cell_20_119 (.BL(BL119),.BLN(BLN119),.WL(WL20));
sram_cell_6t_5 inst_cell_20_120 (.BL(BL120),.BLN(BLN120),.WL(WL20));
sram_cell_6t_5 inst_cell_20_121 (.BL(BL121),.BLN(BLN121),.WL(WL20));
sram_cell_6t_5 inst_cell_20_122 (.BL(BL122),.BLN(BLN122),.WL(WL20));
sram_cell_6t_5 inst_cell_20_123 (.BL(BL123),.BLN(BLN123),.WL(WL20));
sram_cell_6t_5 inst_cell_20_124 (.BL(BL124),.BLN(BLN124),.WL(WL20));
sram_cell_6t_5 inst_cell_20_125 (.BL(BL125),.BLN(BLN125),.WL(WL20));
sram_cell_6t_5 inst_cell_20_126 (.BL(BL126),.BLN(BLN126),.WL(WL20));
sram_cell_6t_5 inst_cell_20_127 (.BL(BL127),.BLN(BLN127),.WL(WL20));
sram_cell_6t_5 inst_cell_21_0 (.BL(BL0),.BLN(BLN0),.WL(WL21));
sram_cell_6t_5 inst_cell_21_1 (.BL(BL1),.BLN(BLN1),.WL(WL21));
sram_cell_6t_5 inst_cell_21_2 (.BL(BL2),.BLN(BLN2),.WL(WL21));
sram_cell_6t_5 inst_cell_21_3 (.BL(BL3),.BLN(BLN3),.WL(WL21));
sram_cell_6t_5 inst_cell_21_4 (.BL(BL4),.BLN(BLN4),.WL(WL21));
sram_cell_6t_5 inst_cell_21_5 (.BL(BL5),.BLN(BLN5),.WL(WL21));
sram_cell_6t_5 inst_cell_21_6 (.BL(BL6),.BLN(BLN6),.WL(WL21));
sram_cell_6t_5 inst_cell_21_7 (.BL(BL7),.BLN(BLN7),.WL(WL21));
sram_cell_6t_5 inst_cell_21_8 (.BL(BL8),.BLN(BLN8),.WL(WL21));
sram_cell_6t_5 inst_cell_21_9 (.BL(BL9),.BLN(BLN9),.WL(WL21));
sram_cell_6t_5 inst_cell_21_10 (.BL(BL10),.BLN(BLN10),.WL(WL21));
sram_cell_6t_5 inst_cell_21_11 (.BL(BL11),.BLN(BLN11),.WL(WL21));
sram_cell_6t_5 inst_cell_21_12 (.BL(BL12),.BLN(BLN12),.WL(WL21));
sram_cell_6t_5 inst_cell_21_13 (.BL(BL13),.BLN(BLN13),.WL(WL21));
sram_cell_6t_5 inst_cell_21_14 (.BL(BL14),.BLN(BLN14),.WL(WL21));
sram_cell_6t_5 inst_cell_21_15 (.BL(BL15),.BLN(BLN15),.WL(WL21));
sram_cell_6t_5 inst_cell_21_16 (.BL(BL16),.BLN(BLN16),.WL(WL21));
sram_cell_6t_5 inst_cell_21_17 (.BL(BL17),.BLN(BLN17),.WL(WL21));
sram_cell_6t_5 inst_cell_21_18 (.BL(BL18),.BLN(BLN18),.WL(WL21));
sram_cell_6t_5 inst_cell_21_19 (.BL(BL19),.BLN(BLN19),.WL(WL21));
sram_cell_6t_5 inst_cell_21_20 (.BL(BL20),.BLN(BLN20),.WL(WL21));
sram_cell_6t_5 inst_cell_21_21 (.BL(BL21),.BLN(BLN21),.WL(WL21));
sram_cell_6t_5 inst_cell_21_22 (.BL(BL22),.BLN(BLN22),.WL(WL21));
sram_cell_6t_5 inst_cell_21_23 (.BL(BL23),.BLN(BLN23),.WL(WL21));
sram_cell_6t_5 inst_cell_21_24 (.BL(BL24),.BLN(BLN24),.WL(WL21));
sram_cell_6t_5 inst_cell_21_25 (.BL(BL25),.BLN(BLN25),.WL(WL21));
sram_cell_6t_5 inst_cell_21_26 (.BL(BL26),.BLN(BLN26),.WL(WL21));
sram_cell_6t_5 inst_cell_21_27 (.BL(BL27),.BLN(BLN27),.WL(WL21));
sram_cell_6t_5 inst_cell_21_28 (.BL(BL28),.BLN(BLN28),.WL(WL21));
sram_cell_6t_5 inst_cell_21_29 (.BL(BL29),.BLN(BLN29),.WL(WL21));
sram_cell_6t_5 inst_cell_21_30 (.BL(BL30),.BLN(BLN30),.WL(WL21));
sram_cell_6t_5 inst_cell_21_31 (.BL(BL31),.BLN(BLN31),.WL(WL21));
sram_cell_6t_5 inst_cell_21_32 (.BL(BL32),.BLN(BLN32),.WL(WL21));
sram_cell_6t_5 inst_cell_21_33 (.BL(BL33),.BLN(BLN33),.WL(WL21));
sram_cell_6t_5 inst_cell_21_34 (.BL(BL34),.BLN(BLN34),.WL(WL21));
sram_cell_6t_5 inst_cell_21_35 (.BL(BL35),.BLN(BLN35),.WL(WL21));
sram_cell_6t_5 inst_cell_21_36 (.BL(BL36),.BLN(BLN36),.WL(WL21));
sram_cell_6t_5 inst_cell_21_37 (.BL(BL37),.BLN(BLN37),.WL(WL21));
sram_cell_6t_5 inst_cell_21_38 (.BL(BL38),.BLN(BLN38),.WL(WL21));
sram_cell_6t_5 inst_cell_21_39 (.BL(BL39),.BLN(BLN39),.WL(WL21));
sram_cell_6t_5 inst_cell_21_40 (.BL(BL40),.BLN(BLN40),.WL(WL21));
sram_cell_6t_5 inst_cell_21_41 (.BL(BL41),.BLN(BLN41),.WL(WL21));
sram_cell_6t_5 inst_cell_21_42 (.BL(BL42),.BLN(BLN42),.WL(WL21));
sram_cell_6t_5 inst_cell_21_43 (.BL(BL43),.BLN(BLN43),.WL(WL21));
sram_cell_6t_5 inst_cell_21_44 (.BL(BL44),.BLN(BLN44),.WL(WL21));
sram_cell_6t_5 inst_cell_21_45 (.BL(BL45),.BLN(BLN45),.WL(WL21));
sram_cell_6t_5 inst_cell_21_46 (.BL(BL46),.BLN(BLN46),.WL(WL21));
sram_cell_6t_5 inst_cell_21_47 (.BL(BL47),.BLN(BLN47),.WL(WL21));
sram_cell_6t_5 inst_cell_21_48 (.BL(BL48),.BLN(BLN48),.WL(WL21));
sram_cell_6t_5 inst_cell_21_49 (.BL(BL49),.BLN(BLN49),.WL(WL21));
sram_cell_6t_5 inst_cell_21_50 (.BL(BL50),.BLN(BLN50),.WL(WL21));
sram_cell_6t_5 inst_cell_21_51 (.BL(BL51),.BLN(BLN51),.WL(WL21));
sram_cell_6t_5 inst_cell_21_52 (.BL(BL52),.BLN(BLN52),.WL(WL21));
sram_cell_6t_5 inst_cell_21_53 (.BL(BL53),.BLN(BLN53),.WL(WL21));
sram_cell_6t_5 inst_cell_21_54 (.BL(BL54),.BLN(BLN54),.WL(WL21));
sram_cell_6t_5 inst_cell_21_55 (.BL(BL55),.BLN(BLN55),.WL(WL21));
sram_cell_6t_5 inst_cell_21_56 (.BL(BL56),.BLN(BLN56),.WL(WL21));
sram_cell_6t_5 inst_cell_21_57 (.BL(BL57),.BLN(BLN57),.WL(WL21));
sram_cell_6t_5 inst_cell_21_58 (.BL(BL58),.BLN(BLN58),.WL(WL21));
sram_cell_6t_5 inst_cell_21_59 (.BL(BL59),.BLN(BLN59),.WL(WL21));
sram_cell_6t_5 inst_cell_21_60 (.BL(BL60),.BLN(BLN60),.WL(WL21));
sram_cell_6t_5 inst_cell_21_61 (.BL(BL61),.BLN(BLN61),.WL(WL21));
sram_cell_6t_5 inst_cell_21_62 (.BL(BL62),.BLN(BLN62),.WL(WL21));
sram_cell_6t_5 inst_cell_21_63 (.BL(BL63),.BLN(BLN63),.WL(WL21));
sram_cell_6t_5 inst_cell_21_64 (.BL(BL64),.BLN(BLN64),.WL(WL21));
sram_cell_6t_5 inst_cell_21_65 (.BL(BL65),.BLN(BLN65),.WL(WL21));
sram_cell_6t_5 inst_cell_21_66 (.BL(BL66),.BLN(BLN66),.WL(WL21));
sram_cell_6t_5 inst_cell_21_67 (.BL(BL67),.BLN(BLN67),.WL(WL21));
sram_cell_6t_5 inst_cell_21_68 (.BL(BL68),.BLN(BLN68),.WL(WL21));
sram_cell_6t_5 inst_cell_21_69 (.BL(BL69),.BLN(BLN69),.WL(WL21));
sram_cell_6t_5 inst_cell_21_70 (.BL(BL70),.BLN(BLN70),.WL(WL21));
sram_cell_6t_5 inst_cell_21_71 (.BL(BL71),.BLN(BLN71),.WL(WL21));
sram_cell_6t_5 inst_cell_21_72 (.BL(BL72),.BLN(BLN72),.WL(WL21));
sram_cell_6t_5 inst_cell_21_73 (.BL(BL73),.BLN(BLN73),.WL(WL21));
sram_cell_6t_5 inst_cell_21_74 (.BL(BL74),.BLN(BLN74),.WL(WL21));
sram_cell_6t_5 inst_cell_21_75 (.BL(BL75),.BLN(BLN75),.WL(WL21));
sram_cell_6t_5 inst_cell_21_76 (.BL(BL76),.BLN(BLN76),.WL(WL21));
sram_cell_6t_5 inst_cell_21_77 (.BL(BL77),.BLN(BLN77),.WL(WL21));
sram_cell_6t_5 inst_cell_21_78 (.BL(BL78),.BLN(BLN78),.WL(WL21));
sram_cell_6t_5 inst_cell_21_79 (.BL(BL79),.BLN(BLN79),.WL(WL21));
sram_cell_6t_5 inst_cell_21_80 (.BL(BL80),.BLN(BLN80),.WL(WL21));
sram_cell_6t_5 inst_cell_21_81 (.BL(BL81),.BLN(BLN81),.WL(WL21));
sram_cell_6t_5 inst_cell_21_82 (.BL(BL82),.BLN(BLN82),.WL(WL21));
sram_cell_6t_5 inst_cell_21_83 (.BL(BL83),.BLN(BLN83),.WL(WL21));
sram_cell_6t_5 inst_cell_21_84 (.BL(BL84),.BLN(BLN84),.WL(WL21));
sram_cell_6t_5 inst_cell_21_85 (.BL(BL85),.BLN(BLN85),.WL(WL21));
sram_cell_6t_5 inst_cell_21_86 (.BL(BL86),.BLN(BLN86),.WL(WL21));
sram_cell_6t_5 inst_cell_21_87 (.BL(BL87),.BLN(BLN87),.WL(WL21));
sram_cell_6t_5 inst_cell_21_88 (.BL(BL88),.BLN(BLN88),.WL(WL21));
sram_cell_6t_5 inst_cell_21_89 (.BL(BL89),.BLN(BLN89),.WL(WL21));
sram_cell_6t_5 inst_cell_21_90 (.BL(BL90),.BLN(BLN90),.WL(WL21));
sram_cell_6t_5 inst_cell_21_91 (.BL(BL91),.BLN(BLN91),.WL(WL21));
sram_cell_6t_5 inst_cell_21_92 (.BL(BL92),.BLN(BLN92),.WL(WL21));
sram_cell_6t_5 inst_cell_21_93 (.BL(BL93),.BLN(BLN93),.WL(WL21));
sram_cell_6t_5 inst_cell_21_94 (.BL(BL94),.BLN(BLN94),.WL(WL21));
sram_cell_6t_5 inst_cell_21_95 (.BL(BL95),.BLN(BLN95),.WL(WL21));
sram_cell_6t_5 inst_cell_21_96 (.BL(BL96),.BLN(BLN96),.WL(WL21));
sram_cell_6t_5 inst_cell_21_97 (.BL(BL97),.BLN(BLN97),.WL(WL21));
sram_cell_6t_5 inst_cell_21_98 (.BL(BL98),.BLN(BLN98),.WL(WL21));
sram_cell_6t_5 inst_cell_21_99 (.BL(BL99),.BLN(BLN99),.WL(WL21));
sram_cell_6t_5 inst_cell_21_100 (.BL(BL100),.BLN(BLN100),.WL(WL21));
sram_cell_6t_5 inst_cell_21_101 (.BL(BL101),.BLN(BLN101),.WL(WL21));
sram_cell_6t_5 inst_cell_21_102 (.BL(BL102),.BLN(BLN102),.WL(WL21));
sram_cell_6t_5 inst_cell_21_103 (.BL(BL103),.BLN(BLN103),.WL(WL21));
sram_cell_6t_5 inst_cell_21_104 (.BL(BL104),.BLN(BLN104),.WL(WL21));
sram_cell_6t_5 inst_cell_21_105 (.BL(BL105),.BLN(BLN105),.WL(WL21));
sram_cell_6t_5 inst_cell_21_106 (.BL(BL106),.BLN(BLN106),.WL(WL21));
sram_cell_6t_5 inst_cell_21_107 (.BL(BL107),.BLN(BLN107),.WL(WL21));
sram_cell_6t_5 inst_cell_21_108 (.BL(BL108),.BLN(BLN108),.WL(WL21));
sram_cell_6t_5 inst_cell_21_109 (.BL(BL109),.BLN(BLN109),.WL(WL21));
sram_cell_6t_5 inst_cell_21_110 (.BL(BL110),.BLN(BLN110),.WL(WL21));
sram_cell_6t_5 inst_cell_21_111 (.BL(BL111),.BLN(BLN111),.WL(WL21));
sram_cell_6t_5 inst_cell_21_112 (.BL(BL112),.BLN(BLN112),.WL(WL21));
sram_cell_6t_5 inst_cell_21_113 (.BL(BL113),.BLN(BLN113),.WL(WL21));
sram_cell_6t_5 inst_cell_21_114 (.BL(BL114),.BLN(BLN114),.WL(WL21));
sram_cell_6t_5 inst_cell_21_115 (.BL(BL115),.BLN(BLN115),.WL(WL21));
sram_cell_6t_5 inst_cell_21_116 (.BL(BL116),.BLN(BLN116),.WL(WL21));
sram_cell_6t_5 inst_cell_21_117 (.BL(BL117),.BLN(BLN117),.WL(WL21));
sram_cell_6t_5 inst_cell_21_118 (.BL(BL118),.BLN(BLN118),.WL(WL21));
sram_cell_6t_5 inst_cell_21_119 (.BL(BL119),.BLN(BLN119),.WL(WL21));
sram_cell_6t_5 inst_cell_21_120 (.BL(BL120),.BLN(BLN120),.WL(WL21));
sram_cell_6t_5 inst_cell_21_121 (.BL(BL121),.BLN(BLN121),.WL(WL21));
sram_cell_6t_5 inst_cell_21_122 (.BL(BL122),.BLN(BLN122),.WL(WL21));
sram_cell_6t_5 inst_cell_21_123 (.BL(BL123),.BLN(BLN123),.WL(WL21));
sram_cell_6t_5 inst_cell_21_124 (.BL(BL124),.BLN(BLN124),.WL(WL21));
sram_cell_6t_5 inst_cell_21_125 (.BL(BL125),.BLN(BLN125),.WL(WL21));
sram_cell_6t_5 inst_cell_21_126 (.BL(BL126),.BLN(BLN126),.WL(WL21));
sram_cell_6t_5 inst_cell_21_127 (.BL(BL127),.BLN(BLN127),.WL(WL21));
sram_cell_6t_5 inst_cell_22_0 (.BL(BL0),.BLN(BLN0),.WL(WL22));
sram_cell_6t_5 inst_cell_22_1 (.BL(BL1),.BLN(BLN1),.WL(WL22));
sram_cell_6t_5 inst_cell_22_2 (.BL(BL2),.BLN(BLN2),.WL(WL22));
sram_cell_6t_5 inst_cell_22_3 (.BL(BL3),.BLN(BLN3),.WL(WL22));
sram_cell_6t_5 inst_cell_22_4 (.BL(BL4),.BLN(BLN4),.WL(WL22));
sram_cell_6t_5 inst_cell_22_5 (.BL(BL5),.BLN(BLN5),.WL(WL22));
sram_cell_6t_5 inst_cell_22_6 (.BL(BL6),.BLN(BLN6),.WL(WL22));
sram_cell_6t_5 inst_cell_22_7 (.BL(BL7),.BLN(BLN7),.WL(WL22));
sram_cell_6t_5 inst_cell_22_8 (.BL(BL8),.BLN(BLN8),.WL(WL22));
sram_cell_6t_5 inst_cell_22_9 (.BL(BL9),.BLN(BLN9),.WL(WL22));
sram_cell_6t_5 inst_cell_22_10 (.BL(BL10),.BLN(BLN10),.WL(WL22));
sram_cell_6t_5 inst_cell_22_11 (.BL(BL11),.BLN(BLN11),.WL(WL22));
sram_cell_6t_5 inst_cell_22_12 (.BL(BL12),.BLN(BLN12),.WL(WL22));
sram_cell_6t_5 inst_cell_22_13 (.BL(BL13),.BLN(BLN13),.WL(WL22));
sram_cell_6t_5 inst_cell_22_14 (.BL(BL14),.BLN(BLN14),.WL(WL22));
sram_cell_6t_5 inst_cell_22_15 (.BL(BL15),.BLN(BLN15),.WL(WL22));
sram_cell_6t_5 inst_cell_22_16 (.BL(BL16),.BLN(BLN16),.WL(WL22));
sram_cell_6t_5 inst_cell_22_17 (.BL(BL17),.BLN(BLN17),.WL(WL22));
sram_cell_6t_5 inst_cell_22_18 (.BL(BL18),.BLN(BLN18),.WL(WL22));
sram_cell_6t_5 inst_cell_22_19 (.BL(BL19),.BLN(BLN19),.WL(WL22));
sram_cell_6t_5 inst_cell_22_20 (.BL(BL20),.BLN(BLN20),.WL(WL22));
sram_cell_6t_5 inst_cell_22_21 (.BL(BL21),.BLN(BLN21),.WL(WL22));
sram_cell_6t_5 inst_cell_22_22 (.BL(BL22),.BLN(BLN22),.WL(WL22));
sram_cell_6t_5 inst_cell_22_23 (.BL(BL23),.BLN(BLN23),.WL(WL22));
sram_cell_6t_5 inst_cell_22_24 (.BL(BL24),.BLN(BLN24),.WL(WL22));
sram_cell_6t_5 inst_cell_22_25 (.BL(BL25),.BLN(BLN25),.WL(WL22));
sram_cell_6t_5 inst_cell_22_26 (.BL(BL26),.BLN(BLN26),.WL(WL22));
sram_cell_6t_5 inst_cell_22_27 (.BL(BL27),.BLN(BLN27),.WL(WL22));
sram_cell_6t_5 inst_cell_22_28 (.BL(BL28),.BLN(BLN28),.WL(WL22));
sram_cell_6t_5 inst_cell_22_29 (.BL(BL29),.BLN(BLN29),.WL(WL22));
sram_cell_6t_5 inst_cell_22_30 (.BL(BL30),.BLN(BLN30),.WL(WL22));
sram_cell_6t_5 inst_cell_22_31 (.BL(BL31),.BLN(BLN31),.WL(WL22));
sram_cell_6t_5 inst_cell_22_32 (.BL(BL32),.BLN(BLN32),.WL(WL22));
sram_cell_6t_5 inst_cell_22_33 (.BL(BL33),.BLN(BLN33),.WL(WL22));
sram_cell_6t_5 inst_cell_22_34 (.BL(BL34),.BLN(BLN34),.WL(WL22));
sram_cell_6t_5 inst_cell_22_35 (.BL(BL35),.BLN(BLN35),.WL(WL22));
sram_cell_6t_5 inst_cell_22_36 (.BL(BL36),.BLN(BLN36),.WL(WL22));
sram_cell_6t_5 inst_cell_22_37 (.BL(BL37),.BLN(BLN37),.WL(WL22));
sram_cell_6t_5 inst_cell_22_38 (.BL(BL38),.BLN(BLN38),.WL(WL22));
sram_cell_6t_5 inst_cell_22_39 (.BL(BL39),.BLN(BLN39),.WL(WL22));
sram_cell_6t_5 inst_cell_22_40 (.BL(BL40),.BLN(BLN40),.WL(WL22));
sram_cell_6t_5 inst_cell_22_41 (.BL(BL41),.BLN(BLN41),.WL(WL22));
sram_cell_6t_5 inst_cell_22_42 (.BL(BL42),.BLN(BLN42),.WL(WL22));
sram_cell_6t_5 inst_cell_22_43 (.BL(BL43),.BLN(BLN43),.WL(WL22));
sram_cell_6t_5 inst_cell_22_44 (.BL(BL44),.BLN(BLN44),.WL(WL22));
sram_cell_6t_5 inst_cell_22_45 (.BL(BL45),.BLN(BLN45),.WL(WL22));
sram_cell_6t_5 inst_cell_22_46 (.BL(BL46),.BLN(BLN46),.WL(WL22));
sram_cell_6t_5 inst_cell_22_47 (.BL(BL47),.BLN(BLN47),.WL(WL22));
sram_cell_6t_5 inst_cell_22_48 (.BL(BL48),.BLN(BLN48),.WL(WL22));
sram_cell_6t_5 inst_cell_22_49 (.BL(BL49),.BLN(BLN49),.WL(WL22));
sram_cell_6t_5 inst_cell_22_50 (.BL(BL50),.BLN(BLN50),.WL(WL22));
sram_cell_6t_5 inst_cell_22_51 (.BL(BL51),.BLN(BLN51),.WL(WL22));
sram_cell_6t_5 inst_cell_22_52 (.BL(BL52),.BLN(BLN52),.WL(WL22));
sram_cell_6t_5 inst_cell_22_53 (.BL(BL53),.BLN(BLN53),.WL(WL22));
sram_cell_6t_5 inst_cell_22_54 (.BL(BL54),.BLN(BLN54),.WL(WL22));
sram_cell_6t_5 inst_cell_22_55 (.BL(BL55),.BLN(BLN55),.WL(WL22));
sram_cell_6t_5 inst_cell_22_56 (.BL(BL56),.BLN(BLN56),.WL(WL22));
sram_cell_6t_5 inst_cell_22_57 (.BL(BL57),.BLN(BLN57),.WL(WL22));
sram_cell_6t_5 inst_cell_22_58 (.BL(BL58),.BLN(BLN58),.WL(WL22));
sram_cell_6t_5 inst_cell_22_59 (.BL(BL59),.BLN(BLN59),.WL(WL22));
sram_cell_6t_5 inst_cell_22_60 (.BL(BL60),.BLN(BLN60),.WL(WL22));
sram_cell_6t_5 inst_cell_22_61 (.BL(BL61),.BLN(BLN61),.WL(WL22));
sram_cell_6t_5 inst_cell_22_62 (.BL(BL62),.BLN(BLN62),.WL(WL22));
sram_cell_6t_5 inst_cell_22_63 (.BL(BL63),.BLN(BLN63),.WL(WL22));
sram_cell_6t_5 inst_cell_22_64 (.BL(BL64),.BLN(BLN64),.WL(WL22));
sram_cell_6t_5 inst_cell_22_65 (.BL(BL65),.BLN(BLN65),.WL(WL22));
sram_cell_6t_5 inst_cell_22_66 (.BL(BL66),.BLN(BLN66),.WL(WL22));
sram_cell_6t_5 inst_cell_22_67 (.BL(BL67),.BLN(BLN67),.WL(WL22));
sram_cell_6t_5 inst_cell_22_68 (.BL(BL68),.BLN(BLN68),.WL(WL22));
sram_cell_6t_5 inst_cell_22_69 (.BL(BL69),.BLN(BLN69),.WL(WL22));
sram_cell_6t_5 inst_cell_22_70 (.BL(BL70),.BLN(BLN70),.WL(WL22));
sram_cell_6t_5 inst_cell_22_71 (.BL(BL71),.BLN(BLN71),.WL(WL22));
sram_cell_6t_5 inst_cell_22_72 (.BL(BL72),.BLN(BLN72),.WL(WL22));
sram_cell_6t_5 inst_cell_22_73 (.BL(BL73),.BLN(BLN73),.WL(WL22));
sram_cell_6t_5 inst_cell_22_74 (.BL(BL74),.BLN(BLN74),.WL(WL22));
sram_cell_6t_5 inst_cell_22_75 (.BL(BL75),.BLN(BLN75),.WL(WL22));
sram_cell_6t_5 inst_cell_22_76 (.BL(BL76),.BLN(BLN76),.WL(WL22));
sram_cell_6t_5 inst_cell_22_77 (.BL(BL77),.BLN(BLN77),.WL(WL22));
sram_cell_6t_5 inst_cell_22_78 (.BL(BL78),.BLN(BLN78),.WL(WL22));
sram_cell_6t_5 inst_cell_22_79 (.BL(BL79),.BLN(BLN79),.WL(WL22));
sram_cell_6t_5 inst_cell_22_80 (.BL(BL80),.BLN(BLN80),.WL(WL22));
sram_cell_6t_5 inst_cell_22_81 (.BL(BL81),.BLN(BLN81),.WL(WL22));
sram_cell_6t_5 inst_cell_22_82 (.BL(BL82),.BLN(BLN82),.WL(WL22));
sram_cell_6t_5 inst_cell_22_83 (.BL(BL83),.BLN(BLN83),.WL(WL22));
sram_cell_6t_5 inst_cell_22_84 (.BL(BL84),.BLN(BLN84),.WL(WL22));
sram_cell_6t_5 inst_cell_22_85 (.BL(BL85),.BLN(BLN85),.WL(WL22));
sram_cell_6t_5 inst_cell_22_86 (.BL(BL86),.BLN(BLN86),.WL(WL22));
sram_cell_6t_5 inst_cell_22_87 (.BL(BL87),.BLN(BLN87),.WL(WL22));
sram_cell_6t_5 inst_cell_22_88 (.BL(BL88),.BLN(BLN88),.WL(WL22));
sram_cell_6t_5 inst_cell_22_89 (.BL(BL89),.BLN(BLN89),.WL(WL22));
sram_cell_6t_5 inst_cell_22_90 (.BL(BL90),.BLN(BLN90),.WL(WL22));
sram_cell_6t_5 inst_cell_22_91 (.BL(BL91),.BLN(BLN91),.WL(WL22));
sram_cell_6t_5 inst_cell_22_92 (.BL(BL92),.BLN(BLN92),.WL(WL22));
sram_cell_6t_5 inst_cell_22_93 (.BL(BL93),.BLN(BLN93),.WL(WL22));
sram_cell_6t_5 inst_cell_22_94 (.BL(BL94),.BLN(BLN94),.WL(WL22));
sram_cell_6t_5 inst_cell_22_95 (.BL(BL95),.BLN(BLN95),.WL(WL22));
sram_cell_6t_5 inst_cell_22_96 (.BL(BL96),.BLN(BLN96),.WL(WL22));
sram_cell_6t_5 inst_cell_22_97 (.BL(BL97),.BLN(BLN97),.WL(WL22));
sram_cell_6t_5 inst_cell_22_98 (.BL(BL98),.BLN(BLN98),.WL(WL22));
sram_cell_6t_5 inst_cell_22_99 (.BL(BL99),.BLN(BLN99),.WL(WL22));
sram_cell_6t_5 inst_cell_22_100 (.BL(BL100),.BLN(BLN100),.WL(WL22));
sram_cell_6t_5 inst_cell_22_101 (.BL(BL101),.BLN(BLN101),.WL(WL22));
sram_cell_6t_5 inst_cell_22_102 (.BL(BL102),.BLN(BLN102),.WL(WL22));
sram_cell_6t_5 inst_cell_22_103 (.BL(BL103),.BLN(BLN103),.WL(WL22));
sram_cell_6t_5 inst_cell_22_104 (.BL(BL104),.BLN(BLN104),.WL(WL22));
sram_cell_6t_5 inst_cell_22_105 (.BL(BL105),.BLN(BLN105),.WL(WL22));
sram_cell_6t_5 inst_cell_22_106 (.BL(BL106),.BLN(BLN106),.WL(WL22));
sram_cell_6t_5 inst_cell_22_107 (.BL(BL107),.BLN(BLN107),.WL(WL22));
sram_cell_6t_5 inst_cell_22_108 (.BL(BL108),.BLN(BLN108),.WL(WL22));
sram_cell_6t_5 inst_cell_22_109 (.BL(BL109),.BLN(BLN109),.WL(WL22));
sram_cell_6t_5 inst_cell_22_110 (.BL(BL110),.BLN(BLN110),.WL(WL22));
sram_cell_6t_5 inst_cell_22_111 (.BL(BL111),.BLN(BLN111),.WL(WL22));
sram_cell_6t_5 inst_cell_22_112 (.BL(BL112),.BLN(BLN112),.WL(WL22));
sram_cell_6t_5 inst_cell_22_113 (.BL(BL113),.BLN(BLN113),.WL(WL22));
sram_cell_6t_5 inst_cell_22_114 (.BL(BL114),.BLN(BLN114),.WL(WL22));
sram_cell_6t_5 inst_cell_22_115 (.BL(BL115),.BLN(BLN115),.WL(WL22));
sram_cell_6t_5 inst_cell_22_116 (.BL(BL116),.BLN(BLN116),.WL(WL22));
sram_cell_6t_5 inst_cell_22_117 (.BL(BL117),.BLN(BLN117),.WL(WL22));
sram_cell_6t_5 inst_cell_22_118 (.BL(BL118),.BLN(BLN118),.WL(WL22));
sram_cell_6t_5 inst_cell_22_119 (.BL(BL119),.BLN(BLN119),.WL(WL22));
sram_cell_6t_5 inst_cell_22_120 (.BL(BL120),.BLN(BLN120),.WL(WL22));
sram_cell_6t_5 inst_cell_22_121 (.BL(BL121),.BLN(BLN121),.WL(WL22));
sram_cell_6t_5 inst_cell_22_122 (.BL(BL122),.BLN(BLN122),.WL(WL22));
sram_cell_6t_5 inst_cell_22_123 (.BL(BL123),.BLN(BLN123),.WL(WL22));
sram_cell_6t_5 inst_cell_22_124 (.BL(BL124),.BLN(BLN124),.WL(WL22));
sram_cell_6t_5 inst_cell_22_125 (.BL(BL125),.BLN(BLN125),.WL(WL22));
sram_cell_6t_5 inst_cell_22_126 (.BL(BL126),.BLN(BLN126),.WL(WL22));
sram_cell_6t_5 inst_cell_22_127 (.BL(BL127),.BLN(BLN127),.WL(WL22));
sram_cell_6t_5 inst_cell_23_0 (.BL(BL0),.BLN(BLN0),.WL(WL23));
sram_cell_6t_5 inst_cell_23_1 (.BL(BL1),.BLN(BLN1),.WL(WL23));
sram_cell_6t_5 inst_cell_23_2 (.BL(BL2),.BLN(BLN2),.WL(WL23));
sram_cell_6t_5 inst_cell_23_3 (.BL(BL3),.BLN(BLN3),.WL(WL23));
sram_cell_6t_5 inst_cell_23_4 (.BL(BL4),.BLN(BLN4),.WL(WL23));
sram_cell_6t_5 inst_cell_23_5 (.BL(BL5),.BLN(BLN5),.WL(WL23));
sram_cell_6t_5 inst_cell_23_6 (.BL(BL6),.BLN(BLN6),.WL(WL23));
sram_cell_6t_5 inst_cell_23_7 (.BL(BL7),.BLN(BLN7),.WL(WL23));
sram_cell_6t_5 inst_cell_23_8 (.BL(BL8),.BLN(BLN8),.WL(WL23));
sram_cell_6t_5 inst_cell_23_9 (.BL(BL9),.BLN(BLN9),.WL(WL23));
sram_cell_6t_5 inst_cell_23_10 (.BL(BL10),.BLN(BLN10),.WL(WL23));
sram_cell_6t_5 inst_cell_23_11 (.BL(BL11),.BLN(BLN11),.WL(WL23));
sram_cell_6t_5 inst_cell_23_12 (.BL(BL12),.BLN(BLN12),.WL(WL23));
sram_cell_6t_5 inst_cell_23_13 (.BL(BL13),.BLN(BLN13),.WL(WL23));
sram_cell_6t_5 inst_cell_23_14 (.BL(BL14),.BLN(BLN14),.WL(WL23));
sram_cell_6t_5 inst_cell_23_15 (.BL(BL15),.BLN(BLN15),.WL(WL23));
sram_cell_6t_5 inst_cell_23_16 (.BL(BL16),.BLN(BLN16),.WL(WL23));
sram_cell_6t_5 inst_cell_23_17 (.BL(BL17),.BLN(BLN17),.WL(WL23));
sram_cell_6t_5 inst_cell_23_18 (.BL(BL18),.BLN(BLN18),.WL(WL23));
sram_cell_6t_5 inst_cell_23_19 (.BL(BL19),.BLN(BLN19),.WL(WL23));
sram_cell_6t_5 inst_cell_23_20 (.BL(BL20),.BLN(BLN20),.WL(WL23));
sram_cell_6t_5 inst_cell_23_21 (.BL(BL21),.BLN(BLN21),.WL(WL23));
sram_cell_6t_5 inst_cell_23_22 (.BL(BL22),.BLN(BLN22),.WL(WL23));
sram_cell_6t_5 inst_cell_23_23 (.BL(BL23),.BLN(BLN23),.WL(WL23));
sram_cell_6t_5 inst_cell_23_24 (.BL(BL24),.BLN(BLN24),.WL(WL23));
sram_cell_6t_5 inst_cell_23_25 (.BL(BL25),.BLN(BLN25),.WL(WL23));
sram_cell_6t_5 inst_cell_23_26 (.BL(BL26),.BLN(BLN26),.WL(WL23));
sram_cell_6t_5 inst_cell_23_27 (.BL(BL27),.BLN(BLN27),.WL(WL23));
sram_cell_6t_5 inst_cell_23_28 (.BL(BL28),.BLN(BLN28),.WL(WL23));
sram_cell_6t_5 inst_cell_23_29 (.BL(BL29),.BLN(BLN29),.WL(WL23));
sram_cell_6t_5 inst_cell_23_30 (.BL(BL30),.BLN(BLN30),.WL(WL23));
sram_cell_6t_5 inst_cell_23_31 (.BL(BL31),.BLN(BLN31),.WL(WL23));
sram_cell_6t_5 inst_cell_23_32 (.BL(BL32),.BLN(BLN32),.WL(WL23));
sram_cell_6t_5 inst_cell_23_33 (.BL(BL33),.BLN(BLN33),.WL(WL23));
sram_cell_6t_5 inst_cell_23_34 (.BL(BL34),.BLN(BLN34),.WL(WL23));
sram_cell_6t_5 inst_cell_23_35 (.BL(BL35),.BLN(BLN35),.WL(WL23));
sram_cell_6t_5 inst_cell_23_36 (.BL(BL36),.BLN(BLN36),.WL(WL23));
sram_cell_6t_5 inst_cell_23_37 (.BL(BL37),.BLN(BLN37),.WL(WL23));
sram_cell_6t_5 inst_cell_23_38 (.BL(BL38),.BLN(BLN38),.WL(WL23));
sram_cell_6t_5 inst_cell_23_39 (.BL(BL39),.BLN(BLN39),.WL(WL23));
sram_cell_6t_5 inst_cell_23_40 (.BL(BL40),.BLN(BLN40),.WL(WL23));
sram_cell_6t_5 inst_cell_23_41 (.BL(BL41),.BLN(BLN41),.WL(WL23));
sram_cell_6t_5 inst_cell_23_42 (.BL(BL42),.BLN(BLN42),.WL(WL23));
sram_cell_6t_5 inst_cell_23_43 (.BL(BL43),.BLN(BLN43),.WL(WL23));
sram_cell_6t_5 inst_cell_23_44 (.BL(BL44),.BLN(BLN44),.WL(WL23));
sram_cell_6t_5 inst_cell_23_45 (.BL(BL45),.BLN(BLN45),.WL(WL23));
sram_cell_6t_5 inst_cell_23_46 (.BL(BL46),.BLN(BLN46),.WL(WL23));
sram_cell_6t_5 inst_cell_23_47 (.BL(BL47),.BLN(BLN47),.WL(WL23));
sram_cell_6t_5 inst_cell_23_48 (.BL(BL48),.BLN(BLN48),.WL(WL23));
sram_cell_6t_5 inst_cell_23_49 (.BL(BL49),.BLN(BLN49),.WL(WL23));
sram_cell_6t_5 inst_cell_23_50 (.BL(BL50),.BLN(BLN50),.WL(WL23));
sram_cell_6t_5 inst_cell_23_51 (.BL(BL51),.BLN(BLN51),.WL(WL23));
sram_cell_6t_5 inst_cell_23_52 (.BL(BL52),.BLN(BLN52),.WL(WL23));
sram_cell_6t_5 inst_cell_23_53 (.BL(BL53),.BLN(BLN53),.WL(WL23));
sram_cell_6t_5 inst_cell_23_54 (.BL(BL54),.BLN(BLN54),.WL(WL23));
sram_cell_6t_5 inst_cell_23_55 (.BL(BL55),.BLN(BLN55),.WL(WL23));
sram_cell_6t_5 inst_cell_23_56 (.BL(BL56),.BLN(BLN56),.WL(WL23));
sram_cell_6t_5 inst_cell_23_57 (.BL(BL57),.BLN(BLN57),.WL(WL23));
sram_cell_6t_5 inst_cell_23_58 (.BL(BL58),.BLN(BLN58),.WL(WL23));
sram_cell_6t_5 inst_cell_23_59 (.BL(BL59),.BLN(BLN59),.WL(WL23));
sram_cell_6t_5 inst_cell_23_60 (.BL(BL60),.BLN(BLN60),.WL(WL23));
sram_cell_6t_5 inst_cell_23_61 (.BL(BL61),.BLN(BLN61),.WL(WL23));
sram_cell_6t_5 inst_cell_23_62 (.BL(BL62),.BLN(BLN62),.WL(WL23));
sram_cell_6t_5 inst_cell_23_63 (.BL(BL63),.BLN(BLN63),.WL(WL23));
sram_cell_6t_5 inst_cell_23_64 (.BL(BL64),.BLN(BLN64),.WL(WL23));
sram_cell_6t_5 inst_cell_23_65 (.BL(BL65),.BLN(BLN65),.WL(WL23));
sram_cell_6t_5 inst_cell_23_66 (.BL(BL66),.BLN(BLN66),.WL(WL23));
sram_cell_6t_5 inst_cell_23_67 (.BL(BL67),.BLN(BLN67),.WL(WL23));
sram_cell_6t_5 inst_cell_23_68 (.BL(BL68),.BLN(BLN68),.WL(WL23));
sram_cell_6t_5 inst_cell_23_69 (.BL(BL69),.BLN(BLN69),.WL(WL23));
sram_cell_6t_5 inst_cell_23_70 (.BL(BL70),.BLN(BLN70),.WL(WL23));
sram_cell_6t_5 inst_cell_23_71 (.BL(BL71),.BLN(BLN71),.WL(WL23));
sram_cell_6t_5 inst_cell_23_72 (.BL(BL72),.BLN(BLN72),.WL(WL23));
sram_cell_6t_5 inst_cell_23_73 (.BL(BL73),.BLN(BLN73),.WL(WL23));
sram_cell_6t_5 inst_cell_23_74 (.BL(BL74),.BLN(BLN74),.WL(WL23));
sram_cell_6t_5 inst_cell_23_75 (.BL(BL75),.BLN(BLN75),.WL(WL23));
sram_cell_6t_5 inst_cell_23_76 (.BL(BL76),.BLN(BLN76),.WL(WL23));
sram_cell_6t_5 inst_cell_23_77 (.BL(BL77),.BLN(BLN77),.WL(WL23));
sram_cell_6t_5 inst_cell_23_78 (.BL(BL78),.BLN(BLN78),.WL(WL23));
sram_cell_6t_5 inst_cell_23_79 (.BL(BL79),.BLN(BLN79),.WL(WL23));
sram_cell_6t_5 inst_cell_23_80 (.BL(BL80),.BLN(BLN80),.WL(WL23));
sram_cell_6t_5 inst_cell_23_81 (.BL(BL81),.BLN(BLN81),.WL(WL23));
sram_cell_6t_5 inst_cell_23_82 (.BL(BL82),.BLN(BLN82),.WL(WL23));
sram_cell_6t_5 inst_cell_23_83 (.BL(BL83),.BLN(BLN83),.WL(WL23));
sram_cell_6t_5 inst_cell_23_84 (.BL(BL84),.BLN(BLN84),.WL(WL23));
sram_cell_6t_5 inst_cell_23_85 (.BL(BL85),.BLN(BLN85),.WL(WL23));
sram_cell_6t_5 inst_cell_23_86 (.BL(BL86),.BLN(BLN86),.WL(WL23));
sram_cell_6t_5 inst_cell_23_87 (.BL(BL87),.BLN(BLN87),.WL(WL23));
sram_cell_6t_5 inst_cell_23_88 (.BL(BL88),.BLN(BLN88),.WL(WL23));
sram_cell_6t_5 inst_cell_23_89 (.BL(BL89),.BLN(BLN89),.WL(WL23));
sram_cell_6t_5 inst_cell_23_90 (.BL(BL90),.BLN(BLN90),.WL(WL23));
sram_cell_6t_5 inst_cell_23_91 (.BL(BL91),.BLN(BLN91),.WL(WL23));
sram_cell_6t_5 inst_cell_23_92 (.BL(BL92),.BLN(BLN92),.WL(WL23));
sram_cell_6t_5 inst_cell_23_93 (.BL(BL93),.BLN(BLN93),.WL(WL23));
sram_cell_6t_5 inst_cell_23_94 (.BL(BL94),.BLN(BLN94),.WL(WL23));
sram_cell_6t_5 inst_cell_23_95 (.BL(BL95),.BLN(BLN95),.WL(WL23));
sram_cell_6t_5 inst_cell_23_96 (.BL(BL96),.BLN(BLN96),.WL(WL23));
sram_cell_6t_5 inst_cell_23_97 (.BL(BL97),.BLN(BLN97),.WL(WL23));
sram_cell_6t_5 inst_cell_23_98 (.BL(BL98),.BLN(BLN98),.WL(WL23));
sram_cell_6t_5 inst_cell_23_99 (.BL(BL99),.BLN(BLN99),.WL(WL23));
sram_cell_6t_5 inst_cell_23_100 (.BL(BL100),.BLN(BLN100),.WL(WL23));
sram_cell_6t_5 inst_cell_23_101 (.BL(BL101),.BLN(BLN101),.WL(WL23));
sram_cell_6t_5 inst_cell_23_102 (.BL(BL102),.BLN(BLN102),.WL(WL23));
sram_cell_6t_5 inst_cell_23_103 (.BL(BL103),.BLN(BLN103),.WL(WL23));
sram_cell_6t_5 inst_cell_23_104 (.BL(BL104),.BLN(BLN104),.WL(WL23));
sram_cell_6t_5 inst_cell_23_105 (.BL(BL105),.BLN(BLN105),.WL(WL23));
sram_cell_6t_5 inst_cell_23_106 (.BL(BL106),.BLN(BLN106),.WL(WL23));
sram_cell_6t_5 inst_cell_23_107 (.BL(BL107),.BLN(BLN107),.WL(WL23));
sram_cell_6t_5 inst_cell_23_108 (.BL(BL108),.BLN(BLN108),.WL(WL23));
sram_cell_6t_5 inst_cell_23_109 (.BL(BL109),.BLN(BLN109),.WL(WL23));
sram_cell_6t_5 inst_cell_23_110 (.BL(BL110),.BLN(BLN110),.WL(WL23));
sram_cell_6t_5 inst_cell_23_111 (.BL(BL111),.BLN(BLN111),.WL(WL23));
sram_cell_6t_5 inst_cell_23_112 (.BL(BL112),.BLN(BLN112),.WL(WL23));
sram_cell_6t_5 inst_cell_23_113 (.BL(BL113),.BLN(BLN113),.WL(WL23));
sram_cell_6t_5 inst_cell_23_114 (.BL(BL114),.BLN(BLN114),.WL(WL23));
sram_cell_6t_5 inst_cell_23_115 (.BL(BL115),.BLN(BLN115),.WL(WL23));
sram_cell_6t_5 inst_cell_23_116 (.BL(BL116),.BLN(BLN116),.WL(WL23));
sram_cell_6t_5 inst_cell_23_117 (.BL(BL117),.BLN(BLN117),.WL(WL23));
sram_cell_6t_5 inst_cell_23_118 (.BL(BL118),.BLN(BLN118),.WL(WL23));
sram_cell_6t_5 inst_cell_23_119 (.BL(BL119),.BLN(BLN119),.WL(WL23));
sram_cell_6t_5 inst_cell_23_120 (.BL(BL120),.BLN(BLN120),.WL(WL23));
sram_cell_6t_5 inst_cell_23_121 (.BL(BL121),.BLN(BLN121),.WL(WL23));
sram_cell_6t_5 inst_cell_23_122 (.BL(BL122),.BLN(BLN122),.WL(WL23));
sram_cell_6t_5 inst_cell_23_123 (.BL(BL123),.BLN(BLN123),.WL(WL23));
sram_cell_6t_5 inst_cell_23_124 (.BL(BL124),.BLN(BLN124),.WL(WL23));
sram_cell_6t_5 inst_cell_23_125 (.BL(BL125),.BLN(BLN125),.WL(WL23));
sram_cell_6t_5 inst_cell_23_126 (.BL(BL126),.BLN(BLN126),.WL(WL23));
sram_cell_6t_5 inst_cell_23_127 (.BL(BL127),.BLN(BLN127),.WL(WL23));
sram_cell_6t_5 inst_cell_24_0 (.BL(BL0),.BLN(BLN0),.WL(WL24));
sram_cell_6t_5 inst_cell_24_1 (.BL(BL1),.BLN(BLN1),.WL(WL24));
sram_cell_6t_5 inst_cell_24_2 (.BL(BL2),.BLN(BLN2),.WL(WL24));
sram_cell_6t_5 inst_cell_24_3 (.BL(BL3),.BLN(BLN3),.WL(WL24));
sram_cell_6t_5 inst_cell_24_4 (.BL(BL4),.BLN(BLN4),.WL(WL24));
sram_cell_6t_5 inst_cell_24_5 (.BL(BL5),.BLN(BLN5),.WL(WL24));
sram_cell_6t_5 inst_cell_24_6 (.BL(BL6),.BLN(BLN6),.WL(WL24));
sram_cell_6t_5 inst_cell_24_7 (.BL(BL7),.BLN(BLN7),.WL(WL24));
sram_cell_6t_5 inst_cell_24_8 (.BL(BL8),.BLN(BLN8),.WL(WL24));
sram_cell_6t_5 inst_cell_24_9 (.BL(BL9),.BLN(BLN9),.WL(WL24));
sram_cell_6t_5 inst_cell_24_10 (.BL(BL10),.BLN(BLN10),.WL(WL24));
sram_cell_6t_5 inst_cell_24_11 (.BL(BL11),.BLN(BLN11),.WL(WL24));
sram_cell_6t_5 inst_cell_24_12 (.BL(BL12),.BLN(BLN12),.WL(WL24));
sram_cell_6t_5 inst_cell_24_13 (.BL(BL13),.BLN(BLN13),.WL(WL24));
sram_cell_6t_5 inst_cell_24_14 (.BL(BL14),.BLN(BLN14),.WL(WL24));
sram_cell_6t_5 inst_cell_24_15 (.BL(BL15),.BLN(BLN15),.WL(WL24));
sram_cell_6t_5 inst_cell_24_16 (.BL(BL16),.BLN(BLN16),.WL(WL24));
sram_cell_6t_5 inst_cell_24_17 (.BL(BL17),.BLN(BLN17),.WL(WL24));
sram_cell_6t_5 inst_cell_24_18 (.BL(BL18),.BLN(BLN18),.WL(WL24));
sram_cell_6t_5 inst_cell_24_19 (.BL(BL19),.BLN(BLN19),.WL(WL24));
sram_cell_6t_5 inst_cell_24_20 (.BL(BL20),.BLN(BLN20),.WL(WL24));
sram_cell_6t_5 inst_cell_24_21 (.BL(BL21),.BLN(BLN21),.WL(WL24));
sram_cell_6t_5 inst_cell_24_22 (.BL(BL22),.BLN(BLN22),.WL(WL24));
sram_cell_6t_5 inst_cell_24_23 (.BL(BL23),.BLN(BLN23),.WL(WL24));
sram_cell_6t_5 inst_cell_24_24 (.BL(BL24),.BLN(BLN24),.WL(WL24));
sram_cell_6t_5 inst_cell_24_25 (.BL(BL25),.BLN(BLN25),.WL(WL24));
sram_cell_6t_5 inst_cell_24_26 (.BL(BL26),.BLN(BLN26),.WL(WL24));
sram_cell_6t_5 inst_cell_24_27 (.BL(BL27),.BLN(BLN27),.WL(WL24));
sram_cell_6t_5 inst_cell_24_28 (.BL(BL28),.BLN(BLN28),.WL(WL24));
sram_cell_6t_5 inst_cell_24_29 (.BL(BL29),.BLN(BLN29),.WL(WL24));
sram_cell_6t_5 inst_cell_24_30 (.BL(BL30),.BLN(BLN30),.WL(WL24));
sram_cell_6t_5 inst_cell_24_31 (.BL(BL31),.BLN(BLN31),.WL(WL24));
sram_cell_6t_5 inst_cell_24_32 (.BL(BL32),.BLN(BLN32),.WL(WL24));
sram_cell_6t_5 inst_cell_24_33 (.BL(BL33),.BLN(BLN33),.WL(WL24));
sram_cell_6t_5 inst_cell_24_34 (.BL(BL34),.BLN(BLN34),.WL(WL24));
sram_cell_6t_5 inst_cell_24_35 (.BL(BL35),.BLN(BLN35),.WL(WL24));
sram_cell_6t_5 inst_cell_24_36 (.BL(BL36),.BLN(BLN36),.WL(WL24));
sram_cell_6t_5 inst_cell_24_37 (.BL(BL37),.BLN(BLN37),.WL(WL24));
sram_cell_6t_5 inst_cell_24_38 (.BL(BL38),.BLN(BLN38),.WL(WL24));
sram_cell_6t_5 inst_cell_24_39 (.BL(BL39),.BLN(BLN39),.WL(WL24));
sram_cell_6t_5 inst_cell_24_40 (.BL(BL40),.BLN(BLN40),.WL(WL24));
sram_cell_6t_5 inst_cell_24_41 (.BL(BL41),.BLN(BLN41),.WL(WL24));
sram_cell_6t_5 inst_cell_24_42 (.BL(BL42),.BLN(BLN42),.WL(WL24));
sram_cell_6t_5 inst_cell_24_43 (.BL(BL43),.BLN(BLN43),.WL(WL24));
sram_cell_6t_5 inst_cell_24_44 (.BL(BL44),.BLN(BLN44),.WL(WL24));
sram_cell_6t_5 inst_cell_24_45 (.BL(BL45),.BLN(BLN45),.WL(WL24));
sram_cell_6t_5 inst_cell_24_46 (.BL(BL46),.BLN(BLN46),.WL(WL24));
sram_cell_6t_5 inst_cell_24_47 (.BL(BL47),.BLN(BLN47),.WL(WL24));
sram_cell_6t_5 inst_cell_24_48 (.BL(BL48),.BLN(BLN48),.WL(WL24));
sram_cell_6t_5 inst_cell_24_49 (.BL(BL49),.BLN(BLN49),.WL(WL24));
sram_cell_6t_5 inst_cell_24_50 (.BL(BL50),.BLN(BLN50),.WL(WL24));
sram_cell_6t_5 inst_cell_24_51 (.BL(BL51),.BLN(BLN51),.WL(WL24));
sram_cell_6t_5 inst_cell_24_52 (.BL(BL52),.BLN(BLN52),.WL(WL24));
sram_cell_6t_5 inst_cell_24_53 (.BL(BL53),.BLN(BLN53),.WL(WL24));
sram_cell_6t_5 inst_cell_24_54 (.BL(BL54),.BLN(BLN54),.WL(WL24));
sram_cell_6t_5 inst_cell_24_55 (.BL(BL55),.BLN(BLN55),.WL(WL24));
sram_cell_6t_5 inst_cell_24_56 (.BL(BL56),.BLN(BLN56),.WL(WL24));
sram_cell_6t_5 inst_cell_24_57 (.BL(BL57),.BLN(BLN57),.WL(WL24));
sram_cell_6t_5 inst_cell_24_58 (.BL(BL58),.BLN(BLN58),.WL(WL24));
sram_cell_6t_5 inst_cell_24_59 (.BL(BL59),.BLN(BLN59),.WL(WL24));
sram_cell_6t_5 inst_cell_24_60 (.BL(BL60),.BLN(BLN60),.WL(WL24));
sram_cell_6t_5 inst_cell_24_61 (.BL(BL61),.BLN(BLN61),.WL(WL24));
sram_cell_6t_5 inst_cell_24_62 (.BL(BL62),.BLN(BLN62),.WL(WL24));
sram_cell_6t_5 inst_cell_24_63 (.BL(BL63),.BLN(BLN63),.WL(WL24));
sram_cell_6t_5 inst_cell_24_64 (.BL(BL64),.BLN(BLN64),.WL(WL24));
sram_cell_6t_5 inst_cell_24_65 (.BL(BL65),.BLN(BLN65),.WL(WL24));
sram_cell_6t_5 inst_cell_24_66 (.BL(BL66),.BLN(BLN66),.WL(WL24));
sram_cell_6t_5 inst_cell_24_67 (.BL(BL67),.BLN(BLN67),.WL(WL24));
sram_cell_6t_5 inst_cell_24_68 (.BL(BL68),.BLN(BLN68),.WL(WL24));
sram_cell_6t_5 inst_cell_24_69 (.BL(BL69),.BLN(BLN69),.WL(WL24));
sram_cell_6t_5 inst_cell_24_70 (.BL(BL70),.BLN(BLN70),.WL(WL24));
sram_cell_6t_5 inst_cell_24_71 (.BL(BL71),.BLN(BLN71),.WL(WL24));
sram_cell_6t_5 inst_cell_24_72 (.BL(BL72),.BLN(BLN72),.WL(WL24));
sram_cell_6t_5 inst_cell_24_73 (.BL(BL73),.BLN(BLN73),.WL(WL24));
sram_cell_6t_5 inst_cell_24_74 (.BL(BL74),.BLN(BLN74),.WL(WL24));
sram_cell_6t_5 inst_cell_24_75 (.BL(BL75),.BLN(BLN75),.WL(WL24));
sram_cell_6t_5 inst_cell_24_76 (.BL(BL76),.BLN(BLN76),.WL(WL24));
sram_cell_6t_5 inst_cell_24_77 (.BL(BL77),.BLN(BLN77),.WL(WL24));
sram_cell_6t_5 inst_cell_24_78 (.BL(BL78),.BLN(BLN78),.WL(WL24));
sram_cell_6t_5 inst_cell_24_79 (.BL(BL79),.BLN(BLN79),.WL(WL24));
sram_cell_6t_5 inst_cell_24_80 (.BL(BL80),.BLN(BLN80),.WL(WL24));
sram_cell_6t_5 inst_cell_24_81 (.BL(BL81),.BLN(BLN81),.WL(WL24));
sram_cell_6t_5 inst_cell_24_82 (.BL(BL82),.BLN(BLN82),.WL(WL24));
sram_cell_6t_5 inst_cell_24_83 (.BL(BL83),.BLN(BLN83),.WL(WL24));
sram_cell_6t_5 inst_cell_24_84 (.BL(BL84),.BLN(BLN84),.WL(WL24));
sram_cell_6t_5 inst_cell_24_85 (.BL(BL85),.BLN(BLN85),.WL(WL24));
sram_cell_6t_5 inst_cell_24_86 (.BL(BL86),.BLN(BLN86),.WL(WL24));
sram_cell_6t_5 inst_cell_24_87 (.BL(BL87),.BLN(BLN87),.WL(WL24));
sram_cell_6t_5 inst_cell_24_88 (.BL(BL88),.BLN(BLN88),.WL(WL24));
sram_cell_6t_5 inst_cell_24_89 (.BL(BL89),.BLN(BLN89),.WL(WL24));
sram_cell_6t_5 inst_cell_24_90 (.BL(BL90),.BLN(BLN90),.WL(WL24));
sram_cell_6t_5 inst_cell_24_91 (.BL(BL91),.BLN(BLN91),.WL(WL24));
sram_cell_6t_5 inst_cell_24_92 (.BL(BL92),.BLN(BLN92),.WL(WL24));
sram_cell_6t_5 inst_cell_24_93 (.BL(BL93),.BLN(BLN93),.WL(WL24));
sram_cell_6t_5 inst_cell_24_94 (.BL(BL94),.BLN(BLN94),.WL(WL24));
sram_cell_6t_5 inst_cell_24_95 (.BL(BL95),.BLN(BLN95),.WL(WL24));
sram_cell_6t_5 inst_cell_24_96 (.BL(BL96),.BLN(BLN96),.WL(WL24));
sram_cell_6t_5 inst_cell_24_97 (.BL(BL97),.BLN(BLN97),.WL(WL24));
sram_cell_6t_5 inst_cell_24_98 (.BL(BL98),.BLN(BLN98),.WL(WL24));
sram_cell_6t_5 inst_cell_24_99 (.BL(BL99),.BLN(BLN99),.WL(WL24));
sram_cell_6t_5 inst_cell_24_100 (.BL(BL100),.BLN(BLN100),.WL(WL24));
sram_cell_6t_5 inst_cell_24_101 (.BL(BL101),.BLN(BLN101),.WL(WL24));
sram_cell_6t_5 inst_cell_24_102 (.BL(BL102),.BLN(BLN102),.WL(WL24));
sram_cell_6t_5 inst_cell_24_103 (.BL(BL103),.BLN(BLN103),.WL(WL24));
sram_cell_6t_5 inst_cell_24_104 (.BL(BL104),.BLN(BLN104),.WL(WL24));
sram_cell_6t_5 inst_cell_24_105 (.BL(BL105),.BLN(BLN105),.WL(WL24));
sram_cell_6t_5 inst_cell_24_106 (.BL(BL106),.BLN(BLN106),.WL(WL24));
sram_cell_6t_5 inst_cell_24_107 (.BL(BL107),.BLN(BLN107),.WL(WL24));
sram_cell_6t_5 inst_cell_24_108 (.BL(BL108),.BLN(BLN108),.WL(WL24));
sram_cell_6t_5 inst_cell_24_109 (.BL(BL109),.BLN(BLN109),.WL(WL24));
sram_cell_6t_5 inst_cell_24_110 (.BL(BL110),.BLN(BLN110),.WL(WL24));
sram_cell_6t_5 inst_cell_24_111 (.BL(BL111),.BLN(BLN111),.WL(WL24));
sram_cell_6t_5 inst_cell_24_112 (.BL(BL112),.BLN(BLN112),.WL(WL24));
sram_cell_6t_5 inst_cell_24_113 (.BL(BL113),.BLN(BLN113),.WL(WL24));
sram_cell_6t_5 inst_cell_24_114 (.BL(BL114),.BLN(BLN114),.WL(WL24));
sram_cell_6t_5 inst_cell_24_115 (.BL(BL115),.BLN(BLN115),.WL(WL24));
sram_cell_6t_5 inst_cell_24_116 (.BL(BL116),.BLN(BLN116),.WL(WL24));
sram_cell_6t_5 inst_cell_24_117 (.BL(BL117),.BLN(BLN117),.WL(WL24));
sram_cell_6t_5 inst_cell_24_118 (.BL(BL118),.BLN(BLN118),.WL(WL24));
sram_cell_6t_5 inst_cell_24_119 (.BL(BL119),.BLN(BLN119),.WL(WL24));
sram_cell_6t_5 inst_cell_24_120 (.BL(BL120),.BLN(BLN120),.WL(WL24));
sram_cell_6t_5 inst_cell_24_121 (.BL(BL121),.BLN(BLN121),.WL(WL24));
sram_cell_6t_5 inst_cell_24_122 (.BL(BL122),.BLN(BLN122),.WL(WL24));
sram_cell_6t_5 inst_cell_24_123 (.BL(BL123),.BLN(BLN123),.WL(WL24));
sram_cell_6t_5 inst_cell_24_124 (.BL(BL124),.BLN(BLN124),.WL(WL24));
sram_cell_6t_5 inst_cell_24_125 (.BL(BL125),.BLN(BLN125),.WL(WL24));
sram_cell_6t_5 inst_cell_24_126 (.BL(BL126),.BLN(BLN126),.WL(WL24));
sram_cell_6t_5 inst_cell_24_127 (.BL(BL127),.BLN(BLN127),.WL(WL24));
sram_cell_6t_5 inst_cell_25_0 (.BL(BL0),.BLN(BLN0),.WL(WL25));
sram_cell_6t_5 inst_cell_25_1 (.BL(BL1),.BLN(BLN1),.WL(WL25));
sram_cell_6t_5 inst_cell_25_2 (.BL(BL2),.BLN(BLN2),.WL(WL25));
sram_cell_6t_5 inst_cell_25_3 (.BL(BL3),.BLN(BLN3),.WL(WL25));
sram_cell_6t_5 inst_cell_25_4 (.BL(BL4),.BLN(BLN4),.WL(WL25));
sram_cell_6t_5 inst_cell_25_5 (.BL(BL5),.BLN(BLN5),.WL(WL25));
sram_cell_6t_5 inst_cell_25_6 (.BL(BL6),.BLN(BLN6),.WL(WL25));
sram_cell_6t_5 inst_cell_25_7 (.BL(BL7),.BLN(BLN7),.WL(WL25));
sram_cell_6t_5 inst_cell_25_8 (.BL(BL8),.BLN(BLN8),.WL(WL25));
sram_cell_6t_5 inst_cell_25_9 (.BL(BL9),.BLN(BLN9),.WL(WL25));
sram_cell_6t_5 inst_cell_25_10 (.BL(BL10),.BLN(BLN10),.WL(WL25));
sram_cell_6t_5 inst_cell_25_11 (.BL(BL11),.BLN(BLN11),.WL(WL25));
sram_cell_6t_5 inst_cell_25_12 (.BL(BL12),.BLN(BLN12),.WL(WL25));
sram_cell_6t_5 inst_cell_25_13 (.BL(BL13),.BLN(BLN13),.WL(WL25));
sram_cell_6t_5 inst_cell_25_14 (.BL(BL14),.BLN(BLN14),.WL(WL25));
sram_cell_6t_5 inst_cell_25_15 (.BL(BL15),.BLN(BLN15),.WL(WL25));
sram_cell_6t_5 inst_cell_25_16 (.BL(BL16),.BLN(BLN16),.WL(WL25));
sram_cell_6t_5 inst_cell_25_17 (.BL(BL17),.BLN(BLN17),.WL(WL25));
sram_cell_6t_5 inst_cell_25_18 (.BL(BL18),.BLN(BLN18),.WL(WL25));
sram_cell_6t_5 inst_cell_25_19 (.BL(BL19),.BLN(BLN19),.WL(WL25));
sram_cell_6t_5 inst_cell_25_20 (.BL(BL20),.BLN(BLN20),.WL(WL25));
sram_cell_6t_5 inst_cell_25_21 (.BL(BL21),.BLN(BLN21),.WL(WL25));
sram_cell_6t_5 inst_cell_25_22 (.BL(BL22),.BLN(BLN22),.WL(WL25));
sram_cell_6t_5 inst_cell_25_23 (.BL(BL23),.BLN(BLN23),.WL(WL25));
sram_cell_6t_5 inst_cell_25_24 (.BL(BL24),.BLN(BLN24),.WL(WL25));
sram_cell_6t_5 inst_cell_25_25 (.BL(BL25),.BLN(BLN25),.WL(WL25));
sram_cell_6t_5 inst_cell_25_26 (.BL(BL26),.BLN(BLN26),.WL(WL25));
sram_cell_6t_5 inst_cell_25_27 (.BL(BL27),.BLN(BLN27),.WL(WL25));
sram_cell_6t_5 inst_cell_25_28 (.BL(BL28),.BLN(BLN28),.WL(WL25));
sram_cell_6t_5 inst_cell_25_29 (.BL(BL29),.BLN(BLN29),.WL(WL25));
sram_cell_6t_5 inst_cell_25_30 (.BL(BL30),.BLN(BLN30),.WL(WL25));
sram_cell_6t_5 inst_cell_25_31 (.BL(BL31),.BLN(BLN31),.WL(WL25));
sram_cell_6t_5 inst_cell_25_32 (.BL(BL32),.BLN(BLN32),.WL(WL25));
sram_cell_6t_5 inst_cell_25_33 (.BL(BL33),.BLN(BLN33),.WL(WL25));
sram_cell_6t_5 inst_cell_25_34 (.BL(BL34),.BLN(BLN34),.WL(WL25));
sram_cell_6t_5 inst_cell_25_35 (.BL(BL35),.BLN(BLN35),.WL(WL25));
sram_cell_6t_5 inst_cell_25_36 (.BL(BL36),.BLN(BLN36),.WL(WL25));
sram_cell_6t_5 inst_cell_25_37 (.BL(BL37),.BLN(BLN37),.WL(WL25));
sram_cell_6t_5 inst_cell_25_38 (.BL(BL38),.BLN(BLN38),.WL(WL25));
sram_cell_6t_5 inst_cell_25_39 (.BL(BL39),.BLN(BLN39),.WL(WL25));
sram_cell_6t_5 inst_cell_25_40 (.BL(BL40),.BLN(BLN40),.WL(WL25));
sram_cell_6t_5 inst_cell_25_41 (.BL(BL41),.BLN(BLN41),.WL(WL25));
sram_cell_6t_5 inst_cell_25_42 (.BL(BL42),.BLN(BLN42),.WL(WL25));
sram_cell_6t_5 inst_cell_25_43 (.BL(BL43),.BLN(BLN43),.WL(WL25));
sram_cell_6t_5 inst_cell_25_44 (.BL(BL44),.BLN(BLN44),.WL(WL25));
sram_cell_6t_5 inst_cell_25_45 (.BL(BL45),.BLN(BLN45),.WL(WL25));
sram_cell_6t_5 inst_cell_25_46 (.BL(BL46),.BLN(BLN46),.WL(WL25));
sram_cell_6t_5 inst_cell_25_47 (.BL(BL47),.BLN(BLN47),.WL(WL25));
sram_cell_6t_5 inst_cell_25_48 (.BL(BL48),.BLN(BLN48),.WL(WL25));
sram_cell_6t_5 inst_cell_25_49 (.BL(BL49),.BLN(BLN49),.WL(WL25));
sram_cell_6t_5 inst_cell_25_50 (.BL(BL50),.BLN(BLN50),.WL(WL25));
sram_cell_6t_5 inst_cell_25_51 (.BL(BL51),.BLN(BLN51),.WL(WL25));
sram_cell_6t_5 inst_cell_25_52 (.BL(BL52),.BLN(BLN52),.WL(WL25));
sram_cell_6t_5 inst_cell_25_53 (.BL(BL53),.BLN(BLN53),.WL(WL25));
sram_cell_6t_5 inst_cell_25_54 (.BL(BL54),.BLN(BLN54),.WL(WL25));
sram_cell_6t_5 inst_cell_25_55 (.BL(BL55),.BLN(BLN55),.WL(WL25));
sram_cell_6t_5 inst_cell_25_56 (.BL(BL56),.BLN(BLN56),.WL(WL25));
sram_cell_6t_5 inst_cell_25_57 (.BL(BL57),.BLN(BLN57),.WL(WL25));
sram_cell_6t_5 inst_cell_25_58 (.BL(BL58),.BLN(BLN58),.WL(WL25));
sram_cell_6t_5 inst_cell_25_59 (.BL(BL59),.BLN(BLN59),.WL(WL25));
sram_cell_6t_5 inst_cell_25_60 (.BL(BL60),.BLN(BLN60),.WL(WL25));
sram_cell_6t_5 inst_cell_25_61 (.BL(BL61),.BLN(BLN61),.WL(WL25));
sram_cell_6t_5 inst_cell_25_62 (.BL(BL62),.BLN(BLN62),.WL(WL25));
sram_cell_6t_5 inst_cell_25_63 (.BL(BL63),.BLN(BLN63),.WL(WL25));
sram_cell_6t_5 inst_cell_25_64 (.BL(BL64),.BLN(BLN64),.WL(WL25));
sram_cell_6t_5 inst_cell_25_65 (.BL(BL65),.BLN(BLN65),.WL(WL25));
sram_cell_6t_5 inst_cell_25_66 (.BL(BL66),.BLN(BLN66),.WL(WL25));
sram_cell_6t_5 inst_cell_25_67 (.BL(BL67),.BLN(BLN67),.WL(WL25));
sram_cell_6t_5 inst_cell_25_68 (.BL(BL68),.BLN(BLN68),.WL(WL25));
sram_cell_6t_5 inst_cell_25_69 (.BL(BL69),.BLN(BLN69),.WL(WL25));
sram_cell_6t_5 inst_cell_25_70 (.BL(BL70),.BLN(BLN70),.WL(WL25));
sram_cell_6t_5 inst_cell_25_71 (.BL(BL71),.BLN(BLN71),.WL(WL25));
sram_cell_6t_5 inst_cell_25_72 (.BL(BL72),.BLN(BLN72),.WL(WL25));
sram_cell_6t_5 inst_cell_25_73 (.BL(BL73),.BLN(BLN73),.WL(WL25));
sram_cell_6t_5 inst_cell_25_74 (.BL(BL74),.BLN(BLN74),.WL(WL25));
sram_cell_6t_5 inst_cell_25_75 (.BL(BL75),.BLN(BLN75),.WL(WL25));
sram_cell_6t_5 inst_cell_25_76 (.BL(BL76),.BLN(BLN76),.WL(WL25));
sram_cell_6t_5 inst_cell_25_77 (.BL(BL77),.BLN(BLN77),.WL(WL25));
sram_cell_6t_5 inst_cell_25_78 (.BL(BL78),.BLN(BLN78),.WL(WL25));
sram_cell_6t_5 inst_cell_25_79 (.BL(BL79),.BLN(BLN79),.WL(WL25));
sram_cell_6t_5 inst_cell_25_80 (.BL(BL80),.BLN(BLN80),.WL(WL25));
sram_cell_6t_5 inst_cell_25_81 (.BL(BL81),.BLN(BLN81),.WL(WL25));
sram_cell_6t_5 inst_cell_25_82 (.BL(BL82),.BLN(BLN82),.WL(WL25));
sram_cell_6t_5 inst_cell_25_83 (.BL(BL83),.BLN(BLN83),.WL(WL25));
sram_cell_6t_5 inst_cell_25_84 (.BL(BL84),.BLN(BLN84),.WL(WL25));
sram_cell_6t_5 inst_cell_25_85 (.BL(BL85),.BLN(BLN85),.WL(WL25));
sram_cell_6t_5 inst_cell_25_86 (.BL(BL86),.BLN(BLN86),.WL(WL25));
sram_cell_6t_5 inst_cell_25_87 (.BL(BL87),.BLN(BLN87),.WL(WL25));
sram_cell_6t_5 inst_cell_25_88 (.BL(BL88),.BLN(BLN88),.WL(WL25));
sram_cell_6t_5 inst_cell_25_89 (.BL(BL89),.BLN(BLN89),.WL(WL25));
sram_cell_6t_5 inst_cell_25_90 (.BL(BL90),.BLN(BLN90),.WL(WL25));
sram_cell_6t_5 inst_cell_25_91 (.BL(BL91),.BLN(BLN91),.WL(WL25));
sram_cell_6t_5 inst_cell_25_92 (.BL(BL92),.BLN(BLN92),.WL(WL25));
sram_cell_6t_5 inst_cell_25_93 (.BL(BL93),.BLN(BLN93),.WL(WL25));
sram_cell_6t_5 inst_cell_25_94 (.BL(BL94),.BLN(BLN94),.WL(WL25));
sram_cell_6t_5 inst_cell_25_95 (.BL(BL95),.BLN(BLN95),.WL(WL25));
sram_cell_6t_5 inst_cell_25_96 (.BL(BL96),.BLN(BLN96),.WL(WL25));
sram_cell_6t_5 inst_cell_25_97 (.BL(BL97),.BLN(BLN97),.WL(WL25));
sram_cell_6t_5 inst_cell_25_98 (.BL(BL98),.BLN(BLN98),.WL(WL25));
sram_cell_6t_5 inst_cell_25_99 (.BL(BL99),.BLN(BLN99),.WL(WL25));
sram_cell_6t_5 inst_cell_25_100 (.BL(BL100),.BLN(BLN100),.WL(WL25));
sram_cell_6t_5 inst_cell_25_101 (.BL(BL101),.BLN(BLN101),.WL(WL25));
sram_cell_6t_5 inst_cell_25_102 (.BL(BL102),.BLN(BLN102),.WL(WL25));
sram_cell_6t_5 inst_cell_25_103 (.BL(BL103),.BLN(BLN103),.WL(WL25));
sram_cell_6t_5 inst_cell_25_104 (.BL(BL104),.BLN(BLN104),.WL(WL25));
sram_cell_6t_5 inst_cell_25_105 (.BL(BL105),.BLN(BLN105),.WL(WL25));
sram_cell_6t_5 inst_cell_25_106 (.BL(BL106),.BLN(BLN106),.WL(WL25));
sram_cell_6t_5 inst_cell_25_107 (.BL(BL107),.BLN(BLN107),.WL(WL25));
sram_cell_6t_5 inst_cell_25_108 (.BL(BL108),.BLN(BLN108),.WL(WL25));
sram_cell_6t_5 inst_cell_25_109 (.BL(BL109),.BLN(BLN109),.WL(WL25));
sram_cell_6t_5 inst_cell_25_110 (.BL(BL110),.BLN(BLN110),.WL(WL25));
sram_cell_6t_5 inst_cell_25_111 (.BL(BL111),.BLN(BLN111),.WL(WL25));
sram_cell_6t_5 inst_cell_25_112 (.BL(BL112),.BLN(BLN112),.WL(WL25));
sram_cell_6t_5 inst_cell_25_113 (.BL(BL113),.BLN(BLN113),.WL(WL25));
sram_cell_6t_5 inst_cell_25_114 (.BL(BL114),.BLN(BLN114),.WL(WL25));
sram_cell_6t_5 inst_cell_25_115 (.BL(BL115),.BLN(BLN115),.WL(WL25));
sram_cell_6t_5 inst_cell_25_116 (.BL(BL116),.BLN(BLN116),.WL(WL25));
sram_cell_6t_5 inst_cell_25_117 (.BL(BL117),.BLN(BLN117),.WL(WL25));
sram_cell_6t_5 inst_cell_25_118 (.BL(BL118),.BLN(BLN118),.WL(WL25));
sram_cell_6t_5 inst_cell_25_119 (.BL(BL119),.BLN(BLN119),.WL(WL25));
sram_cell_6t_5 inst_cell_25_120 (.BL(BL120),.BLN(BLN120),.WL(WL25));
sram_cell_6t_5 inst_cell_25_121 (.BL(BL121),.BLN(BLN121),.WL(WL25));
sram_cell_6t_5 inst_cell_25_122 (.BL(BL122),.BLN(BLN122),.WL(WL25));
sram_cell_6t_5 inst_cell_25_123 (.BL(BL123),.BLN(BLN123),.WL(WL25));
sram_cell_6t_5 inst_cell_25_124 (.BL(BL124),.BLN(BLN124),.WL(WL25));
sram_cell_6t_5 inst_cell_25_125 (.BL(BL125),.BLN(BLN125),.WL(WL25));
sram_cell_6t_5 inst_cell_25_126 (.BL(BL126),.BLN(BLN126),.WL(WL25));
sram_cell_6t_5 inst_cell_25_127 (.BL(BL127),.BLN(BLN127),.WL(WL25));
sram_cell_6t_5 inst_cell_26_0 (.BL(BL0),.BLN(BLN0),.WL(WL26));
sram_cell_6t_5 inst_cell_26_1 (.BL(BL1),.BLN(BLN1),.WL(WL26));
sram_cell_6t_5 inst_cell_26_2 (.BL(BL2),.BLN(BLN2),.WL(WL26));
sram_cell_6t_5 inst_cell_26_3 (.BL(BL3),.BLN(BLN3),.WL(WL26));
sram_cell_6t_5 inst_cell_26_4 (.BL(BL4),.BLN(BLN4),.WL(WL26));
sram_cell_6t_5 inst_cell_26_5 (.BL(BL5),.BLN(BLN5),.WL(WL26));
sram_cell_6t_5 inst_cell_26_6 (.BL(BL6),.BLN(BLN6),.WL(WL26));
sram_cell_6t_5 inst_cell_26_7 (.BL(BL7),.BLN(BLN7),.WL(WL26));
sram_cell_6t_5 inst_cell_26_8 (.BL(BL8),.BLN(BLN8),.WL(WL26));
sram_cell_6t_5 inst_cell_26_9 (.BL(BL9),.BLN(BLN9),.WL(WL26));
sram_cell_6t_5 inst_cell_26_10 (.BL(BL10),.BLN(BLN10),.WL(WL26));
sram_cell_6t_5 inst_cell_26_11 (.BL(BL11),.BLN(BLN11),.WL(WL26));
sram_cell_6t_5 inst_cell_26_12 (.BL(BL12),.BLN(BLN12),.WL(WL26));
sram_cell_6t_5 inst_cell_26_13 (.BL(BL13),.BLN(BLN13),.WL(WL26));
sram_cell_6t_5 inst_cell_26_14 (.BL(BL14),.BLN(BLN14),.WL(WL26));
sram_cell_6t_5 inst_cell_26_15 (.BL(BL15),.BLN(BLN15),.WL(WL26));
sram_cell_6t_5 inst_cell_26_16 (.BL(BL16),.BLN(BLN16),.WL(WL26));
sram_cell_6t_5 inst_cell_26_17 (.BL(BL17),.BLN(BLN17),.WL(WL26));
sram_cell_6t_5 inst_cell_26_18 (.BL(BL18),.BLN(BLN18),.WL(WL26));
sram_cell_6t_5 inst_cell_26_19 (.BL(BL19),.BLN(BLN19),.WL(WL26));
sram_cell_6t_5 inst_cell_26_20 (.BL(BL20),.BLN(BLN20),.WL(WL26));
sram_cell_6t_5 inst_cell_26_21 (.BL(BL21),.BLN(BLN21),.WL(WL26));
sram_cell_6t_5 inst_cell_26_22 (.BL(BL22),.BLN(BLN22),.WL(WL26));
sram_cell_6t_5 inst_cell_26_23 (.BL(BL23),.BLN(BLN23),.WL(WL26));
sram_cell_6t_5 inst_cell_26_24 (.BL(BL24),.BLN(BLN24),.WL(WL26));
sram_cell_6t_5 inst_cell_26_25 (.BL(BL25),.BLN(BLN25),.WL(WL26));
sram_cell_6t_5 inst_cell_26_26 (.BL(BL26),.BLN(BLN26),.WL(WL26));
sram_cell_6t_5 inst_cell_26_27 (.BL(BL27),.BLN(BLN27),.WL(WL26));
sram_cell_6t_5 inst_cell_26_28 (.BL(BL28),.BLN(BLN28),.WL(WL26));
sram_cell_6t_5 inst_cell_26_29 (.BL(BL29),.BLN(BLN29),.WL(WL26));
sram_cell_6t_5 inst_cell_26_30 (.BL(BL30),.BLN(BLN30),.WL(WL26));
sram_cell_6t_5 inst_cell_26_31 (.BL(BL31),.BLN(BLN31),.WL(WL26));
sram_cell_6t_5 inst_cell_26_32 (.BL(BL32),.BLN(BLN32),.WL(WL26));
sram_cell_6t_5 inst_cell_26_33 (.BL(BL33),.BLN(BLN33),.WL(WL26));
sram_cell_6t_5 inst_cell_26_34 (.BL(BL34),.BLN(BLN34),.WL(WL26));
sram_cell_6t_5 inst_cell_26_35 (.BL(BL35),.BLN(BLN35),.WL(WL26));
sram_cell_6t_5 inst_cell_26_36 (.BL(BL36),.BLN(BLN36),.WL(WL26));
sram_cell_6t_5 inst_cell_26_37 (.BL(BL37),.BLN(BLN37),.WL(WL26));
sram_cell_6t_5 inst_cell_26_38 (.BL(BL38),.BLN(BLN38),.WL(WL26));
sram_cell_6t_5 inst_cell_26_39 (.BL(BL39),.BLN(BLN39),.WL(WL26));
sram_cell_6t_5 inst_cell_26_40 (.BL(BL40),.BLN(BLN40),.WL(WL26));
sram_cell_6t_5 inst_cell_26_41 (.BL(BL41),.BLN(BLN41),.WL(WL26));
sram_cell_6t_5 inst_cell_26_42 (.BL(BL42),.BLN(BLN42),.WL(WL26));
sram_cell_6t_5 inst_cell_26_43 (.BL(BL43),.BLN(BLN43),.WL(WL26));
sram_cell_6t_5 inst_cell_26_44 (.BL(BL44),.BLN(BLN44),.WL(WL26));
sram_cell_6t_5 inst_cell_26_45 (.BL(BL45),.BLN(BLN45),.WL(WL26));
sram_cell_6t_5 inst_cell_26_46 (.BL(BL46),.BLN(BLN46),.WL(WL26));
sram_cell_6t_5 inst_cell_26_47 (.BL(BL47),.BLN(BLN47),.WL(WL26));
sram_cell_6t_5 inst_cell_26_48 (.BL(BL48),.BLN(BLN48),.WL(WL26));
sram_cell_6t_5 inst_cell_26_49 (.BL(BL49),.BLN(BLN49),.WL(WL26));
sram_cell_6t_5 inst_cell_26_50 (.BL(BL50),.BLN(BLN50),.WL(WL26));
sram_cell_6t_5 inst_cell_26_51 (.BL(BL51),.BLN(BLN51),.WL(WL26));
sram_cell_6t_5 inst_cell_26_52 (.BL(BL52),.BLN(BLN52),.WL(WL26));
sram_cell_6t_5 inst_cell_26_53 (.BL(BL53),.BLN(BLN53),.WL(WL26));
sram_cell_6t_5 inst_cell_26_54 (.BL(BL54),.BLN(BLN54),.WL(WL26));
sram_cell_6t_5 inst_cell_26_55 (.BL(BL55),.BLN(BLN55),.WL(WL26));
sram_cell_6t_5 inst_cell_26_56 (.BL(BL56),.BLN(BLN56),.WL(WL26));
sram_cell_6t_5 inst_cell_26_57 (.BL(BL57),.BLN(BLN57),.WL(WL26));
sram_cell_6t_5 inst_cell_26_58 (.BL(BL58),.BLN(BLN58),.WL(WL26));
sram_cell_6t_5 inst_cell_26_59 (.BL(BL59),.BLN(BLN59),.WL(WL26));
sram_cell_6t_5 inst_cell_26_60 (.BL(BL60),.BLN(BLN60),.WL(WL26));
sram_cell_6t_5 inst_cell_26_61 (.BL(BL61),.BLN(BLN61),.WL(WL26));
sram_cell_6t_5 inst_cell_26_62 (.BL(BL62),.BLN(BLN62),.WL(WL26));
sram_cell_6t_5 inst_cell_26_63 (.BL(BL63),.BLN(BLN63),.WL(WL26));
sram_cell_6t_5 inst_cell_26_64 (.BL(BL64),.BLN(BLN64),.WL(WL26));
sram_cell_6t_5 inst_cell_26_65 (.BL(BL65),.BLN(BLN65),.WL(WL26));
sram_cell_6t_5 inst_cell_26_66 (.BL(BL66),.BLN(BLN66),.WL(WL26));
sram_cell_6t_5 inst_cell_26_67 (.BL(BL67),.BLN(BLN67),.WL(WL26));
sram_cell_6t_5 inst_cell_26_68 (.BL(BL68),.BLN(BLN68),.WL(WL26));
sram_cell_6t_5 inst_cell_26_69 (.BL(BL69),.BLN(BLN69),.WL(WL26));
sram_cell_6t_5 inst_cell_26_70 (.BL(BL70),.BLN(BLN70),.WL(WL26));
sram_cell_6t_5 inst_cell_26_71 (.BL(BL71),.BLN(BLN71),.WL(WL26));
sram_cell_6t_5 inst_cell_26_72 (.BL(BL72),.BLN(BLN72),.WL(WL26));
sram_cell_6t_5 inst_cell_26_73 (.BL(BL73),.BLN(BLN73),.WL(WL26));
sram_cell_6t_5 inst_cell_26_74 (.BL(BL74),.BLN(BLN74),.WL(WL26));
sram_cell_6t_5 inst_cell_26_75 (.BL(BL75),.BLN(BLN75),.WL(WL26));
sram_cell_6t_5 inst_cell_26_76 (.BL(BL76),.BLN(BLN76),.WL(WL26));
sram_cell_6t_5 inst_cell_26_77 (.BL(BL77),.BLN(BLN77),.WL(WL26));
sram_cell_6t_5 inst_cell_26_78 (.BL(BL78),.BLN(BLN78),.WL(WL26));
sram_cell_6t_5 inst_cell_26_79 (.BL(BL79),.BLN(BLN79),.WL(WL26));
sram_cell_6t_5 inst_cell_26_80 (.BL(BL80),.BLN(BLN80),.WL(WL26));
sram_cell_6t_5 inst_cell_26_81 (.BL(BL81),.BLN(BLN81),.WL(WL26));
sram_cell_6t_5 inst_cell_26_82 (.BL(BL82),.BLN(BLN82),.WL(WL26));
sram_cell_6t_5 inst_cell_26_83 (.BL(BL83),.BLN(BLN83),.WL(WL26));
sram_cell_6t_5 inst_cell_26_84 (.BL(BL84),.BLN(BLN84),.WL(WL26));
sram_cell_6t_5 inst_cell_26_85 (.BL(BL85),.BLN(BLN85),.WL(WL26));
sram_cell_6t_5 inst_cell_26_86 (.BL(BL86),.BLN(BLN86),.WL(WL26));
sram_cell_6t_5 inst_cell_26_87 (.BL(BL87),.BLN(BLN87),.WL(WL26));
sram_cell_6t_5 inst_cell_26_88 (.BL(BL88),.BLN(BLN88),.WL(WL26));
sram_cell_6t_5 inst_cell_26_89 (.BL(BL89),.BLN(BLN89),.WL(WL26));
sram_cell_6t_5 inst_cell_26_90 (.BL(BL90),.BLN(BLN90),.WL(WL26));
sram_cell_6t_5 inst_cell_26_91 (.BL(BL91),.BLN(BLN91),.WL(WL26));
sram_cell_6t_5 inst_cell_26_92 (.BL(BL92),.BLN(BLN92),.WL(WL26));
sram_cell_6t_5 inst_cell_26_93 (.BL(BL93),.BLN(BLN93),.WL(WL26));
sram_cell_6t_5 inst_cell_26_94 (.BL(BL94),.BLN(BLN94),.WL(WL26));
sram_cell_6t_5 inst_cell_26_95 (.BL(BL95),.BLN(BLN95),.WL(WL26));
sram_cell_6t_5 inst_cell_26_96 (.BL(BL96),.BLN(BLN96),.WL(WL26));
sram_cell_6t_5 inst_cell_26_97 (.BL(BL97),.BLN(BLN97),.WL(WL26));
sram_cell_6t_5 inst_cell_26_98 (.BL(BL98),.BLN(BLN98),.WL(WL26));
sram_cell_6t_5 inst_cell_26_99 (.BL(BL99),.BLN(BLN99),.WL(WL26));
sram_cell_6t_5 inst_cell_26_100 (.BL(BL100),.BLN(BLN100),.WL(WL26));
sram_cell_6t_5 inst_cell_26_101 (.BL(BL101),.BLN(BLN101),.WL(WL26));
sram_cell_6t_5 inst_cell_26_102 (.BL(BL102),.BLN(BLN102),.WL(WL26));
sram_cell_6t_5 inst_cell_26_103 (.BL(BL103),.BLN(BLN103),.WL(WL26));
sram_cell_6t_5 inst_cell_26_104 (.BL(BL104),.BLN(BLN104),.WL(WL26));
sram_cell_6t_5 inst_cell_26_105 (.BL(BL105),.BLN(BLN105),.WL(WL26));
sram_cell_6t_5 inst_cell_26_106 (.BL(BL106),.BLN(BLN106),.WL(WL26));
sram_cell_6t_5 inst_cell_26_107 (.BL(BL107),.BLN(BLN107),.WL(WL26));
sram_cell_6t_5 inst_cell_26_108 (.BL(BL108),.BLN(BLN108),.WL(WL26));
sram_cell_6t_5 inst_cell_26_109 (.BL(BL109),.BLN(BLN109),.WL(WL26));
sram_cell_6t_5 inst_cell_26_110 (.BL(BL110),.BLN(BLN110),.WL(WL26));
sram_cell_6t_5 inst_cell_26_111 (.BL(BL111),.BLN(BLN111),.WL(WL26));
sram_cell_6t_5 inst_cell_26_112 (.BL(BL112),.BLN(BLN112),.WL(WL26));
sram_cell_6t_5 inst_cell_26_113 (.BL(BL113),.BLN(BLN113),.WL(WL26));
sram_cell_6t_5 inst_cell_26_114 (.BL(BL114),.BLN(BLN114),.WL(WL26));
sram_cell_6t_5 inst_cell_26_115 (.BL(BL115),.BLN(BLN115),.WL(WL26));
sram_cell_6t_5 inst_cell_26_116 (.BL(BL116),.BLN(BLN116),.WL(WL26));
sram_cell_6t_5 inst_cell_26_117 (.BL(BL117),.BLN(BLN117),.WL(WL26));
sram_cell_6t_5 inst_cell_26_118 (.BL(BL118),.BLN(BLN118),.WL(WL26));
sram_cell_6t_5 inst_cell_26_119 (.BL(BL119),.BLN(BLN119),.WL(WL26));
sram_cell_6t_5 inst_cell_26_120 (.BL(BL120),.BLN(BLN120),.WL(WL26));
sram_cell_6t_5 inst_cell_26_121 (.BL(BL121),.BLN(BLN121),.WL(WL26));
sram_cell_6t_5 inst_cell_26_122 (.BL(BL122),.BLN(BLN122),.WL(WL26));
sram_cell_6t_5 inst_cell_26_123 (.BL(BL123),.BLN(BLN123),.WL(WL26));
sram_cell_6t_5 inst_cell_26_124 (.BL(BL124),.BLN(BLN124),.WL(WL26));
sram_cell_6t_5 inst_cell_26_125 (.BL(BL125),.BLN(BLN125),.WL(WL26));
sram_cell_6t_5 inst_cell_26_126 (.BL(BL126),.BLN(BLN126),.WL(WL26));
sram_cell_6t_5 inst_cell_26_127 (.BL(BL127),.BLN(BLN127),.WL(WL26));
sram_cell_6t_5 inst_cell_27_0 (.BL(BL0),.BLN(BLN0),.WL(WL27));
sram_cell_6t_5 inst_cell_27_1 (.BL(BL1),.BLN(BLN1),.WL(WL27));
sram_cell_6t_5 inst_cell_27_2 (.BL(BL2),.BLN(BLN2),.WL(WL27));
sram_cell_6t_5 inst_cell_27_3 (.BL(BL3),.BLN(BLN3),.WL(WL27));
sram_cell_6t_5 inst_cell_27_4 (.BL(BL4),.BLN(BLN4),.WL(WL27));
sram_cell_6t_5 inst_cell_27_5 (.BL(BL5),.BLN(BLN5),.WL(WL27));
sram_cell_6t_5 inst_cell_27_6 (.BL(BL6),.BLN(BLN6),.WL(WL27));
sram_cell_6t_5 inst_cell_27_7 (.BL(BL7),.BLN(BLN7),.WL(WL27));
sram_cell_6t_5 inst_cell_27_8 (.BL(BL8),.BLN(BLN8),.WL(WL27));
sram_cell_6t_5 inst_cell_27_9 (.BL(BL9),.BLN(BLN9),.WL(WL27));
sram_cell_6t_5 inst_cell_27_10 (.BL(BL10),.BLN(BLN10),.WL(WL27));
sram_cell_6t_5 inst_cell_27_11 (.BL(BL11),.BLN(BLN11),.WL(WL27));
sram_cell_6t_5 inst_cell_27_12 (.BL(BL12),.BLN(BLN12),.WL(WL27));
sram_cell_6t_5 inst_cell_27_13 (.BL(BL13),.BLN(BLN13),.WL(WL27));
sram_cell_6t_5 inst_cell_27_14 (.BL(BL14),.BLN(BLN14),.WL(WL27));
sram_cell_6t_5 inst_cell_27_15 (.BL(BL15),.BLN(BLN15),.WL(WL27));
sram_cell_6t_5 inst_cell_27_16 (.BL(BL16),.BLN(BLN16),.WL(WL27));
sram_cell_6t_5 inst_cell_27_17 (.BL(BL17),.BLN(BLN17),.WL(WL27));
sram_cell_6t_5 inst_cell_27_18 (.BL(BL18),.BLN(BLN18),.WL(WL27));
sram_cell_6t_5 inst_cell_27_19 (.BL(BL19),.BLN(BLN19),.WL(WL27));
sram_cell_6t_5 inst_cell_27_20 (.BL(BL20),.BLN(BLN20),.WL(WL27));
sram_cell_6t_5 inst_cell_27_21 (.BL(BL21),.BLN(BLN21),.WL(WL27));
sram_cell_6t_5 inst_cell_27_22 (.BL(BL22),.BLN(BLN22),.WL(WL27));
sram_cell_6t_5 inst_cell_27_23 (.BL(BL23),.BLN(BLN23),.WL(WL27));
sram_cell_6t_5 inst_cell_27_24 (.BL(BL24),.BLN(BLN24),.WL(WL27));
sram_cell_6t_5 inst_cell_27_25 (.BL(BL25),.BLN(BLN25),.WL(WL27));
sram_cell_6t_5 inst_cell_27_26 (.BL(BL26),.BLN(BLN26),.WL(WL27));
sram_cell_6t_5 inst_cell_27_27 (.BL(BL27),.BLN(BLN27),.WL(WL27));
sram_cell_6t_5 inst_cell_27_28 (.BL(BL28),.BLN(BLN28),.WL(WL27));
sram_cell_6t_5 inst_cell_27_29 (.BL(BL29),.BLN(BLN29),.WL(WL27));
sram_cell_6t_5 inst_cell_27_30 (.BL(BL30),.BLN(BLN30),.WL(WL27));
sram_cell_6t_5 inst_cell_27_31 (.BL(BL31),.BLN(BLN31),.WL(WL27));
sram_cell_6t_5 inst_cell_27_32 (.BL(BL32),.BLN(BLN32),.WL(WL27));
sram_cell_6t_5 inst_cell_27_33 (.BL(BL33),.BLN(BLN33),.WL(WL27));
sram_cell_6t_5 inst_cell_27_34 (.BL(BL34),.BLN(BLN34),.WL(WL27));
sram_cell_6t_5 inst_cell_27_35 (.BL(BL35),.BLN(BLN35),.WL(WL27));
sram_cell_6t_5 inst_cell_27_36 (.BL(BL36),.BLN(BLN36),.WL(WL27));
sram_cell_6t_5 inst_cell_27_37 (.BL(BL37),.BLN(BLN37),.WL(WL27));
sram_cell_6t_5 inst_cell_27_38 (.BL(BL38),.BLN(BLN38),.WL(WL27));
sram_cell_6t_5 inst_cell_27_39 (.BL(BL39),.BLN(BLN39),.WL(WL27));
sram_cell_6t_5 inst_cell_27_40 (.BL(BL40),.BLN(BLN40),.WL(WL27));
sram_cell_6t_5 inst_cell_27_41 (.BL(BL41),.BLN(BLN41),.WL(WL27));
sram_cell_6t_5 inst_cell_27_42 (.BL(BL42),.BLN(BLN42),.WL(WL27));
sram_cell_6t_5 inst_cell_27_43 (.BL(BL43),.BLN(BLN43),.WL(WL27));
sram_cell_6t_5 inst_cell_27_44 (.BL(BL44),.BLN(BLN44),.WL(WL27));
sram_cell_6t_5 inst_cell_27_45 (.BL(BL45),.BLN(BLN45),.WL(WL27));
sram_cell_6t_5 inst_cell_27_46 (.BL(BL46),.BLN(BLN46),.WL(WL27));
sram_cell_6t_5 inst_cell_27_47 (.BL(BL47),.BLN(BLN47),.WL(WL27));
sram_cell_6t_5 inst_cell_27_48 (.BL(BL48),.BLN(BLN48),.WL(WL27));
sram_cell_6t_5 inst_cell_27_49 (.BL(BL49),.BLN(BLN49),.WL(WL27));
sram_cell_6t_5 inst_cell_27_50 (.BL(BL50),.BLN(BLN50),.WL(WL27));
sram_cell_6t_5 inst_cell_27_51 (.BL(BL51),.BLN(BLN51),.WL(WL27));
sram_cell_6t_5 inst_cell_27_52 (.BL(BL52),.BLN(BLN52),.WL(WL27));
sram_cell_6t_5 inst_cell_27_53 (.BL(BL53),.BLN(BLN53),.WL(WL27));
sram_cell_6t_5 inst_cell_27_54 (.BL(BL54),.BLN(BLN54),.WL(WL27));
sram_cell_6t_5 inst_cell_27_55 (.BL(BL55),.BLN(BLN55),.WL(WL27));
sram_cell_6t_5 inst_cell_27_56 (.BL(BL56),.BLN(BLN56),.WL(WL27));
sram_cell_6t_5 inst_cell_27_57 (.BL(BL57),.BLN(BLN57),.WL(WL27));
sram_cell_6t_5 inst_cell_27_58 (.BL(BL58),.BLN(BLN58),.WL(WL27));
sram_cell_6t_5 inst_cell_27_59 (.BL(BL59),.BLN(BLN59),.WL(WL27));
sram_cell_6t_5 inst_cell_27_60 (.BL(BL60),.BLN(BLN60),.WL(WL27));
sram_cell_6t_5 inst_cell_27_61 (.BL(BL61),.BLN(BLN61),.WL(WL27));
sram_cell_6t_5 inst_cell_27_62 (.BL(BL62),.BLN(BLN62),.WL(WL27));
sram_cell_6t_5 inst_cell_27_63 (.BL(BL63),.BLN(BLN63),.WL(WL27));
sram_cell_6t_5 inst_cell_27_64 (.BL(BL64),.BLN(BLN64),.WL(WL27));
sram_cell_6t_5 inst_cell_27_65 (.BL(BL65),.BLN(BLN65),.WL(WL27));
sram_cell_6t_5 inst_cell_27_66 (.BL(BL66),.BLN(BLN66),.WL(WL27));
sram_cell_6t_5 inst_cell_27_67 (.BL(BL67),.BLN(BLN67),.WL(WL27));
sram_cell_6t_5 inst_cell_27_68 (.BL(BL68),.BLN(BLN68),.WL(WL27));
sram_cell_6t_5 inst_cell_27_69 (.BL(BL69),.BLN(BLN69),.WL(WL27));
sram_cell_6t_5 inst_cell_27_70 (.BL(BL70),.BLN(BLN70),.WL(WL27));
sram_cell_6t_5 inst_cell_27_71 (.BL(BL71),.BLN(BLN71),.WL(WL27));
sram_cell_6t_5 inst_cell_27_72 (.BL(BL72),.BLN(BLN72),.WL(WL27));
sram_cell_6t_5 inst_cell_27_73 (.BL(BL73),.BLN(BLN73),.WL(WL27));
sram_cell_6t_5 inst_cell_27_74 (.BL(BL74),.BLN(BLN74),.WL(WL27));
sram_cell_6t_5 inst_cell_27_75 (.BL(BL75),.BLN(BLN75),.WL(WL27));
sram_cell_6t_5 inst_cell_27_76 (.BL(BL76),.BLN(BLN76),.WL(WL27));
sram_cell_6t_5 inst_cell_27_77 (.BL(BL77),.BLN(BLN77),.WL(WL27));
sram_cell_6t_5 inst_cell_27_78 (.BL(BL78),.BLN(BLN78),.WL(WL27));
sram_cell_6t_5 inst_cell_27_79 (.BL(BL79),.BLN(BLN79),.WL(WL27));
sram_cell_6t_5 inst_cell_27_80 (.BL(BL80),.BLN(BLN80),.WL(WL27));
sram_cell_6t_5 inst_cell_27_81 (.BL(BL81),.BLN(BLN81),.WL(WL27));
sram_cell_6t_5 inst_cell_27_82 (.BL(BL82),.BLN(BLN82),.WL(WL27));
sram_cell_6t_5 inst_cell_27_83 (.BL(BL83),.BLN(BLN83),.WL(WL27));
sram_cell_6t_5 inst_cell_27_84 (.BL(BL84),.BLN(BLN84),.WL(WL27));
sram_cell_6t_5 inst_cell_27_85 (.BL(BL85),.BLN(BLN85),.WL(WL27));
sram_cell_6t_5 inst_cell_27_86 (.BL(BL86),.BLN(BLN86),.WL(WL27));
sram_cell_6t_5 inst_cell_27_87 (.BL(BL87),.BLN(BLN87),.WL(WL27));
sram_cell_6t_5 inst_cell_27_88 (.BL(BL88),.BLN(BLN88),.WL(WL27));
sram_cell_6t_5 inst_cell_27_89 (.BL(BL89),.BLN(BLN89),.WL(WL27));
sram_cell_6t_5 inst_cell_27_90 (.BL(BL90),.BLN(BLN90),.WL(WL27));
sram_cell_6t_5 inst_cell_27_91 (.BL(BL91),.BLN(BLN91),.WL(WL27));
sram_cell_6t_5 inst_cell_27_92 (.BL(BL92),.BLN(BLN92),.WL(WL27));
sram_cell_6t_5 inst_cell_27_93 (.BL(BL93),.BLN(BLN93),.WL(WL27));
sram_cell_6t_5 inst_cell_27_94 (.BL(BL94),.BLN(BLN94),.WL(WL27));
sram_cell_6t_5 inst_cell_27_95 (.BL(BL95),.BLN(BLN95),.WL(WL27));
sram_cell_6t_5 inst_cell_27_96 (.BL(BL96),.BLN(BLN96),.WL(WL27));
sram_cell_6t_5 inst_cell_27_97 (.BL(BL97),.BLN(BLN97),.WL(WL27));
sram_cell_6t_5 inst_cell_27_98 (.BL(BL98),.BLN(BLN98),.WL(WL27));
sram_cell_6t_5 inst_cell_27_99 (.BL(BL99),.BLN(BLN99),.WL(WL27));
sram_cell_6t_5 inst_cell_27_100 (.BL(BL100),.BLN(BLN100),.WL(WL27));
sram_cell_6t_5 inst_cell_27_101 (.BL(BL101),.BLN(BLN101),.WL(WL27));
sram_cell_6t_5 inst_cell_27_102 (.BL(BL102),.BLN(BLN102),.WL(WL27));
sram_cell_6t_5 inst_cell_27_103 (.BL(BL103),.BLN(BLN103),.WL(WL27));
sram_cell_6t_5 inst_cell_27_104 (.BL(BL104),.BLN(BLN104),.WL(WL27));
sram_cell_6t_5 inst_cell_27_105 (.BL(BL105),.BLN(BLN105),.WL(WL27));
sram_cell_6t_5 inst_cell_27_106 (.BL(BL106),.BLN(BLN106),.WL(WL27));
sram_cell_6t_5 inst_cell_27_107 (.BL(BL107),.BLN(BLN107),.WL(WL27));
sram_cell_6t_5 inst_cell_27_108 (.BL(BL108),.BLN(BLN108),.WL(WL27));
sram_cell_6t_5 inst_cell_27_109 (.BL(BL109),.BLN(BLN109),.WL(WL27));
sram_cell_6t_5 inst_cell_27_110 (.BL(BL110),.BLN(BLN110),.WL(WL27));
sram_cell_6t_5 inst_cell_27_111 (.BL(BL111),.BLN(BLN111),.WL(WL27));
sram_cell_6t_5 inst_cell_27_112 (.BL(BL112),.BLN(BLN112),.WL(WL27));
sram_cell_6t_5 inst_cell_27_113 (.BL(BL113),.BLN(BLN113),.WL(WL27));
sram_cell_6t_5 inst_cell_27_114 (.BL(BL114),.BLN(BLN114),.WL(WL27));
sram_cell_6t_5 inst_cell_27_115 (.BL(BL115),.BLN(BLN115),.WL(WL27));
sram_cell_6t_5 inst_cell_27_116 (.BL(BL116),.BLN(BLN116),.WL(WL27));
sram_cell_6t_5 inst_cell_27_117 (.BL(BL117),.BLN(BLN117),.WL(WL27));
sram_cell_6t_5 inst_cell_27_118 (.BL(BL118),.BLN(BLN118),.WL(WL27));
sram_cell_6t_5 inst_cell_27_119 (.BL(BL119),.BLN(BLN119),.WL(WL27));
sram_cell_6t_5 inst_cell_27_120 (.BL(BL120),.BLN(BLN120),.WL(WL27));
sram_cell_6t_5 inst_cell_27_121 (.BL(BL121),.BLN(BLN121),.WL(WL27));
sram_cell_6t_5 inst_cell_27_122 (.BL(BL122),.BLN(BLN122),.WL(WL27));
sram_cell_6t_5 inst_cell_27_123 (.BL(BL123),.BLN(BLN123),.WL(WL27));
sram_cell_6t_5 inst_cell_27_124 (.BL(BL124),.BLN(BLN124),.WL(WL27));
sram_cell_6t_5 inst_cell_27_125 (.BL(BL125),.BLN(BLN125),.WL(WL27));
sram_cell_6t_5 inst_cell_27_126 (.BL(BL126),.BLN(BLN126),.WL(WL27));
sram_cell_6t_5 inst_cell_27_127 (.BL(BL127),.BLN(BLN127),.WL(WL27));
sram_cell_6t_5 inst_cell_28_0 (.BL(BL0),.BLN(BLN0),.WL(WL28));
sram_cell_6t_5 inst_cell_28_1 (.BL(BL1),.BLN(BLN1),.WL(WL28));
sram_cell_6t_5 inst_cell_28_2 (.BL(BL2),.BLN(BLN2),.WL(WL28));
sram_cell_6t_5 inst_cell_28_3 (.BL(BL3),.BLN(BLN3),.WL(WL28));
sram_cell_6t_5 inst_cell_28_4 (.BL(BL4),.BLN(BLN4),.WL(WL28));
sram_cell_6t_5 inst_cell_28_5 (.BL(BL5),.BLN(BLN5),.WL(WL28));
sram_cell_6t_5 inst_cell_28_6 (.BL(BL6),.BLN(BLN6),.WL(WL28));
sram_cell_6t_5 inst_cell_28_7 (.BL(BL7),.BLN(BLN7),.WL(WL28));
sram_cell_6t_5 inst_cell_28_8 (.BL(BL8),.BLN(BLN8),.WL(WL28));
sram_cell_6t_5 inst_cell_28_9 (.BL(BL9),.BLN(BLN9),.WL(WL28));
sram_cell_6t_5 inst_cell_28_10 (.BL(BL10),.BLN(BLN10),.WL(WL28));
sram_cell_6t_5 inst_cell_28_11 (.BL(BL11),.BLN(BLN11),.WL(WL28));
sram_cell_6t_5 inst_cell_28_12 (.BL(BL12),.BLN(BLN12),.WL(WL28));
sram_cell_6t_5 inst_cell_28_13 (.BL(BL13),.BLN(BLN13),.WL(WL28));
sram_cell_6t_5 inst_cell_28_14 (.BL(BL14),.BLN(BLN14),.WL(WL28));
sram_cell_6t_5 inst_cell_28_15 (.BL(BL15),.BLN(BLN15),.WL(WL28));
sram_cell_6t_5 inst_cell_28_16 (.BL(BL16),.BLN(BLN16),.WL(WL28));
sram_cell_6t_5 inst_cell_28_17 (.BL(BL17),.BLN(BLN17),.WL(WL28));
sram_cell_6t_5 inst_cell_28_18 (.BL(BL18),.BLN(BLN18),.WL(WL28));
sram_cell_6t_5 inst_cell_28_19 (.BL(BL19),.BLN(BLN19),.WL(WL28));
sram_cell_6t_5 inst_cell_28_20 (.BL(BL20),.BLN(BLN20),.WL(WL28));
sram_cell_6t_5 inst_cell_28_21 (.BL(BL21),.BLN(BLN21),.WL(WL28));
sram_cell_6t_5 inst_cell_28_22 (.BL(BL22),.BLN(BLN22),.WL(WL28));
sram_cell_6t_5 inst_cell_28_23 (.BL(BL23),.BLN(BLN23),.WL(WL28));
sram_cell_6t_5 inst_cell_28_24 (.BL(BL24),.BLN(BLN24),.WL(WL28));
sram_cell_6t_5 inst_cell_28_25 (.BL(BL25),.BLN(BLN25),.WL(WL28));
sram_cell_6t_5 inst_cell_28_26 (.BL(BL26),.BLN(BLN26),.WL(WL28));
sram_cell_6t_5 inst_cell_28_27 (.BL(BL27),.BLN(BLN27),.WL(WL28));
sram_cell_6t_5 inst_cell_28_28 (.BL(BL28),.BLN(BLN28),.WL(WL28));
sram_cell_6t_5 inst_cell_28_29 (.BL(BL29),.BLN(BLN29),.WL(WL28));
sram_cell_6t_5 inst_cell_28_30 (.BL(BL30),.BLN(BLN30),.WL(WL28));
sram_cell_6t_5 inst_cell_28_31 (.BL(BL31),.BLN(BLN31),.WL(WL28));
sram_cell_6t_5 inst_cell_28_32 (.BL(BL32),.BLN(BLN32),.WL(WL28));
sram_cell_6t_5 inst_cell_28_33 (.BL(BL33),.BLN(BLN33),.WL(WL28));
sram_cell_6t_5 inst_cell_28_34 (.BL(BL34),.BLN(BLN34),.WL(WL28));
sram_cell_6t_5 inst_cell_28_35 (.BL(BL35),.BLN(BLN35),.WL(WL28));
sram_cell_6t_5 inst_cell_28_36 (.BL(BL36),.BLN(BLN36),.WL(WL28));
sram_cell_6t_5 inst_cell_28_37 (.BL(BL37),.BLN(BLN37),.WL(WL28));
sram_cell_6t_5 inst_cell_28_38 (.BL(BL38),.BLN(BLN38),.WL(WL28));
sram_cell_6t_5 inst_cell_28_39 (.BL(BL39),.BLN(BLN39),.WL(WL28));
sram_cell_6t_5 inst_cell_28_40 (.BL(BL40),.BLN(BLN40),.WL(WL28));
sram_cell_6t_5 inst_cell_28_41 (.BL(BL41),.BLN(BLN41),.WL(WL28));
sram_cell_6t_5 inst_cell_28_42 (.BL(BL42),.BLN(BLN42),.WL(WL28));
sram_cell_6t_5 inst_cell_28_43 (.BL(BL43),.BLN(BLN43),.WL(WL28));
sram_cell_6t_5 inst_cell_28_44 (.BL(BL44),.BLN(BLN44),.WL(WL28));
sram_cell_6t_5 inst_cell_28_45 (.BL(BL45),.BLN(BLN45),.WL(WL28));
sram_cell_6t_5 inst_cell_28_46 (.BL(BL46),.BLN(BLN46),.WL(WL28));
sram_cell_6t_5 inst_cell_28_47 (.BL(BL47),.BLN(BLN47),.WL(WL28));
sram_cell_6t_5 inst_cell_28_48 (.BL(BL48),.BLN(BLN48),.WL(WL28));
sram_cell_6t_5 inst_cell_28_49 (.BL(BL49),.BLN(BLN49),.WL(WL28));
sram_cell_6t_5 inst_cell_28_50 (.BL(BL50),.BLN(BLN50),.WL(WL28));
sram_cell_6t_5 inst_cell_28_51 (.BL(BL51),.BLN(BLN51),.WL(WL28));
sram_cell_6t_5 inst_cell_28_52 (.BL(BL52),.BLN(BLN52),.WL(WL28));
sram_cell_6t_5 inst_cell_28_53 (.BL(BL53),.BLN(BLN53),.WL(WL28));
sram_cell_6t_5 inst_cell_28_54 (.BL(BL54),.BLN(BLN54),.WL(WL28));
sram_cell_6t_5 inst_cell_28_55 (.BL(BL55),.BLN(BLN55),.WL(WL28));
sram_cell_6t_5 inst_cell_28_56 (.BL(BL56),.BLN(BLN56),.WL(WL28));
sram_cell_6t_5 inst_cell_28_57 (.BL(BL57),.BLN(BLN57),.WL(WL28));
sram_cell_6t_5 inst_cell_28_58 (.BL(BL58),.BLN(BLN58),.WL(WL28));
sram_cell_6t_5 inst_cell_28_59 (.BL(BL59),.BLN(BLN59),.WL(WL28));
sram_cell_6t_5 inst_cell_28_60 (.BL(BL60),.BLN(BLN60),.WL(WL28));
sram_cell_6t_5 inst_cell_28_61 (.BL(BL61),.BLN(BLN61),.WL(WL28));
sram_cell_6t_5 inst_cell_28_62 (.BL(BL62),.BLN(BLN62),.WL(WL28));
sram_cell_6t_5 inst_cell_28_63 (.BL(BL63),.BLN(BLN63),.WL(WL28));
sram_cell_6t_5 inst_cell_28_64 (.BL(BL64),.BLN(BLN64),.WL(WL28));
sram_cell_6t_5 inst_cell_28_65 (.BL(BL65),.BLN(BLN65),.WL(WL28));
sram_cell_6t_5 inst_cell_28_66 (.BL(BL66),.BLN(BLN66),.WL(WL28));
sram_cell_6t_5 inst_cell_28_67 (.BL(BL67),.BLN(BLN67),.WL(WL28));
sram_cell_6t_5 inst_cell_28_68 (.BL(BL68),.BLN(BLN68),.WL(WL28));
sram_cell_6t_5 inst_cell_28_69 (.BL(BL69),.BLN(BLN69),.WL(WL28));
sram_cell_6t_5 inst_cell_28_70 (.BL(BL70),.BLN(BLN70),.WL(WL28));
sram_cell_6t_5 inst_cell_28_71 (.BL(BL71),.BLN(BLN71),.WL(WL28));
sram_cell_6t_5 inst_cell_28_72 (.BL(BL72),.BLN(BLN72),.WL(WL28));
sram_cell_6t_5 inst_cell_28_73 (.BL(BL73),.BLN(BLN73),.WL(WL28));
sram_cell_6t_5 inst_cell_28_74 (.BL(BL74),.BLN(BLN74),.WL(WL28));
sram_cell_6t_5 inst_cell_28_75 (.BL(BL75),.BLN(BLN75),.WL(WL28));
sram_cell_6t_5 inst_cell_28_76 (.BL(BL76),.BLN(BLN76),.WL(WL28));
sram_cell_6t_5 inst_cell_28_77 (.BL(BL77),.BLN(BLN77),.WL(WL28));
sram_cell_6t_5 inst_cell_28_78 (.BL(BL78),.BLN(BLN78),.WL(WL28));
sram_cell_6t_5 inst_cell_28_79 (.BL(BL79),.BLN(BLN79),.WL(WL28));
sram_cell_6t_5 inst_cell_28_80 (.BL(BL80),.BLN(BLN80),.WL(WL28));
sram_cell_6t_5 inst_cell_28_81 (.BL(BL81),.BLN(BLN81),.WL(WL28));
sram_cell_6t_5 inst_cell_28_82 (.BL(BL82),.BLN(BLN82),.WL(WL28));
sram_cell_6t_5 inst_cell_28_83 (.BL(BL83),.BLN(BLN83),.WL(WL28));
sram_cell_6t_5 inst_cell_28_84 (.BL(BL84),.BLN(BLN84),.WL(WL28));
sram_cell_6t_5 inst_cell_28_85 (.BL(BL85),.BLN(BLN85),.WL(WL28));
sram_cell_6t_5 inst_cell_28_86 (.BL(BL86),.BLN(BLN86),.WL(WL28));
sram_cell_6t_5 inst_cell_28_87 (.BL(BL87),.BLN(BLN87),.WL(WL28));
sram_cell_6t_5 inst_cell_28_88 (.BL(BL88),.BLN(BLN88),.WL(WL28));
sram_cell_6t_5 inst_cell_28_89 (.BL(BL89),.BLN(BLN89),.WL(WL28));
sram_cell_6t_5 inst_cell_28_90 (.BL(BL90),.BLN(BLN90),.WL(WL28));
sram_cell_6t_5 inst_cell_28_91 (.BL(BL91),.BLN(BLN91),.WL(WL28));
sram_cell_6t_5 inst_cell_28_92 (.BL(BL92),.BLN(BLN92),.WL(WL28));
sram_cell_6t_5 inst_cell_28_93 (.BL(BL93),.BLN(BLN93),.WL(WL28));
sram_cell_6t_5 inst_cell_28_94 (.BL(BL94),.BLN(BLN94),.WL(WL28));
sram_cell_6t_5 inst_cell_28_95 (.BL(BL95),.BLN(BLN95),.WL(WL28));
sram_cell_6t_5 inst_cell_28_96 (.BL(BL96),.BLN(BLN96),.WL(WL28));
sram_cell_6t_5 inst_cell_28_97 (.BL(BL97),.BLN(BLN97),.WL(WL28));
sram_cell_6t_5 inst_cell_28_98 (.BL(BL98),.BLN(BLN98),.WL(WL28));
sram_cell_6t_5 inst_cell_28_99 (.BL(BL99),.BLN(BLN99),.WL(WL28));
sram_cell_6t_5 inst_cell_28_100 (.BL(BL100),.BLN(BLN100),.WL(WL28));
sram_cell_6t_5 inst_cell_28_101 (.BL(BL101),.BLN(BLN101),.WL(WL28));
sram_cell_6t_5 inst_cell_28_102 (.BL(BL102),.BLN(BLN102),.WL(WL28));
sram_cell_6t_5 inst_cell_28_103 (.BL(BL103),.BLN(BLN103),.WL(WL28));
sram_cell_6t_5 inst_cell_28_104 (.BL(BL104),.BLN(BLN104),.WL(WL28));
sram_cell_6t_5 inst_cell_28_105 (.BL(BL105),.BLN(BLN105),.WL(WL28));
sram_cell_6t_5 inst_cell_28_106 (.BL(BL106),.BLN(BLN106),.WL(WL28));
sram_cell_6t_5 inst_cell_28_107 (.BL(BL107),.BLN(BLN107),.WL(WL28));
sram_cell_6t_5 inst_cell_28_108 (.BL(BL108),.BLN(BLN108),.WL(WL28));
sram_cell_6t_5 inst_cell_28_109 (.BL(BL109),.BLN(BLN109),.WL(WL28));
sram_cell_6t_5 inst_cell_28_110 (.BL(BL110),.BLN(BLN110),.WL(WL28));
sram_cell_6t_5 inst_cell_28_111 (.BL(BL111),.BLN(BLN111),.WL(WL28));
sram_cell_6t_5 inst_cell_28_112 (.BL(BL112),.BLN(BLN112),.WL(WL28));
sram_cell_6t_5 inst_cell_28_113 (.BL(BL113),.BLN(BLN113),.WL(WL28));
sram_cell_6t_5 inst_cell_28_114 (.BL(BL114),.BLN(BLN114),.WL(WL28));
sram_cell_6t_5 inst_cell_28_115 (.BL(BL115),.BLN(BLN115),.WL(WL28));
sram_cell_6t_5 inst_cell_28_116 (.BL(BL116),.BLN(BLN116),.WL(WL28));
sram_cell_6t_5 inst_cell_28_117 (.BL(BL117),.BLN(BLN117),.WL(WL28));
sram_cell_6t_5 inst_cell_28_118 (.BL(BL118),.BLN(BLN118),.WL(WL28));
sram_cell_6t_5 inst_cell_28_119 (.BL(BL119),.BLN(BLN119),.WL(WL28));
sram_cell_6t_5 inst_cell_28_120 (.BL(BL120),.BLN(BLN120),.WL(WL28));
sram_cell_6t_5 inst_cell_28_121 (.BL(BL121),.BLN(BLN121),.WL(WL28));
sram_cell_6t_5 inst_cell_28_122 (.BL(BL122),.BLN(BLN122),.WL(WL28));
sram_cell_6t_5 inst_cell_28_123 (.BL(BL123),.BLN(BLN123),.WL(WL28));
sram_cell_6t_5 inst_cell_28_124 (.BL(BL124),.BLN(BLN124),.WL(WL28));
sram_cell_6t_5 inst_cell_28_125 (.BL(BL125),.BLN(BLN125),.WL(WL28));
sram_cell_6t_5 inst_cell_28_126 (.BL(BL126),.BLN(BLN126),.WL(WL28));
sram_cell_6t_5 inst_cell_28_127 (.BL(BL127),.BLN(BLN127),.WL(WL28));
sram_cell_6t_5 inst_cell_29_0 (.BL(BL0),.BLN(BLN0),.WL(WL29));
sram_cell_6t_5 inst_cell_29_1 (.BL(BL1),.BLN(BLN1),.WL(WL29));
sram_cell_6t_5 inst_cell_29_2 (.BL(BL2),.BLN(BLN2),.WL(WL29));
sram_cell_6t_5 inst_cell_29_3 (.BL(BL3),.BLN(BLN3),.WL(WL29));
sram_cell_6t_5 inst_cell_29_4 (.BL(BL4),.BLN(BLN4),.WL(WL29));
sram_cell_6t_5 inst_cell_29_5 (.BL(BL5),.BLN(BLN5),.WL(WL29));
sram_cell_6t_5 inst_cell_29_6 (.BL(BL6),.BLN(BLN6),.WL(WL29));
sram_cell_6t_5 inst_cell_29_7 (.BL(BL7),.BLN(BLN7),.WL(WL29));
sram_cell_6t_5 inst_cell_29_8 (.BL(BL8),.BLN(BLN8),.WL(WL29));
sram_cell_6t_5 inst_cell_29_9 (.BL(BL9),.BLN(BLN9),.WL(WL29));
sram_cell_6t_5 inst_cell_29_10 (.BL(BL10),.BLN(BLN10),.WL(WL29));
sram_cell_6t_5 inst_cell_29_11 (.BL(BL11),.BLN(BLN11),.WL(WL29));
sram_cell_6t_5 inst_cell_29_12 (.BL(BL12),.BLN(BLN12),.WL(WL29));
sram_cell_6t_5 inst_cell_29_13 (.BL(BL13),.BLN(BLN13),.WL(WL29));
sram_cell_6t_5 inst_cell_29_14 (.BL(BL14),.BLN(BLN14),.WL(WL29));
sram_cell_6t_5 inst_cell_29_15 (.BL(BL15),.BLN(BLN15),.WL(WL29));
sram_cell_6t_5 inst_cell_29_16 (.BL(BL16),.BLN(BLN16),.WL(WL29));
sram_cell_6t_5 inst_cell_29_17 (.BL(BL17),.BLN(BLN17),.WL(WL29));
sram_cell_6t_5 inst_cell_29_18 (.BL(BL18),.BLN(BLN18),.WL(WL29));
sram_cell_6t_5 inst_cell_29_19 (.BL(BL19),.BLN(BLN19),.WL(WL29));
sram_cell_6t_5 inst_cell_29_20 (.BL(BL20),.BLN(BLN20),.WL(WL29));
sram_cell_6t_5 inst_cell_29_21 (.BL(BL21),.BLN(BLN21),.WL(WL29));
sram_cell_6t_5 inst_cell_29_22 (.BL(BL22),.BLN(BLN22),.WL(WL29));
sram_cell_6t_5 inst_cell_29_23 (.BL(BL23),.BLN(BLN23),.WL(WL29));
sram_cell_6t_5 inst_cell_29_24 (.BL(BL24),.BLN(BLN24),.WL(WL29));
sram_cell_6t_5 inst_cell_29_25 (.BL(BL25),.BLN(BLN25),.WL(WL29));
sram_cell_6t_5 inst_cell_29_26 (.BL(BL26),.BLN(BLN26),.WL(WL29));
sram_cell_6t_5 inst_cell_29_27 (.BL(BL27),.BLN(BLN27),.WL(WL29));
sram_cell_6t_5 inst_cell_29_28 (.BL(BL28),.BLN(BLN28),.WL(WL29));
sram_cell_6t_5 inst_cell_29_29 (.BL(BL29),.BLN(BLN29),.WL(WL29));
sram_cell_6t_5 inst_cell_29_30 (.BL(BL30),.BLN(BLN30),.WL(WL29));
sram_cell_6t_5 inst_cell_29_31 (.BL(BL31),.BLN(BLN31),.WL(WL29));
sram_cell_6t_5 inst_cell_29_32 (.BL(BL32),.BLN(BLN32),.WL(WL29));
sram_cell_6t_5 inst_cell_29_33 (.BL(BL33),.BLN(BLN33),.WL(WL29));
sram_cell_6t_5 inst_cell_29_34 (.BL(BL34),.BLN(BLN34),.WL(WL29));
sram_cell_6t_5 inst_cell_29_35 (.BL(BL35),.BLN(BLN35),.WL(WL29));
sram_cell_6t_5 inst_cell_29_36 (.BL(BL36),.BLN(BLN36),.WL(WL29));
sram_cell_6t_5 inst_cell_29_37 (.BL(BL37),.BLN(BLN37),.WL(WL29));
sram_cell_6t_5 inst_cell_29_38 (.BL(BL38),.BLN(BLN38),.WL(WL29));
sram_cell_6t_5 inst_cell_29_39 (.BL(BL39),.BLN(BLN39),.WL(WL29));
sram_cell_6t_5 inst_cell_29_40 (.BL(BL40),.BLN(BLN40),.WL(WL29));
sram_cell_6t_5 inst_cell_29_41 (.BL(BL41),.BLN(BLN41),.WL(WL29));
sram_cell_6t_5 inst_cell_29_42 (.BL(BL42),.BLN(BLN42),.WL(WL29));
sram_cell_6t_5 inst_cell_29_43 (.BL(BL43),.BLN(BLN43),.WL(WL29));
sram_cell_6t_5 inst_cell_29_44 (.BL(BL44),.BLN(BLN44),.WL(WL29));
sram_cell_6t_5 inst_cell_29_45 (.BL(BL45),.BLN(BLN45),.WL(WL29));
sram_cell_6t_5 inst_cell_29_46 (.BL(BL46),.BLN(BLN46),.WL(WL29));
sram_cell_6t_5 inst_cell_29_47 (.BL(BL47),.BLN(BLN47),.WL(WL29));
sram_cell_6t_5 inst_cell_29_48 (.BL(BL48),.BLN(BLN48),.WL(WL29));
sram_cell_6t_5 inst_cell_29_49 (.BL(BL49),.BLN(BLN49),.WL(WL29));
sram_cell_6t_5 inst_cell_29_50 (.BL(BL50),.BLN(BLN50),.WL(WL29));
sram_cell_6t_5 inst_cell_29_51 (.BL(BL51),.BLN(BLN51),.WL(WL29));
sram_cell_6t_5 inst_cell_29_52 (.BL(BL52),.BLN(BLN52),.WL(WL29));
sram_cell_6t_5 inst_cell_29_53 (.BL(BL53),.BLN(BLN53),.WL(WL29));
sram_cell_6t_5 inst_cell_29_54 (.BL(BL54),.BLN(BLN54),.WL(WL29));
sram_cell_6t_5 inst_cell_29_55 (.BL(BL55),.BLN(BLN55),.WL(WL29));
sram_cell_6t_5 inst_cell_29_56 (.BL(BL56),.BLN(BLN56),.WL(WL29));
sram_cell_6t_5 inst_cell_29_57 (.BL(BL57),.BLN(BLN57),.WL(WL29));
sram_cell_6t_5 inst_cell_29_58 (.BL(BL58),.BLN(BLN58),.WL(WL29));
sram_cell_6t_5 inst_cell_29_59 (.BL(BL59),.BLN(BLN59),.WL(WL29));
sram_cell_6t_5 inst_cell_29_60 (.BL(BL60),.BLN(BLN60),.WL(WL29));
sram_cell_6t_5 inst_cell_29_61 (.BL(BL61),.BLN(BLN61),.WL(WL29));
sram_cell_6t_5 inst_cell_29_62 (.BL(BL62),.BLN(BLN62),.WL(WL29));
sram_cell_6t_5 inst_cell_29_63 (.BL(BL63),.BLN(BLN63),.WL(WL29));
sram_cell_6t_5 inst_cell_29_64 (.BL(BL64),.BLN(BLN64),.WL(WL29));
sram_cell_6t_5 inst_cell_29_65 (.BL(BL65),.BLN(BLN65),.WL(WL29));
sram_cell_6t_5 inst_cell_29_66 (.BL(BL66),.BLN(BLN66),.WL(WL29));
sram_cell_6t_5 inst_cell_29_67 (.BL(BL67),.BLN(BLN67),.WL(WL29));
sram_cell_6t_5 inst_cell_29_68 (.BL(BL68),.BLN(BLN68),.WL(WL29));
sram_cell_6t_5 inst_cell_29_69 (.BL(BL69),.BLN(BLN69),.WL(WL29));
sram_cell_6t_5 inst_cell_29_70 (.BL(BL70),.BLN(BLN70),.WL(WL29));
sram_cell_6t_5 inst_cell_29_71 (.BL(BL71),.BLN(BLN71),.WL(WL29));
sram_cell_6t_5 inst_cell_29_72 (.BL(BL72),.BLN(BLN72),.WL(WL29));
sram_cell_6t_5 inst_cell_29_73 (.BL(BL73),.BLN(BLN73),.WL(WL29));
sram_cell_6t_5 inst_cell_29_74 (.BL(BL74),.BLN(BLN74),.WL(WL29));
sram_cell_6t_5 inst_cell_29_75 (.BL(BL75),.BLN(BLN75),.WL(WL29));
sram_cell_6t_5 inst_cell_29_76 (.BL(BL76),.BLN(BLN76),.WL(WL29));
sram_cell_6t_5 inst_cell_29_77 (.BL(BL77),.BLN(BLN77),.WL(WL29));
sram_cell_6t_5 inst_cell_29_78 (.BL(BL78),.BLN(BLN78),.WL(WL29));
sram_cell_6t_5 inst_cell_29_79 (.BL(BL79),.BLN(BLN79),.WL(WL29));
sram_cell_6t_5 inst_cell_29_80 (.BL(BL80),.BLN(BLN80),.WL(WL29));
sram_cell_6t_5 inst_cell_29_81 (.BL(BL81),.BLN(BLN81),.WL(WL29));
sram_cell_6t_5 inst_cell_29_82 (.BL(BL82),.BLN(BLN82),.WL(WL29));
sram_cell_6t_5 inst_cell_29_83 (.BL(BL83),.BLN(BLN83),.WL(WL29));
sram_cell_6t_5 inst_cell_29_84 (.BL(BL84),.BLN(BLN84),.WL(WL29));
sram_cell_6t_5 inst_cell_29_85 (.BL(BL85),.BLN(BLN85),.WL(WL29));
sram_cell_6t_5 inst_cell_29_86 (.BL(BL86),.BLN(BLN86),.WL(WL29));
sram_cell_6t_5 inst_cell_29_87 (.BL(BL87),.BLN(BLN87),.WL(WL29));
sram_cell_6t_5 inst_cell_29_88 (.BL(BL88),.BLN(BLN88),.WL(WL29));
sram_cell_6t_5 inst_cell_29_89 (.BL(BL89),.BLN(BLN89),.WL(WL29));
sram_cell_6t_5 inst_cell_29_90 (.BL(BL90),.BLN(BLN90),.WL(WL29));
sram_cell_6t_5 inst_cell_29_91 (.BL(BL91),.BLN(BLN91),.WL(WL29));
sram_cell_6t_5 inst_cell_29_92 (.BL(BL92),.BLN(BLN92),.WL(WL29));
sram_cell_6t_5 inst_cell_29_93 (.BL(BL93),.BLN(BLN93),.WL(WL29));
sram_cell_6t_5 inst_cell_29_94 (.BL(BL94),.BLN(BLN94),.WL(WL29));
sram_cell_6t_5 inst_cell_29_95 (.BL(BL95),.BLN(BLN95),.WL(WL29));
sram_cell_6t_5 inst_cell_29_96 (.BL(BL96),.BLN(BLN96),.WL(WL29));
sram_cell_6t_5 inst_cell_29_97 (.BL(BL97),.BLN(BLN97),.WL(WL29));
sram_cell_6t_5 inst_cell_29_98 (.BL(BL98),.BLN(BLN98),.WL(WL29));
sram_cell_6t_5 inst_cell_29_99 (.BL(BL99),.BLN(BLN99),.WL(WL29));
sram_cell_6t_5 inst_cell_29_100 (.BL(BL100),.BLN(BLN100),.WL(WL29));
sram_cell_6t_5 inst_cell_29_101 (.BL(BL101),.BLN(BLN101),.WL(WL29));
sram_cell_6t_5 inst_cell_29_102 (.BL(BL102),.BLN(BLN102),.WL(WL29));
sram_cell_6t_5 inst_cell_29_103 (.BL(BL103),.BLN(BLN103),.WL(WL29));
sram_cell_6t_5 inst_cell_29_104 (.BL(BL104),.BLN(BLN104),.WL(WL29));
sram_cell_6t_5 inst_cell_29_105 (.BL(BL105),.BLN(BLN105),.WL(WL29));
sram_cell_6t_5 inst_cell_29_106 (.BL(BL106),.BLN(BLN106),.WL(WL29));
sram_cell_6t_5 inst_cell_29_107 (.BL(BL107),.BLN(BLN107),.WL(WL29));
sram_cell_6t_5 inst_cell_29_108 (.BL(BL108),.BLN(BLN108),.WL(WL29));
sram_cell_6t_5 inst_cell_29_109 (.BL(BL109),.BLN(BLN109),.WL(WL29));
sram_cell_6t_5 inst_cell_29_110 (.BL(BL110),.BLN(BLN110),.WL(WL29));
sram_cell_6t_5 inst_cell_29_111 (.BL(BL111),.BLN(BLN111),.WL(WL29));
sram_cell_6t_5 inst_cell_29_112 (.BL(BL112),.BLN(BLN112),.WL(WL29));
sram_cell_6t_5 inst_cell_29_113 (.BL(BL113),.BLN(BLN113),.WL(WL29));
sram_cell_6t_5 inst_cell_29_114 (.BL(BL114),.BLN(BLN114),.WL(WL29));
sram_cell_6t_5 inst_cell_29_115 (.BL(BL115),.BLN(BLN115),.WL(WL29));
sram_cell_6t_5 inst_cell_29_116 (.BL(BL116),.BLN(BLN116),.WL(WL29));
sram_cell_6t_5 inst_cell_29_117 (.BL(BL117),.BLN(BLN117),.WL(WL29));
sram_cell_6t_5 inst_cell_29_118 (.BL(BL118),.BLN(BLN118),.WL(WL29));
sram_cell_6t_5 inst_cell_29_119 (.BL(BL119),.BLN(BLN119),.WL(WL29));
sram_cell_6t_5 inst_cell_29_120 (.BL(BL120),.BLN(BLN120),.WL(WL29));
sram_cell_6t_5 inst_cell_29_121 (.BL(BL121),.BLN(BLN121),.WL(WL29));
sram_cell_6t_5 inst_cell_29_122 (.BL(BL122),.BLN(BLN122),.WL(WL29));
sram_cell_6t_5 inst_cell_29_123 (.BL(BL123),.BLN(BLN123),.WL(WL29));
sram_cell_6t_5 inst_cell_29_124 (.BL(BL124),.BLN(BLN124),.WL(WL29));
sram_cell_6t_5 inst_cell_29_125 (.BL(BL125),.BLN(BLN125),.WL(WL29));
sram_cell_6t_5 inst_cell_29_126 (.BL(BL126),.BLN(BLN126),.WL(WL29));
sram_cell_6t_5 inst_cell_29_127 (.BL(BL127),.BLN(BLN127),.WL(WL29));
sram_cell_6t_5 inst_cell_30_0 (.BL(BL0),.BLN(BLN0),.WL(WL30));
sram_cell_6t_5 inst_cell_30_1 (.BL(BL1),.BLN(BLN1),.WL(WL30));
sram_cell_6t_5 inst_cell_30_2 (.BL(BL2),.BLN(BLN2),.WL(WL30));
sram_cell_6t_5 inst_cell_30_3 (.BL(BL3),.BLN(BLN3),.WL(WL30));
sram_cell_6t_5 inst_cell_30_4 (.BL(BL4),.BLN(BLN4),.WL(WL30));
sram_cell_6t_5 inst_cell_30_5 (.BL(BL5),.BLN(BLN5),.WL(WL30));
sram_cell_6t_5 inst_cell_30_6 (.BL(BL6),.BLN(BLN6),.WL(WL30));
sram_cell_6t_5 inst_cell_30_7 (.BL(BL7),.BLN(BLN7),.WL(WL30));
sram_cell_6t_5 inst_cell_30_8 (.BL(BL8),.BLN(BLN8),.WL(WL30));
sram_cell_6t_5 inst_cell_30_9 (.BL(BL9),.BLN(BLN9),.WL(WL30));
sram_cell_6t_5 inst_cell_30_10 (.BL(BL10),.BLN(BLN10),.WL(WL30));
sram_cell_6t_5 inst_cell_30_11 (.BL(BL11),.BLN(BLN11),.WL(WL30));
sram_cell_6t_5 inst_cell_30_12 (.BL(BL12),.BLN(BLN12),.WL(WL30));
sram_cell_6t_5 inst_cell_30_13 (.BL(BL13),.BLN(BLN13),.WL(WL30));
sram_cell_6t_5 inst_cell_30_14 (.BL(BL14),.BLN(BLN14),.WL(WL30));
sram_cell_6t_5 inst_cell_30_15 (.BL(BL15),.BLN(BLN15),.WL(WL30));
sram_cell_6t_5 inst_cell_30_16 (.BL(BL16),.BLN(BLN16),.WL(WL30));
sram_cell_6t_5 inst_cell_30_17 (.BL(BL17),.BLN(BLN17),.WL(WL30));
sram_cell_6t_5 inst_cell_30_18 (.BL(BL18),.BLN(BLN18),.WL(WL30));
sram_cell_6t_5 inst_cell_30_19 (.BL(BL19),.BLN(BLN19),.WL(WL30));
sram_cell_6t_5 inst_cell_30_20 (.BL(BL20),.BLN(BLN20),.WL(WL30));
sram_cell_6t_5 inst_cell_30_21 (.BL(BL21),.BLN(BLN21),.WL(WL30));
sram_cell_6t_5 inst_cell_30_22 (.BL(BL22),.BLN(BLN22),.WL(WL30));
sram_cell_6t_5 inst_cell_30_23 (.BL(BL23),.BLN(BLN23),.WL(WL30));
sram_cell_6t_5 inst_cell_30_24 (.BL(BL24),.BLN(BLN24),.WL(WL30));
sram_cell_6t_5 inst_cell_30_25 (.BL(BL25),.BLN(BLN25),.WL(WL30));
sram_cell_6t_5 inst_cell_30_26 (.BL(BL26),.BLN(BLN26),.WL(WL30));
sram_cell_6t_5 inst_cell_30_27 (.BL(BL27),.BLN(BLN27),.WL(WL30));
sram_cell_6t_5 inst_cell_30_28 (.BL(BL28),.BLN(BLN28),.WL(WL30));
sram_cell_6t_5 inst_cell_30_29 (.BL(BL29),.BLN(BLN29),.WL(WL30));
sram_cell_6t_5 inst_cell_30_30 (.BL(BL30),.BLN(BLN30),.WL(WL30));
sram_cell_6t_5 inst_cell_30_31 (.BL(BL31),.BLN(BLN31),.WL(WL30));
sram_cell_6t_5 inst_cell_30_32 (.BL(BL32),.BLN(BLN32),.WL(WL30));
sram_cell_6t_5 inst_cell_30_33 (.BL(BL33),.BLN(BLN33),.WL(WL30));
sram_cell_6t_5 inst_cell_30_34 (.BL(BL34),.BLN(BLN34),.WL(WL30));
sram_cell_6t_5 inst_cell_30_35 (.BL(BL35),.BLN(BLN35),.WL(WL30));
sram_cell_6t_5 inst_cell_30_36 (.BL(BL36),.BLN(BLN36),.WL(WL30));
sram_cell_6t_5 inst_cell_30_37 (.BL(BL37),.BLN(BLN37),.WL(WL30));
sram_cell_6t_5 inst_cell_30_38 (.BL(BL38),.BLN(BLN38),.WL(WL30));
sram_cell_6t_5 inst_cell_30_39 (.BL(BL39),.BLN(BLN39),.WL(WL30));
sram_cell_6t_5 inst_cell_30_40 (.BL(BL40),.BLN(BLN40),.WL(WL30));
sram_cell_6t_5 inst_cell_30_41 (.BL(BL41),.BLN(BLN41),.WL(WL30));
sram_cell_6t_5 inst_cell_30_42 (.BL(BL42),.BLN(BLN42),.WL(WL30));
sram_cell_6t_5 inst_cell_30_43 (.BL(BL43),.BLN(BLN43),.WL(WL30));
sram_cell_6t_5 inst_cell_30_44 (.BL(BL44),.BLN(BLN44),.WL(WL30));
sram_cell_6t_5 inst_cell_30_45 (.BL(BL45),.BLN(BLN45),.WL(WL30));
sram_cell_6t_5 inst_cell_30_46 (.BL(BL46),.BLN(BLN46),.WL(WL30));
sram_cell_6t_5 inst_cell_30_47 (.BL(BL47),.BLN(BLN47),.WL(WL30));
sram_cell_6t_5 inst_cell_30_48 (.BL(BL48),.BLN(BLN48),.WL(WL30));
sram_cell_6t_5 inst_cell_30_49 (.BL(BL49),.BLN(BLN49),.WL(WL30));
sram_cell_6t_5 inst_cell_30_50 (.BL(BL50),.BLN(BLN50),.WL(WL30));
sram_cell_6t_5 inst_cell_30_51 (.BL(BL51),.BLN(BLN51),.WL(WL30));
sram_cell_6t_5 inst_cell_30_52 (.BL(BL52),.BLN(BLN52),.WL(WL30));
sram_cell_6t_5 inst_cell_30_53 (.BL(BL53),.BLN(BLN53),.WL(WL30));
sram_cell_6t_5 inst_cell_30_54 (.BL(BL54),.BLN(BLN54),.WL(WL30));
sram_cell_6t_5 inst_cell_30_55 (.BL(BL55),.BLN(BLN55),.WL(WL30));
sram_cell_6t_5 inst_cell_30_56 (.BL(BL56),.BLN(BLN56),.WL(WL30));
sram_cell_6t_5 inst_cell_30_57 (.BL(BL57),.BLN(BLN57),.WL(WL30));
sram_cell_6t_5 inst_cell_30_58 (.BL(BL58),.BLN(BLN58),.WL(WL30));
sram_cell_6t_5 inst_cell_30_59 (.BL(BL59),.BLN(BLN59),.WL(WL30));
sram_cell_6t_5 inst_cell_30_60 (.BL(BL60),.BLN(BLN60),.WL(WL30));
sram_cell_6t_5 inst_cell_30_61 (.BL(BL61),.BLN(BLN61),.WL(WL30));
sram_cell_6t_5 inst_cell_30_62 (.BL(BL62),.BLN(BLN62),.WL(WL30));
sram_cell_6t_5 inst_cell_30_63 (.BL(BL63),.BLN(BLN63),.WL(WL30));
sram_cell_6t_5 inst_cell_30_64 (.BL(BL64),.BLN(BLN64),.WL(WL30));
sram_cell_6t_5 inst_cell_30_65 (.BL(BL65),.BLN(BLN65),.WL(WL30));
sram_cell_6t_5 inst_cell_30_66 (.BL(BL66),.BLN(BLN66),.WL(WL30));
sram_cell_6t_5 inst_cell_30_67 (.BL(BL67),.BLN(BLN67),.WL(WL30));
sram_cell_6t_5 inst_cell_30_68 (.BL(BL68),.BLN(BLN68),.WL(WL30));
sram_cell_6t_5 inst_cell_30_69 (.BL(BL69),.BLN(BLN69),.WL(WL30));
sram_cell_6t_5 inst_cell_30_70 (.BL(BL70),.BLN(BLN70),.WL(WL30));
sram_cell_6t_5 inst_cell_30_71 (.BL(BL71),.BLN(BLN71),.WL(WL30));
sram_cell_6t_5 inst_cell_30_72 (.BL(BL72),.BLN(BLN72),.WL(WL30));
sram_cell_6t_5 inst_cell_30_73 (.BL(BL73),.BLN(BLN73),.WL(WL30));
sram_cell_6t_5 inst_cell_30_74 (.BL(BL74),.BLN(BLN74),.WL(WL30));
sram_cell_6t_5 inst_cell_30_75 (.BL(BL75),.BLN(BLN75),.WL(WL30));
sram_cell_6t_5 inst_cell_30_76 (.BL(BL76),.BLN(BLN76),.WL(WL30));
sram_cell_6t_5 inst_cell_30_77 (.BL(BL77),.BLN(BLN77),.WL(WL30));
sram_cell_6t_5 inst_cell_30_78 (.BL(BL78),.BLN(BLN78),.WL(WL30));
sram_cell_6t_5 inst_cell_30_79 (.BL(BL79),.BLN(BLN79),.WL(WL30));
sram_cell_6t_5 inst_cell_30_80 (.BL(BL80),.BLN(BLN80),.WL(WL30));
sram_cell_6t_5 inst_cell_30_81 (.BL(BL81),.BLN(BLN81),.WL(WL30));
sram_cell_6t_5 inst_cell_30_82 (.BL(BL82),.BLN(BLN82),.WL(WL30));
sram_cell_6t_5 inst_cell_30_83 (.BL(BL83),.BLN(BLN83),.WL(WL30));
sram_cell_6t_5 inst_cell_30_84 (.BL(BL84),.BLN(BLN84),.WL(WL30));
sram_cell_6t_5 inst_cell_30_85 (.BL(BL85),.BLN(BLN85),.WL(WL30));
sram_cell_6t_5 inst_cell_30_86 (.BL(BL86),.BLN(BLN86),.WL(WL30));
sram_cell_6t_5 inst_cell_30_87 (.BL(BL87),.BLN(BLN87),.WL(WL30));
sram_cell_6t_5 inst_cell_30_88 (.BL(BL88),.BLN(BLN88),.WL(WL30));
sram_cell_6t_5 inst_cell_30_89 (.BL(BL89),.BLN(BLN89),.WL(WL30));
sram_cell_6t_5 inst_cell_30_90 (.BL(BL90),.BLN(BLN90),.WL(WL30));
sram_cell_6t_5 inst_cell_30_91 (.BL(BL91),.BLN(BLN91),.WL(WL30));
sram_cell_6t_5 inst_cell_30_92 (.BL(BL92),.BLN(BLN92),.WL(WL30));
sram_cell_6t_5 inst_cell_30_93 (.BL(BL93),.BLN(BLN93),.WL(WL30));
sram_cell_6t_5 inst_cell_30_94 (.BL(BL94),.BLN(BLN94),.WL(WL30));
sram_cell_6t_5 inst_cell_30_95 (.BL(BL95),.BLN(BLN95),.WL(WL30));
sram_cell_6t_5 inst_cell_30_96 (.BL(BL96),.BLN(BLN96),.WL(WL30));
sram_cell_6t_5 inst_cell_30_97 (.BL(BL97),.BLN(BLN97),.WL(WL30));
sram_cell_6t_5 inst_cell_30_98 (.BL(BL98),.BLN(BLN98),.WL(WL30));
sram_cell_6t_5 inst_cell_30_99 (.BL(BL99),.BLN(BLN99),.WL(WL30));
sram_cell_6t_5 inst_cell_30_100 (.BL(BL100),.BLN(BLN100),.WL(WL30));
sram_cell_6t_5 inst_cell_30_101 (.BL(BL101),.BLN(BLN101),.WL(WL30));
sram_cell_6t_5 inst_cell_30_102 (.BL(BL102),.BLN(BLN102),.WL(WL30));
sram_cell_6t_5 inst_cell_30_103 (.BL(BL103),.BLN(BLN103),.WL(WL30));
sram_cell_6t_5 inst_cell_30_104 (.BL(BL104),.BLN(BLN104),.WL(WL30));
sram_cell_6t_5 inst_cell_30_105 (.BL(BL105),.BLN(BLN105),.WL(WL30));
sram_cell_6t_5 inst_cell_30_106 (.BL(BL106),.BLN(BLN106),.WL(WL30));
sram_cell_6t_5 inst_cell_30_107 (.BL(BL107),.BLN(BLN107),.WL(WL30));
sram_cell_6t_5 inst_cell_30_108 (.BL(BL108),.BLN(BLN108),.WL(WL30));
sram_cell_6t_5 inst_cell_30_109 (.BL(BL109),.BLN(BLN109),.WL(WL30));
sram_cell_6t_5 inst_cell_30_110 (.BL(BL110),.BLN(BLN110),.WL(WL30));
sram_cell_6t_5 inst_cell_30_111 (.BL(BL111),.BLN(BLN111),.WL(WL30));
sram_cell_6t_5 inst_cell_30_112 (.BL(BL112),.BLN(BLN112),.WL(WL30));
sram_cell_6t_5 inst_cell_30_113 (.BL(BL113),.BLN(BLN113),.WL(WL30));
sram_cell_6t_5 inst_cell_30_114 (.BL(BL114),.BLN(BLN114),.WL(WL30));
sram_cell_6t_5 inst_cell_30_115 (.BL(BL115),.BLN(BLN115),.WL(WL30));
sram_cell_6t_5 inst_cell_30_116 (.BL(BL116),.BLN(BLN116),.WL(WL30));
sram_cell_6t_5 inst_cell_30_117 (.BL(BL117),.BLN(BLN117),.WL(WL30));
sram_cell_6t_5 inst_cell_30_118 (.BL(BL118),.BLN(BLN118),.WL(WL30));
sram_cell_6t_5 inst_cell_30_119 (.BL(BL119),.BLN(BLN119),.WL(WL30));
sram_cell_6t_5 inst_cell_30_120 (.BL(BL120),.BLN(BLN120),.WL(WL30));
sram_cell_6t_5 inst_cell_30_121 (.BL(BL121),.BLN(BLN121),.WL(WL30));
sram_cell_6t_5 inst_cell_30_122 (.BL(BL122),.BLN(BLN122),.WL(WL30));
sram_cell_6t_5 inst_cell_30_123 (.BL(BL123),.BLN(BLN123),.WL(WL30));
sram_cell_6t_5 inst_cell_30_124 (.BL(BL124),.BLN(BLN124),.WL(WL30));
sram_cell_6t_5 inst_cell_30_125 (.BL(BL125),.BLN(BLN125),.WL(WL30));
sram_cell_6t_5 inst_cell_30_126 (.BL(BL126),.BLN(BLN126),.WL(WL30));
sram_cell_6t_5 inst_cell_30_127 (.BL(BL127),.BLN(BLN127),.WL(WL30));
sram_cell_6t_5 inst_cell_31_0 (.BL(BL0),.BLN(BLN0),.WL(WL31));
sram_cell_6t_5 inst_cell_31_1 (.BL(BL1),.BLN(BLN1),.WL(WL31));
sram_cell_6t_5 inst_cell_31_2 (.BL(BL2),.BLN(BLN2),.WL(WL31));
sram_cell_6t_5 inst_cell_31_3 (.BL(BL3),.BLN(BLN3),.WL(WL31));
sram_cell_6t_5 inst_cell_31_4 (.BL(BL4),.BLN(BLN4),.WL(WL31));
sram_cell_6t_5 inst_cell_31_5 (.BL(BL5),.BLN(BLN5),.WL(WL31));
sram_cell_6t_5 inst_cell_31_6 (.BL(BL6),.BLN(BLN6),.WL(WL31));
sram_cell_6t_5 inst_cell_31_7 (.BL(BL7),.BLN(BLN7),.WL(WL31));
sram_cell_6t_5 inst_cell_31_8 (.BL(BL8),.BLN(BLN8),.WL(WL31));
sram_cell_6t_5 inst_cell_31_9 (.BL(BL9),.BLN(BLN9),.WL(WL31));
sram_cell_6t_5 inst_cell_31_10 (.BL(BL10),.BLN(BLN10),.WL(WL31));
sram_cell_6t_5 inst_cell_31_11 (.BL(BL11),.BLN(BLN11),.WL(WL31));
sram_cell_6t_5 inst_cell_31_12 (.BL(BL12),.BLN(BLN12),.WL(WL31));
sram_cell_6t_5 inst_cell_31_13 (.BL(BL13),.BLN(BLN13),.WL(WL31));
sram_cell_6t_5 inst_cell_31_14 (.BL(BL14),.BLN(BLN14),.WL(WL31));
sram_cell_6t_5 inst_cell_31_15 (.BL(BL15),.BLN(BLN15),.WL(WL31));
sram_cell_6t_5 inst_cell_31_16 (.BL(BL16),.BLN(BLN16),.WL(WL31));
sram_cell_6t_5 inst_cell_31_17 (.BL(BL17),.BLN(BLN17),.WL(WL31));
sram_cell_6t_5 inst_cell_31_18 (.BL(BL18),.BLN(BLN18),.WL(WL31));
sram_cell_6t_5 inst_cell_31_19 (.BL(BL19),.BLN(BLN19),.WL(WL31));
sram_cell_6t_5 inst_cell_31_20 (.BL(BL20),.BLN(BLN20),.WL(WL31));
sram_cell_6t_5 inst_cell_31_21 (.BL(BL21),.BLN(BLN21),.WL(WL31));
sram_cell_6t_5 inst_cell_31_22 (.BL(BL22),.BLN(BLN22),.WL(WL31));
sram_cell_6t_5 inst_cell_31_23 (.BL(BL23),.BLN(BLN23),.WL(WL31));
sram_cell_6t_5 inst_cell_31_24 (.BL(BL24),.BLN(BLN24),.WL(WL31));
sram_cell_6t_5 inst_cell_31_25 (.BL(BL25),.BLN(BLN25),.WL(WL31));
sram_cell_6t_5 inst_cell_31_26 (.BL(BL26),.BLN(BLN26),.WL(WL31));
sram_cell_6t_5 inst_cell_31_27 (.BL(BL27),.BLN(BLN27),.WL(WL31));
sram_cell_6t_5 inst_cell_31_28 (.BL(BL28),.BLN(BLN28),.WL(WL31));
sram_cell_6t_5 inst_cell_31_29 (.BL(BL29),.BLN(BLN29),.WL(WL31));
sram_cell_6t_5 inst_cell_31_30 (.BL(BL30),.BLN(BLN30),.WL(WL31));
sram_cell_6t_5 inst_cell_31_31 (.BL(BL31),.BLN(BLN31),.WL(WL31));
sram_cell_6t_5 inst_cell_31_32 (.BL(BL32),.BLN(BLN32),.WL(WL31));
sram_cell_6t_5 inst_cell_31_33 (.BL(BL33),.BLN(BLN33),.WL(WL31));
sram_cell_6t_5 inst_cell_31_34 (.BL(BL34),.BLN(BLN34),.WL(WL31));
sram_cell_6t_5 inst_cell_31_35 (.BL(BL35),.BLN(BLN35),.WL(WL31));
sram_cell_6t_5 inst_cell_31_36 (.BL(BL36),.BLN(BLN36),.WL(WL31));
sram_cell_6t_5 inst_cell_31_37 (.BL(BL37),.BLN(BLN37),.WL(WL31));
sram_cell_6t_5 inst_cell_31_38 (.BL(BL38),.BLN(BLN38),.WL(WL31));
sram_cell_6t_5 inst_cell_31_39 (.BL(BL39),.BLN(BLN39),.WL(WL31));
sram_cell_6t_5 inst_cell_31_40 (.BL(BL40),.BLN(BLN40),.WL(WL31));
sram_cell_6t_5 inst_cell_31_41 (.BL(BL41),.BLN(BLN41),.WL(WL31));
sram_cell_6t_5 inst_cell_31_42 (.BL(BL42),.BLN(BLN42),.WL(WL31));
sram_cell_6t_5 inst_cell_31_43 (.BL(BL43),.BLN(BLN43),.WL(WL31));
sram_cell_6t_5 inst_cell_31_44 (.BL(BL44),.BLN(BLN44),.WL(WL31));
sram_cell_6t_5 inst_cell_31_45 (.BL(BL45),.BLN(BLN45),.WL(WL31));
sram_cell_6t_5 inst_cell_31_46 (.BL(BL46),.BLN(BLN46),.WL(WL31));
sram_cell_6t_5 inst_cell_31_47 (.BL(BL47),.BLN(BLN47),.WL(WL31));
sram_cell_6t_5 inst_cell_31_48 (.BL(BL48),.BLN(BLN48),.WL(WL31));
sram_cell_6t_5 inst_cell_31_49 (.BL(BL49),.BLN(BLN49),.WL(WL31));
sram_cell_6t_5 inst_cell_31_50 (.BL(BL50),.BLN(BLN50),.WL(WL31));
sram_cell_6t_5 inst_cell_31_51 (.BL(BL51),.BLN(BLN51),.WL(WL31));
sram_cell_6t_5 inst_cell_31_52 (.BL(BL52),.BLN(BLN52),.WL(WL31));
sram_cell_6t_5 inst_cell_31_53 (.BL(BL53),.BLN(BLN53),.WL(WL31));
sram_cell_6t_5 inst_cell_31_54 (.BL(BL54),.BLN(BLN54),.WL(WL31));
sram_cell_6t_5 inst_cell_31_55 (.BL(BL55),.BLN(BLN55),.WL(WL31));
sram_cell_6t_5 inst_cell_31_56 (.BL(BL56),.BLN(BLN56),.WL(WL31));
sram_cell_6t_5 inst_cell_31_57 (.BL(BL57),.BLN(BLN57),.WL(WL31));
sram_cell_6t_5 inst_cell_31_58 (.BL(BL58),.BLN(BLN58),.WL(WL31));
sram_cell_6t_5 inst_cell_31_59 (.BL(BL59),.BLN(BLN59),.WL(WL31));
sram_cell_6t_5 inst_cell_31_60 (.BL(BL60),.BLN(BLN60),.WL(WL31));
sram_cell_6t_5 inst_cell_31_61 (.BL(BL61),.BLN(BLN61),.WL(WL31));
sram_cell_6t_5 inst_cell_31_62 (.BL(BL62),.BLN(BLN62),.WL(WL31));
sram_cell_6t_5 inst_cell_31_63 (.BL(BL63),.BLN(BLN63),.WL(WL31));
sram_cell_6t_5 inst_cell_31_64 (.BL(BL64),.BLN(BLN64),.WL(WL31));
sram_cell_6t_5 inst_cell_31_65 (.BL(BL65),.BLN(BLN65),.WL(WL31));
sram_cell_6t_5 inst_cell_31_66 (.BL(BL66),.BLN(BLN66),.WL(WL31));
sram_cell_6t_5 inst_cell_31_67 (.BL(BL67),.BLN(BLN67),.WL(WL31));
sram_cell_6t_5 inst_cell_31_68 (.BL(BL68),.BLN(BLN68),.WL(WL31));
sram_cell_6t_5 inst_cell_31_69 (.BL(BL69),.BLN(BLN69),.WL(WL31));
sram_cell_6t_5 inst_cell_31_70 (.BL(BL70),.BLN(BLN70),.WL(WL31));
sram_cell_6t_5 inst_cell_31_71 (.BL(BL71),.BLN(BLN71),.WL(WL31));
sram_cell_6t_5 inst_cell_31_72 (.BL(BL72),.BLN(BLN72),.WL(WL31));
sram_cell_6t_5 inst_cell_31_73 (.BL(BL73),.BLN(BLN73),.WL(WL31));
sram_cell_6t_5 inst_cell_31_74 (.BL(BL74),.BLN(BLN74),.WL(WL31));
sram_cell_6t_5 inst_cell_31_75 (.BL(BL75),.BLN(BLN75),.WL(WL31));
sram_cell_6t_5 inst_cell_31_76 (.BL(BL76),.BLN(BLN76),.WL(WL31));
sram_cell_6t_5 inst_cell_31_77 (.BL(BL77),.BLN(BLN77),.WL(WL31));
sram_cell_6t_5 inst_cell_31_78 (.BL(BL78),.BLN(BLN78),.WL(WL31));
sram_cell_6t_5 inst_cell_31_79 (.BL(BL79),.BLN(BLN79),.WL(WL31));
sram_cell_6t_5 inst_cell_31_80 (.BL(BL80),.BLN(BLN80),.WL(WL31));
sram_cell_6t_5 inst_cell_31_81 (.BL(BL81),.BLN(BLN81),.WL(WL31));
sram_cell_6t_5 inst_cell_31_82 (.BL(BL82),.BLN(BLN82),.WL(WL31));
sram_cell_6t_5 inst_cell_31_83 (.BL(BL83),.BLN(BLN83),.WL(WL31));
sram_cell_6t_5 inst_cell_31_84 (.BL(BL84),.BLN(BLN84),.WL(WL31));
sram_cell_6t_5 inst_cell_31_85 (.BL(BL85),.BLN(BLN85),.WL(WL31));
sram_cell_6t_5 inst_cell_31_86 (.BL(BL86),.BLN(BLN86),.WL(WL31));
sram_cell_6t_5 inst_cell_31_87 (.BL(BL87),.BLN(BLN87),.WL(WL31));
sram_cell_6t_5 inst_cell_31_88 (.BL(BL88),.BLN(BLN88),.WL(WL31));
sram_cell_6t_5 inst_cell_31_89 (.BL(BL89),.BLN(BLN89),.WL(WL31));
sram_cell_6t_5 inst_cell_31_90 (.BL(BL90),.BLN(BLN90),.WL(WL31));
sram_cell_6t_5 inst_cell_31_91 (.BL(BL91),.BLN(BLN91),.WL(WL31));
sram_cell_6t_5 inst_cell_31_92 (.BL(BL92),.BLN(BLN92),.WL(WL31));
sram_cell_6t_5 inst_cell_31_93 (.BL(BL93),.BLN(BLN93),.WL(WL31));
sram_cell_6t_5 inst_cell_31_94 (.BL(BL94),.BLN(BLN94),.WL(WL31));
sram_cell_6t_5 inst_cell_31_95 (.BL(BL95),.BLN(BLN95),.WL(WL31));
sram_cell_6t_5 inst_cell_31_96 (.BL(BL96),.BLN(BLN96),.WL(WL31));
sram_cell_6t_5 inst_cell_31_97 (.BL(BL97),.BLN(BLN97),.WL(WL31));
sram_cell_6t_5 inst_cell_31_98 (.BL(BL98),.BLN(BLN98),.WL(WL31));
sram_cell_6t_5 inst_cell_31_99 (.BL(BL99),.BLN(BLN99),.WL(WL31));
sram_cell_6t_5 inst_cell_31_100 (.BL(BL100),.BLN(BLN100),.WL(WL31));
sram_cell_6t_5 inst_cell_31_101 (.BL(BL101),.BLN(BLN101),.WL(WL31));
sram_cell_6t_5 inst_cell_31_102 (.BL(BL102),.BLN(BLN102),.WL(WL31));
sram_cell_6t_5 inst_cell_31_103 (.BL(BL103),.BLN(BLN103),.WL(WL31));
sram_cell_6t_5 inst_cell_31_104 (.BL(BL104),.BLN(BLN104),.WL(WL31));
sram_cell_6t_5 inst_cell_31_105 (.BL(BL105),.BLN(BLN105),.WL(WL31));
sram_cell_6t_5 inst_cell_31_106 (.BL(BL106),.BLN(BLN106),.WL(WL31));
sram_cell_6t_5 inst_cell_31_107 (.BL(BL107),.BLN(BLN107),.WL(WL31));
sram_cell_6t_5 inst_cell_31_108 (.BL(BL108),.BLN(BLN108),.WL(WL31));
sram_cell_6t_5 inst_cell_31_109 (.BL(BL109),.BLN(BLN109),.WL(WL31));
sram_cell_6t_5 inst_cell_31_110 (.BL(BL110),.BLN(BLN110),.WL(WL31));
sram_cell_6t_5 inst_cell_31_111 (.BL(BL111),.BLN(BLN111),.WL(WL31));
sram_cell_6t_5 inst_cell_31_112 (.BL(BL112),.BLN(BLN112),.WL(WL31));
sram_cell_6t_5 inst_cell_31_113 (.BL(BL113),.BLN(BLN113),.WL(WL31));
sram_cell_6t_5 inst_cell_31_114 (.BL(BL114),.BLN(BLN114),.WL(WL31));
sram_cell_6t_5 inst_cell_31_115 (.BL(BL115),.BLN(BLN115),.WL(WL31));
sram_cell_6t_5 inst_cell_31_116 (.BL(BL116),.BLN(BLN116),.WL(WL31));
sram_cell_6t_5 inst_cell_31_117 (.BL(BL117),.BLN(BLN117),.WL(WL31));
sram_cell_6t_5 inst_cell_31_118 (.BL(BL118),.BLN(BLN118),.WL(WL31));
sram_cell_6t_5 inst_cell_31_119 (.BL(BL119),.BLN(BLN119),.WL(WL31));
sram_cell_6t_5 inst_cell_31_120 (.BL(BL120),.BLN(BLN120),.WL(WL31));
sram_cell_6t_5 inst_cell_31_121 (.BL(BL121),.BLN(BLN121),.WL(WL31));
sram_cell_6t_5 inst_cell_31_122 (.BL(BL122),.BLN(BLN122),.WL(WL31));
sram_cell_6t_5 inst_cell_31_123 (.BL(BL123),.BLN(BLN123),.WL(WL31));
sram_cell_6t_5 inst_cell_31_124 (.BL(BL124),.BLN(BLN124),.WL(WL31));
sram_cell_6t_5 inst_cell_31_125 (.BL(BL125),.BLN(BLN125),.WL(WL31));
sram_cell_6t_5 inst_cell_31_126 (.BL(BL126),.BLN(BLN126),.WL(WL31));
sram_cell_6t_5 inst_cell_31_127 (.BL(BL127),.BLN(BLN127),.WL(WL31));
sram_cell_6t_5 inst_cell_32_0 (.BL(BL0),.BLN(BLN0),.WL(WL32));
sram_cell_6t_5 inst_cell_32_1 (.BL(BL1),.BLN(BLN1),.WL(WL32));
sram_cell_6t_5 inst_cell_32_2 (.BL(BL2),.BLN(BLN2),.WL(WL32));
sram_cell_6t_5 inst_cell_32_3 (.BL(BL3),.BLN(BLN3),.WL(WL32));
sram_cell_6t_5 inst_cell_32_4 (.BL(BL4),.BLN(BLN4),.WL(WL32));
sram_cell_6t_5 inst_cell_32_5 (.BL(BL5),.BLN(BLN5),.WL(WL32));
sram_cell_6t_5 inst_cell_32_6 (.BL(BL6),.BLN(BLN6),.WL(WL32));
sram_cell_6t_5 inst_cell_32_7 (.BL(BL7),.BLN(BLN7),.WL(WL32));
sram_cell_6t_5 inst_cell_32_8 (.BL(BL8),.BLN(BLN8),.WL(WL32));
sram_cell_6t_5 inst_cell_32_9 (.BL(BL9),.BLN(BLN9),.WL(WL32));
sram_cell_6t_5 inst_cell_32_10 (.BL(BL10),.BLN(BLN10),.WL(WL32));
sram_cell_6t_5 inst_cell_32_11 (.BL(BL11),.BLN(BLN11),.WL(WL32));
sram_cell_6t_5 inst_cell_32_12 (.BL(BL12),.BLN(BLN12),.WL(WL32));
sram_cell_6t_5 inst_cell_32_13 (.BL(BL13),.BLN(BLN13),.WL(WL32));
sram_cell_6t_5 inst_cell_32_14 (.BL(BL14),.BLN(BLN14),.WL(WL32));
sram_cell_6t_5 inst_cell_32_15 (.BL(BL15),.BLN(BLN15),.WL(WL32));
sram_cell_6t_5 inst_cell_32_16 (.BL(BL16),.BLN(BLN16),.WL(WL32));
sram_cell_6t_5 inst_cell_32_17 (.BL(BL17),.BLN(BLN17),.WL(WL32));
sram_cell_6t_5 inst_cell_32_18 (.BL(BL18),.BLN(BLN18),.WL(WL32));
sram_cell_6t_5 inst_cell_32_19 (.BL(BL19),.BLN(BLN19),.WL(WL32));
sram_cell_6t_5 inst_cell_32_20 (.BL(BL20),.BLN(BLN20),.WL(WL32));
sram_cell_6t_5 inst_cell_32_21 (.BL(BL21),.BLN(BLN21),.WL(WL32));
sram_cell_6t_5 inst_cell_32_22 (.BL(BL22),.BLN(BLN22),.WL(WL32));
sram_cell_6t_5 inst_cell_32_23 (.BL(BL23),.BLN(BLN23),.WL(WL32));
sram_cell_6t_5 inst_cell_32_24 (.BL(BL24),.BLN(BLN24),.WL(WL32));
sram_cell_6t_5 inst_cell_32_25 (.BL(BL25),.BLN(BLN25),.WL(WL32));
sram_cell_6t_5 inst_cell_32_26 (.BL(BL26),.BLN(BLN26),.WL(WL32));
sram_cell_6t_5 inst_cell_32_27 (.BL(BL27),.BLN(BLN27),.WL(WL32));
sram_cell_6t_5 inst_cell_32_28 (.BL(BL28),.BLN(BLN28),.WL(WL32));
sram_cell_6t_5 inst_cell_32_29 (.BL(BL29),.BLN(BLN29),.WL(WL32));
sram_cell_6t_5 inst_cell_32_30 (.BL(BL30),.BLN(BLN30),.WL(WL32));
sram_cell_6t_5 inst_cell_32_31 (.BL(BL31),.BLN(BLN31),.WL(WL32));
sram_cell_6t_5 inst_cell_32_32 (.BL(BL32),.BLN(BLN32),.WL(WL32));
sram_cell_6t_5 inst_cell_32_33 (.BL(BL33),.BLN(BLN33),.WL(WL32));
sram_cell_6t_5 inst_cell_32_34 (.BL(BL34),.BLN(BLN34),.WL(WL32));
sram_cell_6t_5 inst_cell_32_35 (.BL(BL35),.BLN(BLN35),.WL(WL32));
sram_cell_6t_5 inst_cell_32_36 (.BL(BL36),.BLN(BLN36),.WL(WL32));
sram_cell_6t_5 inst_cell_32_37 (.BL(BL37),.BLN(BLN37),.WL(WL32));
sram_cell_6t_5 inst_cell_32_38 (.BL(BL38),.BLN(BLN38),.WL(WL32));
sram_cell_6t_5 inst_cell_32_39 (.BL(BL39),.BLN(BLN39),.WL(WL32));
sram_cell_6t_5 inst_cell_32_40 (.BL(BL40),.BLN(BLN40),.WL(WL32));
sram_cell_6t_5 inst_cell_32_41 (.BL(BL41),.BLN(BLN41),.WL(WL32));
sram_cell_6t_5 inst_cell_32_42 (.BL(BL42),.BLN(BLN42),.WL(WL32));
sram_cell_6t_5 inst_cell_32_43 (.BL(BL43),.BLN(BLN43),.WL(WL32));
sram_cell_6t_5 inst_cell_32_44 (.BL(BL44),.BLN(BLN44),.WL(WL32));
sram_cell_6t_5 inst_cell_32_45 (.BL(BL45),.BLN(BLN45),.WL(WL32));
sram_cell_6t_5 inst_cell_32_46 (.BL(BL46),.BLN(BLN46),.WL(WL32));
sram_cell_6t_5 inst_cell_32_47 (.BL(BL47),.BLN(BLN47),.WL(WL32));
sram_cell_6t_5 inst_cell_32_48 (.BL(BL48),.BLN(BLN48),.WL(WL32));
sram_cell_6t_5 inst_cell_32_49 (.BL(BL49),.BLN(BLN49),.WL(WL32));
sram_cell_6t_5 inst_cell_32_50 (.BL(BL50),.BLN(BLN50),.WL(WL32));
sram_cell_6t_5 inst_cell_32_51 (.BL(BL51),.BLN(BLN51),.WL(WL32));
sram_cell_6t_5 inst_cell_32_52 (.BL(BL52),.BLN(BLN52),.WL(WL32));
sram_cell_6t_5 inst_cell_32_53 (.BL(BL53),.BLN(BLN53),.WL(WL32));
sram_cell_6t_5 inst_cell_32_54 (.BL(BL54),.BLN(BLN54),.WL(WL32));
sram_cell_6t_5 inst_cell_32_55 (.BL(BL55),.BLN(BLN55),.WL(WL32));
sram_cell_6t_5 inst_cell_32_56 (.BL(BL56),.BLN(BLN56),.WL(WL32));
sram_cell_6t_5 inst_cell_32_57 (.BL(BL57),.BLN(BLN57),.WL(WL32));
sram_cell_6t_5 inst_cell_32_58 (.BL(BL58),.BLN(BLN58),.WL(WL32));
sram_cell_6t_5 inst_cell_32_59 (.BL(BL59),.BLN(BLN59),.WL(WL32));
sram_cell_6t_5 inst_cell_32_60 (.BL(BL60),.BLN(BLN60),.WL(WL32));
sram_cell_6t_5 inst_cell_32_61 (.BL(BL61),.BLN(BLN61),.WL(WL32));
sram_cell_6t_5 inst_cell_32_62 (.BL(BL62),.BLN(BLN62),.WL(WL32));
sram_cell_6t_5 inst_cell_32_63 (.BL(BL63),.BLN(BLN63),.WL(WL32));
sram_cell_6t_5 inst_cell_32_64 (.BL(BL64),.BLN(BLN64),.WL(WL32));
sram_cell_6t_5 inst_cell_32_65 (.BL(BL65),.BLN(BLN65),.WL(WL32));
sram_cell_6t_5 inst_cell_32_66 (.BL(BL66),.BLN(BLN66),.WL(WL32));
sram_cell_6t_5 inst_cell_32_67 (.BL(BL67),.BLN(BLN67),.WL(WL32));
sram_cell_6t_5 inst_cell_32_68 (.BL(BL68),.BLN(BLN68),.WL(WL32));
sram_cell_6t_5 inst_cell_32_69 (.BL(BL69),.BLN(BLN69),.WL(WL32));
sram_cell_6t_5 inst_cell_32_70 (.BL(BL70),.BLN(BLN70),.WL(WL32));
sram_cell_6t_5 inst_cell_32_71 (.BL(BL71),.BLN(BLN71),.WL(WL32));
sram_cell_6t_5 inst_cell_32_72 (.BL(BL72),.BLN(BLN72),.WL(WL32));
sram_cell_6t_5 inst_cell_32_73 (.BL(BL73),.BLN(BLN73),.WL(WL32));
sram_cell_6t_5 inst_cell_32_74 (.BL(BL74),.BLN(BLN74),.WL(WL32));
sram_cell_6t_5 inst_cell_32_75 (.BL(BL75),.BLN(BLN75),.WL(WL32));
sram_cell_6t_5 inst_cell_32_76 (.BL(BL76),.BLN(BLN76),.WL(WL32));
sram_cell_6t_5 inst_cell_32_77 (.BL(BL77),.BLN(BLN77),.WL(WL32));
sram_cell_6t_5 inst_cell_32_78 (.BL(BL78),.BLN(BLN78),.WL(WL32));
sram_cell_6t_5 inst_cell_32_79 (.BL(BL79),.BLN(BLN79),.WL(WL32));
sram_cell_6t_5 inst_cell_32_80 (.BL(BL80),.BLN(BLN80),.WL(WL32));
sram_cell_6t_5 inst_cell_32_81 (.BL(BL81),.BLN(BLN81),.WL(WL32));
sram_cell_6t_5 inst_cell_32_82 (.BL(BL82),.BLN(BLN82),.WL(WL32));
sram_cell_6t_5 inst_cell_32_83 (.BL(BL83),.BLN(BLN83),.WL(WL32));
sram_cell_6t_5 inst_cell_32_84 (.BL(BL84),.BLN(BLN84),.WL(WL32));
sram_cell_6t_5 inst_cell_32_85 (.BL(BL85),.BLN(BLN85),.WL(WL32));
sram_cell_6t_5 inst_cell_32_86 (.BL(BL86),.BLN(BLN86),.WL(WL32));
sram_cell_6t_5 inst_cell_32_87 (.BL(BL87),.BLN(BLN87),.WL(WL32));
sram_cell_6t_5 inst_cell_32_88 (.BL(BL88),.BLN(BLN88),.WL(WL32));
sram_cell_6t_5 inst_cell_32_89 (.BL(BL89),.BLN(BLN89),.WL(WL32));
sram_cell_6t_5 inst_cell_32_90 (.BL(BL90),.BLN(BLN90),.WL(WL32));
sram_cell_6t_5 inst_cell_32_91 (.BL(BL91),.BLN(BLN91),.WL(WL32));
sram_cell_6t_5 inst_cell_32_92 (.BL(BL92),.BLN(BLN92),.WL(WL32));
sram_cell_6t_5 inst_cell_32_93 (.BL(BL93),.BLN(BLN93),.WL(WL32));
sram_cell_6t_5 inst_cell_32_94 (.BL(BL94),.BLN(BLN94),.WL(WL32));
sram_cell_6t_5 inst_cell_32_95 (.BL(BL95),.BLN(BLN95),.WL(WL32));
sram_cell_6t_5 inst_cell_32_96 (.BL(BL96),.BLN(BLN96),.WL(WL32));
sram_cell_6t_5 inst_cell_32_97 (.BL(BL97),.BLN(BLN97),.WL(WL32));
sram_cell_6t_5 inst_cell_32_98 (.BL(BL98),.BLN(BLN98),.WL(WL32));
sram_cell_6t_5 inst_cell_32_99 (.BL(BL99),.BLN(BLN99),.WL(WL32));
sram_cell_6t_5 inst_cell_32_100 (.BL(BL100),.BLN(BLN100),.WL(WL32));
sram_cell_6t_5 inst_cell_32_101 (.BL(BL101),.BLN(BLN101),.WL(WL32));
sram_cell_6t_5 inst_cell_32_102 (.BL(BL102),.BLN(BLN102),.WL(WL32));
sram_cell_6t_5 inst_cell_32_103 (.BL(BL103),.BLN(BLN103),.WL(WL32));
sram_cell_6t_5 inst_cell_32_104 (.BL(BL104),.BLN(BLN104),.WL(WL32));
sram_cell_6t_5 inst_cell_32_105 (.BL(BL105),.BLN(BLN105),.WL(WL32));
sram_cell_6t_5 inst_cell_32_106 (.BL(BL106),.BLN(BLN106),.WL(WL32));
sram_cell_6t_5 inst_cell_32_107 (.BL(BL107),.BLN(BLN107),.WL(WL32));
sram_cell_6t_5 inst_cell_32_108 (.BL(BL108),.BLN(BLN108),.WL(WL32));
sram_cell_6t_5 inst_cell_32_109 (.BL(BL109),.BLN(BLN109),.WL(WL32));
sram_cell_6t_5 inst_cell_32_110 (.BL(BL110),.BLN(BLN110),.WL(WL32));
sram_cell_6t_5 inst_cell_32_111 (.BL(BL111),.BLN(BLN111),.WL(WL32));
sram_cell_6t_5 inst_cell_32_112 (.BL(BL112),.BLN(BLN112),.WL(WL32));
sram_cell_6t_5 inst_cell_32_113 (.BL(BL113),.BLN(BLN113),.WL(WL32));
sram_cell_6t_5 inst_cell_32_114 (.BL(BL114),.BLN(BLN114),.WL(WL32));
sram_cell_6t_5 inst_cell_32_115 (.BL(BL115),.BLN(BLN115),.WL(WL32));
sram_cell_6t_5 inst_cell_32_116 (.BL(BL116),.BLN(BLN116),.WL(WL32));
sram_cell_6t_5 inst_cell_32_117 (.BL(BL117),.BLN(BLN117),.WL(WL32));
sram_cell_6t_5 inst_cell_32_118 (.BL(BL118),.BLN(BLN118),.WL(WL32));
sram_cell_6t_5 inst_cell_32_119 (.BL(BL119),.BLN(BLN119),.WL(WL32));
sram_cell_6t_5 inst_cell_32_120 (.BL(BL120),.BLN(BLN120),.WL(WL32));
sram_cell_6t_5 inst_cell_32_121 (.BL(BL121),.BLN(BLN121),.WL(WL32));
sram_cell_6t_5 inst_cell_32_122 (.BL(BL122),.BLN(BLN122),.WL(WL32));
sram_cell_6t_5 inst_cell_32_123 (.BL(BL123),.BLN(BLN123),.WL(WL32));
sram_cell_6t_5 inst_cell_32_124 (.BL(BL124),.BLN(BLN124),.WL(WL32));
sram_cell_6t_5 inst_cell_32_125 (.BL(BL125),.BLN(BLN125),.WL(WL32));
sram_cell_6t_5 inst_cell_32_126 (.BL(BL126),.BLN(BLN126),.WL(WL32));
sram_cell_6t_5 inst_cell_32_127 (.BL(BL127),.BLN(BLN127),.WL(WL32));
sram_cell_6t_5 inst_cell_33_0 (.BL(BL0),.BLN(BLN0),.WL(WL33));
sram_cell_6t_5 inst_cell_33_1 (.BL(BL1),.BLN(BLN1),.WL(WL33));
sram_cell_6t_5 inst_cell_33_2 (.BL(BL2),.BLN(BLN2),.WL(WL33));
sram_cell_6t_5 inst_cell_33_3 (.BL(BL3),.BLN(BLN3),.WL(WL33));
sram_cell_6t_5 inst_cell_33_4 (.BL(BL4),.BLN(BLN4),.WL(WL33));
sram_cell_6t_5 inst_cell_33_5 (.BL(BL5),.BLN(BLN5),.WL(WL33));
sram_cell_6t_5 inst_cell_33_6 (.BL(BL6),.BLN(BLN6),.WL(WL33));
sram_cell_6t_5 inst_cell_33_7 (.BL(BL7),.BLN(BLN7),.WL(WL33));
sram_cell_6t_5 inst_cell_33_8 (.BL(BL8),.BLN(BLN8),.WL(WL33));
sram_cell_6t_5 inst_cell_33_9 (.BL(BL9),.BLN(BLN9),.WL(WL33));
sram_cell_6t_5 inst_cell_33_10 (.BL(BL10),.BLN(BLN10),.WL(WL33));
sram_cell_6t_5 inst_cell_33_11 (.BL(BL11),.BLN(BLN11),.WL(WL33));
sram_cell_6t_5 inst_cell_33_12 (.BL(BL12),.BLN(BLN12),.WL(WL33));
sram_cell_6t_5 inst_cell_33_13 (.BL(BL13),.BLN(BLN13),.WL(WL33));
sram_cell_6t_5 inst_cell_33_14 (.BL(BL14),.BLN(BLN14),.WL(WL33));
sram_cell_6t_5 inst_cell_33_15 (.BL(BL15),.BLN(BLN15),.WL(WL33));
sram_cell_6t_5 inst_cell_33_16 (.BL(BL16),.BLN(BLN16),.WL(WL33));
sram_cell_6t_5 inst_cell_33_17 (.BL(BL17),.BLN(BLN17),.WL(WL33));
sram_cell_6t_5 inst_cell_33_18 (.BL(BL18),.BLN(BLN18),.WL(WL33));
sram_cell_6t_5 inst_cell_33_19 (.BL(BL19),.BLN(BLN19),.WL(WL33));
sram_cell_6t_5 inst_cell_33_20 (.BL(BL20),.BLN(BLN20),.WL(WL33));
sram_cell_6t_5 inst_cell_33_21 (.BL(BL21),.BLN(BLN21),.WL(WL33));
sram_cell_6t_5 inst_cell_33_22 (.BL(BL22),.BLN(BLN22),.WL(WL33));
sram_cell_6t_5 inst_cell_33_23 (.BL(BL23),.BLN(BLN23),.WL(WL33));
sram_cell_6t_5 inst_cell_33_24 (.BL(BL24),.BLN(BLN24),.WL(WL33));
sram_cell_6t_5 inst_cell_33_25 (.BL(BL25),.BLN(BLN25),.WL(WL33));
sram_cell_6t_5 inst_cell_33_26 (.BL(BL26),.BLN(BLN26),.WL(WL33));
sram_cell_6t_5 inst_cell_33_27 (.BL(BL27),.BLN(BLN27),.WL(WL33));
sram_cell_6t_5 inst_cell_33_28 (.BL(BL28),.BLN(BLN28),.WL(WL33));
sram_cell_6t_5 inst_cell_33_29 (.BL(BL29),.BLN(BLN29),.WL(WL33));
sram_cell_6t_5 inst_cell_33_30 (.BL(BL30),.BLN(BLN30),.WL(WL33));
sram_cell_6t_5 inst_cell_33_31 (.BL(BL31),.BLN(BLN31),.WL(WL33));
sram_cell_6t_5 inst_cell_33_32 (.BL(BL32),.BLN(BLN32),.WL(WL33));
sram_cell_6t_5 inst_cell_33_33 (.BL(BL33),.BLN(BLN33),.WL(WL33));
sram_cell_6t_5 inst_cell_33_34 (.BL(BL34),.BLN(BLN34),.WL(WL33));
sram_cell_6t_5 inst_cell_33_35 (.BL(BL35),.BLN(BLN35),.WL(WL33));
sram_cell_6t_5 inst_cell_33_36 (.BL(BL36),.BLN(BLN36),.WL(WL33));
sram_cell_6t_5 inst_cell_33_37 (.BL(BL37),.BLN(BLN37),.WL(WL33));
sram_cell_6t_5 inst_cell_33_38 (.BL(BL38),.BLN(BLN38),.WL(WL33));
sram_cell_6t_5 inst_cell_33_39 (.BL(BL39),.BLN(BLN39),.WL(WL33));
sram_cell_6t_5 inst_cell_33_40 (.BL(BL40),.BLN(BLN40),.WL(WL33));
sram_cell_6t_5 inst_cell_33_41 (.BL(BL41),.BLN(BLN41),.WL(WL33));
sram_cell_6t_5 inst_cell_33_42 (.BL(BL42),.BLN(BLN42),.WL(WL33));
sram_cell_6t_5 inst_cell_33_43 (.BL(BL43),.BLN(BLN43),.WL(WL33));
sram_cell_6t_5 inst_cell_33_44 (.BL(BL44),.BLN(BLN44),.WL(WL33));
sram_cell_6t_5 inst_cell_33_45 (.BL(BL45),.BLN(BLN45),.WL(WL33));
sram_cell_6t_5 inst_cell_33_46 (.BL(BL46),.BLN(BLN46),.WL(WL33));
sram_cell_6t_5 inst_cell_33_47 (.BL(BL47),.BLN(BLN47),.WL(WL33));
sram_cell_6t_5 inst_cell_33_48 (.BL(BL48),.BLN(BLN48),.WL(WL33));
sram_cell_6t_5 inst_cell_33_49 (.BL(BL49),.BLN(BLN49),.WL(WL33));
sram_cell_6t_5 inst_cell_33_50 (.BL(BL50),.BLN(BLN50),.WL(WL33));
sram_cell_6t_5 inst_cell_33_51 (.BL(BL51),.BLN(BLN51),.WL(WL33));
sram_cell_6t_5 inst_cell_33_52 (.BL(BL52),.BLN(BLN52),.WL(WL33));
sram_cell_6t_5 inst_cell_33_53 (.BL(BL53),.BLN(BLN53),.WL(WL33));
sram_cell_6t_5 inst_cell_33_54 (.BL(BL54),.BLN(BLN54),.WL(WL33));
sram_cell_6t_5 inst_cell_33_55 (.BL(BL55),.BLN(BLN55),.WL(WL33));
sram_cell_6t_5 inst_cell_33_56 (.BL(BL56),.BLN(BLN56),.WL(WL33));
sram_cell_6t_5 inst_cell_33_57 (.BL(BL57),.BLN(BLN57),.WL(WL33));
sram_cell_6t_5 inst_cell_33_58 (.BL(BL58),.BLN(BLN58),.WL(WL33));
sram_cell_6t_5 inst_cell_33_59 (.BL(BL59),.BLN(BLN59),.WL(WL33));
sram_cell_6t_5 inst_cell_33_60 (.BL(BL60),.BLN(BLN60),.WL(WL33));
sram_cell_6t_5 inst_cell_33_61 (.BL(BL61),.BLN(BLN61),.WL(WL33));
sram_cell_6t_5 inst_cell_33_62 (.BL(BL62),.BLN(BLN62),.WL(WL33));
sram_cell_6t_5 inst_cell_33_63 (.BL(BL63),.BLN(BLN63),.WL(WL33));
sram_cell_6t_5 inst_cell_33_64 (.BL(BL64),.BLN(BLN64),.WL(WL33));
sram_cell_6t_5 inst_cell_33_65 (.BL(BL65),.BLN(BLN65),.WL(WL33));
sram_cell_6t_5 inst_cell_33_66 (.BL(BL66),.BLN(BLN66),.WL(WL33));
sram_cell_6t_5 inst_cell_33_67 (.BL(BL67),.BLN(BLN67),.WL(WL33));
sram_cell_6t_5 inst_cell_33_68 (.BL(BL68),.BLN(BLN68),.WL(WL33));
sram_cell_6t_5 inst_cell_33_69 (.BL(BL69),.BLN(BLN69),.WL(WL33));
sram_cell_6t_5 inst_cell_33_70 (.BL(BL70),.BLN(BLN70),.WL(WL33));
sram_cell_6t_5 inst_cell_33_71 (.BL(BL71),.BLN(BLN71),.WL(WL33));
sram_cell_6t_5 inst_cell_33_72 (.BL(BL72),.BLN(BLN72),.WL(WL33));
sram_cell_6t_5 inst_cell_33_73 (.BL(BL73),.BLN(BLN73),.WL(WL33));
sram_cell_6t_5 inst_cell_33_74 (.BL(BL74),.BLN(BLN74),.WL(WL33));
sram_cell_6t_5 inst_cell_33_75 (.BL(BL75),.BLN(BLN75),.WL(WL33));
sram_cell_6t_5 inst_cell_33_76 (.BL(BL76),.BLN(BLN76),.WL(WL33));
sram_cell_6t_5 inst_cell_33_77 (.BL(BL77),.BLN(BLN77),.WL(WL33));
sram_cell_6t_5 inst_cell_33_78 (.BL(BL78),.BLN(BLN78),.WL(WL33));
sram_cell_6t_5 inst_cell_33_79 (.BL(BL79),.BLN(BLN79),.WL(WL33));
sram_cell_6t_5 inst_cell_33_80 (.BL(BL80),.BLN(BLN80),.WL(WL33));
sram_cell_6t_5 inst_cell_33_81 (.BL(BL81),.BLN(BLN81),.WL(WL33));
sram_cell_6t_5 inst_cell_33_82 (.BL(BL82),.BLN(BLN82),.WL(WL33));
sram_cell_6t_5 inst_cell_33_83 (.BL(BL83),.BLN(BLN83),.WL(WL33));
sram_cell_6t_5 inst_cell_33_84 (.BL(BL84),.BLN(BLN84),.WL(WL33));
sram_cell_6t_5 inst_cell_33_85 (.BL(BL85),.BLN(BLN85),.WL(WL33));
sram_cell_6t_5 inst_cell_33_86 (.BL(BL86),.BLN(BLN86),.WL(WL33));
sram_cell_6t_5 inst_cell_33_87 (.BL(BL87),.BLN(BLN87),.WL(WL33));
sram_cell_6t_5 inst_cell_33_88 (.BL(BL88),.BLN(BLN88),.WL(WL33));
sram_cell_6t_5 inst_cell_33_89 (.BL(BL89),.BLN(BLN89),.WL(WL33));
sram_cell_6t_5 inst_cell_33_90 (.BL(BL90),.BLN(BLN90),.WL(WL33));
sram_cell_6t_5 inst_cell_33_91 (.BL(BL91),.BLN(BLN91),.WL(WL33));
sram_cell_6t_5 inst_cell_33_92 (.BL(BL92),.BLN(BLN92),.WL(WL33));
sram_cell_6t_5 inst_cell_33_93 (.BL(BL93),.BLN(BLN93),.WL(WL33));
sram_cell_6t_5 inst_cell_33_94 (.BL(BL94),.BLN(BLN94),.WL(WL33));
sram_cell_6t_5 inst_cell_33_95 (.BL(BL95),.BLN(BLN95),.WL(WL33));
sram_cell_6t_5 inst_cell_33_96 (.BL(BL96),.BLN(BLN96),.WL(WL33));
sram_cell_6t_5 inst_cell_33_97 (.BL(BL97),.BLN(BLN97),.WL(WL33));
sram_cell_6t_5 inst_cell_33_98 (.BL(BL98),.BLN(BLN98),.WL(WL33));
sram_cell_6t_5 inst_cell_33_99 (.BL(BL99),.BLN(BLN99),.WL(WL33));
sram_cell_6t_5 inst_cell_33_100 (.BL(BL100),.BLN(BLN100),.WL(WL33));
sram_cell_6t_5 inst_cell_33_101 (.BL(BL101),.BLN(BLN101),.WL(WL33));
sram_cell_6t_5 inst_cell_33_102 (.BL(BL102),.BLN(BLN102),.WL(WL33));
sram_cell_6t_5 inst_cell_33_103 (.BL(BL103),.BLN(BLN103),.WL(WL33));
sram_cell_6t_5 inst_cell_33_104 (.BL(BL104),.BLN(BLN104),.WL(WL33));
sram_cell_6t_5 inst_cell_33_105 (.BL(BL105),.BLN(BLN105),.WL(WL33));
sram_cell_6t_5 inst_cell_33_106 (.BL(BL106),.BLN(BLN106),.WL(WL33));
sram_cell_6t_5 inst_cell_33_107 (.BL(BL107),.BLN(BLN107),.WL(WL33));
sram_cell_6t_5 inst_cell_33_108 (.BL(BL108),.BLN(BLN108),.WL(WL33));
sram_cell_6t_5 inst_cell_33_109 (.BL(BL109),.BLN(BLN109),.WL(WL33));
sram_cell_6t_5 inst_cell_33_110 (.BL(BL110),.BLN(BLN110),.WL(WL33));
sram_cell_6t_5 inst_cell_33_111 (.BL(BL111),.BLN(BLN111),.WL(WL33));
sram_cell_6t_5 inst_cell_33_112 (.BL(BL112),.BLN(BLN112),.WL(WL33));
sram_cell_6t_5 inst_cell_33_113 (.BL(BL113),.BLN(BLN113),.WL(WL33));
sram_cell_6t_5 inst_cell_33_114 (.BL(BL114),.BLN(BLN114),.WL(WL33));
sram_cell_6t_5 inst_cell_33_115 (.BL(BL115),.BLN(BLN115),.WL(WL33));
sram_cell_6t_5 inst_cell_33_116 (.BL(BL116),.BLN(BLN116),.WL(WL33));
sram_cell_6t_5 inst_cell_33_117 (.BL(BL117),.BLN(BLN117),.WL(WL33));
sram_cell_6t_5 inst_cell_33_118 (.BL(BL118),.BLN(BLN118),.WL(WL33));
sram_cell_6t_5 inst_cell_33_119 (.BL(BL119),.BLN(BLN119),.WL(WL33));
sram_cell_6t_5 inst_cell_33_120 (.BL(BL120),.BLN(BLN120),.WL(WL33));
sram_cell_6t_5 inst_cell_33_121 (.BL(BL121),.BLN(BLN121),.WL(WL33));
sram_cell_6t_5 inst_cell_33_122 (.BL(BL122),.BLN(BLN122),.WL(WL33));
sram_cell_6t_5 inst_cell_33_123 (.BL(BL123),.BLN(BLN123),.WL(WL33));
sram_cell_6t_5 inst_cell_33_124 (.BL(BL124),.BLN(BLN124),.WL(WL33));
sram_cell_6t_5 inst_cell_33_125 (.BL(BL125),.BLN(BLN125),.WL(WL33));
sram_cell_6t_5 inst_cell_33_126 (.BL(BL126),.BLN(BLN126),.WL(WL33));
sram_cell_6t_5 inst_cell_33_127 (.BL(BL127),.BLN(BLN127),.WL(WL33));
sram_cell_6t_5 inst_cell_34_0 (.BL(BL0),.BLN(BLN0),.WL(WL34));
sram_cell_6t_5 inst_cell_34_1 (.BL(BL1),.BLN(BLN1),.WL(WL34));
sram_cell_6t_5 inst_cell_34_2 (.BL(BL2),.BLN(BLN2),.WL(WL34));
sram_cell_6t_5 inst_cell_34_3 (.BL(BL3),.BLN(BLN3),.WL(WL34));
sram_cell_6t_5 inst_cell_34_4 (.BL(BL4),.BLN(BLN4),.WL(WL34));
sram_cell_6t_5 inst_cell_34_5 (.BL(BL5),.BLN(BLN5),.WL(WL34));
sram_cell_6t_5 inst_cell_34_6 (.BL(BL6),.BLN(BLN6),.WL(WL34));
sram_cell_6t_5 inst_cell_34_7 (.BL(BL7),.BLN(BLN7),.WL(WL34));
sram_cell_6t_5 inst_cell_34_8 (.BL(BL8),.BLN(BLN8),.WL(WL34));
sram_cell_6t_5 inst_cell_34_9 (.BL(BL9),.BLN(BLN9),.WL(WL34));
sram_cell_6t_5 inst_cell_34_10 (.BL(BL10),.BLN(BLN10),.WL(WL34));
sram_cell_6t_5 inst_cell_34_11 (.BL(BL11),.BLN(BLN11),.WL(WL34));
sram_cell_6t_5 inst_cell_34_12 (.BL(BL12),.BLN(BLN12),.WL(WL34));
sram_cell_6t_5 inst_cell_34_13 (.BL(BL13),.BLN(BLN13),.WL(WL34));
sram_cell_6t_5 inst_cell_34_14 (.BL(BL14),.BLN(BLN14),.WL(WL34));
sram_cell_6t_5 inst_cell_34_15 (.BL(BL15),.BLN(BLN15),.WL(WL34));
sram_cell_6t_5 inst_cell_34_16 (.BL(BL16),.BLN(BLN16),.WL(WL34));
sram_cell_6t_5 inst_cell_34_17 (.BL(BL17),.BLN(BLN17),.WL(WL34));
sram_cell_6t_5 inst_cell_34_18 (.BL(BL18),.BLN(BLN18),.WL(WL34));
sram_cell_6t_5 inst_cell_34_19 (.BL(BL19),.BLN(BLN19),.WL(WL34));
sram_cell_6t_5 inst_cell_34_20 (.BL(BL20),.BLN(BLN20),.WL(WL34));
sram_cell_6t_5 inst_cell_34_21 (.BL(BL21),.BLN(BLN21),.WL(WL34));
sram_cell_6t_5 inst_cell_34_22 (.BL(BL22),.BLN(BLN22),.WL(WL34));
sram_cell_6t_5 inst_cell_34_23 (.BL(BL23),.BLN(BLN23),.WL(WL34));
sram_cell_6t_5 inst_cell_34_24 (.BL(BL24),.BLN(BLN24),.WL(WL34));
sram_cell_6t_5 inst_cell_34_25 (.BL(BL25),.BLN(BLN25),.WL(WL34));
sram_cell_6t_5 inst_cell_34_26 (.BL(BL26),.BLN(BLN26),.WL(WL34));
sram_cell_6t_5 inst_cell_34_27 (.BL(BL27),.BLN(BLN27),.WL(WL34));
sram_cell_6t_5 inst_cell_34_28 (.BL(BL28),.BLN(BLN28),.WL(WL34));
sram_cell_6t_5 inst_cell_34_29 (.BL(BL29),.BLN(BLN29),.WL(WL34));
sram_cell_6t_5 inst_cell_34_30 (.BL(BL30),.BLN(BLN30),.WL(WL34));
sram_cell_6t_5 inst_cell_34_31 (.BL(BL31),.BLN(BLN31),.WL(WL34));
sram_cell_6t_5 inst_cell_34_32 (.BL(BL32),.BLN(BLN32),.WL(WL34));
sram_cell_6t_5 inst_cell_34_33 (.BL(BL33),.BLN(BLN33),.WL(WL34));
sram_cell_6t_5 inst_cell_34_34 (.BL(BL34),.BLN(BLN34),.WL(WL34));
sram_cell_6t_5 inst_cell_34_35 (.BL(BL35),.BLN(BLN35),.WL(WL34));
sram_cell_6t_5 inst_cell_34_36 (.BL(BL36),.BLN(BLN36),.WL(WL34));
sram_cell_6t_5 inst_cell_34_37 (.BL(BL37),.BLN(BLN37),.WL(WL34));
sram_cell_6t_5 inst_cell_34_38 (.BL(BL38),.BLN(BLN38),.WL(WL34));
sram_cell_6t_5 inst_cell_34_39 (.BL(BL39),.BLN(BLN39),.WL(WL34));
sram_cell_6t_5 inst_cell_34_40 (.BL(BL40),.BLN(BLN40),.WL(WL34));
sram_cell_6t_5 inst_cell_34_41 (.BL(BL41),.BLN(BLN41),.WL(WL34));
sram_cell_6t_5 inst_cell_34_42 (.BL(BL42),.BLN(BLN42),.WL(WL34));
sram_cell_6t_5 inst_cell_34_43 (.BL(BL43),.BLN(BLN43),.WL(WL34));
sram_cell_6t_5 inst_cell_34_44 (.BL(BL44),.BLN(BLN44),.WL(WL34));
sram_cell_6t_5 inst_cell_34_45 (.BL(BL45),.BLN(BLN45),.WL(WL34));
sram_cell_6t_5 inst_cell_34_46 (.BL(BL46),.BLN(BLN46),.WL(WL34));
sram_cell_6t_5 inst_cell_34_47 (.BL(BL47),.BLN(BLN47),.WL(WL34));
sram_cell_6t_5 inst_cell_34_48 (.BL(BL48),.BLN(BLN48),.WL(WL34));
sram_cell_6t_5 inst_cell_34_49 (.BL(BL49),.BLN(BLN49),.WL(WL34));
sram_cell_6t_5 inst_cell_34_50 (.BL(BL50),.BLN(BLN50),.WL(WL34));
sram_cell_6t_5 inst_cell_34_51 (.BL(BL51),.BLN(BLN51),.WL(WL34));
sram_cell_6t_5 inst_cell_34_52 (.BL(BL52),.BLN(BLN52),.WL(WL34));
sram_cell_6t_5 inst_cell_34_53 (.BL(BL53),.BLN(BLN53),.WL(WL34));
sram_cell_6t_5 inst_cell_34_54 (.BL(BL54),.BLN(BLN54),.WL(WL34));
sram_cell_6t_5 inst_cell_34_55 (.BL(BL55),.BLN(BLN55),.WL(WL34));
sram_cell_6t_5 inst_cell_34_56 (.BL(BL56),.BLN(BLN56),.WL(WL34));
sram_cell_6t_5 inst_cell_34_57 (.BL(BL57),.BLN(BLN57),.WL(WL34));
sram_cell_6t_5 inst_cell_34_58 (.BL(BL58),.BLN(BLN58),.WL(WL34));
sram_cell_6t_5 inst_cell_34_59 (.BL(BL59),.BLN(BLN59),.WL(WL34));
sram_cell_6t_5 inst_cell_34_60 (.BL(BL60),.BLN(BLN60),.WL(WL34));
sram_cell_6t_5 inst_cell_34_61 (.BL(BL61),.BLN(BLN61),.WL(WL34));
sram_cell_6t_5 inst_cell_34_62 (.BL(BL62),.BLN(BLN62),.WL(WL34));
sram_cell_6t_5 inst_cell_34_63 (.BL(BL63),.BLN(BLN63),.WL(WL34));
sram_cell_6t_5 inst_cell_34_64 (.BL(BL64),.BLN(BLN64),.WL(WL34));
sram_cell_6t_5 inst_cell_34_65 (.BL(BL65),.BLN(BLN65),.WL(WL34));
sram_cell_6t_5 inst_cell_34_66 (.BL(BL66),.BLN(BLN66),.WL(WL34));
sram_cell_6t_5 inst_cell_34_67 (.BL(BL67),.BLN(BLN67),.WL(WL34));
sram_cell_6t_5 inst_cell_34_68 (.BL(BL68),.BLN(BLN68),.WL(WL34));
sram_cell_6t_5 inst_cell_34_69 (.BL(BL69),.BLN(BLN69),.WL(WL34));
sram_cell_6t_5 inst_cell_34_70 (.BL(BL70),.BLN(BLN70),.WL(WL34));
sram_cell_6t_5 inst_cell_34_71 (.BL(BL71),.BLN(BLN71),.WL(WL34));
sram_cell_6t_5 inst_cell_34_72 (.BL(BL72),.BLN(BLN72),.WL(WL34));
sram_cell_6t_5 inst_cell_34_73 (.BL(BL73),.BLN(BLN73),.WL(WL34));
sram_cell_6t_5 inst_cell_34_74 (.BL(BL74),.BLN(BLN74),.WL(WL34));
sram_cell_6t_5 inst_cell_34_75 (.BL(BL75),.BLN(BLN75),.WL(WL34));
sram_cell_6t_5 inst_cell_34_76 (.BL(BL76),.BLN(BLN76),.WL(WL34));
sram_cell_6t_5 inst_cell_34_77 (.BL(BL77),.BLN(BLN77),.WL(WL34));
sram_cell_6t_5 inst_cell_34_78 (.BL(BL78),.BLN(BLN78),.WL(WL34));
sram_cell_6t_5 inst_cell_34_79 (.BL(BL79),.BLN(BLN79),.WL(WL34));
sram_cell_6t_5 inst_cell_34_80 (.BL(BL80),.BLN(BLN80),.WL(WL34));
sram_cell_6t_5 inst_cell_34_81 (.BL(BL81),.BLN(BLN81),.WL(WL34));
sram_cell_6t_5 inst_cell_34_82 (.BL(BL82),.BLN(BLN82),.WL(WL34));
sram_cell_6t_5 inst_cell_34_83 (.BL(BL83),.BLN(BLN83),.WL(WL34));
sram_cell_6t_5 inst_cell_34_84 (.BL(BL84),.BLN(BLN84),.WL(WL34));
sram_cell_6t_5 inst_cell_34_85 (.BL(BL85),.BLN(BLN85),.WL(WL34));
sram_cell_6t_5 inst_cell_34_86 (.BL(BL86),.BLN(BLN86),.WL(WL34));
sram_cell_6t_5 inst_cell_34_87 (.BL(BL87),.BLN(BLN87),.WL(WL34));
sram_cell_6t_5 inst_cell_34_88 (.BL(BL88),.BLN(BLN88),.WL(WL34));
sram_cell_6t_5 inst_cell_34_89 (.BL(BL89),.BLN(BLN89),.WL(WL34));
sram_cell_6t_5 inst_cell_34_90 (.BL(BL90),.BLN(BLN90),.WL(WL34));
sram_cell_6t_5 inst_cell_34_91 (.BL(BL91),.BLN(BLN91),.WL(WL34));
sram_cell_6t_5 inst_cell_34_92 (.BL(BL92),.BLN(BLN92),.WL(WL34));
sram_cell_6t_5 inst_cell_34_93 (.BL(BL93),.BLN(BLN93),.WL(WL34));
sram_cell_6t_5 inst_cell_34_94 (.BL(BL94),.BLN(BLN94),.WL(WL34));
sram_cell_6t_5 inst_cell_34_95 (.BL(BL95),.BLN(BLN95),.WL(WL34));
sram_cell_6t_5 inst_cell_34_96 (.BL(BL96),.BLN(BLN96),.WL(WL34));
sram_cell_6t_5 inst_cell_34_97 (.BL(BL97),.BLN(BLN97),.WL(WL34));
sram_cell_6t_5 inst_cell_34_98 (.BL(BL98),.BLN(BLN98),.WL(WL34));
sram_cell_6t_5 inst_cell_34_99 (.BL(BL99),.BLN(BLN99),.WL(WL34));
sram_cell_6t_5 inst_cell_34_100 (.BL(BL100),.BLN(BLN100),.WL(WL34));
sram_cell_6t_5 inst_cell_34_101 (.BL(BL101),.BLN(BLN101),.WL(WL34));
sram_cell_6t_5 inst_cell_34_102 (.BL(BL102),.BLN(BLN102),.WL(WL34));
sram_cell_6t_5 inst_cell_34_103 (.BL(BL103),.BLN(BLN103),.WL(WL34));
sram_cell_6t_5 inst_cell_34_104 (.BL(BL104),.BLN(BLN104),.WL(WL34));
sram_cell_6t_5 inst_cell_34_105 (.BL(BL105),.BLN(BLN105),.WL(WL34));
sram_cell_6t_5 inst_cell_34_106 (.BL(BL106),.BLN(BLN106),.WL(WL34));
sram_cell_6t_5 inst_cell_34_107 (.BL(BL107),.BLN(BLN107),.WL(WL34));
sram_cell_6t_5 inst_cell_34_108 (.BL(BL108),.BLN(BLN108),.WL(WL34));
sram_cell_6t_5 inst_cell_34_109 (.BL(BL109),.BLN(BLN109),.WL(WL34));
sram_cell_6t_5 inst_cell_34_110 (.BL(BL110),.BLN(BLN110),.WL(WL34));
sram_cell_6t_5 inst_cell_34_111 (.BL(BL111),.BLN(BLN111),.WL(WL34));
sram_cell_6t_5 inst_cell_34_112 (.BL(BL112),.BLN(BLN112),.WL(WL34));
sram_cell_6t_5 inst_cell_34_113 (.BL(BL113),.BLN(BLN113),.WL(WL34));
sram_cell_6t_5 inst_cell_34_114 (.BL(BL114),.BLN(BLN114),.WL(WL34));
sram_cell_6t_5 inst_cell_34_115 (.BL(BL115),.BLN(BLN115),.WL(WL34));
sram_cell_6t_5 inst_cell_34_116 (.BL(BL116),.BLN(BLN116),.WL(WL34));
sram_cell_6t_5 inst_cell_34_117 (.BL(BL117),.BLN(BLN117),.WL(WL34));
sram_cell_6t_5 inst_cell_34_118 (.BL(BL118),.BLN(BLN118),.WL(WL34));
sram_cell_6t_5 inst_cell_34_119 (.BL(BL119),.BLN(BLN119),.WL(WL34));
sram_cell_6t_5 inst_cell_34_120 (.BL(BL120),.BLN(BLN120),.WL(WL34));
sram_cell_6t_5 inst_cell_34_121 (.BL(BL121),.BLN(BLN121),.WL(WL34));
sram_cell_6t_5 inst_cell_34_122 (.BL(BL122),.BLN(BLN122),.WL(WL34));
sram_cell_6t_5 inst_cell_34_123 (.BL(BL123),.BLN(BLN123),.WL(WL34));
sram_cell_6t_5 inst_cell_34_124 (.BL(BL124),.BLN(BLN124),.WL(WL34));
sram_cell_6t_5 inst_cell_34_125 (.BL(BL125),.BLN(BLN125),.WL(WL34));
sram_cell_6t_5 inst_cell_34_126 (.BL(BL126),.BLN(BLN126),.WL(WL34));
sram_cell_6t_5 inst_cell_34_127 (.BL(BL127),.BLN(BLN127),.WL(WL34));
sram_cell_6t_5 inst_cell_35_0 (.BL(BL0),.BLN(BLN0),.WL(WL35));
sram_cell_6t_5 inst_cell_35_1 (.BL(BL1),.BLN(BLN1),.WL(WL35));
sram_cell_6t_5 inst_cell_35_2 (.BL(BL2),.BLN(BLN2),.WL(WL35));
sram_cell_6t_5 inst_cell_35_3 (.BL(BL3),.BLN(BLN3),.WL(WL35));
sram_cell_6t_5 inst_cell_35_4 (.BL(BL4),.BLN(BLN4),.WL(WL35));
sram_cell_6t_5 inst_cell_35_5 (.BL(BL5),.BLN(BLN5),.WL(WL35));
sram_cell_6t_5 inst_cell_35_6 (.BL(BL6),.BLN(BLN6),.WL(WL35));
sram_cell_6t_5 inst_cell_35_7 (.BL(BL7),.BLN(BLN7),.WL(WL35));
sram_cell_6t_5 inst_cell_35_8 (.BL(BL8),.BLN(BLN8),.WL(WL35));
sram_cell_6t_5 inst_cell_35_9 (.BL(BL9),.BLN(BLN9),.WL(WL35));
sram_cell_6t_5 inst_cell_35_10 (.BL(BL10),.BLN(BLN10),.WL(WL35));
sram_cell_6t_5 inst_cell_35_11 (.BL(BL11),.BLN(BLN11),.WL(WL35));
sram_cell_6t_5 inst_cell_35_12 (.BL(BL12),.BLN(BLN12),.WL(WL35));
sram_cell_6t_5 inst_cell_35_13 (.BL(BL13),.BLN(BLN13),.WL(WL35));
sram_cell_6t_5 inst_cell_35_14 (.BL(BL14),.BLN(BLN14),.WL(WL35));
sram_cell_6t_5 inst_cell_35_15 (.BL(BL15),.BLN(BLN15),.WL(WL35));
sram_cell_6t_5 inst_cell_35_16 (.BL(BL16),.BLN(BLN16),.WL(WL35));
sram_cell_6t_5 inst_cell_35_17 (.BL(BL17),.BLN(BLN17),.WL(WL35));
sram_cell_6t_5 inst_cell_35_18 (.BL(BL18),.BLN(BLN18),.WL(WL35));
sram_cell_6t_5 inst_cell_35_19 (.BL(BL19),.BLN(BLN19),.WL(WL35));
sram_cell_6t_5 inst_cell_35_20 (.BL(BL20),.BLN(BLN20),.WL(WL35));
sram_cell_6t_5 inst_cell_35_21 (.BL(BL21),.BLN(BLN21),.WL(WL35));
sram_cell_6t_5 inst_cell_35_22 (.BL(BL22),.BLN(BLN22),.WL(WL35));
sram_cell_6t_5 inst_cell_35_23 (.BL(BL23),.BLN(BLN23),.WL(WL35));
sram_cell_6t_5 inst_cell_35_24 (.BL(BL24),.BLN(BLN24),.WL(WL35));
sram_cell_6t_5 inst_cell_35_25 (.BL(BL25),.BLN(BLN25),.WL(WL35));
sram_cell_6t_5 inst_cell_35_26 (.BL(BL26),.BLN(BLN26),.WL(WL35));
sram_cell_6t_5 inst_cell_35_27 (.BL(BL27),.BLN(BLN27),.WL(WL35));
sram_cell_6t_5 inst_cell_35_28 (.BL(BL28),.BLN(BLN28),.WL(WL35));
sram_cell_6t_5 inst_cell_35_29 (.BL(BL29),.BLN(BLN29),.WL(WL35));
sram_cell_6t_5 inst_cell_35_30 (.BL(BL30),.BLN(BLN30),.WL(WL35));
sram_cell_6t_5 inst_cell_35_31 (.BL(BL31),.BLN(BLN31),.WL(WL35));
sram_cell_6t_5 inst_cell_35_32 (.BL(BL32),.BLN(BLN32),.WL(WL35));
sram_cell_6t_5 inst_cell_35_33 (.BL(BL33),.BLN(BLN33),.WL(WL35));
sram_cell_6t_5 inst_cell_35_34 (.BL(BL34),.BLN(BLN34),.WL(WL35));
sram_cell_6t_5 inst_cell_35_35 (.BL(BL35),.BLN(BLN35),.WL(WL35));
sram_cell_6t_5 inst_cell_35_36 (.BL(BL36),.BLN(BLN36),.WL(WL35));
sram_cell_6t_5 inst_cell_35_37 (.BL(BL37),.BLN(BLN37),.WL(WL35));
sram_cell_6t_5 inst_cell_35_38 (.BL(BL38),.BLN(BLN38),.WL(WL35));
sram_cell_6t_5 inst_cell_35_39 (.BL(BL39),.BLN(BLN39),.WL(WL35));
sram_cell_6t_5 inst_cell_35_40 (.BL(BL40),.BLN(BLN40),.WL(WL35));
sram_cell_6t_5 inst_cell_35_41 (.BL(BL41),.BLN(BLN41),.WL(WL35));
sram_cell_6t_5 inst_cell_35_42 (.BL(BL42),.BLN(BLN42),.WL(WL35));
sram_cell_6t_5 inst_cell_35_43 (.BL(BL43),.BLN(BLN43),.WL(WL35));
sram_cell_6t_5 inst_cell_35_44 (.BL(BL44),.BLN(BLN44),.WL(WL35));
sram_cell_6t_5 inst_cell_35_45 (.BL(BL45),.BLN(BLN45),.WL(WL35));
sram_cell_6t_5 inst_cell_35_46 (.BL(BL46),.BLN(BLN46),.WL(WL35));
sram_cell_6t_5 inst_cell_35_47 (.BL(BL47),.BLN(BLN47),.WL(WL35));
sram_cell_6t_5 inst_cell_35_48 (.BL(BL48),.BLN(BLN48),.WL(WL35));
sram_cell_6t_5 inst_cell_35_49 (.BL(BL49),.BLN(BLN49),.WL(WL35));
sram_cell_6t_5 inst_cell_35_50 (.BL(BL50),.BLN(BLN50),.WL(WL35));
sram_cell_6t_5 inst_cell_35_51 (.BL(BL51),.BLN(BLN51),.WL(WL35));
sram_cell_6t_5 inst_cell_35_52 (.BL(BL52),.BLN(BLN52),.WL(WL35));
sram_cell_6t_5 inst_cell_35_53 (.BL(BL53),.BLN(BLN53),.WL(WL35));
sram_cell_6t_5 inst_cell_35_54 (.BL(BL54),.BLN(BLN54),.WL(WL35));
sram_cell_6t_5 inst_cell_35_55 (.BL(BL55),.BLN(BLN55),.WL(WL35));
sram_cell_6t_5 inst_cell_35_56 (.BL(BL56),.BLN(BLN56),.WL(WL35));
sram_cell_6t_5 inst_cell_35_57 (.BL(BL57),.BLN(BLN57),.WL(WL35));
sram_cell_6t_5 inst_cell_35_58 (.BL(BL58),.BLN(BLN58),.WL(WL35));
sram_cell_6t_5 inst_cell_35_59 (.BL(BL59),.BLN(BLN59),.WL(WL35));
sram_cell_6t_5 inst_cell_35_60 (.BL(BL60),.BLN(BLN60),.WL(WL35));
sram_cell_6t_5 inst_cell_35_61 (.BL(BL61),.BLN(BLN61),.WL(WL35));
sram_cell_6t_5 inst_cell_35_62 (.BL(BL62),.BLN(BLN62),.WL(WL35));
sram_cell_6t_5 inst_cell_35_63 (.BL(BL63),.BLN(BLN63),.WL(WL35));
sram_cell_6t_5 inst_cell_35_64 (.BL(BL64),.BLN(BLN64),.WL(WL35));
sram_cell_6t_5 inst_cell_35_65 (.BL(BL65),.BLN(BLN65),.WL(WL35));
sram_cell_6t_5 inst_cell_35_66 (.BL(BL66),.BLN(BLN66),.WL(WL35));
sram_cell_6t_5 inst_cell_35_67 (.BL(BL67),.BLN(BLN67),.WL(WL35));
sram_cell_6t_5 inst_cell_35_68 (.BL(BL68),.BLN(BLN68),.WL(WL35));
sram_cell_6t_5 inst_cell_35_69 (.BL(BL69),.BLN(BLN69),.WL(WL35));
sram_cell_6t_5 inst_cell_35_70 (.BL(BL70),.BLN(BLN70),.WL(WL35));
sram_cell_6t_5 inst_cell_35_71 (.BL(BL71),.BLN(BLN71),.WL(WL35));
sram_cell_6t_5 inst_cell_35_72 (.BL(BL72),.BLN(BLN72),.WL(WL35));
sram_cell_6t_5 inst_cell_35_73 (.BL(BL73),.BLN(BLN73),.WL(WL35));
sram_cell_6t_5 inst_cell_35_74 (.BL(BL74),.BLN(BLN74),.WL(WL35));
sram_cell_6t_5 inst_cell_35_75 (.BL(BL75),.BLN(BLN75),.WL(WL35));
sram_cell_6t_5 inst_cell_35_76 (.BL(BL76),.BLN(BLN76),.WL(WL35));
sram_cell_6t_5 inst_cell_35_77 (.BL(BL77),.BLN(BLN77),.WL(WL35));
sram_cell_6t_5 inst_cell_35_78 (.BL(BL78),.BLN(BLN78),.WL(WL35));
sram_cell_6t_5 inst_cell_35_79 (.BL(BL79),.BLN(BLN79),.WL(WL35));
sram_cell_6t_5 inst_cell_35_80 (.BL(BL80),.BLN(BLN80),.WL(WL35));
sram_cell_6t_5 inst_cell_35_81 (.BL(BL81),.BLN(BLN81),.WL(WL35));
sram_cell_6t_5 inst_cell_35_82 (.BL(BL82),.BLN(BLN82),.WL(WL35));
sram_cell_6t_5 inst_cell_35_83 (.BL(BL83),.BLN(BLN83),.WL(WL35));
sram_cell_6t_5 inst_cell_35_84 (.BL(BL84),.BLN(BLN84),.WL(WL35));
sram_cell_6t_5 inst_cell_35_85 (.BL(BL85),.BLN(BLN85),.WL(WL35));
sram_cell_6t_5 inst_cell_35_86 (.BL(BL86),.BLN(BLN86),.WL(WL35));
sram_cell_6t_5 inst_cell_35_87 (.BL(BL87),.BLN(BLN87),.WL(WL35));
sram_cell_6t_5 inst_cell_35_88 (.BL(BL88),.BLN(BLN88),.WL(WL35));
sram_cell_6t_5 inst_cell_35_89 (.BL(BL89),.BLN(BLN89),.WL(WL35));
sram_cell_6t_5 inst_cell_35_90 (.BL(BL90),.BLN(BLN90),.WL(WL35));
sram_cell_6t_5 inst_cell_35_91 (.BL(BL91),.BLN(BLN91),.WL(WL35));
sram_cell_6t_5 inst_cell_35_92 (.BL(BL92),.BLN(BLN92),.WL(WL35));
sram_cell_6t_5 inst_cell_35_93 (.BL(BL93),.BLN(BLN93),.WL(WL35));
sram_cell_6t_5 inst_cell_35_94 (.BL(BL94),.BLN(BLN94),.WL(WL35));
sram_cell_6t_5 inst_cell_35_95 (.BL(BL95),.BLN(BLN95),.WL(WL35));
sram_cell_6t_5 inst_cell_35_96 (.BL(BL96),.BLN(BLN96),.WL(WL35));
sram_cell_6t_5 inst_cell_35_97 (.BL(BL97),.BLN(BLN97),.WL(WL35));
sram_cell_6t_5 inst_cell_35_98 (.BL(BL98),.BLN(BLN98),.WL(WL35));
sram_cell_6t_5 inst_cell_35_99 (.BL(BL99),.BLN(BLN99),.WL(WL35));
sram_cell_6t_5 inst_cell_35_100 (.BL(BL100),.BLN(BLN100),.WL(WL35));
sram_cell_6t_5 inst_cell_35_101 (.BL(BL101),.BLN(BLN101),.WL(WL35));
sram_cell_6t_5 inst_cell_35_102 (.BL(BL102),.BLN(BLN102),.WL(WL35));
sram_cell_6t_5 inst_cell_35_103 (.BL(BL103),.BLN(BLN103),.WL(WL35));
sram_cell_6t_5 inst_cell_35_104 (.BL(BL104),.BLN(BLN104),.WL(WL35));
sram_cell_6t_5 inst_cell_35_105 (.BL(BL105),.BLN(BLN105),.WL(WL35));
sram_cell_6t_5 inst_cell_35_106 (.BL(BL106),.BLN(BLN106),.WL(WL35));
sram_cell_6t_5 inst_cell_35_107 (.BL(BL107),.BLN(BLN107),.WL(WL35));
sram_cell_6t_5 inst_cell_35_108 (.BL(BL108),.BLN(BLN108),.WL(WL35));
sram_cell_6t_5 inst_cell_35_109 (.BL(BL109),.BLN(BLN109),.WL(WL35));
sram_cell_6t_5 inst_cell_35_110 (.BL(BL110),.BLN(BLN110),.WL(WL35));
sram_cell_6t_5 inst_cell_35_111 (.BL(BL111),.BLN(BLN111),.WL(WL35));
sram_cell_6t_5 inst_cell_35_112 (.BL(BL112),.BLN(BLN112),.WL(WL35));
sram_cell_6t_5 inst_cell_35_113 (.BL(BL113),.BLN(BLN113),.WL(WL35));
sram_cell_6t_5 inst_cell_35_114 (.BL(BL114),.BLN(BLN114),.WL(WL35));
sram_cell_6t_5 inst_cell_35_115 (.BL(BL115),.BLN(BLN115),.WL(WL35));
sram_cell_6t_5 inst_cell_35_116 (.BL(BL116),.BLN(BLN116),.WL(WL35));
sram_cell_6t_5 inst_cell_35_117 (.BL(BL117),.BLN(BLN117),.WL(WL35));
sram_cell_6t_5 inst_cell_35_118 (.BL(BL118),.BLN(BLN118),.WL(WL35));
sram_cell_6t_5 inst_cell_35_119 (.BL(BL119),.BLN(BLN119),.WL(WL35));
sram_cell_6t_5 inst_cell_35_120 (.BL(BL120),.BLN(BLN120),.WL(WL35));
sram_cell_6t_5 inst_cell_35_121 (.BL(BL121),.BLN(BLN121),.WL(WL35));
sram_cell_6t_5 inst_cell_35_122 (.BL(BL122),.BLN(BLN122),.WL(WL35));
sram_cell_6t_5 inst_cell_35_123 (.BL(BL123),.BLN(BLN123),.WL(WL35));
sram_cell_6t_5 inst_cell_35_124 (.BL(BL124),.BLN(BLN124),.WL(WL35));
sram_cell_6t_5 inst_cell_35_125 (.BL(BL125),.BLN(BLN125),.WL(WL35));
sram_cell_6t_5 inst_cell_35_126 (.BL(BL126),.BLN(BLN126),.WL(WL35));
sram_cell_6t_5 inst_cell_35_127 (.BL(BL127),.BLN(BLN127),.WL(WL35));
sram_cell_6t_5 inst_cell_36_0 (.BL(BL0),.BLN(BLN0),.WL(WL36));
sram_cell_6t_5 inst_cell_36_1 (.BL(BL1),.BLN(BLN1),.WL(WL36));
sram_cell_6t_5 inst_cell_36_2 (.BL(BL2),.BLN(BLN2),.WL(WL36));
sram_cell_6t_5 inst_cell_36_3 (.BL(BL3),.BLN(BLN3),.WL(WL36));
sram_cell_6t_5 inst_cell_36_4 (.BL(BL4),.BLN(BLN4),.WL(WL36));
sram_cell_6t_5 inst_cell_36_5 (.BL(BL5),.BLN(BLN5),.WL(WL36));
sram_cell_6t_5 inst_cell_36_6 (.BL(BL6),.BLN(BLN6),.WL(WL36));
sram_cell_6t_5 inst_cell_36_7 (.BL(BL7),.BLN(BLN7),.WL(WL36));
sram_cell_6t_5 inst_cell_36_8 (.BL(BL8),.BLN(BLN8),.WL(WL36));
sram_cell_6t_5 inst_cell_36_9 (.BL(BL9),.BLN(BLN9),.WL(WL36));
sram_cell_6t_5 inst_cell_36_10 (.BL(BL10),.BLN(BLN10),.WL(WL36));
sram_cell_6t_5 inst_cell_36_11 (.BL(BL11),.BLN(BLN11),.WL(WL36));
sram_cell_6t_5 inst_cell_36_12 (.BL(BL12),.BLN(BLN12),.WL(WL36));
sram_cell_6t_5 inst_cell_36_13 (.BL(BL13),.BLN(BLN13),.WL(WL36));
sram_cell_6t_5 inst_cell_36_14 (.BL(BL14),.BLN(BLN14),.WL(WL36));
sram_cell_6t_5 inst_cell_36_15 (.BL(BL15),.BLN(BLN15),.WL(WL36));
sram_cell_6t_5 inst_cell_36_16 (.BL(BL16),.BLN(BLN16),.WL(WL36));
sram_cell_6t_5 inst_cell_36_17 (.BL(BL17),.BLN(BLN17),.WL(WL36));
sram_cell_6t_5 inst_cell_36_18 (.BL(BL18),.BLN(BLN18),.WL(WL36));
sram_cell_6t_5 inst_cell_36_19 (.BL(BL19),.BLN(BLN19),.WL(WL36));
sram_cell_6t_5 inst_cell_36_20 (.BL(BL20),.BLN(BLN20),.WL(WL36));
sram_cell_6t_5 inst_cell_36_21 (.BL(BL21),.BLN(BLN21),.WL(WL36));
sram_cell_6t_5 inst_cell_36_22 (.BL(BL22),.BLN(BLN22),.WL(WL36));
sram_cell_6t_5 inst_cell_36_23 (.BL(BL23),.BLN(BLN23),.WL(WL36));
sram_cell_6t_5 inst_cell_36_24 (.BL(BL24),.BLN(BLN24),.WL(WL36));
sram_cell_6t_5 inst_cell_36_25 (.BL(BL25),.BLN(BLN25),.WL(WL36));
sram_cell_6t_5 inst_cell_36_26 (.BL(BL26),.BLN(BLN26),.WL(WL36));
sram_cell_6t_5 inst_cell_36_27 (.BL(BL27),.BLN(BLN27),.WL(WL36));
sram_cell_6t_5 inst_cell_36_28 (.BL(BL28),.BLN(BLN28),.WL(WL36));
sram_cell_6t_5 inst_cell_36_29 (.BL(BL29),.BLN(BLN29),.WL(WL36));
sram_cell_6t_5 inst_cell_36_30 (.BL(BL30),.BLN(BLN30),.WL(WL36));
sram_cell_6t_5 inst_cell_36_31 (.BL(BL31),.BLN(BLN31),.WL(WL36));
sram_cell_6t_5 inst_cell_36_32 (.BL(BL32),.BLN(BLN32),.WL(WL36));
sram_cell_6t_5 inst_cell_36_33 (.BL(BL33),.BLN(BLN33),.WL(WL36));
sram_cell_6t_5 inst_cell_36_34 (.BL(BL34),.BLN(BLN34),.WL(WL36));
sram_cell_6t_5 inst_cell_36_35 (.BL(BL35),.BLN(BLN35),.WL(WL36));
sram_cell_6t_5 inst_cell_36_36 (.BL(BL36),.BLN(BLN36),.WL(WL36));
sram_cell_6t_5 inst_cell_36_37 (.BL(BL37),.BLN(BLN37),.WL(WL36));
sram_cell_6t_5 inst_cell_36_38 (.BL(BL38),.BLN(BLN38),.WL(WL36));
sram_cell_6t_5 inst_cell_36_39 (.BL(BL39),.BLN(BLN39),.WL(WL36));
sram_cell_6t_5 inst_cell_36_40 (.BL(BL40),.BLN(BLN40),.WL(WL36));
sram_cell_6t_5 inst_cell_36_41 (.BL(BL41),.BLN(BLN41),.WL(WL36));
sram_cell_6t_5 inst_cell_36_42 (.BL(BL42),.BLN(BLN42),.WL(WL36));
sram_cell_6t_5 inst_cell_36_43 (.BL(BL43),.BLN(BLN43),.WL(WL36));
sram_cell_6t_5 inst_cell_36_44 (.BL(BL44),.BLN(BLN44),.WL(WL36));
sram_cell_6t_5 inst_cell_36_45 (.BL(BL45),.BLN(BLN45),.WL(WL36));
sram_cell_6t_5 inst_cell_36_46 (.BL(BL46),.BLN(BLN46),.WL(WL36));
sram_cell_6t_5 inst_cell_36_47 (.BL(BL47),.BLN(BLN47),.WL(WL36));
sram_cell_6t_5 inst_cell_36_48 (.BL(BL48),.BLN(BLN48),.WL(WL36));
sram_cell_6t_5 inst_cell_36_49 (.BL(BL49),.BLN(BLN49),.WL(WL36));
sram_cell_6t_5 inst_cell_36_50 (.BL(BL50),.BLN(BLN50),.WL(WL36));
sram_cell_6t_5 inst_cell_36_51 (.BL(BL51),.BLN(BLN51),.WL(WL36));
sram_cell_6t_5 inst_cell_36_52 (.BL(BL52),.BLN(BLN52),.WL(WL36));
sram_cell_6t_5 inst_cell_36_53 (.BL(BL53),.BLN(BLN53),.WL(WL36));
sram_cell_6t_5 inst_cell_36_54 (.BL(BL54),.BLN(BLN54),.WL(WL36));
sram_cell_6t_5 inst_cell_36_55 (.BL(BL55),.BLN(BLN55),.WL(WL36));
sram_cell_6t_5 inst_cell_36_56 (.BL(BL56),.BLN(BLN56),.WL(WL36));
sram_cell_6t_5 inst_cell_36_57 (.BL(BL57),.BLN(BLN57),.WL(WL36));
sram_cell_6t_5 inst_cell_36_58 (.BL(BL58),.BLN(BLN58),.WL(WL36));
sram_cell_6t_5 inst_cell_36_59 (.BL(BL59),.BLN(BLN59),.WL(WL36));
sram_cell_6t_5 inst_cell_36_60 (.BL(BL60),.BLN(BLN60),.WL(WL36));
sram_cell_6t_5 inst_cell_36_61 (.BL(BL61),.BLN(BLN61),.WL(WL36));
sram_cell_6t_5 inst_cell_36_62 (.BL(BL62),.BLN(BLN62),.WL(WL36));
sram_cell_6t_5 inst_cell_36_63 (.BL(BL63),.BLN(BLN63),.WL(WL36));
sram_cell_6t_5 inst_cell_36_64 (.BL(BL64),.BLN(BLN64),.WL(WL36));
sram_cell_6t_5 inst_cell_36_65 (.BL(BL65),.BLN(BLN65),.WL(WL36));
sram_cell_6t_5 inst_cell_36_66 (.BL(BL66),.BLN(BLN66),.WL(WL36));
sram_cell_6t_5 inst_cell_36_67 (.BL(BL67),.BLN(BLN67),.WL(WL36));
sram_cell_6t_5 inst_cell_36_68 (.BL(BL68),.BLN(BLN68),.WL(WL36));
sram_cell_6t_5 inst_cell_36_69 (.BL(BL69),.BLN(BLN69),.WL(WL36));
sram_cell_6t_5 inst_cell_36_70 (.BL(BL70),.BLN(BLN70),.WL(WL36));
sram_cell_6t_5 inst_cell_36_71 (.BL(BL71),.BLN(BLN71),.WL(WL36));
sram_cell_6t_5 inst_cell_36_72 (.BL(BL72),.BLN(BLN72),.WL(WL36));
sram_cell_6t_5 inst_cell_36_73 (.BL(BL73),.BLN(BLN73),.WL(WL36));
sram_cell_6t_5 inst_cell_36_74 (.BL(BL74),.BLN(BLN74),.WL(WL36));
sram_cell_6t_5 inst_cell_36_75 (.BL(BL75),.BLN(BLN75),.WL(WL36));
sram_cell_6t_5 inst_cell_36_76 (.BL(BL76),.BLN(BLN76),.WL(WL36));
sram_cell_6t_5 inst_cell_36_77 (.BL(BL77),.BLN(BLN77),.WL(WL36));
sram_cell_6t_5 inst_cell_36_78 (.BL(BL78),.BLN(BLN78),.WL(WL36));
sram_cell_6t_5 inst_cell_36_79 (.BL(BL79),.BLN(BLN79),.WL(WL36));
sram_cell_6t_5 inst_cell_36_80 (.BL(BL80),.BLN(BLN80),.WL(WL36));
sram_cell_6t_5 inst_cell_36_81 (.BL(BL81),.BLN(BLN81),.WL(WL36));
sram_cell_6t_5 inst_cell_36_82 (.BL(BL82),.BLN(BLN82),.WL(WL36));
sram_cell_6t_5 inst_cell_36_83 (.BL(BL83),.BLN(BLN83),.WL(WL36));
sram_cell_6t_5 inst_cell_36_84 (.BL(BL84),.BLN(BLN84),.WL(WL36));
sram_cell_6t_5 inst_cell_36_85 (.BL(BL85),.BLN(BLN85),.WL(WL36));
sram_cell_6t_5 inst_cell_36_86 (.BL(BL86),.BLN(BLN86),.WL(WL36));
sram_cell_6t_5 inst_cell_36_87 (.BL(BL87),.BLN(BLN87),.WL(WL36));
sram_cell_6t_5 inst_cell_36_88 (.BL(BL88),.BLN(BLN88),.WL(WL36));
sram_cell_6t_5 inst_cell_36_89 (.BL(BL89),.BLN(BLN89),.WL(WL36));
sram_cell_6t_5 inst_cell_36_90 (.BL(BL90),.BLN(BLN90),.WL(WL36));
sram_cell_6t_5 inst_cell_36_91 (.BL(BL91),.BLN(BLN91),.WL(WL36));
sram_cell_6t_5 inst_cell_36_92 (.BL(BL92),.BLN(BLN92),.WL(WL36));
sram_cell_6t_5 inst_cell_36_93 (.BL(BL93),.BLN(BLN93),.WL(WL36));
sram_cell_6t_5 inst_cell_36_94 (.BL(BL94),.BLN(BLN94),.WL(WL36));
sram_cell_6t_5 inst_cell_36_95 (.BL(BL95),.BLN(BLN95),.WL(WL36));
sram_cell_6t_5 inst_cell_36_96 (.BL(BL96),.BLN(BLN96),.WL(WL36));
sram_cell_6t_5 inst_cell_36_97 (.BL(BL97),.BLN(BLN97),.WL(WL36));
sram_cell_6t_5 inst_cell_36_98 (.BL(BL98),.BLN(BLN98),.WL(WL36));
sram_cell_6t_5 inst_cell_36_99 (.BL(BL99),.BLN(BLN99),.WL(WL36));
sram_cell_6t_5 inst_cell_36_100 (.BL(BL100),.BLN(BLN100),.WL(WL36));
sram_cell_6t_5 inst_cell_36_101 (.BL(BL101),.BLN(BLN101),.WL(WL36));
sram_cell_6t_5 inst_cell_36_102 (.BL(BL102),.BLN(BLN102),.WL(WL36));
sram_cell_6t_5 inst_cell_36_103 (.BL(BL103),.BLN(BLN103),.WL(WL36));
sram_cell_6t_5 inst_cell_36_104 (.BL(BL104),.BLN(BLN104),.WL(WL36));
sram_cell_6t_5 inst_cell_36_105 (.BL(BL105),.BLN(BLN105),.WL(WL36));
sram_cell_6t_5 inst_cell_36_106 (.BL(BL106),.BLN(BLN106),.WL(WL36));
sram_cell_6t_5 inst_cell_36_107 (.BL(BL107),.BLN(BLN107),.WL(WL36));
sram_cell_6t_5 inst_cell_36_108 (.BL(BL108),.BLN(BLN108),.WL(WL36));
sram_cell_6t_5 inst_cell_36_109 (.BL(BL109),.BLN(BLN109),.WL(WL36));
sram_cell_6t_5 inst_cell_36_110 (.BL(BL110),.BLN(BLN110),.WL(WL36));
sram_cell_6t_5 inst_cell_36_111 (.BL(BL111),.BLN(BLN111),.WL(WL36));
sram_cell_6t_5 inst_cell_36_112 (.BL(BL112),.BLN(BLN112),.WL(WL36));
sram_cell_6t_5 inst_cell_36_113 (.BL(BL113),.BLN(BLN113),.WL(WL36));
sram_cell_6t_5 inst_cell_36_114 (.BL(BL114),.BLN(BLN114),.WL(WL36));
sram_cell_6t_5 inst_cell_36_115 (.BL(BL115),.BLN(BLN115),.WL(WL36));
sram_cell_6t_5 inst_cell_36_116 (.BL(BL116),.BLN(BLN116),.WL(WL36));
sram_cell_6t_5 inst_cell_36_117 (.BL(BL117),.BLN(BLN117),.WL(WL36));
sram_cell_6t_5 inst_cell_36_118 (.BL(BL118),.BLN(BLN118),.WL(WL36));
sram_cell_6t_5 inst_cell_36_119 (.BL(BL119),.BLN(BLN119),.WL(WL36));
sram_cell_6t_5 inst_cell_36_120 (.BL(BL120),.BLN(BLN120),.WL(WL36));
sram_cell_6t_5 inst_cell_36_121 (.BL(BL121),.BLN(BLN121),.WL(WL36));
sram_cell_6t_5 inst_cell_36_122 (.BL(BL122),.BLN(BLN122),.WL(WL36));
sram_cell_6t_5 inst_cell_36_123 (.BL(BL123),.BLN(BLN123),.WL(WL36));
sram_cell_6t_5 inst_cell_36_124 (.BL(BL124),.BLN(BLN124),.WL(WL36));
sram_cell_6t_5 inst_cell_36_125 (.BL(BL125),.BLN(BLN125),.WL(WL36));
sram_cell_6t_5 inst_cell_36_126 (.BL(BL126),.BLN(BLN126),.WL(WL36));
sram_cell_6t_5 inst_cell_36_127 (.BL(BL127),.BLN(BLN127),.WL(WL36));
sram_cell_6t_5 inst_cell_37_0 (.BL(BL0),.BLN(BLN0),.WL(WL37));
sram_cell_6t_5 inst_cell_37_1 (.BL(BL1),.BLN(BLN1),.WL(WL37));
sram_cell_6t_5 inst_cell_37_2 (.BL(BL2),.BLN(BLN2),.WL(WL37));
sram_cell_6t_5 inst_cell_37_3 (.BL(BL3),.BLN(BLN3),.WL(WL37));
sram_cell_6t_5 inst_cell_37_4 (.BL(BL4),.BLN(BLN4),.WL(WL37));
sram_cell_6t_5 inst_cell_37_5 (.BL(BL5),.BLN(BLN5),.WL(WL37));
sram_cell_6t_5 inst_cell_37_6 (.BL(BL6),.BLN(BLN6),.WL(WL37));
sram_cell_6t_5 inst_cell_37_7 (.BL(BL7),.BLN(BLN7),.WL(WL37));
sram_cell_6t_5 inst_cell_37_8 (.BL(BL8),.BLN(BLN8),.WL(WL37));
sram_cell_6t_5 inst_cell_37_9 (.BL(BL9),.BLN(BLN9),.WL(WL37));
sram_cell_6t_5 inst_cell_37_10 (.BL(BL10),.BLN(BLN10),.WL(WL37));
sram_cell_6t_5 inst_cell_37_11 (.BL(BL11),.BLN(BLN11),.WL(WL37));
sram_cell_6t_5 inst_cell_37_12 (.BL(BL12),.BLN(BLN12),.WL(WL37));
sram_cell_6t_5 inst_cell_37_13 (.BL(BL13),.BLN(BLN13),.WL(WL37));
sram_cell_6t_5 inst_cell_37_14 (.BL(BL14),.BLN(BLN14),.WL(WL37));
sram_cell_6t_5 inst_cell_37_15 (.BL(BL15),.BLN(BLN15),.WL(WL37));
sram_cell_6t_5 inst_cell_37_16 (.BL(BL16),.BLN(BLN16),.WL(WL37));
sram_cell_6t_5 inst_cell_37_17 (.BL(BL17),.BLN(BLN17),.WL(WL37));
sram_cell_6t_5 inst_cell_37_18 (.BL(BL18),.BLN(BLN18),.WL(WL37));
sram_cell_6t_5 inst_cell_37_19 (.BL(BL19),.BLN(BLN19),.WL(WL37));
sram_cell_6t_5 inst_cell_37_20 (.BL(BL20),.BLN(BLN20),.WL(WL37));
sram_cell_6t_5 inst_cell_37_21 (.BL(BL21),.BLN(BLN21),.WL(WL37));
sram_cell_6t_5 inst_cell_37_22 (.BL(BL22),.BLN(BLN22),.WL(WL37));
sram_cell_6t_5 inst_cell_37_23 (.BL(BL23),.BLN(BLN23),.WL(WL37));
sram_cell_6t_5 inst_cell_37_24 (.BL(BL24),.BLN(BLN24),.WL(WL37));
sram_cell_6t_5 inst_cell_37_25 (.BL(BL25),.BLN(BLN25),.WL(WL37));
sram_cell_6t_5 inst_cell_37_26 (.BL(BL26),.BLN(BLN26),.WL(WL37));
sram_cell_6t_5 inst_cell_37_27 (.BL(BL27),.BLN(BLN27),.WL(WL37));
sram_cell_6t_5 inst_cell_37_28 (.BL(BL28),.BLN(BLN28),.WL(WL37));
sram_cell_6t_5 inst_cell_37_29 (.BL(BL29),.BLN(BLN29),.WL(WL37));
sram_cell_6t_5 inst_cell_37_30 (.BL(BL30),.BLN(BLN30),.WL(WL37));
sram_cell_6t_5 inst_cell_37_31 (.BL(BL31),.BLN(BLN31),.WL(WL37));
sram_cell_6t_5 inst_cell_37_32 (.BL(BL32),.BLN(BLN32),.WL(WL37));
sram_cell_6t_5 inst_cell_37_33 (.BL(BL33),.BLN(BLN33),.WL(WL37));
sram_cell_6t_5 inst_cell_37_34 (.BL(BL34),.BLN(BLN34),.WL(WL37));
sram_cell_6t_5 inst_cell_37_35 (.BL(BL35),.BLN(BLN35),.WL(WL37));
sram_cell_6t_5 inst_cell_37_36 (.BL(BL36),.BLN(BLN36),.WL(WL37));
sram_cell_6t_5 inst_cell_37_37 (.BL(BL37),.BLN(BLN37),.WL(WL37));
sram_cell_6t_5 inst_cell_37_38 (.BL(BL38),.BLN(BLN38),.WL(WL37));
sram_cell_6t_5 inst_cell_37_39 (.BL(BL39),.BLN(BLN39),.WL(WL37));
sram_cell_6t_5 inst_cell_37_40 (.BL(BL40),.BLN(BLN40),.WL(WL37));
sram_cell_6t_5 inst_cell_37_41 (.BL(BL41),.BLN(BLN41),.WL(WL37));
sram_cell_6t_5 inst_cell_37_42 (.BL(BL42),.BLN(BLN42),.WL(WL37));
sram_cell_6t_5 inst_cell_37_43 (.BL(BL43),.BLN(BLN43),.WL(WL37));
sram_cell_6t_5 inst_cell_37_44 (.BL(BL44),.BLN(BLN44),.WL(WL37));
sram_cell_6t_5 inst_cell_37_45 (.BL(BL45),.BLN(BLN45),.WL(WL37));
sram_cell_6t_5 inst_cell_37_46 (.BL(BL46),.BLN(BLN46),.WL(WL37));
sram_cell_6t_5 inst_cell_37_47 (.BL(BL47),.BLN(BLN47),.WL(WL37));
sram_cell_6t_5 inst_cell_37_48 (.BL(BL48),.BLN(BLN48),.WL(WL37));
sram_cell_6t_5 inst_cell_37_49 (.BL(BL49),.BLN(BLN49),.WL(WL37));
sram_cell_6t_5 inst_cell_37_50 (.BL(BL50),.BLN(BLN50),.WL(WL37));
sram_cell_6t_5 inst_cell_37_51 (.BL(BL51),.BLN(BLN51),.WL(WL37));
sram_cell_6t_5 inst_cell_37_52 (.BL(BL52),.BLN(BLN52),.WL(WL37));
sram_cell_6t_5 inst_cell_37_53 (.BL(BL53),.BLN(BLN53),.WL(WL37));
sram_cell_6t_5 inst_cell_37_54 (.BL(BL54),.BLN(BLN54),.WL(WL37));
sram_cell_6t_5 inst_cell_37_55 (.BL(BL55),.BLN(BLN55),.WL(WL37));
sram_cell_6t_5 inst_cell_37_56 (.BL(BL56),.BLN(BLN56),.WL(WL37));
sram_cell_6t_5 inst_cell_37_57 (.BL(BL57),.BLN(BLN57),.WL(WL37));
sram_cell_6t_5 inst_cell_37_58 (.BL(BL58),.BLN(BLN58),.WL(WL37));
sram_cell_6t_5 inst_cell_37_59 (.BL(BL59),.BLN(BLN59),.WL(WL37));
sram_cell_6t_5 inst_cell_37_60 (.BL(BL60),.BLN(BLN60),.WL(WL37));
sram_cell_6t_5 inst_cell_37_61 (.BL(BL61),.BLN(BLN61),.WL(WL37));
sram_cell_6t_5 inst_cell_37_62 (.BL(BL62),.BLN(BLN62),.WL(WL37));
sram_cell_6t_5 inst_cell_37_63 (.BL(BL63),.BLN(BLN63),.WL(WL37));
sram_cell_6t_5 inst_cell_37_64 (.BL(BL64),.BLN(BLN64),.WL(WL37));
sram_cell_6t_5 inst_cell_37_65 (.BL(BL65),.BLN(BLN65),.WL(WL37));
sram_cell_6t_5 inst_cell_37_66 (.BL(BL66),.BLN(BLN66),.WL(WL37));
sram_cell_6t_5 inst_cell_37_67 (.BL(BL67),.BLN(BLN67),.WL(WL37));
sram_cell_6t_5 inst_cell_37_68 (.BL(BL68),.BLN(BLN68),.WL(WL37));
sram_cell_6t_5 inst_cell_37_69 (.BL(BL69),.BLN(BLN69),.WL(WL37));
sram_cell_6t_5 inst_cell_37_70 (.BL(BL70),.BLN(BLN70),.WL(WL37));
sram_cell_6t_5 inst_cell_37_71 (.BL(BL71),.BLN(BLN71),.WL(WL37));
sram_cell_6t_5 inst_cell_37_72 (.BL(BL72),.BLN(BLN72),.WL(WL37));
sram_cell_6t_5 inst_cell_37_73 (.BL(BL73),.BLN(BLN73),.WL(WL37));
sram_cell_6t_5 inst_cell_37_74 (.BL(BL74),.BLN(BLN74),.WL(WL37));
sram_cell_6t_5 inst_cell_37_75 (.BL(BL75),.BLN(BLN75),.WL(WL37));
sram_cell_6t_5 inst_cell_37_76 (.BL(BL76),.BLN(BLN76),.WL(WL37));
sram_cell_6t_5 inst_cell_37_77 (.BL(BL77),.BLN(BLN77),.WL(WL37));
sram_cell_6t_5 inst_cell_37_78 (.BL(BL78),.BLN(BLN78),.WL(WL37));
sram_cell_6t_5 inst_cell_37_79 (.BL(BL79),.BLN(BLN79),.WL(WL37));
sram_cell_6t_5 inst_cell_37_80 (.BL(BL80),.BLN(BLN80),.WL(WL37));
sram_cell_6t_5 inst_cell_37_81 (.BL(BL81),.BLN(BLN81),.WL(WL37));
sram_cell_6t_5 inst_cell_37_82 (.BL(BL82),.BLN(BLN82),.WL(WL37));
sram_cell_6t_5 inst_cell_37_83 (.BL(BL83),.BLN(BLN83),.WL(WL37));
sram_cell_6t_5 inst_cell_37_84 (.BL(BL84),.BLN(BLN84),.WL(WL37));
sram_cell_6t_5 inst_cell_37_85 (.BL(BL85),.BLN(BLN85),.WL(WL37));
sram_cell_6t_5 inst_cell_37_86 (.BL(BL86),.BLN(BLN86),.WL(WL37));
sram_cell_6t_5 inst_cell_37_87 (.BL(BL87),.BLN(BLN87),.WL(WL37));
sram_cell_6t_5 inst_cell_37_88 (.BL(BL88),.BLN(BLN88),.WL(WL37));
sram_cell_6t_5 inst_cell_37_89 (.BL(BL89),.BLN(BLN89),.WL(WL37));
sram_cell_6t_5 inst_cell_37_90 (.BL(BL90),.BLN(BLN90),.WL(WL37));
sram_cell_6t_5 inst_cell_37_91 (.BL(BL91),.BLN(BLN91),.WL(WL37));
sram_cell_6t_5 inst_cell_37_92 (.BL(BL92),.BLN(BLN92),.WL(WL37));
sram_cell_6t_5 inst_cell_37_93 (.BL(BL93),.BLN(BLN93),.WL(WL37));
sram_cell_6t_5 inst_cell_37_94 (.BL(BL94),.BLN(BLN94),.WL(WL37));
sram_cell_6t_5 inst_cell_37_95 (.BL(BL95),.BLN(BLN95),.WL(WL37));
sram_cell_6t_5 inst_cell_37_96 (.BL(BL96),.BLN(BLN96),.WL(WL37));
sram_cell_6t_5 inst_cell_37_97 (.BL(BL97),.BLN(BLN97),.WL(WL37));
sram_cell_6t_5 inst_cell_37_98 (.BL(BL98),.BLN(BLN98),.WL(WL37));
sram_cell_6t_5 inst_cell_37_99 (.BL(BL99),.BLN(BLN99),.WL(WL37));
sram_cell_6t_5 inst_cell_37_100 (.BL(BL100),.BLN(BLN100),.WL(WL37));
sram_cell_6t_5 inst_cell_37_101 (.BL(BL101),.BLN(BLN101),.WL(WL37));
sram_cell_6t_5 inst_cell_37_102 (.BL(BL102),.BLN(BLN102),.WL(WL37));
sram_cell_6t_5 inst_cell_37_103 (.BL(BL103),.BLN(BLN103),.WL(WL37));
sram_cell_6t_5 inst_cell_37_104 (.BL(BL104),.BLN(BLN104),.WL(WL37));
sram_cell_6t_5 inst_cell_37_105 (.BL(BL105),.BLN(BLN105),.WL(WL37));
sram_cell_6t_5 inst_cell_37_106 (.BL(BL106),.BLN(BLN106),.WL(WL37));
sram_cell_6t_5 inst_cell_37_107 (.BL(BL107),.BLN(BLN107),.WL(WL37));
sram_cell_6t_5 inst_cell_37_108 (.BL(BL108),.BLN(BLN108),.WL(WL37));
sram_cell_6t_5 inst_cell_37_109 (.BL(BL109),.BLN(BLN109),.WL(WL37));
sram_cell_6t_5 inst_cell_37_110 (.BL(BL110),.BLN(BLN110),.WL(WL37));
sram_cell_6t_5 inst_cell_37_111 (.BL(BL111),.BLN(BLN111),.WL(WL37));
sram_cell_6t_5 inst_cell_37_112 (.BL(BL112),.BLN(BLN112),.WL(WL37));
sram_cell_6t_5 inst_cell_37_113 (.BL(BL113),.BLN(BLN113),.WL(WL37));
sram_cell_6t_5 inst_cell_37_114 (.BL(BL114),.BLN(BLN114),.WL(WL37));
sram_cell_6t_5 inst_cell_37_115 (.BL(BL115),.BLN(BLN115),.WL(WL37));
sram_cell_6t_5 inst_cell_37_116 (.BL(BL116),.BLN(BLN116),.WL(WL37));
sram_cell_6t_5 inst_cell_37_117 (.BL(BL117),.BLN(BLN117),.WL(WL37));
sram_cell_6t_5 inst_cell_37_118 (.BL(BL118),.BLN(BLN118),.WL(WL37));
sram_cell_6t_5 inst_cell_37_119 (.BL(BL119),.BLN(BLN119),.WL(WL37));
sram_cell_6t_5 inst_cell_37_120 (.BL(BL120),.BLN(BLN120),.WL(WL37));
sram_cell_6t_5 inst_cell_37_121 (.BL(BL121),.BLN(BLN121),.WL(WL37));
sram_cell_6t_5 inst_cell_37_122 (.BL(BL122),.BLN(BLN122),.WL(WL37));
sram_cell_6t_5 inst_cell_37_123 (.BL(BL123),.BLN(BLN123),.WL(WL37));
sram_cell_6t_5 inst_cell_37_124 (.BL(BL124),.BLN(BLN124),.WL(WL37));
sram_cell_6t_5 inst_cell_37_125 (.BL(BL125),.BLN(BLN125),.WL(WL37));
sram_cell_6t_5 inst_cell_37_126 (.BL(BL126),.BLN(BLN126),.WL(WL37));
sram_cell_6t_5 inst_cell_37_127 (.BL(BL127),.BLN(BLN127),.WL(WL37));
sram_cell_6t_5 inst_cell_38_0 (.BL(BL0),.BLN(BLN0),.WL(WL38));
sram_cell_6t_5 inst_cell_38_1 (.BL(BL1),.BLN(BLN1),.WL(WL38));
sram_cell_6t_5 inst_cell_38_2 (.BL(BL2),.BLN(BLN2),.WL(WL38));
sram_cell_6t_5 inst_cell_38_3 (.BL(BL3),.BLN(BLN3),.WL(WL38));
sram_cell_6t_5 inst_cell_38_4 (.BL(BL4),.BLN(BLN4),.WL(WL38));
sram_cell_6t_5 inst_cell_38_5 (.BL(BL5),.BLN(BLN5),.WL(WL38));
sram_cell_6t_5 inst_cell_38_6 (.BL(BL6),.BLN(BLN6),.WL(WL38));
sram_cell_6t_5 inst_cell_38_7 (.BL(BL7),.BLN(BLN7),.WL(WL38));
sram_cell_6t_5 inst_cell_38_8 (.BL(BL8),.BLN(BLN8),.WL(WL38));
sram_cell_6t_5 inst_cell_38_9 (.BL(BL9),.BLN(BLN9),.WL(WL38));
sram_cell_6t_5 inst_cell_38_10 (.BL(BL10),.BLN(BLN10),.WL(WL38));
sram_cell_6t_5 inst_cell_38_11 (.BL(BL11),.BLN(BLN11),.WL(WL38));
sram_cell_6t_5 inst_cell_38_12 (.BL(BL12),.BLN(BLN12),.WL(WL38));
sram_cell_6t_5 inst_cell_38_13 (.BL(BL13),.BLN(BLN13),.WL(WL38));
sram_cell_6t_5 inst_cell_38_14 (.BL(BL14),.BLN(BLN14),.WL(WL38));
sram_cell_6t_5 inst_cell_38_15 (.BL(BL15),.BLN(BLN15),.WL(WL38));
sram_cell_6t_5 inst_cell_38_16 (.BL(BL16),.BLN(BLN16),.WL(WL38));
sram_cell_6t_5 inst_cell_38_17 (.BL(BL17),.BLN(BLN17),.WL(WL38));
sram_cell_6t_5 inst_cell_38_18 (.BL(BL18),.BLN(BLN18),.WL(WL38));
sram_cell_6t_5 inst_cell_38_19 (.BL(BL19),.BLN(BLN19),.WL(WL38));
sram_cell_6t_5 inst_cell_38_20 (.BL(BL20),.BLN(BLN20),.WL(WL38));
sram_cell_6t_5 inst_cell_38_21 (.BL(BL21),.BLN(BLN21),.WL(WL38));
sram_cell_6t_5 inst_cell_38_22 (.BL(BL22),.BLN(BLN22),.WL(WL38));
sram_cell_6t_5 inst_cell_38_23 (.BL(BL23),.BLN(BLN23),.WL(WL38));
sram_cell_6t_5 inst_cell_38_24 (.BL(BL24),.BLN(BLN24),.WL(WL38));
sram_cell_6t_5 inst_cell_38_25 (.BL(BL25),.BLN(BLN25),.WL(WL38));
sram_cell_6t_5 inst_cell_38_26 (.BL(BL26),.BLN(BLN26),.WL(WL38));
sram_cell_6t_5 inst_cell_38_27 (.BL(BL27),.BLN(BLN27),.WL(WL38));
sram_cell_6t_5 inst_cell_38_28 (.BL(BL28),.BLN(BLN28),.WL(WL38));
sram_cell_6t_5 inst_cell_38_29 (.BL(BL29),.BLN(BLN29),.WL(WL38));
sram_cell_6t_5 inst_cell_38_30 (.BL(BL30),.BLN(BLN30),.WL(WL38));
sram_cell_6t_5 inst_cell_38_31 (.BL(BL31),.BLN(BLN31),.WL(WL38));
sram_cell_6t_5 inst_cell_38_32 (.BL(BL32),.BLN(BLN32),.WL(WL38));
sram_cell_6t_5 inst_cell_38_33 (.BL(BL33),.BLN(BLN33),.WL(WL38));
sram_cell_6t_5 inst_cell_38_34 (.BL(BL34),.BLN(BLN34),.WL(WL38));
sram_cell_6t_5 inst_cell_38_35 (.BL(BL35),.BLN(BLN35),.WL(WL38));
sram_cell_6t_5 inst_cell_38_36 (.BL(BL36),.BLN(BLN36),.WL(WL38));
sram_cell_6t_5 inst_cell_38_37 (.BL(BL37),.BLN(BLN37),.WL(WL38));
sram_cell_6t_5 inst_cell_38_38 (.BL(BL38),.BLN(BLN38),.WL(WL38));
sram_cell_6t_5 inst_cell_38_39 (.BL(BL39),.BLN(BLN39),.WL(WL38));
sram_cell_6t_5 inst_cell_38_40 (.BL(BL40),.BLN(BLN40),.WL(WL38));
sram_cell_6t_5 inst_cell_38_41 (.BL(BL41),.BLN(BLN41),.WL(WL38));
sram_cell_6t_5 inst_cell_38_42 (.BL(BL42),.BLN(BLN42),.WL(WL38));
sram_cell_6t_5 inst_cell_38_43 (.BL(BL43),.BLN(BLN43),.WL(WL38));
sram_cell_6t_5 inst_cell_38_44 (.BL(BL44),.BLN(BLN44),.WL(WL38));
sram_cell_6t_5 inst_cell_38_45 (.BL(BL45),.BLN(BLN45),.WL(WL38));
sram_cell_6t_5 inst_cell_38_46 (.BL(BL46),.BLN(BLN46),.WL(WL38));
sram_cell_6t_5 inst_cell_38_47 (.BL(BL47),.BLN(BLN47),.WL(WL38));
sram_cell_6t_5 inst_cell_38_48 (.BL(BL48),.BLN(BLN48),.WL(WL38));
sram_cell_6t_5 inst_cell_38_49 (.BL(BL49),.BLN(BLN49),.WL(WL38));
sram_cell_6t_5 inst_cell_38_50 (.BL(BL50),.BLN(BLN50),.WL(WL38));
sram_cell_6t_5 inst_cell_38_51 (.BL(BL51),.BLN(BLN51),.WL(WL38));
sram_cell_6t_5 inst_cell_38_52 (.BL(BL52),.BLN(BLN52),.WL(WL38));
sram_cell_6t_5 inst_cell_38_53 (.BL(BL53),.BLN(BLN53),.WL(WL38));
sram_cell_6t_5 inst_cell_38_54 (.BL(BL54),.BLN(BLN54),.WL(WL38));
sram_cell_6t_5 inst_cell_38_55 (.BL(BL55),.BLN(BLN55),.WL(WL38));
sram_cell_6t_5 inst_cell_38_56 (.BL(BL56),.BLN(BLN56),.WL(WL38));
sram_cell_6t_5 inst_cell_38_57 (.BL(BL57),.BLN(BLN57),.WL(WL38));
sram_cell_6t_5 inst_cell_38_58 (.BL(BL58),.BLN(BLN58),.WL(WL38));
sram_cell_6t_5 inst_cell_38_59 (.BL(BL59),.BLN(BLN59),.WL(WL38));
sram_cell_6t_5 inst_cell_38_60 (.BL(BL60),.BLN(BLN60),.WL(WL38));
sram_cell_6t_5 inst_cell_38_61 (.BL(BL61),.BLN(BLN61),.WL(WL38));
sram_cell_6t_5 inst_cell_38_62 (.BL(BL62),.BLN(BLN62),.WL(WL38));
sram_cell_6t_5 inst_cell_38_63 (.BL(BL63),.BLN(BLN63),.WL(WL38));
sram_cell_6t_5 inst_cell_38_64 (.BL(BL64),.BLN(BLN64),.WL(WL38));
sram_cell_6t_5 inst_cell_38_65 (.BL(BL65),.BLN(BLN65),.WL(WL38));
sram_cell_6t_5 inst_cell_38_66 (.BL(BL66),.BLN(BLN66),.WL(WL38));
sram_cell_6t_5 inst_cell_38_67 (.BL(BL67),.BLN(BLN67),.WL(WL38));
sram_cell_6t_5 inst_cell_38_68 (.BL(BL68),.BLN(BLN68),.WL(WL38));
sram_cell_6t_5 inst_cell_38_69 (.BL(BL69),.BLN(BLN69),.WL(WL38));
sram_cell_6t_5 inst_cell_38_70 (.BL(BL70),.BLN(BLN70),.WL(WL38));
sram_cell_6t_5 inst_cell_38_71 (.BL(BL71),.BLN(BLN71),.WL(WL38));
sram_cell_6t_5 inst_cell_38_72 (.BL(BL72),.BLN(BLN72),.WL(WL38));
sram_cell_6t_5 inst_cell_38_73 (.BL(BL73),.BLN(BLN73),.WL(WL38));
sram_cell_6t_5 inst_cell_38_74 (.BL(BL74),.BLN(BLN74),.WL(WL38));
sram_cell_6t_5 inst_cell_38_75 (.BL(BL75),.BLN(BLN75),.WL(WL38));
sram_cell_6t_5 inst_cell_38_76 (.BL(BL76),.BLN(BLN76),.WL(WL38));
sram_cell_6t_5 inst_cell_38_77 (.BL(BL77),.BLN(BLN77),.WL(WL38));
sram_cell_6t_5 inst_cell_38_78 (.BL(BL78),.BLN(BLN78),.WL(WL38));
sram_cell_6t_5 inst_cell_38_79 (.BL(BL79),.BLN(BLN79),.WL(WL38));
sram_cell_6t_5 inst_cell_38_80 (.BL(BL80),.BLN(BLN80),.WL(WL38));
sram_cell_6t_5 inst_cell_38_81 (.BL(BL81),.BLN(BLN81),.WL(WL38));
sram_cell_6t_5 inst_cell_38_82 (.BL(BL82),.BLN(BLN82),.WL(WL38));
sram_cell_6t_5 inst_cell_38_83 (.BL(BL83),.BLN(BLN83),.WL(WL38));
sram_cell_6t_5 inst_cell_38_84 (.BL(BL84),.BLN(BLN84),.WL(WL38));
sram_cell_6t_5 inst_cell_38_85 (.BL(BL85),.BLN(BLN85),.WL(WL38));
sram_cell_6t_5 inst_cell_38_86 (.BL(BL86),.BLN(BLN86),.WL(WL38));
sram_cell_6t_5 inst_cell_38_87 (.BL(BL87),.BLN(BLN87),.WL(WL38));
sram_cell_6t_5 inst_cell_38_88 (.BL(BL88),.BLN(BLN88),.WL(WL38));
sram_cell_6t_5 inst_cell_38_89 (.BL(BL89),.BLN(BLN89),.WL(WL38));
sram_cell_6t_5 inst_cell_38_90 (.BL(BL90),.BLN(BLN90),.WL(WL38));
sram_cell_6t_5 inst_cell_38_91 (.BL(BL91),.BLN(BLN91),.WL(WL38));
sram_cell_6t_5 inst_cell_38_92 (.BL(BL92),.BLN(BLN92),.WL(WL38));
sram_cell_6t_5 inst_cell_38_93 (.BL(BL93),.BLN(BLN93),.WL(WL38));
sram_cell_6t_5 inst_cell_38_94 (.BL(BL94),.BLN(BLN94),.WL(WL38));
sram_cell_6t_5 inst_cell_38_95 (.BL(BL95),.BLN(BLN95),.WL(WL38));
sram_cell_6t_5 inst_cell_38_96 (.BL(BL96),.BLN(BLN96),.WL(WL38));
sram_cell_6t_5 inst_cell_38_97 (.BL(BL97),.BLN(BLN97),.WL(WL38));
sram_cell_6t_5 inst_cell_38_98 (.BL(BL98),.BLN(BLN98),.WL(WL38));
sram_cell_6t_5 inst_cell_38_99 (.BL(BL99),.BLN(BLN99),.WL(WL38));
sram_cell_6t_5 inst_cell_38_100 (.BL(BL100),.BLN(BLN100),.WL(WL38));
sram_cell_6t_5 inst_cell_38_101 (.BL(BL101),.BLN(BLN101),.WL(WL38));
sram_cell_6t_5 inst_cell_38_102 (.BL(BL102),.BLN(BLN102),.WL(WL38));
sram_cell_6t_5 inst_cell_38_103 (.BL(BL103),.BLN(BLN103),.WL(WL38));
sram_cell_6t_5 inst_cell_38_104 (.BL(BL104),.BLN(BLN104),.WL(WL38));
sram_cell_6t_5 inst_cell_38_105 (.BL(BL105),.BLN(BLN105),.WL(WL38));
sram_cell_6t_5 inst_cell_38_106 (.BL(BL106),.BLN(BLN106),.WL(WL38));
sram_cell_6t_5 inst_cell_38_107 (.BL(BL107),.BLN(BLN107),.WL(WL38));
sram_cell_6t_5 inst_cell_38_108 (.BL(BL108),.BLN(BLN108),.WL(WL38));
sram_cell_6t_5 inst_cell_38_109 (.BL(BL109),.BLN(BLN109),.WL(WL38));
sram_cell_6t_5 inst_cell_38_110 (.BL(BL110),.BLN(BLN110),.WL(WL38));
sram_cell_6t_5 inst_cell_38_111 (.BL(BL111),.BLN(BLN111),.WL(WL38));
sram_cell_6t_5 inst_cell_38_112 (.BL(BL112),.BLN(BLN112),.WL(WL38));
sram_cell_6t_5 inst_cell_38_113 (.BL(BL113),.BLN(BLN113),.WL(WL38));
sram_cell_6t_5 inst_cell_38_114 (.BL(BL114),.BLN(BLN114),.WL(WL38));
sram_cell_6t_5 inst_cell_38_115 (.BL(BL115),.BLN(BLN115),.WL(WL38));
sram_cell_6t_5 inst_cell_38_116 (.BL(BL116),.BLN(BLN116),.WL(WL38));
sram_cell_6t_5 inst_cell_38_117 (.BL(BL117),.BLN(BLN117),.WL(WL38));
sram_cell_6t_5 inst_cell_38_118 (.BL(BL118),.BLN(BLN118),.WL(WL38));
sram_cell_6t_5 inst_cell_38_119 (.BL(BL119),.BLN(BLN119),.WL(WL38));
sram_cell_6t_5 inst_cell_38_120 (.BL(BL120),.BLN(BLN120),.WL(WL38));
sram_cell_6t_5 inst_cell_38_121 (.BL(BL121),.BLN(BLN121),.WL(WL38));
sram_cell_6t_5 inst_cell_38_122 (.BL(BL122),.BLN(BLN122),.WL(WL38));
sram_cell_6t_5 inst_cell_38_123 (.BL(BL123),.BLN(BLN123),.WL(WL38));
sram_cell_6t_5 inst_cell_38_124 (.BL(BL124),.BLN(BLN124),.WL(WL38));
sram_cell_6t_5 inst_cell_38_125 (.BL(BL125),.BLN(BLN125),.WL(WL38));
sram_cell_6t_5 inst_cell_38_126 (.BL(BL126),.BLN(BLN126),.WL(WL38));
sram_cell_6t_5 inst_cell_38_127 (.BL(BL127),.BLN(BLN127),.WL(WL38));
sram_cell_6t_5 inst_cell_39_0 (.BL(BL0),.BLN(BLN0),.WL(WL39));
sram_cell_6t_5 inst_cell_39_1 (.BL(BL1),.BLN(BLN1),.WL(WL39));
sram_cell_6t_5 inst_cell_39_2 (.BL(BL2),.BLN(BLN2),.WL(WL39));
sram_cell_6t_5 inst_cell_39_3 (.BL(BL3),.BLN(BLN3),.WL(WL39));
sram_cell_6t_5 inst_cell_39_4 (.BL(BL4),.BLN(BLN4),.WL(WL39));
sram_cell_6t_5 inst_cell_39_5 (.BL(BL5),.BLN(BLN5),.WL(WL39));
sram_cell_6t_5 inst_cell_39_6 (.BL(BL6),.BLN(BLN6),.WL(WL39));
sram_cell_6t_5 inst_cell_39_7 (.BL(BL7),.BLN(BLN7),.WL(WL39));
sram_cell_6t_5 inst_cell_39_8 (.BL(BL8),.BLN(BLN8),.WL(WL39));
sram_cell_6t_5 inst_cell_39_9 (.BL(BL9),.BLN(BLN9),.WL(WL39));
sram_cell_6t_5 inst_cell_39_10 (.BL(BL10),.BLN(BLN10),.WL(WL39));
sram_cell_6t_5 inst_cell_39_11 (.BL(BL11),.BLN(BLN11),.WL(WL39));
sram_cell_6t_5 inst_cell_39_12 (.BL(BL12),.BLN(BLN12),.WL(WL39));
sram_cell_6t_5 inst_cell_39_13 (.BL(BL13),.BLN(BLN13),.WL(WL39));
sram_cell_6t_5 inst_cell_39_14 (.BL(BL14),.BLN(BLN14),.WL(WL39));
sram_cell_6t_5 inst_cell_39_15 (.BL(BL15),.BLN(BLN15),.WL(WL39));
sram_cell_6t_5 inst_cell_39_16 (.BL(BL16),.BLN(BLN16),.WL(WL39));
sram_cell_6t_5 inst_cell_39_17 (.BL(BL17),.BLN(BLN17),.WL(WL39));
sram_cell_6t_5 inst_cell_39_18 (.BL(BL18),.BLN(BLN18),.WL(WL39));
sram_cell_6t_5 inst_cell_39_19 (.BL(BL19),.BLN(BLN19),.WL(WL39));
sram_cell_6t_5 inst_cell_39_20 (.BL(BL20),.BLN(BLN20),.WL(WL39));
sram_cell_6t_5 inst_cell_39_21 (.BL(BL21),.BLN(BLN21),.WL(WL39));
sram_cell_6t_5 inst_cell_39_22 (.BL(BL22),.BLN(BLN22),.WL(WL39));
sram_cell_6t_5 inst_cell_39_23 (.BL(BL23),.BLN(BLN23),.WL(WL39));
sram_cell_6t_5 inst_cell_39_24 (.BL(BL24),.BLN(BLN24),.WL(WL39));
sram_cell_6t_5 inst_cell_39_25 (.BL(BL25),.BLN(BLN25),.WL(WL39));
sram_cell_6t_5 inst_cell_39_26 (.BL(BL26),.BLN(BLN26),.WL(WL39));
sram_cell_6t_5 inst_cell_39_27 (.BL(BL27),.BLN(BLN27),.WL(WL39));
sram_cell_6t_5 inst_cell_39_28 (.BL(BL28),.BLN(BLN28),.WL(WL39));
sram_cell_6t_5 inst_cell_39_29 (.BL(BL29),.BLN(BLN29),.WL(WL39));
sram_cell_6t_5 inst_cell_39_30 (.BL(BL30),.BLN(BLN30),.WL(WL39));
sram_cell_6t_5 inst_cell_39_31 (.BL(BL31),.BLN(BLN31),.WL(WL39));
sram_cell_6t_5 inst_cell_39_32 (.BL(BL32),.BLN(BLN32),.WL(WL39));
sram_cell_6t_5 inst_cell_39_33 (.BL(BL33),.BLN(BLN33),.WL(WL39));
sram_cell_6t_5 inst_cell_39_34 (.BL(BL34),.BLN(BLN34),.WL(WL39));
sram_cell_6t_5 inst_cell_39_35 (.BL(BL35),.BLN(BLN35),.WL(WL39));
sram_cell_6t_5 inst_cell_39_36 (.BL(BL36),.BLN(BLN36),.WL(WL39));
sram_cell_6t_5 inst_cell_39_37 (.BL(BL37),.BLN(BLN37),.WL(WL39));
sram_cell_6t_5 inst_cell_39_38 (.BL(BL38),.BLN(BLN38),.WL(WL39));
sram_cell_6t_5 inst_cell_39_39 (.BL(BL39),.BLN(BLN39),.WL(WL39));
sram_cell_6t_5 inst_cell_39_40 (.BL(BL40),.BLN(BLN40),.WL(WL39));
sram_cell_6t_5 inst_cell_39_41 (.BL(BL41),.BLN(BLN41),.WL(WL39));
sram_cell_6t_5 inst_cell_39_42 (.BL(BL42),.BLN(BLN42),.WL(WL39));
sram_cell_6t_5 inst_cell_39_43 (.BL(BL43),.BLN(BLN43),.WL(WL39));
sram_cell_6t_5 inst_cell_39_44 (.BL(BL44),.BLN(BLN44),.WL(WL39));
sram_cell_6t_5 inst_cell_39_45 (.BL(BL45),.BLN(BLN45),.WL(WL39));
sram_cell_6t_5 inst_cell_39_46 (.BL(BL46),.BLN(BLN46),.WL(WL39));
sram_cell_6t_5 inst_cell_39_47 (.BL(BL47),.BLN(BLN47),.WL(WL39));
sram_cell_6t_5 inst_cell_39_48 (.BL(BL48),.BLN(BLN48),.WL(WL39));
sram_cell_6t_5 inst_cell_39_49 (.BL(BL49),.BLN(BLN49),.WL(WL39));
sram_cell_6t_5 inst_cell_39_50 (.BL(BL50),.BLN(BLN50),.WL(WL39));
sram_cell_6t_5 inst_cell_39_51 (.BL(BL51),.BLN(BLN51),.WL(WL39));
sram_cell_6t_5 inst_cell_39_52 (.BL(BL52),.BLN(BLN52),.WL(WL39));
sram_cell_6t_5 inst_cell_39_53 (.BL(BL53),.BLN(BLN53),.WL(WL39));
sram_cell_6t_5 inst_cell_39_54 (.BL(BL54),.BLN(BLN54),.WL(WL39));
sram_cell_6t_5 inst_cell_39_55 (.BL(BL55),.BLN(BLN55),.WL(WL39));
sram_cell_6t_5 inst_cell_39_56 (.BL(BL56),.BLN(BLN56),.WL(WL39));
sram_cell_6t_5 inst_cell_39_57 (.BL(BL57),.BLN(BLN57),.WL(WL39));
sram_cell_6t_5 inst_cell_39_58 (.BL(BL58),.BLN(BLN58),.WL(WL39));
sram_cell_6t_5 inst_cell_39_59 (.BL(BL59),.BLN(BLN59),.WL(WL39));
sram_cell_6t_5 inst_cell_39_60 (.BL(BL60),.BLN(BLN60),.WL(WL39));
sram_cell_6t_5 inst_cell_39_61 (.BL(BL61),.BLN(BLN61),.WL(WL39));
sram_cell_6t_5 inst_cell_39_62 (.BL(BL62),.BLN(BLN62),.WL(WL39));
sram_cell_6t_5 inst_cell_39_63 (.BL(BL63),.BLN(BLN63),.WL(WL39));
sram_cell_6t_5 inst_cell_39_64 (.BL(BL64),.BLN(BLN64),.WL(WL39));
sram_cell_6t_5 inst_cell_39_65 (.BL(BL65),.BLN(BLN65),.WL(WL39));
sram_cell_6t_5 inst_cell_39_66 (.BL(BL66),.BLN(BLN66),.WL(WL39));
sram_cell_6t_5 inst_cell_39_67 (.BL(BL67),.BLN(BLN67),.WL(WL39));
sram_cell_6t_5 inst_cell_39_68 (.BL(BL68),.BLN(BLN68),.WL(WL39));
sram_cell_6t_5 inst_cell_39_69 (.BL(BL69),.BLN(BLN69),.WL(WL39));
sram_cell_6t_5 inst_cell_39_70 (.BL(BL70),.BLN(BLN70),.WL(WL39));
sram_cell_6t_5 inst_cell_39_71 (.BL(BL71),.BLN(BLN71),.WL(WL39));
sram_cell_6t_5 inst_cell_39_72 (.BL(BL72),.BLN(BLN72),.WL(WL39));
sram_cell_6t_5 inst_cell_39_73 (.BL(BL73),.BLN(BLN73),.WL(WL39));
sram_cell_6t_5 inst_cell_39_74 (.BL(BL74),.BLN(BLN74),.WL(WL39));
sram_cell_6t_5 inst_cell_39_75 (.BL(BL75),.BLN(BLN75),.WL(WL39));
sram_cell_6t_5 inst_cell_39_76 (.BL(BL76),.BLN(BLN76),.WL(WL39));
sram_cell_6t_5 inst_cell_39_77 (.BL(BL77),.BLN(BLN77),.WL(WL39));
sram_cell_6t_5 inst_cell_39_78 (.BL(BL78),.BLN(BLN78),.WL(WL39));
sram_cell_6t_5 inst_cell_39_79 (.BL(BL79),.BLN(BLN79),.WL(WL39));
sram_cell_6t_5 inst_cell_39_80 (.BL(BL80),.BLN(BLN80),.WL(WL39));
sram_cell_6t_5 inst_cell_39_81 (.BL(BL81),.BLN(BLN81),.WL(WL39));
sram_cell_6t_5 inst_cell_39_82 (.BL(BL82),.BLN(BLN82),.WL(WL39));
sram_cell_6t_5 inst_cell_39_83 (.BL(BL83),.BLN(BLN83),.WL(WL39));
sram_cell_6t_5 inst_cell_39_84 (.BL(BL84),.BLN(BLN84),.WL(WL39));
sram_cell_6t_5 inst_cell_39_85 (.BL(BL85),.BLN(BLN85),.WL(WL39));
sram_cell_6t_5 inst_cell_39_86 (.BL(BL86),.BLN(BLN86),.WL(WL39));
sram_cell_6t_5 inst_cell_39_87 (.BL(BL87),.BLN(BLN87),.WL(WL39));
sram_cell_6t_5 inst_cell_39_88 (.BL(BL88),.BLN(BLN88),.WL(WL39));
sram_cell_6t_5 inst_cell_39_89 (.BL(BL89),.BLN(BLN89),.WL(WL39));
sram_cell_6t_5 inst_cell_39_90 (.BL(BL90),.BLN(BLN90),.WL(WL39));
sram_cell_6t_5 inst_cell_39_91 (.BL(BL91),.BLN(BLN91),.WL(WL39));
sram_cell_6t_5 inst_cell_39_92 (.BL(BL92),.BLN(BLN92),.WL(WL39));
sram_cell_6t_5 inst_cell_39_93 (.BL(BL93),.BLN(BLN93),.WL(WL39));
sram_cell_6t_5 inst_cell_39_94 (.BL(BL94),.BLN(BLN94),.WL(WL39));
sram_cell_6t_5 inst_cell_39_95 (.BL(BL95),.BLN(BLN95),.WL(WL39));
sram_cell_6t_5 inst_cell_39_96 (.BL(BL96),.BLN(BLN96),.WL(WL39));
sram_cell_6t_5 inst_cell_39_97 (.BL(BL97),.BLN(BLN97),.WL(WL39));
sram_cell_6t_5 inst_cell_39_98 (.BL(BL98),.BLN(BLN98),.WL(WL39));
sram_cell_6t_5 inst_cell_39_99 (.BL(BL99),.BLN(BLN99),.WL(WL39));
sram_cell_6t_5 inst_cell_39_100 (.BL(BL100),.BLN(BLN100),.WL(WL39));
sram_cell_6t_5 inst_cell_39_101 (.BL(BL101),.BLN(BLN101),.WL(WL39));
sram_cell_6t_5 inst_cell_39_102 (.BL(BL102),.BLN(BLN102),.WL(WL39));
sram_cell_6t_5 inst_cell_39_103 (.BL(BL103),.BLN(BLN103),.WL(WL39));
sram_cell_6t_5 inst_cell_39_104 (.BL(BL104),.BLN(BLN104),.WL(WL39));
sram_cell_6t_5 inst_cell_39_105 (.BL(BL105),.BLN(BLN105),.WL(WL39));
sram_cell_6t_5 inst_cell_39_106 (.BL(BL106),.BLN(BLN106),.WL(WL39));
sram_cell_6t_5 inst_cell_39_107 (.BL(BL107),.BLN(BLN107),.WL(WL39));
sram_cell_6t_5 inst_cell_39_108 (.BL(BL108),.BLN(BLN108),.WL(WL39));
sram_cell_6t_5 inst_cell_39_109 (.BL(BL109),.BLN(BLN109),.WL(WL39));
sram_cell_6t_5 inst_cell_39_110 (.BL(BL110),.BLN(BLN110),.WL(WL39));
sram_cell_6t_5 inst_cell_39_111 (.BL(BL111),.BLN(BLN111),.WL(WL39));
sram_cell_6t_5 inst_cell_39_112 (.BL(BL112),.BLN(BLN112),.WL(WL39));
sram_cell_6t_5 inst_cell_39_113 (.BL(BL113),.BLN(BLN113),.WL(WL39));
sram_cell_6t_5 inst_cell_39_114 (.BL(BL114),.BLN(BLN114),.WL(WL39));
sram_cell_6t_5 inst_cell_39_115 (.BL(BL115),.BLN(BLN115),.WL(WL39));
sram_cell_6t_5 inst_cell_39_116 (.BL(BL116),.BLN(BLN116),.WL(WL39));
sram_cell_6t_5 inst_cell_39_117 (.BL(BL117),.BLN(BLN117),.WL(WL39));
sram_cell_6t_5 inst_cell_39_118 (.BL(BL118),.BLN(BLN118),.WL(WL39));
sram_cell_6t_5 inst_cell_39_119 (.BL(BL119),.BLN(BLN119),.WL(WL39));
sram_cell_6t_5 inst_cell_39_120 (.BL(BL120),.BLN(BLN120),.WL(WL39));
sram_cell_6t_5 inst_cell_39_121 (.BL(BL121),.BLN(BLN121),.WL(WL39));
sram_cell_6t_5 inst_cell_39_122 (.BL(BL122),.BLN(BLN122),.WL(WL39));
sram_cell_6t_5 inst_cell_39_123 (.BL(BL123),.BLN(BLN123),.WL(WL39));
sram_cell_6t_5 inst_cell_39_124 (.BL(BL124),.BLN(BLN124),.WL(WL39));
sram_cell_6t_5 inst_cell_39_125 (.BL(BL125),.BLN(BLN125),.WL(WL39));
sram_cell_6t_5 inst_cell_39_126 (.BL(BL126),.BLN(BLN126),.WL(WL39));
sram_cell_6t_5 inst_cell_39_127 (.BL(BL127),.BLN(BLN127),.WL(WL39));
sram_cell_6t_5 inst_cell_40_0 (.BL(BL0),.BLN(BLN0),.WL(WL40));
sram_cell_6t_5 inst_cell_40_1 (.BL(BL1),.BLN(BLN1),.WL(WL40));
sram_cell_6t_5 inst_cell_40_2 (.BL(BL2),.BLN(BLN2),.WL(WL40));
sram_cell_6t_5 inst_cell_40_3 (.BL(BL3),.BLN(BLN3),.WL(WL40));
sram_cell_6t_5 inst_cell_40_4 (.BL(BL4),.BLN(BLN4),.WL(WL40));
sram_cell_6t_5 inst_cell_40_5 (.BL(BL5),.BLN(BLN5),.WL(WL40));
sram_cell_6t_5 inst_cell_40_6 (.BL(BL6),.BLN(BLN6),.WL(WL40));
sram_cell_6t_5 inst_cell_40_7 (.BL(BL7),.BLN(BLN7),.WL(WL40));
sram_cell_6t_5 inst_cell_40_8 (.BL(BL8),.BLN(BLN8),.WL(WL40));
sram_cell_6t_5 inst_cell_40_9 (.BL(BL9),.BLN(BLN9),.WL(WL40));
sram_cell_6t_5 inst_cell_40_10 (.BL(BL10),.BLN(BLN10),.WL(WL40));
sram_cell_6t_5 inst_cell_40_11 (.BL(BL11),.BLN(BLN11),.WL(WL40));
sram_cell_6t_5 inst_cell_40_12 (.BL(BL12),.BLN(BLN12),.WL(WL40));
sram_cell_6t_5 inst_cell_40_13 (.BL(BL13),.BLN(BLN13),.WL(WL40));
sram_cell_6t_5 inst_cell_40_14 (.BL(BL14),.BLN(BLN14),.WL(WL40));
sram_cell_6t_5 inst_cell_40_15 (.BL(BL15),.BLN(BLN15),.WL(WL40));
sram_cell_6t_5 inst_cell_40_16 (.BL(BL16),.BLN(BLN16),.WL(WL40));
sram_cell_6t_5 inst_cell_40_17 (.BL(BL17),.BLN(BLN17),.WL(WL40));
sram_cell_6t_5 inst_cell_40_18 (.BL(BL18),.BLN(BLN18),.WL(WL40));
sram_cell_6t_5 inst_cell_40_19 (.BL(BL19),.BLN(BLN19),.WL(WL40));
sram_cell_6t_5 inst_cell_40_20 (.BL(BL20),.BLN(BLN20),.WL(WL40));
sram_cell_6t_5 inst_cell_40_21 (.BL(BL21),.BLN(BLN21),.WL(WL40));
sram_cell_6t_5 inst_cell_40_22 (.BL(BL22),.BLN(BLN22),.WL(WL40));
sram_cell_6t_5 inst_cell_40_23 (.BL(BL23),.BLN(BLN23),.WL(WL40));
sram_cell_6t_5 inst_cell_40_24 (.BL(BL24),.BLN(BLN24),.WL(WL40));
sram_cell_6t_5 inst_cell_40_25 (.BL(BL25),.BLN(BLN25),.WL(WL40));
sram_cell_6t_5 inst_cell_40_26 (.BL(BL26),.BLN(BLN26),.WL(WL40));
sram_cell_6t_5 inst_cell_40_27 (.BL(BL27),.BLN(BLN27),.WL(WL40));
sram_cell_6t_5 inst_cell_40_28 (.BL(BL28),.BLN(BLN28),.WL(WL40));
sram_cell_6t_5 inst_cell_40_29 (.BL(BL29),.BLN(BLN29),.WL(WL40));
sram_cell_6t_5 inst_cell_40_30 (.BL(BL30),.BLN(BLN30),.WL(WL40));
sram_cell_6t_5 inst_cell_40_31 (.BL(BL31),.BLN(BLN31),.WL(WL40));
sram_cell_6t_5 inst_cell_40_32 (.BL(BL32),.BLN(BLN32),.WL(WL40));
sram_cell_6t_5 inst_cell_40_33 (.BL(BL33),.BLN(BLN33),.WL(WL40));
sram_cell_6t_5 inst_cell_40_34 (.BL(BL34),.BLN(BLN34),.WL(WL40));
sram_cell_6t_5 inst_cell_40_35 (.BL(BL35),.BLN(BLN35),.WL(WL40));
sram_cell_6t_5 inst_cell_40_36 (.BL(BL36),.BLN(BLN36),.WL(WL40));
sram_cell_6t_5 inst_cell_40_37 (.BL(BL37),.BLN(BLN37),.WL(WL40));
sram_cell_6t_5 inst_cell_40_38 (.BL(BL38),.BLN(BLN38),.WL(WL40));
sram_cell_6t_5 inst_cell_40_39 (.BL(BL39),.BLN(BLN39),.WL(WL40));
sram_cell_6t_5 inst_cell_40_40 (.BL(BL40),.BLN(BLN40),.WL(WL40));
sram_cell_6t_5 inst_cell_40_41 (.BL(BL41),.BLN(BLN41),.WL(WL40));
sram_cell_6t_5 inst_cell_40_42 (.BL(BL42),.BLN(BLN42),.WL(WL40));
sram_cell_6t_5 inst_cell_40_43 (.BL(BL43),.BLN(BLN43),.WL(WL40));
sram_cell_6t_5 inst_cell_40_44 (.BL(BL44),.BLN(BLN44),.WL(WL40));
sram_cell_6t_5 inst_cell_40_45 (.BL(BL45),.BLN(BLN45),.WL(WL40));
sram_cell_6t_5 inst_cell_40_46 (.BL(BL46),.BLN(BLN46),.WL(WL40));
sram_cell_6t_5 inst_cell_40_47 (.BL(BL47),.BLN(BLN47),.WL(WL40));
sram_cell_6t_5 inst_cell_40_48 (.BL(BL48),.BLN(BLN48),.WL(WL40));
sram_cell_6t_5 inst_cell_40_49 (.BL(BL49),.BLN(BLN49),.WL(WL40));
sram_cell_6t_5 inst_cell_40_50 (.BL(BL50),.BLN(BLN50),.WL(WL40));
sram_cell_6t_5 inst_cell_40_51 (.BL(BL51),.BLN(BLN51),.WL(WL40));
sram_cell_6t_5 inst_cell_40_52 (.BL(BL52),.BLN(BLN52),.WL(WL40));
sram_cell_6t_5 inst_cell_40_53 (.BL(BL53),.BLN(BLN53),.WL(WL40));
sram_cell_6t_5 inst_cell_40_54 (.BL(BL54),.BLN(BLN54),.WL(WL40));
sram_cell_6t_5 inst_cell_40_55 (.BL(BL55),.BLN(BLN55),.WL(WL40));
sram_cell_6t_5 inst_cell_40_56 (.BL(BL56),.BLN(BLN56),.WL(WL40));
sram_cell_6t_5 inst_cell_40_57 (.BL(BL57),.BLN(BLN57),.WL(WL40));
sram_cell_6t_5 inst_cell_40_58 (.BL(BL58),.BLN(BLN58),.WL(WL40));
sram_cell_6t_5 inst_cell_40_59 (.BL(BL59),.BLN(BLN59),.WL(WL40));
sram_cell_6t_5 inst_cell_40_60 (.BL(BL60),.BLN(BLN60),.WL(WL40));
sram_cell_6t_5 inst_cell_40_61 (.BL(BL61),.BLN(BLN61),.WL(WL40));
sram_cell_6t_5 inst_cell_40_62 (.BL(BL62),.BLN(BLN62),.WL(WL40));
sram_cell_6t_5 inst_cell_40_63 (.BL(BL63),.BLN(BLN63),.WL(WL40));
sram_cell_6t_5 inst_cell_40_64 (.BL(BL64),.BLN(BLN64),.WL(WL40));
sram_cell_6t_5 inst_cell_40_65 (.BL(BL65),.BLN(BLN65),.WL(WL40));
sram_cell_6t_5 inst_cell_40_66 (.BL(BL66),.BLN(BLN66),.WL(WL40));
sram_cell_6t_5 inst_cell_40_67 (.BL(BL67),.BLN(BLN67),.WL(WL40));
sram_cell_6t_5 inst_cell_40_68 (.BL(BL68),.BLN(BLN68),.WL(WL40));
sram_cell_6t_5 inst_cell_40_69 (.BL(BL69),.BLN(BLN69),.WL(WL40));
sram_cell_6t_5 inst_cell_40_70 (.BL(BL70),.BLN(BLN70),.WL(WL40));
sram_cell_6t_5 inst_cell_40_71 (.BL(BL71),.BLN(BLN71),.WL(WL40));
sram_cell_6t_5 inst_cell_40_72 (.BL(BL72),.BLN(BLN72),.WL(WL40));
sram_cell_6t_5 inst_cell_40_73 (.BL(BL73),.BLN(BLN73),.WL(WL40));
sram_cell_6t_5 inst_cell_40_74 (.BL(BL74),.BLN(BLN74),.WL(WL40));
sram_cell_6t_5 inst_cell_40_75 (.BL(BL75),.BLN(BLN75),.WL(WL40));
sram_cell_6t_5 inst_cell_40_76 (.BL(BL76),.BLN(BLN76),.WL(WL40));
sram_cell_6t_5 inst_cell_40_77 (.BL(BL77),.BLN(BLN77),.WL(WL40));
sram_cell_6t_5 inst_cell_40_78 (.BL(BL78),.BLN(BLN78),.WL(WL40));
sram_cell_6t_5 inst_cell_40_79 (.BL(BL79),.BLN(BLN79),.WL(WL40));
sram_cell_6t_5 inst_cell_40_80 (.BL(BL80),.BLN(BLN80),.WL(WL40));
sram_cell_6t_5 inst_cell_40_81 (.BL(BL81),.BLN(BLN81),.WL(WL40));
sram_cell_6t_5 inst_cell_40_82 (.BL(BL82),.BLN(BLN82),.WL(WL40));
sram_cell_6t_5 inst_cell_40_83 (.BL(BL83),.BLN(BLN83),.WL(WL40));
sram_cell_6t_5 inst_cell_40_84 (.BL(BL84),.BLN(BLN84),.WL(WL40));
sram_cell_6t_5 inst_cell_40_85 (.BL(BL85),.BLN(BLN85),.WL(WL40));
sram_cell_6t_5 inst_cell_40_86 (.BL(BL86),.BLN(BLN86),.WL(WL40));
sram_cell_6t_5 inst_cell_40_87 (.BL(BL87),.BLN(BLN87),.WL(WL40));
sram_cell_6t_5 inst_cell_40_88 (.BL(BL88),.BLN(BLN88),.WL(WL40));
sram_cell_6t_5 inst_cell_40_89 (.BL(BL89),.BLN(BLN89),.WL(WL40));
sram_cell_6t_5 inst_cell_40_90 (.BL(BL90),.BLN(BLN90),.WL(WL40));
sram_cell_6t_5 inst_cell_40_91 (.BL(BL91),.BLN(BLN91),.WL(WL40));
sram_cell_6t_5 inst_cell_40_92 (.BL(BL92),.BLN(BLN92),.WL(WL40));
sram_cell_6t_5 inst_cell_40_93 (.BL(BL93),.BLN(BLN93),.WL(WL40));
sram_cell_6t_5 inst_cell_40_94 (.BL(BL94),.BLN(BLN94),.WL(WL40));
sram_cell_6t_5 inst_cell_40_95 (.BL(BL95),.BLN(BLN95),.WL(WL40));
sram_cell_6t_5 inst_cell_40_96 (.BL(BL96),.BLN(BLN96),.WL(WL40));
sram_cell_6t_5 inst_cell_40_97 (.BL(BL97),.BLN(BLN97),.WL(WL40));
sram_cell_6t_5 inst_cell_40_98 (.BL(BL98),.BLN(BLN98),.WL(WL40));
sram_cell_6t_5 inst_cell_40_99 (.BL(BL99),.BLN(BLN99),.WL(WL40));
sram_cell_6t_5 inst_cell_40_100 (.BL(BL100),.BLN(BLN100),.WL(WL40));
sram_cell_6t_5 inst_cell_40_101 (.BL(BL101),.BLN(BLN101),.WL(WL40));
sram_cell_6t_5 inst_cell_40_102 (.BL(BL102),.BLN(BLN102),.WL(WL40));
sram_cell_6t_5 inst_cell_40_103 (.BL(BL103),.BLN(BLN103),.WL(WL40));
sram_cell_6t_5 inst_cell_40_104 (.BL(BL104),.BLN(BLN104),.WL(WL40));
sram_cell_6t_5 inst_cell_40_105 (.BL(BL105),.BLN(BLN105),.WL(WL40));
sram_cell_6t_5 inst_cell_40_106 (.BL(BL106),.BLN(BLN106),.WL(WL40));
sram_cell_6t_5 inst_cell_40_107 (.BL(BL107),.BLN(BLN107),.WL(WL40));
sram_cell_6t_5 inst_cell_40_108 (.BL(BL108),.BLN(BLN108),.WL(WL40));
sram_cell_6t_5 inst_cell_40_109 (.BL(BL109),.BLN(BLN109),.WL(WL40));
sram_cell_6t_5 inst_cell_40_110 (.BL(BL110),.BLN(BLN110),.WL(WL40));
sram_cell_6t_5 inst_cell_40_111 (.BL(BL111),.BLN(BLN111),.WL(WL40));
sram_cell_6t_5 inst_cell_40_112 (.BL(BL112),.BLN(BLN112),.WL(WL40));
sram_cell_6t_5 inst_cell_40_113 (.BL(BL113),.BLN(BLN113),.WL(WL40));
sram_cell_6t_5 inst_cell_40_114 (.BL(BL114),.BLN(BLN114),.WL(WL40));
sram_cell_6t_5 inst_cell_40_115 (.BL(BL115),.BLN(BLN115),.WL(WL40));
sram_cell_6t_5 inst_cell_40_116 (.BL(BL116),.BLN(BLN116),.WL(WL40));
sram_cell_6t_5 inst_cell_40_117 (.BL(BL117),.BLN(BLN117),.WL(WL40));
sram_cell_6t_5 inst_cell_40_118 (.BL(BL118),.BLN(BLN118),.WL(WL40));
sram_cell_6t_5 inst_cell_40_119 (.BL(BL119),.BLN(BLN119),.WL(WL40));
sram_cell_6t_5 inst_cell_40_120 (.BL(BL120),.BLN(BLN120),.WL(WL40));
sram_cell_6t_5 inst_cell_40_121 (.BL(BL121),.BLN(BLN121),.WL(WL40));
sram_cell_6t_5 inst_cell_40_122 (.BL(BL122),.BLN(BLN122),.WL(WL40));
sram_cell_6t_5 inst_cell_40_123 (.BL(BL123),.BLN(BLN123),.WL(WL40));
sram_cell_6t_5 inst_cell_40_124 (.BL(BL124),.BLN(BLN124),.WL(WL40));
sram_cell_6t_5 inst_cell_40_125 (.BL(BL125),.BLN(BLN125),.WL(WL40));
sram_cell_6t_5 inst_cell_40_126 (.BL(BL126),.BLN(BLN126),.WL(WL40));
sram_cell_6t_5 inst_cell_40_127 (.BL(BL127),.BLN(BLN127),.WL(WL40));
sram_cell_6t_5 inst_cell_41_0 (.BL(BL0),.BLN(BLN0),.WL(WL41));
sram_cell_6t_5 inst_cell_41_1 (.BL(BL1),.BLN(BLN1),.WL(WL41));
sram_cell_6t_5 inst_cell_41_2 (.BL(BL2),.BLN(BLN2),.WL(WL41));
sram_cell_6t_5 inst_cell_41_3 (.BL(BL3),.BLN(BLN3),.WL(WL41));
sram_cell_6t_5 inst_cell_41_4 (.BL(BL4),.BLN(BLN4),.WL(WL41));
sram_cell_6t_5 inst_cell_41_5 (.BL(BL5),.BLN(BLN5),.WL(WL41));
sram_cell_6t_5 inst_cell_41_6 (.BL(BL6),.BLN(BLN6),.WL(WL41));
sram_cell_6t_5 inst_cell_41_7 (.BL(BL7),.BLN(BLN7),.WL(WL41));
sram_cell_6t_5 inst_cell_41_8 (.BL(BL8),.BLN(BLN8),.WL(WL41));
sram_cell_6t_5 inst_cell_41_9 (.BL(BL9),.BLN(BLN9),.WL(WL41));
sram_cell_6t_5 inst_cell_41_10 (.BL(BL10),.BLN(BLN10),.WL(WL41));
sram_cell_6t_5 inst_cell_41_11 (.BL(BL11),.BLN(BLN11),.WL(WL41));
sram_cell_6t_5 inst_cell_41_12 (.BL(BL12),.BLN(BLN12),.WL(WL41));
sram_cell_6t_5 inst_cell_41_13 (.BL(BL13),.BLN(BLN13),.WL(WL41));
sram_cell_6t_5 inst_cell_41_14 (.BL(BL14),.BLN(BLN14),.WL(WL41));
sram_cell_6t_5 inst_cell_41_15 (.BL(BL15),.BLN(BLN15),.WL(WL41));
sram_cell_6t_5 inst_cell_41_16 (.BL(BL16),.BLN(BLN16),.WL(WL41));
sram_cell_6t_5 inst_cell_41_17 (.BL(BL17),.BLN(BLN17),.WL(WL41));
sram_cell_6t_5 inst_cell_41_18 (.BL(BL18),.BLN(BLN18),.WL(WL41));
sram_cell_6t_5 inst_cell_41_19 (.BL(BL19),.BLN(BLN19),.WL(WL41));
sram_cell_6t_5 inst_cell_41_20 (.BL(BL20),.BLN(BLN20),.WL(WL41));
sram_cell_6t_5 inst_cell_41_21 (.BL(BL21),.BLN(BLN21),.WL(WL41));
sram_cell_6t_5 inst_cell_41_22 (.BL(BL22),.BLN(BLN22),.WL(WL41));
sram_cell_6t_5 inst_cell_41_23 (.BL(BL23),.BLN(BLN23),.WL(WL41));
sram_cell_6t_5 inst_cell_41_24 (.BL(BL24),.BLN(BLN24),.WL(WL41));
sram_cell_6t_5 inst_cell_41_25 (.BL(BL25),.BLN(BLN25),.WL(WL41));
sram_cell_6t_5 inst_cell_41_26 (.BL(BL26),.BLN(BLN26),.WL(WL41));
sram_cell_6t_5 inst_cell_41_27 (.BL(BL27),.BLN(BLN27),.WL(WL41));
sram_cell_6t_5 inst_cell_41_28 (.BL(BL28),.BLN(BLN28),.WL(WL41));
sram_cell_6t_5 inst_cell_41_29 (.BL(BL29),.BLN(BLN29),.WL(WL41));
sram_cell_6t_5 inst_cell_41_30 (.BL(BL30),.BLN(BLN30),.WL(WL41));
sram_cell_6t_5 inst_cell_41_31 (.BL(BL31),.BLN(BLN31),.WL(WL41));
sram_cell_6t_5 inst_cell_41_32 (.BL(BL32),.BLN(BLN32),.WL(WL41));
sram_cell_6t_5 inst_cell_41_33 (.BL(BL33),.BLN(BLN33),.WL(WL41));
sram_cell_6t_5 inst_cell_41_34 (.BL(BL34),.BLN(BLN34),.WL(WL41));
sram_cell_6t_5 inst_cell_41_35 (.BL(BL35),.BLN(BLN35),.WL(WL41));
sram_cell_6t_5 inst_cell_41_36 (.BL(BL36),.BLN(BLN36),.WL(WL41));
sram_cell_6t_5 inst_cell_41_37 (.BL(BL37),.BLN(BLN37),.WL(WL41));
sram_cell_6t_5 inst_cell_41_38 (.BL(BL38),.BLN(BLN38),.WL(WL41));
sram_cell_6t_5 inst_cell_41_39 (.BL(BL39),.BLN(BLN39),.WL(WL41));
sram_cell_6t_5 inst_cell_41_40 (.BL(BL40),.BLN(BLN40),.WL(WL41));
sram_cell_6t_5 inst_cell_41_41 (.BL(BL41),.BLN(BLN41),.WL(WL41));
sram_cell_6t_5 inst_cell_41_42 (.BL(BL42),.BLN(BLN42),.WL(WL41));
sram_cell_6t_5 inst_cell_41_43 (.BL(BL43),.BLN(BLN43),.WL(WL41));
sram_cell_6t_5 inst_cell_41_44 (.BL(BL44),.BLN(BLN44),.WL(WL41));
sram_cell_6t_5 inst_cell_41_45 (.BL(BL45),.BLN(BLN45),.WL(WL41));
sram_cell_6t_5 inst_cell_41_46 (.BL(BL46),.BLN(BLN46),.WL(WL41));
sram_cell_6t_5 inst_cell_41_47 (.BL(BL47),.BLN(BLN47),.WL(WL41));
sram_cell_6t_5 inst_cell_41_48 (.BL(BL48),.BLN(BLN48),.WL(WL41));
sram_cell_6t_5 inst_cell_41_49 (.BL(BL49),.BLN(BLN49),.WL(WL41));
sram_cell_6t_5 inst_cell_41_50 (.BL(BL50),.BLN(BLN50),.WL(WL41));
sram_cell_6t_5 inst_cell_41_51 (.BL(BL51),.BLN(BLN51),.WL(WL41));
sram_cell_6t_5 inst_cell_41_52 (.BL(BL52),.BLN(BLN52),.WL(WL41));
sram_cell_6t_5 inst_cell_41_53 (.BL(BL53),.BLN(BLN53),.WL(WL41));
sram_cell_6t_5 inst_cell_41_54 (.BL(BL54),.BLN(BLN54),.WL(WL41));
sram_cell_6t_5 inst_cell_41_55 (.BL(BL55),.BLN(BLN55),.WL(WL41));
sram_cell_6t_5 inst_cell_41_56 (.BL(BL56),.BLN(BLN56),.WL(WL41));
sram_cell_6t_5 inst_cell_41_57 (.BL(BL57),.BLN(BLN57),.WL(WL41));
sram_cell_6t_5 inst_cell_41_58 (.BL(BL58),.BLN(BLN58),.WL(WL41));
sram_cell_6t_5 inst_cell_41_59 (.BL(BL59),.BLN(BLN59),.WL(WL41));
sram_cell_6t_5 inst_cell_41_60 (.BL(BL60),.BLN(BLN60),.WL(WL41));
sram_cell_6t_5 inst_cell_41_61 (.BL(BL61),.BLN(BLN61),.WL(WL41));
sram_cell_6t_5 inst_cell_41_62 (.BL(BL62),.BLN(BLN62),.WL(WL41));
sram_cell_6t_5 inst_cell_41_63 (.BL(BL63),.BLN(BLN63),.WL(WL41));
sram_cell_6t_5 inst_cell_41_64 (.BL(BL64),.BLN(BLN64),.WL(WL41));
sram_cell_6t_5 inst_cell_41_65 (.BL(BL65),.BLN(BLN65),.WL(WL41));
sram_cell_6t_5 inst_cell_41_66 (.BL(BL66),.BLN(BLN66),.WL(WL41));
sram_cell_6t_5 inst_cell_41_67 (.BL(BL67),.BLN(BLN67),.WL(WL41));
sram_cell_6t_5 inst_cell_41_68 (.BL(BL68),.BLN(BLN68),.WL(WL41));
sram_cell_6t_5 inst_cell_41_69 (.BL(BL69),.BLN(BLN69),.WL(WL41));
sram_cell_6t_5 inst_cell_41_70 (.BL(BL70),.BLN(BLN70),.WL(WL41));
sram_cell_6t_5 inst_cell_41_71 (.BL(BL71),.BLN(BLN71),.WL(WL41));
sram_cell_6t_5 inst_cell_41_72 (.BL(BL72),.BLN(BLN72),.WL(WL41));
sram_cell_6t_5 inst_cell_41_73 (.BL(BL73),.BLN(BLN73),.WL(WL41));
sram_cell_6t_5 inst_cell_41_74 (.BL(BL74),.BLN(BLN74),.WL(WL41));
sram_cell_6t_5 inst_cell_41_75 (.BL(BL75),.BLN(BLN75),.WL(WL41));
sram_cell_6t_5 inst_cell_41_76 (.BL(BL76),.BLN(BLN76),.WL(WL41));
sram_cell_6t_5 inst_cell_41_77 (.BL(BL77),.BLN(BLN77),.WL(WL41));
sram_cell_6t_5 inst_cell_41_78 (.BL(BL78),.BLN(BLN78),.WL(WL41));
sram_cell_6t_5 inst_cell_41_79 (.BL(BL79),.BLN(BLN79),.WL(WL41));
sram_cell_6t_5 inst_cell_41_80 (.BL(BL80),.BLN(BLN80),.WL(WL41));
sram_cell_6t_5 inst_cell_41_81 (.BL(BL81),.BLN(BLN81),.WL(WL41));
sram_cell_6t_5 inst_cell_41_82 (.BL(BL82),.BLN(BLN82),.WL(WL41));
sram_cell_6t_5 inst_cell_41_83 (.BL(BL83),.BLN(BLN83),.WL(WL41));
sram_cell_6t_5 inst_cell_41_84 (.BL(BL84),.BLN(BLN84),.WL(WL41));
sram_cell_6t_5 inst_cell_41_85 (.BL(BL85),.BLN(BLN85),.WL(WL41));
sram_cell_6t_5 inst_cell_41_86 (.BL(BL86),.BLN(BLN86),.WL(WL41));
sram_cell_6t_5 inst_cell_41_87 (.BL(BL87),.BLN(BLN87),.WL(WL41));
sram_cell_6t_5 inst_cell_41_88 (.BL(BL88),.BLN(BLN88),.WL(WL41));
sram_cell_6t_5 inst_cell_41_89 (.BL(BL89),.BLN(BLN89),.WL(WL41));
sram_cell_6t_5 inst_cell_41_90 (.BL(BL90),.BLN(BLN90),.WL(WL41));
sram_cell_6t_5 inst_cell_41_91 (.BL(BL91),.BLN(BLN91),.WL(WL41));
sram_cell_6t_5 inst_cell_41_92 (.BL(BL92),.BLN(BLN92),.WL(WL41));
sram_cell_6t_5 inst_cell_41_93 (.BL(BL93),.BLN(BLN93),.WL(WL41));
sram_cell_6t_5 inst_cell_41_94 (.BL(BL94),.BLN(BLN94),.WL(WL41));
sram_cell_6t_5 inst_cell_41_95 (.BL(BL95),.BLN(BLN95),.WL(WL41));
sram_cell_6t_5 inst_cell_41_96 (.BL(BL96),.BLN(BLN96),.WL(WL41));
sram_cell_6t_5 inst_cell_41_97 (.BL(BL97),.BLN(BLN97),.WL(WL41));
sram_cell_6t_5 inst_cell_41_98 (.BL(BL98),.BLN(BLN98),.WL(WL41));
sram_cell_6t_5 inst_cell_41_99 (.BL(BL99),.BLN(BLN99),.WL(WL41));
sram_cell_6t_5 inst_cell_41_100 (.BL(BL100),.BLN(BLN100),.WL(WL41));
sram_cell_6t_5 inst_cell_41_101 (.BL(BL101),.BLN(BLN101),.WL(WL41));
sram_cell_6t_5 inst_cell_41_102 (.BL(BL102),.BLN(BLN102),.WL(WL41));
sram_cell_6t_5 inst_cell_41_103 (.BL(BL103),.BLN(BLN103),.WL(WL41));
sram_cell_6t_5 inst_cell_41_104 (.BL(BL104),.BLN(BLN104),.WL(WL41));
sram_cell_6t_5 inst_cell_41_105 (.BL(BL105),.BLN(BLN105),.WL(WL41));
sram_cell_6t_5 inst_cell_41_106 (.BL(BL106),.BLN(BLN106),.WL(WL41));
sram_cell_6t_5 inst_cell_41_107 (.BL(BL107),.BLN(BLN107),.WL(WL41));
sram_cell_6t_5 inst_cell_41_108 (.BL(BL108),.BLN(BLN108),.WL(WL41));
sram_cell_6t_5 inst_cell_41_109 (.BL(BL109),.BLN(BLN109),.WL(WL41));
sram_cell_6t_5 inst_cell_41_110 (.BL(BL110),.BLN(BLN110),.WL(WL41));
sram_cell_6t_5 inst_cell_41_111 (.BL(BL111),.BLN(BLN111),.WL(WL41));
sram_cell_6t_5 inst_cell_41_112 (.BL(BL112),.BLN(BLN112),.WL(WL41));
sram_cell_6t_5 inst_cell_41_113 (.BL(BL113),.BLN(BLN113),.WL(WL41));
sram_cell_6t_5 inst_cell_41_114 (.BL(BL114),.BLN(BLN114),.WL(WL41));
sram_cell_6t_5 inst_cell_41_115 (.BL(BL115),.BLN(BLN115),.WL(WL41));
sram_cell_6t_5 inst_cell_41_116 (.BL(BL116),.BLN(BLN116),.WL(WL41));
sram_cell_6t_5 inst_cell_41_117 (.BL(BL117),.BLN(BLN117),.WL(WL41));
sram_cell_6t_5 inst_cell_41_118 (.BL(BL118),.BLN(BLN118),.WL(WL41));
sram_cell_6t_5 inst_cell_41_119 (.BL(BL119),.BLN(BLN119),.WL(WL41));
sram_cell_6t_5 inst_cell_41_120 (.BL(BL120),.BLN(BLN120),.WL(WL41));
sram_cell_6t_5 inst_cell_41_121 (.BL(BL121),.BLN(BLN121),.WL(WL41));
sram_cell_6t_5 inst_cell_41_122 (.BL(BL122),.BLN(BLN122),.WL(WL41));
sram_cell_6t_5 inst_cell_41_123 (.BL(BL123),.BLN(BLN123),.WL(WL41));
sram_cell_6t_5 inst_cell_41_124 (.BL(BL124),.BLN(BLN124),.WL(WL41));
sram_cell_6t_5 inst_cell_41_125 (.BL(BL125),.BLN(BLN125),.WL(WL41));
sram_cell_6t_5 inst_cell_41_126 (.BL(BL126),.BLN(BLN126),.WL(WL41));
sram_cell_6t_5 inst_cell_41_127 (.BL(BL127),.BLN(BLN127),.WL(WL41));
sram_cell_6t_5 inst_cell_42_0 (.BL(BL0),.BLN(BLN0),.WL(WL42));
sram_cell_6t_5 inst_cell_42_1 (.BL(BL1),.BLN(BLN1),.WL(WL42));
sram_cell_6t_5 inst_cell_42_2 (.BL(BL2),.BLN(BLN2),.WL(WL42));
sram_cell_6t_5 inst_cell_42_3 (.BL(BL3),.BLN(BLN3),.WL(WL42));
sram_cell_6t_5 inst_cell_42_4 (.BL(BL4),.BLN(BLN4),.WL(WL42));
sram_cell_6t_5 inst_cell_42_5 (.BL(BL5),.BLN(BLN5),.WL(WL42));
sram_cell_6t_5 inst_cell_42_6 (.BL(BL6),.BLN(BLN6),.WL(WL42));
sram_cell_6t_5 inst_cell_42_7 (.BL(BL7),.BLN(BLN7),.WL(WL42));
sram_cell_6t_5 inst_cell_42_8 (.BL(BL8),.BLN(BLN8),.WL(WL42));
sram_cell_6t_5 inst_cell_42_9 (.BL(BL9),.BLN(BLN9),.WL(WL42));
sram_cell_6t_5 inst_cell_42_10 (.BL(BL10),.BLN(BLN10),.WL(WL42));
sram_cell_6t_5 inst_cell_42_11 (.BL(BL11),.BLN(BLN11),.WL(WL42));
sram_cell_6t_5 inst_cell_42_12 (.BL(BL12),.BLN(BLN12),.WL(WL42));
sram_cell_6t_5 inst_cell_42_13 (.BL(BL13),.BLN(BLN13),.WL(WL42));
sram_cell_6t_5 inst_cell_42_14 (.BL(BL14),.BLN(BLN14),.WL(WL42));
sram_cell_6t_5 inst_cell_42_15 (.BL(BL15),.BLN(BLN15),.WL(WL42));
sram_cell_6t_5 inst_cell_42_16 (.BL(BL16),.BLN(BLN16),.WL(WL42));
sram_cell_6t_5 inst_cell_42_17 (.BL(BL17),.BLN(BLN17),.WL(WL42));
sram_cell_6t_5 inst_cell_42_18 (.BL(BL18),.BLN(BLN18),.WL(WL42));
sram_cell_6t_5 inst_cell_42_19 (.BL(BL19),.BLN(BLN19),.WL(WL42));
sram_cell_6t_5 inst_cell_42_20 (.BL(BL20),.BLN(BLN20),.WL(WL42));
sram_cell_6t_5 inst_cell_42_21 (.BL(BL21),.BLN(BLN21),.WL(WL42));
sram_cell_6t_5 inst_cell_42_22 (.BL(BL22),.BLN(BLN22),.WL(WL42));
sram_cell_6t_5 inst_cell_42_23 (.BL(BL23),.BLN(BLN23),.WL(WL42));
sram_cell_6t_5 inst_cell_42_24 (.BL(BL24),.BLN(BLN24),.WL(WL42));
sram_cell_6t_5 inst_cell_42_25 (.BL(BL25),.BLN(BLN25),.WL(WL42));
sram_cell_6t_5 inst_cell_42_26 (.BL(BL26),.BLN(BLN26),.WL(WL42));
sram_cell_6t_5 inst_cell_42_27 (.BL(BL27),.BLN(BLN27),.WL(WL42));
sram_cell_6t_5 inst_cell_42_28 (.BL(BL28),.BLN(BLN28),.WL(WL42));
sram_cell_6t_5 inst_cell_42_29 (.BL(BL29),.BLN(BLN29),.WL(WL42));
sram_cell_6t_5 inst_cell_42_30 (.BL(BL30),.BLN(BLN30),.WL(WL42));
sram_cell_6t_5 inst_cell_42_31 (.BL(BL31),.BLN(BLN31),.WL(WL42));
sram_cell_6t_5 inst_cell_42_32 (.BL(BL32),.BLN(BLN32),.WL(WL42));
sram_cell_6t_5 inst_cell_42_33 (.BL(BL33),.BLN(BLN33),.WL(WL42));
sram_cell_6t_5 inst_cell_42_34 (.BL(BL34),.BLN(BLN34),.WL(WL42));
sram_cell_6t_5 inst_cell_42_35 (.BL(BL35),.BLN(BLN35),.WL(WL42));
sram_cell_6t_5 inst_cell_42_36 (.BL(BL36),.BLN(BLN36),.WL(WL42));
sram_cell_6t_5 inst_cell_42_37 (.BL(BL37),.BLN(BLN37),.WL(WL42));
sram_cell_6t_5 inst_cell_42_38 (.BL(BL38),.BLN(BLN38),.WL(WL42));
sram_cell_6t_5 inst_cell_42_39 (.BL(BL39),.BLN(BLN39),.WL(WL42));
sram_cell_6t_5 inst_cell_42_40 (.BL(BL40),.BLN(BLN40),.WL(WL42));
sram_cell_6t_5 inst_cell_42_41 (.BL(BL41),.BLN(BLN41),.WL(WL42));
sram_cell_6t_5 inst_cell_42_42 (.BL(BL42),.BLN(BLN42),.WL(WL42));
sram_cell_6t_5 inst_cell_42_43 (.BL(BL43),.BLN(BLN43),.WL(WL42));
sram_cell_6t_5 inst_cell_42_44 (.BL(BL44),.BLN(BLN44),.WL(WL42));
sram_cell_6t_5 inst_cell_42_45 (.BL(BL45),.BLN(BLN45),.WL(WL42));
sram_cell_6t_5 inst_cell_42_46 (.BL(BL46),.BLN(BLN46),.WL(WL42));
sram_cell_6t_5 inst_cell_42_47 (.BL(BL47),.BLN(BLN47),.WL(WL42));
sram_cell_6t_5 inst_cell_42_48 (.BL(BL48),.BLN(BLN48),.WL(WL42));
sram_cell_6t_5 inst_cell_42_49 (.BL(BL49),.BLN(BLN49),.WL(WL42));
sram_cell_6t_5 inst_cell_42_50 (.BL(BL50),.BLN(BLN50),.WL(WL42));
sram_cell_6t_5 inst_cell_42_51 (.BL(BL51),.BLN(BLN51),.WL(WL42));
sram_cell_6t_5 inst_cell_42_52 (.BL(BL52),.BLN(BLN52),.WL(WL42));
sram_cell_6t_5 inst_cell_42_53 (.BL(BL53),.BLN(BLN53),.WL(WL42));
sram_cell_6t_5 inst_cell_42_54 (.BL(BL54),.BLN(BLN54),.WL(WL42));
sram_cell_6t_5 inst_cell_42_55 (.BL(BL55),.BLN(BLN55),.WL(WL42));
sram_cell_6t_5 inst_cell_42_56 (.BL(BL56),.BLN(BLN56),.WL(WL42));
sram_cell_6t_5 inst_cell_42_57 (.BL(BL57),.BLN(BLN57),.WL(WL42));
sram_cell_6t_5 inst_cell_42_58 (.BL(BL58),.BLN(BLN58),.WL(WL42));
sram_cell_6t_5 inst_cell_42_59 (.BL(BL59),.BLN(BLN59),.WL(WL42));
sram_cell_6t_5 inst_cell_42_60 (.BL(BL60),.BLN(BLN60),.WL(WL42));
sram_cell_6t_5 inst_cell_42_61 (.BL(BL61),.BLN(BLN61),.WL(WL42));
sram_cell_6t_5 inst_cell_42_62 (.BL(BL62),.BLN(BLN62),.WL(WL42));
sram_cell_6t_5 inst_cell_42_63 (.BL(BL63),.BLN(BLN63),.WL(WL42));
sram_cell_6t_5 inst_cell_42_64 (.BL(BL64),.BLN(BLN64),.WL(WL42));
sram_cell_6t_5 inst_cell_42_65 (.BL(BL65),.BLN(BLN65),.WL(WL42));
sram_cell_6t_5 inst_cell_42_66 (.BL(BL66),.BLN(BLN66),.WL(WL42));
sram_cell_6t_5 inst_cell_42_67 (.BL(BL67),.BLN(BLN67),.WL(WL42));
sram_cell_6t_5 inst_cell_42_68 (.BL(BL68),.BLN(BLN68),.WL(WL42));
sram_cell_6t_5 inst_cell_42_69 (.BL(BL69),.BLN(BLN69),.WL(WL42));
sram_cell_6t_5 inst_cell_42_70 (.BL(BL70),.BLN(BLN70),.WL(WL42));
sram_cell_6t_5 inst_cell_42_71 (.BL(BL71),.BLN(BLN71),.WL(WL42));
sram_cell_6t_5 inst_cell_42_72 (.BL(BL72),.BLN(BLN72),.WL(WL42));
sram_cell_6t_5 inst_cell_42_73 (.BL(BL73),.BLN(BLN73),.WL(WL42));
sram_cell_6t_5 inst_cell_42_74 (.BL(BL74),.BLN(BLN74),.WL(WL42));
sram_cell_6t_5 inst_cell_42_75 (.BL(BL75),.BLN(BLN75),.WL(WL42));
sram_cell_6t_5 inst_cell_42_76 (.BL(BL76),.BLN(BLN76),.WL(WL42));
sram_cell_6t_5 inst_cell_42_77 (.BL(BL77),.BLN(BLN77),.WL(WL42));
sram_cell_6t_5 inst_cell_42_78 (.BL(BL78),.BLN(BLN78),.WL(WL42));
sram_cell_6t_5 inst_cell_42_79 (.BL(BL79),.BLN(BLN79),.WL(WL42));
sram_cell_6t_5 inst_cell_42_80 (.BL(BL80),.BLN(BLN80),.WL(WL42));
sram_cell_6t_5 inst_cell_42_81 (.BL(BL81),.BLN(BLN81),.WL(WL42));
sram_cell_6t_5 inst_cell_42_82 (.BL(BL82),.BLN(BLN82),.WL(WL42));
sram_cell_6t_5 inst_cell_42_83 (.BL(BL83),.BLN(BLN83),.WL(WL42));
sram_cell_6t_5 inst_cell_42_84 (.BL(BL84),.BLN(BLN84),.WL(WL42));
sram_cell_6t_5 inst_cell_42_85 (.BL(BL85),.BLN(BLN85),.WL(WL42));
sram_cell_6t_5 inst_cell_42_86 (.BL(BL86),.BLN(BLN86),.WL(WL42));
sram_cell_6t_5 inst_cell_42_87 (.BL(BL87),.BLN(BLN87),.WL(WL42));
sram_cell_6t_5 inst_cell_42_88 (.BL(BL88),.BLN(BLN88),.WL(WL42));
sram_cell_6t_5 inst_cell_42_89 (.BL(BL89),.BLN(BLN89),.WL(WL42));
sram_cell_6t_5 inst_cell_42_90 (.BL(BL90),.BLN(BLN90),.WL(WL42));
sram_cell_6t_5 inst_cell_42_91 (.BL(BL91),.BLN(BLN91),.WL(WL42));
sram_cell_6t_5 inst_cell_42_92 (.BL(BL92),.BLN(BLN92),.WL(WL42));
sram_cell_6t_5 inst_cell_42_93 (.BL(BL93),.BLN(BLN93),.WL(WL42));
sram_cell_6t_5 inst_cell_42_94 (.BL(BL94),.BLN(BLN94),.WL(WL42));
sram_cell_6t_5 inst_cell_42_95 (.BL(BL95),.BLN(BLN95),.WL(WL42));
sram_cell_6t_5 inst_cell_42_96 (.BL(BL96),.BLN(BLN96),.WL(WL42));
sram_cell_6t_5 inst_cell_42_97 (.BL(BL97),.BLN(BLN97),.WL(WL42));
sram_cell_6t_5 inst_cell_42_98 (.BL(BL98),.BLN(BLN98),.WL(WL42));
sram_cell_6t_5 inst_cell_42_99 (.BL(BL99),.BLN(BLN99),.WL(WL42));
sram_cell_6t_5 inst_cell_42_100 (.BL(BL100),.BLN(BLN100),.WL(WL42));
sram_cell_6t_5 inst_cell_42_101 (.BL(BL101),.BLN(BLN101),.WL(WL42));
sram_cell_6t_5 inst_cell_42_102 (.BL(BL102),.BLN(BLN102),.WL(WL42));
sram_cell_6t_5 inst_cell_42_103 (.BL(BL103),.BLN(BLN103),.WL(WL42));
sram_cell_6t_5 inst_cell_42_104 (.BL(BL104),.BLN(BLN104),.WL(WL42));
sram_cell_6t_5 inst_cell_42_105 (.BL(BL105),.BLN(BLN105),.WL(WL42));
sram_cell_6t_5 inst_cell_42_106 (.BL(BL106),.BLN(BLN106),.WL(WL42));
sram_cell_6t_5 inst_cell_42_107 (.BL(BL107),.BLN(BLN107),.WL(WL42));
sram_cell_6t_5 inst_cell_42_108 (.BL(BL108),.BLN(BLN108),.WL(WL42));
sram_cell_6t_5 inst_cell_42_109 (.BL(BL109),.BLN(BLN109),.WL(WL42));
sram_cell_6t_5 inst_cell_42_110 (.BL(BL110),.BLN(BLN110),.WL(WL42));
sram_cell_6t_5 inst_cell_42_111 (.BL(BL111),.BLN(BLN111),.WL(WL42));
sram_cell_6t_5 inst_cell_42_112 (.BL(BL112),.BLN(BLN112),.WL(WL42));
sram_cell_6t_5 inst_cell_42_113 (.BL(BL113),.BLN(BLN113),.WL(WL42));
sram_cell_6t_5 inst_cell_42_114 (.BL(BL114),.BLN(BLN114),.WL(WL42));
sram_cell_6t_5 inst_cell_42_115 (.BL(BL115),.BLN(BLN115),.WL(WL42));
sram_cell_6t_5 inst_cell_42_116 (.BL(BL116),.BLN(BLN116),.WL(WL42));
sram_cell_6t_5 inst_cell_42_117 (.BL(BL117),.BLN(BLN117),.WL(WL42));
sram_cell_6t_5 inst_cell_42_118 (.BL(BL118),.BLN(BLN118),.WL(WL42));
sram_cell_6t_5 inst_cell_42_119 (.BL(BL119),.BLN(BLN119),.WL(WL42));
sram_cell_6t_5 inst_cell_42_120 (.BL(BL120),.BLN(BLN120),.WL(WL42));
sram_cell_6t_5 inst_cell_42_121 (.BL(BL121),.BLN(BLN121),.WL(WL42));
sram_cell_6t_5 inst_cell_42_122 (.BL(BL122),.BLN(BLN122),.WL(WL42));
sram_cell_6t_5 inst_cell_42_123 (.BL(BL123),.BLN(BLN123),.WL(WL42));
sram_cell_6t_5 inst_cell_42_124 (.BL(BL124),.BLN(BLN124),.WL(WL42));
sram_cell_6t_5 inst_cell_42_125 (.BL(BL125),.BLN(BLN125),.WL(WL42));
sram_cell_6t_5 inst_cell_42_126 (.BL(BL126),.BLN(BLN126),.WL(WL42));
sram_cell_6t_5 inst_cell_42_127 (.BL(BL127),.BLN(BLN127),.WL(WL42));
sram_cell_6t_5 inst_cell_43_0 (.BL(BL0),.BLN(BLN0),.WL(WL43));
sram_cell_6t_5 inst_cell_43_1 (.BL(BL1),.BLN(BLN1),.WL(WL43));
sram_cell_6t_5 inst_cell_43_2 (.BL(BL2),.BLN(BLN2),.WL(WL43));
sram_cell_6t_5 inst_cell_43_3 (.BL(BL3),.BLN(BLN3),.WL(WL43));
sram_cell_6t_5 inst_cell_43_4 (.BL(BL4),.BLN(BLN4),.WL(WL43));
sram_cell_6t_5 inst_cell_43_5 (.BL(BL5),.BLN(BLN5),.WL(WL43));
sram_cell_6t_5 inst_cell_43_6 (.BL(BL6),.BLN(BLN6),.WL(WL43));
sram_cell_6t_5 inst_cell_43_7 (.BL(BL7),.BLN(BLN7),.WL(WL43));
sram_cell_6t_5 inst_cell_43_8 (.BL(BL8),.BLN(BLN8),.WL(WL43));
sram_cell_6t_5 inst_cell_43_9 (.BL(BL9),.BLN(BLN9),.WL(WL43));
sram_cell_6t_5 inst_cell_43_10 (.BL(BL10),.BLN(BLN10),.WL(WL43));
sram_cell_6t_5 inst_cell_43_11 (.BL(BL11),.BLN(BLN11),.WL(WL43));
sram_cell_6t_5 inst_cell_43_12 (.BL(BL12),.BLN(BLN12),.WL(WL43));
sram_cell_6t_5 inst_cell_43_13 (.BL(BL13),.BLN(BLN13),.WL(WL43));
sram_cell_6t_5 inst_cell_43_14 (.BL(BL14),.BLN(BLN14),.WL(WL43));
sram_cell_6t_5 inst_cell_43_15 (.BL(BL15),.BLN(BLN15),.WL(WL43));
sram_cell_6t_5 inst_cell_43_16 (.BL(BL16),.BLN(BLN16),.WL(WL43));
sram_cell_6t_5 inst_cell_43_17 (.BL(BL17),.BLN(BLN17),.WL(WL43));
sram_cell_6t_5 inst_cell_43_18 (.BL(BL18),.BLN(BLN18),.WL(WL43));
sram_cell_6t_5 inst_cell_43_19 (.BL(BL19),.BLN(BLN19),.WL(WL43));
sram_cell_6t_5 inst_cell_43_20 (.BL(BL20),.BLN(BLN20),.WL(WL43));
sram_cell_6t_5 inst_cell_43_21 (.BL(BL21),.BLN(BLN21),.WL(WL43));
sram_cell_6t_5 inst_cell_43_22 (.BL(BL22),.BLN(BLN22),.WL(WL43));
sram_cell_6t_5 inst_cell_43_23 (.BL(BL23),.BLN(BLN23),.WL(WL43));
sram_cell_6t_5 inst_cell_43_24 (.BL(BL24),.BLN(BLN24),.WL(WL43));
sram_cell_6t_5 inst_cell_43_25 (.BL(BL25),.BLN(BLN25),.WL(WL43));
sram_cell_6t_5 inst_cell_43_26 (.BL(BL26),.BLN(BLN26),.WL(WL43));
sram_cell_6t_5 inst_cell_43_27 (.BL(BL27),.BLN(BLN27),.WL(WL43));
sram_cell_6t_5 inst_cell_43_28 (.BL(BL28),.BLN(BLN28),.WL(WL43));
sram_cell_6t_5 inst_cell_43_29 (.BL(BL29),.BLN(BLN29),.WL(WL43));
sram_cell_6t_5 inst_cell_43_30 (.BL(BL30),.BLN(BLN30),.WL(WL43));
sram_cell_6t_5 inst_cell_43_31 (.BL(BL31),.BLN(BLN31),.WL(WL43));
sram_cell_6t_5 inst_cell_43_32 (.BL(BL32),.BLN(BLN32),.WL(WL43));
sram_cell_6t_5 inst_cell_43_33 (.BL(BL33),.BLN(BLN33),.WL(WL43));
sram_cell_6t_5 inst_cell_43_34 (.BL(BL34),.BLN(BLN34),.WL(WL43));
sram_cell_6t_5 inst_cell_43_35 (.BL(BL35),.BLN(BLN35),.WL(WL43));
sram_cell_6t_5 inst_cell_43_36 (.BL(BL36),.BLN(BLN36),.WL(WL43));
sram_cell_6t_5 inst_cell_43_37 (.BL(BL37),.BLN(BLN37),.WL(WL43));
sram_cell_6t_5 inst_cell_43_38 (.BL(BL38),.BLN(BLN38),.WL(WL43));
sram_cell_6t_5 inst_cell_43_39 (.BL(BL39),.BLN(BLN39),.WL(WL43));
sram_cell_6t_5 inst_cell_43_40 (.BL(BL40),.BLN(BLN40),.WL(WL43));
sram_cell_6t_5 inst_cell_43_41 (.BL(BL41),.BLN(BLN41),.WL(WL43));
sram_cell_6t_5 inst_cell_43_42 (.BL(BL42),.BLN(BLN42),.WL(WL43));
sram_cell_6t_5 inst_cell_43_43 (.BL(BL43),.BLN(BLN43),.WL(WL43));
sram_cell_6t_5 inst_cell_43_44 (.BL(BL44),.BLN(BLN44),.WL(WL43));
sram_cell_6t_5 inst_cell_43_45 (.BL(BL45),.BLN(BLN45),.WL(WL43));
sram_cell_6t_5 inst_cell_43_46 (.BL(BL46),.BLN(BLN46),.WL(WL43));
sram_cell_6t_5 inst_cell_43_47 (.BL(BL47),.BLN(BLN47),.WL(WL43));
sram_cell_6t_5 inst_cell_43_48 (.BL(BL48),.BLN(BLN48),.WL(WL43));
sram_cell_6t_5 inst_cell_43_49 (.BL(BL49),.BLN(BLN49),.WL(WL43));
sram_cell_6t_5 inst_cell_43_50 (.BL(BL50),.BLN(BLN50),.WL(WL43));
sram_cell_6t_5 inst_cell_43_51 (.BL(BL51),.BLN(BLN51),.WL(WL43));
sram_cell_6t_5 inst_cell_43_52 (.BL(BL52),.BLN(BLN52),.WL(WL43));
sram_cell_6t_5 inst_cell_43_53 (.BL(BL53),.BLN(BLN53),.WL(WL43));
sram_cell_6t_5 inst_cell_43_54 (.BL(BL54),.BLN(BLN54),.WL(WL43));
sram_cell_6t_5 inst_cell_43_55 (.BL(BL55),.BLN(BLN55),.WL(WL43));
sram_cell_6t_5 inst_cell_43_56 (.BL(BL56),.BLN(BLN56),.WL(WL43));
sram_cell_6t_5 inst_cell_43_57 (.BL(BL57),.BLN(BLN57),.WL(WL43));
sram_cell_6t_5 inst_cell_43_58 (.BL(BL58),.BLN(BLN58),.WL(WL43));
sram_cell_6t_5 inst_cell_43_59 (.BL(BL59),.BLN(BLN59),.WL(WL43));
sram_cell_6t_5 inst_cell_43_60 (.BL(BL60),.BLN(BLN60),.WL(WL43));
sram_cell_6t_5 inst_cell_43_61 (.BL(BL61),.BLN(BLN61),.WL(WL43));
sram_cell_6t_5 inst_cell_43_62 (.BL(BL62),.BLN(BLN62),.WL(WL43));
sram_cell_6t_5 inst_cell_43_63 (.BL(BL63),.BLN(BLN63),.WL(WL43));
sram_cell_6t_5 inst_cell_43_64 (.BL(BL64),.BLN(BLN64),.WL(WL43));
sram_cell_6t_5 inst_cell_43_65 (.BL(BL65),.BLN(BLN65),.WL(WL43));
sram_cell_6t_5 inst_cell_43_66 (.BL(BL66),.BLN(BLN66),.WL(WL43));
sram_cell_6t_5 inst_cell_43_67 (.BL(BL67),.BLN(BLN67),.WL(WL43));
sram_cell_6t_5 inst_cell_43_68 (.BL(BL68),.BLN(BLN68),.WL(WL43));
sram_cell_6t_5 inst_cell_43_69 (.BL(BL69),.BLN(BLN69),.WL(WL43));
sram_cell_6t_5 inst_cell_43_70 (.BL(BL70),.BLN(BLN70),.WL(WL43));
sram_cell_6t_5 inst_cell_43_71 (.BL(BL71),.BLN(BLN71),.WL(WL43));
sram_cell_6t_5 inst_cell_43_72 (.BL(BL72),.BLN(BLN72),.WL(WL43));
sram_cell_6t_5 inst_cell_43_73 (.BL(BL73),.BLN(BLN73),.WL(WL43));
sram_cell_6t_5 inst_cell_43_74 (.BL(BL74),.BLN(BLN74),.WL(WL43));
sram_cell_6t_5 inst_cell_43_75 (.BL(BL75),.BLN(BLN75),.WL(WL43));
sram_cell_6t_5 inst_cell_43_76 (.BL(BL76),.BLN(BLN76),.WL(WL43));
sram_cell_6t_5 inst_cell_43_77 (.BL(BL77),.BLN(BLN77),.WL(WL43));
sram_cell_6t_5 inst_cell_43_78 (.BL(BL78),.BLN(BLN78),.WL(WL43));
sram_cell_6t_5 inst_cell_43_79 (.BL(BL79),.BLN(BLN79),.WL(WL43));
sram_cell_6t_5 inst_cell_43_80 (.BL(BL80),.BLN(BLN80),.WL(WL43));
sram_cell_6t_5 inst_cell_43_81 (.BL(BL81),.BLN(BLN81),.WL(WL43));
sram_cell_6t_5 inst_cell_43_82 (.BL(BL82),.BLN(BLN82),.WL(WL43));
sram_cell_6t_5 inst_cell_43_83 (.BL(BL83),.BLN(BLN83),.WL(WL43));
sram_cell_6t_5 inst_cell_43_84 (.BL(BL84),.BLN(BLN84),.WL(WL43));
sram_cell_6t_5 inst_cell_43_85 (.BL(BL85),.BLN(BLN85),.WL(WL43));
sram_cell_6t_5 inst_cell_43_86 (.BL(BL86),.BLN(BLN86),.WL(WL43));
sram_cell_6t_5 inst_cell_43_87 (.BL(BL87),.BLN(BLN87),.WL(WL43));
sram_cell_6t_5 inst_cell_43_88 (.BL(BL88),.BLN(BLN88),.WL(WL43));
sram_cell_6t_5 inst_cell_43_89 (.BL(BL89),.BLN(BLN89),.WL(WL43));
sram_cell_6t_5 inst_cell_43_90 (.BL(BL90),.BLN(BLN90),.WL(WL43));
sram_cell_6t_5 inst_cell_43_91 (.BL(BL91),.BLN(BLN91),.WL(WL43));
sram_cell_6t_5 inst_cell_43_92 (.BL(BL92),.BLN(BLN92),.WL(WL43));
sram_cell_6t_5 inst_cell_43_93 (.BL(BL93),.BLN(BLN93),.WL(WL43));
sram_cell_6t_5 inst_cell_43_94 (.BL(BL94),.BLN(BLN94),.WL(WL43));
sram_cell_6t_5 inst_cell_43_95 (.BL(BL95),.BLN(BLN95),.WL(WL43));
sram_cell_6t_5 inst_cell_43_96 (.BL(BL96),.BLN(BLN96),.WL(WL43));
sram_cell_6t_5 inst_cell_43_97 (.BL(BL97),.BLN(BLN97),.WL(WL43));
sram_cell_6t_5 inst_cell_43_98 (.BL(BL98),.BLN(BLN98),.WL(WL43));
sram_cell_6t_5 inst_cell_43_99 (.BL(BL99),.BLN(BLN99),.WL(WL43));
sram_cell_6t_5 inst_cell_43_100 (.BL(BL100),.BLN(BLN100),.WL(WL43));
sram_cell_6t_5 inst_cell_43_101 (.BL(BL101),.BLN(BLN101),.WL(WL43));
sram_cell_6t_5 inst_cell_43_102 (.BL(BL102),.BLN(BLN102),.WL(WL43));
sram_cell_6t_5 inst_cell_43_103 (.BL(BL103),.BLN(BLN103),.WL(WL43));
sram_cell_6t_5 inst_cell_43_104 (.BL(BL104),.BLN(BLN104),.WL(WL43));
sram_cell_6t_5 inst_cell_43_105 (.BL(BL105),.BLN(BLN105),.WL(WL43));
sram_cell_6t_5 inst_cell_43_106 (.BL(BL106),.BLN(BLN106),.WL(WL43));
sram_cell_6t_5 inst_cell_43_107 (.BL(BL107),.BLN(BLN107),.WL(WL43));
sram_cell_6t_5 inst_cell_43_108 (.BL(BL108),.BLN(BLN108),.WL(WL43));
sram_cell_6t_5 inst_cell_43_109 (.BL(BL109),.BLN(BLN109),.WL(WL43));
sram_cell_6t_5 inst_cell_43_110 (.BL(BL110),.BLN(BLN110),.WL(WL43));
sram_cell_6t_5 inst_cell_43_111 (.BL(BL111),.BLN(BLN111),.WL(WL43));
sram_cell_6t_5 inst_cell_43_112 (.BL(BL112),.BLN(BLN112),.WL(WL43));
sram_cell_6t_5 inst_cell_43_113 (.BL(BL113),.BLN(BLN113),.WL(WL43));
sram_cell_6t_5 inst_cell_43_114 (.BL(BL114),.BLN(BLN114),.WL(WL43));
sram_cell_6t_5 inst_cell_43_115 (.BL(BL115),.BLN(BLN115),.WL(WL43));
sram_cell_6t_5 inst_cell_43_116 (.BL(BL116),.BLN(BLN116),.WL(WL43));
sram_cell_6t_5 inst_cell_43_117 (.BL(BL117),.BLN(BLN117),.WL(WL43));
sram_cell_6t_5 inst_cell_43_118 (.BL(BL118),.BLN(BLN118),.WL(WL43));
sram_cell_6t_5 inst_cell_43_119 (.BL(BL119),.BLN(BLN119),.WL(WL43));
sram_cell_6t_5 inst_cell_43_120 (.BL(BL120),.BLN(BLN120),.WL(WL43));
sram_cell_6t_5 inst_cell_43_121 (.BL(BL121),.BLN(BLN121),.WL(WL43));
sram_cell_6t_5 inst_cell_43_122 (.BL(BL122),.BLN(BLN122),.WL(WL43));
sram_cell_6t_5 inst_cell_43_123 (.BL(BL123),.BLN(BLN123),.WL(WL43));
sram_cell_6t_5 inst_cell_43_124 (.BL(BL124),.BLN(BLN124),.WL(WL43));
sram_cell_6t_5 inst_cell_43_125 (.BL(BL125),.BLN(BLN125),.WL(WL43));
sram_cell_6t_5 inst_cell_43_126 (.BL(BL126),.BLN(BLN126),.WL(WL43));
sram_cell_6t_5 inst_cell_43_127 (.BL(BL127),.BLN(BLN127),.WL(WL43));
sram_cell_6t_5 inst_cell_44_0 (.BL(BL0),.BLN(BLN0),.WL(WL44));
sram_cell_6t_5 inst_cell_44_1 (.BL(BL1),.BLN(BLN1),.WL(WL44));
sram_cell_6t_5 inst_cell_44_2 (.BL(BL2),.BLN(BLN2),.WL(WL44));
sram_cell_6t_5 inst_cell_44_3 (.BL(BL3),.BLN(BLN3),.WL(WL44));
sram_cell_6t_5 inst_cell_44_4 (.BL(BL4),.BLN(BLN4),.WL(WL44));
sram_cell_6t_5 inst_cell_44_5 (.BL(BL5),.BLN(BLN5),.WL(WL44));
sram_cell_6t_5 inst_cell_44_6 (.BL(BL6),.BLN(BLN6),.WL(WL44));
sram_cell_6t_5 inst_cell_44_7 (.BL(BL7),.BLN(BLN7),.WL(WL44));
sram_cell_6t_5 inst_cell_44_8 (.BL(BL8),.BLN(BLN8),.WL(WL44));
sram_cell_6t_5 inst_cell_44_9 (.BL(BL9),.BLN(BLN9),.WL(WL44));
sram_cell_6t_5 inst_cell_44_10 (.BL(BL10),.BLN(BLN10),.WL(WL44));
sram_cell_6t_5 inst_cell_44_11 (.BL(BL11),.BLN(BLN11),.WL(WL44));
sram_cell_6t_5 inst_cell_44_12 (.BL(BL12),.BLN(BLN12),.WL(WL44));
sram_cell_6t_5 inst_cell_44_13 (.BL(BL13),.BLN(BLN13),.WL(WL44));
sram_cell_6t_5 inst_cell_44_14 (.BL(BL14),.BLN(BLN14),.WL(WL44));
sram_cell_6t_5 inst_cell_44_15 (.BL(BL15),.BLN(BLN15),.WL(WL44));
sram_cell_6t_5 inst_cell_44_16 (.BL(BL16),.BLN(BLN16),.WL(WL44));
sram_cell_6t_5 inst_cell_44_17 (.BL(BL17),.BLN(BLN17),.WL(WL44));
sram_cell_6t_5 inst_cell_44_18 (.BL(BL18),.BLN(BLN18),.WL(WL44));
sram_cell_6t_5 inst_cell_44_19 (.BL(BL19),.BLN(BLN19),.WL(WL44));
sram_cell_6t_5 inst_cell_44_20 (.BL(BL20),.BLN(BLN20),.WL(WL44));
sram_cell_6t_5 inst_cell_44_21 (.BL(BL21),.BLN(BLN21),.WL(WL44));
sram_cell_6t_5 inst_cell_44_22 (.BL(BL22),.BLN(BLN22),.WL(WL44));
sram_cell_6t_5 inst_cell_44_23 (.BL(BL23),.BLN(BLN23),.WL(WL44));
sram_cell_6t_5 inst_cell_44_24 (.BL(BL24),.BLN(BLN24),.WL(WL44));
sram_cell_6t_5 inst_cell_44_25 (.BL(BL25),.BLN(BLN25),.WL(WL44));
sram_cell_6t_5 inst_cell_44_26 (.BL(BL26),.BLN(BLN26),.WL(WL44));
sram_cell_6t_5 inst_cell_44_27 (.BL(BL27),.BLN(BLN27),.WL(WL44));
sram_cell_6t_5 inst_cell_44_28 (.BL(BL28),.BLN(BLN28),.WL(WL44));
sram_cell_6t_5 inst_cell_44_29 (.BL(BL29),.BLN(BLN29),.WL(WL44));
sram_cell_6t_5 inst_cell_44_30 (.BL(BL30),.BLN(BLN30),.WL(WL44));
sram_cell_6t_5 inst_cell_44_31 (.BL(BL31),.BLN(BLN31),.WL(WL44));
sram_cell_6t_5 inst_cell_44_32 (.BL(BL32),.BLN(BLN32),.WL(WL44));
sram_cell_6t_5 inst_cell_44_33 (.BL(BL33),.BLN(BLN33),.WL(WL44));
sram_cell_6t_5 inst_cell_44_34 (.BL(BL34),.BLN(BLN34),.WL(WL44));
sram_cell_6t_5 inst_cell_44_35 (.BL(BL35),.BLN(BLN35),.WL(WL44));
sram_cell_6t_5 inst_cell_44_36 (.BL(BL36),.BLN(BLN36),.WL(WL44));
sram_cell_6t_5 inst_cell_44_37 (.BL(BL37),.BLN(BLN37),.WL(WL44));
sram_cell_6t_5 inst_cell_44_38 (.BL(BL38),.BLN(BLN38),.WL(WL44));
sram_cell_6t_5 inst_cell_44_39 (.BL(BL39),.BLN(BLN39),.WL(WL44));
sram_cell_6t_5 inst_cell_44_40 (.BL(BL40),.BLN(BLN40),.WL(WL44));
sram_cell_6t_5 inst_cell_44_41 (.BL(BL41),.BLN(BLN41),.WL(WL44));
sram_cell_6t_5 inst_cell_44_42 (.BL(BL42),.BLN(BLN42),.WL(WL44));
sram_cell_6t_5 inst_cell_44_43 (.BL(BL43),.BLN(BLN43),.WL(WL44));
sram_cell_6t_5 inst_cell_44_44 (.BL(BL44),.BLN(BLN44),.WL(WL44));
sram_cell_6t_5 inst_cell_44_45 (.BL(BL45),.BLN(BLN45),.WL(WL44));
sram_cell_6t_5 inst_cell_44_46 (.BL(BL46),.BLN(BLN46),.WL(WL44));
sram_cell_6t_5 inst_cell_44_47 (.BL(BL47),.BLN(BLN47),.WL(WL44));
sram_cell_6t_5 inst_cell_44_48 (.BL(BL48),.BLN(BLN48),.WL(WL44));
sram_cell_6t_5 inst_cell_44_49 (.BL(BL49),.BLN(BLN49),.WL(WL44));
sram_cell_6t_5 inst_cell_44_50 (.BL(BL50),.BLN(BLN50),.WL(WL44));
sram_cell_6t_5 inst_cell_44_51 (.BL(BL51),.BLN(BLN51),.WL(WL44));
sram_cell_6t_5 inst_cell_44_52 (.BL(BL52),.BLN(BLN52),.WL(WL44));
sram_cell_6t_5 inst_cell_44_53 (.BL(BL53),.BLN(BLN53),.WL(WL44));
sram_cell_6t_5 inst_cell_44_54 (.BL(BL54),.BLN(BLN54),.WL(WL44));
sram_cell_6t_5 inst_cell_44_55 (.BL(BL55),.BLN(BLN55),.WL(WL44));
sram_cell_6t_5 inst_cell_44_56 (.BL(BL56),.BLN(BLN56),.WL(WL44));
sram_cell_6t_5 inst_cell_44_57 (.BL(BL57),.BLN(BLN57),.WL(WL44));
sram_cell_6t_5 inst_cell_44_58 (.BL(BL58),.BLN(BLN58),.WL(WL44));
sram_cell_6t_5 inst_cell_44_59 (.BL(BL59),.BLN(BLN59),.WL(WL44));
sram_cell_6t_5 inst_cell_44_60 (.BL(BL60),.BLN(BLN60),.WL(WL44));
sram_cell_6t_5 inst_cell_44_61 (.BL(BL61),.BLN(BLN61),.WL(WL44));
sram_cell_6t_5 inst_cell_44_62 (.BL(BL62),.BLN(BLN62),.WL(WL44));
sram_cell_6t_5 inst_cell_44_63 (.BL(BL63),.BLN(BLN63),.WL(WL44));
sram_cell_6t_5 inst_cell_44_64 (.BL(BL64),.BLN(BLN64),.WL(WL44));
sram_cell_6t_5 inst_cell_44_65 (.BL(BL65),.BLN(BLN65),.WL(WL44));
sram_cell_6t_5 inst_cell_44_66 (.BL(BL66),.BLN(BLN66),.WL(WL44));
sram_cell_6t_5 inst_cell_44_67 (.BL(BL67),.BLN(BLN67),.WL(WL44));
sram_cell_6t_5 inst_cell_44_68 (.BL(BL68),.BLN(BLN68),.WL(WL44));
sram_cell_6t_5 inst_cell_44_69 (.BL(BL69),.BLN(BLN69),.WL(WL44));
sram_cell_6t_5 inst_cell_44_70 (.BL(BL70),.BLN(BLN70),.WL(WL44));
sram_cell_6t_5 inst_cell_44_71 (.BL(BL71),.BLN(BLN71),.WL(WL44));
sram_cell_6t_5 inst_cell_44_72 (.BL(BL72),.BLN(BLN72),.WL(WL44));
sram_cell_6t_5 inst_cell_44_73 (.BL(BL73),.BLN(BLN73),.WL(WL44));
sram_cell_6t_5 inst_cell_44_74 (.BL(BL74),.BLN(BLN74),.WL(WL44));
sram_cell_6t_5 inst_cell_44_75 (.BL(BL75),.BLN(BLN75),.WL(WL44));
sram_cell_6t_5 inst_cell_44_76 (.BL(BL76),.BLN(BLN76),.WL(WL44));
sram_cell_6t_5 inst_cell_44_77 (.BL(BL77),.BLN(BLN77),.WL(WL44));
sram_cell_6t_5 inst_cell_44_78 (.BL(BL78),.BLN(BLN78),.WL(WL44));
sram_cell_6t_5 inst_cell_44_79 (.BL(BL79),.BLN(BLN79),.WL(WL44));
sram_cell_6t_5 inst_cell_44_80 (.BL(BL80),.BLN(BLN80),.WL(WL44));
sram_cell_6t_5 inst_cell_44_81 (.BL(BL81),.BLN(BLN81),.WL(WL44));
sram_cell_6t_5 inst_cell_44_82 (.BL(BL82),.BLN(BLN82),.WL(WL44));
sram_cell_6t_5 inst_cell_44_83 (.BL(BL83),.BLN(BLN83),.WL(WL44));
sram_cell_6t_5 inst_cell_44_84 (.BL(BL84),.BLN(BLN84),.WL(WL44));
sram_cell_6t_5 inst_cell_44_85 (.BL(BL85),.BLN(BLN85),.WL(WL44));
sram_cell_6t_5 inst_cell_44_86 (.BL(BL86),.BLN(BLN86),.WL(WL44));
sram_cell_6t_5 inst_cell_44_87 (.BL(BL87),.BLN(BLN87),.WL(WL44));
sram_cell_6t_5 inst_cell_44_88 (.BL(BL88),.BLN(BLN88),.WL(WL44));
sram_cell_6t_5 inst_cell_44_89 (.BL(BL89),.BLN(BLN89),.WL(WL44));
sram_cell_6t_5 inst_cell_44_90 (.BL(BL90),.BLN(BLN90),.WL(WL44));
sram_cell_6t_5 inst_cell_44_91 (.BL(BL91),.BLN(BLN91),.WL(WL44));
sram_cell_6t_5 inst_cell_44_92 (.BL(BL92),.BLN(BLN92),.WL(WL44));
sram_cell_6t_5 inst_cell_44_93 (.BL(BL93),.BLN(BLN93),.WL(WL44));
sram_cell_6t_5 inst_cell_44_94 (.BL(BL94),.BLN(BLN94),.WL(WL44));
sram_cell_6t_5 inst_cell_44_95 (.BL(BL95),.BLN(BLN95),.WL(WL44));
sram_cell_6t_5 inst_cell_44_96 (.BL(BL96),.BLN(BLN96),.WL(WL44));
sram_cell_6t_5 inst_cell_44_97 (.BL(BL97),.BLN(BLN97),.WL(WL44));
sram_cell_6t_5 inst_cell_44_98 (.BL(BL98),.BLN(BLN98),.WL(WL44));
sram_cell_6t_5 inst_cell_44_99 (.BL(BL99),.BLN(BLN99),.WL(WL44));
sram_cell_6t_5 inst_cell_44_100 (.BL(BL100),.BLN(BLN100),.WL(WL44));
sram_cell_6t_5 inst_cell_44_101 (.BL(BL101),.BLN(BLN101),.WL(WL44));
sram_cell_6t_5 inst_cell_44_102 (.BL(BL102),.BLN(BLN102),.WL(WL44));
sram_cell_6t_5 inst_cell_44_103 (.BL(BL103),.BLN(BLN103),.WL(WL44));
sram_cell_6t_5 inst_cell_44_104 (.BL(BL104),.BLN(BLN104),.WL(WL44));
sram_cell_6t_5 inst_cell_44_105 (.BL(BL105),.BLN(BLN105),.WL(WL44));
sram_cell_6t_5 inst_cell_44_106 (.BL(BL106),.BLN(BLN106),.WL(WL44));
sram_cell_6t_5 inst_cell_44_107 (.BL(BL107),.BLN(BLN107),.WL(WL44));
sram_cell_6t_5 inst_cell_44_108 (.BL(BL108),.BLN(BLN108),.WL(WL44));
sram_cell_6t_5 inst_cell_44_109 (.BL(BL109),.BLN(BLN109),.WL(WL44));
sram_cell_6t_5 inst_cell_44_110 (.BL(BL110),.BLN(BLN110),.WL(WL44));
sram_cell_6t_5 inst_cell_44_111 (.BL(BL111),.BLN(BLN111),.WL(WL44));
sram_cell_6t_5 inst_cell_44_112 (.BL(BL112),.BLN(BLN112),.WL(WL44));
sram_cell_6t_5 inst_cell_44_113 (.BL(BL113),.BLN(BLN113),.WL(WL44));
sram_cell_6t_5 inst_cell_44_114 (.BL(BL114),.BLN(BLN114),.WL(WL44));
sram_cell_6t_5 inst_cell_44_115 (.BL(BL115),.BLN(BLN115),.WL(WL44));
sram_cell_6t_5 inst_cell_44_116 (.BL(BL116),.BLN(BLN116),.WL(WL44));
sram_cell_6t_5 inst_cell_44_117 (.BL(BL117),.BLN(BLN117),.WL(WL44));
sram_cell_6t_5 inst_cell_44_118 (.BL(BL118),.BLN(BLN118),.WL(WL44));
sram_cell_6t_5 inst_cell_44_119 (.BL(BL119),.BLN(BLN119),.WL(WL44));
sram_cell_6t_5 inst_cell_44_120 (.BL(BL120),.BLN(BLN120),.WL(WL44));
sram_cell_6t_5 inst_cell_44_121 (.BL(BL121),.BLN(BLN121),.WL(WL44));
sram_cell_6t_5 inst_cell_44_122 (.BL(BL122),.BLN(BLN122),.WL(WL44));
sram_cell_6t_5 inst_cell_44_123 (.BL(BL123),.BLN(BLN123),.WL(WL44));
sram_cell_6t_5 inst_cell_44_124 (.BL(BL124),.BLN(BLN124),.WL(WL44));
sram_cell_6t_5 inst_cell_44_125 (.BL(BL125),.BLN(BLN125),.WL(WL44));
sram_cell_6t_5 inst_cell_44_126 (.BL(BL126),.BLN(BLN126),.WL(WL44));
sram_cell_6t_5 inst_cell_44_127 (.BL(BL127),.BLN(BLN127),.WL(WL44));
sram_cell_6t_5 inst_cell_45_0 (.BL(BL0),.BLN(BLN0),.WL(WL45));
sram_cell_6t_5 inst_cell_45_1 (.BL(BL1),.BLN(BLN1),.WL(WL45));
sram_cell_6t_5 inst_cell_45_2 (.BL(BL2),.BLN(BLN2),.WL(WL45));
sram_cell_6t_5 inst_cell_45_3 (.BL(BL3),.BLN(BLN3),.WL(WL45));
sram_cell_6t_5 inst_cell_45_4 (.BL(BL4),.BLN(BLN4),.WL(WL45));
sram_cell_6t_5 inst_cell_45_5 (.BL(BL5),.BLN(BLN5),.WL(WL45));
sram_cell_6t_5 inst_cell_45_6 (.BL(BL6),.BLN(BLN6),.WL(WL45));
sram_cell_6t_5 inst_cell_45_7 (.BL(BL7),.BLN(BLN7),.WL(WL45));
sram_cell_6t_5 inst_cell_45_8 (.BL(BL8),.BLN(BLN8),.WL(WL45));
sram_cell_6t_5 inst_cell_45_9 (.BL(BL9),.BLN(BLN9),.WL(WL45));
sram_cell_6t_5 inst_cell_45_10 (.BL(BL10),.BLN(BLN10),.WL(WL45));
sram_cell_6t_5 inst_cell_45_11 (.BL(BL11),.BLN(BLN11),.WL(WL45));
sram_cell_6t_5 inst_cell_45_12 (.BL(BL12),.BLN(BLN12),.WL(WL45));
sram_cell_6t_5 inst_cell_45_13 (.BL(BL13),.BLN(BLN13),.WL(WL45));
sram_cell_6t_5 inst_cell_45_14 (.BL(BL14),.BLN(BLN14),.WL(WL45));
sram_cell_6t_5 inst_cell_45_15 (.BL(BL15),.BLN(BLN15),.WL(WL45));
sram_cell_6t_5 inst_cell_45_16 (.BL(BL16),.BLN(BLN16),.WL(WL45));
sram_cell_6t_5 inst_cell_45_17 (.BL(BL17),.BLN(BLN17),.WL(WL45));
sram_cell_6t_5 inst_cell_45_18 (.BL(BL18),.BLN(BLN18),.WL(WL45));
sram_cell_6t_5 inst_cell_45_19 (.BL(BL19),.BLN(BLN19),.WL(WL45));
sram_cell_6t_5 inst_cell_45_20 (.BL(BL20),.BLN(BLN20),.WL(WL45));
sram_cell_6t_5 inst_cell_45_21 (.BL(BL21),.BLN(BLN21),.WL(WL45));
sram_cell_6t_5 inst_cell_45_22 (.BL(BL22),.BLN(BLN22),.WL(WL45));
sram_cell_6t_5 inst_cell_45_23 (.BL(BL23),.BLN(BLN23),.WL(WL45));
sram_cell_6t_5 inst_cell_45_24 (.BL(BL24),.BLN(BLN24),.WL(WL45));
sram_cell_6t_5 inst_cell_45_25 (.BL(BL25),.BLN(BLN25),.WL(WL45));
sram_cell_6t_5 inst_cell_45_26 (.BL(BL26),.BLN(BLN26),.WL(WL45));
sram_cell_6t_5 inst_cell_45_27 (.BL(BL27),.BLN(BLN27),.WL(WL45));
sram_cell_6t_5 inst_cell_45_28 (.BL(BL28),.BLN(BLN28),.WL(WL45));
sram_cell_6t_5 inst_cell_45_29 (.BL(BL29),.BLN(BLN29),.WL(WL45));
sram_cell_6t_5 inst_cell_45_30 (.BL(BL30),.BLN(BLN30),.WL(WL45));
sram_cell_6t_5 inst_cell_45_31 (.BL(BL31),.BLN(BLN31),.WL(WL45));
sram_cell_6t_5 inst_cell_45_32 (.BL(BL32),.BLN(BLN32),.WL(WL45));
sram_cell_6t_5 inst_cell_45_33 (.BL(BL33),.BLN(BLN33),.WL(WL45));
sram_cell_6t_5 inst_cell_45_34 (.BL(BL34),.BLN(BLN34),.WL(WL45));
sram_cell_6t_5 inst_cell_45_35 (.BL(BL35),.BLN(BLN35),.WL(WL45));
sram_cell_6t_5 inst_cell_45_36 (.BL(BL36),.BLN(BLN36),.WL(WL45));
sram_cell_6t_5 inst_cell_45_37 (.BL(BL37),.BLN(BLN37),.WL(WL45));
sram_cell_6t_5 inst_cell_45_38 (.BL(BL38),.BLN(BLN38),.WL(WL45));
sram_cell_6t_5 inst_cell_45_39 (.BL(BL39),.BLN(BLN39),.WL(WL45));
sram_cell_6t_5 inst_cell_45_40 (.BL(BL40),.BLN(BLN40),.WL(WL45));
sram_cell_6t_5 inst_cell_45_41 (.BL(BL41),.BLN(BLN41),.WL(WL45));
sram_cell_6t_5 inst_cell_45_42 (.BL(BL42),.BLN(BLN42),.WL(WL45));
sram_cell_6t_5 inst_cell_45_43 (.BL(BL43),.BLN(BLN43),.WL(WL45));
sram_cell_6t_5 inst_cell_45_44 (.BL(BL44),.BLN(BLN44),.WL(WL45));
sram_cell_6t_5 inst_cell_45_45 (.BL(BL45),.BLN(BLN45),.WL(WL45));
sram_cell_6t_5 inst_cell_45_46 (.BL(BL46),.BLN(BLN46),.WL(WL45));
sram_cell_6t_5 inst_cell_45_47 (.BL(BL47),.BLN(BLN47),.WL(WL45));
sram_cell_6t_5 inst_cell_45_48 (.BL(BL48),.BLN(BLN48),.WL(WL45));
sram_cell_6t_5 inst_cell_45_49 (.BL(BL49),.BLN(BLN49),.WL(WL45));
sram_cell_6t_5 inst_cell_45_50 (.BL(BL50),.BLN(BLN50),.WL(WL45));
sram_cell_6t_5 inst_cell_45_51 (.BL(BL51),.BLN(BLN51),.WL(WL45));
sram_cell_6t_5 inst_cell_45_52 (.BL(BL52),.BLN(BLN52),.WL(WL45));
sram_cell_6t_5 inst_cell_45_53 (.BL(BL53),.BLN(BLN53),.WL(WL45));
sram_cell_6t_5 inst_cell_45_54 (.BL(BL54),.BLN(BLN54),.WL(WL45));
sram_cell_6t_5 inst_cell_45_55 (.BL(BL55),.BLN(BLN55),.WL(WL45));
sram_cell_6t_5 inst_cell_45_56 (.BL(BL56),.BLN(BLN56),.WL(WL45));
sram_cell_6t_5 inst_cell_45_57 (.BL(BL57),.BLN(BLN57),.WL(WL45));
sram_cell_6t_5 inst_cell_45_58 (.BL(BL58),.BLN(BLN58),.WL(WL45));
sram_cell_6t_5 inst_cell_45_59 (.BL(BL59),.BLN(BLN59),.WL(WL45));
sram_cell_6t_5 inst_cell_45_60 (.BL(BL60),.BLN(BLN60),.WL(WL45));
sram_cell_6t_5 inst_cell_45_61 (.BL(BL61),.BLN(BLN61),.WL(WL45));
sram_cell_6t_5 inst_cell_45_62 (.BL(BL62),.BLN(BLN62),.WL(WL45));
sram_cell_6t_5 inst_cell_45_63 (.BL(BL63),.BLN(BLN63),.WL(WL45));
sram_cell_6t_5 inst_cell_45_64 (.BL(BL64),.BLN(BLN64),.WL(WL45));
sram_cell_6t_5 inst_cell_45_65 (.BL(BL65),.BLN(BLN65),.WL(WL45));
sram_cell_6t_5 inst_cell_45_66 (.BL(BL66),.BLN(BLN66),.WL(WL45));
sram_cell_6t_5 inst_cell_45_67 (.BL(BL67),.BLN(BLN67),.WL(WL45));
sram_cell_6t_5 inst_cell_45_68 (.BL(BL68),.BLN(BLN68),.WL(WL45));
sram_cell_6t_5 inst_cell_45_69 (.BL(BL69),.BLN(BLN69),.WL(WL45));
sram_cell_6t_5 inst_cell_45_70 (.BL(BL70),.BLN(BLN70),.WL(WL45));
sram_cell_6t_5 inst_cell_45_71 (.BL(BL71),.BLN(BLN71),.WL(WL45));
sram_cell_6t_5 inst_cell_45_72 (.BL(BL72),.BLN(BLN72),.WL(WL45));
sram_cell_6t_5 inst_cell_45_73 (.BL(BL73),.BLN(BLN73),.WL(WL45));
sram_cell_6t_5 inst_cell_45_74 (.BL(BL74),.BLN(BLN74),.WL(WL45));
sram_cell_6t_5 inst_cell_45_75 (.BL(BL75),.BLN(BLN75),.WL(WL45));
sram_cell_6t_5 inst_cell_45_76 (.BL(BL76),.BLN(BLN76),.WL(WL45));
sram_cell_6t_5 inst_cell_45_77 (.BL(BL77),.BLN(BLN77),.WL(WL45));
sram_cell_6t_5 inst_cell_45_78 (.BL(BL78),.BLN(BLN78),.WL(WL45));
sram_cell_6t_5 inst_cell_45_79 (.BL(BL79),.BLN(BLN79),.WL(WL45));
sram_cell_6t_5 inst_cell_45_80 (.BL(BL80),.BLN(BLN80),.WL(WL45));
sram_cell_6t_5 inst_cell_45_81 (.BL(BL81),.BLN(BLN81),.WL(WL45));
sram_cell_6t_5 inst_cell_45_82 (.BL(BL82),.BLN(BLN82),.WL(WL45));
sram_cell_6t_5 inst_cell_45_83 (.BL(BL83),.BLN(BLN83),.WL(WL45));
sram_cell_6t_5 inst_cell_45_84 (.BL(BL84),.BLN(BLN84),.WL(WL45));
sram_cell_6t_5 inst_cell_45_85 (.BL(BL85),.BLN(BLN85),.WL(WL45));
sram_cell_6t_5 inst_cell_45_86 (.BL(BL86),.BLN(BLN86),.WL(WL45));
sram_cell_6t_5 inst_cell_45_87 (.BL(BL87),.BLN(BLN87),.WL(WL45));
sram_cell_6t_5 inst_cell_45_88 (.BL(BL88),.BLN(BLN88),.WL(WL45));
sram_cell_6t_5 inst_cell_45_89 (.BL(BL89),.BLN(BLN89),.WL(WL45));
sram_cell_6t_5 inst_cell_45_90 (.BL(BL90),.BLN(BLN90),.WL(WL45));
sram_cell_6t_5 inst_cell_45_91 (.BL(BL91),.BLN(BLN91),.WL(WL45));
sram_cell_6t_5 inst_cell_45_92 (.BL(BL92),.BLN(BLN92),.WL(WL45));
sram_cell_6t_5 inst_cell_45_93 (.BL(BL93),.BLN(BLN93),.WL(WL45));
sram_cell_6t_5 inst_cell_45_94 (.BL(BL94),.BLN(BLN94),.WL(WL45));
sram_cell_6t_5 inst_cell_45_95 (.BL(BL95),.BLN(BLN95),.WL(WL45));
sram_cell_6t_5 inst_cell_45_96 (.BL(BL96),.BLN(BLN96),.WL(WL45));
sram_cell_6t_5 inst_cell_45_97 (.BL(BL97),.BLN(BLN97),.WL(WL45));
sram_cell_6t_5 inst_cell_45_98 (.BL(BL98),.BLN(BLN98),.WL(WL45));
sram_cell_6t_5 inst_cell_45_99 (.BL(BL99),.BLN(BLN99),.WL(WL45));
sram_cell_6t_5 inst_cell_45_100 (.BL(BL100),.BLN(BLN100),.WL(WL45));
sram_cell_6t_5 inst_cell_45_101 (.BL(BL101),.BLN(BLN101),.WL(WL45));
sram_cell_6t_5 inst_cell_45_102 (.BL(BL102),.BLN(BLN102),.WL(WL45));
sram_cell_6t_5 inst_cell_45_103 (.BL(BL103),.BLN(BLN103),.WL(WL45));
sram_cell_6t_5 inst_cell_45_104 (.BL(BL104),.BLN(BLN104),.WL(WL45));
sram_cell_6t_5 inst_cell_45_105 (.BL(BL105),.BLN(BLN105),.WL(WL45));
sram_cell_6t_5 inst_cell_45_106 (.BL(BL106),.BLN(BLN106),.WL(WL45));
sram_cell_6t_5 inst_cell_45_107 (.BL(BL107),.BLN(BLN107),.WL(WL45));
sram_cell_6t_5 inst_cell_45_108 (.BL(BL108),.BLN(BLN108),.WL(WL45));
sram_cell_6t_5 inst_cell_45_109 (.BL(BL109),.BLN(BLN109),.WL(WL45));
sram_cell_6t_5 inst_cell_45_110 (.BL(BL110),.BLN(BLN110),.WL(WL45));
sram_cell_6t_5 inst_cell_45_111 (.BL(BL111),.BLN(BLN111),.WL(WL45));
sram_cell_6t_5 inst_cell_45_112 (.BL(BL112),.BLN(BLN112),.WL(WL45));
sram_cell_6t_5 inst_cell_45_113 (.BL(BL113),.BLN(BLN113),.WL(WL45));
sram_cell_6t_5 inst_cell_45_114 (.BL(BL114),.BLN(BLN114),.WL(WL45));
sram_cell_6t_5 inst_cell_45_115 (.BL(BL115),.BLN(BLN115),.WL(WL45));
sram_cell_6t_5 inst_cell_45_116 (.BL(BL116),.BLN(BLN116),.WL(WL45));
sram_cell_6t_5 inst_cell_45_117 (.BL(BL117),.BLN(BLN117),.WL(WL45));
sram_cell_6t_5 inst_cell_45_118 (.BL(BL118),.BLN(BLN118),.WL(WL45));
sram_cell_6t_5 inst_cell_45_119 (.BL(BL119),.BLN(BLN119),.WL(WL45));
sram_cell_6t_5 inst_cell_45_120 (.BL(BL120),.BLN(BLN120),.WL(WL45));
sram_cell_6t_5 inst_cell_45_121 (.BL(BL121),.BLN(BLN121),.WL(WL45));
sram_cell_6t_5 inst_cell_45_122 (.BL(BL122),.BLN(BLN122),.WL(WL45));
sram_cell_6t_5 inst_cell_45_123 (.BL(BL123),.BLN(BLN123),.WL(WL45));
sram_cell_6t_5 inst_cell_45_124 (.BL(BL124),.BLN(BLN124),.WL(WL45));
sram_cell_6t_5 inst_cell_45_125 (.BL(BL125),.BLN(BLN125),.WL(WL45));
sram_cell_6t_5 inst_cell_45_126 (.BL(BL126),.BLN(BLN126),.WL(WL45));
sram_cell_6t_5 inst_cell_45_127 (.BL(BL127),.BLN(BLN127),.WL(WL45));
sram_cell_6t_5 inst_cell_46_0 (.BL(BL0),.BLN(BLN0),.WL(WL46));
sram_cell_6t_5 inst_cell_46_1 (.BL(BL1),.BLN(BLN1),.WL(WL46));
sram_cell_6t_5 inst_cell_46_2 (.BL(BL2),.BLN(BLN2),.WL(WL46));
sram_cell_6t_5 inst_cell_46_3 (.BL(BL3),.BLN(BLN3),.WL(WL46));
sram_cell_6t_5 inst_cell_46_4 (.BL(BL4),.BLN(BLN4),.WL(WL46));
sram_cell_6t_5 inst_cell_46_5 (.BL(BL5),.BLN(BLN5),.WL(WL46));
sram_cell_6t_5 inst_cell_46_6 (.BL(BL6),.BLN(BLN6),.WL(WL46));
sram_cell_6t_5 inst_cell_46_7 (.BL(BL7),.BLN(BLN7),.WL(WL46));
sram_cell_6t_5 inst_cell_46_8 (.BL(BL8),.BLN(BLN8),.WL(WL46));
sram_cell_6t_5 inst_cell_46_9 (.BL(BL9),.BLN(BLN9),.WL(WL46));
sram_cell_6t_5 inst_cell_46_10 (.BL(BL10),.BLN(BLN10),.WL(WL46));
sram_cell_6t_5 inst_cell_46_11 (.BL(BL11),.BLN(BLN11),.WL(WL46));
sram_cell_6t_5 inst_cell_46_12 (.BL(BL12),.BLN(BLN12),.WL(WL46));
sram_cell_6t_5 inst_cell_46_13 (.BL(BL13),.BLN(BLN13),.WL(WL46));
sram_cell_6t_5 inst_cell_46_14 (.BL(BL14),.BLN(BLN14),.WL(WL46));
sram_cell_6t_5 inst_cell_46_15 (.BL(BL15),.BLN(BLN15),.WL(WL46));
sram_cell_6t_5 inst_cell_46_16 (.BL(BL16),.BLN(BLN16),.WL(WL46));
sram_cell_6t_5 inst_cell_46_17 (.BL(BL17),.BLN(BLN17),.WL(WL46));
sram_cell_6t_5 inst_cell_46_18 (.BL(BL18),.BLN(BLN18),.WL(WL46));
sram_cell_6t_5 inst_cell_46_19 (.BL(BL19),.BLN(BLN19),.WL(WL46));
sram_cell_6t_5 inst_cell_46_20 (.BL(BL20),.BLN(BLN20),.WL(WL46));
sram_cell_6t_5 inst_cell_46_21 (.BL(BL21),.BLN(BLN21),.WL(WL46));
sram_cell_6t_5 inst_cell_46_22 (.BL(BL22),.BLN(BLN22),.WL(WL46));
sram_cell_6t_5 inst_cell_46_23 (.BL(BL23),.BLN(BLN23),.WL(WL46));
sram_cell_6t_5 inst_cell_46_24 (.BL(BL24),.BLN(BLN24),.WL(WL46));
sram_cell_6t_5 inst_cell_46_25 (.BL(BL25),.BLN(BLN25),.WL(WL46));
sram_cell_6t_5 inst_cell_46_26 (.BL(BL26),.BLN(BLN26),.WL(WL46));
sram_cell_6t_5 inst_cell_46_27 (.BL(BL27),.BLN(BLN27),.WL(WL46));
sram_cell_6t_5 inst_cell_46_28 (.BL(BL28),.BLN(BLN28),.WL(WL46));
sram_cell_6t_5 inst_cell_46_29 (.BL(BL29),.BLN(BLN29),.WL(WL46));
sram_cell_6t_5 inst_cell_46_30 (.BL(BL30),.BLN(BLN30),.WL(WL46));
sram_cell_6t_5 inst_cell_46_31 (.BL(BL31),.BLN(BLN31),.WL(WL46));
sram_cell_6t_5 inst_cell_46_32 (.BL(BL32),.BLN(BLN32),.WL(WL46));
sram_cell_6t_5 inst_cell_46_33 (.BL(BL33),.BLN(BLN33),.WL(WL46));
sram_cell_6t_5 inst_cell_46_34 (.BL(BL34),.BLN(BLN34),.WL(WL46));
sram_cell_6t_5 inst_cell_46_35 (.BL(BL35),.BLN(BLN35),.WL(WL46));
sram_cell_6t_5 inst_cell_46_36 (.BL(BL36),.BLN(BLN36),.WL(WL46));
sram_cell_6t_5 inst_cell_46_37 (.BL(BL37),.BLN(BLN37),.WL(WL46));
sram_cell_6t_5 inst_cell_46_38 (.BL(BL38),.BLN(BLN38),.WL(WL46));
sram_cell_6t_5 inst_cell_46_39 (.BL(BL39),.BLN(BLN39),.WL(WL46));
sram_cell_6t_5 inst_cell_46_40 (.BL(BL40),.BLN(BLN40),.WL(WL46));
sram_cell_6t_5 inst_cell_46_41 (.BL(BL41),.BLN(BLN41),.WL(WL46));
sram_cell_6t_5 inst_cell_46_42 (.BL(BL42),.BLN(BLN42),.WL(WL46));
sram_cell_6t_5 inst_cell_46_43 (.BL(BL43),.BLN(BLN43),.WL(WL46));
sram_cell_6t_5 inst_cell_46_44 (.BL(BL44),.BLN(BLN44),.WL(WL46));
sram_cell_6t_5 inst_cell_46_45 (.BL(BL45),.BLN(BLN45),.WL(WL46));
sram_cell_6t_5 inst_cell_46_46 (.BL(BL46),.BLN(BLN46),.WL(WL46));
sram_cell_6t_5 inst_cell_46_47 (.BL(BL47),.BLN(BLN47),.WL(WL46));
sram_cell_6t_5 inst_cell_46_48 (.BL(BL48),.BLN(BLN48),.WL(WL46));
sram_cell_6t_5 inst_cell_46_49 (.BL(BL49),.BLN(BLN49),.WL(WL46));
sram_cell_6t_5 inst_cell_46_50 (.BL(BL50),.BLN(BLN50),.WL(WL46));
sram_cell_6t_5 inst_cell_46_51 (.BL(BL51),.BLN(BLN51),.WL(WL46));
sram_cell_6t_5 inst_cell_46_52 (.BL(BL52),.BLN(BLN52),.WL(WL46));
sram_cell_6t_5 inst_cell_46_53 (.BL(BL53),.BLN(BLN53),.WL(WL46));
sram_cell_6t_5 inst_cell_46_54 (.BL(BL54),.BLN(BLN54),.WL(WL46));
sram_cell_6t_5 inst_cell_46_55 (.BL(BL55),.BLN(BLN55),.WL(WL46));
sram_cell_6t_5 inst_cell_46_56 (.BL(BL56),.BLN(BLN56),.WL(WL46));
sram_cell_6t_5 inst_cell_46_57 (.BL(BL57),.BLN(BLN57),.WL(WL46));
sram_cell_6t_5 inst_cell_46_58 (.BL(BL58),.BLN(BLN58),.WL(WL46));
sram_cell_6t_5 inst_cell_46_59 (.BL(BL59),.BLN(BLN59),.WL(WL46));
sram_cell_6t_5 inst_cell_46_60 (.BL(BL60),.BLN(BLN60),.WL(WL46));
sram_cell_6t_5 inst_cell_46_61 (.BL(BL61),.BLN(BLN61),.WL(WL46));
sram_cell_6t_5 inst_cell_46_62 (.BL(BL62),.BLN(BLN62),.WL(WL46));
sram_cell_6t_5 inst_cell_46_63 (.BL(BL63),.BLN(BLN63),.WL(WL46));
sram_cell_6t_5 inst_cell_46_64 (.BL(BL64),.BLN(BLN64),.WL(WL46));
sram_cell_6t_5 inst_cell_46_65 (.BL(BL65),.BLN(BLN65),.WL(WL46));
sram_cell_6t_5 inst_cell_46_66 (.BL(BL66),.BLN(BLN66),.WL(WL46));
sram_cell_6t_5 inst_cell_46_67 (.BL(BL67),.BLN(BLN67),.WL(WL46));
sram_cell_6t_5 inst_cell_46_68 (.BL(BL68),.BLN(BLN68),.WL(WL46));
sram_cell_6t_5 inst_cell_46_69 (.BL(BL69),.BLN(BLN69),.WL(WL46));
sram_cell_6t_5 inst_cell_46_70 (.BL(BL70),.BLN(BLN70),.WL(WL46));
sram_cell_6t_5 inst_cell_46_71 (.BL(BL71),.BLN(BLN71),.WL(WL46));
sram_cell_6t_5 inst_cell_46_72 (.BL(BL72),.BLN(BLN72),.WL(WL46));
sram_cell_6t_5 inst_cell_46_73 (.BL(BL73),.BLN(BLN73),.WL(WL46));
sram_cell_6t_5 inst_cell_46_74 (.BL(BL74),.BLN(BLN74),.WL(WL46));
sram_cell_6t_5 inst_cell_46_75 (.BL(BL75),.BLN(BLN75),.WL(WL46));
sram_cell_6t_5 inst_cell_46_76 (.BL(BL76),.BLN(BLN76),.WL(WL46));
sram_cell_6t_5 inst_cell_46_77 (.BL(BL77),.BLN(BLN77),.WL(WL46));
sram_cell_6t_5 inst_cell_46_78 (.BL(BL78),.BLN(BLN78),.WL(WL46));
sram_cell_6t_5 inst_cell_46_79 (.BL(BL79),.BLN(BLN79),.WL(WL46));
sram_cell_6t_5 inst_cell_46_80 (.BL(BL80),.BLN(BLN80),.WL(WL46));
sram_cell_6t_5 inst_cell_46_81 (.BL(BL81),.BLN(BLN81),.WL(WL46));
sram_cell_6t_5 inst_cell_46_82 (.BL(BL82),.BLN(BLN82),.WL(WL46));
sram_cell_6t_5 inst_cell_46_83 (.BL(BL83),.BLN(BLN83),.WL(WL46));
sram_cell_6t_5 inst_cell_46_84 (.BL(BL84),.BLN(BLN84),.WL(WL46));
sram_cell_6t_5 inst_cell_46_85 (.BL(BL85),.BLN(BLN85),.WL(WL46));
sram_cell_6t_5 inst_cell_46_86 (.BL(BL86),.BLN(BLN86),.WL(WL46));
sram_cell_6t_5 inst_cell_46_87 (.BL(BL87),.BLN(BLN87),.WL(WL46));
sram_cell_6t_5 inst_cell_46_88 (.BL(BL88),.BLN(BLN88),.WL(WL46));
sram_cell_6t_5 inst_cell_46_89 (.BL(BL89),.BLN(BLN89),.WL(WL46));
sram_cell_6t_5 inst_cell_46_90 (.BL(BL90),.BLN(BLN90),.WL(WL46));
sram_cell_6t_5 inst_cell_46_91 (.BL(BL91),.BLN(BLN91),.WL(WL46));
sram_cell_6t_5 inst_cell_46_92 (.BL(BL92),.BLN(BLN92),.WL(WL46));
sram_cell_6t_5 inst_cell_46_93 (.BL(BL93),.BLN(BLN93),.WL(WL46));
sram_cell_6t_5 inst_cell_46_94 (.BL(BL94),.BLN(BLN94),.WL(WL46));
sram_cell_6t_5 inst_cell_46_95 (.BL(BL95),.BLN(BLN95),.WL(WL46));
sram_cell_6t_5 inst_cell_46_96 (.BL(BL96),.BLN(BLN96),.WL(WL46));
sram_cell_6t_5 inst_cell_46_97 (.BL(BL97),.BLN(BLN97),.WL(WL46));
sram_cell_6t_5 inst_cell_46_98 (.BL(BL98),.BLN(BLN98),.WL(WL46));
sram_cell_6t_5 inst_cell_46_99 (.BL(BL99),.BLN(BLN99),.WL(WL46));
sram_cell_6t_5 inst_cell_46_100 (.BL(BL100),.BLN(BLN100),.WL(WL46));
sram_cell_6t_5 inst_cell_46_101 (.BL(BL101),.BLN(BLN101),.WL(WL46));
sram_cell_6t_5 inst_cell_46_102 (.BL(BL102),.BLN(BLN102),.WL(WL46));
sram_cell_6t_5 inst_cell_46_103 (.BL(BL103),.BLN(BLN103),.WL(WL46));
sram_cell_6t_5 inst_cell_46_104 (.BL(BL104),.BLN(BLN104),.WL(WL46));
sram_cell_6t_5 inst_cell_46_105 (.BL(BL105),.BLN(BLN105),.WL(WL46));
sram_cell_6t_5 inst_cell_46_106 (.BL(BL106),.BLN(BLN106),.WL(WL46));
sram_cell_6t_5 inst_cell_46_107 (.BL(BL107),.BLN(BLN107),.WL(WL46));
sram_cell_6t_5 inst_cell_46_108 (.BL(BL108),.BLN(BLN108),.WL(WL46));
sram_cell_6t_5 inst_cell_46_109 (.BL(BL109),.BLN(BLN109),.WL(WL46));
sram_cell_6t_5 inst_cell_46_110 (.BL(BL110),.BLN(BLN110),.WL(WL46));
sram_cell_6t_5 inst_cell_46_111 (.BL(BL111),.BLN(BLN111),.WL(WL46));
sram_cell_6t_5 inst_cell_46_112 (.BL(BL112),.BLN(BLN112),.WL(WL46));
sram_cell_6t_5 inst_cell_46_113 (.BL(BL113),.BLN(BLN113),.WL(WL46));
sram_cell_6t_5 inst_cell_46_114 (.BL(BL114),.BLN(BLN114),.WL(WL46));
sram_cell_6t_5 inst_cell_46_115 (.BL(BL115),.BLN(BLN115),.WL(WL46));
sram_cell_6t_5 inst_cell_46_116 (.BL(BL116),.BLN(BLN116),.WL(WL46));
sram_cell_6t_5 inst_cell_46_117 (.BL(BL117),.BLN(BLN117),.WL(WL46));
sram_cell_6t_5 inst_cell_46_118 (.BL(BL118),.BLN(BLN118),.WL(WL46));
sram_cell_6t_5 inst_cell_46_119 (.BL(BL119),.BLN(BLN119),.WL(WL46));
sram_cell_6t_5 inst_cell_46_120 (.BL(BL120),.BLN(BLN120),.WL(WL46));
sram_cell_6t_5 inst_cell_46_121 (.BL(BL121),.BLN(BLN121),.WL(WL46));
sram_cell_6t_5 inst_cell_46_122 (.BL(BL122),.BLN(BLN122),.WL(WL46));
sram_cell_6t_5 inst_cell_46_123 (.BL(BL123),.BLN(BLN123),.WL(WL46));
sram_cell_6t_5 inst_cell_46_124 (.BL(BL124),.BLN(BLN124),.WL(WL46));
sram_cell_6t_5 inst_cell_46_125 (.BL(BL125),.BLN(BLN125),.WL(WL46));
sram_cell_6t_5 inst_cell_46_126 (.BL(BL126),.BLN(BLN126),.WL(WL46));
sram_cell_6t_5 inst_cell_46_127 (.BL(BL127),.BLN(BLN127),.WL(WL46));
sram_cell_6t_5 inst_cell_47_0 (.BL(BL0),.BLN(BLN0),.WL(WL47));
sram_cell_6t_5 inst_cell_47_1 (.BL(BL1),.BLN(BLN1),.WL(WL47));
sram_cell_6t_5 inst_cell_47_2 (.BL(BL2),.BLN(BLN2),.WL(WL47));
sram_cell_6t_5 inst_cell_47_3 (.BL(BL3),.BLN(BLN3),.WL(WL47));
sram_cell_6t_5 inst_cell_47_4 (.BL(BL4),.BLN(BLN4),.WL(WL47));
sram_cell_6t_5 inst_cell_47_5 (.BL(BL5),.BLN(BLN5),.WL(WL47));
sram_cell_6t_5 inst_cell_47_6 (.BL(BL6),.BLN(BLN6),.WL(WL47));
sram_cell_6t_5 inst_cell_47_7 (.BL(BL7),.BLN(BLN7),.WL(WL47));
sram_cell_6t_5 inst_cell_47_8 (.BL(BL8),.BLN(BLN8),.WL(WL47));
sram_cell_6t_5 inst_cell_47_9 (.BL(BL9),.BLN(BLN9),.WL(WL47));
sram_cell_6t_5 inst_cell_47_10 (.BL(BL10),.BLN(BLN10),.WL(WL47));
sram_cell_6t_5 inst_cell_47_11 (.BL(BL11),.BLN(BLN11),.WL(WL47));
sram_cell_6t_5 inst_cell_47_12 (.BL(BL12),.BLN(BLN12),.WL(WL47));
sram_cell_6t_5 inst_cell_47_13 (.BL(BL13),.BLN(BLN13),.WL(WL47));
sram_cell_6t_5 inst_cell_47_14 (.BL(BL14),.BLN(BLN14),.WL(WL47));
sram_cell_6t_5 inst_cell_47_15 (.BL(BL15),.BLN(BLN15),.WL(WL47));
sram_cell_6t_5 inst_cell_47_16 (.BL(BL16),.BLN(BLN16),.WL(WL47));
sram_cell_6t_5 inst_cell_47_17 (.BL(BL17),.BLN(BLN17),.WL(WL47));
sram_cell_6t_5 inst_cell_47_18 (.BL(BL18),.BLN(BLN18),.WL(WL47));
sram_cell_6t_5 inst_cell_47_19 (.BL(BL19),.BLN(BLN19),.WL(WL47));
sram_cell_6t_5 inst_cell_47_20 (.BL(BL20),.BLN(BLN20),.WL(WL47));
sram_cell_6t_5 inst_cell_47_21 (.BL(BL21),.BLN(BLN21),.WL(WL47));
sram_cell_6t_5 inst_cell_47_22 (.BL(BL22),.BLN(BLN22),.WL(WL47));
sram_cell_6t_5 inst_cell_47_23 (.BL(BL23),.BLN(BLN23),.WL(WL47));
sram_cell_6t_5 inst_cell_47_24 (.BL(BL24),.BLN(BLN24),.WL(WL47));
sram_cell_6t_5 inst_cell_47_25 (.BL(BL25),.BLN(BLN25),.WL(WL47));
sram_cell_6t_5 inst_cell_47_26 (.BL(BL26),.BLN(BLN26),.WL(WL47));
sram_cell_6t_5 inst_cell_47_27 (.BL(BL27),.BLN(BLN27),.WL(WL47));
sram_cell_6t_5 inst_cell_47_28 (.BL(BL28),.BLN(BLN28),.WL(WL47));
sram_cell_6t_5 inst_cell_47_29 (.BL(BL29),.BLN(BLN29),.WL(WL47));
sram_cell_6t_5 inst_cell_47_30 (.BL(BL30),.BLN(BLN30),.WL(WL47));
sram_cell_6t_5 inst_cell_47_31 (.BL(BL31),.BLN(BLN31),.WL(WL47));
sram_cell_6t_5 inst_cell_47_32 (.BL(BL32),.BLN(BLN32),.WL(WL47));
sram_cell_6t_5 inst_cell_47_33 (.BL(BL33),.BLN(BLN33),.WL(WL47));
sram_cell_6t_5 inst_cell_47_34 (.BL(BL34),.BLN(BLN34),.WL(WL47));
sram_cell_6t_5 inst_cell_47_35 (.BL(BL35),.BLN(BLN35),.WL(WL47));
sram_cell_6t_5 inst_cell_47_36 (.BL(BL36),.BLN(BLN36),.WL(WL47));
sram_cell_6t_5 inst_cell_47_37 (.BL(BL37),.BLN(BLN37),.WL(WL47));
sram_cell_6t_5 inst_cell_47_38 (.BL(BL38),.BLN(BLN38),.WL(WL47));
sram_cell_6t_5 inst_cell_47_39 (.BL(BL39),.BLN(BLN39),.WL(WL47));
sram_cell_6t_5 inst_cell_47_40 (.BL(BL40),.BLN(BLN40),.WL(WL47));
sram_cell_6t_5 inst_cell_47_41 (.BL(BL41),.BLN(BLN41),.WL(WL47));
sram_cell_6t_5 inst_cell_47_42 (.BL(BL42),.BLN(BLN42),.WL(WL47));
sram_cell_6t_5 inst_cell_47_43 (.BL(BL43),.BLN(BLN43),.WL(WL47));
sram_cell_6t_5 inst_cell_47_44 (.BL(BL44),.BLN(BLN44),.WL(WL47));
sram_cell_6t_5 inst_cell_47_45 (.BL(BL45),.BLN(BLN45),.WL(WL47));
sram_cell_6t_5 inst_cell_47_46 (.BL(BL46),.BLN(BLN46),.WL(WL47));
sram_cell_6t_5 inst_cell_47_47 (.BL(BL47),.BLN(BLN47),.WL(WL47));
sram_cell_6t_5 inst_cell_47_48 (.BL(BL48),.BLN(BLN48),.WL(WL47));
sram_cell_6t_5 inst_cell_47_49 (.BL(BL49),.BLN(BLN49),.WL(WL47));
sram_cell_6t_5 inst_cell_47_50 (.BL(BL50),.BLN(BLN50),.WL(WL47));
sram_cell_6t_5 inst_cell_47_51 (.BL(BL51),.BLN(BLN51),.WL(WL47));
sram_cell_6t_5 inst_cell_47_52 (.BL(BL52),.BLN(BLN52),.WL(WL47));
sram_cell_6t_5 inst_cell_47_53 (.BL(BL53),.BLN(BLN53),.WL(WL47));
sram_cell_6t_5 inst_cell_47_54 (.BL(BL54),.BLN(BLN54),.WL(WL47));
sram_cell_6t_5 inst_cell_47_55 (.BL(BL55),.BLN(BLN55),.WL(WL47));
sram_cell_6t_5 inst_cell_47_56 (.BL(BL56),.BLN(BLN56),.WL(WL47));
sram_cell_6t_5 inst_cell_47_57 (.BL(BL57),.BLN(BLN57),.WL(WL47));
sram_cell_6t_5 inst_cell_47_58 (.BL(BL58),.BLN(BLN58),.WL(WL47));
sram_cell_6t_5 inst_cell_47_59 (.BL(BL59),.BLN(BLN59),.WL(WL47));
sram_cell_6t_5 inst_cell_47_60 (.BL(BL60),.BLN(BLN60),.WL(WL47));
sram_cell_6t_5 inst_cell_47_61 (.BL(BL61),.BLN(BLN61),.WL(WL47));
sram_cell_6t_5 inst_cell_47_62 (.BL(BL62),.BLN(BLN62),.WL(WL47));
sram_cell_6t_5 inst_cell_47_63 (.BL(BL63),.BLN(BLN63),.WL(WL47));
sram_cell_6t_5 inst_cell_47_64 (.BL(BL64),.BLN(BLN64),.WL(WL47));
sram_cell_6t_5 inst_cell_47_65 (.BL(BL65),.BLN(BLN65),.WL(WL47));
sram_cell_6t_5 inst_cell_47_66 (.BL(BL66),.BLN(BLN66),.WL(WL47));
sram_cell_6t_5 inst_cell_47_67 (.BL(BL67),.BLN(BLN67),.WL(WL47));
sram_cell_6t_5 inst_cell_47_68 (.BL(BL68),.BLN(BLN68),.WL(WL47));
sram_cell_6t_5 inst_cell_47_69 (.BL(BL69),.BLN(BLN69),.WL(WL47));
sram_cell_6t_5 inst_cell_47_70 (.BL(BL70),.BLN(BLN70),.WL(WL47));
sram_cell_6t_5 inst_cell_47_71 (.BL(BL71),.BLN(BLN71),.WL(WL47));
sram_cell_6t_5 inst_cell_47_72 (.BL(BL72),.BLN(BLN72),.WL(WL47));
sram_cell_6t_5 inst_cell_47_73 (.BL(BL73),.BLN(BLN73),.WL(WL47));
sram_cell_6t_5 inst_cell_47_74 (.BL(BL74),.BLN(BLN74),.WL(WL47));
sram_cell_6t_5 inst_cell_47_75 (.BL(BL75),.BLN(BLN75),.WL(WL47));
sram_cell_6t_5 inst_cell_47_76 (.BL(BL76),.BLN(BLN76),.WL(WL47));
sram_cell_6t_5 inst_cell_47_77 (.BL(BL77),.BLN(BLN77),.WL(WL47));
sram_cell_6t_5 inst_cell_47_78 (.BL(BL78),.BLN(BLN78),.WL(WL47));
sram_cell_6t_5 inst_cell_47_79 (.BL(BL79),.BLN(BLN79),.WL(WL47));
sram_cell_6t_5 inst_cell_47_80 (.BL(BL80),.BLN(BLN80),.WL(WL47));
sram_cell_6t_5 inst_cell_47_81 (.BL(BL81),.BLN(BLN81),.WL(WL47));
sram_cell_6t_5 inst_cell_47_82 (.BL(BL82),.BLN(BLN82),.WL(WL47));
sram_cell_6t_5 inst_cell_47_83 (.BL(BL83),.BLN(BLN83),.WL(WL47));
sram_cell_6t_5 inst_cell_47_84 (.BL(BL84),.BLN(BLN84),.WL(WL47));
sram_cell_6t_5 inst_cell_47_85 (.BL(BL85),.BLN(BLN85),.WL(WL47));
sram_cell_6t_5 inst_cell_47_86 (.BL(BL86),.BLN(BLN86),.WL(WL47));
sram_cell_6t_5 inst_cell_47_87 (.BL(BL87),.BLN(BLN87),.WL(WL47));
sram_cell_6t_5 inst_cell_47_88 (.BL(BL88),.BLN(BLN88),.WL(WL47));
sram_cell_6t_5 inst_cell_47_89 (.BL(BL89),.BLN(BLN89),.WL(WL47));
sram_cell_6t_5 inst_cell_47_90 (.BL(BL90),.BLN(BLN90),.WL(WL47));
sram_cell_6t_5 inst_cell_47_91 (.BL(BL91),.BLN(BLN91),.WL(WL47));
sram_cell_6t_5 inst_cell_47_92 (.BL(BL92),.BLN(BLN92),.WL(WL47));
sram_cell_6t_5 inst_cell_47_93 (.BL(BL93),.BLN(BLN93),.WL(WL47));
sram_cell_6t_5 inst_cell_47_94 (.BL(BL94),.BLN(BLN94),.WL(WL47));
sram_cell_6t_5 inst_cell_47_95 (.BL(BL95),.BLN(BLN95),.WL(WL47));
sram_cell_6t_5 inst_cell_47_96 (.BL(BL96),.BLN(BLN96),.WL(WL47));
sram_cell_6t_5 inst_cell_47_97 (.BL(BL97),.BLN(BLN97),.WL(WL47));
sram_cell_6t_5 inst_cell_47_98 (.BL(BL98),.BLN(BLN98),.WL(WL47));
sram_cell_6t_5 inst_cell_47_99 (.BL(BL99),.BLN(BLN99),.WL(WL47));
sram_cell_6t_5 inst_cell_47_100 (.BL(BL100),.BLN(BLN100),.WL(WL47));
sram_cell_6t_5 inst_cell_47_101 (.BL(BL101),.BLN(BLN101),.WL(WL47));
sram_cell_6t_5 inst_cell_47_102 (.BL(BL102),.BLN(BLN102),.WL(WL47));
sram_cell_6t_5 inst_cell_47_103 (.BL(BL103),.BLN(BLN103),.WL(WL47));
sram_cell_6t_5 inst_cell_47_104 (.BL(BL104),.BLN(BLN104),.WL(WL47));
sram_cell_6t_5 inst_cell_47_105 (.BL(BL105),.BLN(BLN105),.WL(WL47));
sram_cell_6t_5 inst_cell_47_106 (.BL(BL106),.BLN(BLN106),.WL(WL47));
sram_cell_6t_5 inst_cell_47_107 (.BL(BL107),.BLN(BLN107),.WL(WL47));
sram_cell_6t_5 inst_cell_47_108 (.BL(BL108),.BLN(BLN108),.WL(WL47));
sram_cell_6t_5 inst_cell_47_109 (.BL(BL109),.BLN(BLN109),.WL(WL47));
sram_cell_6t_5 inst_cell_47_110 (.BL(BL110),.BLN(BLN110),.WL(WL47));
sram_cell_6t_5 inst_cell_47_111 (.BL(BL111),.BLN(BLN111),.WL(WL47));
sram_cell_6t_5 inst_cell_47_112 (.BL(BL112),.BLN(BLN112),.WL(WL47));
sram_cell_6t_5 inst_cell_47_113 (.BL(BL113),.BLN(BLN113),.WL(WL47));
sram_cell_6t_5 inst_cell_47_114 (.BL(BL114),.BLN(BLN114),.WL(WL47));
sram_cell_6t_5 inst_cell_47_115 (.BL(BL115),.BLN(BLN115),.WL(WL47));
sram_cell_6t_5 inst_cell_47_116 (.BL(BL116),.BLN(BLN116),.WL(WL47));
sram_cell_6t_5 inst_cell_47_117 (.BL(BL117),.BLN(BLN117),.WL(WL47));
sram_cell_6t_5 inst_cell_47_118 (.BL(BL118),.BLN(BLN118),.WL(WL47));
sram_cell_6t_5 inst_cell_47_119 (.BL(BL119),.BLN(BLN119),.WL(WL47));
sram_cell_6t_5 inst_cell_47_120 (.BL(BL120),.BLN(BLN120),.WL(WL47));
sram_cell_6t_5 inst_cell_47_121 (.BL(BL121),.BLN(BLN121),.WL(WL47));
sram_cell_6t_5 inst_cell_47_122 (.BL(BL122),.BLN(BLN122),.WL(WL47));
sram_cell_6t_5 inst_cell_47_123 (.BL(BL123),.BLN(BLN123),.WL(WL47));
sram_cell_6t_5 inst_cell_47_124 (.BL(BL124),.BLN(BLN124),.WL(WL47));
sram_cell_6t_5 inst_cell_47_125 (.BL(BL125),.BLN(BLN125),.WL(WL47));
sram_cell_6t_5 inst_cell_47_126 (.BL(BL126),.BLN(BLN126),.WL(WL47));
sram_cell_6t_5 inst_cell_47_127 (.BL(BL127),.BLN(BLN127),.WL(WL47));
sram_cell_6t_5 inst_cell_48_0 (.BL(BL0),.BLN(BLN0),.WL(WL48));
sram_cell_6t_5 inst_cell_48_1 (.BL(BL1),.BLN(BLN1),.WL(WL48));
sram_cell_6t_5 inst_cell_48_2 (.BL(BL2),.BLN(BLN2),.WL(WL48));
sram_cell_6t_5 inst_cell_48_3 (.BL(BL3),.BLN(BLN3),.WL(WL48));
sram_cell_6t_5 inst_cell_48_4 (.BL(BL4),.BLN(BLN4),.WL(WL48));
sram_cell_6t_5 inst_cell_48_5 (.BL(BL5),.BLN(BLN5),.WL(WL48));
sram_cell_6t_5 inst_cell_48_6 (.BL(BL6),.BLN(BLN6),.WL(WL48));
sram_cell_6t_5 inst_cell_48_7 (.BL(BL7),.BLN(BLN7),.WL(WL48));
sram_cell_6t_5 inst_cell_48_8 (.BL(BL8),.BLN(BLN8),.WL(WL48));
sram_cell_6t_5 inst_cell_48_9 (.BL(BL9),.BLN(BLN9),.WL(WL48));
sram_cell_6t_5 inst_cell_48_10 (.BL(BL10),.BLN(BLN10),.WL(WL48));
sram_cell_6t_5 inst_cell_48_11 (.BL(BL11),.BLN(BLN11),.WL(WL48));
sram_cell_6t_5 inst_cell_48_12 (.BL(BL12),.BLN(BLN12),.WL(WL48));
sram_cell_6t_5 inst_cell_48_13 (.BL(BL13),.BLN(BLN13),.WL(WL48));
sram_cell_6t_5 inst_cell_48_14 (.BL(BL14),.BLN(BLN14),.WL(WL48));
sram_cell_6t_5 inst_cell_48_15 (.BL(BL15),.BLN(BLN15),.WL(WL48));
sram_cell_6t_5 inst_cell_48_16 (.BL(BL16),.BLN(BLN16),.WL(WL48));
sram_cell_6t_5 inst_cell_48_17 (.BL(BL17),.BLN(BLN17),.WL(WL48));
sram_cell_6t_5 inst_cell_48_18 (.BL(BL18),.BLN(BLN18),.WL(WL48));
sram_cell_6t_5 inst_cell_48_19 (.BL(BL19),.BLN(BLN19),.WL(WL48));
sram_cell_6t_5 inst_cell_48_20 (.BL(BL20),.BLN(BLN20),.WL(WL48));
sram_cell_6t_5 inst_cell_48_21 (.BL(BL21),.BLN(BLN21),.WL(WL48));
sram_cell_6t_5 inst_cell_48_22 (.BL(BL22),.BLN(BLN22),.WL(WL48));
sram_cell_6t_5 inst_cell_48_23 (.BL(BL23),.BLN(BLN23),.WL(WL48));
sram_cell_6t_5 inst_cell_48_24 (.BL(BL24),.BLN(BLN24),.WL(WL48));
sram_cell_6t_5 inst_cell_48_25 (.BL(BL25),.BLN(BLN25),.WL(WL48));
sram_cell_6t_5 inst_cell_48_26 (.BL(BL26),.BLN(BLN26),.WL(WL48));
sram_cell_6t_5 inst_cell_48_27 (.BL(BL27),.BLN(BLN27),.WL(WL48));
sram_cell_6t_5 inst_cell_48_28 (.BL(BL28),.BLN(BLN28),.WL(WL48));
sram_cell_6t_5 inst_cell_48_29 (.BL(BL29),.BLN(BLN29),.WL(WL48));
sram_cell_6t_5 inst_cell_48_30 (.BL(BL30),.BLN(BLN30),.WL(WL48));
sram_cell_6t_5 inst_cell_48_31 (.BL(BL31),.BLN(BLN31),.WL(WL48));
sram_cell_6t_5 inst_cell_48_32 (.BL(BL32),.BLN(BLN32),.WL(WL48));
sram_cell_6t_5 inst_cell_48_33 (.BL(BL33),.BLN(BLN33),.WL(WL48));
sram_cell_6t_5 inst_cell_48_34 (.BL(BL34),.BLN(BLN34),.WL(WL48));
sram_cell_6t_5 inst_cell_48_35 (.BL(BL35),.BLN(BLN35),.WL(WL48));
sram_cell_6t_5 inst_cell_48_36 (.BL(BL36),.BLN(BLN36),.WL(WL48));
sram_cell_6t_5 inst_cell_48_37 (.BL(BL37),.BLN(BLN37),.WL(WL48));
sram_cell_6t_5 inst_cell_48_38 (.BL(BL38),.BLN(BLN38),.WL(WL48));
sram_cell_6t_5 inst_cell_48_39 (.BL(BL39),.BLN(BLN39),.WL(WL48));
sram_cell_6t_5 inst_cell_48_40 (.BL(BL40),.BLN(BLN40),.WL(WL48));
sram_cell_6t_5 inst_cell_48_41 (.BL(BL41),.BLN(BLN41),.WL(WL48));
sram_cell_6t_5 inst_cell_48_42 (.BL(BL42),.BLN(BLN42),.WL(WL48));
sram_cell_6t_5 inst_cell_48_43 (.BL(BL43),.BLN(BLN43),.WL(WL48));
sram_cell_6t_5 inst_cell_48_44 (.BL(BL44),.BLN(BLN44),.WL(WL48));
sram_cell_6t_5 inst_cell_48_45 (.BL(BL45),.BLN(BLN45),.WL(WL48));
sram_cell_6t_5 inst_cell_48_46 (.BL(BL46),.BLN(BLN46),.WL(WL48));
sram_cell_6t_5 inst_cell_48_47 (.BL(BL47),.BLN(BLN47),.WL(WL48));
sram_cell_6t_5 inst_cell_48_48 (.BL(BL48),.BLN(BLN48),.WL(WL48));
sram_cell_6t_5 inst_cell_48_49 (.BL(BL49),.BLN(BLN49),.WL(WL48));
sram_cell_6t_5 inst_cell_48_50 (.BL(BL50),.BLN(BLN50),.WL(WL48));
sram_cell_6t_5 inst_cell_48_51 (.BL(BL51),.BLN(BLN51),.WL(WL48));
sram_cell_6t_5 inst_cell_48_52 (.BL(BL52),.BLN(BLN52),.WL(WL48));
sram_cell_6t_5 inst_cell_48_53 (.BL(BL53),.BLN(BLN53),.WL(WL48));
sram_cell_6t_5 inst_cell_48_54 (.BL(BL54),.BLN(BLN54),.WL(WL48));
sram_cell_6t_5 inst_cell_48_55 (.BL(BL55),.BLN(BLN55),.WL(WL48));
sram_cell_6t_5 inst_cell_48_56 (.BL(BL56),.BLN(BLN56),.WL(WL48));
sram_cell_6t_5 inst_cell_48_57 (.BL(BL57),.BLN(BLN57),.WL(WL48));
sram_cell_6t_5 inst_cell_48_58 (.BL(BL58),.BLN(BLN58),.WL(WL48));
sram_cell_6t_5 inst_cell_48_59 (.BL(BL59),.BLN(BLN59),.WL(WL48));
sram_cell_6t_5 inst_cell_48_60 (.BL(BL60),.BLN(BLN60),.WL(WL48));
sram_cell_6t_5 inst_cell_48_61 (.BL(BL61),.BLN(BLN61),.WL(WL48));
sram_cell_6t_5 inst_cell_48_62 (.BL(BL62),.BLN(BLN62),.WL(WL48));
sram_cell_6t_5 inst_cell_48_63 (.BL(BL63),.BLN(BLN63),.WL(WL48));
sram_cell_6t_5 inst_cell_48_64 (.BL(BL64),.BLN(BLN64),.WL(WL48));
sram_cell_6t_5 inst_cell_48_65 (.BL(BL65),.BLN(BLN65),.WL(WL48));
sram_cell_6t_5 inst_cell_48_66 (.BL(BL66),.BLN(BLN66),.WL(WL48));
sram_cell_6t_5 inst_cell_48_67 (.BL(BL67),.BLN(BLN67),.WL(WL48));
sram_cell_6t_5 inst_cell_48_68 (.BL(BL68),.BLN(BLN68),.WL(WL48));
sram_cell_6t_5 inst_cell_48_69 (.BL(BL69),.BLN(BLN69),.WL(WL48));
sram_cell_6t_5 inst_cell_48_70 (.BL(BL70),.BLN(BLN70),.WL(WL48));
sram_cell_6t_5 inst_cell_48_71 (.BL(BL71),.BLN(BLN71),.WL(WL48));
sram_cell_6t_5 inst_cell_48_72 (.BL(BL72),.BLN(BLN72),.WL(WL48));
sram_cell_6t_5 inst_cell_48_73 (.BL(BL73),.BLN(BLN73),.WL(WL48));
sram_cell_6t_5 inst_cell_48_74 (.BL(BL74),.BLN(BLN74),.WL(WL48));
sram_cell_6t_5 inst_cell_48_75 (.BL(BL75),.BLN(BLN75),.WL(WL48));
sram_cell_6t_5 inst_cell_48_76 (.BL(BL76),.BLN(BLN76),.WL(WL48));
sram_cell_6t_5 inst_cell_48_77 (.BL(BL77),.BLN(BLN77),.WL(WL48));
sram_cell_6t_5 inst_cell_48_78 (.BL(BL78),.BLN(BLN78),.WL(WL48));
sram_cell_6t_5 inst_cell_48_79 (.BL(BL79),.BLN(BLN79),.WL(WL48));
sram_cell_6t_5 inst_cell_48_80 (.BL(BL80),.BLN(BLN80),.WL(WL48));
sram_cell_6t_5 inst_cell_48_81 (.BL(BL81),.BLN(BLN81),.WL(WL48));
sram_cell_6t_5 inst_cell_48_82 (.BL(BL82),.BLN(BLN82),.WL(WL48));
sram_cell_6t_5 inst_cell_48_83 (.BL(BL83),.BLN(BLN83),.WL(WL48));
sram_cell_6t_5 inst_cell_48_84 (.BL(BL84),.BLN(BLN84),.WL(WL48));
sram_cell_6t_5 inst_cell_48_85 (.BL(BL85),.BLN(BLN85),.WL(WL48));
sram_cell_6t_5 inst_cell_48_86 (.BL(BL86),.BLN(BLN86),.WL(WL48));
sram_cell_6t_5 inst_cell_48_87 (.BL(BL87),.BLN(BLN87),.WL(WL48));
sram_cell_6t_5 inst_cell_48_88 (.BL(BL88),.BLN(BLN88),.WL(WL48));
sram_cell_6t_5 inst_cell_48_89 (.BL(BL89),.BLN(BLN89),.WL(WL48));
sram_cell_6t_5 inst_cell_48_90 (.BL(BL90),.BLN(BLN90),.WL(WL48));
sram_cell_6t_5 inst_cell_48_91 (.BL(BL91),.BLN(BLN91),.WL(WL48));
sram_cell_6t_5 inst_cell_48_92 (.BL(BL92),.BLN(BLN92),.WL(WL48));
sram_cell_6t_5 inst_cell_48_93 (.BL(BL93),.BLN(BLN93),.WL(WL48));
sram_cell_6t_5 inst_cell_48_94 (.BL(BL94),.BLN(BLN94),.WL(WL48));
sram_cell_6t_5 inst_cell_48_95 (.BL(BL95),.BLN(BLN95),.WL(WL48));
sram_cell_6t_5 inst_cell_48_96 (.BL(BL96),.BLN(BLN96),.WL(WL48));
sram_cell_6t_5 inst_cell_48_97 (.BL(BL97),.BLN(BLN97),.WL(WL48));
sram_cell_6t_5 inst_cell_48_98 (.BL(BL98),.BLN(BLN98),.WL(WL48));
sram_cell_6t_5 inst_cell_48_99 (.BL(BL99),.BLN(BLN99),.WL(WL48));
sram_cell_6t_5 inst_cell_48_100 (.BL(BL100),.BLN(BLN100),.WL(WL48));
sram_cell_6t_5 inst_cell_48_101 (.BL(BL101),.BLN(BLN101),.WL(WL48));
sram_cell_6t_5 inst_cell_48_102 (.BL(BL102),.BLN(BLN102),.WL(WL48));
sram_cell_6t_5 inst_cell_48_103 (.BL(BL103),.BLN(BLN103),.WL(WL48));
sram_cell_6t_5 inst_cell_48_104 (.BL(BL104),.BLN(BLN104),.WL(WL48));
sram_cell_6t_5 inst_cell_48_105 (.BL(BL105),.BLN(BLN105),.WL(WL48));
sram_cell_6t_5 inst_cell_48_106 (.BL(BL106),.BLN(BLN106),.WL(WL48));
sram_cell_6t_5 inst_cell_48_107 (.BL(BL107),.BLN(BLN107),.WL(WL48));
sram_cell_6t_5 inst_cell_48_108 (.BL(BL108),.BLN(BLN108),.WL(WL48));
sram_cell_6t_5 inst_cell_48_109 (.BL(BL109),.BLN(BLN109),.WL(WL48));
sram_cell_6t_5 inst_cell_48_110 (.BL(BL110),.BLN(BLN110),.WL(WL48));
sram_cell_6t_5 inst_cell_48_111 (.BL(BL111),.BLN(BLN111),.WL(WL48));
sram_cell_6t_5 inst_cell_48_112 (.BL(BL112),.BLN(BLN112),.WL(WL48));
sram_cell_6t_5 inst_cell_48_113 (.BL(BL113),.BLN(BLN113),.WL(WL48));
sram_cell_6t_5 inst_cell_48_114 (.BL(BL114),.BLN(BLN114),.WL(WL48));
sram_cell_6t_5 inst_cell_48_115 (.BL(BL115),.BLN(BLN115),.WL(WL48));
sram_cell_6t_5 inst_cell_48_116 (.BL(BL116),.BLN(BLN116),.WL(WL48));
sram_cell_6t_5 inst_cell_48_117 (.BL(BL117),.BLN(BLN117),.WL(WL48));
sram_cell_6t_5 inst_cell_48_118 (.BL(BL118),.BLN(BLN118),.WL(WL48));
sram_cell_6t_5 inst_cell_48_119 (.BL(BL119),.BLN(BLN119),.WL(WL48));
sram_cell_6t_5 inst_cell_48_120 (.BL(BL120),.BLN(BLN120),.WL(WL48));
sram_cell_6t_5 inst_cell_48_121 (.BL(BL121),.BLN(BLN121),.WL(WL48));
sram_cell_6t_5 inst_cell_48_122 (.BL(BL122),.BLN(BLN122),.WL(WL48));
sram_cell_6t_5 inst_cell_48_123 (.BL(BL123),.BLN(BLN123),.WL(WL48));
sram_cell_6t_5 inst_cell_48_124 (.BL(BL124),.BLN(BLN124),.WL(WL48));
sram_cell_6t_5 inst_cell_48_125 (.BL(BL125),.BLN(BLN125),.WL(WL48));
sram_cell_6t_5 inst_cell_48_126 (.BL(BL126),.BLN(BLN126),.WL(WL48));
sram_cell_6t_5 inst_cell_48_127 (.BL(BL127),.BLN(BLN127),.WL(WL48));
sram_cell_6t_5 inst_cell_49_0 (.BL(BL0),.BLN(BLN0),.WL(WL49));
sram_cell_6t_5 inst_cell_49_1 (.BL(BL1),.BLN(BLN1),.WL(WL49));
sram_cell_6t_5 inst_cell_49_2 (.BL(BL2),.BLN(BLN2),.WL(WL49));
sram_cell_6t_5 inst_cell_49_3 (.BL(BL3),.BLN(BLN3),.WL(WL49));
sram_cell_6t_5 inst_cell_49_4 (.BL(BL4),.BLN(BLN4),.WL(WL49));
sram_cell_6t_5 inst_cell_49_5 (.BL(BL5),.BLN(BLN5),.WL(WL49));
sram_cell_6t_5 inst_cell_49_6 (.BL(BL6),.BLN(BLN6),.WL(WL49));
sram_cell_6t_5 inst_cell_49_7 (.BL(BL7),.BLN(BLN7),.WL(WL49));
sram_cell_6t_5 inst_cell_49_8 (.BL(BL8),.BLN(BLN8),.WL(WL49));
sram_cell_6t_5 inst_cell_49_9 (.BL(BL9),.BLN(BLN9),.WL(WL49));
sram_cell_6t_5 inst_cell_49_10 (.BL(BL10),.BLN(BLN10),.WL(WL49));
sram_cell_6t_5 inst_cell_49_11 (.BL(BL11),.BLN(BLN11),.WL(WL49));
sram_cell_6t_5 inst_cell_49_12 (.BL(BL12),.BLN(BLN12),.WL(WL49));
sram_cell_6t_5 inst_cell_49_13 (.BL(BL13),.BLN(BLN13),.WL(WL49));
sram_cell_6t_5 inst_cell_49_14 (.BL(BL14),.BLN(BLN14),.WL(WL49));
sram_cell_6t_5 inst_cell_49_15 (.BL(BL15),.BLN(BLN15),.WL(WL49));
sram_cell_6t_5 inst_cell_49_16 (.BL(BL16),.BLN(BLN16),.WL(WL49));
sram_cell_6t_5 inst_cell_49_17 (.BL(BL17),.BLN(BLN17),.WL(WL49));
sram_cell_6t_5 inst_cell_49_18 (.BL(BL18),.BLN(BLN18),.WL(WL49));
sram_cell_6t_5 inst_cell_49_19 (.BL(BL19),.BLN(BLN19),.WL(WL49));
sram_cell_6t_5 inst_cell_49_20 (.BL(BL20),.BLN(BLN20),.WL(WL49));
sram_cell_6t_5 inst_cell_49_21 (.BL(BL21),.BLN(BLN21),.WL(WL49));
sram_cell_6t_5 inst_cell_49_22 (.BL(BL22),.BLN(BLN22),.WL(WL49));
sram_cell_6t_5 inst_cell_49_23 (.BL(BL23),.BLN(BLN23),.WL(WL49));
sram_cell_6t_5 inst_cell_49_24 (.BL(BL24),.BLN(BLN24),.WL(WL49));
sram_cell_6t_5 inst_cell_49_25 (.BL(BL25),.BLN(BLN25),.WL(WL49));
sram_cell_6t_5 inst_cell_49_26 (.BL(BL26),.BLN(BLN26),.WL(WL49));
sram_cell_6t_5 inst_cell_49_27 (.BL(BL27),.BLN(BLN27),.WL(WL49));
sram_cell_6t_5 inst_cell_49_28 (.BL(BL28),.BLN(BLN28),.WL(WL49));
sram_cell_6t_5 inst_cell_49_29 (.BL(BL29),.BLN(BLN29),.WL(WL49));
sram_cell_6t_5 inst_cell_49_30 (.BL(BL30),.BLN(BLN30),.WL(WL49));
sram_cell_6t_5 inst_cell_49_31 (.BL(BL31),.BLN(BLN31),.WL(WL49));
sram_cell_6t_5 inst_cell_49_32 (.BL(BL32),.BLN(BLN32),.WL(WL49));
sram_cell_6t_5 inst_cell_49_33 (.BL(BL33),.BLN(BLN33),.WL(WL49));
sram_cell_6t_5 inst_cell_49_34 (.BL(BL34),.BLN(BLN34),.WL(WL49));
sram_cell_6t_5 inst_cell_49_35 (.BL(BL35),.BLN(BLN35),.WL(WL49));
sram_cell_6t_5 inst_cell_49_36 (.BL(BL36),.BLN(BLN36),.WL(WL49));
sram_cell_6t_5 inst_cell_49_37 (.BL(BL37),.BLN(BLN37),.WL(WL49));
sram_cell_6t_5 inst_cell_49_38 (.BL(BL38),.BLN(BLN38),.WL(WL49));
sram_cell_6t_5 inst_cell_49_39 (.BL(BL39),.BLN(BLN39),.WL(WL49));
sram_cell_6t_5 inst_cell_49_40 (.BL(BL40),.BLN(BLN40),.WL(WL49));
sram_cell_6t_5 inst_cell_49_41 (.BL(BL41),.BLN(BLN41),.WL(WL49));
sram_cell_6t_5 inst_cell_49_42 (.BL(BL42),.BLN(BLN42),.WL(WL49));
sram_cell_6t_5 inst_cell_49_43 (.BL(BL43),.BLN(BLN43),.WL(WL49));
sram_cell_6t_5 inst_cell_49_44 (.BL(BL44),.BLN(BLN44),.WL(WL49));
sram_cell_6t_5 inst_cell_49_45 (.BL(BL45),.BLN(BLN45),.WL(WL49));
sram_cell_6t_5 inst_cell_49_46 (.BL(BL46),.BLN(BLN46),.WL(WL49));
sram_cell_6t_5 inst_cell_49_47 (.BL(BL47),.BLN(BLN47),.WL(WL49));
sram_cell_6t_5 inst_cell_49_48 (.BL(BL48),.BLN(BLN48),.WL(WL49));
sram_cell_6t_5 inst_cell_49_49 (.BL(BL49),.BLN(BLN49),.WL(WL49));
sram_cell_6t_5 inst_cell_49_50 (.BL(BL50),.BLN(BLN50),.WL(WL49));
sram_cell_6t_5 inst_cell_49_51 (.BL(BL51),.BLN(BLN51),.WL(WL49));
sram_cell_6t_5 inst_cell_49_52 (.BL(BL52),.BLN(BLN52),.WL(WL49));
sram_cell_6t_5 inst_cell_49_53 (.BL(BL53),.BLN(BLN53),.WL(WL49));
sram_cell_6t_5 inst_cell_49_54 (.BL(BL54),.BLN(BLN54),.WL(WL49));
sram_cell_6t_5 inst_cell_49_55 (.BL(BL55),.BLN(BLN55),.WL(WL49));
sram_cell_6t_5 inst_cell_49_56 (.BL(BL56),.BLN(BLN56),.WL(WL49));
sram_cell_6t_5 inst_cell_49_57 (.BL(BL57),.BLN(BLN57),.WL(WL49));
sram_cell_6t_5 inst_cell_49_58 (.BL(BL58),.BLN(BLN58),.WL(WL49));
sram_cell_6t_5 inst_cell_49_59 (.BL(BL59),.BLN(BLN59),.WL(WL49));
sram_cell_6t_5 inst_cell_49_60 (.BL(BL60),.BLN(BLN60),.WL(WL49));
sram_cell_6t_5 inst_cell_49_61 (.BL(BL61),.BLN(BLN61),.WL(WL49));
sram_cell_6t_5 inst_cell_49_62 (.BL(BL62),.BLN(BLN62),.WL(WL49));
sram_cell_6t_5 inst_cell_49_63 (.BL(BL63),.BLN(BLN63),.WL(WL49));
sram_cell_6t_5 inst_cell_49_64 (.BL(BL64),.BLN(BLN64),.WL(WL49));
sram_cell_6t_5 inst_cell_49_65 (.BL(BL65),.BLN(BLN65),.WL(WL49));
sram_cell_6t_5 inst_cell_49_66 (.BL(BL66),.BLN(BLN66),.WL(WL49));
sram_cell_6t_5 inst_cell_49_67 (.BL(BL67),.BLN(BLN67),.WL(WL49));
sram_cell_6t_5 inst_cell_49_68 (.BL(BL68),.BLN(BLN68),.WL(WL49));
sram_cell_6t_5 inst_cell_49_69 (.BL(BL69),.BLN(BLN69),.WL(WL49));
sram_cell_6t_5 inst_cell_49_70 (.BL(BL70),.BLN(BLN70),.WL(WL49));
sram_cell_6t_5 inst_cell_49_71 (.BL(BL71),.BLN(BLN71),.WL(WL49));
sram_cell_6t_5 inst_cell_49_72 (.BL(BL72),.BLN(BLN72),.WL(WL49));
sram_cell_6t_5 inst_cell_49_73 (.BL(BL73),.BLN(BLN73),.WL(WL49));
sram_cell_6t_5 inst_cell_49_74 (.BL(BL74),.BLN(BLN74),.WL(WL49));
sram_cell_6t_5 inst_cell_49_75 (.BL(BL75),.BLN(BLN75),.WL(WL49));
sram_cell_6t_5 inst_cell_49_76 (.BL(BL76),.BLN(BLN76),.WL(WL49));
sram_cell_6t_5 inst_cell_49_77 (.BL(BL77),.BLN(BLN77),.WL(WL49));
sram_cell_6t_5 inst_cell_49_78 (.BL(BL78),.BLN(BLN78),.WL(WL49));
sram_cell_6t_5 inst_cell_49_79 (.BL(BL79),.BLN(BLN79),.WL(WL49));
sram_cell_6t_5 inst_cell_49_80 (.BL(BL80),.BLN(BLN80),.WL(WL49));
sram_cell_6t_5 inst_cell_49_81 (.BL(BL81),.BLN(BLN81),.WL(WL49));
sram_cell_6t_5 inst_cell_49_82 (.BL(BL82),.BLN(BLN82),.WL(WL49));
sram_cell_6t_5 inst_cell_49_83 (.BL(BL83),.BLN(BLN83),.WL(WL49));
sram_cell_6t_5 inst_cell_49_84 (.BL(BL84),.BLN(BLN84),.WL(WL49));
sram_cell_6t_5 inst_cell_49_85 (.BL(BL85),.BLN(BLN85),.WL(WL49));
sram_cell_6t_5 inst_cell_49_86 (.BL(BL86),.BLN(BLN86),.WL(WL49));
sram_cell_6t_5 inst_cell_49_87 (.BL(BL87),.BLN(BLN87),.WL(WL49));
sram_cell_6t_5 inst_cell_49_88 (.BL(BL88),.BLN(BLN88),.WL(WL49));
sram_cell_6t_5 inst_cell_49_89 (.BL(BL89),.BLN(BLN89),.WL(WL49));
sram_cell_6t_5 inst_cell_49_90 (.BL(BL90),.BLN(BLN90),.WL(WL49));
sram_cell_6t_5 inst_cell_49_91 (.BL(BL91),.BLN(BLN91),.WL(WL49));
sram_cell_6t_5 inst_cell_49_92 (.BL(BL92),.BLN(BLN92),.WL(WL49));
sram_cell_6t_5 inst_cell_49_93 (.BL(BL93),.BLN(BLN93),.WL(WL49));
sram_cell_6t_5 inst_cell_49_94 (.BL(BL94),.BLN(BLN94),.WL(WL49));
sram_cell_6t_5 inst_cell_49_95 (.BL(BL95),.BLN(BLN95),.WL(WL49));
sram_cell_6t_5 inst_cell_49_96 (.BL(BL96),.BLN(BLN96),.WL(WL49));
sram_cell_6t_5 inst_cell_49_97 (.BL(BL97),.BLN(BLN97),.WL(WL49));
sram_cell_6t_5 inst_cell_49_98 (.BL(BL98),.BLN(BLN98),.WL(WL49));
sram_cell_6t_5 inst_cell_49_99 (.BL(BL99),.BLN(BLN99),.WL(WL49));
sram_cell_6t_5 inst_cell_49_100 (.BL(BL100),.BLN(BLN100),.WL(WL49));
sram_cell_6t_5 inst_cell_49_101 (.BL(BL101),.BLN(BLN101),.WL(WL49));
sram_cell_6t_5 inst_cell_49_102 (.BL(BL102),.BLN(BLN102),.WL(WL49));
sram_cell_6t_5 inst_cell_49_103 (.BL(BL103),.BLN(BLN103),.WL(WL49));
sram_cell_6t_5 inst_cell_49_104 (.BL(BL104),.BLN(BLN104),.WL(WL49));
sram_cell_6t_5 inst_cell_49_105 (.BL(BL105),.BLN(BLN105),.WL(WL49));
sram_cell_6t_5 inst_cell_49_106 (.BL(BL106),.BLN(BLN106),.WL(WL49));
sram_cell_6t_5 inst_cell_49_107 (.BL(BL107),.BLN(BLN107),.WL(WL49));
sram_cell_6t_5 inst_cell_49_108 (.BL(BL108),.BLN(BLN108),.WL(WL49));
sram_cell_6t_5 inst_cell_49_109 (.BL(BL109),.BLN(BLN109),.WL(WL49));
sram_cell_6t_5 inst_cell_49_110 (.BL(BL110),.BLN(BLN110),.WL(WL49));
sram_cell_6t_5 inst_cell_49_111 (.BL(BL111),.BLN(BLN111),.WL(WL49));
sram_cell_6t_5 inst_cell_49_112 (.BL(BL112),.BLN(BLN112),.WL(WL49));
sram_cell_6t_5 inst_cell_49_113 (.BL(BL113),.BLN(BLN113),.WL(WL49));
sram_cell_6t_5 inst_cell_49_114 (.BL(BL114),.BLN(BLN114),.WL(WL49));
sram_cell_6t_5 inst_cell_49_115 (.BL(BL115),.BLN(BLN115),.WL(WL49));
sram_cell_6t_5 inst_cell_49_116 (.BL(BL116),.BLN(BLN116),.WL(WL49));
sram_cell_6t_5 inst_cell_49_117 (.BL(BL117),.BLN(BLN117),.WL(WL49));
sram_cell_6t_5 inst_cell_49_118 (.BL(BL118),.BLN(BLN118),.WL(WL49));
sram_cell_6t_5 inst_cell_49_119 (.BL(BL119),.BLN(BLN119),.WL(WL49));
sram_cell_6t_5 inst_cell_49_120 (.BL(BL120),.BLN(BLN120),.WL(WL49));
sram_cell_6t_5 inst_cell_49_121 (.BL(BL121),.BLN(BLN121),.WL(WL49));
sram_cell_6t_5 inst_cell_49_122 (.BL(BL122),.BLN(BLN122),.WL(WL49));
sram_cell_6t_5 inst_cell_49_123 (.BL(BL123),.BLN(BLN123),.WL(WL49));
sram_cell_6t_5 inst_cell_49_124 (.BL(BL124),.BLN(BLN124),.WL(WL49));
sram_cell_6t_5 inst_cell_49_125 (.BL(BL125),.BLN(BLN125),.WL(WL49));
sram_cell_6t_5 inst_cell_49_126 (.BL(BL126),.BLN(BLN126),.WL(WL49));
sram_cell_6t_5 inst_cell_49_127 (.BL(BL127),.BLN(BLN127),.WL(WL49));
sram_cell_6t_5 inst_cell_50_0 (.BL(BL0),.BLN(BLN0),.WL(WL50));
sram_cell_6t_5 inst_cell_50_1 (.BL(BL1),.BLN(BLN1),.WL(WL50));
sram_cell_6t_5 inst_cell_50_2 (.BL(BL2),.BLN(BLN2),.WL(WL50));
sram_cell_6t_5 inst_cell_50_3 (.BL(BL3),.BLN(BLN3),.WL(WL50));
sram_cell_6t_5 inst_cell_50_4 (.BL(BL4),.BLN(BLN4),.WL(WL50));
sram_cell_6t_5 inst_cell_50_5 (.BL(BL5),.BLN(BLN5),.WL(WL50));
sram_cell_6t_5 inst_cell_50_6 (.BL(BL6),.BLN(BLN6),.WL(WL50));
sram_cell_6t_5 inst_cell_50_7 (.BL(BL7),.BLN(BLN7),.WL(WL50));
sram_cell_6t_5 inst_cell_50_8 (.BL(BL8),.BLN(BLN8),.WL(WL50));
sram_cell_6t_5 inst_cell_50_9 (.BL(BL9),.BLN(BLN9),.WL(WL50));
sram_cell_6t_5 inst_cell_50_10 (.BL(BL10),.BLN(BLN10),.WL(WL50));
sram_cell_6t_5 inst_cell_50_11 (.BL(BL11),.BLN(BLN11),.WL(WL50));
sram_cell_6t_5 inst_cell_50_12 (.BL(BL12),.BLN(BLN12),.WL(WL50));
sram_cell_6t_5 inst_cell_50_13 (.BL(BL13),.BLN(BLN13),.WL(WL50));
sram_cell_6t_5 inst_cell_50_14 (.BL(BL14),.BLN(BLN14),.WL(WL50));
sram_cell_6t_5 inst_cell_50_15 (.BL(BL15),.BLN(BLN15),.WL(WL50));
sram_cell_6t_5 inst_cell_50_16 (.BL(BL16),.BLN(BLN16),.WL(WL50));
sram_cell_6t_5 inst_cell_50_17 (.BL(BL17),.BLN(BLN17),.WL(WL50));
sram_cell_6t_5 inst_cell_50_18 (.BL(BL18),.BLN(BLN18),.WL(WL50));
sram_cell_6t_5 inst_cell_50_19 (.BL(BL19),.BLN(BLN19),.WL(WL50));
sram_cell_6t_5 inst_cell_50_20 (.BL(BL20),.BLN(BLN20),.WL(WL50));
sram_cell_6t_5 inst_cell_50_21 (.BL(BL21),.BLN(BLN21),.WL(WL50));
sram_cell_6t_5 inst_cell_50_22 (.BL(BL22),.BLN(BLN22),.WL(WL50));
sram_cell_6t_5 inst_cell_50_23 (.BL(BL23),.BLN(BLN23),.WL(WL50));
sram_cell_6t_5 inst_cell_50_24 (.BL(BL24),.BLN(BLN24),.WL(WL50));
sram_cell_6t_5 inst_cell_50_25 (.BL(BL25),.BLN(BLN25),.WL(WL50));
sram_cell_6t_5 inst_cell_50_26 (.BL(BL26),.BLN(BLN26),.WL(WL50));
sram_cell_6t_5 inst_cell_50_27 (.BL(BL27),.BLN(BLN27),.WL(WL50));
sram_cell_6t_5 inst_cell_50_28 (.BL(BL28),.BLN(BLN28),.WL(WL50));
sram_cell_6t_5 inst_cell_50_29 (.BL(BL29),.BLN(BLN29),.WL(WL50));
sram_cell_6t_5 inst_cell_50_30 (.BL(BL30),.BLN(BLN30),.WL(WL50));
sram_cell_6t_5 inst_cell_50_31 (.BL(BL31),.BLN(BLN31),.WL(WL50));
sram_cell_6t_5 inst_cell_50_32 (.BL(BL32),.BLN(BLN32),.WL(WL50));
sram_cell_6t_5 inst_cell_50_33 (.BL(BL33),.BLN(BLN33),.WL(WL50));
sram_cell_6t_5 inst_cell_50_34 (.BL(BL34),.BLN(BLN34),.WL(WL50));
sram_cell_6t_5 inst_cell_50_35 (.BL(BL35),.BLN(BLN35),.WL(WL50));
sram_cell_6t_5 inst_cell_50_36 (.BL(BL36),.BLN(BLN36),.WL(WL50));
sram_cell_6t_5 inst_cell_50_37 (.BL(BL37),.BLN(BLN37),.WL(WL50));
sram_cell_6t_5 inst_cell_50_38 (.BL(BL38),.BLN(BLN38),.WL(WL50));
sram_cell_6t_5 inst_cell_50_39 (.BL(BL39),.BLN(BLN39),.WL(WL50));
sram_cell_6t_5 inst_cell_50_40 (.BL(BL40),.BLN(BLN40),.WL(WL50));
sram_cell_6t_5 inst_cell_50_41 (.BL(BL41),.BLN(BLN41),.WL(WL50));
sram_cell_6t_5 inst_cell_50_42 (.BL(BL42),.BLN(BLN42),.WL(WL50));
sram_cell_6t_5 inst_cell_50_43 (.BL(BL43),.BLN(BLN43),.WL(WL50));
sram_cell_6t_5 inst_cell_50_44 (.BL(BL44),.BLN(BLN44),.WL(WL50));
sram_cell_6t_5 inst_cell_50_45 (.BL(BL45),.BLN(BLN45),.WL(WL50));
sram_cell_6t_5 inst_cell_50_46 (.BL(BL46),.BLN(BLN46),.WL(WL50));
sram_cell_6t_5 inst_cell_50_47 (.BL(BL47),.BLN(BLN47),.WL(WL50));
sram_cell_6t_5 inst_cell_50_48 (.BL(BL48),.BLN(BLN48),.WL(WL50));
sram_cell_6t_5 inst_cell_50_49 (.BL(BL49),.BLN(BLN49),.WL(WL50));
sram_cell_6t_5 inst_cell_50_50 (.BL(BL50),.BLN(BLN50),.WL(WL50));
sram_cell_6t_5 inst_cell_50_51 (.BL(BL51),.BLN(BLN51),.WL(WL50));
sram_cell_6t_5 inst_cell_50_52 (.BL(BL52),.BLN(BLN52),.WL(WL50));
sram_cell_6t_5 inst_cell_50_53 (.BL(BL53),.BLN(BLN53),.WL(WL50));
sram_cell_6t_5 inst_cell_50_54 (.BL(BL54),.BLN(BLN54),.WL(WL50));
sram_cell_6t_5 inst_cell_50_55 (.BL(BL55),.BLN(BLN55),.WL(WL50));
sram_cell_6t_5 inst_cell_50_56 (.BL(BL56),.BLN(BLN56),.WL(WL50));
sram_cell_6t_5 inst_cell_50_57 (.BL(BL57),.BLN(BLN57),.WL(WL50));
sram_cell_6t_5 inst_cell_50_58 (.BL(BL58),.BLN(BLN58),.WL(WL50));
sram_cell_6t_5 inst_cell_50_59 (.BL(BL59),.BLN(BLN59),.WL(WL50));
sram_cell_6t_5 inst_cell_50_60 (.BL(BL60),.BLN(BLN60),.WL(WL50));
sram_cell_6t_5 inst_cell_50_61 (.BL(BL61),.BLN(BLN61),.WL(WL50));
sram_cell_6t_5 inst_cell_50_62 (.BL(BL62),.BLN(BLN62),.WL(WL50));
sram_cell_6t_5 inst_cell_50_63 (.BL(BL63),.BLN(BLN63),.WL(WL50));
sram_cell_6t_5 inst_cell_50_64 (.BL(BL64),.BLN(BLN64),.WL(WL50));
sram_cell_6t_5 inst_cell_50_65 (.BL(BL65),.BLN(BLN65),.WL(WL50));
sram_cell_6t_5 inst_cell_50_66 (.BL(BL66),.BLN(BLN66),.WL(WL50));
sram_cell_6t_5 inst_cell_50_67 (.BL(BL67),.BLN(BLN67),.WL(WL50));
sram_cell_6t_5 inst_cell_50_68 (.BL(BL68),.BLN(BLN68),.WL(WL50));
sram_cell_6t_5 inst_cell_50_69 (.BL(BL69),.BLN(BLN69),.WL(WL50));
sram_cell_6t_5 inst_cell_50_70 (.BL(BL70),.BLN(BLN70),.WL(WL50));
sram_cell_6t_5 inst_cell_50_71 (.BL(BL71),.BLN(BLN71),.WL(WL50));
sram_cell_6t_5 inst_cell_50_72 (.BL(BL72),.BLN(BLN72),.WL(WL50));
sram_cell_6t_5 inst_cell_50_73 (.BL(BL73),.BLN(BLN73),.WL(WL50));
sram_cell_6t_5 inst_cell_50_74 (.BL(BL74),.BLN(BLN74),.WL(WL50));
sram_cell_6t_5 inst_cell_50_75 (.BL(BL75),.BLN(BLN75),.WL(WL50));
sram_cell_6t_5 inst_cell_50_76 (.BL(BL76),.BLN(BLN76),.WL(WL50));
sram_cell_6t_5 inst_cell_50_77 (.BL(BL77),.BLN(BLN77),.WL(WL50));
sram_cell_6t_5 inst_cell_50_78 (.BL(BL78),.BLN(BLN78),.WL(WL50));
sram_cell_6t_5 inst_cell_50_79 (.BL(BL79),.BLN(BLN79),.WL(WL50));
sram_cell_6t_5 inst_cell_50_80 (.BL(BL80),.BLN(BLN80),.WL(WL50));
sram_cell_6t_5 inst_cell_50_81 (.BL(BL81),.BLN(BLN81),.WL(WL50));
sram_cell_6t_5 inst_cell_50_82 (.BL(BL82),.BLN(BLN82),.WL(WL50));
sram_cell_6t_5 inst_cell_50_83 (.BL(BL83),.BLN(BLN83),.WL(WL50));
sram_cell_6t_5 inst_cell_50_84 (.BL(BL84),.BLN(BLN84),.WL(WL50));
sram_cell_6t_5 inst_cell_50_85 (.BL(BL85),.BLN(BLN85),.WL(WL50));
sram_cell_6t_5 inst_cell_50_86 (.BL(BL86),.BLN(BLN86),.WL(WL50));
sram_cell_6t_5 inst_cell_50_87 (.BL(BL87),.BLN(BLN87),.WL(WL50));
sram_cell_6t_5 inst_cell_50_88 (.BL(BL88),.BLN(BLN88),.WL(WL50));
sram_cell_6t_5 inst_cell_50_89 (.BL(BL89),.BLN(BLN89),.WL(WL50));
sram_cell_6t_5 inst_cell_50_90 (.BL(BL90),.BLN(BLN90),.WL(WL50));
sram_cell_6t_5 inst_cell_50_91 (.BL(BL91),.BLN(BLN91),.WL(WL50));
sram_cell_6t_5 inst_cell_50_92 (.BL(BL92),.BLN(BLN92),.WL(WL50));
sram_cell_6t_5 inst_cell_50_93 (.BL(BL93),.BLN(BLN93),.WL(WL50));
sram_cell_6t_5 inst_cell_50_94 (.BL(BL94),.BLN(BLN94),.WL(WL50));
sram_cell_6t_5 inst_cell_50_95 (.BL(BL95),.BLN(BLN95),.WL(WL50));
sram_cell_6t_5 inst_cell_50_96 (.BL(BL96),.BLN(BLN96),.WL(WL50));
sram_cell_6t_5 inst_cell_50_97 (.BL(BL97),.BLN(BLN97),.WL(WL50));
sram_cell_6t_5 inst_cell_50_98 (.BL(BL98),.BLN(BLN98),.WL(WL50));
sram_cell_6t_5 inst_cell_50_99 (.BL(BL99),.BLN(BLN99),.WL(WL50));
sram_cell_6t_5 inst_cell_50_100 (.BL(BL100),.BLN(BLN100),.WL(WL50));
sram_cell_6t_5 inst_cell_50_101 (.BL(BL101),.BLN(BLN101),.WL(WL50));
sram_cell_6t_5 inst_cell_50_102 (.BL(BL102),.BLN(BLN102),.WL(WL50));
sram_cell_6t_5 inst_cell_50_103 (.BL(BL103),.BLN(BLN103),.WL(WL50));
sram_cell_6t_5 inst_cell_50_104 (.BL(BL104),.BLN(BLN104),.WL(WL50));
sram_cell_6t_5 inst_cell_50_105 (.BL(BL105),.BLN(BLN105),.WL(WL50));
sram_cell_6t_5 inst_cell_50_106 (.BL(BL106),.BLN(BLN106),.WL(WL50));
sram_cell_6t_5 inst_cell_50_107 (.BL(BL107),.BLN(BLN107),.WL(WL50));
sram_cell_6t_5 inst_cell_50_108 (.BL(BL108),.BLN(BLN108),.WL(WL50));
sram_cell_6t_5 inst_cell_50_109 (.BL(BL109),.BLN(BLN109),.WL(WL50));
sram_cell_6t_5 inst_cell_50_110 (.BL(BL110),.BLN(BLN110),.WL(WL50));
sram_cell_6t_5 inst_cell_50_111 (.BL(BL111),.BLN(BLN111),.WL(WL50));
sram_cell_6t_5 inst_cell_50_112 (.BL(BL112),.BLN(BLN112),.WL(WL50));
sram_cell_6t_5 inst_cell_50_113 (.BL(BL113),.BLN(BLN113),.WL(WL50));
sram_cell_6t_5 inst_cell_50_114 (.BL(BL114),.BLN(BLN114),.WL(WL50));
sram_cell_6t_5 inst_cell_50_115 (.BL(BL115),.BLN(BLN115),.WL(WL50));
sram_cell_6t_5 inst_cell_50_116 (.BL(BL116),.BLN(BLN116),.WL(WL50));
sram_cell_6t_5 inst_cell_50_117 (.BL(BL117),.BLN(BLN117),.WL(WL50));
sram_cell_6t_5 inst_cell_50_118 (.BL(BL118),.BLN(BLN118),.WL(WL50));
sram_cell_6t_5 inst_cell_50_119 (.BL(BL119),.BLN(BLN119),.WL(WL50));
sram_cell_6t_5 inst_cell_50_120 (.BL(BL120),.BLN(BLN120),.WL(WL50));
sram_cell_6t_5 inst_cell_50_121 (.BL(BL121),.BLN(BLN121),.WL(WL50));
sram_cell_6t_5 inst_cell_50_122 (.BL(BL122),.BLN(BLN122),.WL(WL50));
sram_cell_6t_5 inst_cell_50_123 (.BL(BL123),.BLN(BLN123),.WL(WL50));
sram_cell_6t_5 inst_cell_50_124 (.BL(BL124),.BLN(BLN124),.WL(WL50));
sram_cell_6t_5 inst_cell_50_125 (.BL(BL125),.BLN(BLN125),.WL(WL50));
sram_cell_6t_5 inst_cell_50_126 (.BL(BL126),.BLN(BLN126),.WL(WL50));
sram_cell_6t_5 inst_cell_50_127 (.BL(BL127),.BLN(BLN127),.WL(WL50));
sram_cell_6t_5 inst_cell_51_0 (.BL(BL0),.BLN(BLN0),.WL(WL51));
sram_cell_6t_5 inst_cell_51_1 (.BL(BL1),.BLN(BLN1),.WL(WL51));
sram_cell_6t_5 inst_cell_51_2 (.BL(BL2),.BLN(BLN2),.WL(WL51));
sram_cell_6t_5 inst_cell_51_3 (.BL(BL3),.BLN(BLN3),.WL(WL51));
sram_cell_6t_5 inst_cell_51_4 (.BL(BL4),.BLN(BLN4),.WL(WL51));
sram_cell_6t_5 inst_cell_51_5 (.BL(BL5),.BLN(BLN5),.WL(WL51));
sram_cell_6t_5 inst_cell_51_6 (.BL(BL6),.BLN(BLN6),.WL(WL51));
sram_cell_6t_5 inst_cell_51_7 (.BL(BL7),.BLN(BLN7),.WL(WL51));
sram_cell_6t_5 inst_cell_51_8 (.BL(BL8),.BLN(BLN8),.WL(WL51));
sram_cell_6t_5 inst_cell_51_9 (.BL(BL9),.BLN(BLN9),.WL(WL51));
sram_cell_6t_5 inst_cell_51_10 (.BL(BL10),.BLN(BLN10),.WL(WL51));
sram_cell_6t_5 inst_cell_51_11 (.BL(BL11),.BLN(BLN11),.WL(WL51));
sram_cell_6t_5 inst_cell_51_12 (.BL(BL12),.BLN(BLN12),.WL(WL51));
sram_cell_6t_5 inst_cell_51_13 (.BL(BL13),.BLN(BLN13),.WL(WL51));
sram_cell_6t_5 inst_cell_51_14 (.BL(BL14),.BLN(BLN14),.WL(WL51));
sram_cell_6t_5 inst_cell_51_15 (.BL(BL15),.BLN(BLN15),.WL(WL51));
sram_cell_6t_5 inst_cell_51_16 (.BL(BL16),.BLN(BLN16),.WL(WL51));
sram_cell_6t_5 inst_cell_51_17 (.BL(BL17),.BLN(BLN17),.WL(WL51));
sram_cell_6t_5 inst_cell_51_18 (.BL(BL18),.BLN(BLN18),.WL(WL51));
sram_cell_6t_5 inst_cell_51_19 (.BL(BL19),.BLN(BLN19),.WL(WL51));
sram_cell_6t_5 inst_cell_51_20 (.BL(BL20),.BLN(BLN20),.WL(WL51));
sram_cell_6t_5 inst_cell_51_21 (.BL(BL21),.BLN(BLN21),.WL(WL51));
sram_cell_6t_5 inst_cell_51_22 (.BL(BL22),.BLN(BLN22),.WL(WL51));
sram_cell_6t_5 inst_cell_51_23 (.BL(BL23),.BLN(BLN23),.WL(WL51));
sram_cell_6t_5 inst_cell_51_24 (.BL(BL24),.BLN(BLN24),.WL(WL51));
sram_cell_6t_5 inst_cell_51_25 (.BL(BL25),.BLN(BLN25),.WL(WL51));
sram_cell_6t_5 inst_cell_51_26 (.BL(BL26),.BLN(BLN26),.WL(WL51));
sram_cell_6t_5 inst_cell_51_27 (.BL(BL27),.BLN(BLN27),.WL(WL51));
sram_cell_6t_5 inst_cell_51_28 (.BL(BL28),.BLN(BLN28),.WL(WL51));
sram_cell_6t_5 inst_cell_51_29 (.BL(BL29),.BLN(BLN29),.WL(WL51));
sram_cell_6t_5 inst_cell_51_30 (.BL(BL30),.BLN(BLN30),.WL(WL51));
sram_cell_6t_5 inst_cell_51_31 (.BL(BL31),.BLN(BLN31),.WL(WL51));
sram_cell_6t_5 inst_cell_51_32 (.BL(BL32),.BLN(BLN32),.WL(WL51));
sram_cell_6t_5 inst_cell_51_33 (.BL(BL33),.BLN(BLN33),.WL(WL51));
sram_cell_6t_5 inst_cell_51_34 (.BL(BL34),.BLN(BLN34),.WL(WL51));
sram_cell_6t_5 inst_cell_51_35 (.BL(BL35),.BLN(BLN35),.WL(WL51));
sram_cell_6t_5 inst_cell_51_36 (.BL(BL36),.BLN(BLN36),.WL(WL51));
sram_cell_6t_5 inst_cell_51_37 (.BL(BL37),.BLN(BLN37),.WL(WL51));
sram_cell_6t_5 inst_cell_51_38 (.BL(BL38),.BLN(BLN38),.WL(WL51));
sram_cell_6t_5 inst_cell_51_39 (.BL(BL39),.BLN(BLN39),.WL(WL51));
sram_cell_6t_5 inst_cell_51_40 (.BL(BL40),.BLN(BLN40),.WL(WL51));
sram_cell_6t_5 inst_cell_51_41 (.BL(BL41),.BLN(BLN41),.WL(WL51));
sram_cell_6t_5 inst_cell_51_42 (.BL(BL42),.BLN(BLN42),.WL(WL51));
sram_cell_6t_5 inst_cell_51_43 (.BL(BL43),.BLN(BLN43),.WL(WL51));
sram_cell_6t_5 inst_cell_51_44 (.BL(BL44),.BLN(BLN44),.WL(WL51));
sram_cell_6t_5 inst_cell_51_45 (.BL(BL45),.BLN(BLN45),.WL(WL51));
sram_cell_6t_5 inst_cell_51_46 (.BL(BL46),.BLN(BLN46),.WL(WL51));
sram_cell_6t_5 inst_cell_51_47 (.BL(BL47),.BLN(BLN47),.WL(WL51));
sram_cell_6t_5 inst_cell_51_48 (.BL(BL48),.BLN(BLN48),.WL(WL51));
sram_cell_6t_5 inst_cell_51_49 (.BL(BL49),.BLN(BLN49),.WL(WL51));
sram_cell_6t_5 inst_cell_51_50 (.BL(BL50),.BLN(BLN50),.WL(WL51));
sram_cell_6t_5 inst_cell_51_51 (.BL(BL51),.BLN(BLN51),.WL(WL51));
sram_cell_6t_5 inst_cell_51_52 (.BL(BL52),.BLN(BLN52),.WL(WL51));
sram_cell_6t_5 inst_cell_51_53 (.BL(BL53),.BLN(BLN53),.WL(WL51));
sram_cell_6t_5 inst_cell_51_54 (.BL(BL54),.BLN(BLN54),.WL(WL51));
sram_cell_6t_5 inst_cell_51_55 (.BL(BL55),.BLN(BLN55),.WL(WL51));
sram_cell_6t_5 inst_cell_51_56 (.BL(BL56),.BLN(BLN56),.WL(WL51));
sram_cell_6t_5 inst_cell_51_57 (.BL(BL57),.BLN(BLN57),.WL(WL51));
sram_cell_6t_5 inst_cell_51_58 (.BL(BL58),.BLN(BLN58),.WL(WL51));
sram_cell_6t_5 inst_cell_51_59 (.BL(BL59),.BLN(BLN59),.WL(WL51));
sram_cell_6t_5 inst_cell_51_60 (.BL(BL60),.BLN(BLN60),.WL(WL51));
sram_cell_6t_5 inst_cell_51_61 (.BL(BL61),.BLN(BLN61),.WL(WL51));
sram_cell_6t_5 inst_cell_51_62 (.BL(BL62),.BLN(BLN62),.WL(WL51));
sram_cell_6t_5 inst_cell_51_63 (.BL(BL63),.BLN(BLN63),.WL(WL51));
sram_cell_6t_5 inst_cell_51_64 (.BL(BL64),.BLN(BLN64),.WL(WL51));
sram_cell_6t_5 inst_cell_51_65 (.BL(BL65),.BLN(BLN65),.WL(WL51));
sram_cell_6t_5 inst_cell_51_66 (.BL(BL66),.BLN(BLN66),.WL(WL51));
sram_cell_6t_5 inst_cell_51_67 (.BL(BL67),.BLN(BLN67),.WL(WL51));
sram_cell_6t_5 inst_cell_51_68 (.BL(BL68),.BLN(BLN68),.WL(WL51));
sram_cell_6t_5 inst_cell_51_69 (.BL(BL69),.BLN(BLN69),.WL(WL51));
sram_cell_6t_5 inst_cell_51_70 (.BL(BL70),.BLN(BLN70),.WL(WL51));
sram_cell_6t_5 inst_cell_51_71 (.BL(BL71),.BLN(BLN71),.WL(WL51));
sram_cell_6t_5 inst_cell_51_72 (.BL(BL72),.BLN(BLN72),.WL(WL51));
sram_cell_6t_5 inst_cell_51_73 (.BL(BL73),.BLN(BLN73),.WL(WL51));
sram_cell_6t_5 inst_cell_51_74 (.BL(BL74),.BLN(BLN74),.WL(WL51));
sram_cell_6t_5 inst_cell_51_75 (.BL(BL75),.BLN(BLN75),.WL(WL51));
sram_cell_6t_5 inst_cell_51_76 (.BL(BL76),.BLN(BLN76),.WL(WL51));
sram_cell_6t_5 inst_cell_51_77 (.BL(BL77),.BLN(BLN77),.WL(WL51));
sram_cell_6t_5 inst_cell_51_78 (.BL(BL78),.BLN(BLN78),.WL(WL51));
sram_cell_6t_5 inst_cell_51_79 (.BL(BL79),.BLN(BLN79),.WL(WL51));
sram_cell_6t_5 inst_cell_51_80 (.BL(BL80),.BLN(BLN80),.WL(WL51));
sram_cell_6t_5 inst_cell_51_81 (.BL(BL81),.BLN(BLN81),.WL(WL51));
sram_cell_6t_5 inst_cell_51_82 (.BL(BL82),.BLN(BLN82),.WL(WL51));
sram_cell_6t_5 inst_cell_51_83 (.BL(BL83),.BLN(BLN83),.WL(WL51));
sram_cell_6t_5 inst_cell_51_84 (.BL(BL84),.BLN(BLN84),.WL(WL51));
sram_cell_6t_5 inst_cell_51_85 (.BL(BL85),.BLN(BLN85),.WL(WL51));
sram_cell_6t_5 inst_cell_51_86 (.BL(BL86),.BLN(BLN86),.WL(WL51));
sram_cell_6t_5 inst_cell_51_87 (.BL(BL87),.BLN(BLN87),.WL(WL51));
sram_cell_6t_5 inst_cell_51_88 (.BL(BL88),.BLN(BLN88),.WL(WL51));
sram_cell_6t_5 inst_cell_51_89 (.BL(BL89),.BLN(BLN89),.WL(WL51));
sram_cell_6t_5 inst_cell_51_90 (.BL(BL90),.BLN(BLN90),.WL(WL51));
sram_cell_6t_5 inst_cell_51_91 (.BL(BL91),.BLN(BLN91),.WL(WL51));
sram_cell_6t_5 inst_cell_51_92 (.BL(BL92),.BLN(BLN92),.WL(WL51));
sram_cell_6t_5 inst_cell_51_93 (.BL(BL93),.BLN(BLN93),.WL(WL51));
sram_cell_6t_5 inst_cell_51_94 (.BL(BL94),.BLN(BLN94),.WL(WL51));
sram_cell_6t_5 inst_cell_51_95 (.BL(BL95),.BLN(BLN95),.WL(WL51));
sram_cell_6t_5 inst_cell_51_96 (.BL(BL96),.BLN(BLN96),.WL(WL51));
sram_cell_6t_5 inst_cell_51_97 (.BL(BL97),.BLN(BLN97),.WL(WL51));
sram_cell_6t_5 inst_cell_51_98 (.BL(BL98),.BLN(BLN98),.WL(WL51));
sram_cell_6t_5 inst_cell_51_99 (.BL(BL99),.BLN(BLN99),.WL(WL51));
sram_cell_6t_5 inst_cell_51_100 (.BL(BL100),.BLN(BLN100),.WL(WL51));
sram_cell_6t_5 inst_cell_51_101 (.BL(BL101),.BLN(BLN101),.WL(WL51));
sram_cell_6t_5 inst_cell_51_102 (.BL(BL102),.BLN(BLN102),.WL(WL51));
sram_cell_6t_5 inst_cell_51_103 (.BL(BL103),.BLN(BLN103),.WL(WL51));
sram_cell_6t_5 inst_cell_51_104 (.BL(BL104),.BLN(BLN104),.WL(WL51));
sram_cell_6t_5 inst_cell_51_105 (.BL(BL105),.BLN(BLN105),.WL(WL51));
sram_cell_6t_5 inst_cell_51_106 (.BL(BL106),.BLN(BLN106),.WL(WL51));
sram_cell_6t_5 inst_cell_51_107 (.BL(BL107),.BLN(BLN107),.WL(WL51));
sram_cell_6t_5 inst_cell_51_108 (.BL(BL108),.BLN(BLN108),.WL(WL51));
sram_cell_6t_5 inst_cell_51_109 (.BL(BL109),.BLN(BLN109),.WL(WL51));
sram_cell_6t_5 inst_cell_51_110 (.BL(BL110),.BLN(BLN110),.WL(WL51));
sram_cell_6t_5 inst_cell_51_111 (.BL(BL111),.BLN(BLN111),.WL(WL51));
sram_cell_6t_5 inst_cell_51_112 (.BL(BL112),.BLN(BLN112),.WL(WL51));
sram_cell_6t_5 inst_cell_51_113 (.BL(BL113),.BLN(BLN113),.WL(WL51));
sram_cell_6t_5 inst_cell_51_114 (.BL(BL114),.BLN(BLN114),.WL(WL51));
sram_cell_6t_5 inst_cell_51_115 (.BL(BL115),.BLN(BLN115),.WL(WL51));
sram_cell_6t_5 inst_cell_51_116 (.BL(BL116),.BLN(BLN116),.WL(WL51));
sram_cell_6t_5 inst_cell_51_117 (.BL(BL117),.BLN(BLN117),.WL(WL51));
sram_cell_6t_5 inst_cell_51_118 (.BL(BL118),.BLN(BLN118),.WL(WL51));
sram_cell_6t_5 inst_cell_51_119 (.BL(BL119),.BLN(BLN119),.WL(WL51));
sram_cell_6t_5 inst_cell_51_120 (.BL(BL120),.BLN(BLN120),.WL(WL51));
sram_cell_6t_5 inst_cell_51_121 (.BL(BL121),.BLN(BLN121),.WL(WL51));
sram_cell_6t_5 inst_cell_51_122 (.BL(BL122),.BLN(BLN122),.WL(WL51));
sram_cell_6t_5 inst_cell_51_123 (.BL(BL123),.BLN(BLN123),.WL(WL51));
sram_cell_6t_5 inst_cell_51_124 (.BL(BL124),.BLN(BLN124),.WL(WL51));
sram_cell_6t_5 inst_cell_51_125 (.BL(BL125),.BLN(BLN125),.WL(WL51));
sram_cell_6t_5 inst_cell_51_126 (.BL(BL126),.BLN(BLN126),.WL(WL51));
sram_cell_6t_5 inst_cell_51_127 (.BL(BL127),.BLN(BLN127),.WL(WL51));
sram_cell_6t_5 inst_cell_52_0 (.BL(BL0),.BLN(BLN0),.WL(WL52));
sram_cell_6t_5 inst_cell_52_1 (.BL(BL1),.BLN(BLN1),.WL(WL52));
sram_cell_6t_5 inst_cell_52_2 (.BL(BL2),.BLN(BLN2),.WL(WL52));
sram_cell_6t_5 inst_cell_52_3 (.BL(BL3),.BLN(BLN3),.WL(WL52));
sram_cell_6t_5 inst_cell_52_4 (.BL(BL4),.BLN(BLN4),.WL(WL52));
sram_cell_6t_5 inst_cell_52_5 (.BL(BL5),.BLN(BLN5),.WL(WL52));
sram_cell_6t_5 inst_cell_52_6 (.BL(BL6),.BLN(BLN6),.WL(WL52));
sram_cell_6t_5 inst_cell_52_7 (.BL(BL7),.BLN(BLN7),.WL(WL52));
sram_cell_6t_5 inst_cell_52_8 (.BL(BL8),.BLN(BLN8),.WL(WL52));
sram_cell_6t_5 inst_cell_52_9 (.BL(BL9),.BLN(BLN9),.WL(WL52));
sram_cell_6t_5 inst_cell_52_10 (.BL(BL10),.BLN(BLN10),.WL(WL52));
sram_cell_6t_5 inst_cell_52_11 (.BL(BL11),.BLN(BLN11),.WL(WL52));
sram_cell_6t_5 inst_cell_52_12 (.BL(BL12),.BLN(BLN12),.WL(WL52));
sram_cell_6t_5 inst_cell_52_13 (.BL(BL13),.BLN(BLN13),.WL(WL52));
sram_cell_6t_5 inst_cell_52_14 (.BL(BL14),.BLN(BLN14),.WL(WL52));
sram_cell_6t_5 inst_cell_52_15 (.BL(BL15),.BLN(BLN15),.WL(WL52));
sram_cell_6t_5 inst_cell_52_16 (.BL(BL16),.BLN(BLN16),.WL(WL52));
sram_cell_6t_5 inst_cell_52_17 (.BL(BL17),.BLN(BLN17),.WL(WL52));
sram_cell_6t_5 inst_cell_52_18 (.BL(BL18),.BLN(BLN18),.WL(WL52));
sram_cell_6t_5 inst_cell_52_19 (.BL(BL19),.BLN(BLN19),.WL(WL52));
sram_cell_6t_5 inst_cell_52_20 (.BL(BL20),.BLN(BLN20),.WL(WL52));
sram_cell_6t_5 inst_cell_52_21 (.BL(BL21),.BLN(BLN21),.WL(WL52));
sram_cell_6t_5 inst_cell_52_22 (.BL(BL22),.BLN(BLN22),.WL(WL52));
sram_cell_6t_5 inst_cell_52_23 (.BL(BL23),.BLN(BLN23),.WL(WL52));
sram_cell_6t_5 inst_cell_52_24 (.BL(BL24),.BLN(BLN24),.WL(WL52));
sram_cell_6t_5 inst_cell_52_25 (.BL(BL25),.BLN(BLN25),.WL(WL52));
sram_cell_6t_5 inst_cell_52_26 (.BL(BL26),.BLN(BLN26),.WL(WL52));
sram_cell_6t_5 inst_cell_52_27 (.BL(BL27),.BLN(BLN27),.WL(WL52));
sram_cell_6t_5 inst_cell_52_28 (.BL(BL28),.BLN(BLN28),.WL(WL52));
sram_cell_6t_5 inst_cell_52_29 (.BL(BL29),.BLN(BLN29),.WL(WL52));
sram_cell_6t_5 inst_cell_52_30 (.BL(BL30),.BLN(BLN30),.WL(WL52));
sram_cell_6t_5 inst_cell_52_31 (.BL(BL31),.BLN(BLN31),.WL(WL52));
sram_cell_6t_5 inst_cell_52_32 (.BL(BL32),.BLN(BLN32),.WL(WL52));
sram_cell_6t_5 inst_cell_52_33 (.BL(BL33),.BLN(BLN33),.WL(WL52));
sram_cell_6t_5 inst_cell_52_34 (.BL(BL34),.BLN(BLN34),.WL(WL52));
sram_cell_6t_5 inst_cell_52_35 (.BL(BL35),.BLN(BLN35),.WL(WL52));
sram_cell_6t_5 inst_cell_52_36 (.BL(BL36),.BLN(BLN36),.WL(WL52));
sram_cell_6t_5 inst_cell_52_37 (.BL(BL37),.BLN(BLN37),.WL(WL52));
sram_cell_6t_5 inst_cell_52_38 (.BL(BL38),.BLN(BLN38),.WL(WL52));
sram_cell_6t_5 inst_cell_52_39 (.BL(BL39),.BLN(BLN39),.WL(WL52));
sram_cell_6t_5 inst_cell_52_40 (.BL(BL40),.BLN(BLN40),.WL(WL52));
sram_cell_6t_5 inst_cell_52_41 (.BL(BL41),.BLN(BLN41),.WL(WL52));
sram_cell_6t_5 inst_cell_52_42 (.BL(BL42),.BLN(BLN42),.WL(WL52));
sram_cell_6t_5 inst_cell_52_43 (.BL(BL43),.BLN(BLN43),.WL(WL52));
sram_cell_6t_5 inst_cell_52_44 (.BL(BL44),.BLN(BLN44),.WL(WL52));
sram_cell_6t_5 inst_cell_52_45 (.BL(BL45),.BLN(BLN45),.WL(WL52));
sram_cell_6t_5 inst_cell_52_46 (.BL(BL46),.BLN(BLN46),.WL(WL52));
sram_cell_6t_5 inst_cell_52_47 (.BL(BL47),.BLN(BLN47),.WL(WL52));
sram_cell_6t_5 inst_cell_52_48 (.BL(BL48),.BLN(BLN48),.WL(WL52));
sram_cell_6t_5 inst_cell_52_49 (.BL(BL49),.BLN(BLN49),.WL(WL52));
sram_cell_6t_5 inst_cell_52_50 (.BL(BL50),.BLN(BLN50),.WL(WL52));
sram_cell_6t_5 inst_cell_52_51 (.BL(BL51),.BLN(BLN51),.WL(WL52));
sram_cell_6t_5 inst_cell_52_52 (.BL(BL52),.BLN(BLN52),.WL(WL52));
sram_cell_6t_5 inst_cell_52_53 (.BL(BL53),.BLN(BLN53),.WL(WL52));
sram_cell_6t_5 inst_cell_52_54 (.BL(BL54),.BLN(BLN54),.WL(WL52));
sram_cell_6t_5 inst_cell_52_55 (.BL(BL55),.BLN(BLN55),.WL(WL52));
sram_cell_6t_5 inst_cell_52_56 (.BL(BL56),.BLN(BLN56),.WL(WL52));
sram_cell_6t_5 inst_cell_52_57 (.BL(BL57),.BLN(BLN57),.WL(WL52));
sram_cell_6t_5 inst_cell_52_58 (.BL(BL58),.BLN(BLN58),.WL(WL52));
sram_cell_6t_5 inst_cell_52_59 (.BL(BL59),.BLN(BLN59),.WL(WL52));
sram_cell_6t_5 inst_cell_52_60 (.BL(BL60),.BLN(BLN60),.WL(WL52));
sram_cell_6t_5 inst_cell_52_61 (.BL(BL61),.BLN(BLN61),.WL(WL52));
sram_cell_6t_5 inst_cell_52_62 (.BL(BL62),.BLN(BLN62),.WL(WL52));
sram_cell_6t_5 inst_cell_52_63 (.BL(BL63),.BLN(BLN63),.WL(WL52));
sram_cell_6t_5 inst_cell_52_64 (.BL(BL64),.BLN(BLN64),.WL(WL52));
sram_cell_6t_5 inst_cell_52_65 (.BL(BL65),.BLN(BLN65),.WL(WL52));
sram_cell_6t_5 inst_cell_52_66 (.BL(BL66),.BLN(BLN66),.WL(WL52));
sram_cell_6t_5 inst_cell_52_67 (.BL(BL67),.BLN(BLN67),.WL(WL52));
sram_cell_6t_5 inst_cell_52_68 (.BL(BL68),.BLN(BLN68),.WL(WL52));
sram_cell_6t_5 inst_cell_52_69 (.BL(BL69),.BLN(BLN69),.WL(WL52));
sram_cell_6t_5 inst_cell_52_70 (.BL(BL70),.BLN(BLN70),.WL(WL52));
sram_cell_6t_5 inst_cell_52_71 (.BL(BL71),.BLN(BLN71),.WL(WL52));
sram_cell_6t_5 inst_cell_52_72 (.BL(BL72),.BLN(BLN72),.WL(WL52));
sram_cell_6t_5 inst_cell_52_73 (.BL(BL73),.BLN(BLN73),.WL(WL52));
sram_cell_6t_5 inst_cell_52_74 (.BL(BL74),.BLN(BLN74),.WL(WL52));
sram_cell_6t_5 inst_cell_52_75 (.BL(BL75),.BLN(BLN75),.WL(WL52));
sram_cell_6t_5 inst_cell_52_76 (.BL(BL76),.BLN(BLN76),.WL(WL52));
sram_cell_6t_5 inst_cell_52_77 (.BL(BL77),.BLN(BLN77),.WL(WL52));
sram_cell_6t_5 inst_cell_52_78 (.BL(BL78),.BLN(BLN78),.WL(WL52));
sram_cell_6t_5 inst_cell_52_79 (.BL(BL79),.BLN(BLN79),.WL(WL52));
sram_cell_6t_5 inst_cell_52_80 (.BL(BL80),.BLN(BLN80),.WL(WL52));
sram_cell_6t_5 inst_cell_52_81 (.BL(BL81),.BLN(BLN81),.WL(WL52));
sram_cell_6t_5 inst_cell_52_82 (.BL(BL82),.BLN(BLN82),.WL(WL52));
sram_cell_6t_5 inst_cell_52_83 (.BL(BL83),.BLN(BLN83),.WL(WL52));
sram_cell_6t_5 inst_cell_52_84 (.BL(BL84),.BLN(BLN84),.WL(WL52));
sram_cell_6t_5 inst_cell_52_85 (.BL(BL85),.BLN(BLN85),.WL(WL52));
sram_cell_6t_5 inst_cell_52_86 (.BL(BL86),.BLN(BLN86),.WL(WL52));
sram_cell_6t_5 inst_cell_52_87 (.BL(BL87),.BLN(BLN87),.WL(WL52));
sram_cell_6t_5 inst_cell_52_88 (.BL(BL88),.BLN(BLN88),.WL(WL52));
sram_cell_6t_5 inst_cell_52_89 (.BL(BL89),.BLN(BLN89),.WL(WL52));
sram_cell_6t_5 inst_cell_52_90 (.BL(BL90),.BLN(BLN90),.WL(WL52));
sram_cell_6t_5 inst_cell_52_91 (.BL(BL91),.BLN(BLN91),.WL(WL52));
sram_cell_6t_5 inst_cell_52_92 (.BL(BL92),.BLN(BLN92),.WL(WL52));
sram_cell_6t_5 inst_cell_52_93 (.BL(BL93),.BLN(BLN93),.WL(WL52));
sram_cell_6t_5 inst_cell_52_94 (.BL(BL94),.BLN(BLN94),.WL(WL52));
sram_cell_6t_5 inst_cell_52_95 (.BL(BL95),.BLN(BLN95),.WL(WL52));
sram_cell_6t_5 inst_cell_52_96 (.BL(BL96),.BLN(BLN96),.WL(WL52));
sram_cell_6t_5 inst_cell_52_97 (.BL(BL97),.BLN(BLN97),.WL(WL52));
sram_cell_6t_5 inst_cell_52_98 (.BL(BL98),.BLN(BLN98),.WL(WL52));
sram_cell_6t_5 inst_cell_52_99 (.BL(BL99),.BLN(BLN99),.WL(WL52));
sram_cell_6t_5 inst_cell_52_100 (.BL(BL100),.BLN(BLN100),.WL(WL52));
sram_cell_6t_5 inst_cell_52_101 (.BL(BL101),.BLN(BLN101),.WL(WL52));
sram_cell_6t_5 inst_cell_52_102 (.BL(BL102),.BLN(BLN102),.WL(WL52));
sram_cell_6t_5 inst_cell_52_103 (.BL(BL103),.BLN(BLN103),.WL(WL52));
sram_cell_6t_5 inst_cell_52_104 (.BL(BL104),.BLN(BLN104),.WL(WL52));
sram_cell_6t_5 inst_cell_52_105 (.BL(BL105),.BLN(BLN105),.WL(WL52));
sram_cell_6t_5 inst_cell_52_106 (.BL(BL106),.BLN(BLN106),.WL(WL52));
sram_cell_6t_5 inst_cell_52_107 (.BL(BL107),.BLN(BLN107),.WL(WL52));
sram_cell_6t_5 inst_cell_52_108 (.BL(BL108),.BLN(BLN108),.WL(WL52));
sram_cell_6t_5 inst_cell_52_109 (.BL(BL109),.BLN(BLN109),.WL(WL52));
sram_cell_6t_5 inst_cell_52_110 (.BL(BL110),.BLN(BLN110),.WL(WL52));
sram_cell_6t_5 inst_cell_52_111 (.BL(BL111),.BLN(BLN111),.WL(WL52));
sram_cell_6t_5 inst_cell_52_112 (.BL(BL112),.BLN(BLN112),.WL(WL52));
sram_cell_6t_5 inst_cell_52_113 (.BL(BL113),.BLN(BLN113),.WL(WL52));
sram_cell_6t_5 inst_cell_52_114 (.BL(BL114),.BLN(BLN114),.WL(WL52));
sram_cell_6t_5 inst_cell_52_115 (.BL(BL115),.BLN(BLN115),.WL(WL52));
sram_cell_6t_5 inst_cell_52_116 (.BL(BL116),.BLN(BLN116),.WL(WL52));
sram_cell_6t_5 inst_cell_52_117 (.BL(BL117),.BLN(BLN117),.WL(WL52));
sram_cell_6t_5 inst_cell_52_118 (.BL(BL118),.BLN(BLN118),.WL(WL52));
sram_cell_6t_5 inst_cell_52_119 (.BL(BL119),.BLN(BLN119),.WL(WL52));
sram_cell_6t_5 inst_cell_52_120 (.BL(BL120),.BLN(BLN120),.WL(WL52));
sram_cell_6t_5 inst_cell_52_121 (.BL(BL121),.BLN(BLN121),.WL(WL52));
sram_cell_6t_5 inst_cell_52_122 (.BL(BL122),.BLN(BLN122),.WL(WL52));
sram_cell_6t_5 inst_cell_52_123 (.BL(BL123),.BLN(BLN123),.WL(WL52));
sram_cell_6t_5 inst_cell_52_124 (.BL(BL124),.BLN(BLN124),.WL(WL52));
sram_cell_6t_5 inst_cell_52_125 (.BL(BL125),.BLN(BLN125),.WL(WL52));
sram_cell_6t_5 inst_cell_52_126 (.BL(BL126),.BLN(BLN126),.WL(WL52));
sram_cell_6t_5 inst_cell_52_127 (.BL(BL127),.BLN(BLN127),.WL(WL52));
sram_cell_6t_5 inst_cell_53_0 (.BL(BL0),.BLN(BLN0),.WL(WL53));
sram_cell_6t_5 inst_cell_53_1 (.BL(BL1),.BLN(BLN1),.WL(WL53));
sram_cell_6t_5 inst_cell_53_2 (.BL(BL2),.BLN(BLN2),.WL(WL53));
sram_cell_6t_5 inst_cell_53_3 (.BL(BL3),.BLN(BLN3),.WL(WL53));
sram_cell_6t_5 inst_cell_53_4 (.BL(BL4),.BLN(BLN4),.WL(WL53));
sram_cell_6t_5 inst_cell_53_5 (.BL(BL5),.BLN(BLN5),.WL(WL53));
sram_cell_6t_5 inst_cell_53_6 (.BL(BL6),.BLN(BLN6),.WL(WL53));
sram_cell_6t_5 inst_cell_53_7 (.BL(BL7),.BLN(BLN7),.WL(WL53));
sram_cell_6t_5 inst_cell_53_8 (.BL(BL8),.BLN(BLN8),.WL(WL53));
sram_cell_6t_5 inst_cell_53_9 (.BL(BL9),.BLN(BLN9),.WL(WL53));
sram_cell_6t_5 inst_cell_53_10 (.BL(BL10),.BLN(BLN10),.WL(WL53));
sram_cell_6t_5 inst_cell_53_11 (.BL(BL11),.BLN(BLN11),.WL(WL53));
sram_cell_6t_5 inst_cell_53_12 (.BL(BL12),.BLN(BLN12),.WL(WL53));
sram_cell_6t_5 inst_cell_53_13 (.BL(BL13),.BLN(BLN13),.WL(WL53));
sram_cell_6t_5 inst_cell_53_14 (.BL(BL14),.BLN(BLN14),.WL(WL53));
sram_cell_6t_5 inst_cell_53_15 (.BL(BL15),.BLN(BLN15),.WL(WL53));
sram_cell_6t_5 inst_cell_53_16 (.BL(BL16),.BLN(BLN16),.WL(WL53));
sram_cell_6t_5 inst_cell_53_17 (.BL(BL17),.BLN(BLN17),.WL(WL53));
sram_cell_6t_5 inst_cell_53_18 (.BL(BL18),.BLN(BLN18),.WL(WL53));
sram_cell_6t_5 inst_cell_53_19 (.BL(BL19),.BLN(BLN19),.WL(WL53));
sram_cell_6t_5 inst_cell_53_20 (.BL(BL20),.BLN(BLN20),.WL(WL53));
sram_cell_6t_5 inst_cell_53_21 (.BL(BL21),.BLN(BLN21),.WL(WL53));
sram_cell_6t_5 inst_cell_53_22 (.BL(BL22),.BLN(BLN22),.WL(WL53));
sram_cell_6t_5 inst_cell_53_23 (.BL(BL23),.BLN(BLN23),.WL(WL53));
sram_cell_6t_5 inst_cell_53_24 (.BL(BL24),.BLN(BLN24),.WL(WL53));
sram_cell_6t_5 inst_cell_53_25 (.BL(BL25),.BLN(BLN25),.WL(WL53));
sram_cell_6t_5 inst_cell_53_26 (.BL(BL26),.BLN(BLN26),.WL(WL53));
sram_cell_6t_5 inst_cell_53_27 (.BL(BL27),.BLN(BLN27),.WL(WL53));
sram_cell_6t_5 inst_cell_53_28 (.BL(BL28),.BLN(BLN28),.WL(WL53));
sram_cell_6t_5 inst_cell_53_29 (.BL(BL29),.BLN(BLN29),.WL(WL53));
sram_cell_6t_5 inst_cell_53_30 (.BL(BL30),.BLN(BLN30),.WL(WL53));
sram_cell_6t_5 inst_cell_53_31 (.BL(BL31),.BLN(BLN31),.WL(WL53));
sram_cell_6t_5 inst_cell_53_32 (.BL(BL32),.BLN(BLN32),.WL(WL53));
sram_cell_6t_5 inst_cell_53_33 (.BL(BL33),.BLN(BLN33),.WL(WL53));
sram_cell_6t_5 inst_cell_53_34 (.BL(BL34),.BLN(BLN34),.WL(WL53));
sram_cell_6t_5 inst_cell_53_35 (.BL(BL35),.BLN(BLN35),.WL(WL53));
sram_cell_6t_5 inst_cell_53_36 (.BL(BL36),.BLN(BLN36),.WL(WL53));
sram_cell_6t_5 inst_cell_53_37 (.BL(BL37),.BLN(BLN37),.WL(WL53));
sram_cell_6t_5 inst_cell_53_38 (.BL(BL38),.BLN(BLN38),.WL(WL53));
sram_cell_6t_5 inst_cell_53_39 (.BL(BL39),.BLN(BLN39),.WL(WL53));
sram_cell_6t_5 inst_cell_53_40 (.BL(BL40),.BLN(BLN40),.WL(WL53));
sram_cell_6t_5 inst_cell_53_41 (.BL(BL41),.BLN(BLN41),.WL(WL53));
sram_cell_6t_5 inst_cell_53_42 (.BL(BL42),.BLN(BLN42),.WL(WL53));
sram_cell_6t_5 inst_cell_53_43 (.BL(BL43),.BLN(BLN43),.WL(WL53));
sram_cell_6t_5 inst_cell_53_44 (.BL(BL44),.BLN(BLN44),.WL(WL53));
sram_cell_6t_5 inst_cell_53_45 (.BL(BL45),.BLN(BLN45),.WL(WL53));
sram_cell_6t_5 inst_cell_53_46 (.BL(BL46),.BLN(BLN46),.WL(WL53));
sram_cell_6t_5 inst_cell_53_47 (.BL(BL47),.BLN(BLN47),.WL(WL53));
sram_cell_6t_5 inst_cell_53_48 (.BL(BL48),.BLN(BLN48),.WL(WL53));
sram_cell_6t_5 inst_cell_53_49 (.BL(BL49),.BLN(BLN49),.WL(WL53));
sram_cell_6t_5 inst_cell_53_50 (.BL(BL50),.BLN(BLN50),.WL(WL53));
sram_cell_6t_5 inst_cell_53_51 (.BL(BL51),.BLN(BLN51),.WL(WL53));
sram_cell_6t_5 inst_cell_53_52 (.BL(BL52),.BLN(BLN52),.WL(WL53));
sram_cell_6t_5 inst_cell_53_53 (.BL(BL53),.BLN(BLN53),.WL(WL53));
sram_cell_6t_5 inst_cell_53_54 (.BL(BL54),.BLN(BLN54),.WL(WL53));
sram_cell_6t_5 inst_cell_53_55 (.BL(BL55),.BLN(BLN55),.WL(WL53));
sram_cell_6t_5 inst_cell_53_56 (.BL(BL56),.BLN(BLN56),.WL(WL53));
sram_cell_6t_5 inst_cell_53_57 (.BL(BL57),.BLN(BLN57),.WL(WL53));
sram_cell_6t_5 inst_cell_53_58 (.BL(BL58),.BLN(BLN58),.WL(WL53));
sram_cell_6t_5 inst_cell_53_59 (.BL(BL59),.BLN(BLN59),.WL(WL53));
sram_cell_6t_5 inst_cell_53_60 (.BL(BL60),.BLN(BLN60),.WL(WL53));
sram_cell_6t_5 inst_cell_53_61 (.BL(BL61),.BLN(BLN61),.WL(WL53));
sram_cell_6t_5 inst_cell_53_62 (.BL(BL62),.BLN(BLN62),.WL(WL53));
sram_cell_6t_5 inst_cell_53_63 (.BL(BL63),.BLN(BLN63),.WL(WL53));
sram_cell_6t_5 inst_cell_53_64 (.BL(BL64),.BLN(BLN64),.WL(WL53));
sram_cell_6t_5 inst_cell_53_65 (.BL(BL65),.BLN(BLN65),.WL(WL53));
sram_cell_6t_5 inst_cell_53_66 (.BL(BL66),.BLN(BLN66),.WL(WL53));
sram_cell_6t_5 inst_cell_53_67 (.BL(BL67),.BLN(BLN67),.WL(WL53));
sram_cell_6t_5 inst_cell_53_68 (.BL(BL68),.BLN(BLN68),.WL(WL53));
sram_cell_6t_5 inst_cell_53_69 (.BL(BL69),.BLN(BLN69),.WL(WL53));
sram_cell_6t_5 inst_cell_53_70 (.BL(BL70),.BLN(BLN70),.WL(WL53));
sram_cell_6t_5 inst_cell_53_71 (.BL(BL71),.BLN(BLN71),.WL(WL53));
sram_cell_6t_5 inst_cell_53_72 (.BL(BL72),.BLN(BLN72),.WL(WL53));
sram_cell_6t_5 inst_cell_53_73 (.BL(BL73),.BLN(BLN73),.WL(WL53));
sram_cell_6t_5 inst_cell_53_74 (.BL(BL74),.BLN(BLN74),.WL(WL53));
sram_cell_6t_5 inst_cell_53_75 (.BL(BL75),.BLN(BLN75),.WL(WL53));
sram_cell_6t_5 inst_cell_53_76 (.BL(BL76),.BLN(BLN76),.WL(WL53));
sram_cell_6t_5 inst_cell_53_77 (.BL(BL77),.BLN(BLN77),.WL(WL53));
sram_cell_6t_5 inst_cell_53_78 (.BL(BL78),.BLN(BLN78),.WL(WL53));
sram_cell_6t_5 inst_cell_53_79 (.BL(BL79),.BLN(BLN79),.WL(WL53));
sram_cell_6t_5 inst_cell_53_80 (.BL(BL80),.BLN(BLN80),.WL(WL53));
sram_cell_6t_5 inst_cell_53_81 (.BL(BL81),.BLN(BLN81),.WL(WL53));
sram_cell_6t_5 inst_cell_53_82 (.BL(BL82),.BLN(BLN82),.WL(WL53));
sram_cell_6t_5 inst_cell_53_83 (.BL(BL83),.BLN(BLN83),.WL(WL53));
sram_cell_6t_5 inst_cell_53_84 (.BL(BL84),.BLN(BLN84),.WL(WL53));
sram_cell_6t_5 inst_cell_53_85 (.BL(BL85),.BLN(BLN85),.WL(WL53));
sram_cell_6t_5 inst_cell_53_86 (.BL(BL86),.BLN(BLN86),.WL(WL53));
sram_cell_6t_5 inst_cell_53_87 (.BL(BL87),.BLN(BLN87),.WL(WL53));
sram_cell_6t_5 inst_cell_53_88 (.BL(BL88),.BLN(BLN88),.WL(WL53));
sram_cell_6t_5 inst_cell_53_89 (.BL(BL89),.BLN(BLN89),.WL(WL53));
sram_cell_6t_5 inst_cell_53_90 (.BL(BL90),.BLN(BLN90),.WL(WL53));
sram_cell_6t_5 inst_cell_53_91 (.BL(BL91),.BLN(BLN91),.WL(WL53));
sram_cell_6t_5 inst_cell_53_92 (.BL(BL92),.BLN(BLN92),.WL(WL53));
sram_cell_6t_5 inst_cell_53_93 (.BL(BL93),.BLN(BLN93),.WL(WL53));
sram_cell_6t_5 inst_cell_53_94 (.BL(BL94),.BLN(BLN94),.WL(WL53));
sram_cell_6t_5 inst_cell_53_95 (.BL(BL95),.BLN(BLN95),.WL(WL53));
sram_cell_6t_5 inst_cell_53_96 (.BL(BL96),.BLN(BLN96),.WL(WL53));
sram_cell_6t_5 inst_cell_53_97 (.BL(BL97),.BLN(BLN97),.WL(WL53));
sram_cell_6t_5 inst_cell_53_98 (.BL(BL98),.BLN(BLN98),.WL(WL53));
sram_cell_6t_5 inst_cell_53_99 (.BL(BL99),.BLN(BLN99),.WL(WL53));
sram_cell_6t_5 inst_cell_53_100 (.BL(BL100),.BLN(BLN100),.WL(WL53));
sram_cell_6t_5 inst_cell_53_101 (.BL(BL101),.BLN(BLN101),.WL(WL53));
sram_cell_6t_5 inst_cell_53_102 (.BL(BL102),.BLN(BLN102),.WL(WL53));
sram_cell_6t_5 inst_cell_53_103 (.BL(BL103),.BLN(BLN103),.WL(WL53));
sram_cell_6t_5 inst_cell_53_104 (.BL(BL104),.BLN(BLN104),.WL(WL53));
sram_cell_6t_5 inst_cell_53_105 (.BL(BL105),.BLN(BLN105),.WL(WL53));
sram_cell_6t_5 inst_cell_53_106 (.BL(BL106),.BLN(BLN106),.WL(WL53));
sram_cell_6t_5 inst_cell_53_107 (.BL(BL107),.BLN(BLN107),.WL(WL53));
sram_cell_6t_5 inst_cell_53_108 (.BL(BL108),.BLN(BLN108),.WL(WL53));
sram_cell_6t_5 inst_cell_53_109 (.BL(BL109),.BLN(BLN109),.WL(WL53));
sram_cell_6t_5 inst_cell_53_110 (.BL(BL110),.BLN(BLN110),.WL(WL53));
sram_cell_6t_5 inst_cell_53_111 (.BL(BL111),.BLN(BLN111),.WL(WL53));
sram_cell_6t_5 inst_cell_53_112 (.BL(BL112),.BLN(BLN112),.WL(WL53));
sram_cell_6t_5 inst_cell_53_113 (.BL(BL113),.BLN(BLN113),.WL(WL53));
sram_cell_6t_5 inst_cell_53_114 (.BL(BL114),.BLN(BLN114),.WL(WL53));
sram_cell_6t_5 inst_cell_53_115 (.BL(BL115),.BLN(BLN115),.WL(WL53));
sram_cell_6t_5 inst_cell_53_116 (.BL(BL116),.BLN(BLN116),.WL(WL53));
sram_cell_6t_5 inst_cell_53_117 (.BL(BL117),.BLN(BLN117),.WL(WL53));
sram_cell_6t_5 inst_cell_53_118 (.BL(BL118),.BLN(BLN118),.WL(WL53));
sram_cell_6t_5 inst_cell_53_119 (.BL(BL119),.BLN(BLN119),.WL(WL53));
sram_cell_6t_5 inst_cell_53_120 (.BL(BL120),.BLN(BLN120),.WL(WL53));
sram_cell_6t_5 inst_cell_53_121 (.BL(BL121),.BLN(BLN121),.WL(WL53));
sram_cell_6t_5 inst_cell_53_122 (.BL(BL122),.BLN(BLN122),.WL(WL53));
sram_cell_6t_5 inst_cell_53_123 (.BL(BL123),.BLN(BLN123),.WL(WL53));
sram_cell_6t_5 inst_cell_53_124 (.BL(BL124),.BLN(BLN124),.WL(WL53));
sram_cell_6t_5 inst_cell_53_125 (.BL(BL125),.BLN(BLN125),.WL(WL53));
sram_cell_6t_5 inst_cell_53_126 (.BL(BL126),.BLN(BLN126),.WL(WL53));
sram_cell_6t_5 inst_cell_53_127 (.BL(BL127),.BLN(BLN127),.WL(WL53));
sram_cell_6t_5 inst_cell_54_0 (.BL(BL0),.BLN(BLN0),.WL(WL54));
sram_cell_6t_5 inst_cell_54_1 (.BL(BL1),.BLN(BLN1),.WL(WL54));
sram_cell_6t_5 inst_cell_54_2 (.BL(BL2),.BLN(BLN2),.WL(WL54));
sram_cell_6t_5 inst_cell_54_3 (.BL(BL3),.BLN(BLN3),.WL(WL54));
sram_cell_6t_5 inst_cell_54_4 (.BL(BL4),.BLN(BLN4),.WL(WL54));
sram_cell_6t_5 inst_cell_54_5 (.BL(BL5),.BLN(BLN5),.WL(WL54));
sram_cell_6t_5 inst_cell_54_6 (.BL(BL6),.BLN(BLN6),.WL(WL54));
sram_cell_6t_5 inst_cell_54_7 (.BL(BL7),.BLN(BLN7),.WL(WL54));
sram_cell_6t_5 inst_cell_54_8 (.BL(BL8),.BLN(BLN8),.WL(WL54));
sram_cell_6t_5 inst_cell_54_9 (.BL(BL9),.BLN(BLN9),.WL(WL54));
sram_cell_6t_5 inst_cell_54_10 (.BL(BL10),.BLN(BLN10),.WL(WL54));
sram_cell_6t_5 inst_cell_54_11 (.BL(BL11),.BLN(BLN11),.WL(WL54));
sram_cell_6t_5 inst_cell_54_12 (.BL(BL12),.BLN(BLN12),.WL(WL54));
sram_cell_6t_5 inst_cell_54_13 (.BL(BL13),.BLN(BLN13),.WL(WL54));
sram_cell_6t_5 inst_cell_54_14 (.BL(BL14),.BLN(BLN14),.WL(WL54));
sram_cell_6t_5 inst_cell_54_15 (.BL(BL15),.BLN(BLN15),.WL(WL54));
sram_cell_6t_5 inst_cell_54_16 (.BL(BL16),.BLN(BLN16),.WL(WL54));
sram_cell_6t_5 inst_cell_54_17 (.BL(BL17),.BLN(BLN17),.WL(WL54));
sram_cell_6t_5 inst_cell_54_18 (.BL(BL18),.BLN(BLN18),.WL(WL54));
sram_cell_6t_5 inst_cell_54_19 (.BL(BL19),.BLN(BLN19),.WL(WL54));
sram_cell_6t_5 inst_cell_54_20 (.BL(BL20),.BLN(BLN20),.WL(WL54));
sram_cell_6t_5 inst_cell_54_21 (.BL(BL21),.BLN(BLN21),.WL(WL54));
sram_cell_6t_5 inst_cell_54_22 (.BL(BL22),.BLN(BLN22),.WL(WL54));
sram_cell_6t_5 inst_cell_54_23 (.BL(BL23),.BLN(BLN23),.WL(WL54));
sram_cell_6t_5 inst_cell_54_24 (.BL(BL24),.BLN(BLN24),.WL(WL54));
sram_cell_6t_5 inst_cell_54_25 (.BL(BL25),.BLN(BLN25),.WL(WL54));
sram_cell_6t_5 inst_cell_54_26 (.BL(BL26),.BLN(BLN26),.WL(WL54));
sram_cell_6t_5 inst_cell_54_27 (.BL(BL27),.BLN(BLN27),.WL(WL54));
sram_cell_6t_5 inst_cell_54_28 (.BL(BL28),.BLN(BLN28),.WL(WL54));
sram_cell_6t_5 inst_cell_54_29 (.BL(BL29),.BLN(BLN29),.WL(WL54));
sram_cell_6t_5 inst_cell_54_30 (.BL(BL30),.BLN(BLN30),.WL(WL54));
sram_cell_6t_5 inst_cell_54_31 (.BL(BL31),.BLN(BLN31),.WL(WL54));
sram_cell_6t_5 inst_cell_54_32 (.BL(BL32),.BLN(BLN32),.WL(WL54));
sram_cell_6t_5 inst_cell_54_33 (.BL(BL33),.BLN(BLN33),.WL(WL54));
sram_cell_6t_5 inst_cell_54_34 (.BL(BL34),.BLN(BLN34),.WL(WL54));
sram_cell_6t_5 inst_cell_54_35 (.BL(BL35),.BLN(BLN35),.WL(WL54));
sram_cell_6t_5 inst_cell_54_36 (.BL(BL36),.BLN(BLN36),.WL(WL54));
sram_cell_6t_5 inst_cell_54_37 (.BL(BL37),.BLN(BLN37),.WL(WL54));
sram_cell_6t_5 inst_cell_54_38 (.BL(BL38),.BLN(BLN38),.WL(WL54));
sram_cell_6t_5 inst_cell_54_39 (.BL(BL39),.BLN(BLN39),.WL(WL54));
sram_cell_6t_5 inst_cell_54_40 (.BL(BL40),.BLN(BLN40),.WL(WL54));
sram_cell_6t_5 inst_cell_54_41 (.BL(BL41),.BLN(BLN41),.WL(WL54));
sram_cell_6t_5 inst_cell_54_42 (.BL(BL42),.BLN(BLN42),.WL(WL54));
sram_cell_6t_5 inst_cell_54_43 (.BL(BL43),.BLN(BLN43),.WL(WL54));
sram_cell_6t_5 inst_cell_54_44 (.BL(BL44),.BLN(BLN44),.WL(WL54));
sram_cell_6t_5 inst_cell_54_45 (.BL(BL45),.BLN(BLN45),.WL(WL54));
sram_cell_6t_5 inst_cell_54_46 (.BL(BL46),.BLN(BLN46),.WL(WL54));
sram_cell_6t_5 inst_cell_54_47 (.BL(BL47),.BLN(BLN47),.WL(WL54));
sram_cell_6t_5 inst_cell_54_48 (.BL(BL48),.BLN(BLN48),.WL(WL54));
sram_cell_6t_5 inst_cell_54_49 (.BL(BL49),.BLN(BLN49),.WL(WL54));
sram_cell_6t_5 inst_cell_54_50 (.BL(BL50),.BLN(BLN50),.WL(WL54));
sram_cell_6t_5 inst_cell_54_51 (.BL(BL51),.BLN(BLN51),.WL(WL54));
sram_cell_6t_5 inst_cell_54_52 (.BL(BL52),.BLN(BLN52),.WL(WL54));
sram_cell_6t_5 inst_cell_54_53 (.BL(BL53),.BLN(BLN53),.WL(WL54));
sram_cell_6t_5 inst_cell_54_54 (.BL(BL54),.BLN(BLN54),.WL(WL54));
sram_cell_6t_5 inst_cell_54_55 (.BL(BL55),.BLN(BLN55),.WL(WL54));
sram_cell_6t_5 inst_cell_54_56 (.BL(BL56),.BLN(BLN56),.WL(WL54));
sram_cell_6t_5 inst_cell_54_57 (.BL(BL57),.BLN(BLN57),.WL(WL54));
sram_cell_6t_5 inst_cell_54_58 (.BL(BL58),.BLN(BLN58),.WL(WL54));
sram_cell_6t_5 inst_cell_54_59 (.BL(BL59),.BLN(BLN59),.WL(WL54));
sram_cell_6t_5 inst_cell_54_60 (.BL(BL60),.BLN(BLN60),.WL(WL54));
sram_cell_6t_5 inst_cell_54_61 (.BL(BL61),.BLN(BLN61),.WL(WL54));
sram_cell_6t_5 inst_cell_54_62 (.BL(BL62),.BLN(BLN62),.WL(WL54));
sram_cell_6t_5 inst_cell_54_63 (.BL(BL63),.BLN(BLN63),.WL(WL54));
sram_cell_6t_5 inst_cell_54_64 (.BL(BL64),.BLN(BLN64),.WL(WL54));
sram_cell_6t_5 inst_cell_54_65 (.BL(BL65),.BLN(BLN65),.WL(WL54));
sram_cell_6t_5 inst_cell_54_66 (.BL(BL66),.BLN(BLN66),.WL(WL54));
sram_cell_6t_5 inst_cell_54_67 (.BL(BL67),.BLN(BLN67),.WL(WL54));
sram_cell_6t_5 inst_cell_54_68 (.BL(BL68),.BLN(BLN68),.WL(WL54));
sram_cell_6t_5 inst_cell_54_69 (.BL(BL69),.BLN(BLN69),.WL(WL54));
sram_cell_6t_5 inst_cell_54_70 (.BL(BL70),.BLN(BLN70),.WL(WL54));
sram_cell_6t_5 inst_cell_54_71 (.BL(BL71),.BLN(BLN71),.WL(WL54));
sram_cell_6t_5 inst_cell_54_72 (.BL(BL72),.BLN(BLN72),.WL(WL54));
sram_cell_6t_5 inst_cell_54_73 (.BL(BL73),.BLN(BLN73),.WL(WL54));
sram_cell_6t_5 inst_cell_54_74 (.BL(BL74),.BLN(BLN74),.WL(WL54));
sram_cell_6t_5 inst_cell_54_75 (.BL(BL75),.BLN(BLN75),.WL(WL54));
sram_cell_6t_5 inst_cell_54_76 (.BL(BL76),.BLN(BLN76),.WL(WL54));
sram_cell_6t_5 inst_cell_54_77 (.BL(BL77),.BLN(BLN77),.WL(WL54));
sram_cell_6t_5 inst_cell_54_78 (.BL(BL78),.BLN(BLN78),.WL(WL54));
sram_cell_6t_5 inst_cell_54_79 (.BL(BL79),.BLN(BLN79),.WL(WL54));
sram_cell_6t_5 inst_cell_54_80 (.BL(BL80),.BLN(BLN80),.WL(WL54));
sram_cell_6t_5 inst_cell_54_81 (.BL(BL81),.BLN(BLN81),.WL(WL54));
sram_cell_6t_5 inst_cell_54_82 (.BL(BL82),.BLN(BLN82),.WL(WL54));
sram_cell_6t_5 inst_cell_54_83 (.BL(BL83),.BLN(BLN83),.WL(WL54));
sram_cell_6t_5 inst_cell_54_84 (.BL(BL84),.BLN(BLN84),.WL(WL54));
sram_cell_6t_5 inst_cell_54_85 (.BL(BL85),.BLN(BLN85),.WL(WL54));
sram_cell_6t_5 inst_cell_54_86 (.BL(BL86),.BLN(BLN86),.WL(WL54));
sram_cell_6t_5 inst_cell_54_87 (.BL(BL87),.BLN(BLN87),.WL(WL54));
sram_cell_6t_5 inst_cell_54_88 (.BL(BL88),.BLN(BLN88),.WL(WL54));
sram_cell_6t_5 inst_cell_54_89 (.BL(BL89),.BLN(BLN89),.WL(WL54));
sram_cell_6t_5 inst_cell_54_90 (.BL(BL90),.BLN(BLN90),.WL(WL54));
sram_cell_6t_5 inst_cell_54_91 (.BL(BL91),.BLN(BLN91),.WL(WL54));
sram_cell_6t_5 inst_cell_54_92 (.BL(BL92),.BLN(BLN92),.WL(WL54));
sram_cell_6t_5 inst_cell_54_93 (.BL(BL93),.BLN(BLN93),.WL(WL54));
sram_cell_6t_5 inst_cell_54_94 (.BL(BL94),.BLN(BLN94),.WL(WL54));
sram_cell_6t_5 inst_cell_54_95 (.BL(BL95),.BLN(BLN95),.WL(WL54));
sram_cell_6t_5 inst_cell_54_96 (.BL(BL96),.BLN(BLN96),.WL(WL54));
sram_cell_6t_5 inst_cell_54_97 (.BL(BL97),.BLN(BLN97),.WL(WL54));
sram_cell_6t_5 inst_cell_54_98 (.BL(BL98),.BLN(BLN98),.WL(WL54));
sram_cell_6t_5 inst_cell_54_99 (.BL(BL99),.BLN(BLN99),.WL(WL54));
sram_cell_6t_5 inst_cell_54_100 (.BL(BL100),.BLN(BLN100),.WL(WL54));
sram_cell_6t_5 inst_cell_54_101 (.BL(BL101),.BLN(BLN101),.WL(WL54));
sram_cell_6t_5 inst_cell_54_102 (.BL(BL102),.BLN(BLN102),.WL(WL54));
sram_cell_6t_5 inst_cell_54_103 (.BL(BL103),.BLN(BLN103),.WL(WL54));
sram_cell_6t_5 inst_cell_54_104 (.BL(BL104),.BLN(BLN104),.WL(WL54));
sram_cell_6t_5 inst_cell_54_105 (.BL(BL105),.BLN(BLN105),.WL(WL54));
sram_cell_6t_5 inst_cell_54_106 (.BL(BL106),.BLN(BLN106),.WL(WL54));
sram_cell_6t_5 inst_cell_54_107 (.BL(BL107),.BLN(BLN107),.WL(WL54));
sram_cell_6t_5 inst_cell_54_108 (.BL(BL108),.BLN(BLN108),.WL(WL54));
sram_cell_6t_5 inst_cell_54_109 (.BL(BL109),.BLN(BLN109),.WL(WL54));
sram_cell_6t_5 inst_cell_54_110 (.BL(BL110),.BLN(BLN110),.WL(WL54));
sram_cell_6t_5 inst_cell_54_111 (.BL(BL111),.BLN(BLN111),.WL(WL54));
sram_cell_6t_5 inst_cell_54_112 (.BL(BL112),.BLN(BLN112),.WL(WL54));
sram_cell_6t_5 inst_cell_54_113 (.BL(BL113),.BLN(BLN113),.WL(WL54));
sram_cell_6t_5 inst_cell_54_114 (.BL(BL114),.BLN(BLN114),.WL(WL54));
sram_cell_6t_5 inst_cell_54_115 (.BL(BL115),.BLN(BLN115),.WL(WL54));
sram_cell_6t_5 inst_cell_54_116 (.BL(BL116),.BLN(BLN116),.WL(WL54));
sram_cell_6t_5 inst_cell_54_117 (.BL(BL117),.BLN(BLN117),.WL(WL54));
sram_cell_6t_5 inst_cell_54_118 (.BL(BL118),.BLN(BLN118),.WL(WL54));
sram_cell_6t_5 inst_cell_54_119 (.BL(BL119),.BLN(BLN119),.WL(WL54));
sram_cell_6t_5 inst_cell_54_120 (.BL(BL120),.BLN(BLN120),.WL(WL54));
sram_cell_6t_5 inst_cell_54_121 (.BL(BL121),.BLN(BLN121),.WL(WL54));
sram_cell_6t_5 inst_cell_54_122 (.BL(BL122),.BLN(BLN122),.WL(WL54));
sram_cell_6t_5 inst_cell_54_123 (.BL(BL123),.BLN(BLN123),.WL(WL54));
sram_cell_6t_5 inst_cell_54_124 (.BL(BL124),.BLN(BLN124),.WL(WL54));
sram_cell_6t_5 inst_cell_54_125 (.BL(BL125),.BLN(BLN125),.WL(WL54));
sram_cell_6t_5 inst_cell_54_126 (.BL(BL126),.BLN(BLN126),.WL(WL54));
sram_cell_6t_5 inst_cell_54_127 (.BL(BL127),.BLN(BLN127),.WL(WL54));
sram_cell_6t_5 inst_cell_55_0 (.BL(BL0),.BLN(BLN0),.WL(WL55));
sram_cell_6t_5 inst_cell_55_1 (.BL(BL1),.BLN(BLN1),.WL(WL55));
sram_cell_6t_5 inst_cell_55_2 (.BL(BL2),.BLN(BLN2),.WL(WL55));
sram_cell_6t_5 inst_cell_55_3 (.BL(BL3),.BLN(BLN3),.WL(WL55));
sram_cell_6t_5 inst_cell_55_4 (.BL(BL4),.BLN(BLN4),.WL(WL55));
sram_cell_6t_5 inst_cell_55_5 (.BL(BL5),.BLN(BLN5),.WL(WL55));
sram_cell_6t_5 inst_cell_55_6 (.BL(BL6),.BLN(BLN6),.WL(WL55));
sram_cell_6t_5 inst_cell_55_7 (.BL(BL7),.BLN(BLN7),.WL(WL55));
sram_cell_6t_5 inst_cell_55_8 (.BL(BL8),.BLN(BLN8),.WL(WL55));
sram_cell_6t_5 inst_cell_55_9 (.BL(BL9),.BLN(BLN9),.WL(WL55));
sram_cell_6t_5 inst_cell_55_10 (.BL(BL10),.BLN(BLN10),.WL(WL55));
sram_cell_6t_5 inst_cell_55_11 (.BL(BL11),.BLN(BLN11),.WL(WL55));
sram_cell_6t_5 inst_cell_55_12 (.BL(BL12),.BLN(BLN12),.WL(WL55));
sram_cell_6t_5 inst_cell_55_13 (.BL(BL13),.BLN(BLN13),.WL(WL55));
sram_cell_6t_5 inst_cell_55_14 (.BL(BL14),.BLN(BLN14),.WL(WL55));
sram_cell_6t_5 inst_cell_55_15 (.BL(BL15),.BLN(BLN15),.WL(WL55));
sram_cell_6t_5 inst_cell_55_16 (.BL(BL16),.BLN(BLN16),.WL(WL55));
sram_cell_6t_5 inst_cell_55_17 (.BL(BL17),.BLN(BLN17),.WL(WL55));
sram_cell_6t_5 inst_cell_55_18 (.BL(BL18),.BLN(BLN18),.WL(WL55));
sram_cell_6t_5 inst_cell_55_19 (.BL(BL19),.BLN(BLN19),.WL(WL55));
sram_cell_6t_5 inst_cell_55_20 (.BL(BL20),.BLN(BLN20),.WL(WL55));
sram_cell_6t_5 inst_cell_55_21 (.BL(BL21),.BLN(BLN21),.WL(WL55));
sram_cell_6t_5 inst_cell_55_22 (.BL(BL22),.BLN(BLN22),.WL(WL55));
sram_cell_6t_5 inst_cell_55_23 (.BL(BL23),.BLN(BLN23),.WL(WL55));
sram_cell_6t_5 inst_cell_55_24 (.BL(BL24),.BLN(BLN24),.WL(WL55));
sram_cell_6t_5 inst_cell_55_25 (.BL(BL25),.BLN(BLN25),.WL(WL55));
sram_cell_6t_5 inst_cell_55_26 (.BL(BL26),.BLN(BLN26),.WL(WL55));
sram_cell_6t_5 inst_cell_55_27 (.BL(BL27),.BLN(BLN27),.WL(WL55));
sram_cell_6t_5 inst_cell_55_28 (.BL(BL28),.BLN(BLN28),.WL(WL55));
sram_cell_6t_5 inst_cell_55_29 (.BL(BL29),.BLN(BLN29),.WL(WL55));
sram_cell_6t_5 inst_cell_55_30 (.BL(BL30),.BLN(BLN30),.WL(WL55));
sram_cell_6t_5 inst_cell_55_31 (.BL(BL31),.BLN(BLN31),.WL(WL55));
sram_cell_6t_5 inst_cell_55_32 (.BL(BL32),.BLN(BLN32),.WL(WL55));
sram_cell_6t_5 inst_cell_55_33 (.BL(BL33),.BLN(BLN33),.WL(WL55));
sram_cell_6t_5 inst_cell_55_34 (.BL(BL34),.BLN(BLN34),.WL(WL55));
sram_cell_6t_5 inst_cell_55_35 (.BL(BL35),.BLN(BLN35),.WL(WL55));
sram_cell_6t_5 inst_cell_55_36 (.BL(BL36),.BLN(BLN36),.WL(WL55));
sram_cell_6t_5 inst_cell_55_37 (.BL(BL37),.BLN(BLN37),.WL(WL55));
sram_cell_6t_5 inst_cell_55_38 (.BL(BL38),.BLN(BLN38),.WL(WL55));
sram_cell_6t_5 inst_cell_55_39 (.BL(BL39),.BLN(BLN39),.WL(WL55));
sram_cell_6t_5 inst_cell_55_40 (.BL(BL40),.BLN(BLN40),.WL(WL55));
sram_cell_6t_5 inst_cell_55_41 (.BL(BL41),.BLN(BLN41),.WL(WL55));
sram_cell_6t_5 inst_cell_55_42 (.BL(BL42),.BLN(BLN42),.WL(WL55));
sram_cell_6t_5 inst_cell_55_43 (.BL(BL43),.BLN(BLN43),.WL(WL55));
sram_cell_6t_5 inst_cell_55_44 (.BL(BL44),.BLN(BLN44),.WL(WL55));
sram_cell_6t_5 inst_cell_55_45 (.BL(BL45),.BLN(BLN45),.WL(WL55));
sram_cell_6t_5 inst_cell_55_46 (.BL(BL46),.BLN(BLN46),.WL(WL55));
sram_cell_6t_5 inst_cell_55_47 (.BL(BL47),.BLN(BLN47),.WL(WL55));
sram_cell_6t_5 inst_cell_55_48 (.BL(BL48),.BLN(BLN48),.WL(WL55));
sram_cell_6t_5 inst_cell_55_49 (.BL(BL49),.BLN(BLN49),.WL(WL55));
sram_cell_6t_5 inst_cell_55_50 (.BL(BL50),.BLN(BLN50),.WL(WL55));
sram_cell_6t_5 inst_cell_55_51 (.BL(BL51),.BLN(BLN51),.WL(WL55));
sram_cell_6t_5 inst_cell_55_52 (.BL(BL52),.BLN(BLN52),.WL(WL55));
sram_cell_6t_5 inst_cell_55_53 (.BL(BL53),.BLN(BLN53),.WL(WL55));
sram_cell_6t_5 inst_cell_55_54 (.BL(BL54),.BLN(BLN54),.WL(WL55));
sram_cell_6t_5 inst_cell_55_55 (.BL(BL55),.BLN(BLN55),.WL(WL55));
sram_cell_6t_5 inst_cell_55_56 (.BL(BL56),.BLN(BLN56),.WL(WL55));
sram_cell_6t_5 inst_cell_55_57 (.BL(BL57),.BLN(BLN57),.WL(WL55));
sram_cell_6t_5 inst_cell_55_58 (.BL(BL58),.BLN(BLN58),.WL(WL55));
sram_cell_6t_5 inst_cell_55_59 (.BL(BL59),.BLN(BLN59),.WL(WL55));
sram_cell_6t_5 inst_cell_55_60 (.BL(BL60),.BLN(BLN60),.WL(WL55));
sram_cell_6t_5 inst_cell_55_61 (.BL(BL61),.BLN(BLN61),.WL(WL55));
sram_cell_6t_5 inst_cell_55_62 (.BL(BL62),.BLN(BLN62),.WL(WL55));
sram_cell_6t_5 inst_cell_55_63 (.BL(BL63),.BLN(BLN63),.WL(WL55));
sram_cell_6t_5 inst_cell_55_64 (.BL(BL64),.BLN(BLN64),.WL(WL55));
sram_cell_6t_5 inst_cell_55_65 (.BL(BL65),.BLN(BLN65),.WL(WL55));
sram_cell_6t_5 inst_cell_55_66 (.BL(BL66),.BLN(BLN66),.WL(WL55));
sram_cell_6t_5 inst_cell_55_67 (.BL(BL67),.BLN(BLN67),.WL(WL55));
sram_cell_6t_5 inst_cell_55_68 (.BL(BL68),.BLN(BLN68),.WL(WL55));
sram_cell_6t_5 inst_cell_55_69 (.BL(BL69),.BLN(BLN69),.WL(WL55));
sram_cell_6t_5 inst_cell_55_70 (.BL(BL70),.BLN(BLN70),.WL(WL55));
sram_cell_6t_5 inst_cell_55_71 (.BL(BL71),.BLN(BLN71),.WL(WL55));
sram_cell_6t_5 inst_cell_55_72 (.BL(BL72),.BLN(BLN72),.WL(WL55));
sram_cell_6t_5 inst_cell_55_73 (.BL(BL73),.BLN(BLN73),.WL(WL55));
sram_cell_6t_5 inst_cell_55_74 (.BL(BL74),.BLN(BLN74),.WL(WL55));
sram_cell_6t_5 inst_cell_55_75 (.BL(BL75),.BLN(BLN75),.WL(WL55));
sram_cell_6t_5 inst_cell_55_76 (.BL(BL76),.BLN(BLN76),.WL(WL55));
sram_cell_6t_5 inst_cell_55_77 (.BL(BL77),.BLN(BLN77),.WL(WL55));
sram_cell_6t_5 inst_cell_55_78 (.BL(BL78),.BLN(BLN78),.WL(WL55));
sram_cell_6t_5 inst_cell_55_79 (.BL(BL79),.BLN(BLN79),.WL(WL55));
sram_cell_6t_5 inst_cell_55_80 (.BL(BL80),.BLN(BLN80),.WL(WL55));
sram_cell_6t_5 inst_cell_55_81 (.BL(BL81),.BLN(BLN81),.WL(WL55));
sram_cell_6t_5 inst_cell_55_82 (.BL(BL82),.BLN(BLN82),.WL(WL55));
sram_cell_6t_5 inst_cell_55_83 (.BL(BL83),.BLN(BLN83),.WL(WL55));
sram_cell_6t_5 inst_cell_55_84 (.BL(BL84),.BLN(BLN84),.WL(WL55));
sram_cell_6t_5 inst_cell_55_85 (.BL(BL85),.BLN(BLN85),.WL(WL55));
sram_cell_6t_5 inst_cell_55_86 (.BL(BL86),.BLN(BLN86),.WL(WL55));
sram_cell_6t_5 inst_cell_55_87 (.BL(BL87),.BLN(BLN87),.WL(WL55));
sram_cell_6t_5 inst_cell_55_88 (.BL(BL88),.BLN(BLN88),.WL(WL55));
sram_cell_6t_5 inst_cell_55_89 (.BL(BL89),.BLN(BLN89),.WL(WL55));
sram_cell_6t_5 inst_cell_55_90 (.BL(BL90),.BLN(BLN90),.WL(WL55));
sram_cell_6t_5 inst_cell_55_91 (.BL(BL91),.BLN(BLN91),.WL(WL55));
sram_cell_6t_5 inst_cell_55_92 (.BL(BL92),.BLN(BLN92),.WL(WL55));
sram_cell_6t_5 inst_cell_55_93 (.BL(BL93),.BLN(BLN93),.WL(WL55));
sram_cell_6t_5 inst_cell_55_94 (.BL(BL94),.BLN(BLN94),.WL(WL55));
sram_cell_6t_5 inst_cell_55_95 (.BL(BL95),.BLN(BLN95),.WL(WL55));
sram_cell_6t_5 inst_cell_55_96 (.BL(BL96),.BLN(BLN96),.WL(WL55));
sram_cell_6t_5 inst_cell_55_97 (.BL(BL97),.BLN(BLN97),.WL(WL55));
sram_cell_6t_5 inst_cell_55_98 (.BL(BL98),.BLN(BLN98),.WL(WL55));
sram_cell_6t_5 inst_cell_55_99 (.BL(BL99),.BLN(BLN99),.WL(WL55));
sram_cell_6t_5 inst_cell_55_100 (.BL(BL100),.BLN(BLN100),.WL(WL55));
sram_cell_6t_5 inst_cell_55_101 (.BL(BL101),.BLN(BLN101),.WL(WL55));
sram_cell_6t_5 inst_cell_55_102 (.BL(BL102),.BLN(BLN102),.WL(WL55));
sram_cell_6t_5 inst_cell_55_103 (.BL(BL103),.BLN(BLN103),.WL(WL55));
sram_cell_6t_5 inst_cell_55_104 (.BL(BL104),.BLN(BLN104),.WL(WL55));
sram_cell_6t_5 inst_cell_55_105 (.BL(BL105),.BLN(BLN105),.WL(WL55));
sram_cell_6t_5 inst_cell_55_106 (.BL(BL106),.BLN(BLN106),.WL(WL55));
sram_cell_6t_5 inst_cell_55_107 (.BL(BL107),.BLN(BLN107),.WL(WL55));
sram_cell_6t_5 inst_cell_55_108 (.BL(BL108),.BLN(BLN108),.WL(WL55));
sram_cell_6t_5 inst_cell_55_109 (.BL(BL109),.BLN(BLN109),.WL(WL55));
sram_cell_6t_5 inst_cell_55_110 (.BL(BL110),.BLN(BLN110),.WL(WL55));
sram_cell_6t_5 inst_cell_55_111 (.BL(BL111),.BLN(BLN111),.WL(WL55));
sram_cell_6t_5 inst_cell_55_112 (.BL(BL112),.BLN(BLN112),.WL(WL55));
sram_cell_6t_5 inst_cell_55_113 (.BL(BL113),.BLN(BLN113),.WL(WL55));
sram_cell_6t_5 inst_cell_55_114 (.BL(BL114),.BLN(BLN114),.WL(WL55));
sram_cell_6t_5 inst_cell_55_115 (.BL(BL115),.BLN(BLN115),.WL(WL55));
sram_cell_6t_5 inst_cell_55_116 (.BL(BL116),.BLN(BLN116),.WL(WL55));
sram_cell_6t_5 inst_cell_55_117 (.BL(BL117),.BLN(BLN117),.WL(WL55));
sram_cell_6t_5 inst_cell_55_118 (.BL(BL118),.BLN(BLN118),.WL(WL55));
sram_cell_6t_5 inst_cell_55_119 (.BL(BL119),.BLN(BLN119),.WL(WL55));
sram_cell_6t_5 inst_cell_55_120 (.BL(BL120),.BLN(BLN120),.WL(WL55));
sram_cell_6t_5 inst_cell_55_121 (.BL(BL121),.BLN(BLN121),.WL(WL55));
sram_cell_6t_5 inst_cell_55_122 (.BL(BL122),.BLN(BLN122),.WL(WL55));
sram_cell_6t_5 inst_cell_55_123 (.BL(BL123),.BLN(BLN123),.WL(WL55));
sram_cell_6t_5 inst_cell_55_124 (.BL(BL124),.BLN(BLN124),.WL(WL55));
sram_cell_6t_5 inst_cell_55_125 (.BL(BL125),.BLN(BLN125),.WL(WL55));
sram_cell_6t_5 inst_cell_55_126 (.BL(BL126),.BLN(BLN126),.WL(WL55));
sram_cell_6t_5 inst_cell_55_127 (.BL(BL127),.BLN(BLN127),.WL(WL55));
sram_cell_6t_5 inst_cell_56_0 (.BL(BL0),.BLN(BLN0),.WL(WL56));
sram_cell_6t_5 inst_cell_56_1 (.BL(BL1),.BLN(BLN1),.WL(WL56));
sram_cell_6t_5 inst_cell_56_2 (.BL(BL2),.BLN(BLN2),.WL(WL56));
sram_cell_6t_5 inst_cell_56_3 (.BL(BL3),.BLN(BLN3),.WL(WL56));
sram_cell_6t_5 inst_cell_56_4 (.BL(BL4),.BLN(BLN4),.WL(WL56));
sram_cell_6t_5 inst_cell_56_5 (.BL(BL5),.BLN(BLN5),.WL(WL56));
sram_cell_6t_5 inst_cell_56_6 (.BL(BL6),.BLN(BLN6),.WL(WL56));
sram_cell_6t_5 inst_cell_56_7 (.BL(BL7),.BLN(BLN7),.WL(WL56));
sram_cell_6t_5 inst_cell_56_8 (.BL(BL8),.BLN(BLN8),.WL(WL56));
sram_cell_6t_5 inst_cell_56_9 (.BL(BL9),.BLN(BLN9),.WL(WL56));
sram_cell_6t_5 inst_cell_56_10 (.BL(BL10),.BLN(BLN10),.WL(WL56));
sram_cell_6t_5 inst_cell_56_11 (.BL(BL11),.BLN(BLN11),.WL(WL56));
sram_cell_6t_5 inst_cell_56_12 (.BL(BL12),.BLN(BLN12),.WL(WL56));
sram_cell_6t_5 inst_cell_56_13 (.BL(BL13),.BLN(BLN13),.WL(WL56));
sram_cell_6t_5 inst_cell_56_14 (.BL(BL14),.BLN(BLN14),.WL(WL56));
sram_cell_6t_5 inst_cell_56_15 (.BL(BL15),.BLN(BLN15),.WL(WL56));
sram_cell_6t_5 inst_cell_56_16 (.BL(BL16),.BLN(BLN16),.WL(WL56));
sram_cell_6t_5 inst_cell_56_17 (.BL(BL17),.BLN(BLN17),.WL(WL56));
sram_cell_6t_5 inst_cell_56_18 (.BL(BL18),.BLN(BLN18),.WL(WL56));
sram_cell_6t_5 inst_cell_56_19 (.BL(BL19),.BLN(BLN19),.WL(WL56));
sram_cell_6t_5 inst_cell_56_20 (.BL(BL20),.BLN(BLN20),.WL(WL56));
sram_cell_6t_5 inst_cell_56_21 (.BL(BL21),.BLN(BLN21),.WL(WL56));
sram_cell_6t_5 inst_cell_56_22 (.BL(BL22),.BLN(BLN22),.WL(WL56));
sram_cell_6t_5 inst_cell_56_23 (.BL(BL23),.BLN(BLN23),.WL(WL56));
sram_cell_6t_5 inst_cell_56_24 (.BL(BL24),.BLN(BLN24),.WL(WL56));
sram_cell_6t_5 inst_cell_56_25 (.BL(BL25),.BLN(BLN25),.WL(WL56));
sram_cell_6t_5 inst_cell_56_26 (.BL(BL26),.BLN(BLN26),.WL(WL56));
sram_cell_6t_5 inst_cell_56_27 (.BL(BL27),.BLN(BLN27),.WL(WL56));
sram_cell_6t_5 inst_cell_56_28 (.BL(BL28),.BLN(BLN28),.WL(WL56));
sram_cell_6t_5 inst_cell_56_29 (.BL(BL29),.BLN(BLN29),.WL(WL56));
sram_cell_6t_5 inst_cell_56_30 (.BL(BL30),.BLN(BLN30),.WL(WL56));
sram_cell_6t_5 inst_cell_56_31 (.BL(BL31),.BLN(BLN31),.WL(WL56));
sram_cell_6t_5 inst_cell_56_32 (.BL(BL32),.BLN(BLN32),.WL(WL56));
sram_cell_6t_5 inst_cell_56_33 (.BL(BL33),.BLN(BLN33),.WL(WL56));
sram_cell_6t_5 inst_cell_56_34 (.BL(BL34),.BLN(BLN34),.WL(WL56));
sram_cell_6t_5 inst_cell_56_35 (.BL(BL35),.BLN(BLN35),.WL(WL56));
sram_cell_6t_5 inst_cell_56_36 (.BL(BL36),.BLN(BLN36),.WL(WL56));
sram_cell_6t_5 inst_cell_56_37 (.BL(BL37),.BLN(BLN37),.WL(WL56));
sram_cell_6t_5 inst_cell_56_38 (.BL(BL38),.BLN(BLN38),.WL(WL56));
sram_cell_6t_5 inst_cell_56_39 (.BL(BL39),.BLN(BLN39),.WL(WL56));
sram_cell_6t_5 inst_cell_56_40 (.BL(BL40),.BLN(BLN40),.WL(WL56));
sram_cell_6t_5 inst_cell_56_41 (.BL(BL41),.BLN(BLN41),.WL(WL56));
sram_cell_6t_5 inst_cell_56_42 (.BL(BL42),.BLN(BLN42),.WL(WL56));
sram_cell_6t_5 inst_cell_56_43 (.BL(BL43),.BLN(BLN43),.WL(WL56));
sram_cell_6t_5 inst_cell_56_44 (.BL(BL44),.BLN(BLN44),.WL(WL56));
sram_cell_6t_5 inst_cell_56_45 (.BL(BL45),.BLN(BLN45),.WL(WL56));
sram_cell_6t_5 inst_cell_56_46 (.BL(BL46),.BLN(BLN46),.WL(WL56));
sram_cell_6t_5 inst_cell_56_47 (.BL(BL47),.BLN(BLN47),.WL(WL56));
sram_cell_6t_5 inst_cell_56_48 (.BL(BL48),.BLN(BLN48),.WL(WL56));
sram_cell_6t_5 inst_cell_56_49 (.BL(BL49),.BLN(BLN49),.WL(WL56));
sram_cell_6t_5 inst_cell_56_50 (.BL(BL50),.BLN(BLN50),.WL(WL56));
sram_cell_6t_5 inst_cell_56_51 (.BL(BL51),.BLN(BLN51),.WL(WL56));
sram_cell_6t_5 inst_cell_56_52 (.BL(BL52),.BLN(BLN52),.WL(WL56));
sram_cell_6t_5 inst_cell_56_53 (.BL(BL53),.BLN(BLN53),.WL(WL56));
sram_cell_6t_5 inst_cell_56_54 (.BL(BL54),.BLN(BLN54),.WL(WL56));
sram_cell_6t_5 inst_cell_56_55 (.BL(BL55),.BLN(BLN55),.WL(WL56));
sram_cell_6t_5 inst_cell_56_56 (.BL(BL56),.BLN(BLN56),.WL(WL56));
sram_cell_6t_5 inst_cell_56_57 (.BL(BL57),.BLN(BLN57),.WL(WL56));
sram_cell_6t_5 inst_cell_56_58 (.BL(BL58),.BLN(BLN58),.WL(WL56));
sram_cell_6t_5 inst_cell_56_59 (.BL(BL59),.BLN(BLN59),.WL(WL56));
sram_cell_6t_5 inst_cell_56_60 (.BL(BL60),.BLN(BLN60),.WL(WL56));
sram_cell_6t_5 inst_cell_56_61 (.BL(BL61),.BLN(BLN61),.WL(WL56));
sram_cell_6t_5 inst_cell_56_62 (.BL(BL62),.BLN(BLN62),.WL(WL56));
sram_cell_6t_5 inst_cell_56_63 (.BL(BL63),.BLN(BLN63),.WL(WL56));
sram_cell_6t_5 inst_cell_56_64 (.BL(BL64),.BLN(BLN64),.WL(WL56));
sram_cell_6t_5 inst_cell_56_65 (.BL(BL65),.BLN(BLN65),.WL(WL56));
sram_cell_6t_5 inst_cell_56_66 (.BL(BL66),.BLN(BLN66),.WL(WL56));
sram_cell_6t_5 inst_cell_56_67 (.BL(BL67),.BLN(BLN67),.WL(WL56));
sram_cell_6t_5 inst_cell_56_68 (.BL(BL68),.BLN(BLN68),.WL(WL56));
sram_cell_6t_5 inst_cell_56_69 (.BL(BL69),.BLN(BLN69),.WL(WL56));
sram_cell_6t_5 inst_cell_56_70 (.BL(BL70),.BLN(BLN70),.WL(WL56));
sram_cell_6t_5 inst_cell_56_71 (.BL(BL71),.BLN(BLN71),.WL(WL56));
sram_cell_6t_5 inst_cell_56_72 (.BL(BL72),.BLN(BLN72),.WL(WL56));
sram_cell_6t_5 inst_cell_56_73 (.BL(BL73),.BLN(BLN73),.WL(WL56));
sram_cell_6t_5 inst_cell_56_74 (.BL(BL74),.BLN(BLN74),.WL(WL56));
sram_cell_6t_5 inst_cell_56_75 (.BL(BL75),.BLN(BLN75),.WL(WL56));
sram_cell_6t_5 inst_cell_56_76 (.BL(BL76),.BLN(BLN76),.WL(WL56));
sram_cell_6t_5 inst_cell_56_77 (.BL(BL77),.BLN(BLN77),.WL(WL56));
sram_cell_6t_5 inst_cell_56_78 (.BL(BL78),.BLN(BLN78),.WL(WL56));
sram_cell_6t_5 inst_cell_56_79 (.BL(BL79),.BLN(BLN79),.WL(WL56));
sram_cell_6t_5 inst_cell_56_80 (.BL(BL80),.BLN(BLN80),.WL(WL56));
sram_cell_6t_5 inst_cell_56_81 (.BL(BL81),.BLN(BLN81),.WL(WL56));
sram_cell_6t_5 inst_cell_56_82 (.BL(BL82),.BLN(BLN82),.WL(WL56));
sram_cell_6t_5 inst_cell_56_83 (.BL(BL83),.BLN(BLN83),.WL(WL56));
sram_cell_6t_5 inst_cell_56_84 (.BL(BL84),.BLN(BLN84),.WL(WL56));
sram_cell_6t_5 inst_cell_56_85 (.BL(BL85),.BLN(BLN85),.WL(WL56));
sram_cell_6t_5 inst_cell_56_86 (.BL(BL86),.BLN(BLN86),.WL(WL56));
sram_cell_6t_5 inst_cell_56_87 (.BL(BL87),.BLN(BLN87),.WL(WL56));
sram_cell_6t_5 inst_cell_56_88 (.BL(BL88),.BLN(BLN88),.WL(WL56));
sram_cell_6t_5 inst_cell_56_89 (.BL(BL89),.BLN(BLN89),.WL(WL56));
sram_cell_6t_5 inst_cell_56_90 (.BL(BL90),.BLN(BLN90),.WL(WL56));
sram_cell_6t_5 inst_cell_56_91 (.BL(BL91),.BLN(BLN91),.WL(WL56));
sram_cell_6t_5 inst_cell_56_92 (.BL(BL92),.BLN(BLN92),.WL(WL56));
sram_cell_6t_5 inst_cell_56_93 (.BL(BL93),.BLN(BLN93),.WL(WL56));
sram_cell_6t_5 inst_cell_56_94 (.BL(BL94),.BLN(BLN94),.WL(WL56));
sram_cell_6t_5 inst_cell_56_95 (.BL(BL95),.BLN(BLN95),.WL(WL56));
sram_cell_6t_5 inst_cell_56_96 (.BL(BL96),.BLN(BLN96),.WL(WL56));
sram_cell_6t_5 inst_cell_56_97 (.BL(BL97),.BLN(BLN97),.WL(WL56));
sram_cell_6t_5 inst_cell_56_98 (.BL(BL98),.BLN(BLN98),.WL(WL56));
sram_cell_6t_5 inst_cell_56_99 (.BL(BL99),.BLN(BLN99),.WL(WL56));
sram_cell_6t_5 inst_cell_56_100 (.BL(BL100),.BLN(BLN100),.WL(WL56));
sram_cell_6t_5 inst_cell_56_101 (.BL(BL101),.BLN(BLN101),.WL(WL56));
sram_cell_6t_5 inst_cell_56_102 (.BL(BL102),.BLN(BLN102),.WL(WL56));
sram_cell_6t_5 inst_cell_56_103 (.BL(BL103),.BLN(BLN103),.WL(WL56));
sram_cell_6t_5 inst_cell_56_104 (.BL(BL104),.BLN(BLN104),.WL(WL56));
sram_cell_6t_5 inst_cell_56_105 (.BL(BL105),.BLN(BLN105),.WL(WL56));
sram_cell_6t_5 inst_cell_56_106 (.BL(BL106),.BLN(BLN106),.WL(WL56));
sram_cell_6t_5 inst_cell_56_107 (.BL(BL107),.BLN(BLN107),.WL(WL56));
sram_cell_6t_5 inst_cell_56_108 (.BL(BL108),.BLN(BLN108),.WL(WL56));
sram_cell_6t_5 inst_cell_56_109 (.BL(BL109),.BLN(BLN109),.WL(WL56));
sram_cell_6t_5 inst_cell_56_110 (.BL(BL110),.BLN(BLN110),.WL(WL56));
sram_cell_6t_5 inst_cell_56_111 (.BL(BL111),.BLN(BLN111),.WL(WL56));
sram_cell_6t_5 inst_cell_56_112 (.BL(BL112),.BLN(BLN112),.WL(WL56));
sram_cell_6t_5 inst_cell_56_113 (.BL(BL113),.BLN(BLN113),.WL(WL56));
sram_cell_6t_5 inst_cell_56_114 (.BL(BL114),.BLN(BLN114),.WL(WL56));
sram_cell_6t_5 inst_cell_56_115 (.BL(BL115),.BLN(BLN115),.WL(WL56));
sram_cell_6t_5 inst_cell_56_116 (.BL(BL116),.BLN(BLN116),.WL(WL56));
sram_cell_6t_5 inst_cell_56_117 (.BL(BL117),.BLN(BLN117),.WL(WL56));
sram_cell_6t_5 inst_cell_56_118 (.BL(BL118),.BLN(BLN118),.WL(WL56));
sram_cell_6t_5 inst_cell_56_119 (.BL(BL119),.BLN(BLN119),.WL(WL56));
sram_cell_6t_5 inst_cell_56_120 (.BL(BL120),.BLN(BLN120),.WL(WL56));
sram_cell_6t_5 inst_cell_56_121 (.BL(BL121),.BLN(BLN121),.WL(WL56));
sram_cell_6t_5 inst_cell_56_122 (.BL(BL122),.BLN(BLN122),.WL(WL56));
sram_cell_6t_5 inst_cell_56_123 (.BL(BL123),.BLN(BLN123),.WL(WL56));
sram_cell_6t_5 inst_cell_56_124 (.BL(BL124),.BLN(BLN124),.WL(WL56));
sram_cell_6t_5 inst_cell_56_125 (.BL(BL125),.BLN(BLN125),.WL(WL56));
sram_cell_6t_5 inst_cell_56_126 (.BL(BL126),.BLN(BLN126),.WL(WL56));
sram_cell_6t_5 inst_cell_56_127 (.BL(BL127),.BLN(BLN127),.WL(WL56));
sram_cell_6t_5 inst_cell_57_0 (.BL(BL0),.BLN(BLN0),.WL(WL57));
sram_cell_6t_5 inst_cell_57_1 (.BL(BL1),.BLN(BLN1),.WL(WL57));
sram_cell_6t_5 inst_cell_57_2 (.BL(BL2),.BLN(BLN2),.WL(WL57));
sram_cell_6t_5 inst_cell_57_3 (.BL(BL3),.BLN(BLN3),.WL(WL57));
sram_cell_6t_5 inst_cell_57_4 (.BL(BL4),.BLN(BLN4),.WL(WL57));
sram_cell_6t_5 inst_cell_57_5 (.BL(BL5),.BLN(BLN5),.WL(WL57));
sram_cell_6t_5 inst_cell_57_6 (.BL(BL6),.BLN(BLN6),.WL(WL57));
sram_cell_6t_5 inst_cell_57_7 (.BL(BL7),.BLN(BLN7),.WL(WL57));
sram_cell_6t_5 inst_cell_57_8 (.BL(BL8),.BLN(BLN8),.WL(WL57));
sram_cell_6t_5 inst_cell_57_9 (.BL(BL9),.BLN(BLN9),.WL(WL57));
sram_cell_6t_5 inst_cell_57_10 (.BL(BL10),.BLN(BLN10),.WL(WL57));
sram_cell_6t_5 inst_cell_57_11 (.BL(BL11),.BLN(BLN11),.WL(WL57));
sram_cell_6t_5 inst_cell_57_12 (.BL(BL12),.BLN(BLN12),.WL(WL57));
sram_cell_6t_5 inst_cell_57_13 (.BL(BL13),.BLN(BLN13),.WL(WL57));
sram_cell_6t_5 inst_cell_57_14 (.BL(BL14),.BLN(BLN14),.WL(WL57));
sram_cell_6t_5 inst_cell_57_15 (.BL(BL15),.BLN(BLN15),.WL(WL57));
sram_cell_6t_5 inst_cell_57_16 (.BL(BL16),.BLN(BLN16),.WL(WL57));
sram_cell_6t_5 inst_cell_57_17 (.BL(BL17),.BLN(BLN17),.WL(WL57));
sram_cell_6t_5 inst_cell_57_18 (.BL(BL18),.BLN(BLN18),.WL(WL57));
sram_cell_6t_5 inst_cell_57_19 (.BL(BL19),.BLN(BLN19),.WL(WL57));
sram_cell_6t_5 inst_cell_57_20 (.BL(BL20),.BLN(BLN20),.WL(WL57));
sram_cell_6t_5 inst_cell_57_21 (.BL(BL21),.BLN(BLN21),.WL(WL57));
sram_cell_6t_5 inst_cell_57_22 (.BL(BL22),.BLN(BLN22),.WL(WL57));
sram_cell_6t_5 inst_cell_57_23 (.BL(BL23),.BLN(BLN23),.WL(WL57));
sram_cell_6t_5 inst_cell_57_24 (.BL(BL24),.BLN(BLN24),.WL(WL57));
sram_cell_6t_5 inst_cell_57_25 (.BL(BL25),.BLN(BLN25),.WL(WL57));
sram_cell_6t_5 inst_cell_57_26 (.BL(BL26),.BLN(BLN26),.WL(WL57));
sram_cell_6t_5 inst_cell_57_27 (.BL(BL27),.BLN(BLN27),.WL(WL57));
sram_cell_6t_5 inst_cell_57_28 (.BL(BL28),.BLN(BLN28),.WL(WL57));
sram_cell_6t_5 inst_cell_57_29 (.BL(BL29),.BLN(BLN29),.WL(WL57));
sram_cell_6t_5 inst_cell_57_30 (.BL(BL30),.BLN(BLN30),.WL(WL57));
sram_cell_6t_5 inst_cell_57_31 (.BL(BL31),.BLN(BLN31),.WL(WL57));
sram_cell_6t_5 inst_cell_57_32 (.BL(BL32),.BLN(BLN32),.WL(WL57));
sram_cell_6t_5 inst_cell_57_33 (.BL(BL33),.BLN(BLN33),.WL(WL57));
sram_cell_6t_5 inst_cell_57_34 (.BL(BL34),.BLN(BLN34),.WL(WL57));
sram_cell_6t_5 inst_cell_57_35 (.BL(BL35),.BLN(BLN35),.WL(WL57));
sram_cell_6t_5 inst_cell_57_36 (.BL(BL36),.BLN(BLN36),.WL(WL57));
sram_cell_6t_5 inst_cell_57_37 (.BL(BL37),.BLN(BLN37),.WL(WL57));
sram_cell_6t_5 inst_cell_57_38 (.BL(BL38),.BLN(BLN38),.WL(WL57));
sram_cell_6t_5 inst_cell_57_39 (.BL(BL39),.BLN(BLN39),.WL(WL57));
sram_cell_6t_5 inst_cell_57_40 (.BL(BL40),.BLN(BLN40),.WL(WL57));
sram_cell_6t_5 inst_cell_57_41 (.BL(BL41),.BLN(BLN41),.WL(WL57));
sram_cell_6t_5 inst_cell_57_42 (.BL(BL42),.BLN(BLN42),.WL(WL57));
sram_cell_6t_5 inst_cell_57_43 (.BL(BL43),.BLN(BLN43),.WL(WL57));
sram_cell_6t_5 inst_cell_57_44 (.BL(BL44),.BLN(BLN44),.WL(WL57));
sram_cell_6t_5 inst_cell_57_45 (.BL(BL45),.BLN(BLN45),.WL(WL57));
sram_cell_6t_5 inst_cell_57_46 (.BL(BL46),.BLN(BLN46),.WL(WL57));
sram_cell_6t_5 inst_cell_57_47 (.BL(BL47),.BLN(BLN47),.WL(WL57));
sram_cell_6t_5 inst_cell_57_48 (.BL(BL48),.BLN(BLN48),.WL(WL57));
sram_cell_6t_5 inst_cell_57_49 (.BL(BL49),.BLN(BLN49),.WL(WL57));
sram_cell_6t_5 inst_cell_57_50 (.BL(BL50),.BLN(BLN50),.WL(WL57));
sram_cell_6t_5 inst_cell_57_51 (.BL(BL51),.BLN(BLN51),.WL(WL57));
sram_cell_6t_5 inst_cell_57_52 (.BL(BL52),.BLN(BLN52),.WL(WL57));
sram_cell_6t_5 inst_cell_57_53 (.BL(BL53),.BLN(BLN53),.WL(WL57));
sram_cell_6t_5 inst_cell_57_54 (.BL(BL54),.BLN(BLN54),.WL(WL57));
sram_cell_6t_5 inst_cell_57_55 (.BL(BL55),.BLN(BLN55),.WL(WL57));
sram_cell_6t_5 inst_cell_57_56 (.BL(BL56),.BLN(BLN56),.WL(WL57));
sram_cell_6t_5 inst_cell_57_57 (.BL(BL57),.BLN(BLN57),.WL(WL57));
sram_cell_6t_5 inst_cell_57_58 (.BL(BL58),.BLN(BLN58),.WL(WL57));
sram_cell_6t_5 inst_cell_57_59 (.BL(BL59),.BLN(BLN59),.WL(WL57));
sram_cell_6t_5 inst_cell_57_60 (.BL(BL60),.BLN(BLN60),.WL(WL57));
sram_cell_6t_5 inst_cell_57_61 (.BL(BL61),.BLN(BLN61),.WL(WL57));
sram_cell_6t_5 inst_cell_57_62 (.BL(BL62),.BLN(BLN62),.WL(WL57));
sram_cell_6t_5 inst_cell_57_63 (.BL(BL63),.BLN(BLN63),.WL(WL57));
sram_cell_6t_5 inst_cell_57_64 (.BL(BL64),.BLN(BLN64),.WL(WL57));
sram_cell_6t_5 inst_cell_57_65 (.BL(BL65),.BLN(BLN65),.WL(WL57));
sram_cell_6t_5 inst_cell_57_66 (.BL(BL66),.BLN(BLN66),.WL(WL57));
sram_cell_6t_5 inst_cell_57_67 (.BL(BL67),.BLN(BLN67),.WL(WL57));
sram_cell_6t_5 inst_cell_57_68 (.BL(BL68),.BLN(BLN68),.WL(WL57));
sram_cell_6t_5 inst_cell_57_69 (.BL(BL69),.BLN(BLN69),.WL(WL57));
sram_cell_6t_5 inst_cell_57_70 (.BL(BL70),.BLN(BLN70),.WL(WL57));
sram_cell_6t_5 inst_cell_57_71 (.BL(BL71),.BLN(BLN71),.WL(WL57));
sram_cell_6t_5 inst_cell_57_72 (.BL(BL72),.BLN(BLN72),.WL(WL57));
sram_cell_6t_5 inst_cell_57_73 (.BL(BL73),.BLN(BLN73),.WL(WL57));
sram_cell_6t_5 inst_cell_57_74 (.BL(BL74),.BLN(BLN74),.WL(WL57));
sram_cell_6t_5 inst_cell_57_75 (.BL(BL75),.BLN(BLN75),.WL(WL57));
sram_cell_6t_5 inst_cell_57_76 (.BL(BL76),.BLN(BLN76),.WL(WL57));
sram_cell_6t_5 inst_cell_57_77 (.BL(BL77),.BLN(BLN77),.WL(WL57));
sram_cell_6t_5 inst_cell_57_78 (.BL(BL78),.BLN(BLN78),.WL(WL57));
sram_cell_6t_5 inst_cell_57_79 (.BL(BL79),.BLN(BLN79),.WL(WL57));
sram_cell_6t_5 inst_cell_57_80 (.BL(BL80),.BLN(BLN80),.WL(WL57));
sram_cell_6t_5 inst_cell_57_81 (.BL(BL81),.BLN(BLN81),.WL(WL57));
sram_cell_6t_5 inst_cell_57_82 (.BL(BL82),.BLN(BLN82),.WL(WL57));
sram_cell_6t_5 inst_cell_57_83 (.BL(BL83),.BLN(BLN83),.WL(WL57));
sram_cell_6t_5 inst_cell_57_84 (.BL(BL84),.BLN(BLN84),.WL(WL57));
sram_cell_6t_5 inst_cell_57_85 (.BL(BL85),.BLN(BLN85),.WL(WL57));
sram_cell_6t_5 inst_cell_57_86 (.BL(BL86),.BLN(BLN86),.WL(WL57));
sram_cell_6t_5 inst_cell_57_87 (.BL(BL87),.BLN(BLN87),.WL(WL57));
sram_cell_6t_5 inst_cell_57_88 (.BL(BL88),.BLN(BLN88),.WL(WL57));
sram_cell_6t_5 inst_cell_57_89 (.BL(BL89),.BLN(BLN89),.WL(WL57));
sram_cell_6t_5 inst_cell_57_90 (.BL(BL90),.BLN(BLN90),.WL(WL57));
sram_cell_6t_5 inst_cell_57_91 (.BL(BL91),.BLN(BLN91),.WL(WL57));
sram_cell_6t_5 inst_cell_57_92 (.BL(BL92),.BLN(BLN92),.WL(WL57));
sram_cell_6t_5 inst_cell_57_93 (.BL(BL93),.BLN(BLN93),.WL(WL57));
sram_cell_6t_5 inst_cell_57_94 (.BL(BL94),.BLN(BLN94),.WL(WL57));
sram_cell_6t_5 inst_cell_57_95 (.BL(BL95),.BLN(BLN95),.WL(WL57));
sram_cell_6t_5 inst_cell_57_96 (.BL(BL96),.BLN(BLN96),.WL(WL57));
sram_cell_6t_5 inst_cell_57_97 (.BL(BL97),.BLN(BLN97),.WL(WL57));
sram_cell_6t_5 inst_cell_57_98 (.BL(BL98),.BLN(BLN98),.WL(WL57));
sram_cell_6t_5 inst_cell_57_99 (.BL(BL99),.BLN(BLN99),.WL(WL57));
sram_cell_6t_5 inst_cell_57_100 (.BL(BL100),.BLN(BLN100),.WL(WL57));
sram_cell_6t_5 inst_cell_57_101 (.BL(BL101),.BLN(BLN101),.WL(WL57));
sram_cell_6t_5 inst_cell_57_102 (.BL(BL102),.BLN(BLN102),.WL(WL57));
sram_cell_6t_5 inst_cell_57_103 (.BL(BL103),.BLN(BLN103),.WL(WL57));
sram_cell_6t_5 inst_cell_57_104 (.BL(BL104),.BLN(BLN104),.WL(WL57));
sram_cell_6t_5 inst_cell_57_105 (.BL(BL105),.BLN(BLN105),.WL(WL57));
sram_cell_6t_5 inst_cell_57_106 (.BL(BL106),.BLN(BLN106),.WL(WL57));
sram_cell_6t_5 inst_cell_57_107 (.BL(BL107),.BLN(BLN107),.WL(WL57));
sram_cell_6t_5 inst_cell_57_108 (.BL(BL108),.BLN(BLN108),.WL(WL57));
sram_cell_6t_5 inst_cell_57_109 (.BL(BL109),.BLN(BLN109),.WL(WL57));
sram_cell_6t_5 inst_cell_57_110 (.BL(BL110),.BLN(BLN110),.WL(WL57));
sram_cell_6t_5 inst_cell_57_111 (.BL(BL111),.BLN(BLN111),.WL(WL57));
sram_cell_6t_5 inst_cell_57_112 (.BL(BL112),.BLN(BLN112),.WL(WL57));
sram_cell_6t_5 inst_cell_57_113 (.BL(BL113),.BLN(BLN113),.WL(WL57));
sram_cell_6t_5 inst_cell_57_114 (.BL(BL114),.BLN(BLN114),.WL(WL57));
sram_cell_6t_5 inst_cell_57_115 (.BL(BL115),.BLN(BLN115),.WL(WL57));
sram_cell_6t_5 inst_cell_57_116 (.BL(BL116),.BLN(BLN116),.WL(WL57));
sram_cell_6t_5 inst_cell_57_117 (.BL(BL117),.BLN(BLN117),.WL(WL57));
sram_cell_6t_5 inst_cell_57_118 (.BL(BL118),.BLN(BLN118),.WL(WL57));
sram_cell_6t_5 inst_cell_57_119 (.BL(BL119),.BLN(BLN119),.WL(WL57));
sram_cell_6t_5 inst_cell_57_120 (.BL(BL120),.BLN(BLN120),.WL(WL57));
sram_cell_6t_5 inst_cell_57_121 (.BL(BL121),.BLN(BLN121),.WL(WL57));
sram_cell_6t_5 inst_cell_57_122 (.BL(BL122),.BLN(BLN122),.WL(WL57));
sram_cell_6t_5 inst_cell_57_123 (.BL(BL123),.BLN(BLN123),.WL(WL57));
sram_cell_6t_5 inst_cell_57_124 (.BL(BL124),.BLN(BLN124),.WL(WL57));
sram_cell_6t_5 inst_cell_57_125 (.BL(BL125),.BLN(BLN125),.WL(WL57));
sram_cell_6t_5 inst_cell_57_126 (.BL(BL126),.BLN(BLN126),.WL(WL57));
sram_cell_6t_5 inst_cell_57_127 (.BL(BL127),.BLN(BLN127),.WL(WL57));
sram_cell_6t_5 inst_cell_58_0 (.BL(BL0),.BLN(BLN0),.WL(WL58));
sram_cell_6t_5 inst_cell_58_1 (.BL(BL1),.BLN(BLN1),.WL(WL58));
sram_cell_6t_5 inst_cell_58_2 (.BL(BL2),.BLN(BLN2),.WL(WL58));
sram_cell_6t_5 inst_cell_58_3 (.BL(BL3),.BLN(BLN3),.WL(WL58));
sram_cell_6t_5 inst_cell_58_4 (.BL(BL4),.BLN(BLN4),.WL(WL58));
sram_cell_6t_5 inst_cell_58_5 (.BL(BL5),.BLN(BLN5),.WL(WL58));
sram_cell_6t_5 inst_cell_58_6 (.BL(BL6),.BLN(BLN6),.WL(WL58));
sram_cell_6t_5 inst_cell_58_7 (.BL(BL7),.BLN(BLN7),.WL(WL58));
sram_cell_6t_5 inst_cell_58_8 (.BL(BL8),.BLN(BLN8),.WL(WL58));
sram_cell_6t_5 inst_cell_58_9 (.BL(BL9),.BLN(BLN9),.WL(WL58));
sram_cell_6t_5 inst_cell_58_10 (.BL(BL10),.BLN(BLN10),.WL(WL58));
sram_cell_6t_5 inst_cell_58_11 (.BL(BL11),.BLN(BLN11),.WL(WL58));
sram_cell_6t_5 inst_cell_58_12 (.BL(BL12),.BLN(BLN12),.WL(WL58));
sram_cell_6t_5 inst_cell_58_13 (.BL(BL13),.BLN(BLN13),.WL(WL58));
sram_cell_6t_5 inst_cell_58_14 (.BL(BL14),.BLN(BLN14),.WL(WL58));
sram_cell_6t_5 inst_cell_58_15 (.BL(BL15),.BLN(BLN15),.WL(WL58));
sram_cell_6t_5 inst_cell_58_16 (.BL(BL16),.BLN(BLN16),.WL(WL58));
sram_cell_6t_5 inst_cell_58_17 (.BL(BL17),.BLN(BLN17),.WL(WL58));
sram_cell_6t_5 inst_cell_58_18 (.BL(BL18),.BLN(BLN18),.WL(WL58));
sram_cell_6t_5 inst_cell_58_19 (.BL(BL19),.BLN(BLN19),.WL(WL58));
sram_cell_6t_5 inst_cell_58_20 (.BL(BL20),.BLN(BLN20),.WL(WL58));
sram_cell_6t_5 inst_cell_58_21 (.BL(BL21),.BLN(BLN21),.WL(WL58));
sram_cell_6t_5 inst_cell_58_22 (.BL(BL22),.BLN(BLN22),.WL(WL58));
sram_cell_6t_5 inst_cell_58_23 (.BL(BL23),.BLN(BLN23),.WL(WL58));
sram_cell_6t_5 inst_cell_58_24 (.BL(BL24),.BLN(BLN24),.WL(WL58));
sram_cell_6t_5 inst_cell_58_25 (.BL(BL25),.BLN(BLN25),.WL(WL58));
sram_cell_6t_5 inst_cell_58_26 (.BL(BL26),.BLN(BLN26),.WL(WL58));
sram_cell_6t_5 inst_cell_58_27 (.BL(BL27),.BLN(BLN27),.WL(WL58));
sram_cell_6t_5 inst_cell_58_28 (.BL(BL28),.BLN(BLN28),.WL(WL58));
sram_cell_6t_5 inst_cell_58_29 (.BL(BL29),.BLN(BLN29),.WL(WL58));
sram_cell_6t_5 inst_cell_58_30 (.BL(BL30),.BLN(BLN30),.WL(WL58));
sram_cell_6t_5 inst_cell_58_31 (.BL(BL31),.BLN(BLN31),.WL(WL58));
sram_cell_6t_5 inst_cell_58_32 (.BL(BL32),.BLN(BLN32),.WL(WL58));
sram_cell_6t_5 inst_cell_58_33 (.BL(BL33),.BLN(BLN33),.WL(WL58));
sram_cell_6t_5 inst_cell_58_34 (.BL(BL34),.BLN(BLN34),.WL(WL58));
sram_cell_6t_5 inst_cell_58_35 (.BL(BL35),.BLN(BLN35),.WL(WL58));
sram_cell_6t_5 inst_cell_58_36 (.BL(BL36),.BLN(BLN36),.WL(WL58));
sram_cell_6t_5 inst_cell_58_37 (.BL(BL37),.BLN(BLN37),.WL(WL58));
sram_cell_6t_5 inst_cell_58_38 (.BL(BL38),.BLN(BLN38),.WL(WL58));
sram_cell_6t_5 inst_cell_58_39 (.BL(BL39),.BLN(BLN39),.WL(WL58));
sram_cell_6t_5 inst_cell_58_40 (.BL(BL40),.BLN(BLN40),.WL(WL58));
sram_cell_6t_5 inst_cell_58_41 (.BL(BL41),.BLN(BLN41),.WL(WL58));
sram_cell_6t_5 inst_cell_58_42 (.BL(BL42),.BLN(BLN42),.WL(WL58));
sram_cell_6t_5 inst_cell_58_43 (.BL(BL43),.BLN(BLN43),.WL(WL58));
sram_cell_6t_5 inst_cell_58_44 (.BL(BL44),.BLN(BLN44),.WL(WL58));
sram_cell_6t_5 inst_cell_58_45 (.BL(BL45),.BLN(BLN45),.WL(WL58));
sram_cell_6t_5 inst_cell_58_46 (.BL(BL46),.BLN(BLN46),.WL(WL58));
sram_cell_6t_5 inst_cell_58_47 (.BL(BL47),.BLN(BLN47),.WL(WL58));
sram_cell_6t_5 inst_cell_58_48 (.BL(BL48),.BLN(BLN48),.WL(WL58));
sram_cell_6t_5 inst_cell_58_49 (.BL(BL49),.BLN(BLN49),.WL(WL58));
sram_cell_6t_5 inst_cell_58_50 (.BL(BL50),.BLN(BLN50),.WL(WL58));
sram_cell_6t_5 inst_cell_58_51 (.BL(BL51),.BLN(BLN51),.WL(WL58));
sram_cell_6t_5 inst_cell_58_52 (.BL(BL52),.BLN(BLN52),.WL(WL58));
sram_cell_6t_5 inst_cell_58_53 (.BL(BL53),.BLN(BLN53),.WL(WL58));
sram_cell_6t_5 inst_cell_58_54 (.BL(BL54),.BLN(BLN54),.WL(WL58));
sram_cell_6t_5 inst_cell_58_55 (.BL(BL55),.BLN(BLN55),.WL(WL58));
sram_cell_6t_5 inst_cell_58_56 (.BL(BL56),.BLN(BLN56),.WL(WL58));
sram_cell_6t_5 inst_cell_58_57 (.BL(BL57),.BLN(BLN57),.WL(WL58));
sram_cell_6t_5 inst_cell_58_58 (.BL(BL58),.BLN(BLN58),.WL(WL58));
sram_cell_6t_5 inst_cell_58_59 (.BL(BL59),.BLN(BLN59),.WL(WL58));
sram_cell_6t_5 inst_cell_58_60 (.BL(BL60),.BLN(BLN60),.WL(WL58));
sram_cell_6t_5 inst_cell_58_61 (.BL(BL61),.BLN(BLN61),.WL(WL58));
sram_cell_6t_5 inst_cell_58_62 (.BL(BL62),.BLN(BLN62),.WL(WL58));
sram_cell_6t_5 inst_cell_58_63 (.BL(BL63),.BLN(BLN63),.WL(WL58));
sram_cell_6t_5 inst_cell_58_64 (.BL(BL64),.BLN(BLN64),.WL(WL58));
sram_cell_6t_5 inst_cell_58_65 (.BL(BL65),.BLN(BLN65),.WL(WL58));
sram_cell_6t_5 inst_cell_58_66 (.BL(BL66),.BLN(BLN66),.WL(WL58));
sram_cell_6t_5 inst_cell_58_67 (.BL(BL67),.BLN(BLN67),.WL(WL58));
sram_cell_6t_5 inst_cell_58_68 (.BL(BL68),.BLN(BLN68),.WL(WL58));
sram_cell_6t_5 inst_cell_58_69 (.BL(BL69),.BLN(BLN69),.WL(WL58));
sram_cell_6t_5 inst_cell_58_70 (.BL(BL70),.BLN(BLN70),.WL(WL58));
sram_cell_6t_5 inst_cell_58_71 (.BL(BL71),.BLN(BLN71),.WL(WL58));
sram_cell_6t_5 inst_cell_58_72 (.BL(BL72),.BLN(BLN72),.WL(WL58));
sram_cell_6t_5 inst_cell_58_73 (.BL(BL73),.BLN(BLN73),.WL(WL58));
sram_cell_6t_5 inst_cell_58_74 (.BL(BL74),.BLN(BLN74),.WL(WL58));
sram_cell_6t_5 inst_cell_58_75 (.BL(BL75),.BLN(BLN75),.WL(WL58));
sram_cell_6t_5 inst_cell_58_76 (.BL(BL76),.BLN(BLN76),.WL(WL58));
sram_cell_6t_5 inst_cell_58_77 (.BL(BL77),.BLN(BLN77),.WL(WL58));
sram_cell_6t_5 inst_cell_58_78 (.BL(BL78),.BLN(BLN78),.WL(WL58));
sram_cell_6t_5 inst_cell_58_79 (.BL(BL79),.BLN(BLN79),.WL(WL58));
sram_cell_6t_5 inst_cell_58_80 (.BL(BL80),.BLN(BLN80),.WL(WL58));
sram_cell_6t_5 inst_cell_58_81 (.BL(BL81),.BLN(BLN81),.WL(WL58));
sram_cell_6t_5 inst_cell_58_82 (.BL(BL82),.BLN(BLN82),.WL(WL58));
sram_cell_6t_5 inst_cell_58_83 (.BL(BL83),.BLN(BLN83),.WL(WL58));
sram_cell_6t_5 inst_cell_58_84 (.BL(BL84),.BLN(BLN84),.WL(WL58));
sram_cell_6t_5 inst_cell_58_85 (.BL(BL85),.BLN(BLN85),.WL(WL58));
sram_cell_6t_5 inst_cell_58_86 (.BL(BL86),.BLN(BLN86),.WL(WL58));
sram_cell_6t_5 inst_cell_58_87 (.BL(BL87),.BLN(BLN87),.WL(WL58));
sram_cell_6t_5 inst_cell_58_88 (.BL(BL88),.BLN(BLN88),.WL(WL58));
sram_cell_6t_5 inst_cell_58_89 (.BL(BL89),.BLN(BLN89),.WL(WL58));
sram_cell_6t_5 inst_cell_58_90 (.BL(BL90),.BLN(BLN90),.WL(WL58));
sram_cell_6t_5 inst_cell_58_91 (.BL(BL91),.BLN(BLN91),.WL(WL58));
sram_cell_6t_5 inst_cell_58_92 (.BL(BL92),.BLN(BLN92),.WL(WL58));
sram_cell_6t_5 inst_cell_58_93 (.BL(BL93),.BLN(BLN93),.WL(WL58));
sram_cell_6t_5 inst_cell_58_94 (.BL(BL94),.BLN(BLN94),.WL(WL58));
sram_cell_6t_5 inst_cell_58_95 (.BL(BL95),.BLN(BLN95),.WL(WL58));
sram_cell_6t_5 inst_cell_58_96 (.BL(BL96),.BLN(BLN96),.WL(WL58));
sram_cell_6t_5 inst_cell_58_97 (.BL(BL97),.BLN(BLN97),.WL(WL58));
sram_cell_6t_5 inst_cell_58_98 (.BL(BL98),.BLN(BLN98),.WL(WL58));
sram_cell_6t_5 inst_cell_58_99 (.BL(BL99),.BLN(BLN99),.WL(WL58));
sram_cell_6t_5 inst_cell_58_100 (.BL(BL100),.BLN(BLN100),.WL(WL58));
sram_cell_6t_5 inst_cell_58_101 (.BL(BL101),.BLN(BLN101),.WL(WL58));
sram_cell_6t_5 inst_cell_58_102 (.BL(BL102),.BLN(BLN102),.WL(WL58));
sram_cell_6t_5 inst_cell_58_103 (.BL(BL103),.BLN(BLN103),.WL(WL58));
sram_cell_6t_5 inst_cell_58_104 (.BL(BL104),.BLN(BLN104),.WL(WL58));
sram_cell_6t_5 inst_cell_58_105 (.BL(BL105),.BLN(BLN105),.WL(WL58));
sram_cell_6t_5 inst_cell_58_106 (.BL(BL106),.BLN(BLN106),.WL(WL58));
sram_cell_6t_5 inst_cell_58_107 (.BL(BL107),.BLN(BLN107),.WL(WL58));
sram_cell_6t_5 inst_cell_58_108 (.BL(BL108),.BLN(BLN108),.WL(WL58));
sram_cell_6t_5 inst_cell_58_109 (.BL(BL109),.BLN(BLN109),.WL(WL58));
sram_cell_6t_5 inst_cell_58_110 (.BL(BL110),.BLN(BLN110),.WL(WL58));
sram_cell_6t_5 inst_cell_58_111 (.BL(BL111),.BLN(BLN111),.WL(WL58));
sram_cell_6t_5 inst_cell_58_112 (.BL(BL112),.BLN(BLN112),.WL(WL58));
sram_cell_6t_5 inst_cell_58_113 (.BL(BL113),.BLN(BLN113),.WL(WL58));
sram_cell_6t_5 inst_cell_58_114 (.BL(BL114),.BLN(BLN114),.WL(WL58));
sram_cell_6t_5 inst_cell_58_115 (.BL(BL115),.BLN(BLN115),.WL(WL58));
sram_cell_6t_5 inst_cell_58_116 (.BL(BL116),.BLN(BLN116),.WL(WL58));
sram_cell_6t_5 inst_cell_58_117 (.BL(BL117),.BLN(BLN117),.WL(WL58));
sram_cell_6t_5 inst_cell_58_118 (.BL(BL118),.BLN(BLN118),.WL(WL58));
sram_cell_6t_5 inst_cell_58_119 (.BL(BL119),.BLN(BLN119),.WL(WL58));
sram_cell_6t_5 inst_cell_58_120 (.BL(BL120),.BLN(BLN120),.WL(WL58));
sram_cell_6t_5 inst_cell_58_121 (.BL(BL121),.BLN(BLN121),.WL(WL58));
sram_cell_6t_5 inst_cell_58_122 (.BL(BL122),.BLN(BLN122),.WL(WL58));
sram_cell_6t_5 inst_cell_58_123 (.BL(BL123),.BLN(BLN123),.WL(WL58));
sram_cell_6t_5 inst_cell_58_124 (.BL(BL124),.BLN(BLN124),.WL(WL58));
sram_cell_6t_5 inst_cell_58_125 (.BL(BL125),.BLN(BLN125),.WL(WL58));
sram_cell_6t_5 inst_cell_58_126 (.BL(BL126),.BLN(BLN126),.WL(WL58));
sram_cell_6t_5 inst_cell_58_127 (.BL(BL127),.BLN(BLN127),.WL(WL58));
sram_cell_6t_5 inst_cell_59_0 (.BL(BL0),.BLN(BLN0),.WL(WL59));
sram_cell_6t_5 inst_cell_59_1 (.BL(BL1),.BLN(BLN1),.WL(WL59));
sram_cell_6t_5 inst_cell_59_2 (.BL(BL2),.BLN(BLN2),.WL(WL59));
sram_cell_6t_5 inst_cell_59_3 (.BL(BL3),.BLN(BLN3),.WL(WL59));
sram_cell_6t_5 inst_cell_59_4 (.BL(BL4),.BLN(BLN4),.WL(WL59));
sram_cell_6t_5 inst_cell_59_5 (.BL(BL5),.BLN(BLN5),.WL(WL59));
sram_cell_6t_5 inst_cell_59_6 (.BL(BL6),.BLN(BLN6),.WL(WL59));
sram_cell_6t_5 inst_cell_59_7 (.BL(BL7),.BLN(BLN7),.WL(WL59));
sram_cell_6t_5 inst_cell_59_8 (.BL(BL8),.BLN(BLN8),.WL(WL59));
sram_cell_6t_5 inst_cell_59_9 (.BL(BL9),.BLN(BLN9),.WL(WL59));
sram_cell_6t_5 inst_cell_59_10 (.BL(BL10),.BLN(BLN10),.WL(WL59));
sram_cell_6t_5 inst_cell_59_11 (.BL(BL11),.BLN(BLN11),.WL(WL59));
sram_cell_6t_5 inst_cell_59_12 (.BL(BL12),.BLN(BLN12),.WL(WL59));
sram_cell_6t_5 inst_cell_59_13 (.BL(BL13),.BLN(BLN13),.WL(WL59));
sram_cell_6t_5 inst_cell_59_14 (.BL(BL14),.BLN(BLN14),.WL(WL59));
sram_cell_6t_5 inst_cell_59_15 (.BL(BL15),.BLN(BLN15),.WL(WL59));
sram_cell_6t_5 inst_cell_59_16 (.BL(BL16),.BLN(BLN16),.WL(WL59));
sram_cell_6t_5 inst_cell_59_17 (.BL(BL17),.BLN(BLN17),.WL(WL59));
sram_cell_6t_5 inst_cell_59_18 (.BL(BL18),.BLN(BLN18),.WL(WL59));
sram_cell_6t_5 inst_cell_59_19 (.BL(BL19),.BLN(BLN19),.WL(WL59));
sram_cell_6t_5 inst_cell_59_20 (.BL(BL20),.BLN(BLN20),.WL(WL59));
sram_cell_6t_5 inst_cell_59_21 (.BL(BL21),.BLN(BLN21),.WL(WL59));
sram_cell_6t_5 inst_cell_59_22 (.BL(BL22),.BLN(BLN22),.WL(WL59));
sram_cell_6t_5 inst_cell_59_23 (.BL(BL23),.BLN(BLN23),.WL(WL59));
sram_cell_6t_5 inst_cell_59_24 (.BL(BL24),.BLN(BLN24),.WL(WL59));
sram_cell_6t_5 inst_cell_59_25 (.BL(BL25),.BLN(BLN25),.WL(WL59));
sram_cell_6t_5 inst_cell_59_26 (.BL(BL26),.BLN(BLN26),.WL(WL59));
sram_cell_6t_5 inst_cell_59_27 (.BL(BL27),.BLN(BLN27),.WL(WL59));
sram_cell_6t_5 inst_cell_59_28 (.BL(BL28),.BLN(BLN28),.WL(WL59));
sram_cell_6t_5 inst_cell_59_29 (.BL(BL29),.BLN(BLN29),.WL(WL59));
sram_cell_6t_5 inst_cell_59_30 (.BL(BL30),.BLN(BLN30),.WL(WL59));
sram_cell_6t_5 inst_cell_59_31 (.BL(BL31),.BLN(BLN31),.WL(WL59));
sram_cell_6t_5 inst_cell_59_32 (.BL(BL32),.BLN(BLN32),.WL(WL59));
sram_cell_6t_5 inst_cell_59_33 (.BL(BL33),.BLN(BLN33),.WL(WL59));
sram_cell_6t_5 inst_cell_59_34 (.BL(BL34),.BLN(BLN34),.WL(WL59));
sram_cell_6t_5 inst_cell_59_35 (.BL(BL35),.BLN(BLN35),.WL(WL59));
sram_cell_6t_5 inst_cell_59_36 (.BL(BL36),.BLN(BLN36),.WL(WL59));
sram_cell_6t_5 inst_cell_59_37 (.BL(BL37),.BLN(BLN37),.WL(WL59));
sram_cell_6t_5 inst_cell_59_38 (.BL(BL38),.BLN(BLN38),.WL(WL59));
sram_cell_6t_5 inst_cell_59_39 (.BL(BL39),.BLN(BLN39),.WL(WL59));
sram_cell_6t_5 inst_cell_59_40 (.BL(BL40),.BLN(BLN40),.WL(WL59));
sram_cell_6t_5 inst_cell_59_41 (.BL(BL41),.BLN(BLN41),.WL(WL59));
sram_cell_6t_5 inst_cell_59_42 (.BL(BL42),.BLN(BLN42),.WL(WL59));
sram_cell_6t_5 inst_cell_59_43 (.BL(BL43),.BLN(BLN43),.WL(WL59));
sram_cell_6t_5 inst_cell_59_44 (.BL(BL44),.BLN(BLN44),.WL(WL59));
sram_cell_6t_5 inst_cell_59_45 (.BL(BL45),.BLN(BLN45),.WL(WL59));
sram_cell_6t_5 inst_cell_59_46 (.BL(BL46),.BLN(BLN46),.WL(WL59));
sram_cell_6t_5 inst_cell_59_47 (.BL(BL47),.BLN(BLN47),.WL(WL59));
sram_cell_6t_5 inst_cell_59_48 (.BL(BL48),.BLN(BLN48),.WL(WL59));
sram_cell_6t_5 inst_cell_59_49 (.BL(BL49),.BLN(BLN49),.WL(WL59));
sram_cell_6t_5 inst_cell_59_50 (.BL(BL50),.BLN(BLN50),.WL(WL59));
sram_cell_6t_5 inst_cell_59_51 (.BL(BL51),.BLN(BLN51),.WL(WL59));
sram_cell_6t_5 inst_cell_59_52 (.BL(BL52),.BLN(BLN52),.WL(WL59));
sram_cell_6t_5 inst_cell_59_53 (.BL(BL53),.BLN(BLN53),.WL(WL59));
sram_cell_6t_5 inst_cell_59_54 (.BL(BL54),.BLN(BLN54),.WL(WL59));
sram_cell_6t_5 inst_cell_59_55 (.BL(BL55),.BLN(BLN55),.WL(WL59));
sram_cell_6t_5 inst_cell_59_56 (.BL(BL56),.BLN(BLN56),.WL(WL59));
sram_cell_6t_5 inst_cell_59_57 (.BL(BL57),.BLN(BLN57),.WL(WL59));
sram_cell_6t_5 inst_cell_59_58 (.BL(BL58),.BLN(BLN58),.WL(WL59));
sram_cell_6t_5 inst_cell_59_59 (.BL(BL59),.BLN(BLN59),.WL(WL59));
sram_cell_6t_5 inst_cell_59_60 (.BL(BL60),.BLN(BLN60),.WL(WL59));
sram_cell_6t_5 inst_cell_59_61 (.BL(BL61),.BLN(BLN61),.WL(WL59));
sram_cell_6t_5 inst_cell_59_62 (.BL(BL62),.BLN(BLN62),.WL(WL59));
sram_cell_6t_5 inst_cell_59_63 (.BL(BL63),.BLN(BLN63),.WL(WL59));
sram_cell_6t_5 inst_cell_59_64 (.BL(BL64),.BLN(BLN64),.WL(WL59));
sram_cell_6t_5 inst_cell_59_65 (.BL(BL65),.BLN(BLN65),.WL(WL59));
sram_cell_6t_5 inst_cell_59_66 (.BL(BL66),.BLN(BLN66),.WL(WL59));
sram_cell_6t_5 inst_cell_59_67 (.BL(BL67),.BLN(BLN67),.WL(WL59));
sram_cell_6t_5 inst_cell_59_68 (.BL(BL68),.BLN(BLN68),.WL(WL59));
sram_cell_6t_5 inst_cell_59_69 (.BL(BL69),.BLN(BLN69),.WL(WL59));
sram_cell_6t_5 inst_cell_59_70 (.BL(BL70),.BLN(BLN70),.WL(WL59));
sram_cell_6t_5 inst_cell_59_71 (.BL(BL71),.BLN(BLN71),.WL(WL59));
sram_cell_6t_5 inst_cell_59_72 (.BL(BL72),.BLN(BLN72),.WL(WL59));
sram_cell_6t_5 inst_cell_59_73 (.BL(BL73),.BLN(BLN73),.WL(WL59));
sram_cell_6t_5 inst_cell_59_74 (.BL(BL74),.BLN(BLN74),.WL(WL59));
sram_cell_6t_5 inst_cell_59_75 (.BL(BL75),.BLN(BLN75),.WL(WL59));
sram_cell_6t_5 inst_cell_59_76 (.BL(BL76),.BLN(BLN76),.WL(WL59));
sram_cell_6t_5 inst_cell_59_77 (.BL(BL77),.BLN(BLN77),.WL(WL59));
sram_cell_6t_5 inst_cell_59_78 (.BL(BL78),.BLN(BLN78),.WL(WL59));
sram_cell_6t_5 inst_cell_59_79 (.BL(BL79),.BLN(BLN79),.WL(WL59));
sram_cell_6t_5 inst_cell_59_80 (.BL(BL80),.BLN(BLN80),.WL(WL59));
sram_cell_6t_5 inst_cell_59_81 (.BL(BL81),.BLN(BLN81),.WL(WL59));
sram_cell_6t_5 inst_cell_59_82 (.BL(BL82),.BLN(BLN82),.WL(WL59));
sram_cell_6t_5 inst_cell_59_83 (.BL(BL83),.BLN(BLN83),.WL(WL59));
sram_cell_6t_5 inst_cell_59_84 (.BL(BL84),.BLN(BLN84),.WL(WL59));
sram_cell_6t_5 inst_cell_59_85 (.BL(BL85),.BLN(BLN85),.WL(WL59));
sram_cell_6t_5 inst_cell_59_86 (.BL(BL86),.BLN(BLN86),.WL(WL59));
sram_cell_6t_5 inst_cell_59_87 (.BL(BL87),.BLN(BLN87),.WL(WL59));
sram_cell_6t_5 inst_cell_59_88 (.BL(BL88),.BLN(BLN88),.WL(WL59));
sram_cell_6t_5 inst_cell_59_89 (.BL(BL89),.BLN(BLN89),.WL(WL59));
sram_cell_6t_5 inst_cell_59_90 (.BL(BL90),.BLN(BLN90),.WL(WL59));
sram_cell_6t_5 inst_cell_59_91 (.BL(BL91),.BLN(BLN91),.WL(WL59));
sram_cell_6t_5 inst_cell_59_92 (.BL(BL92),.BLN(BLN92),.WL(WL59));
sram_cell_6t_5 inst_cell_59_93 (.BL(BL93),.BLN(BLN93),.WL(WL59));
sram_cell_6t_5 inst_cell_59_94 (.BL(BL94),.BLN(BLN94),.WL(WL59));
sram_cell_6t_5 inst_cell_59_95 (.BL(BL95),.BLN(BLN95),.WL(WL59));
sram_cell_6t_5 inst_cell_59_96 (.BL(BL96),.BLN(BLN96),.WL(WL59));
sram_cell_6t_5 inst_cell_59_97 (.BL(BL97),.BLN(BLN97),.WL(WL59));
sram_cell_6t_5 inst_cell_59_98 (.BL(BL98),.BLN(BLN98),.WL(WL59));
sram_cell_6t_5 inst_cell_59_99 (.BL(BL99),.BLN(BLN99),.WL(WL59));
sram_cell_6t_5 inst_cell_59_100 (.BL(BL100),.BLN(BLN100),.WL(WL59));
sram_cell_6t_5 inst_cell_59_101 (.BL(BL101),.BLN(BLN101),.WL(WL59));
sram_cell_6t_5 inst_cell_59_102 (.BL(BL102),.BLN(BLN102),.WL(WL59));
sram_cell_6t_5 inst_cell_59_103 (.BL(BL103),.BLN(BLN103),.WL(WL59));
sram_cell_6t_5 inst_cell_59_104 (.BL(BL104),.BLN(BLN104),.WL(WL59));
sram_cell_6t_5 inst_cell_59_105 (.BL(BL105),.BLN(BLN105),.WL(WL59));
sram_cell_6t_5 inst_cell_59_106 (.BL(BL106),.BLN(BLN106),.WL(WL59));
sram_cell_6t_5 inst_cell_59_107 (.BL(BL107),.BLN(BLN107),.WL(WL59));
sram_cell_6t_5 inst_cell_59_108 (.BL(BL108),.BLN(BLN108),.WL(WL59));
sram_cell_6t_5 inst_cell_59_109 (.BL(BL109),.BLN(BLN109),.WL(WL59));
sram_cell_6t_5 inst_cell_59_110 (.BL(BL110),.BLN(BLN110),.WL(WL59));
sram_cell_6t_5 inst_cell_59_111 (.BL(BL111),.BLN(BLN111),.WL(WL59));
sram_cell_6t_5 inst_cell_59_112 (.BL(BL112),.BLN(BLN112),.WL(WL59));
sram_cell_6t_5 inst_cell_59_113 (.BL(BL113),.BLN(BLN113),.WL(WL59));
sram_cell_6t_5 inst_cell_59_114 (.BL(BL114),.BLN(BLN114),.WL(WL59));
sram_cell_6t_5 inst_cell_59_115 (.BL(BL115),.BLN(BLN115),.WL(WL59));
sram_cell_6t_5 inst_cell_59_116 (.BL(BL116),.BLN(BLN116),.WL(WL59));
sram_cell_6t_5 inst_cell_59_117 (.BL(BL117),.BLN(BLN117),.WL(WL59));
sram_cell_6t_5 inst_cell_59_118 (.BL(BL118),.BLN(BLN118),.WL(WL59));
sram_cell_6t_5 inst_cell_59_119 (.BL(BL119),.BLN(BLN119),.WL(WL59));
sram_cell_6t_5 inst_cell_59_120 (.BL(BL120),.BLN(BLN120),.WL(WL59));
sram_cell_6t_5 inst_cell_59_121 (.BL(BL121),.BLN(BLN121),.WL(WL59));
sram_cell_6t_5 inst_cell_59_122 (.BL(BL122),.BLN(BLN122),.WL(WL59));
sram_cell_6t_5 inst_cell_59_123 (.BL(BL123),.BLN(BLN123),.WL(WL59));
sram_cell_6t_5 inst_cell_59_124 (.BL(BL124),.BLN(BLN124),.WL(WL59));
sram_cell_6t_5 inst_cell_59_125 (.BL(BL125),.BLN(BLN125),.WL(WL59));
sram_cell_6t_5 inst_cell_59_126 (.BL(BL126),.BLN(BLN126),.WL(WL59));
sram_cell_6t_5 inst_cell_59_127 (.BL(BL127),.BLN(BLN127),.WL(WL59));
sram_cell_6t_5 inst_cell_60_0 (.BL(BL0),.BLN(BLN0),.WL(WL60));
sram_cell_6t_5 inst_cell_60_1 (.BL(BL1),.BLN(BLN1),.WL(WL60));
sram_cell_6t_5 inst_cell_60_2 (.BL(BL2),.BLN(BLN2),.WL(WL60));
sram_cell_6t_5 inst_cell_60_3 (.BL(BL3),.BLN(BLN3),.WL(WL60));
sram_cell_6t_5 inst_cell_60_4 (.BL(BL4),.BLN(BLN4),.WL(WL60));
sram_cell_6t_5 inst_cell_60_5 (.BL(BL5),.BLN(BLN5),.WL(WL60));
sram_cell_6t_5 inst_cell_60_6 (.BL(BL6),.BLN(BLN6),.WL(WL60));
sram_cell_6t_5 inst_cell_60_7 (.BL(BL7),.BLN(BLN7),.WL(WL60));
sram_cell_6t_5 inst_cell_60_8 (.BL(BL8),.BLN(BLN8),.WL(WL60));
sram_cell_6t_5 inst_cell_60_9 (.BL(BL9),.BLN(BLN9),.WL(WL60));
sram_cell_6t_5 inst_cell_60_10 (.BL(BL10),.BLN(BLN10),.WL(WL60));
sram_cell_6t_5 inst_cell_60_11 (.BL(BL11),.BLN(BLN11),.WL(WL60));
sram_cell_6t_5 inst_cell_60_12 (.BL(BL12),.BLN(BLN12),.WL(WL60));
sram_cell_6t_5 inst_cell_60_13 (.BL(BL13),.BLN(BLN13),.WL(WL60));
sram_cell_6t_5 inst_cell_60_14 (.BL(BL14),.BLN(BLN14),.WL(WL60));
sram_cell_6t_5 inst_cell_60_15 (.BL(BL15),.BLN(BLN15),.WL(WL60));
sram_cell_6t_5 inst_cell_60_16 (.BL(BL16),.BLN(BLN16),.WL(WL60));
sram_cell_6t_5 inst_cell_60_17 (.BL(BL17),.BLN(BLN17),.WL(WL60));
sram_cell_6t_5 inst_cell_60_18 (.BL(BL18),.BLN(BLN18),.WL(WL60));
sram_cell_6t_5 inst_cell_60_19 (.BL(BL19),.BLN(BLN19),.WL(WL60));
sram_cell_6t_5 inst_cell_60_20 (.BL(BL20),.BLN(BLN20),.WL(WL60));
sram_cell_6t_5 inst_cell_60_21 (.BL(BL21),.BLN(BLN21),.WL(WL60));
sram_cell_6t_5 inst_cell_60_22 (.BL(BL22),.BLN(BLN22),.WL(WL60));
sram_cell_6t_5 inst_cell_60_23 (.BL(BL23),.BLN(BLN23),.WL(WL60));
sram_cell_6t_5 inst_cell_60_24 (.BL(BL24),.BLN(BLN24),.WL(WL60));
sram_cell_6t_5 inst_cell_60_25 (.BL(BL25),.BLN(BLN25),.WL(WL60));
sram_cell_6t_5 inst_cell_60_26 (.BL(BL26),.BLN(BLN26),.WL(WL60));
sram_cell_6t_5 inst_cell_60_27 (.BL(BL27),.BLN(BLN27),.WL(WL60));
sram_cell_6t_5 inst_cell_60_28 (.BL(BL28),.BLN(BLN28),.WL(WL60));
sram_cell_6t_5 inst_cell_60_29 (.BL(BL29),.BLN(BLN29),.WL(WL60));
sram_cell_6t_5 inst_cell_60_30 (.BL(BL30),.BLN(BLN30),.WL(WL60));
sram_cell_6t_5 inst_cell_60_31 (.BL(BL31),.BLN(BLN31),.WL(WL60));
sram_cell_6t_5 inst_cell_60_32 (.BL(BL32),.BLN(BLN32),.WL(WL60));
sram_cell_6t_5 inst_cell_60_33 (.BL(BL33),.BLN(BLN33),.WL(WL60));
sram_cell_6t_5 inst_cell_60_34 (.BL(BL34),.BLN(BLN34),.WL(WL60));
sram_cell_6t_5 inst_cell_60_35 (.BL(BL35),.BLN(BLN35),.WL(WL60));
sram_cell_6t_5 inst_cell_60_36 (.BL(BL36),.BLN(BLN36),.WL(WL60));
sram_cell_6t_5 inst_cell_60_37 (.BL(BL37),.BLN(BLN37),.WL(WL60));
sram_cell_6t_5 inst_cell_60_38 (.BL(BL38),.BLN(BLN38),.WL(WL60));
sram_cell_6t_5 inst_cell_60_39 (.BL(BL39),.BLN(BLN39),.WL(WL60));
sram_cell_6t_5 inst_cell_60_40 (.BL(BL40),.BLN(BLN40),.WL(WL60));
sram_cell_6t_5 inst_cell_60_41 (.BL(BL41),.BLN(BLN41),.WL(WL60));
sram_cell_6t_5 inst_cell_60_42 (.BL(BL42),.BLN(BLN42),.WL(WL60));
sram_cell_6t_5 inst_cell_60_43 (.BL(BL43),.BLN(BLN43),.WL(WL60));
sram_cell_6t_5 inst_cell_60_44 (.BL(BL44),.BLN(BLN44),.WL(WL60));
sram_cell_6t_5 inst_cell_60_45 (.BL(BL45),.BLN(BLN45),.WL(WL60));
sram_cell_6t_5 inst_cell_60_46 (.BL(BL46),.BLN(BLN46),.WL(WL60));
sram_cell_6t_5 inst_cell_60_47 (.BL(BL47),.BLN(BLN47),.WL(WL60));
sram_cell_6t_5 inst_cell_60_48 (.BL(BL48),.BLN(BLN48),.WL(WL60));
sram_cell_6t_5 inst_cell_60_49 (.BL(BL49),.BLN(BLN49),.WL(WL60));
sram_cell_6t_5 inst_cell_60_50 (.BL(BL50),.BLN(BLN50),.WL(WL60));
sram_cell_6t_5 inst_cell_60_51 (.BL(BL51),.BLN(BLN51),.WL(WL60));
sram_cell_6t_5 inst_cell_60_52 (.BL(BL52),.BLN(BLN52),.WL(WL60));
sram_cell_6t_5 inst_cell_60_53 (.BL(BL53),.BLN(BLN53),.WL(WL60));
sram_cell_6t_5 inst_cell_60_54 (.BL(BL54),.BLN(BLN54),.WL(WL60));
sram_cell_6t_5 inst_cell_60_55 (.BL(BL55),.BLN(BLN55),.WL(WL60));
sram_cell_6t_5 inst_cell_60_56 (.BL(BL56),.BLN(BLN56),.WL(WL60));
sram_cell_6t_5 inst_cell_60_57 (.BL(BL57),.BLN(BLN57),.WL(WL60));
sram_cell_6t_5 inst_cell_60_58 (.BL(BL58),.BLN(BLN58),.WL(WL60));
sram_cell_6t_5 inst_cell_60_59 (.BL(BL59),.BLN(BLN59),.WL(WL60));
sram_cell_6t_5 inst_cell_60_60 (.BL(BL60),.BLN(BLN60),.WL(WL60));
sram_cell_6t_5 inst_cell_60_61 (.BL(BL61),.BLN(BLN61),.WL(WL60));
sram_cell_6t_5 inst_cell_60_62 (.BL(BL62),.BLN(BLN62),.WL(WL60));
sram_cell_6t_5 inst_cell_60_63 (.BL(BL63),.BLN(BLN63),.WL(WL60));
sram_cell_6t_5 inst_cell_60_64 (.BL(BL64),.BLN(BLN64),.WL(WL60));
sram_cell_6t_5 inst_cell_60_65 (.BL(BL65),.BLN(BLN65),.WL(WL60));
sram_cell_6t_5 inst_cell_60_66 (.BL(BL66),.BLN(BLN66),.WL(WL60));
sram_cell_6t_5 inst_cell_60_67 (.BL(BL67),.BLN(BLN67),.WL(WL60));
sram_cell_6t_5 inst_cell_60_68 (.BL(BL68),.BLN(BLN68),.WL(WL60));
sram_cell_6t_5 inst_cell_60_69 (.BL(BL69),.BLN(BLN69),.WL(WL60));
sram_cell_6t_5 inst_cell_60_70 (.BL(BL70),.BLN(BLN70),.WL(WL60));
sram_cell_6t_5 inst_cell_60_71 (.BL(BL71),.BLN(BLN71),.WL(WL60));
sram_cell_6t_5 inst_cell_60_72 (.BL(BL72),.BLN(BLN72),.WL(WL60));
sram_cell_6t_5 inst_cell_60_73 (.BL(BL73),.BLN(BLN73),.WL(WL60));
sram_cell_6t_5 inst_cell_60_74 (.BL(BL74),.BLN(BLN74),.WL(WL60));
sram_cell_6t_5 inst_cell_60_75 (.BL(BL75),.BLN(BLN75),.WL(WL60));
sram_cell_6t_5 inst_cell_60_76 (.BL(BL76),.BLN(BLN76),.WL(WL60));
sram_cell_6t_5 inst_cell_60_77 (.BL(BL77),.BLN(BLN77),.WL(WL60));
sram_cell_6t_5 inst_cell_60_78 (.BL(BL78),.BLN(BLN78),.WL(WL60));
sram_cell_6t_5 inst_cell_60_79 (.BL(BL79),.BLN(BLN79),.WL(WL60));
sram_cell_6t_5 inst_cell_60_80 (.BL(BL80),.BLN(BLN80),.WL(WL60));
sram_cell_6t_5 inst_cell_60_81 (.BL(BL81),.BLN(BLN81),.WL(WL60));
sram_cell_6t_5 inst_cell_60_82 (.BL(BL82),.BLN(BLN82),.WL(WL60));
sram_cell_6t_5 inst_cell_60_83 (.BL(BL83),.BLN(BLN83),.WL(WL60));
sram_cell_6t_5 inst_cell_60_84 (.BL(BL84),.BLN(BLN84),.WL(WL60));
sram_cell_6t_5 inst_cell_60_85 (.BL(BL85),.BLN(BLN85),.WL(WL60));
sram_cell_6t_5 inst_cell_60_86 (.BL(BL86),.BLN(BLN86),.WL(WL60));
sram_cell_6t_5 inst_cell_60_87 (.BL(BL87),.BLN(BLN87),.WL(WL60));
sram_cell_6t_5 inst_cell_60_88 (.BL(BL88),.BLN(BLN88),.WL(WL60));
sram_cell_6t_5 inst_cell_60_89 (.BL(BL89),.BLN(BLN89),.WL(WL60));
sram_cell_6t_5 inst_cell_60_90 (.BL(BL90),.BLN(BLN90),.WL(WL60));
sram_cell_6t_5 inst_cell_60_91 (.BL(BL91),.BLN(BLN91),.WL(WL60));
sram_cell_6t_5 inst_cell_60_92 (.BL(BL92),.BLN(BLN92),.WL(WL60));
sram_cell_6t_5 inst_cell_60_93 (.BL(BL93),.BLN(BLN93),.WL(WL60));
sram_cell_6t_5 inst_cell_60_94 (.BL(BL94),.BLN(BLN94),.WL(WL60));
sram_cell_6t_5 inst_cell_60_95 (.BL(BL95),.BLN(BLN95),.WL(WL60));
sram_cell_6t_5 inst_cell_60_96 (.BL(BL96),.BLN(BLN96),.WL(WL60));
sram_cell_6t_5 inst_cell_60_97 (.BL(BL97),.BLN(BLN97),.WL(WL60));
sram_cell_6t_5 inst_cell_60_98 (.BL(BL98),.BLN(BLN98),.WL(WL60));
sram_cell_6t_5 inst_cell_60_99 (.BL(BL99),.BLN(BLN99),.WL(WL60));
sram_cell_6t_5 inst_cell_60_100 (.BL(BL100),.BLN(BLN100),.WL(WL60));
sram_cell_6t_5 inst_cell_60_101 (.BL(BL101),.BLN(BLN101),.WL(WL60));
sram_cell_6t_5 inst_cell_60_102 (.BL(BL102),.BLN(BLN102),.WL(WL60));
sram_cell_6t_5 inst_cell_60_103 (.BL(BL103),.BLN(BLN103),.WL(WL60));
sram_cell_6t_5 inst_cell_60_104 (.BL(BL104),.BLN(BLN104),.WL(WL60));
sram_cell_6t_5 inst_cell_60_105 (.BL(BL105),.BLN(BLN105),.WL(WL60));
sram_cell_6t_5 inst_cell_60_106 (.BL(BL106),.BLN(BLN106),.WL(WL60));
sram_cell_6t_5 inst_cell_60_107 (.BL(BL107),.BLN(BLN107),.WL(WL60));
sram_cell_6t_5 inst_cell_60_108 (.BL(BL108),.BLN(BLN108),.WL(WL60));
sram_cell_6t_5 inst_cell_60_109 (.BL(BL109),.BLN(BLN109),.WL(WL60));
sram_cell_6t_5 inst_cell_60_110 (.BL(BL110),.BLN(BLN110),.WL(WL60));
sram_cell_6t_5 inst_cell_60_111 (.BL(BL111),.BLN(BLN111),.WL(WL60));
sram_cell_6t_5 inst_cell_60_112 (.BL(BL112),.BLN(BLN112),.WL(WL60));
sram_cell_6t_5 inst_cell_60_113 (.BL(BL113),.BLN(BLN113),.WL(WL60));
sram_cell_6t_5 inst_cell_60_114 (.BL(BL114),.BLN(BLN114),.WL(WL60));
sram_cell_6t_5 inst_cell_60_115 (.BL(BL115),.BLN(BLN115),.WL(WL60));
sram_cell_6t_5 inst_cell_60_116 (.BL(BL116),.BLN(BLN116),.WL(WL60));
sram_cell_6t_5 inst_cell_60_117 (.BL(BL117),.BLN(BLN117),.WL(WL60));
sram_cell_6t_5 inst_cell_60_118 (.BL(BL118),.BLN(BLN118),.WL(WL60));
sram_cell_6t_5 inst_cell_60_119 (.BL(BL119),.BLN(BLN119),.WL(WL60));
sram_cell_6t_5 inst_cell_60_120 (.BL(BL120),.BLN(BLN120),.WL(WL60));
sram_cell_6t_5 inst_cell_60_121 (.BL(BL121),.BLN(BLN121),.WL(WL60));
sram_cell_6t_5 inst_cell_60_122 (.BL(BL122),.BLN(BLN122),.WL(WL60));
sram_cell_6t_5 inst_cell_60_123 (.BL(BL123),.BLN(BLN123),.WL(WL60));
sram_cell_6t_5 inst_cell_60_124 (.BL(BL124),.BLN(BLN124),.WL(WL60));
sram_cell_6t_5 inst_cell_60_125 (.BL(BL125),.BLN(BLN125),.WL(WL60));
sram_cell_6t_5 inst_cell_60_126 (.BL(BL126),.BLN(BLN126),.WL(WL60));
sram_cell_6t_5 inst_cell_60_127 (.BL(BL127),.BLN(BLN127),.WL(WL60));
sram_cell_6t_5 inst_cell_61_0 (.BL(BL0),.BLN(BLN0),.WL(WL61));
sram_cell_6t_5 inst_cell_61_1 (.BL(BL1),.BLN(BLN1),.WL(WL61));
sram_cell_6t_5 inst_cell_61_2 (.BL(BL2),.BLN(BLN2),.WL(WL61));
sram_cell_6t_5 inst_cell_61_3 (.BL(BL3),.BLN(BLN3),.WL(WL61));
sram_cell_6t_5 inst_cell_61_4 (.BL(BL4),.BLN(BLN4),.WL(WL61));
sram_cell_6t_5 inst_cell_61_5 (.BL(BL5),.BLN(BLN5),.WL(WL61));
sram_cell_6t_5 inst_cell_61_6 (.BL(BL6),.BLN(BLN6),.WL(WL61));
sram_cell_6t_5 inst_cell_61_7 (.BL(BL7),.BLN(BLN7),.WL(WL61));
sram_cell_6t_5 inst_cell_61_8 (.BL(BL8),.BLN(BLN8),.WL(WL61));
sram_cell_6t_5 inst_cell_61_9 (.BL(BL9),.BLN(BLN9),.WL(WL61));
sram_cell_6t_5 inst_cell_61_10 (.BL(BL10),.BLN(BLN10),.WL(WL61));
sram_cell_6t_5 inst_cell_61_11 (.BL(BL11),.BLN(BLN11),.WL(WL61));
sram_cell_6t_5 inst_cell_61_12 (.BL(BL12),.BLN(BLN12),.WL(WL61));
sram_cell_6t_5 inst_cell_61_13 (.BL(BL13),.BLN(BLN13),.WL(WL61));
sram_cell_6t_5 inst_cell_61_14 (.BL(BL14),.BLN(BLN14),.WL(WL61));
sram_cell_6t_5 inst_cell_61_15 (.BL(BL15),.BLN(BLN15),.WL(WL61));
sram_cell_6t_5 inst_cell_61_16 (.BL(BL16),.BLN(BLN16),.WL(WL61));
sram_cell_6t_5 inst_cell_61_17 (.BL(BL17),.BLN(BLN17),.WL(WL61));
sram_cell_6t_5 inst_cell_61_18 (.BL(BL18),.BLN(BLN18),.WL(WL61));
sram_cell_6t_5 inst_cell_61_19 (.BL(BL19),.BLN(BLN19),.WL(WL61));
sram_cell_6t_5 inst_cell_61_20 (.BL(BL20),.BLN(BLN20),.WL(WL61));
sram_cell_6t_5 inst_cell_61_21 (.BL(BL21),.BLN(BLN21),.WL(WL61));
sram_cell_6t_5 inst_cell_61_22 (.BL(BL22),.BLN(BLN22),.WL(WL61));
sram_cell_6t_5 inst_cell_61_23 (.BL(BL23),.BLN(BLN23),.WL(WL61));
sram_cell_6t_5 inst_cell_61_24 (.BL(BL24),.BLN(BLN24),.WL(WL61));
sram_cell_6t_5 inst_cell_61_25 (.BL(BL25),.BLN(BLN25),.WL(WL61));
sram_cell_6t_5 inst_cell_61_26 (.BL(BL26),.BLN(BLN26),.WL(WL61));
sram_cell_6t_5 inst_cell_61_27 (.BL(BL27),.BLN(BLN27),.WL(WL61));
sram_cell_6t_5 inst_cell_61_28 (.BL(BL28),.BLN(BLN28),.WL(WL61));
sram_cell_6t_5 inst_cell_61_29 (.BL(BL29),.BLN(BLN29),.WL(WL61));
sram_cell_6t_5 inst_cell_61_30 (.BL(BL30),.BLN(BLN30),.WL(WL61));
sram_cell_6t_5 inst_cell_61_31 (.BL(BL31),.BLN(BLN31),.WL(WL61));
sram_cell_6t_5 inst_cell_61_32 (.BL(BL32),.BLN(BLN32),.WL(WL61));
sram_cell_6t_5 inst_cell_61_33 (.BL(BL33),.BLN(BLN33),.WL(WL61));
sram_cell_6t_5 inst_cell_61_34 (.BL(BL34),.BLN(BLN34),.WL(WL61));
sram_cell_6t_5 inst_cell_61_35 (.BL(BL35),.BLN(BLN35),.WL(WL61));
sram_cell_6t_5 inst_cell_61_36 (.BL(BL36),.BLN(BLN36),.WL(WL61));
sram_cell_6t_5 inst_cell_61_37 (.BL(BL37),.BLN(BLN37),.WL(WL61));
sram_cell_6t_5 inst_cell_61_38 (.BL(BL38),.BLN(BLN38),.WL(WL61));
sram_cell_6t_5 inst_cell_61_39 (.BL(BL39),.BLN(BLN39),.WL(WL61));
sram_cell_6t_5 inst_cell_61_40 (.BL(BL40),.BLN(BLN40),.WL(WL61));
sram_cell_6t_5 inst_cell_61_41 (.BL(BL41),.BLN(BLN41),.WL(WL61));
sram_cell_6t_5 inst_cell_61_42 (.BL(BL42),.BLN(BLN42),.WL(WL61));
sram_cell_6t_5 inst_cell_61_43 (.BL(BL43),.BLN(BLN43),.WL(WL61));
sram_cell_6t_5 inst_cell_61_44 (.BL(BL44),.BLN(BLN44),.WL(WL61));
sram_cell_6t_5 inst_cell_61_45 (.BL(BL45),.BLN(BLN45),.WL(WL61));
sram_cell_6t_5 inst_cell_61_46 (.BL(BL46),.BLN(BLN46),.WL(WL61));
sram_cell_6t_5 inst_cell_61_47 (.BL(BL47),.BLN(BLN47),.WL(WL61));
sram_cell_6t_5 inst_cell_61_48 (.BL(BL48),.BLN(BLN48),.WL(WL61));
sram_cell_6t_5 inst_cell_61_49 (.BL(BL49),.BLN(BLN49),.WL(WL61));
sram_cell_6t_5 inst_cell_61_50 (.BL(BL50),.BLN(BLN50),.WL(WL61));
sram_cell_6t_5 inst_cell_61_51 (.BL(BL51),.BLN(BLN51),.WL(WL61));
sram_cell_6t_5 inst_cell_61_52 (.BL(BL52),.BLN(BLN52),.WL(WL61));
sram_cell_6t_5 inst_cell_61_53 (.BL(BL53),.BLN(BLN53),.WL(WL61));
sram_cell_6t_5 inst_cell_61_54 (.BL(BL54),.BLN(BLN54),.WL(WL61));
sram_cell_6t_5 inst_cell_61_55 (.BL(BL55),.BLN(BLN55),.WL(WL61));
sram_cell_6t_5 inst_cell_61_56 (.BL(BL56),.BLN(BLN56),.WL(WL61));
sram_cell_6t_5 inst_cell_61_57 (.BL(BL57),.BLN(BLN57),.WL(WL61));
sram_cell_6t_5 inst_cell_61_58 (.BL(BL58),.BLN(BLN58),.WL(WL61));
sram_cell_6t_5 inst_cell_61_59 (.BL(BL59),.BLN(BLN59),.WL(WL61));
sram_cell_6t_5 inst_cell_61_60 (.BL(BL60),.BLN(BLN60),.WL(WL61));
sram_cell_6t_5 inst_cell_61_61 (.BL(BL61),.BLN(BLN61),.WL(WL61));
sram_cell_6t_5 inst_cell_61_62 (.BL(BL62),.BLN(BLN62),.WL(WL61));
sram_cell_6t_5 inst_cell_61_63 (.BL(BL63),.BLN(BLN63),.WL(WL61));
sram_cell_6t_5 inst_cell_61_64 (.BL(BL64),.BLN(BLN64),.WL(WL61));
sram_cell_6t_5 inst_cell_61_65 (.BL(BL65),.BLN(BLN65),.WL(WL61));
sram_cell_6t_5 inst_cell_61_66 (.BL(BL66),.BLN(BLN66),.WL(WL61));
sram_cell_6t_5 inst_cell_61_67 (.BL(BL67),.BLN(BLN67),.WL(WL61));
sram_cell_6t_5 inst_cell_61_68 (.BL(BL68),.BLN(BLN68),.WL(WL61));
sram_cell_6t_5 inst_cell_61_69 (.BL(BL69),.BLN(BLN69),.WL(WL61));
sram_cell_6t_5 inst_cell_61_70 (.BL(BL70),.BLN(BLN70),.WL(WL61));
sram_cell_6t_5 inst_cell_61_71 (.BL(BL71),.BLN(BLN71),.WL(WL61));
sram_cell_6t_5 inst_cell_61_72 (.BL(BL72),.BLN(BLN72),.WL(WL61));
sram_cell_6t_5 inst_cell_61_73 (.BL(BL73),.BLN(BLN73),.WL(WL61));
sram_cell_6t_5 inst_cell_61_74 (.BL(BL74),.BLN(BLN74),.WL(WL61));
sram_cell_6t_5 inst_cell_61_75 (.BL(BL75),.BLN(BLN75),.WL(WL61));
sram_cell_6t_5 inst_cell_61_76 (.BL(BL76),.BLN(BLN76),.WL(WL61));
sram_cell_6t_5 inst_cell_61_77 (.BL(BL77),.BLN(BLN77),.WL(WL61));
sram_cell_6t_5 inst_cell_61_78 (.BL(BL78),.BLN(BLN78),.WL(WL61));
sram_cell_6t_5 inst_cell_61_79 (.BL(BL79),.BLN(BLN79),.WL(WL61));
sram_cell_6t_5 inst_cell_61_80 (.BL(BL80),.BLN(BLN80),.WL(WL61));
sram_cell_6t_5 inst_cell_61_81 (.BL(BL81),.BLN(BLN81),.WL(WL61));
sram_cell_6t_5 inst_cell_61_82 (.BL(BL82),.BLN(BLN82),.WL(WL61));
sram_cell_6t_5 inst_cell_61_83 (.BL(BL83),.BLN(BLN83),.WL(WL61));
sram_cell_6t_5 inst_cell_61_84 (.BL(BL84),.BLN(BLN84),.WL(WL61));
sram_cell_6t_5 inst_cell_61_85 (.BL(BL85),.BLN(BLN85),.WL(WL61));
sram_cell_6t_5 inst_cell_61_86 (.BL(BL86),.BLN(BLN86),.WL(WL61));
sram_cell_6t_5 inst_cell_61_87 (.BL(BL87),.BLN(BLN87),.WL(WL61));
sram_cell_6t_5 inst_cell_61_88 (.BL(BL88),.BLN(BLN88),.WL(WL61));
sram_cell_6t_5 inst_cell_61_89 (.BL(BL89),.BLN(BLN89),.WL(WL61));
sram_cell_6t_5 inst_cell_61_90 (.BL(BL90),.BLN(BLN90),.WL(WL61));
sram_cell_6t_5 inst_cell_61_91 (.BL(BL91),.BLN(BLN91),.WL(WL61));
sram_cell_6t_5 inst_cell_61_92 (.BL(BL92),.BLN(BLN92),.WL(WL61));
sram_cell_6t_5 inst_cell_61_93 (.BL(BL93),.BLN(BLN93),.WL(WL61));
sram_cell_6t_5 inst_cell_61_94 (.BL(BL94),.BLN(BLN94),.WL(WL61));
sram_cell_6t_5 inst_cell_61_95 (.BL(BL95),.BLN(BLN95),.WL(WL61));
sram_cell_6t_5 inst_cell_61_96 (.BL(BL96),.BLN(BLN96),.WL(WL61));
sram_cell_6t_5 inst_cell_61_97 (.BL(BL97),.BLN(BLN97),.WL(WL61));
sram_cell_6t_5 inst_cell_61_98 (.BL(BL98),.BLN(BLN98),.WL(WL61));
sram_cell_6t_5 inst_cell_61_99 (.BL(BL99),.BLN(BLN99),.WL(WL61));
sram_cell_6t_5 inst_cell_61_100 (.BL(BL100),.BLN(BLN100),.WL(WL61));
sram_cell_6t_5 inst_cell_61_101 (.BL(BL101),.BLN(BLN101),.WL(WL61));
sram_cell_6t_5 inst_cell_61_102 (.BL(BL102),.BLN(BLN102),.WL(WL61));
sram_cell_6t_5 inst_cell_61_103 (.BL(BL103),.BLN(BLN103),.WL(WL61));
sram_cell_6t_5 inst_cell_61_104 (.BL(BL104),.BLN(BLN104),.WL(WL61));
sram_cell_6t_5 inst_cell_61_105 (.BL(BL105),.BLN(BLN105),.WL(WL61));
sram_cell_6t_5 inst_cell_61_106 (.BL(BL106),.BLN(BLN106),.WL(WL61));
sram_cell_6t_5 inst_cell_61_107 (.BL(BL107),.BLN(BLN107),.WL(WL61));
sram_cell_6t_5 inst_cell_61_108 (.BL(BL108),.BLN(BLN108),.WL(WL61));
sram_cell_6t_5 inst_cell_61_109 (.BL(BL109),.BLN(BLN109),.WL(WL61));
sram_cell_6t_5 inst_cell_61_110 (.BL(BL110),.BLN(BLN110),.WL(WL61));
sram_cell_6t_5 inst_cell_61_111 (.BL(BL111),.BLN(BLN111),.WL(WL61));
sram_cell_6t_5 inst_cell_61_112 (.BL(BL112),.BLN(BLN112),.WL(WL61));
sram_cell_6t_5 inst_cell_61_113 (.BL(BL113),.BLN(BLN113),.WL(WL61));
sram_cell_6t_5 inst_cell_61_114 (.BL(BL114),.BLN(BLN114),.WL(WL61));
sram_cell_6t_5 inst_cell_61_115 (.BL(BL115),.BLN(BLN115),.WL(WL61));
sram_cell_6t_5 inst_cell_61_116 (.BL(BL116),.BLN(BLN116),.WL(WL61));
sram_cell_6t_5 inst_cell_61_117 (.BL(BL117),.BLN(BLN117),.WL(WL61));
sram_cell_6t_5 inst_cell_61_118 (.BL(BL118),.BLN(BLN118),.WL(WL61));
sram_cell_6t_5 inst_cell_61_119 (.BL(BL119),.BLN(BLN119),.WL(WL61));
sram_cell_6t_5 inst_cell_61_120 (.BL(BL120),.BLN(BLN120),.WL(WL61));
sram_cell_6t_5 inst_cell_61_121 (.BL(BL121),.BLN(BLN121),.WL(WL61));
sram_cell_6t_5 inst_cell_61_122 (.BL(BL122),.BLN(BLN122),.WL(WL61));
sram_cell_6t_5 inst_cell_61_123 (.BL(BL123),.BLN(BLN123),.WL(WL61));
sram_cell_6t_5 inst_cell_61_124 (.BL(BL124),.BLN(BLN124),.WL(WL61));
sram_cell_6t_5 inst_cell_61_125 (.BL(BL125),.BLN(BLN125),.WL(WL61));
sram_cell_6t_5 inst_cell_61_126 (.BL(BL126),.BLN(BLN126),.WL(WL61));
sram_cell_6t_5 inst_cell_61_127 (.BL(BL127),.BLN(BLN127),.WL(WL61));
sram_cell_6t_5 inst_cell_62_0 (.BL(BL0),.BLN(BLN0),.WL(WL62));
sram_cell_6t_5 inst_cell_62_1 (.BL(BL1),.BLN(BLN1),.WL(WL62));
sram_cell_6t_5 inst_cell_62_2 (.BL(BL2),.BLN(BLN2),.WL(WL62));
sram_cell_6t_5 inst_cell_62_3 (.BL(BL3),.BLN(BLN3),.WL(WL62));
sram_cell_6t_5 inst_cell_62_4 (.BL(BL4),.BLN(BLN4),.WL(WL62));
sram_cell_6t_5 inst_cell_62_5 (.BL(BL5),.BLN(BLN5),.WL(WL62));
sram_cell_6t_5 inst_cell_62_6 (.BL(BL6),.BLN(BLN6),.WL(WL62));
sram_cell_6t_5 inst_cell_62_7 (.BL(BL7),.BLN(BLN7),.WL(WL62));
sram_cell_6t_5 inst_cell_62_8 (.BL(BL8),.BLN(BLN8),.WL(WL62));
sram_cell_6t_5 inst_cell_62_9 (.BL(BL9),.BLN(BLN9),.WL(WL62));
sram_cell_6t_5 inst_cell_62_10 (.BL(BL10),.BLN(BLN10),.WL(WL62));
sram_cell_6t_5 inst_cell_62_11 (.BL(BL11),.BLN(BLN11),.WL(WL62));
sram_cell_6t_5 inst_cell_62_12 (.BL(BL12),.BLN(BLN12),.WL(WL62));
sram_cell_6t_5 inst_cell_62_13 (.BL(BL13),.BLN(BLN13),.WL(WL62));
sram_cell_6t_5 inst_cell_62_14 (.BL(BL14),.BLN(BLN14),.WL(WL62));
sram_cell_6t_5 inst_cell_62_15 (.BL(BL15),.BLN(BLN15),.WL(WL62));
sram_cell_6t_5 inst_cell_62_16 (.BL(BL16),.BLN(BLN16),.WL(WL62));
sram_cell_6t_5 inst_cell_62_17 (.BL(BL17),.BLN(BLN17),.WL(WL62));
sram_cell_6t_5 inst_cell_62_18 (.BL(BL18),.BLN(BLN18),.WL(WL62));
sram_cell_6t_5 inst_cell_62_19 (.BL(BL19),.BLN(BLN19),.WL(WL62));
sram_cell_6t_5 inst_cell_62_20 (.BL(BL20),.BLN(BLN20),.WL(WL62));
sram_cell_6t_5 inst_cell_62_21 (.BL(BL21),.BLN(BLN21),.WL(WL62));
sram_cell_6t_5 inst_cell_62_22 (.BL(BL22),.BLN(BLN22),.WL(WL62));
sram_cell_6t_5 inst_cell_62_23 (.BL(BL23),.BLN(BLN23),.WL(WL62));
sram_cell_6t_5 inst_cell_62_24 (.BL(BL24),.BLN(BLN24),.WL(WL62));
sram_cell_6t_5 inst_cell_62_25 (.BL(BL25),.BLN(BLN25),.WL(WL62));
sram_cell_6t_5 inst_cell_62_26 (.BL(BL26),.BLN(BLN26),.WL(WL62));
sram_cell_6t_5 inst_cell_62_27 (.BL(BL27),.BLN(BLN27),.WL(WL62));
sram_cell_6t_5 inst_cell_62_28 (.BL(BL28),.BLN(BLN28),.WL(WL62));
sram_cell_6t_5 inst_cell_62_29 (.BL(BL29),.BLN(BLN29),.WL(WL62));
sram_cell_6t_5 inst_cell_62_30 (.BL(BL30),.BLN(BLN30),.WL(WL62));
sram_cell_6t_5 inst_cell_62_31 (.BL(BL31),.BLN(BLN31),.WL(WL62));
sram_cell_6t_5 inst_cell_62_32 (.BL(BL32),.BLN(BLN32),.WL(WL62));
sram_cell_6t_5 inst_cell_62_33 (.BL(BL33),.BLN(BLN33),.WL(WL62));
sram_cell_6t_5 inst_cell_62_34 (.BL(BL34),.BLN(BLN34),.WL(WL62));
sram_cell_6t_5 inst_cell_62_35 (.BL(BL35),.BLN(BLN35),.WL(WL62));
sram_cell_6t_5 inst_cell_62_36 (.BL(BL36),.BLN(BLN36),.WL(WL62));
sram_cell_6t_5 inst_cell_62_37 (.BL(BL37),.BLN(BLN37),.WL(WL62));
sram_cell_6t_5 inst_cell_62_38 (.BL(BL38),.BLN(BLN38),.WL(WL62));
sram_cell_6t_5 inst_cell_62_39 (.BL(BL39),.BLN(BLN39),.WL(WL62));
sram_cell_6t_5 inst_cell_62_40 (.BL(BL40),.BLN(BLN40),.WL(WL62));
sram_cell_6t_5 inst_cell_62_41 (.BL(BL41),.BLN(BLN41),.WL(WL62));
sram_cell_6t_5 inst_cell_62_42 (.BL(BL42),.BLN(BLN42),.WL(WL62));
sram_cell_6t_5 inst_cell_62_43 (.BL(BL43),.BLN(BLN43),.WL(WL62));
sram_cell_6t_5 inst_cell_62_44 (.BL(BL44),.BLN(BLN44),.WL(WL62));
sram_cell_6t_5 inst_cell_62_45 (.BL(BL45),.BLN(BLN45),.WL(WL62));
sram_cell_6t_5 inst_cell_62_46 (.BL(BL46),.BLN(BLN46),.WL(WL62));
sram_cell_6t_5 inst_cell_62_47 (.BL(BL47),.BLN(BLN47),.WL(WL62));
sram_cell_6t_5 inst_cell_62_48 (.BL(BL48),.BLN(BLN48),.WL(WL62));
sram_cell_6t_5 inst_cell_62_49 (.BL(BL49),.BLN(BLN49),.WL(WL62));
sram_cell_6t_5 inst_cell_62_50 (.BL(BL50),.BLN(BLN50),.WL(WL62));
sram_cell_6t_5 inst_cell_62_51 (.BL(BL51),.BLN(BLN51),.WL(WL62));
sram_cell_6t_5 inst_cell_62_52 (.BL(BL52),.BLN(BLN52),.WL(WL62));
sram_cell_6t_5 inst_cell_62_53 (.BL(BL53),.BLN(BLN53),.WL(WL62));
sram_cell_6t_5 inst_cell_62_54 (.BL(BL54),.BLN(BLN54),.WL(WL62));
sram_cell_6t_5 inst_cell_62_55 (.BL(BL55),.BLN(BLN55),.WL(WL62));
sram_cell_6t_5 inst_cell_62_56 (.BL(BL56),.BLN(BLN56),.WL(WL62));
sram_cell_6t_5 inst_cell_62_57 (.BL(BL57),.BLN(BLN57),.WL(WL62));
sram_cell_6t_5 inst_cell_62_58 (.BL(BL58),.BLN(BLN58),.WL(WL62));
sram_cell_6t_5 inst_cell_62_59 (.BL(BL59),.BLN(BLN59),.WL(WL62));
sram_cell_6t_5 inst_cell_62_60 (.BL(BL60),.BLN(BLN60),.WL(WL62));
sram_cell_6t_5 inst_cell_62_61 (.BL(BL61),.BLN(BLN61),.WL(WL62));
sram_cell_6t_5 inst_cell_62_62 (.BL(BL62),.BLN(BLN62),.WL(WL62));
sram_cell_6t_5 inst_cell_62_63 (.BL(BL63),.BLN(BLN63),.WL(WL62));
sram_cell_6t_5 inst_cell_62_64 (.BL(BL64),.BLN(BLN64),.WL(WL62));
sram_cell_6t_5 inst_cell_62_65 (.BL(BL65),.BLN(BLN65),.WL(WL62));
sram_cell_6t_5 inst_cell_62_66 (.BL(BL66),.BLN(BLN66),.WL(WL62));
sram_cell_6t_5 inst_cell_62_67 (.BL(BL67),.BLN(BLN67),.WL(WL62));
sram_cell_6t_5 inst_cell_62_68 (.BL(BL68),.BLN(BLN68),.WL(WL62));
sram_cell_6t_5 inst_cell_62_69 (.BL(BL69),.BLN(BLN69),.WL(WL62));
sram_cell_6t_5 inst_cell_62_70 (.BL(BL70),.BLN(BLN70),.WL(WL62));
sram_cell_6t_5 inst_cell_62_71 (.BL(BL71),.BLN(BLN71),.WL(WL62));
sram_cell_6t_5 inst_cell_62_72 (.BL(BL72),.BLN(BLN72),.WL(WL62));
sram_cell_6t_5 inst_cell_62_73 (.BL(BL73),.BLN(BLN73),.WL(WL62));
sram_cell_6t_5 inst_cell_62_74 (.BL(BL74),.BLN(BLN74),.WL(WL62));
sram_cell_6t_5 inst_cell_62_75 (.BL(BL75),.BLN(BLN75),.WL(WL62));
sram_cell_6t_5 inst_cell_62_76 (.BL(BL76),.BLN(BLN76),.WL(WL62));
sram_cell_6t_5 inst_cell_62_77 (.BL(BL77),.BLN(BLN77),.WL(WL62));
sram_cell_6t_5 inst_cell_62_78 (.BL(BL78),.BLN(BLN78),.WL(WL62));
sram_cell_6t_5 inst_cell_62_79 (.BL(BL79),.BLN(BLN79),.WL(WL62));
sram_cell_6t_5 inst_cell_62_80 (.BL(BL80),.BLN(BLN80),.WL(WL62));
sram_cell_6t_5 inst_cell_62_81 (.BL(BL81),.BLN(BLN81),.WL(WL62));
sram_cell_6t_5 inst_cell_62_82 (.BL(BL82),.BLN(BLN82),.WL(WL62));
sram_cell_6t_5 inst_cell_62_83 (.BL(BL83),.BLN(BLN83),.WL(WL62));
sram_cell_6t_5 inst_cell_62_84 (.BL(BL84),.BLN(BLN84),.WL(WL62));
sram_cell_6t_5 inst_cell_62_85 (.BL(BL85),.BLN(BLN85),.WL(WL62));
sram_cell_6t_5 inst_cell_62_86 (.BL(BL86),.BLN(BLN86),.WL(WL62));
sram_cell_6t_5 inst_cell_62_87 (.BL(BL87),.BLN(BLN87),.WL(WL62));
sram_cell_6t_5 inst_cell_62_88 (.BL(BL88),.BLN(BLN88),.WL(WL62));
sram_cell_6t_5 inst_cell_62_89 (.BL(BL89),.BLN(BLN89),.WL(WL62));
sram_cell_6t_5 inst_cell_62_90 (.BL(BL90),.BLN(BLN90),.WL(WL62));
sram_cell_6t_5 inst_cell_62_91 (.BL(BL91),.BLN(BLN91),.WL(WL62));
sram_cell_6t_5 inst_cell_62_92 (.BL(BL92),.BLN(BLN92),.WL(WL62));
sram_cell_6t_5 inst_cell_62_93 (.BL(BL93),.BLN(BLN93),.WL(WL62));
sram_cell_6t_5 inst_cell_62_94 (.BL(BL94),.BLN(BLN94),.WL(WL62));
sram_cell_6t_5 inst_cell_62_95 (.BL(BL95),.BLN(BLN95),.WL(WL62));
sram_cell_6t_5 inst_cell_62_96 (.BL(BL96),.BLN(BLN96),.WL(WL62));
sram_cell_6t_5 inst_cell_62_97 (.BL(BL97),.BLN(BLN97),.WL(WL62));
sram_cell_6t_5 inst_cell_62_98 (.BL(BL98),.BLN(BLN98),.WL(WL62));
sram_cell_6t_5 inst_cell_62_99 (.BL(BL99),.BLN(BLN99),.WL(WL62));
sram_cell_6t_5 inst_cell_62_100 (.BL(BL100),.BLN(BLN100),.WL(WL62));
sram_cell_6t_5 inst_cell_62_101 (.BL(BL101),.BLN(BLN101),.WL(WL62));
sram_cell_6t_5 inst_cell_62_102 (.BL(BL102),.BLN(BLN102),.WL(WL62));
sram_cell_6t_5 inst_cell_62_103 (.BL(BL103),.BLN(BLN103),.WL(WL62));
sram_cell_6t_5 inst_cell_62_104 (.BL(BL104),.BLN(BLN104),.WL(WL62));
sram_cell_6t_5 inst_cell_62_105 (.BL(BL105),.BLN(BLN105),.WL(WL62));
sram_cell_6t_5 inst_cell_62_106 (.BL(BL106),.BLN(BLN106),.WL(WL62));
sram_cell_6t_5 inst_cell_62_107 (.BL(BL107),.BLN(BLN107),.WL(WL62));
sram_cell_6t_5 inst_cell_62_108 (.BL(BL108),.BLN(BLN108),.WL(WL62));
sram_cell_6t_5 inst_cell_62_109 (.BL(BL109),.BLN(BLN109),.WL(WL62));
sram_cell_6t_5 inst_cell_62_110 (.BL(BL110),.BLN(BLN110),.WL(WL62));
sram_cell_6t_5 inst_cell_62_111 (.BL(BL111),.BLN(BLN111),.WL(WL62));
sram_cell_6t_5 inst_cell_62_112 (.BL(BL112),.BLN(BLN112),.WL(WL62));
sram_cell_6t_5 inst_cell_62_113 (.BL(BL113),.BLN(BLN113),.WL(WL62));
sram_cell_6t_5 inst_cell_62_114 (.BL(BL114),.BLN(BLN114),.WL(WL62));
sram_cell_6t_5 inst_cell_62_115 (.BL(BL115),.BLN(BLN115),.WL(WL62));
sram_cell_6t_5 inst_cell_62_116 (.BL(BL116),.BLN(BLN116),.WL(WL62));
sram_cell_6t_5 inst_cell_62_117 (.BL(BL117),.BLN(BLN117),.WL(WL62));
sram_cell_6t_5 inst_cell_62_118 (.BL(BL118),.BLN(BLN118),.WL(WL62));
sram_cell_6t_5 inst_cell_62_119 (.BL(BL119),.BLN(BLN119),.WL(WL62));
sram_cell_6t_5 inst_cell_62_120 (.BL(BL120),.BLN(BLN120),.WL(WL62));
sram_cell_6t_5 inst_cell_62_121 (.BL(BL121),.BLN(BLN121),.WL(WL62));
sram_cell_6t_5 inst_cell_62_122 (.BL(BL122),.BLN(BLN122),.WL(WL62));
sram_cell_6t_5 inst_cell_62_123 (.BL(BL123),.BLN(BLN123),.WL(WL62));
sram_cell_6t_5 inst_cell_62_124 (.BL(BL124),.BLN(BLN124),.WL(WL62));
sram_cell_6t_5 inst_cell_62_125 (.BL(BL125),.BLN(BLN125),.WL(WL62));
sram_cell_6t_5 inst_cell_62_126 (.BL(BL126),.BLN(BLN126),.WL(WL62));
sram_cell_6t_5 inst_cell_62_127 (.BL(BL127),.BLN(BLN127),.WL(WL62));
sram_cell_6t_5 inst_cell_63_0 (.BL(BL0),.BLN(BLN0),.WL(WL63));
sram_cell_6t_5 inst_cell_63_1 (.BL(BL1),.BLN(BLN1),.WL(WL63));
sram_cell_6t_5 inst_cell_63_2 (.BL(BL2),.BLN(BLN2),.WL(WL63));
sram_cell_6t_5 inst_cell_63_3 (.BL(BL3),.BLN(BLN3),.WL(WL63));
sram_cell_6t_5 inst_cell_63_4 (.BL(BL4),.BLN(BLN4),.WL(WL63));
sram_cell_6t_5 inst_cell_63_5 (.BL(BL5),.BLN(BLN5),.WL(WL63));
sram_cell_6t_5 inst_cell_63_6 (.BL(BL6),.BLN(BLN6),.WL(WL63));
sram_cell_6t_5 inst_cell_63_7 (.BL(BL7),.BLN(BLN7),.WL(WL63));
sram_cell_6t_5 inst_cell_63_8 (.BL(BL8),.BLN(BLN8),.WL(WL63));
sram_cell_6t_5 inst_cell_63_9 (.BL(BL9),.BLN(BLN9),.WL(WL63));
sram_cell_6t_5 inst_cell_63_10 (.BL(BL10),.BLN(BLN10),.WL(WL63));
sram_cell_6t_5 inst_cell_63_11 (.BL(BL11),.BLN(BLN11),.WL(WL63));
sram_cell_6t_5 inst_cell_63_12 (.BL(BL12),.BLN(BLN12),.WL(WL63));
sram_cell_6t_5 inst_cell_63_13 (.BL(BL13),.BLN(BLN13),.WL(WL63));
sram_cell_6t_5 inst_cell_63_14 (.BL(BL14),.BLN(BLN14),.WL(WL63));
sram_cell_6t_5 inst_cell_63_15 (.BL(BL15),.BLN(BLN15),.WL(WL63));
sram_cell_6t_5 inst_cell_63_16 (.BL(BL16),.BLN(BLN16),.WL(WL63));
sram_cell_6t_5 inst_cell_63_17 (.BL(BL17),.BLN(BLN17),.WL(WL63));
sram_cell_6t_5 inst_cell_63_18 (.BL(BL18),.BLN(BLN18),.WL(WL63));
sram_cell_6t_5 inst_cell_63_19 (.BL(BL19),.BLN(BLN19),.WL(WL63));
sram_cell_6t_5 inst_cell_63_20 (.BL(BL20),.BLN(BLN20),.WL(WL63));
sram_cell_6t_5 inst_cell_63_21 (.BL(BL21),.BLN(BLN21),.WL(WL63));
sram_cell_6t_5 inst_cell_63_22 (.BL(BL22),.BLN(BLN22),.WL(WL63));
sram_cell_6t_5 inst_cell_63_23 (.BL(BL23),.BLN(BLN23),.WL(WL63));
sram_cell_6t_5 inst_cell_63_24 (.BL(BL24),.BLN(BLN24),.WL(WL63));
sram_cell_6t_5 inst_cell_63_25 (.BL(BL25),.BLN(BLN25),.WL(WL63));
sram_cell_6t_5 inst_cell_63_26 (.BL(BL26),.BLN(BLN26),.WL(WL63));
sram_cell_6t_5 inst_cell_63_27 (.BL(BL27),.BLN(BLN27),.WL(WL63));
sram_cell_6t_5 inst_cell_63_28 (.BL(BL28),.BLN(BLN28),.WL(WL63));
sram_cell_6t_5 inst_cell_63_29 (.BL(BL29),.BLN(BLN29),.WL(WL63));
sram_cell_6t_5 inst_cell_63_30 (.BL(BL30),.BLN(BLN30),.WL(WL63));
sram_cell_6t_5 inst_cell_63_31 (.BL(BL31),.BLN(BLN31),.WL(WL63));
sram_cell_6t_5 inst_cell_63_32 (.BL(BL32),.BLN(BLN32),.WL(WL63));
sram_cell_6t_5 inst_cell_63_33 (.BL(BL33),.BLN(BLN33),.WL(WL63));
sram_cell_6t_5 inst_cell_63_34 (.BL(BL34),.BLN(BLN34),.WL(WL63));
sram_cell_6t_5 inst_cell_63_35 (.BL(BL35),.BLN(BLN35),.WL(WL63));
sram_cell_6t_5 inst_cell_63_36 (.BL(BL36),.BLN(BLN36),.WL(WL63));
sram_cell_6t_5 inst_cell_63_37 (.BL(BL37),.BLN(BLN37),.WL(WL63));
sram_cell_6t_5 inst_cell_63_38 (.BL(BL38),.BLN(BLN38),.WL(WL63));
sram_cell_6t_5 inst_cell_63_39 (.BL(BL39),.BLN(BLN39),.WL(WL63));
sram_cell_6t_5 inst_cell_63_40 (.BL(BL40),.BLN(BLN40),.WL(WL63));
sram_cell_6t_5 inst_cell_63_41 (.BL(BL41),.BLN(BLN41),.WL(WL63));
sram_cell_6t_5 inst_cell_63_42 (.BL(BL42),.BLN(BLN42),.WL(WL63));
sram_cell_6t_5 inst_cell_63_43 (.BL(BL43),.BLN(BLN43),.WL(WL63));
sram_cell_6t_5 inst_cell_63_44 (.BL(BL44),.BLN(BLN44),.WL(WL63));
sram_cell_6t_5 inst_cell_63_45 (.BL(BL45),.BLN(BLN45),.WL(WL63));
sram_cell_6t_5 inst_cell_63_46 (.BL(BL46),.BLN(BLN46),.WL(WL63));
sram_cell_6t_5 inst_cell_63_47 (.BL(BL47),.BLN(BLN47),.WL(WL63));
sram_cell_6t_5 inst_cell_63_48 (.BL(BL48),.BLN(BLN48),.WL(WL63));
sram_cell_6t_5 inst_cell_63_49 (.BL(BL49),.BLN(BLN49),.WL(WL63));
sram_cell_6t_5 inst_cell_63_50 (.BL(BL50),.BLN(BLN50),.WL(WL63));
sram_cell_6t_5 inst_cell_63_51 (.BL(BL51),.BLN(BLN51),.WL(WL63));
sram_cell_6t_5 inst_cell_63_52 (.BL(BL52),.BLN(BLN52),.WL(WL63));
sram_cell_6t_5 inst_cell_63_53 (.BL(BL53),.BLN(BLN53),.WL(WL63));
sram_cell_6t_5 inst_cell_63_54 (.BL(BL54),.BLN(BLN54),.WL(WL63));
sram_cell_6t_5 inst_cell_63_55 (.BL(BL55),.BLN(BLN55),.WL(WL63));
sram_cell_6t_5 inst_cell_63_56 (.BL(BL56),.BLN(BLN56),.WL(WL63));
sram_cell_6t_5 inst_cell_63_57 (.BL(BL57),.BLN(BLN57),.WL(WL63));
sram_cell_6t_5 inst_cell_63_58 (.BL(BL58),.BLN(BLN58),.WL(WL63));
sram_cell_6t_5 inst_cell_63_59 (.BL(BL59),.BLN(BLN59),.WL(WL63));
sram_cell_6t_5 inst_cell_63_60 (.BL(BL60),.BLN(BLN60),.WL(WL63));
sram_cell_6t_5 inst_cell_63_61 (.BL(BL61),.BLN(BLN61),.WL(WL63));
sram_cell_6t_5 inst_cell_63_62 (.BL(BL62),.BLN(BLN62),.WL(WL63));
sram_cell_6t_5 inst_cell_63_63 (.BL(BL63),.BLN(BLN63),.WL(WL63));
sram_cell_6t_5 inst_cell_63_64 (.BL(BL64),.BLN(BLN64),.WL(WL63));
sram_cell_6t_5 inst_cell_63_65 (.BL(BL65),.BLN(BLN65),.WL(WL63));
sram_cell_6t_5 inst_cell_63_66 (.BL(BL66),.BLN(BLN66),.WL(WL63));
sram_cell_6t_5 inst_cell_63_67 (.BL(BL67),.BLN(BLN67),.WL(WL63));
sram_cell_6t_5 inst_cell_63_68 (.BL(BL68),.BLN(BLN68),.WL(WL63));
sram_cell_6t_5 inst_cell_63_69 (.BL(BL69),.BLN(BLN69),.WL(WL63));
sram_cell_6t_5 inst_cell_63_70 (.BL(BL70),.BLN(BLN70),.WL(WL63));
sram_cell_6t_5 inst_cell_63_71 (.BL(BL71),.BLN(BLN71),.WL(WL63));
sram_cell_6t_5 inst_cell_63_72 (.BL(BL72),.BLN(BLN72),.WL(WL63));
sram_cell_6t_5 inst_cell_63_73 (.BL(BL73),.BLN(BLN73),.WL(WL63));
sram_cell_6t_5 inst_cell_63_74 (.BL(BL74),.BLN(BLN74),.WL(WL63));
sram_cell_6t_5 inst_cell_63_75 (.BL(BL75),.BLN(BLN75),.WL(WL63));
sram_cell_6t_5 inst_cell_63_76 (.BL(BL76),.BLN(BLN76),.WL(WL63));
sram_cell_6t_5 inst_cell_63_77 (.BL(BL77),.BLN(BLN77),.WL(WL63));
sram_cell_6t_5 inst_cell_63_78 (.BL(BL78),.BLN(BLN78),.WL(WL63));
sram_cell_6t_5 inst_cell_63_79 (.BL(BL79),.BLN(BLN79),.WL(WL63));
sram_cell_6t_5 inst_cell_63_80 (.BL(BL80),.BLN(BLN80),.WL(WL63));
sram_cell_6t_5 inst_cell_63_81 (.BL(BL81),.BLN(BLN81),.WL(WL63));
sram_cell_6t_5 inst_cell_63_82 (.BL(BL82),.BLN(BLN82),.WL(WL63));
sram_cell_6t_5 inst_cell_63_83 (.BL(BL83),.BLN(BLN83),.WL(WL63));
sram_cell_6t_5 inst_cell_63_84 (.BL(BL84),.BLN(BLN84),.WL(WL63));
sram_cell_6t_5 inst_cell_63_85 (.BL(BL85),.BLN(BLN85),.WL(WL63));
sram_cell_6t_5 inst_cell_63_86 (.BL(BL86),.BLN(BLN86),.WL(WL63));
sram_cell_6t_5 inst_cell_63_87 (.BL(BL87),.BLN(BLN87),.WL(WL63));
sram_cell_6t_5 inst_cell_63_88 (.BL(BL88),.BLN(BLN88),.WL(WL63));
sram_cell_6t_5 inst_cell_63_89 (.BL(BL89),.BLN(BLN89),.WL(WL63));
sram_cell_6t_5 inst_cell_63_90 (.BL(BL90),.BLN(BLN90),.WL(WL63));
sram_cell_6t_5 inst_cell_63_91 (.BL(BL91),.BLN(BLN91),.WL(WL63));
sram_cell_6t_5 inst_cell_63_92 (.BL(BL92),.BLN(BLN92),.WL(WL63));
sram_cell_6t_5 inst_cell_63_93 (.BL(BL93),.BLN(BLN93),.WL(WL63));
sram_cell_6t_5 inst_cell_63_94 (.BL(BL94),.BLN(BLN94),.WL(WL63));
sram_cell_6t_5 inst_cell_63_95 (.BL(BL95),.BLN(BLN95),.WL(WL63));
sram_cell_6t_5 inst_cell_63_96 (.BL(BL96),.BLN(BLN96),.WL(WL63));
sram_cell_6t_5 inst_cell_63_97 (.BL(BL97),.BLN(BLN97),.WL(WL63));
sram_cell_6t_5 inst_cell_63_98 (.BL(BL98),.BLN(BLN98),.WL(WL63));
sram_cell_6t_5 inst_cell_63_99 (.BL(BL99),.BLN(BLN99),.WL(WL63));
sram_cell_6t_5 inst_cell_63_100 (.BL(BL100),.BLN(BLN100),.WL(WL63));
sram_cell_6t_5 inst_cell_63_101 (.BL(BL101),.BLN(BLN101),.WL(WL63));
sram_cell_6t_5 inst_cell_63_102 (.BL(BL102),.BLN(BLN102),.WL(WL63));
sram_cell_6t_5 inst_cell_63_103 (.BL(BL103),.BLN(BLN103),.WL(WL63));
sram_cell_6t_5 inst_cell_63_104 (.BL(BL104),.BLN(BLN104),.WL(WL63));
sram_cell_6t_5 inst_cell_63_105 (.BL(BL105),.BLN(BLN105),.WL(WL63));
sram_cell_6t_5 inst_cell_63_106 (.BL(BL106),.BLN(BLN106),.WL(WL63));
sram_cell_6t_5 inst_cell_63_107 (.BL(BL107),.BLN(BLN107),.WL(WL63));
sram_cell_6t_5 inst_cell_63_108 (.BL(BL108),.BLN(BLN108),.WL(WL63));
sram_cell_6t_5 inst_cell_63_109 (.BL(BL109),.BLN(BLN109),.WL(WL63));
sram_cell_6t_5 inst_cell_63_110 (.BL(BL110),.BLN(BLN110),.WL(WL63));
sram_cell_6t_5 inst_cell_63_111 (.BL(BL111),.BLN(BLN111),.WL(WL63));
sram_cell_6t_5 inst_cell_63_112 (.BL(BL112),.BLN(BLN112),.WL(WL63));
sram_cell_6t_5 inst_cell_63_113 (.BL(BL113),.BLN(BLN113),.WL(WL63));
sram_cell_6t_5 inst_cell_63_114 (.BL(BL114),.BLN(BLN114),.WL(WL63));
sram_cell_6t_5 inst_cell_63_115 (.BL(BL115),.BLN(BLN115),.WL(WL63));
sram_cell_6t_5 inst_cell_63_116 (.BL(BL116),.BLN(BLN116),.WL(WL63));
sram_cell_6t_5 inst_cell_63_117 (.BL(BL117),.BLN(BLN117),.WL(WL63));
sram_cell_6t_5 inst_cell_63_118 (.BL(BL118),.BLN(BLN118),.WL(WL63));
sram_cell_6t_5 inst_cell_63_119 (.BL(BL119),.BLN(BLN119),.WL(WL63));
sram_cell_6t_5 inst_cell_63_120 (.BL(BL120),.BLN(BLN120),.WL(WL63));
sram_cell_6t_5 inst_cell_63_121 (.BL(BL121),.BLN(BLN121),.WL(WL63));
sram_cell_6t_5 inst_cell_63_122 (.BL(BL122),.BLN(BLN122),.WL(WL63));
sram_cell_6t_5 inst_cell_63_123 (.BL(BL123),.BLN(BLN123),.WL(WL63));
sram_cell_6t_5 inst_cell_63_124 (.BL(BL124),.BLN(BLN124),.WL(WL63));
sram_cell_6t_5 inst_cell_63_125 (.BL(BL125),.BLN(BLN125),.WL(WL63));
sram_cell_6t_5 inst_cell_63_126 (.BL(BL126),.BLN(BLN126),.WL(WL63));
sram_cell_6t_5 inst_cell_63_127 (.BL(BL127),.BLN(BLN127),.WL(WL63));
sram_cell_6t_5 inst_cell_64_0 (.BL(BL0),.BLN(BLN0),.WL(WL64));
sram_cell_6t_5 inst_cell_64_1 (.BL(BL1),.BLN(BLN1),.WL(WL64));
sram_cell_6t_5 inst_cell_64_2 (.BL(BL2),.BLN(BLN2),.WL(WL64));
sram_cell_6t_5 inst_cell_64_3 (.BL(BL3),.BLN(BLN3),.WL(WL64));
sram_cell_6t_5 inst_cell_64_4 (.BL(BL4),.BLN(BLN4),.WL(WL64));
sram_cell_6t_5 inst_cell_64_5 (.BL(BL5),.BLN(BLN5),.WL(WL64));
sram_cell_6t_5 inst_cell_64_6 (.BL(BL6),.BLN(BLN6),.WL(WL64));
sram_cell_6t_5 inst_cell_64_7 (.BL(BL7),.BLN(BLN7),.WL(WL64));
sram_cell_6t_5 inst_cell_64_8 (.BL(BL8),.BLN(BLN8),.WL(WL64));
sram_cell_6t_5 inst_cell_64_9 (.BL(BL9),.BLN(BLN9),.WL(WL64));
sram_cell_6t_5 inst_cell_64_10 (.BL(BL10),.BLN(BLN10),.WL(WL64));
sram_cell_6t_5 inst_cell_64_11 (.BL(BL11),.BLN(BLN11),.WL(WL64));
sram_cell_6t_5 inst_cell_64_12 (.BL(BL12),.BLN(BLN12),.WL(WL64));
sram_cell_6t_5 inst_cell_64_13 (.BL(BL13),.BLN(BLN13),.WL(WL64));
sram_cell_6t_5 inst_cell_64_14 (.BL(BL14),.BLN(BLN14),.WL(WL64));
sram_cell_6t_5 inst_cell_64_15 (.BL(BL15),.BLN(BLN15),.WL(WL64));
sram_cell_6t_5 inst_cell_64_16 (.BL(BL16),.BLN(BLN16),.WL(WL64));
sram_cell_6t_5 inst_cell_64_17 (.BL(BL17),.BLN(BLN17),.WL(WL64));
sram_cell_6t_5 inst_cell_64_18 (.BL(BL18),.BLN(BLN18),.WL(WL64));
sram_cell_6t_5 inst_cell_64_19 (.BL(BL19),.BLN(BLN19),.WL(WL64));
sram_cell_6t_5 inst_cell_64_20 (.BL(BL20),.BLN(BLN20),.WL(WL64));
sram_cell_6t_5 inst_cell_64_21 (.BL(BL21),.BLN(BLN21),.WL(WL64));
sram_cell_6t_5 inst_cell_64_22 (.BL(BL22),.BLN(BLN22),.WL(WL64));
sram_cell_6t_5 inst_cell_64_23 (.BL(BL23),.BLN(BLN23),.WL(WL64));
sram_cell_6t_5 inst_cell_64_24 (.BL(BL24),.BLN(BLN24),.WL(WL64));
sram_cell_6t_5 inst_cell_64_25 (.BL(BL25),.BLN(BLN25),.WL(WL64));
sram_cell_6t_5 inst_cell_64_26 (.BL(BL26),.BLN(BLN26),.WL(WL64));
sram_cell_6t_5 inst_cell_64_27 (.BL(BL27),.BLN(BLN27),.WL(WL64));
sram_cell_6t_5 inst_cell_64_28 (.BL(BL28),.BLN(BLN28),.WL(WL64));
sram_cell_6t_5 inst_cell_64_29 (.BL(BL29),.BLN(BLN29),.WL(WL64));
sram_cell_6t_5 inst_cell_64_30 (.BL(BL30),.BLN(BLN30),.WL(WL64));
sram_cell_6t_5 inst_cell_64_31 (.BL(BL31),.BLN(BLN31),.WL(WL64));
sram_cell_6t_5 inst_cell_64_32 (.BL(BL32),.BLN(BLN32),.WL(WL64));
sram_cell_6t_5 inst_cell_64_33 (.BL(BL33),.BLN(BLN33),.WL(WL64));
sram_cell_6t_5 inst_cell_64_34 (.BL(BL34),.BLN(BLN34),.WL(WL64));
sram_cell_6t_5 inst_cell_64_35 (.BL(BL35),.BLN(BLN35),.WL(WL64));
sram_cell_6t_5 inst_cell_64_36 (.BL(BL36),.BLN(BLN36),.WL(WL64));
sram_cell_6t_5 inst_cell_64_37 (.BL(BL37),.BLN(BLN37),.WL(WL64));
sram_cell_6t_5 inst_cell_64_38 (.BL(BL38),.BLN(BLN38),.WL(WL64));
sram_cell_6t_5 inst_cell_64_39 (.BL(BL39),.BLN(BLN39),.WL(WL64));
sram_cell_6t_5 inst_cell_64_40 (.BL(BL40),.BLN(BLN40),.WL(WL64));
sram_cell_6t_5 inst_cell_64_41 (.BL(BL41),.BLN(BLN41),.WL(WL64));
sram_cell_6t_5 inst_cell_64_42 (.BL(BL42),.BLN(BLN42),.WL(WL64));
sram_cell_6t_5 inst_cell_64_43 (.BL(BL43),.BLN(BLN43),.WL(WL64));
sram_cell_6t_5 inst_cell_64_44 (.BL(BL44),.BLN(BLN44),.WL(WL64));
sram_cell_6t_5 inst_cell_64_45 (.BL(BL45),.BLN(BLN45),.WL(WL64));
sram_cell_6t_5 inst_cell_64_46 (.BL(BL46),.BLN(BLN46),.WL(WL64));
sram_cell_6t_5 inst_cell_64_47 (.BL(BL47),.BLN(BLN47),.WL(WL64));
sram_cell_6t_5 inst_cell_64_48 (.BL(BL48),.BLN(BLN48),.WL(WL64));
sram_cell_6t_5 inst_cell_64_49 (.BL(BL49),.BLN(BLN49),.WL(WL64));
sram_cell_6t_5 inst_cell_64_50 (.BL(BL50),.BLN(BLN50),.WL(WL64));
sram_cell_6t_5 inst_cell_64_51 (.BL(BL51),.BLN(BLN51),.WL(WL64));
sram_cell_6t_5 inst_cell_64_52 (.BL(BL52),.BLN(BLN52),.WL(WL64));
sram_cell_6t_5 inst_cell_64_53 (.BL(BL53),.BLN(BLN53),.WL(WL64));
sram_cell_6t_5 inst_cell_64_54 (.BL(BL54),.BLN(BLN54),.WL(WL64));
sram_cell_6t_5 inst_cell_64_55 (.BL(BL55),.BLN(BLN55),.WL(WL64));
sram_cell_6t_5 inst_cell_64_56 (.BL(BL56),.BLN(BLN56),.WL(WL64));
sram_cell_6t_5 inst_cell_64_57 (.BL(BL57),.BLN(BLN57),.WL(WL64));
sram_cell_6t_5 inst_cell_64_58 (.BL(BL58),.BLN(BLN58),.WL(WL64));
sram_cell_6t_5 inst_cell_64_59 (.BL(BL59),.BLN(BLN59),.WL(WL64));
sram_cell_6t_5 inst_cell_64_60 (.BL(BL60),.BLN(BLN60),.WL(WL64));
sram_cell_6t_5 inst_cell_64_61 (.BL(BL61),.BLN(BLN61),.WL(WL64));
sram_cell_6t_5 inst_cell_64_62 (.BL(BL62),.BLN(BLN62),.WL(WL64));
sram_cell_6t_5 inst_cell_64_63 (.BL(BL63),.BLN(BLN63),.WL(WL64));
sram_cell_6t_5 inst_cell_64_64 (.BL(BL64),.BLN(BLN64),.WL(WL64));
sram_cell_6t_5 inst_cell_64_65 (.BL(BL65),.BLN(BLN65),.WL(WL64));
sram_cell_6t_5 inst_cell_64_66 (.BL(BL66),.BLN(BLN66),.WL(WL64));
sram_cell_6t_5 inst_cell_64_67 (.BL(BL67),.BLN(BLN67),.WL(WL64));
sram_cell_6t_5 inst_cell_64_68 (.BL(BL68),.BLN(BLN68),.WL(WL64));
sram_cell_6t_5 inst_cell_64_69 (.BL(BL69),.BLN(BLN69),.WL(WL64));
sram_cell_6t_5 inst_cell_64_70 (.BL(BL70),.BLN(BLN70),.WL(WL64));
sram_cell_6t_5 inst_cell_64_71 (.BL(BL71),.BLN(BLN71),.WL(WL64));
sram_cell_6t_5 inst_cell_64_72 (.BL(BL72),.BLN(BLN72),.WL(WL64));
sram_cell_6t_5 inst_cell_64_73 (.BL(BL73),.BLN(BLN73),.WL(WL64));
sram_cell_6t_5 inst_cell_64_74 (.BL(BL74),.BLN(BLN74),.WL(WL64));
sram_cell_6t_5 inst_cell_64_75 (.BL(BL75),.BLN(BLN75),.WL(WL64));
sram_cell_6t_5 inst_cell_64_76 (.BL(BL76),.BLN(BLN76),.WL(WL64));
sram_cell_6t_5 inst_cell_64_77 (.BL(BL77),.BLN(BLN77),.WL(WL64));
sram_cell_6t_5 inst_cell_64_78 (.BL(BL78),.BLN(BLN78),.WL(WL64));
sram_cell_6t_5 inst_cell_64_79 (.BL(BL79),.BLN(BLN79),.WL(WL64));
sram_cell_6t_5 inst_cell_64_80 (.BL(BL80),.BLN(BLN80),.WL(WL64));
sram_cell_6t_5 inst_cell_64_81 (.BL(BL81),.BLN(BLN81),.WL(WL64));
sram_cell_6t_5 inst_cell_64_82 (.BL(BL82),.BLN(BLN82),.WL(WL64));
sram_cell_6t_5 inst_cell_64_83 (.BL(BL83),.BLN(BLN83),.WL(WL64));
sram_cell_6t_5 inst_cell_64_84 (.BL(BL84),.BLN(BLN84),.WL(WL64));
sram_cell_6t_5 inst_cell_64_85 (.BL(BL85),.BLN(BLN85),.WL(WL64));
sram_cell_6t_5 inst_cell_64_86 (.BL(BL86),.BLN(BLN86),.WL(WL64));
sram_cell_6t_5 inst_cell_64_87 (.BL(BL87),.BLN(BLN87),.WL(WL64));
sram_cell_6t_5 inst_cell_64_88 (.BL(BL88),.BLN(BLN88),.WL(WL64));
sram_cell_6t_5 inst_cell_64_89 (.BL(BL89),.BLN(BLN89),.WL(WL64));
sram_cell_6t_5 inst_cell_64_90 (.BL(BL90),.BLN(BLN90),.WL(WL64));
sram_cell_6t_5 inst_cell_64_91 (.BL(BL91),.BLN(BLN91),.WL(WL64));
sram_cell_6t_5 inst_cell_64_92 (.BL(BL92),.BLN(BLN92),.WL(WL64));
sram_cell_6t_5 inst_cell_64_93 (.BL(BL93),.BLN(BLN93),.WL(WL64));
sram_cell_6t_5 inst_cell_64_94 (.BL(BL94),.BLN(BLN94),.WL(WL64));
sram_cell_6t_5 inst_cell_64_95 (.BL(BL95),.BLN(BLN95),.WL(WL64));
sram_cell_6t_5 inst_cell_64_96 (.BL(BL96),.BLN(BLN96),.WL(WL64));
sram_cell_6t_5 inst_cell_64_97 (.BL(BL97),.BLN(BLN97),.WL(WL64));
sram_cell_6t_5 inst_cell_64_98 (.BL(BL98),.BLN(BLN98),.WL(WL64));
sram_cell_6t_5 inst_cell_64_99 (.BL(BL99),.BLN(BLN99),.WL(WL64));
sram_cell_6t_5 inst_cell_64_100 (.BL(BL100),.BLN(BLN100),.WL(WL64));
sram_cell_6t_5 inst_cell_64_101 (.BL(BL101),.BLN(BLN101),.WL(WL64));
sram_cell_6t_5 inst_cell_64_102 (.BL(BL102),.BLN(BLN102),.WL(WL64));
sram_cell_6t_5 inst_cell_64_103 (.BL(BL103),.BLN(BLN103),.WL(WL64));
sram_cell_6t_5 inst_cell_64_104 (.BL(BL104),.BLN(BLN104),.WL(WL64));
sram_cell_6t_5 inst_cell_64_105 (.BL(BL105),.BLN(BLN105),.WL(WL64));
sram_cell_6t_5 inst_cell_64_106 (.BL(BL106),.BLN(BLN106),.WL(WL64));
sram_cell_6t_5 inst_cell_64_107 (.BL(BL107),.BLN(BLN107),.WL(WL64));
sram_cell_6t_5 inst_cell_64_108 (.BL(BL108),.BLN(BLN108),.WL(WL64));
sram_cell_6t_5 inst_cell_64_109 (.BL(BL109),.BLN(BLN109),.WL(WL64));
sram_cell_6t_5 inst_cell_64_110 (.BL(BL110),.BLN(BLN110),.WL(WL64));
sram_cell_6t_5 inst_cell_64_111 (.BL(BL111),.BLN(BLN111),.WL(WL64));
sram_cell_6t_5 inst_cell_64_112 (.BL(BL112),.BLN(BLN112),.WL(WL64));
sram_cell_6t_5 inst_cell_64_113 (.BL(BL113),.BLN(BLN113),.WL(WL64));
sram_cell_6t_5 inst_cell_64_114 (.BL(BL114),.BLN(BLN114),.WL(WL64));
sram_cell_6t_5 inst_cell_64_115 (.BL(BL115),.BLN(BLN115),.WL(WL64));
sram_cell_6t_5 inst_cell_64_116 (.BL(BL116),.BLN(BLN116),.WL(WL64));
sram_cell_6t_5 inst_cell_64_117 (.BL(BL117),.BLN(BLN117),.WL(WL64));
sram_cell_6t_5 inst_cell_64_118 (.BL(BL118),.BLN(BLN118),.WL(WL64));
sram_cell_6t_5 inst_cell_64_119 (.BL(BL119),.BLN(BLN119),.WL(WL64));
sram_cell_6t_5 inst_cell_64_120 (.BL(BL120),.BLN(BLN120),.WL(WL64));
sram_cell_6t_5 inst_cell_64_121 (.BL(BL121),.BLN(BLN121),.WL(WL64));
sram_cell_6t_5 inst_cell_64_122 (.BL(BL122),.BLN(BLN122),.WL(WL64));
sram_cell_6t_5 inst_cell_64_123 (.BL(BL123),.BLN(BLN123),.WL(WL64));
sram_cell_6t_5 inst_cell_64_124 (.BL(BL124),.BLN(BLN124),.WL(WL64));
sram_cell_6t_5 inst_cell_64_125 (.BL(BL125),.BLN(BLN125),.WL(WL64));
sram_cell_6t_5 inst_cell_64_126 (.BL(BL126),.BLN(BLN126),.WL(WL64));
sram_cell_6t_5 inst_cell_64_127 (.BL(BL127),.BLN(BLN127),.WL(WL64));
sram_cell_6t_5 inst_cell_65_0 (.BL(BL0),.BLN(BLN0),.WL(WL65));
sram_cell_6t_5 inst_cell_65_1 (.BL(BL1),.BLN(BLN1),.WL(WL65));
sram_cell_6t_5 inst_cell_65_2 (.BL(BL2),.BLN(BLN2),.WL(WL65));
sram_cell_6t_5 inst_cell_65_3 (.BL(BL3),.BLN(BLN3),.WL(WL65));
sram_cell_6t_5 inst_cell_65_4 (.BL(BL4),.BLN(BLN4),.WL(WL65));
sram_cell_6t_5 inst_cell_65_5 (.BL(BL5),.BLN(BLN5),.WL(WL65));
sram_cell_6t_5 inst_cell_65_6 (.BL(BL6),.BLN(BLN6),.WL(WL65));
sram_cell_6t_5 inst_cell_65_7 (.BL(BL7),.BLN(BLN7),.WL(WL65));
sram_cell_6t_5 inst_cell_65_8 (.BL(BL8),.BLN(BLN8),.WL(WL65));
sram_cell_6t_5 inst_cell_65_9 (.BL(BL9),.BLN(BLN9),.WL(WL65));
sram_cell_6t_5 inst_cell_65_10 (.BL(BL10),.BLN(BLN10),.WL(WL65));
sram_cell_6t_5 inst_cell_65_11 (.BL(BL11),.BLN(BLN11),.WL(WL65));
sram_cell_6t_5 inst_cell_65_12 (.BL(BL12),.BLN(BLN12),.WL(WL65));
sram_cell_6t_5 inst_cell_65_13 (.BL(BL13),.BLN(BLN13),.WL(WL65));
sram_cell_6t_5 inst_cell_65_14 (.BL(BL14),.BLN(BLN14),.WL(WL65));
sram_cell_6t_5 inst_cell_65_15 (.BL(BL15),.BLN(BLN15),.WL(WL65));
sram_cell_6t_5 inst_cell_65_16 (.BL(BL16),.BLN(BLN16),.WL(WL65));
sram_cell_6t_5 inst_cell_65_17 (.BL(BL17),.BLN(BLN17),.WL(WL65));
sram_cell_6t_5 inst_cell_65_18 (.BL(BL18),.BLN(BLN18),.WL(WL65));
sram_cell_6t_5 inst_cell_65_19 (.BL(BL19),.BLN(BLN19),.WL(WL65));
sram_cell_6t_5 inst_cell_65_20 (.BL(BL20),.BLN(BLN20),.WL(WL65));
sram_cell_6t_5 inst_cell_65_21 (.BL(BL21),.BLN(BLN21),.WL(WL65));
sram_cell_6t_5 inst_cell_65_22 (.BL(BL22),.BLN(BLN22),.WL(WL65));
sram_cell_6t_5 inst_cell_65_23 (.BL(BL23),.BLN(BLN23),.WL(WL65));
sram_cell_6t_5 inst_cell_65_24 (.BL(BL24),.BLN(BLN24),.WL(WL65));
sram_cell_6t_5 inst_cell_65_25 (.BL(BL25),.BLN(BLN25),.WL(WL65));
sram_cell_6t_5 inst_cell_65_26 (.BL(BL26),.BLN(BLN26),.WL(WL65));
sram_cell_6t_5 inst_cell_65_27 (.BL(BL27),.BLN(BLN27),.WL(WL65));
sram_cell_6t_5 inst_cell_65_28 (.BL(BL28),.BLN(BLN28),.WL(WL65));
sram_cell_6t_5 inst_cell_65_29 (.BL(BL29),.BLN(BLN29),.WL(WL65));
sram_cell_6t_5 inst_cell_65_30 (.BL(BL30),.BLN(BLN30),.WL(WL65));
sram_cell_6t_5 inst_cell_65_31 (.BL(BL31),.BLN(BLN31),.WL(WL65));
sram_cell_6t_5 inst_cell_65_32 (.BL(BL32),.BLN(BLN32),.WL(WL65));
sram_cell_6t_5 inst_cell_65_33 (.BL(BL33),.BLN(BLN33),.WL(WL65));
sram_cell_6t_5 inst_cell_65_34 (.BL(BL34),.BLN(BLN34),.WL(WL65));
sram_cell_6t_5 inst_cell_65_35 (.BL(BL35),.BLN(BLN35),.WL(WL65));
sram_cell_6t_5 inst_cell_65_36 (.BL(BL36),.BLN(BLN36),.WL(WL65));
sram_cell_6t_5 inst_cell_65_37 (.BL(BL37),.BLN(BLN37),.WL(WL65));
sram_cell_6t_5 inst_cell_65_38 (.BL(BL38),.BLN(BLN38),.WL(WL65));
sram_cell_6t_5 inst_cell_65_39 (.BL(BL39),.BLN(BLN39),.WL(WL65));
sram_cell_6t_5 inst_cell_65_40 (.BL(BL40),.BLN(BLN40),.WL(WL65));
sram_cell_6t_5 inst_cell_65_41 (.BL(BL41),.BLN(BLN41),.WL(WL65));
sram_cell_6t_5 inst_cell_65_42 (.BL(BL42),.BLN(BLN42),.WL(WL65));
sram_cell_6t_5 inst_cell_65_43 (.BL(BL43),.BLN(BLN43),.WL(WL65));
sram_cell_6t_5 inst_cell_65_44 (.BL(BL44),.BLN(BLN44),.WL(WL65));
sram_cell_6t_5 inst_cell_65_45 (.BL(BL45),.BLN(BLN45),.WL(WL65));
sram_cell_6t_5 inst_cell_65_46 (.BL(BL46),.BLN(BLN46),.WL(WL65));
sram_cell_6t_5 inst_cell_65_47 (.BL(BL47),.BLN(BLN47),.WL(WL65));
sram_cell_6t_5 inst_cell_65_48 (.BL(BL48),.BLN(BLN48),.WL(WL65));
sram_cell_6t_5 inst_cell_65_49 (.BL(BL49),.BLN(BLN49),.WL(WL65));
sram_cell_6t_5 inst_cell_65_50 (.BL(BL50),.BLN(BLN50),.WL(WL65));
sram_cell_6t_5 inst_cell_65_51 (.BL(BL51),.BLN(BLN51),.WL(WL65));
sram_cell_6t_5 inst_cell_65_52 (.BL(BL52),.BLN(BLN52),.WL(WL65));
sram_cell_6t_5 inst_cell_65_53 (.BL(BL53),.BLN(BLN53),.WL(WL65));
sram_cell_6t_5 inst_cell_65_54 (.BL(BL54),.BLN(BLN54),.WL(WL65));
sram_cell_6t_5 inst_cell_65_55 (.BL(BL55),.BLN(BLN55),.WL(WL65));
sram_cell_6t_5 inst_cell_65_56 (.BL(BL56),.BLN(BLN56),.WL(WL65));
sram_cell_6t_5 inst_cell_65_57 (.BL(BL57),.BLN(BLN57),.WL(WL65));
sram_cell_6t_5 inst_cell_65_58 (.BL(BL58),.BLN(BLN58),.WL(WL65));
sram_cell_6t_5 inst_cell_65_59 (.BL(BL59),.BLN(BLN59),.WL(WL65));
sram_cell_6t_5 inst_cell_65_60 (.BL(BL60),.BLN(BLN60),.WL(WL65));
sram_cell_6t_5 inst_cell_65_61 (.BL(BL61),.BLN(BLN61),.WL(WL65));
sram_cell_6t_5 inst_cell_65_62 (.BL(BL62),.BLN(BLN62),.WL(WL65));
sram_cell_6t_5 inst_cell_65_63 (.BL(BL63),.BLN(BLN63),.WL(WL65));
sram_cell_6t_5 inst_cell_65_64 (.BL(BL64),.BLN(BLN64),.WL(WL65));
sram_cell_6t_5 inst_cell_65_65 (.BL(BL65),.BLN(BLN65),.WL(WL65));
sram_cell_6t_5 inst_cell_65_66 (.BL(BL66),.BLN(BLN66),.WL(WL65));
sram_cell_6t_5 inst_cell_65_67 (.BL(BL67),.BLN(BLN67),.WL(WL65));
sram_cell_6t_5 inst_cell_65_68 (.BL(BL68),.BLN(BLN68),.WL(WL65));
sram_cell_6t_5 inst_cell_65_69 (.BL(BL69),.BLN(BLN69),.WL(WL65));
sram_cell_6t_5 inst_cell_65_70 (.BL(BL70),.BLN(BLN70),.WL(WL65));
sram_cell_6t_5 inst_cell_65_71 (.BL(BL71),.BLN(BLN71),.WL(WL65));
sram_cell_6t_5 inst_cell_65_72 (.BL(BL72),.BLN(BLN72),.WL(WL65));
sram_cell_6t_5 inst_cell_65_73 (.BL(BL73),.BLN(BLN73),.WL(WL65));
sram_cell_6t_5 inst_cell_65_74 (.BL(BL74),.BLN(BLN74),.WL(WL65));
sram_cell_6t_5 inst_cell_65_75 (.BL(BL75),.BLN(BLN75),.WL(WL65));
sram_cell_6t_5 inst_cell_65_76 (.BL(BL76),.BLN(BLN76),.WL(WL65));
sram_cell_6t_5 inst_cell_65_77 (.BL(BL77),.BLN(BLN77),.WL(WL65));
sram_cell_6t_5 inst_cell_65_78 (.BL(BL78),.BLN(BLN78),.WL(WL65));
sram_cell_6t_5 inst_cell_65_79 (.BL(BL79),.BLN(BLN79),.WL(WL65));
sram_cell_6t_5 inst_cell_65_80 (.BL(BL80),.BLN(BLN80),.WL(WL65));
sram_cell_6t_5 inst_cell_65_81 (.BL(BL81),.BLN(BLN81),.WL(WL65));
sram_cell_6t_5 inst_cell_65_82 (.BL(BL82),.BLN(BLN82),.WL(WL65));
sram_cell_6t_5 inst_cell_65_83 (.BL(BL83),.BLN(BLN83),.WL(WL65));
sram_cell_6t_5 inst_cell_65_84 (.BL(BL84),.BLN(BLN84),.WL(WL65));
sram_cell_6t_5 inst_cell_65_85 (.BL(BL85),.BLN(BLN85),.WL(WL65));
sram_cell_6t_5 inst_cell_65_86 (.BL(BL86),.BLN(BLN86),.WL(WL65));
sram_cell_6t_5 inst_cell_65_87 (.BL(BL87),.BLN(BLN87),.WL(WL65));
sram_cell_6t_5 inst_cell_65_88 (.BL(BL88),.BLN(BLN88),.WL(WL65));
sram_cell_6t_5 inst_cell_65_89 (.BL(BL89),.BLN(BLN89),.WL(WL65));
sram_cell_6t_5 inst_cell_65_90 (.BL(BL90),.BLN(BLN90),.WL(WL65));
sram_cell_6t_5 inst_cell_65_91 (.BL(BL91),.BLN(BLN91),.WL(WL65));
sram_cell_6t_5 inst_cell_65_92 (.BL(BL92),.BLN(BLN92),.WL(WL65));
sram_cell_6t_5 inst_cell_65_93 (.BL(BL93),.BLN(BLN93),.WL(WL65));
sram_cell_6t_5 inst_cell_65_94 (.BL(BL94),.BLN(BLN94),.WL(WL65));
sram_cell_6t_5 inst_cell_65_95 (.BL(BL95),.BLN(BLN95),.WL(WL65));
sram_cell_6t_5 inst_cell_65_96 (.BL(BL96),.BLN(BLN96),.WL(WL65));
sram_cell_6t_5 inst_cell_65_97 (.BL(BL97),.BLN(BLN97),.WL(WL65));
sram_cell_6t_5 inst_cell_65_98 (.BL(BL98),.BLN(BLN98),.WL(WL65));
sram_cell_6t_5 inst_cell_65_99 (.BL(BL99),.BLN(BLN99),.WL(WL65));
sram_cell_6t_5 inst_cell_65_100 (.BL(BL100),.BLN(BLN100),.WL(WL65));
sram_cell_6t_5 inst_cell_65_101 (.BL(BL101),.BLN(BLN101),.WL(WL65));
sram_cell_6t_5 inst_cell_65_102 (.BL(BL102),.BLN(BLN102),.WL(WL65));
sram_cell_6t_5 inst_cell_65_103 (.BL(BL103),.BLN(BLN103),.WL(WL65));
sram_cell_6t_5 inst_cell_65_104 (.BL(BL104),.BLN(BLN104),.WL(WL65));
sram_cell_6t_5 inst_cell_65_105 (.BL(BL105),.BLN(BLN105),.WL(WL65));
sram_cell_6t_5 inst_cell_65_106 (.BL(BL106),.BLN(BLN106),.WL(WL65));
sram_cell_6t_5 inst_cell_65_107 (.BL(BL107),.BLN(BLN107),.WL(WL65));
sram_cell_6t_5 inst_cell_65_108 (.BL(BL108),.BLN(BLN108),.WL(WL65));
sram_cell_6t_5 inst_cell_65_109 (.BL(BL109),.BLN(BLN109),.WL(WL65));
sram_cell_6t_5 inst_cell_65_110 (.BL(BL110),.BLN(BLN110),.WL(WL65));
sram_cell_6t_5 inst_cell_65_111 (.BL(BL111),.BLN(BLN111),.WL(WL65));
sram_cell_6t_5 inst_cell_65_112 (.BL(BL112),.BLN(BLN112),.WL(WL65));
sram_cell_6t_5 inst_cell_65_113 (.BL(BL113),.BLN(BLN113),.WL(WL65));
sram_cell_6t_5 inst_cell_65_114 (.BL(BL114),.BLN(BLN114),.WL(WL65));
sram_cell_6t_5 inst_cell_65_115 (.BL(BL115),.BLN(BLN115),.WL(WL65));
sram_cell_6t_5 inst_cell_65_116 (.BL(BL116),.BLN(BLN116),.WL(WL65));
sram_cell_6t_5 inst_cell_65_117 (.BL(BL117),.BLN(BLN117),.WL(WL65));
sram_cell_6t_5 inst_cell_65_118 (.BL(BL118),.BLN(BLN118),.WL(WL65));
sram_cell_6t_5 inst_cell_65_119 (.BL(BL119),.BLN(BLN119),.WL(WL65));
sram_cell_6t_5 inst_cell_65_120 (.BL(BL120),.BLN(BLN120),.WL(WL65));
sram_cell_6t_5 inst_cell_65_121 (.BL(BL121),.BLN(BLN121),.WL(WL65));
sram_cell_6t_5 inst_cell_65_122 (.BL(BL122),.BLN(BLN122),.WL(WL65));
sram_cell_6t_5 inst_cell_65_123 (.BL(BL123),.BLN(BLN123),.WL(WL65));
sram_cell_6t_5 inst_cell_65_124 (.BL(BL124),.BLN(BLN124),.WL(WL65));
sram_cell_6t_5 inst_cell_65_125 (.BL(BL125),.BLN(BLN125),.WL(WL65));
sram_cell_6t_5 inst_cell_65_126 (.BL(BL126),.BLN(BLN126),.WL(WL65));
sram_cell_6t_5 inst_cell_65_127 (.BL(BL127),.BLN(BLN127),.WL(WL65));
sram_cell_6t_5 inst_cell_66_0 (.BL(BL0),.BLN(BLN0),.WL(WL66));
sram_cell_6t_5 inst_cell_66_1 (.BL(BL1),.BLN(BLN1),.WL(WL66));
sram_cell_6t_5 inst_cell_66_2 (.BL(BL2),.BLN(BLN2),.WL(WL66));
sram_cell_6t_5 inst_cell_66_3 (.BL(BL3),.BLN(BLN3),.WL(WL66));
sram_cell_6t_5 inst_cell_66_4 (.BL(BL4),.BLN(BLN4),.WL(WL66));
sram_cell_6t_5 inst_cell_66_5 (.BL(BL5),.BLN(BLN5),.WL(WL66));
sram_cell_6t_5 inst_cell_66_6 (.BL(BL6),.BLN(BLN6),.WL(WL66));
sram_cell_6t_5 inst_cell_66_7 (.BL(BL7),.BLN(BLN7),.WL(WL66));
sram_cell_6t_5 inst_cell_66_8 (.BL(BL8),.BLN(BLN8),.WL(WL66));
sram_cell_6t_5 inst_cell_66_9 (.BL(BL9),.BLN(BLN9),.WL(WL66));
sram_cell_6t_5 inst_cell_66_10 (.BL(BL10),.BLN(BLN10),.WL(WL66));
sram_cell_6t_5 inst_cell_66_11 (.BL(BL11),.BLN(BLN11),.WL(WL66));
sram_cell_6t_5 inst_cell_66_12 (.BL(BL12),.BLN(BLN12),.WL(WL66));
sram_cell_6t_5 inst_cell_66_13 (.BL(BL13),.BLN(BLN13),.WL(WL66));
sram_cell_6t_5 inst_cell_66_14 (.BL(BL14),.BLN(BLN14),.WL(WL66));
sram_cell_6t_5 inst_cell_66_15 (.BL(BL15),.BLN(BLN15),.WL(WL66));
sram_cell_6t_5 inst_cell_66_16 (.BL(BL16),.BLN(BLN16),.WL(WL66));
sram_cell_6t_5 inst_cell_66_17 (.BL(BL17),.BLN(BLN17),.WL(WL66));
sram_cell_6t_5 inst_cell_66_18 (.BL(BL18),.BLN(BLN18),.WL(WL66));
sram_cell_6t_5 inst_cell_66_19 (.BL(BL19),.BLN(BLN19),.WL(WL66));
sram_cell_6t_5 inst_cell_66_20 (.BL(BL20),.BLN(BLN20),.WL(WL66));
sram_cell_6t_5 inst_cell_66_21 (.BL(BL21),.BLN(BLN21),.WL(WL66));
sram_cell_6t_5 inst_cell_66_22 (.BL(BL22),.BLN(BLN22),.WL(WL66));
sram_cell_6t_5 inst_cell_66_23 (.BL(BL23),.BLN(BLN23),.WL(WL66));
sram_cell_6t_5 inst_cell_66_24 (.BL(BL24),.BLN(BLN24),.WL(WL66));
sram_cell_6t_5 inst_cell_66_25 (.BL(BL25),.BLN(BLN25),.WL(WL66));
sram_cell_6t_5 inst_cell_66_26 (.BL(BL26),.BLN(BLN26),.WL(WL66));
sram_cell_6t_5 inst_cell_66_27 (.BL(BL27),.BLN(BLN27),.WL(WL66));
sram_cell_6t_5 inst_cell_66_28 (.BL(BL28),.BLN(BLN28),.WL(WL66));
sram_cell_6t_5 inst_cell_66_29 (.BL(BL29),.BLN(BLN29),.WL(WL66));
sram_cell_6t_5 inst_cell_66_30 (.BL(BL30),.BLN(BLN30),.WL(WL66));
sram_cell_6t_5 inst_cell_66_31 (.BL(BL31),.BLN(BLN31),.WL(WL66));
sram_cell_6t_5 inst_cell_66_32 (.BL(BL32),.BLN(BLN32),.WL(WL66));
sram_cell_6t_5 inst_cell_66_33 (.BL(BL33),.BLN(BLN33),.WL(WL66));
sram_cell_6t_5 inst_cell_66_34 (.BL(BL34),.BLN(BLN34),.WL(WL66));
sram_cell_6t_5 inst_cell_66_35 (.BL(BL35),.BLN(BLN35),.WL(WL66));
sram_cell_6t_5 inst_cell_66_36 (.BL(BL36),.BLN(BLN36),.WL(WL66));
sram_cell_6t_5 inst_cell_66_37 (.BL(BL37),.BLN(BLN37),.WL(WL66));
sram_cell_6t_5 inst_cell_66_38 (.BL(BL38),.BLN(BLN38),.WL(WL66));
sram_cell_6t_5 inst_cell_66_39 (.BL(BL39),.BLN(BLN39),.WL(WL66));
sram_cell_6t_5 inst_cell_66_40 (.BL(BL40),.BLN(BLN40),.WL(WL66));
sram_cell_6t_5 inst_cell_66_41 (.BL(BL41),.BLN(BLN41),.WL(WL66));
sram_cell_6t_5 inst_cell_66_42 (.BL(BL42),.BLN(BLN42),.WL(WL66));
sram_cell_6t_5 inst_cell_66_43 (.BL(BL43),.BLN(BLN43),.WL(WL66));
sram_cell_6t_5 inst_cell_66_44 (.BL(BL44),.BLN(BLN44),.WL(WL66));
sram_cell_6t_5 inst_cell_66_45 (.BL(BL45),.BLN(BLN45),.WL(WL66));
sram_cell_6t_5 inst_cell_66_46 (.BL(BL46),.BLN(BLN46),.WL(WL66));
sram_cell_6t_5 inst_cell_66_47 (.BL(BL47),.BLN(BLN47),.WL(WL66));
sram_cell_6t_5 inst_cell_66_48 (.BL(BL48),.BLN(BLN48),.WL(WL66));
sram_cell_6t_5 inst_cell_66_49 (.BL(BL49),.BLN(BLN49),.WL(WL66));
sram_cell_6t_5 inst_cell_66_50 (.BL(BL50),.BLN(BLN50),.WL(WL66));
sram_cell_6t_5 inst_cell_66_51 (.BL(BL51),.BLN(BLN51),.WL(WL66));
sram_cell_6t_5 inst_cell_66_52 (.BL(BL52),.BLN(BLN52),.WL(WL66));
sram_cell_6t_5 inst_cell_66_53 (.BL(BL53),.BLN(BLN53),.WL(WL66));
sram_cell_6t_5 inst_cell_66_54 (.BL(BL54),.BLN(BLN54),.WL(WL66));
sram_cell_6t_5 inst_cell_66_55 (.BL(BL55),.BLN(BLN55),.WL(WL66));
sram_cell_6t_5 inst_cell_66_56 (.BL(BL56),.BLN(BLN56),.WL(WL66));
sram_cell_6t_5 inst_cell_66_57 (.BL(BL57),.BLN(BLN57),.WL(WL66));
sram_cell_6t_5 inst_cell_66_58 (.BL(BL58),.BLN(BLN58),.WL(WL66));
sram_cell_6t_5 inst_cell_66_59 (.BL(BL59),.BLN(BLN59),.WL(WL66));
sram_cell_6t_5 inst_cell_66_60 (.BL(BL60),.BLN(BLN60),.WL(WL66));
sram_cell_6t_5 inst_cell_66_61 (.BL(BL61),.BLN(BLN61),.WL(WL66));
sram_cell_6t_5 inst_cell_66_62 (.BL(BL62),.BLN(BLN62),.WL(WL66));
sram_cell_6t_5 inst_cell_66_63 (.BL(BL63),.BLN(BLN63),.WL(WL66));
sram_cell_6t_5 inst_cell_66_64 (.BL(BL64),.BLN(BLN64),.WL(WL66));
sram_cell_6t_5 inst_cell_66_65 (.BL(BL65),.BLN(BLN65),.WL(WL66));
sram_cell_6t_5 inst_cell_66_66 (.BL(BL66),.BLN(BLN66),.WL(WL66));
sram_cell_6t_5 inst_cell_66_67 (.BL(BL67),.BLN(BLN67),.WL(WL66));
sram_cell_6t_5 inst_cell_66_68 (.BL(BL68),.BLN(BLN68),.WL(WL66));
sram_cell_6t_5 inst_cell_66_69 (.BL(BL69),.BLN(BLN69),.WL(WL66));
sram_cell_6t_5 inst_cell_66_70 (.BL(BL70),.BLN(BLN70),.WL(WL66));
sram_cell_6t_5 inst_cell_66_71 (.BL(BL71),.BLN(BLN71),.WL(WL66));
sram_cell_6t_5 inst_cell_66_72 (.BL(BL72),.BLN(BLN72),.WL(WL66));
sram_cell_6t_5 inst_cell_66_73 (.BL(BL73),.BLN(BLN73),.WL(WL66));
sram_cell_6t_5 inst_cell_66_74 (.BL(BL74),.BLN(BLN74),.WL(WL66));
sram_cell_6t_5 inst_cell_66_75 (.BL(BL75),.BLN(BLN75),.WL(WL66));
sram_cell_6t_5 inst_cell_66_76 (.BL(BL76),.BLN(BLN76),.WL(WL66));
sram_cell_6t_5 inst_cell_66_77 (.BL(BL77),.BLN(BLN77),.WL(WL66));
sram_cell_6t_5 inst_cell_66_78 (.BL(BL78),.BLN(BLN78),.WL(WL66));
sram_cell_6t_5 inst_cell_66_79 (.BL(BL79),.BLN(BLN79),.WL(WL66));
sram_cell_6t_5 inst_cell_66_80 (.BL(BL80),.BLN(BLN80),.WL(WL66));
sram_cell_6t_5 inst_cell_66_81 (.BL(BL81),.BLN(BLN81),.WL(WL66));
sram_cell_6t_5 inst_cell_66_82 (.BL(BL82),.BLN(BLN82),.WL(WL66));
sram_cell_6t_5 inst_cell_66_83 (.BL(BL83),.BLN(BLN83),.WL(WL66));
sram_cell_6t_5 inst_cell_66_84 (.BL(BL84),.BLN(BLN84),.WL(WL66));
sram_cell_6t_5 inst_cell_66_85 (.BL(BL85),.BLN(BLN85),.WL(WL66));
sram_cell_6t_5 inst_cell_66_86 (.BL(BL86),.BLN(BLN86),.WL(WL66));
sram_cell_6t_5 inst_cell_66_87 (.BL(BL87),.BLN(BLN87),.WL(WL66));
sram_cell_6t_5 inst_cell_66_88 (.BL(BL88),.BLN(BLN88),.WL(WL66));
sram_cell_6t_5 inst_cell_66_89 (.BL(BL89),.BLN(BLN89),.WL(WL66));
sram_cell_6t_5 inst_cell_66_90 (.BL(BL90),.BLN(BLN90),.WL(WL66));
sram_cell_6t_5 inst_cell_66_91 (.BL(BL91),.BLN(BLN91),.WL(WL66));
sram_cell_6t_5 inst_cell_66_92 (.BL(BL92),.BLN(BLN92),.WL(WL66));
sram_cell_6t_5 inst_cell_66_93 (.BL(BL93),.BLN(BLN93),.WL(WL66));
sram_cell_6t_5 inst_cell_66_94 (.BL(BL94),.BLN(BLN94),.WL(WL66));
sram_cell_6t_5 inst_cell_66_95 (.BL(BL95),.BLN(BLN95),.WL(WL66));
sram_cell_6t_5 inst_cell_66_96 (.BL(BL96),.BLN(BLN96),.WL(WL66));
sram_cell_6t_5 inst_cell_66_97 (.BL(BL97),.BLN(BLN97),.WL(WL66));
sram_cell_6t_5 inst_cell_66_98 (.BL(BL98),.BLN(BLN98),.WL(WL66));
sram_cell_6t_5 inst_cell_66_99 (.BL(BL99),.BLN(BLN99),.WL(WL66));
sram_cell_6t_5 inst_cell_66_100 (.BL(BL100),.BLN(BLN100),.WL(WL66));
sram_cell_6t_5 inst_cell_66_101 (.BL(BL101),.BLN(BLN101),.WL(WL66));
sram_cell_6t_5 inst_cell_66_102 (.BL(BL102),.BLN(BLN102),.WL(WL66));
sram_cell_6t_5 inst_cell_66_103 (.BL(BL103),.BLN(BLN103),.WL(WL66));
sram_cell_6t_5 inst_cell_66_104 (.BL(BL104),.BLN(BLN104),.WL(WL66));
sram_cell_6t_5 inst_cell_66_105 (.BL(BL105),.BLN(BLN105),.WL(WL66));
sram_cell_6t_5 inst_cell_66_106 (.BL(BL106),.BLN(BLN106),.WL(WL66));
sram_cell_6t_5 inst_cell_66_107 (.BL(BL107),.BLN(BLN107),.WL(WL66));
sram_cell_6t_5 inst_cell_66_108 (.BL(BL108),.BLN(BLN108),.WL(WL66));
sram_cell_6t_5 inst_cell_66_109 (.BL(BL109),.BLN(BLN109),.WL(WL66));
sram_cell_6t_5 inst_cell_66_110 (.BL(BL110),.BLN(BLN110),.WL(WL66));
sram_cell_6t_5 inst_cell_66_111 (.BL(BL111),.BLN(BLN111),.WL(WL66));
sram_cell_6t_5 inst_cell_66_112 (.BL(BL112),.BLN(BLN112),.WL(WL66));
sram_cell_6t_5 inst_cell_66_113 (.BL(BL113),.BLN(BLN113),.WL(WL66));
sram_cell_6t_5 inst_cell_66_114 (.BL(BL114),.BLN(BLN114),.WL(WL66));
sram_cell_6t_5 inst_cell_66_115 (.BL(BL115),.BLN(BLN115),.WL(WL66));
sram_cell_6t_5 inst_cell_66_116 (.BL(BL116),.BLN(BLN116),.WL(WL66));
sram_cell_6t_5 inst_cell_66_117 (.BL(BL117),.BLN(BLN117),.WL(WL66));
sram_cell_6t_5 inst_cell_66_118 (.BL(BL118),.BLN(BLN118),.WL(WL66));
sram_cell_6t_5 inst_cell_66_119 (.BL(BL119),.BLN(BLN119),.WL(WL66));
sram_cell_6t_5 inst_cell_66_120 (.BL(BL120),.BLN(BLN120),.WL(WL66));
sram_cell_6t_5 inst_cell_66_121 (.BL(BL121),.BLN(BLN121),.WL(WL66));
sram_cell_6t_5 inst_cell_66_122 (.BL(BL122),.BLN(BLN122),.WL(WL66));
sram_cell_6t_5 inst_cell_66_123 (.BL(BL123),.BLN(BLN123),.WL(WL66));
sram_cell_6t_5 inst_cell_66_124 (.BL(BL124),.BLN(BLN124),.WL(WL66));
sram_cell_6t_5 inst_cell_66_125 (.BL(BL125),.BLN(BLN125),.WL(WL66));
sram_cell_6t_5 inst_cell_66_126 (.BL(BL126),.BLN(BLN126),.WL(WL66));
sram_cell_6t_5 inst_cell_66_127 (.BL(BL127),.BLN(BLN127),.WL(WL66));
sram_cell_6t_5 inst_cell_67_0 (.BL(BL0),.BLN(BLN0),.WL(WL67));
sram_cell_6t_5 inst_cell_67_1 (.BL(BL1),.BLN(BLN1),.WL(WL67));
sram_cell_6t_5 inst_cell_67_2 (.BL(BL2),.BLN(BLN2),.WL(WL67));
sram_cell_6t_5 inst_cell_67_3 (.BL(BL3),.BLN(BLN3),.WL(WL67));
sram_cell_6t_5 inst_cell_67_4 (.BL(BL4),.BLN(BLN4),.WL(WL67));
sram_cell_6t_5 inst_cell_67_5 (.BL(BL5),.BLN(BLN5),.WL(WL67));
sram_cell_6t_5 inst_cell_67_6 (.BL(BL6),.BLN(BLN6),.WL(WL67));
sram_cell_6t_5 inst_cell_67_7 (.BL(BL7),.BLN(BLN7),.WL(WL67));
sram_cell_6t_5 inst_cell_67_8 (.BL(BL8),.BLN(BLN8),.WL(WL67));
sram_cell_6t_5 inst_cell_67_9 (.BL(BL9),.BLN(BLN9),.WL(WL67));
sram_cell_6t_5 inst_cell_67_10 (.BL(BL10),.BLN(BLN10),.WL(WL67));
sram_cell_6t_5 inst_cell_67_11 (.BL(BL11),.BLN(BLN11),.WL(WL67));
sram_cell_6t_5 inst_cell_67_12 (.BL(BL12),.BLN(BLN12),.WL(WL67));
sram_cell_6t_5 inst_cell_67_13 (.BL(BL13),.BLN(BLN13),.WL(WL67));
sram_cell_6t_5 inst_cell_67_14 (.BL(BL14),.BLN(BLN14),.WL(WL67));
sram_cell_6t_5 inst_cell_67_15 (.BL(BL15),.BLN(BLN15),.WL(WL67));
sram_cell_6t_5 inst_cell_67_16 (.BL(BL16),.BLN(BLN16),.WL(WL67));
sram_cell_6t_5 inst_cell_67_17 (.BL(BL17),.BLN(BLN17),.WL(WL67));
sram_cell_6t_5 inst_cell_67_18 (.BL(BL18),.BLN(BLN18),.WL(WL67));
sram_cell_6t_5 inst_cell_67_19 (.BL(BL19),.BLN(BLN19),.WL(WL67));
sram_cell_6t_5 inst_cell_67_20 (.BL(BL20),.BLN(BLN20),.WL(WL67));
sram_cell_6t_5 inst_cell_67_21 (.BL(BL21),.BLN(BLN21),.WL(WL67));
sram_cell_6t_5 inst_cell_67_22 (.BL(BL22),.BLN(BLN22),.WL(WL67));
sram_cell_6t_5 inst_cell_67_23 (.BL(BL23),.BLN(BLN23),.WL(WL67));
sram_cell_6t_5 inst_cell_67_24 (.BL(BL24),.BLN(BLN24),.WL(WL67));
sram_cell_6t_5 inst_cell_67_25 (.BL(BL25),.BLN(BLN25),.WL(WL67));
sram_cell_6t_5 inst_cell_67_26 (.BL(BL26),.BLN(BLN26),.WL(WL67));
sram_cell_6t_5 inst_cell_67_27 (.BL(BL27),.BLN(BLN27),.WL(WL67));
sram_cell_6t_5 inst_cell_67_28 (.BL(BL28),.BLN(BLN28),.WL(WL67));
sram_cell_6t_5 inst_cell_67_29 (.BL(BL29),.BLN(BLN29),.WL(WL67));
sram_cell_6t_5 inst_cell_67_30 (.BL(BL30),.BLN(BLN30),.WL(WL67));
sram_cell_6t_5 inst_cell_67_31 (.BL(BL31),.BLN(BLN31),.WL(WL67));
sram_cell_6t_5 inst_cell_67_32 (.BL(BL32),.BLN(BLN32),.WL(WL67));
sram_cell_6t_5 inst_cell_67_33 (.BL(BL33),.BLN(BLN33),.WL(WL67));
sram_cell_6t_5 inst_cell_67_34 (.BL(BL34),.BLN(BLN34),.WL(WL67));
sram_cell_6t_5 inst_cell_67_35 (.BL(BL35),.BLN(BLN35),.WL(WL67));
sram_cell_6t_5 inst_cell_67_36 (.BL(BL36),.BLN(BLN36),.WL(WL67));
sram_cell_6t_5 inst_cell_67_37 (.BL(BL37),.BLN(BLN37),.WL(WL67));
sram_cell_6t_5 inst_cell_67_38 (.BL(BL38),.BLN(BLN38),.WL(WL67));
sram_cell_6t_5 inst_cell_67_39 (.BL(BL39),.BLN(BLN39),.WL(WL67));
sram_cell_6t_5 inst_cell_67_40 (.BL(BL40),.BLN(BLN40),.WL(WL67));
sram_cell_6t_5 inst_cell_67_41 (.BL(BL41),.BLN(BLN41),.WL(WL67));
sram_cell_6t_5 inst_cell_67_42 (.BL(BL42),.BLN(BLN42),.WL(WL67));
sram_cell_6t_5 inst_cell_67_43 (.BL(BL43),.BLN(BLN43),.WL(WL67));
sram_cell_6t_5 inst_cell_67_44 (.BL(BL44),.BLN(BLN44),.WL(WL67));
sram_cell_6t_5 inst_cell_67_45 (.BL(BL45),.BLN(BLN45),.WL(WL67));
sram_cell_6t_5 inst_cell_67_46 (.BL(BL46),.BLN(BLN46),.WL(WL67));
sram_cell_6t_5 inst_cell_67_47 (.BL(BL47),.BLN(BLN47),.WL(WL67));
sram_cell_6t_5 inst_cell_67_48 (.BL(BL48),.BLN(BLN48),.WL(WL67));
sram_cell_6t_5 inst_cell_67_49 (.BL(BL49),.BLN(BLN49),.WL(WL67));
sram_cell_6t_5 inst_cell_67_50 (.BL(BL50),.BLN(BLN50),.WL(WL67));
sram_cell_6t_5 inst_cell_67_51 (.BL(BL51),.BLN(BLN51),.WL(WL67));
sram_cell_6t_5 inst_cell_67_52 (.BL(BL52),.BLN(BLN52),.WL(WL67));
sram_cell_6t_5 inst_cell_67_53 (.BL(BL53),.BLN(BLN53),.WL(WL67));
sram_cell_6t_5 inst_cell_67_54 (.BL(BL54),.BLN(BLN54),.WL(WL67));
sram_cell_6t_5 inst_cell_67_55 (.BL(BL55),.BLN(BLN55),.WL(WL67));
sram_cell_6t_5 inst_cell_67_56 (.BL(BL56),.BLN(BLN56),.WL(WL67));
sram_cell_6t_5 inst_cell_67_57 (.BL(BL57),.BLN(BLN57),.WL(WL67));
sram_cell_6t_5 inst_cell_67_58 (.BL(BL58),.BLN(BLN58),.WL(WL67));
sram_cell_6t_5 inst_cell_67_59 (.BL(BL59),.BLN(BLN59),.WL(WL67));
sram_cell_6t_5 inst_cell_67_60 (.BL(BL60),.BLN(BLN60),.WL(WL67));
sram_cell_6t_5 inst_cell_67_61 (.BL(BL61),.BLN(BLN61),.WL(WL67));
sram_cell_6t_5 inst_cell_67_62 (.BL(BL62),.BLN(BLN62),.WL(WL67));
sram_cell_6t_5 inst_cell_67_63 (.BL(BL63),.BLN(BLN63),.WL(WL67));
sram_cell_6t_5 inst_cell_67_64 (.BL(BL64),.BLN(BLN64),.WL(WL67));
sram_cell_6t_5 inst_cell_67_65 (.BL(BL65),.BLN(BLN65),.WL(WL67));
sram_cell_6t_5 inst_cell_67_66 (.BL(BL66),.BLN(BLN66),.WL(WL67));
sram_cell_6t_5 inst_cell_67_67 (.BL(BL67),.BLN(BLN67),.WL(WL67));
sram_cell_6t_5 inst_cell_67_68 (.BL(BL68),.BLN(BLN68),.WL(WL67));
sram_cell_6t_5 inst_cell_67_69 (.BL(BL69),.BLN(BLN69),.WL(WL67));
sram_cell_6t_5 inst_cell_67_70 (.BL(BL70),.BLN(BLN70),.WL(WL67));
sram_cell_6t_5 inst_cell_67_71 (.BL(BL71),.BLN(BLN71),.WL(WL67));
sram_cell_6t_5 inst_cell_67_72 (.BL(BL72),.BLN(BLN72),.WL(WL67));
sram_cell_6t_5 inst_cell_67_73 (.BL(BL73),.BLN(BLN73),.WL(WL67));
sram_cell_6t_5 inst_cell_67_74 (.BL(BL74),.BLN(BLN74),.WL(WL67));
sram_cell_6t_5 inst_cell_67_75 (.BL(BL75),.BLN(BLN75),.WL(WL67));
sram_cell_6t_5 inst_cell_67_76 (.BL(BL76),.BLN(BLN76),.WL(WL67));
sram_cell_6t_5 inst_cell_67_77 (.BL(BL77),.BLN(BLN77),.WL(WL67));
sram_cell_6t_5 inst_cell_67_78 (.BL(BL78),.BLN(BLN78),.WL(WL67));
sram_cell_6t_5 inst_cell_67_79 (.BL(BL79),.BLN(BLN79),.WL(WL67));
sram_cell_6t_5 inst_cell_67_80 (.BL(BL80),.BLN(BLN80),.WL(WL67));
sram_cell_6t_5 inst_cell_67_81 (.BL(BL81),.BLN(BLN81),.WL(WL67));
sram_cell_6t_5 inst_cell_67_82 (.BL(BL82),.BLN(BLN82),.WL(WL67));
sram_cell_6t_5 inst_cell_67_83 (.BL(BL83),.BLN(BLN83),.WL(WL67));
sram_cell_6t_5 inst_cell_67_84 (.BL(BL84),.BLN(BLN84),.WL(WL67));
sram_cell_6t_5 inst_cell_67_85 (.BL(BL85),.BLN(BLN85),.WL(WL67));
sram_cell_6t_5 inst_cell_67_86 (.BL(BL86),.BLN(BLN86),.WL(WL67));
sram_cell_6t_5 inst_cell_67_87 (.BL(BL87),.BLN(BLN87),.WL(WL67));
sram_cell_6t_5 inst_cell_67_88 (.BL(BL88),.BLN(BLN88),.WL(WL67));
sram_cell_6t_5 inst_cell_67_89 (.BL(BL89),.BLN(BLN89),.WL(WL67));
sram_cell_6t_5 inst_cell_67_90 (.BL(BL90),.BLN(BLN90),.WL(WL67));
sram_cell_6t_5 inst_cell_67_91 (.BL(BL91),.BLN(BLN91),.WL(WL67));
sram_cell_6t_5 inst_cell_67_92 (.BL(BL92),.BLN(BLN92),.WL(WL67));
sram_cell_6t_5 inst_cell_67_93 (.BL(BL93),.BLN(BLN93),.WL(WL67));
sram_cell_6t_5 inst_cell_67_94 (.BL(BL94),.BLN(BLN94),.WL(WL67));
sram_cell_6t_5 inst_cell_67_95 (.BL(BL95),.BLN(BLN95),.WL(WL67));
sram_cell_6t_5 inst_cell_67_96 (.BL(BL96),.BLN(BLN96),.WL(WL67));
sram_cell_6t_5 inst_cell_67_97 (.BL(BL97),.BLN(BLN97),.WL(WL67));
sram_cell_6t_5 inst_cell_67_98 (.BL(BL98),.BLN(BLN98),.WL(WL67));
sram_cell_6t_5 inst_cell_67_99 (.BL(BL99),.BLN(BLN99),.WL(WL67));
sram_cell_6t_5 inst_cell_67_100 (.BL(BL100),.BLN(BLN100),.WL(WL67));
sram_cell_6t_5 inst_cell_67_101 (.BL(BL101),.BLN(BLN101),.WL(WL67));
sram_cell_6t_5 inst_cell_67_102 (.BL(BL102),.BLN(BLN102),.WL(WL67));
sram_cell_6t_5 inst_cell_67_103 (.BL(BL103),.BLN(BLN103),.WL(WL67));
sram_cell_6t_5 inst_cell_67_104 (.BL(BL104),.BLN(BLN104),.WL(WL67));
sram_cell_6t_5 inst_cell_67_105 (.BL(BL105),.BLN(BLN105),.WL(WL67));
sram_cell_6t_5 inst_cell_67_106 (.BL(BL106),.BLN(BLN106),.WL(WL67));
sram_cell_6t_5 inst_cell_67_107 (.BL(BL107),.BLN(BLN107),.WL(WL67));
sram_cell_6t_5 inst_cell_67_108 (.BL(BL108),.BLN(BLN108),.WL(WL67));
sram_cell_6t_5 inst_cell_67_109 (.BL(BL109),.BLN(BLN109),.WL(WL67));
sram_cell_6t_5 inst_cell_67_110 (.BL(BL110),.BLN(BLN110),.WL(WL67));
sram_cell_6t_5 inst_cell_67_111 (.BL(BL111),.BLN(BLN111),.WL(WL67));
sram_cell_6t_5 inst_cell_67_112 (.BL(BL112),.BLN(BLN112),.WL(WL67));
sram_cell_6t_5 inst_cell_67_113 (.BL(BL113),.BLN(BLN113),.WL(WL67));
sram_cell_6t_5 inst_cell_67_114 (.BL(BL114),.BLN(BLN114),.WL(WL67));
sram_cell_6t_5 inst_cell_67_115 (.BL(BL115),.BLN(BLN115),.WL(WL67));
sram_cell_6t_5 inst_cell_67_116 (.BL(BL116),.BLN(BLN116),.WL(WL67));
sram_cell_6t_5 inst_cell_67_117 (.BL(BL117),.BLN(BLN117),.WL(WL67));
sram_cell_6t_5 inst_cell_67_118 (.BL(BL118),.BLN(BLN118),.WL(WL67));
sram_cell_6t_5 inst_cell_67_119 (.BL(BL119),.BLN(BLN119),.WL(WL67));
sram_cell_6t_5 inst_cell_67_120 (.BL(BL120),.BLN(BLN120),.WL(WL67));
sram_cell_6t_5 inst_cell_67_121 (.BL(BL121),.BLN(BLN121),.WL(WL67));
sram_cell_6t_5 inst_cell_67_122 (.BL(BL122),.BLN(BLN122),.WL(WL67));
sram_cell_6t_5 inst_cell_67_123 (.BL(BL123),.BLN(BLN123),.WL(WL67));
sram_cell_6t_5 inst_cell_67_124 (.BL(BL124),.BLN(BLN124),.WL(WL67));
sram_cell_6t_5 inst_cell_67_125 (.BL(BL125),.BLN(BLN125),.WL(WL67));
sram_cell_6t_5 inst_cell_67_126 (.BL(BL126),.BLN(BLN126),.WL(WL67));
sram_cell_6t_5 inst_cell_67_127 (.BL(BL127),.BLN(BLN127),.WL(WL67));
sram_cell_6t_5 inst_cell_68_0 (.BL(BL0),.BLN(BLN0),.WL(WL68));
sram_cell_6t_5 inst_cell_68_1 (.BL(BL1),.BLN(BLN1),.WL(WL68));
sram_cell_6t_5 inst_cell_68_2 (.BL(BL2),.BLN(BLN2),.WL(WL68));
sram_cell_6t_5 inst_cell_68_3 (.BL(BL3),.BLN(BLN3),.WL(WL68));
sram_cell_6t_5 inst_cell_68_4 (.BL(BL4),.BLN(BLN4),.WL(WL68));
sram_cell_6t_5 inst_cell_68_5 (.BL(BL5),.BLN(BLN5),.WL(WL68));
sram_cell_6t_5 inst_cell_68_6 (.BL(BL6),.BLN(BLN6),.WL(WL68));
sram_cell_6t_5 inst_cell_68_7 (.BL(BL7),.BLN(BLN7),.WL(WL68));
sram_cell_6t_5 inst_cell_68_8 (.BL(BL8),.BLN(BLN8),.WL(WL68));
sram_cell_6t_5 inst_cell_68_9 (.BL(BL9),.BLN(BLN9),.WL(WL68));
sram_cell_6t_5 inst_cell_68_10 (.BL(BL10),.BLN(BLN10),.WL(WL68));
sram_cell_6t_5 inst_cell_68_11 (.BL(BL11),.BLN(BLN11),.WL(WL68));
sram_cell_6t_5 inst_cell_68_12 (.BL(BL12),.BLN(BLN12),.WL(WL68));
sram_cell_6t_5 inst_cell_68_13 (.BL(BL13),.BLN(BLN13),.WL(WL68));
sram_cell_6t_5 inst_cell_68_14 (.BL(BL14),.BLN(BLN14),.WL(WL68));
sram_cell_6t_5 inst_cell_68_15 (.BL(BL15),.BLN(BLN15),.WL(WL68));
sram_cell_6t_5 inst_cell_68_16 (.BL(BL16),.BLN(BLN16),.WL(WL68));
sram_cell_6t_5 inst_cell_68_17 (.BL(BL17),.BLN(BLN17),.WL(WL68));
sram_cell_6t_5 inst_cell_68_18 (.BL(BL18),.BLN(BLN18),.WL(WL68));
sram_cell_6t_5 inst_cell_68_19 (.BL(BL19),.BLN(BLN19),.WL(WL68));
sram_cell_6t_5 inst_cell_68_20 (.BL(BL20),.BLN(BLN20),.WL(WL68));
sram_cell_6t_5 inst_cell_68_21 (.BL(BL21),.BLN(BLN21),.WL(WL68));
sram_cell_6t_5 inst_cell_68_22 (.BL(BL22),.BLN(BLN22),.WL(WL68));
sram_cell_6t_5 inst_cell_68_23 (.BL(BL23),.BLN(BLN23),.WL(WL68));
sram_cell_6t_5 inst_cell_68_24 (.BL(BL24),.BLN(BLN24),.WL(WL68));
sram_cell_6t_5 inst_cell_68_25 (.BL(BL25),.BLN(BLN25),.WL(WL68));
sram_cell_6t_5 inst_cell_68_26 (.BL(BL26),.BLN(BLN26),.WL(WL68));
sram_cell_6t_5 inst_cell_68_27 (.BL(BL27),.BLN(BLN27),.WL(WL68));
sram_cell_6t_5 inst_cell_68_28 (.BL(BL28),.BLN(BLN28),.WL(WL68));
sram_cell_6t_5 inst_cell_68_29 (.BL(BL29),.BLN(BLN29),.WL(WL68));
sram_cell_6t_5 inst_cell_68_30 (.BL(BL30),.BLN(BLN30),.WL(WL68));
sram_cell_6t_5 inst_cell_68_31 (.BL(BL31),.BLN(BLN31),.WL(WL68));
sram_cell_6t_5 inst_cell_68_32 (.BL(BL32),.BLN(BLN32),.WL(WL68));
sram_cell_6t_5 inst_cell_68_33 (.BL(BL33),.BLN(BLN33),.WL(WL68));
sram_cell_6t_5 inst_cell_68_34 (.BL(BL34),.BLN(BLN34),.WL(WL68));
sram_cell_6t_5 inst_cell_68_35 (.BL(BL35),.BLN(BLN35),.WL(WL68));
sram_cell_6t_5 inst_cell_68_36 (.BL(BL36),.BLN(BLN36),.WL(WL68));
sram_cell_6t_5 inst_cell_68_37 (.BL(BL37),.BLN(BLN37),.WL(WL68));
sram_cell_6t_5 inst_cell_68_38 (.BL(BL38),.BLN(BLN38),.WL(WL68));
sram_cell_6t_5 inst_cell_68_39 (.BL(BL39),.BLN(BLN39),.WL(WL68));
sram_cell_6t_5 inst_cell_68_40 (.BL(BL40),.BLN(BLN40),.WL(WL68));
sram_cell_6t_5 inst_cell_68_41 (.BL(BL41),.BLN(BLN41),.WL(WL68));
sram_cell_6t_5 inst_cell_68_42 (.BL(BL42),.BLN(BLN42),.WL(WL68));
sram_cell_6t_5 inst_cell_68_43 (.BL(BL43),.BLN(BLN43),.WL(WL68));
sram_cell_6t_5 inst_cell_68_44 (.BL(BL44),.BLN(BLN44),.WL(WL68));
sram_cell_6t_5 inst_cell_68_45 (.BL(BL45),.BLN(BLN45),.WL(WL68));
sram_cell_6t_5 inst_cell_68_46 (.BL(BL46),.BLN(BLN46),.WL(WL68));
sram_cell_6t_5 inst_cell_68_47 (.BL(BL47),.BLN(BLN47),.WL(WL68));
sram_cell_6t_5 inst_cell_68_48 (.BL(BL48),.BLN(BLN48),.WL(WL68));
sram_cell_6t_5 inst_cell_68_49 (.BL(BL49),.BLN(BLN49),.WL(WL68));
sram_cell_6t_5 inst_cell_68_50 (.BL(BL50),.BLN(BLN50),.WL(WL68));
sram_cell_6t_5 inst_cell_68_51 (.BL(BL51),.BLN(BLN51),.WL(WL68));
sram_cell_6t_5 inst_cell_68_52 (.BL(BL52),.BLN(BLN52),.WL(WL68));
sram_cell_6t_5 inst_cell_68_53 (.BL(BL53),.BLN(BLN53),.WL(WL68));
sram_cell_6t_5 inst_cell_68_54 (.BL(BL54),.BLN(BLN54),.WL(WL68));
sram_cell_6t_5 inst_cell_68_55 (.BL(BL55),.BLN(BLN55),.WL(WL68));
sram_cell_6t_5 inst_cell_68_56 (.BL(BL56),.BLN(BLN56),.WL(WL68));
sram_cell_6t_5 inst_cell_68_57 (.BL(BL57),.BLN(BLN57),.WL(WL68));
sram_cell_6t_5 inst_cell_68_58 (.BL(BL58),.BLN(BLN58),.WL(WL68));
sram_cell_6t_5 inst_cell_68_59 (.BL(BL59),.BLN(BLN59),.WL(WL68));
sram_cell_6t_5 inst_cell_68_60 (.BL(BL60),.BLN(BLN60),.WL(WL68));
sram_cell_6t_5 inst_cell_68_61 (.BL(BL61),.BLN(BLN61),.WL(WL68));
sram_cell_6t_5 inst_cell_68_62 (.BL(BL62),.BLN(BLN62),.WL(WL68));
sram_cell_6t_5 inst_cell_68_63 (.BL(BL63),.BLN(BLN63),.WL(WL68));
sram_cell_6t_5 inst_cell_68_64 (.BL(BL64),.BLN(BLN64),.WL(WL68));
sram_cell_6t_5 inst_cell_68_65 (.BL(BL65),.BLN(BLN65),.WL(WL68));
sram_cell_6t_5 inst_cell_68_66 (.BL(BL66),.BLN(BLN66),.WL(WL68));
sram_cell_6t_5 inst_cell_68_67 (.BL(BL67),.BLN(BLN67),.WL(WL68));
sram_cell_6t_5 inst_cell_68_68 (.BL(BL68),.BLN(BLN68),.WL(WL68));
sram_cell_6t_5 inst_cell_68_69 (.BL(BL69),.BLN(BLN69),.WL(WL68));
sram_cell_6t_5 inst_cell_68_70 (.BL(BL70),.BLN(BLN70),.WL(WL68));
sram_cell_6t_5 inst_cell_68_71 (.BL(BL71),.BLN(BLN71),.WL(WL68));
sram_cell_6t_5 inst_cell_68_72 (.BL(BL72),.BLN(BLN72),.WL(WL68));
sram_cell_6t_5 inst_cell_68_73 (.BL(BL73),.BLN(BLN73),.WL(WL68));
sram_cell_6t_5 inst_cell_68_74 (.BL(BL74),.BLN(BLN74),.WL(WL68));
sram_cell_6t_5 inst_cell_68_75 (.BL(BL75),.BLN(BLN75),.WL(WL68));
sram_cell_6t_5 inst_cell_68_76 (.BL(BL76),.BLN(BLN76),.WL(WL68));
sram_cell_6t_5 inst_cell_68_77 (.BL(BL77),.BLN(BLN77),.WL(WL68));
sram_cell_6t_5 inst_cell_68_78 (.BL(BL78),.BLN(BLN78),.WL(WL68));
sram_cell_6t_5 inst_cell_68_79 (.BL(BL79),.BLN(BLN79),.WL(WL68));
sram_cell_6t_5 inst_cell_68_80 (.BL(BL80),.BLN(BLN80),.WL(WL68));
sram_cell_6t_5 inst_cell_68_81 (.BL(BL81),.BLN(BLN81),.WL(WL68));
sram_cell_6t_5 inst_cell_68_82 (.BL(BL82),.BLN(BLN82),.WL(WL68));
sram_cell_6t_5 inst_cell_68_83 (.BL(BL83),.BLN(BLN83),.WL(WL68));
sram_cell_6t_5 inst_cell_68_84 (.BL(BL84),.BLN(BLN84),.WL(WL68));
sram_cell_6t_5 inst_cell_68_85 (.BL(BL85),.BLN(BLN85),.WL(WL68));
sram_cell_6t_5 inst_cell_68_86 (.BL(BL86),.BLN(BLN86),.WL(WL68));
sram_cell_6t_5 inst_cell_68_87 (.BL(BL87),.BLN(BLN87),.WL(WL68));
sram_cell_6t_5 inst_cell_68_88 (.BL(BL88),.BLN(BLN88),.WL(WL68));
sram_cell_6t_5 inst_cell_68_89 (.BL(BL89),.BLN(BLN89),.WL(WL68));
sram_cell_6t_5 inst_cell_68_90 (.BL(BL90),.BLN(BLN90),.WL(WL68));
sram_cell_6t_5 inst_cell_68_91 (.BL(BL91),.BLN(BLN91),.WL(WL68));
sram_cell_6t_5 inst_cell_68_92 (.BL(BL92),.BLN(BLN92),.WL(WL68));
sram_cell_6t_5 inst_cell_68_93 (.BL(BL93),.BLN(BLN93),.WL(WL68));
sram_cell_6t_5 inst_cell_68_94 (.BL(BL94),.BLN(BLN94),.WL(WL68));
sram_cell_6t_5 inst_cell_68_95 (.BL(BL95),.BLN(BLN95),.WL(WL68));
sram_cell_6t_5 inst_cell_68_96 (.BL(BL96),.BLN(BLN96),.WL(WL68));
sram_cell_6t_5 inst_cell_68_97 (.BL(BL97),.BLN(BLN97),.WL(WL68));
sram_cell_6t_5 inst_cell_68_98 (.BL(BL98),.BLN(BLN98),.WL(WL68));
sram_cell_6t_5 inst_cell_68_99 (.BL(BL99),.BLN(BLN99),.WL(WL68));
sram_cell_6t_5 inst_cell_68_100 (.BL(BL100),.BLN(BLN100),.WL(WL68));
sram_cell_6t_5 inst_cell_68_101 (.BL(BL101),.BLN(BLN101),.WL(WL68));
sram_cell_6t_5 inst_cell_68_102 (.BL(BL102),.BLN(BLN102),.WL(WL68));
sram_cell_6t_5 inst_cell_68_103 (.BL(BL103),.BLN(BLN103),.WL(WL68));
sram_cell_6t_5 inst_cell_68_104 (.BL(BL104),.BLN(BLN104),.WL(WL68));
sram_cell_6t_5 inst_cell_68_105 (.BL(BL105),.BLN(BLN105),.WL(WL68));
sram_cell_6t_5 inst_cell_68_106 (.BL(BL106),.BLN(BLN106),.WL(WL68));
sram_cell_6t_5 inst_cell_68_107 (.BL(BL107),.BLN(BLN107),.WL(WL68));
sram_cell_6t_5 inst_cell_68_108 (.BL(BL108),.BLN(BLN108),.WL(WL68));
sram_cell_6t_5 inst_cell_68_109 (.BL(BL109),.BLN(BLN109),.WL(WL68));
sram_cell_6t_5 inst_cell_68_110 (.BL(BL110),.BLN(BLN110),.WL(WL68));
sram_cell_6t_5 inst_cell_68_111 (.BL(BL111),.BLN(BLN111),.WL(WL68));
sram_cell_6t_5 inst_cell_68_112 (.BL(BL112),.BLN(BLN112),.WL(WL68));
sram_cell_6t_5 inst_cell_68_113 (.BL(BL113),.BLN(BLN113),.WL(WL68));
sram_cell_6t_5 inst_cell_68_114 (.BL(BL114),.BLN(BLN114),.WL(WL68));
sram_cell_6t_5 inst_cell_68_115 (.BL(BL115),.BLN(BLN115),.WL(WL68));
sram_cell_6t_5 inst_cell_68_116 (.BL(BL116),.BLN(BLN116),.WL(WL68));
sram_cell_6t_5 inst_cell_68_117 (.BL(BL117),.BLN(BLN117),.WL(WL68));
sram_cell_6t_5 inst_cell_68_118 (.BL(BL118),.BLN(BLN118),.WL(WL68));
sram_cell_6t_5 inst_cell_68_119 (.BL(BL119),.BLN(BLN119),.WL(WL68));
sram_cell_6t_5 inst_cell_68_120 (.BL(BL120),.BLN(BLN120),.WL(WL68));
sram_cell_6t_5 inst_cell_68_121 (.BL(BL121),.BLN(BLN121),.WL(WL68));
sram_cell_6t_5 inst_cell_68_122 (.BL(BL122),.BLN(BLN122),.WL(WL68));
sram_cell_6t_5 inst_cell_68_123 (.BL(BL123),.BLN(BLN123),.WL(WL68));
sram_cell_6t_5 inst_cell_68_124 (.BL(BL124),.BLN(BLN124),.WL(WL68));
sram_cell_6t_5 inst_cell_68_125 (.BL(BL125),.BLN(BLN125),.WL(WL68));
sram_cell_6t_5 inst_cell_68_126 (.BL(BL126),.BLN(BLN126),.WL(WL68));
sram_cell_6t_5 inst_cell_68_127 (.BL(BL127),.BLN(BLN127),.WL(WL68));
sram_cell_6t_5 inst_cell_69_0 (.BL(BL0),.BLN(BLN0),.WL(WL69));
sram_cell_6t_5 inst_cell_69_1 (.BL(BL1),.BLN(BLN1),.WL(WL69));
sram_cell_6t_5 inst_cell_69_2 (.BL(BL2),.BLN(BLN2),.WL(WL69));
sram_cell_6t_5 inst_cell_69_3 (.BL(BL3),.BLN(BLN3),.WL(WL69));
sram_cell_6t_5 inst_cell_69_4 (.BL(BL4),.BLN(BLN4),.WL(WL69));
sram_cell_6t_5 inst_cell_69_5 (.BL(BL5),.BLN(BLN5),.WL(WL69));
sram_cell_6t_5 inst_cell_69_6 (.BL(BL6),.BLN(BLN6),.WL(WL69));
sram_cell_6t_5 inst_cell_69_7 (.BL(BL7),.BLN(BLN7),.WL(WL69));
sram_cell_6t_5 inst_cell_69_8 (.BL(BL8),.BLN(BLN8),.WL(WL69));
sram_cell_6t_5 inst_cell_69_9 (.BL(BL9),.BLN(BLN9),.WL(WL69));
sram_cell_6t_5 inst_cell_69_10 (.BL(BL10),.BLN(BLN10),.WL(WL69));
sram_cell_6t_5 inst_cell_69_11 (.BL(BL11),.BLN(BLN11),.WL(WL69));
sram_cell_6t_5 inst_cell_69_12 (.BL(BL12),.BLN(BLN12),.WL(WL69));
sram_cell_6t_5 inst_cell_69_13 (.BL(BL13),.BLN(BLN13),.WL(WL69));
sram_cell_6t_5 inst_cell_69_14 (.BL(BL14),.BLN(BLN14),.WL(WL69));
sram_cell_6t_5 inst_cell_69_15 (.BL(BL15),.BLN(BLN15),.WL(WL69));
sram_cell_6t_5 inst_cell_69_16 (.BL(BL16),.BLN(BLN16),.WL(WL69));
sram_cell_6t_5 inst_cell_69_17 (.BL(BL17),.BLN(BLN17),.WL(WL69));
sram_cell_6t_5 inst_cell_69_18 (.BL(BL18),.BLN(BLN18),.WL(WL69));
sram_cell_6t_5 inst_cell_69_19 (.BL(BL19),.BLN(BLN19),.WL(WL69));
sram_cell_6t_5 inst_cell_69_20 (.BL(BL20),.BLN(BLN20),.WL(WL69));
sram_cell_6t_5 inst_cell_69_21 (.BL(BL21),.BLN(BLN21),.WL(WL69));
sram_cell_6t_5 inst_cell_69_22 (.BL(BL22),.BLN(BLN22),.WL(WL69));
sram_cell_6t_5 inst_cell_69_23 (.BL(BL23),.BLN(BLN23),.WL(WL69));
sram_cell_6t_5 inst_cell_69_24 (.BL(BL24),.BLN(BLN24),.WL(WL69));
sram_cell_6t_5 inst_cell_69_25 (.BL(BL25),.BLN(BLN25),.WL(WL69));
sram_cell_6t_5 inst_cell_69_26 (.BL(BL26),.BLN(BLN26),.WL(WL69));
sram_cell_6t_5 inst_cell_69_27 (.BL(BL27),.BLN(BLN27),.WL(WL69));
sram_cell_6t_5 inst_cell_69_28 (.BL(BL28),.BLN(BLN28),.WL(WL69));
sram_cell_6t_5 inst_cell_69_29 (.BL(BL29),.BLN(BLN29),.WL(WL69));
sram_cell_6t_5 inst_cell_69_30 (.BL(BL30),.BLN(BLN30),.WL(WL69));
sram_cell_6t_5 inst_cell_69_31 (.BL(BL31),.BLN(BLN31),.WL(WL69));
sram_cell_6t_5 inst_cell_69_32 (.BL(BL32),.BLN(BLN32),.WL(WL69));
sram_cell_6t_5 inst_cell_69_33 (.BL(BL33),.BLN(BLN33),.WL(WL69));
sram_cell_6t_5 inst_cell_69_34 (.BL(BL34),.BLN(BLN34),.WL(WL69));
sram_cell_6t_5 inst_cell_69_35 (.BL(BL35),.BLN(BLN35),.WL(WL69));
sram_cell_6t_5 inst_cell_69_36 (.BL(BL36),.BLN(BLN36),.WL(WL69));
sram_cell_6t_5 inst_cell_69_37 (.BL(BL37),.BLN(BLN37),.WL(WL69));
sram_cell_6t_5 inst_cell_69_38 (.BL(BL38),.BLN(BLN38),.WL(WL69));
sram_cell_6t_5 inst_cell_69_39 (.BL(BL39),.BLN(BLN39),.WL(WL69));
sram_cell_6t_5 inst_cell_69_40 (.BL(BL40),.BLN(BLN40),.WL(WL69));
sram_cell_6t_5 inst_cell_69_41 (.BL(BL41),.BLN(BLN41),.WL(WL69));
sram_cell_6t_5 inst_cell_69_42 (.BL(BL42),.BLN(BLN42),.WL(WL69));
sram_cell_6t_5 inst_cell_69_43 (.BL(BL43),.BLN(BLN43),.WL(WL69));
sram_cell_6t_5 inst_cell_69_44 (.BL(BL44),.BLN(BLN44),.WL(WL69));
sram_cell_6t_5 inst_cell_69_45 (.BL(BL45),.BLN(BLN45),.WL(WL69));
sram_cell_6t_5 inst_cell_69_46 (.BL(BL46),.BLN(BLN46),.WL(WL69));
sram_cell_6t_5 inst_cell_69_47 (.BL(BL47),.BLN(BLN47),.WL(WL69));
sram_cell_6t_5 inst_cell_69_48 (.BL(BL48),.BLN(BLN48),.WL(WL69));
sram_cell_6t_5 inst_cell_69_49 (.BL(BL49),.BLN(BLN49),.WL(WL69));
sram_cell_6t_5 inst_cell_69_50 (.BL(BL50),.BLN(BLN50),.WL(WL69));
sram_cell_6t_5 inst_cell_69_51 (.BL(BL51),.BLN(BLN51),.WL(WL69));
sram_cell_6t_5 inst_cell_69_52 (.BL(BL52),.BLN(BLN52),.WL(WL69));
sram_cell_6t_5 inst_cell_69_53 (.BL(BL53),.BLN(BLN53),.WL(WL69));
sram_cell_6t_5 inst_cell_69_54 (.BL(BL54),.BLN(BLN54),.WL(WL69));
sram_cell_6t_5 inst_cell_69_55 (.BL(BL55),.BLN(BLN55),.WL(WL69));
sram_cell_6t_5 inst_cell_69_56 (.BL(BL56),.BLN(BLN56),.WL(WL69));
sram_cell_6t_5 inst_cell_69_57 (.BL(BL57),.BLN(BLN57),.WL(WL69));
sram_cell_6t_5 inst_cell_69_58 (.BL(BL58),.BLN(BLN58),.WL(WL69));
sram_cell_6t_5 inst_cell_69_59 (.BL(BL59),.BLN(BLN59),.WL(WL69));
sram_cell_6t_5 inst_cell_69_60 (.BL(BL60),.BLN(BLN60),.WL(WL69));
sram_cell_6t_5 inst_cell_69_61 (.BL(BL61),.BLN(BLN61),.WL(WL69));
sram_cell_6t_5 inst_cell_69_62 (.BL(BL62),.BLN(BLN62),.WL(WL69));
sram_cell_6t_5 inst_cell_69_63 (.BL(BL63),.BLN(BLN63),.WL(WL69));
sram_cell_6t_5 inst_cell_69_64 (.BL(BL64),.BLN(BLN64),.WL(WL69));
sram_cell_6t_5 inst_cell_69_65 (.BL(BL65),.BLN(BLN65),.WL(WL69));
sram_cell_6t_5 inst_cell_69_66 (.BL(BL66),.BLN(BLN66),.WL(WL69));
sram_cell_6t_5 inst_cell_69_67 (.BL(BL67),.BLN(BLN67),.WL(WL69));
sram_cell_6t_5 inst_cell_69_68 (.BL(BL68),.BLN(BLN68),.WL(WL69));
sram_cell_6t_5 inst_cell_69_69 (.BL(BL69),.BLN(BLN69),.WL(WL69));
sram_cell_6t_5 inst_cell_69_70 (.BL(BL70),.BLN(BLN70),.WL(WL69));
sram_cell_6t_5 inst_cell_69_71 (.BL(BL71),.BLN(BLN71),.WL(WL69));
sram_cell_6t_5 inst_cell_69_72 (.BL(BL72),.BLN(BLN72),.WL(WL69));
sram_cell_6t_5 inst_cell_69_73 (.BL(BL73),.BLN(BLN73),.WL(WL69));
sram_cell_6t_5 inst_cell_69_74 (.BL(BL74),.BLN(BLN74),.WL(WL69));
sram_cell_6t_5 inst_cell_69_75 (.BL(BL75),.BLN(BLN75),.WL(WL69));
sram_cell_6t_5 inst_cell_69_76 (.BL(BL76),.BLN(BLN76),.WL(WL69));
sram_cell_6t_5 inst_cell_69_77 (.BL(BL77),.BLN(BLN77),.WL(WL69));
sram_cell_6t_5 inst_cell_69_78 (.BL(BL78),.BLN(BLN78),.WL(WL69));
sram_cell_6t_5 inst_cell_69_79 (.BL(BL79),.BLN(BLN79),.WL(WL69));
sram_cell_6t_5 inst_cell_69_80 (.BL(BL80),.BLN(BLN80),.WL(WL69));
sram_cell_6t_5 inst_cell_69_81 (.BL(BL81),.BLN(BLN81),.WL(WL69));
sram_cell_6t_5 inst_cell_69_82 (.BL(BL82),.BLN(BLN82),.WL(WL69));
sram_cell_6t_5 inst_cell_69_83 (.BL(BL83),.BLN(BLN83),.WL(WL69));
sram_cell_6t_5 inst_cell_69_84 (.BL(BL84),.BLN(BLN84),.WL(WL69));
sram_cell_6t_5 inst_cell_69_85 (.BL(BL85),.BLN(BLN85),.WL(WL69));
sram_cell_6t_5 inst_cell_69_86 (.BL(BL86),.BLN(BLN86),.WL(WL69));
sram_cell_6t_5 inst_cell_69_87 (.BL(BL87),.BLN(BLN87),.WL(WL69));
sram_cell_6t_5 inst_cell_69_88 (.BL(BL88),.BLN(BLN88),.WL(WL69));
sram_cell_6t_5 inst_cell_69_89 (.BL(BL89),.BLN(BLN89),.WL(WL69));
sram_cell_6t_5 inst_cell_69_90 (.BL(BL90),.BLN(BLN90),.WL(WL69));
sram_cell_6t_5 inst_cell_69_91 (.BL(BL91),.BLN(BLN91),.WL(WL69));
sram_cell_6t_5 inst_cell_69_92 (.BL(BL92),.BLN(BLN92),.WL(WL69));
sram_cell_6t_5 inst_cell_69_93 (.BL(BL93),.BLN(BLN93),.WL(WL69));
sram_cell_6t_5 inst_cell_69_94 (.BL(BL94),.BLN(BLN94),.WL(WL69));
sram_cell_6t_5 inst_cell_69_95 (.BL(BL95),.BLN(BLN95),.WL(WL69));
sram_cell_6t_5 inst_cell_69_96 (.BL(BL96),.BLN(BLN96),.WL(WL69));
sram_cell_6t_5 inst_cell_69_97 (.BL(BL97),.BLN(BLN97),.WL(WL69));
sram_cell_6t_5 inst_cell_69_98 (.BL(BL98),.BLN(BLN98),.WL(WL69));
sram_cell_6t_5 inst_cell_69_99 (.BL(BL99),.BLN(BLN99),.WL(WL69));
sram_cell_6t_5 inst_cell_69_100 (.BL(BL100),.BLN(BLN100),.WL(WL69));
sram_cell_6t_5 inst_cell_69_101 (.BL(BL101),.BLN(BLN101),.WL(WL69));
sram_cell_6t_5 inst_cell_69_102 (.BL(BL102),.BLN(BLN102),.WL(WL69));
sram_cell_6t_5 inst_cell_69_103 (.BL(BL103),.BLN(BLN103),.WL(WL69));
sram_cell_6t_5 inst_cell_69_104 (.BL(BL104),.BLN(BLN104),.WL(WL69));
sram_cell_6t_5 inst_cell_69_105 (.BL(BL105),.BLN(BLN105),.WL(WL69));
sram_cell_6t_5 inst_cell_69_106 (.BL(BL106),.BLN(BLN106),.WL(WL69));
sram_cell_6t_5 inst_cell_69_107 (.BL(BL107),.BLN(BLN107),.WL(WL69));
sram_cell_6t_5 inst_cell_69_108 (.BL(BL108),.BLN(BLN108),.WL(WL69));
sram_cell_6t_5 inst_cell_69_109 (.BL(BL109),.BLN(BLN109),.WL(WL69));
sram_cell_6t_5 inst_cell_69_110 (.BL(BL110),.BLN(BLN110),.WL(WL69));
sram_cell_6t_5 inst_cell_69_111 (.BL(BL111),.BLN(BLN111),.WL(WL69));
sram_cell_6t_5 inst_cell_69_112 (.BL(BL112),.BLN(BLN112),.WL(WL69));
sram_cell_6t_5 inst_cell_69_113 (.BL(BL113),.BLN(BLN113),.WL(WL69));
sram_cell_6t_5 inst_cell_69_114 (.BL(BL114),.BLN(BLN114),.WL(WL69));
sram_cell_6t_5 inst_cell_69_115 (.BL(BL115),.BLN(BLN115),.WL(WL69));
sram_cell_6t_5 inst_cell_69_116 (.BL(BL116),.BLN(BLN116),.WL(WL69));
sram_cell_6t_5 inst_cell_69_117 (.BL(BL117),.BLN(BLN117),.WL(WL69));
sram_cell_6t_5 inst_cell_69_118 (.BL(BL118),.BLN(BLN118),.WL(WL69));
sram_cell_6t_5 inst_cell_69_119 (.BL(BL119),.BLN(BLN119),.WL(WL69));
sram_cell_6t_5 inst_cell_69_120 (.BL(BL120),.BLN(BLN120),.WL(WL69));
sram_cell_6t_5 inst_cell_69_121 (.BL(BL121),.BLN(BLN121),.WL(WL69));
sram_cell_6t_5 inst_cell_69_122 (.BL(BL122),.BLN(BLN122),.WL(WL69));
sram_cell_6t_5 inst_cell_69_123 (.BL(BL123),.BLN(BLN123),.WL(WL69));
sram_cell_6t_5 inst_cell_69_124 (.BL(BL124),.BLN(BLN124),.WL(WL69));
sram_cell_6t_5 inst_cell_69_125 (.BL(BL125),.BLN(BLN125),.WL(WL69));
sram_cell_6t_5 inst_cell_69_126 (.BL(BL126),.BLN(BLN126),.WL(WL69));
sram_cell_6t_5 inst_cell_69_127 (.BL(BL127),.BLN(BLN127),.WL(WL69));
sram_cell_6t_5 inst_cell_70_0 (.BL(BL0),.BLN(BLN0),.WL(WL70));
sram_cell_6t_5 inst_cell_70_1 (.BL(BL1),.BLN(BLN1),.WL(WL70));
sram_cell_6t_5 inst_cell_70_2 (.BL(BL2),.BLN(BLN2),.WL(WL70));
sram_cell_6t_5 inst_cell_70_3 (.BL(BL3),.BLN(BLN3),.WL(WL70));
sram_cell_6t_5 inst_cell_70_4 (.BL(BL4),.BLN(BLN4),.WL(WL70));
sram_cell_6t_5 inst_cell_70_5 (.BL(BL5),.BLN(BLN5),.WL(WL70));
sram_cell_6t_5 inst_cell_70_6 (.BL(BL6),.BLN(BLN6),.WL(WL70));
sram_cell_6t_5 inst_cell_70_7 (.BL(BL7),.BLN(BLN7),.WL(WL70));
sram_cell_6t_5 inst_cell_70_8 (.BL(BL8),.BLN(BLN8),.WL(WL70));
sram_cell_6t_5 inst_cell_70_9 (.BL(BL9),.BLN(BLN9),.WL(WL70));
sram_cell_6t_5 inst_cell_70_10 (.BL(BL10),.BLN(BLN10),.WL(WL70));
sram_cell_6t_5 inst_cell_70_11 (.BL(BL11),.BLN(BLN11),.WL(WL70));
sram_cell_6t_5 inst_cell_70_12 (.BL(BL12),.BLN(BLN12),.WL(WL70));
sram_cell_6t_5 inst_cell_70_13 (.BL(BL13),.BLN(BLN13),.WL(WL70));
sram_cell_6t_5 inst_cell_70_14 (.BL(BL14),.BLN(BLN14),.WL(WL70));
sram_cell_6t_5 inst_cell_70_15 (.BL(BL15),.BLN(BLN15),.WL(WL70));
sram_cell_6t_5 inst_cell_70_16 (.BL(BL16),.BLN(BLN16),.WL(WL70));
sram_cell_6t_5 inst_cell_70_17 (.BL(BL17),.BLN(BLN17),.WL(WL70));
sram_cell_6t_5 inst_cell_70_18 (.BL(BL18),.BLN(BLN18),.WL(WL70));
sram_cell_6t_5 inst_cell_70_19 (.BL(BL19),.BLN(BLN19),.WL(WL70));
sram_cell_6t_5 inst_cell_70_20 (.BL(BL20),.BLN(BLN20),.WL(WL70));
sram_cell_6t_5 inst_cell_70_21 (.BL(BL21),.BLN(BLN21),.WL(WL70));
sram_cell_6t_5 inst_cell_70_22 (.BL(BL22),.BLN(BLN22),.WL(WL70));
sram_cell_6t_5 inst_cell_70_23 (.BL(BL23),.BLN(BLN23),.WL(WL70));
sram_cell_6t_5 inst_cell_70_24 (.BL(BL24),.BLN(BLN24),.WL(WL70));
sram_cell_6t_5 inst_cell_70_25 (.BL(BL25),.BLN(BLN25),.WL(WL70));
sram_cell_6t_5 inst_cell_70_26 (.BL(BL26),.BLN(BLN26),.WL(WL70));
sram_cell_6t_5 inst_cell_70_27 (.BL(BL27),.BLN(BLN27),.WL(WL70));
sram_cell_6t_5 inst_cell_70_28 (.BL(BL28),.BLN(BLN28),.WL(WL70));
sram_cell_6t_5 inst_cell_70_29 (.BL(BL29),.BLN(BLN29),.WL(WL70));
sram_cell_6t_5 inst_cell_70_30 (.BL(BL30),.BLN(BLN30),.WL(WL70));
sram_cell_6t_5 inst_cell_70_31 (.BL(BL31),.BLN(BLN31),.WL(WL70));
sram_cell_6t_5 inst_cell_70_32 (.BL(BL32),.BLN(BLN32),.WL(WL70));
sram_cell_6t_5 inst_cell_70_33 (.BL(BL33),.BLN(BLN33),.WL(WL70));
sram_cell_6t_5 inst_cell_70_34 (.BL(BL34),.BLN(BLN34),.WL(WL70));
sram_cell_6t_5 inst_cell_70_35 (.BL(BL35),.BLN(BLN35),.WL(WL70));
sram_cell_6t_5 inst_cell_70_36 (.BL(BL36),.BLN(BLN36),.WL(WL70));
sram_cell_6t_5 inst_cell_70_37 (.BL(BL37),.BLN(BLN37),.WL(WL70));
sram_cell_6t_5 inst_cell_70_38 (.BL(BL38),.BLN(BLN38),.WL(WL70));
sram_cell_6t_5 inst_cell_70_39 (.BL(BL39),.BLN(BLN39),.WL(WL70));
sram_cell_6t_5 inst_cell_70_40 (.BL(BL40),.BLN(BLN40),.WL(WL70));
sram_cell_6t_5 inst_cell_70_41 (.BL(BL41),.BLN(BLN41),.WL(WL70));
sram_cell_6t_5 inst_cell_70_42 (.BL(BL42),.BLN(BLN42),.WL(WL70));
sram_cell_6t_5 inst_cell_70_43 (.BL(BL43),.BLN(BLN43),.WL(WL70));
sram_cell_6t_5 inst_cell_70_44 (.BL(BL44),.BLN(BLN44),.WL(WL70));
sram_cell_6t_5 inst_cell_70_45 (.BL(BL45),.BLN(BLN45),.WL(WL70));
sram_cell_6t_5 inst_cell_70_46 (.BL(BL46),.BLN(BLN46),.WL(WL70));
sram_cell_6t_5 inst_cell_70_47 (.BL(BL47),.BLN(BLN47),.WL(WL70));
sram_cell_6t_5 inst_cell_70_48 (.BL(BL48),.BLN(BLN48),.WL(WL70));
sram_cell_6t_5 inst_cell_70_49 (.BL(BL49),.BLN(BLN49),.WL(WL70));
sram_cell_6t_5 inst_cell_70_50 (.BL(BL50),.BLN(BLN50),.WL(WL70));
sram_cell_6t_5 inst_cell_70_51 (.BL(BL51),.BLN(BLN51),.WL(WL70));
sram_cell_6t_5 inst_cell_70_52 (.BL(BL52),.BLN(BLN52),.WL(WL70));
sram_cell_6t_5 inst_cell_70_53 (.BL(BL53),.BLN(BLN53),.WL(WL70));
sram_cell_6t_5 inst_cell_70_54 (.BL(BL54),.BLN(BLN54),.WL(WL70));
sram_cell_6t_5 inst_cell_70_55 (.BL(BL55),.BLN(BLN55),.WL(WL70));
sram_cell_6t_5 inst_cell_70_56 (.BL(BL56),.BLN(BLN56),.WL(WL70));
sram_cell_6t_5 inst_cell_70_57 (.BL(BL57),.BLN(BLN57),.WL(WL70));
sram_cell_6t_5 inst_cell_70_58 (.BL(BL58),.BLN(BLN58),.WL(WL70));
sram_cell_6t_5 inst_cell_70_59 (.BL(BL59),.BLN(BLN59),.WL(WL70));
sram_cell_6t_5 inst_cell_70_60 (.BL(BL60),.BLN(BLN60),.WL(WL70));
sram_cell_6t_5 inst_cell_70_61 (.BL(BL61),.BLN(BLN61),.WL(WL70));
sram_cell_6t_5 inst_cell_70_62 (.BL(BL62),.BLN(BLN62),.WL(WL70));
sram_cell_6t_5 inst_cell_70_63 (.BL(BL63),.BLN(BLN63),.WL(WL70));
sram_cell_6t_5 inst_cell_70_64 (.BL(BL64),.BLN(BLN64),.WL(WL70));
sram_cell_6t_5 inst_cell_70_65 (.BL(BL65),.BLN(BLN65),.WL(WL70));
sram_cell_6t_5 inst_cell_70_66 (.BL(BL66),.BLN(BLN66),.WL(WL70));
sram_cell_6t_5 inst_cell_70_67 (.BL(BL67),.BLN(BLN67),.WL(WL70));
sram_cell_6t_5 inst_cell_70_68 (.BL(BL68),.BLN(BLN68),.WL(WL70));
sram_cell_6t_5 inst_cell_70_69 (.BL(BL69),.BLN(BLN69),.WL(WL70));
sram_cell_6t_5 inst_cell_70_70 (.BL(BL70),.BLN(BLN70),.WL(WL70));
sram_cell_6t_5 inst_cell_70_71 (.BL(BL71),.BLN(BLN71),.WL(WL70));
sram_cell_6t_5 inst_cell_70_72 (.BL(BL72),.BLN(BLN72),.WL(WL70));
sram_cell_6t_5 inst_cell_70_73 (.BL(BL73),.BLN(BLN73),.WL(WL70));
sram_cell_6t_5 inst_cell_70_74 (.BL(BL74),.BLN(BLN74),.WL(WL70));
sram_cell_6t_5 inst_cell_70_75 (.BL(BL75),.BLN(BLN75),.WL(WL70));
sram_cell_6t_5 inst_cell_70_76 (.BL(BL76),.BLN(BLN76),.WL(WL70));
sram_cell_6t_5 inst_cell_70_77 (.BL(BL77),.BLN(BLN77),.WL(WL70));
sram_cell_6t_5 inst_cell_70_78 (.BL(BL78),.BLN(BLN78),.WL(WL70));
sram_cell_6t_5 inst_cell_70_79 (.BL(BL79),.BLN(BLN79),.WL(WL70));
sram_cell_6t_5 inst_cell_70_80 (.BL(BL80),.BLN(BLN80),.WL(WL70));
sram_cell_6t_5 inst_cell_70_81 (.BL(BL81),.BLN(BLN81),.WL(WL70));
sram_cell_6t_5 inst_cell_70_82 (.BL(BL82),.BLN(BLN82),.WL(WL70));
sram_cell_6t_5 inst_cell_70_83 (.BL(BL83),.BLN(BLN83),.WL(WL70));
sram_cell_6t_5 inst_cell_70_84 (.BL(BL84),.BLN(BLN84),.WL(WL70));
sram_cell_6t_5 inst_cell_70_85 (.BL(BL85),.BLN(BLN85),.WL(WL70));
sram_cell_6t_5 inst_cell_70_86 (.BL(BL86),.BLN(BLN86),.WL(WL70));
sram_cell_6t_5 inst_cell_70_87 (.BL(BL87),.BLN(BLN87),.WL(WL70));
sram_cell_6t_5 inst_cell_70_88 (.BL(BL88),.BLN(BLN88),.WL(WL70));
sram_cell_6t_5 inst_cell_70_89 (.BL(BL89),.BLN(BLN89),.WL(WL70));
sram_cell_6t_5 inst_cell_70_90 (.BL(BL90),.BLN(BLN90),.WL(WL70));
sram_cell_6t_5 inst_cell_70_91 (.BL(BL91),.BLN(BLN91),.WL(WL70));
sram_cell_6t_5 inst_cell_70_92 (.BL(BL92),.BLN(BLN92),.WL(WL70));
sram_cell_6t_5 inst_cell_70_93 (.BL(BL93),.BLN(BLN93),.WL(WL70));
sram_cell_6t_5 inst_cell_70_94 (.BL(BL94),.BLN(BLN94),.WL(WL70));
sram_cell_6t_5 inst_cell_70_95 (.BL(BL95),.BLN(BLN95),.WL(WL70));
sram_cell_6t_5 inst_cell_70_96 (.BL(BL96),.BLN(BLN96),.WL(WL70));
sram_cell_6t_5 inst_cell_70_97 (.BL(BL97),.BLN(BLN97),.WL(WL70));
sram_cell_6t_5 inst_cell_70_98 (.BL(BL98),.BLN(BLN98),.WL(WL70));
sram_cell_6t_5 inst_cell_70_99 (.BL(BL99),.BLN(BLN99),.WL(WL70));
sram_cell_6t_5 inst_cell_70_100 (.BL(BL100),.BLN(BLN100),.WL(WL70));
sram_cell_6t_5 inst_cell_70_101 (.BL(BL101),.BLN(BLN101),.WL(WL70));
sram_cell_6t_5 inst_cell_70_102 (.BL(BL102),.BLN(BLN102),.WL(WL70));
sram_cell_6t_5 inst_cell_70_103 (.BL(BL103),.BLN(BLN103),.WL(WL70));
sram_cell_6t_5 inst_cell_70_104 (.BL(BL104),.BLN(BLN104),.WL(WL70));
sram_cell_6t_5 inst_cell_70_105 (.BL(BL105),.BLN(BLN105),.WL(WL70));
sram_cell_6t_5 inst_cell_70_106 (.BL(BL106),.BLN(BLN106),.WL(WL70));
sram_cell_6t_5 inst_cell_70_107 (.BL(BL107),.BLN(BLN107),.WL(WL70));
sram_cell_6t_5 inst_cell_70_108 (.BL(BL108),.BLN(BLN108),.WL(WL70));
sram_cell_6t_5 inst_cell_70_109 (.BL(BL109),.BLN(BLN109),.WL(WL70));
sram_cell_6t_5 inst_cell_70_110 (.BL(BL110),.BLN(BLN110),.WL(WL70));
sram_cell_6t_5 inst_cell_70_111 (.BL(BL111),.BLN(BLN111),.WL(WL70));
sram_cell_6t_5 inst_cell_70_112 (.BL(BL112),.BLN(BLN112),.WL(WL70));
sram_cell_6t_5 inst_cell_70_113 (.BL(BL113),.BLN(BLN113),.WL(WL70));
sram_cell_6t_5 inst_cell_70_114 (.BL(BL114),.BLN(BLN114),.WL(WL70));
sram_cell_6t_5 inst_cell_70_115 (.BL(BL115),.BLN(BLN115),.WL(WL70));
sram_cell_6t_5 inst_cell_70_116 (.BL(BL116),.BLN(BLN116),.WL(WL70));
sram_cell_6t_5 inst_cell_70_117 (.BL(BL117),.BLN(BLN117),.WL(WL70));
sram_cell_6t_5 inst_cell_70_118 (.BL(BL118),.BLN(BLN118),.WL(WL70));
sram_cell_6t_5 inst_cell_70_119 (.BL(BL119),.BLN(BLN119),.WL(WL70));
sram_cell_6t_5 inst_cell_70_120 (.BL(BL120),.BLN(BLN120),.WL(WL70));
sram_cell_6t_5 inst_cell_70_121 (.BL(BL121),.BLN(BLN121),.WL(WL70));
sram_cell_6t_5 inst_cell_70_122 (.BL(BL122),.BLN(BLN122),.WL(WL70));
sram_cell_6t_5 inst_cell_70_123 (.BL(BL123),.BLN(BLN123),.WL(WL70));
sram_cell_6t_5 inst_cell_70_124 (.BL(BL124),.BLN(BLN124),.WL(WL70));
sram_cell_6t_5 inst_cell_70_125 (.BL(BL125),.BLN(BLN125),.WL(WL70));
sram_cell_6t_5 inst_cell_70_126 (.BL(BL126),.BLN(BLN126),.WL(WL70));
sram_cell_6t_5 inst_cell_70_127 (.BL(BL127),.BLN(BLN127),.WL(WL70));
sram_cell_6t_5 inst_cell_71_0 (.BL(BL0),.BLN(BLN0),.WL(WL71));
sram_cell_6t_5 inst_cell_71_1 (.BL(BL1),.BLN(BLN1),.WL(WL71));
sram_cell_6t_5 inst_cell_71_2 (.BL(BL2),.BLN(BLN2),.WL(WL71));
sram_cell_6t_5 inst_cell_71_3 (.BL(BL3),.BLN(BLN3),.WL(WL71));
sram_cell_6t_5 inst_cell_71_4 (.BL(BL4),.BLN(BLN4),.WL(WL71));
sram_cell_6t_5 inst_cell_71_5 (.BL(BL5),.BLN(BLN5),.WL(WL71));
sram_cell_6t_5 inst_cell_71_6 (.BL(BL6),.BLN(BLN6),.WL(WL71));
sram_cell_6t_5 inst_cell_71_7 (.BL(BL7),.BLN(BLN7),.WL(WL71));
sram_cell_6t_5 inst_cell_71_8 (.BL(BL8),.BLN(BLN8),.WL(WL71));
sram_cell_6t_5 inst_cell_71_9 (.BL(BL9),.BLN(BLN9),.WL(WL71));
sram_cell_6t_5 inst_cell_71_10 (.BL(BL10),.BLN(BLN10),.WL(WL71));
sram_cell_6t_5 inst_cell_71_11 (.BL(BL11),.BLN(BLN11),.WL(WL71));
sram_cell_6t_5 inst_cell_71_12 (.BL(BL12),.BLN(BLN12),.WL(WL71));
sram_cell_6t_5 inst_cell_71_13 (.BL(BL13),.BLN(BLN13),.WL(WL71));
sram_cell_6t_5 inst_cell_71_14 (.BL(BL14),.BLN(BLN14),.WL(WL71));
sram_cell_6t_5 inst_cell_71_15 (.BL(BL15),.BLN(BLN15),.WL(WL71));
sram_cell_6t_5 inst_cell_71_16 (.BL(BL16),.BLN(BLN16),.WL(WL71));
sram_cell_6t_5 inst_cell_71_17 (.BL(BL17),.BLN(BLN17),.WL(WL71));
sram_cell_6t_5 inst_cell_71_18 (.BL(BL18),.BLN(BLN18),.WL(WL71));
sram_cell_6t_5 inst_cell_71_19 (.BL(BL19),.BLN(BLN19),.WL(WL71));
sram_cell_6t_5 inst_cell_71_20 (.BL(BL20),.BLN(BLN20),.WL(WL71));
sram_cell_6t_5 inst_cell_71_21 (.BL(BL21),.BLN(BLN21),.WL(WL71));
sram_cell_6t_5 inst_cell_71_22 (.BL(BL22),.BLN(BLN22),.WL(WL71));
sram_cell_6t_5 inst_cell_71_23 (.BL(BL23),.BLN(BLN23),.WL(WL71));
sram_cell_6t_5 inst_cell_71_24 (.BL(BL24),.BLN(BLN24),.WL(WL71));
sram_cell_6t_5 inst_cell_71_25 (.BL(BL25),.BLN(BLN25),.WL(WL71));
sram_cell_6t_5 inst_cell_71_26 (.BL(BL26),.BLN(BLN26),.WL(WL71));
sram_cell_6t_5 inst_cell_71_27 (.BL(BL27),.BLN(BLN27),.WL(WL71));
sram_cell_6t_5 inst_cell_71_28 (.BL(BL28),.BLN(BLN28),.WL(WL71));
sram_cell_6t_5 inst_cell_71_29 (.BL(BL29),.BLN(BLN29),.WL(WL71));
sram_cell_6t_5 inst_cell_71_30 (.BL(BL30),.BLN(BLN30),.WL(WL71));
sram_cell_6t_5 inst_cell_71_31 (.BL(BL31),.BLN(BLN31),.WL(WL71));
sram_cell_6t_5 inst_cell_71_32 (.BL(BL32),.BLN(BLN32),.WL(WL71));
sram_cell_6t_5 inst_cell_71_33 (.BL(BL33),.BLN(BLN33),.WL(WL71));
sram_cell_6t_5 inst_cell_71_34 (.BL(BL34),.BLN(BLN34),.WL(WL71));
sram_cell_6t_5 inst_cell_71_35 (.BL(BL35),.BLN(BLN35),.WL(WL71));
sram_cell_6t_5 inst_cell_71_36 (.BL(BL36),.BLN(BLN36),.WL(WL71));
sram_cell_6t_5 inst_cell_71_37 (.BL(BL37),.BLN(BLN37),.WL(WL71));
sram_cell_6t_5 inst_cell_71_38 (.BL(BL38),.BLN(BLN38),.WL(WL71));
sram_cell_6t_5 inst_cell_71_39 (.BL(BL39),.BLN(BLN39),.WL(WL71));
sram_cell_6t_5 inst_cell_71_40 (.BL(BL40),.BLN(BLN40),.WL(WL71));
sram_cell_6t_5 inst_cell_71_41 (.BL(BL41),.BLN(BLN41),.WL(WL71));
sram_cell_6t_5 inst_cell_71_42 (.BL(BL42),.BLN(BLN42),.WL(WL71));
sram_cell_6t_5 inst_cell_71_43 (.BL(BL43),.BLN(BLN43),.WL(WL71));
sram_cell_6t_5 inst_cell_71_44 (.BL(BL44),.BLN(BLN44),.WL(WL71));
sram_cell_6t_5 inst_cell_71_45 (.BL(BL45),.BLN(BLN45),.WL(WL71));
sram_cell_6t_5 inst_cell_71_46 (.BL(BL46),.BLN(BLN46),.WL(WL71));
sram_cell_6t_5 inst_cell_71_47 (.BL(BL47),.BLN(BLN47),.WL(WL71));
sram_cell_6t_5 inst_cell_71_48 (.BL(BL48),.BLN(BLN48),.WL(WL71));
sram_cell_6t_5 inst_cell_71_49 (.BL(BL49),.BLN(BLN49),.WL(WL71));
sram_cell_6t_5 inst_cell_71_50 (.BL(BL50),.BLN(BLN50),.WL(WL71));
sram_cell_6t_5 inst_cell_71_51 (.BL(BL51),.BLN(BLN51),.WL(WL71));
sram_cell_6t_5 inst_cell_71_52 (.BL(BL52),.BLN(BLN52),.WL(WL71));
sram_cell_6t_5 inst_cell_71_53 (.BL(BL53),.BLN(BLN53),.WL(WL71));
sram_cell_6t_5 inst_cell_71_54 (.BL(BL54),.BLN(BLN54),.WL(WL71));
sram_cell_6t_5 inst_cell_71_55 (.BL(BL55),.BLN(BLN55),.WL(WL71));
sram_cell_6t_5 inst_cell_71_56 (.BL(BL56),.BLN(BLN56),.WL(WL71));
sram_cell_6t_5 inst_cell_71_57 (.BL(BL57),.BLN(BLN57),.WL(WL71));
sram_cell_6t_5 inst_cell_71_58 (.BL(BL58),.BLN(BLN58),.WL(WL71));
sram_cell_6t_5 inst_cell_71_59 (.BL(BL59),.BLN(BLN59),.WL(WL71));
sram_cell_6t_5 inst_cell_71_60 (.BL(BL60),.BLN(BLN60),.WL(WL71));
sram_cell_6t_5 inst_cell_71_61 (.BL(BL61),.BLN(BLN61),.WL(WL71));
sram_cell_6t_5 inst_cell_71_62 (.BL(BL62),.BLN(BLN62),.WL(WL71));
sram_cell_6t_5 inst_cell_71_63 (.BL(BL63),.BLN(BLN63),.WL(WL71));
sram_cell_6t_5 inst_cell_71_64 (.BL(BL64),.BLN(BLN64),.WL(WL71));
sram_cell_6t_5 inst_cell_71_65 (.BL(BL65),.BLN(BLN65),.WL(WL71));
sram_cell_6t_5 inst_cell_71_66 (.BL(BL66),.BLN(BLN66),.WL(WL71));
sram_cell_6t_5 inst_cell_71_67 (.BL(BL67),.BLN(BLN67),.WL(WL71));
sram_cell_6t_5 inst_cell_71_68 (.BL(BL68),.BLN(BLN68),.WL(WL71));
sram_cell_6t_5 inst_cell_71_69 (.BL(BL69),.BLN(BLN69),.WL(WL71));
sram_cell_6t_5 inst_cell_71_70 (.BL(BL70),.BLN(BLN70),.WL(WL71));
sram_cell_6t_5 inst_cell_71_71 (.BL(BL71),.BLN(BLN71),.WL(WL71));
sram_cell_6t_5 inst_cell_71_72 (.BL(BL72),.BLN(BLN72),.WL(WL71));
sram_cell_6t_5 inst_cell_71_73 (.BL(BL73),.BLN(BLN73),.WL(WL71));
sram_cell_6t_5 inst_cell_71_74 (.BL(BL74),.BLN(BLN74),.WL(WL71));
sram_cell_6t_5 inst_cell_71_75 (.BL(BL75),.BLN(BLN75),.WL(WL71));
sram_cell_6t_5 inst_cell_71_76 (.BL(BL76),.BLN(BLN76),.WL(WL71));
sram_cell_6t_5 inst_cell_71_77 (.BL(BL77),.BLN(BLN77),.WL(WL71));
sram_cell_6t_5 inst_cell_71_78 (.BL(BL78),.BLN(BLN78),.WL(WL71));
sram_cell_6t_5 inst_cell_71_79 (.BL(BL79),.BLN(BLN79),.WL(WL71));
sram_cell_6t_5 inst_cell_71_80 (.BL(BL80),.BLN(BLN80),.WL(WL71));
sram_cell_6t_5 inst_cell_71_81 (.BL(BL81),.BLN(BLN81),.WL(WL71));
sram_cell_6t_5 inst_cell_71_82 (.BL(BL82),.BLN(BLN82),.WL(WL71));
sram_cell_6t_5 inst_cell_71_83 (.BL(BL83),.BLN(BLN83),.WL(WL71));
sram_cell_6t_5 inst_cell_71_84 (.BL(BL84),.BLN(BLN84),.WL(WL71));
sram_cell_6t_5 inst_cell_71_85 (.BL(BL85),.BLN(BLN85),.WL(WL71));
sram_cell_6t_5 inst_cell_71_86 (.BL(BL86),.BLN(BLN86),.WL(WL71));
sram_cell_6t_5 inst_cell_71_87 (.BL(BL87),.BLN(BLN87),.WL(WL71));
sram_cell_6t_5 inst_cell_71_88 (.BL(BL88),.BLN(BLN88),.WL(WL71));
sram_cell_6t_5 inst_cell_71_89 (.BL(BL89),.BLN(BLN89),.WL(WL71));
sram_cell_6t_5 inst_cell_71_90 (.BL(BL90),.BLN(BLN90),.WL(WL71));
sram_cell_6t_5 inst_cell_71_91 (.BL(BL91),.BLN(BLN91),.WL(WL71));
sram_cell_6t_5 inst_cell_71_92 (.BL(BL92),.BLN(BLN92),.WL(WL71));
sram_cell_6t_5 inst_cell_71_93 (.BL(BL93),.BLN(BLN93),.WL(WL71));
sram_cell_6t_5 inst_cell_71_94 (.BL(BL94),.BLN(BLN94),.WL(WL71));
sram_cell_6t_5 inst_cell_71_95 (.BL(BL95),.BLN(BLN95),.WL(WL71));
sram_cell_6t_5 inst_cell_71_96 (.BL(BL96),.BLN(BLN96),.WL(WL71));
sram_cell_6t_5 inst_cell_71_97 (.BL(BL97),.BLN(BLN97),.WL(WL71));
sram_cell_6t_5 inst_cell_71_98 (.BL(BL98),.BLN(BLN98),.WL(WL71));
sram_cell_6t_5 inst_cell_71_99 (.BL(BL99),.BLN(BLN99),.WL(WL71));
sram_cell_6t_5 inst_cell_71_100 (.BL(BL100),.BLN(BLN100),.WL(WL71));
sram_cell_6t_5 inst_cell_71_101 (.BL(BL101),.BLN(BLN101),.WL(WL71));
sram_cell_6t_5 inst_cell_71_102 (.BL(BL102),.BLN(BLN102),.WL(WL71));
sram_cell_6t_5 inst_cell_71_103 (.BL(BL103),.BLN(BLN103),.WL(WL71));
sram_cell_6t_5 inst_cell_71_104 (.BL(BL104),.BLN(BLN104),.WL(WL71));
sram_cell_6t_5 inst_cell_71_105 (.BL(BL105),.BLN(BLN105),.WL(WL71));
sram_cell_6t_5 inst_cell_71_106 (.BL(BL106),.BLN(BLN106),.WL(WL71));
sram_cell_6t_5 inst_cell_71_107 (.BL(BL107),.BLN(BLN107),.WL(WL71));
sram_cell_6t_5 inst_cell_71_108 (.BL(BL108),.BLN(BLN108),.WL(WL71));
sram_cell_6t_5 inst_cell_71_109 (.BL(BL109),.BLN(BLN109),.WL(WL71));
sram_cell_6t_5 inst_cell_71_110 (.BL(BL110),.BLN(BLN110),.WL(WL71));
sram_cell_6t_5 inst_cell_71_111 (.BL(BL111),.BLN(BLN111),.WL(WL71));
sram_cell_6t_5 inst_cell_71_112 (.BL(BL112),.BLN(BLN112),.WL(WL71));
sram_cell_6t_5 inst_cell_71_113 (.BL(BL113),.BLN(BLN113),.WL(WL71));
sram_cell_6t_5 inst_cell_71_114 (.BL(BL114),.BLN(BLN114),.WL(WL71));
sram_cell_6t_5 inst_cell_71_115 (.BL(BL115),.BLN(BLN115),.WL(WL71));
sram_cell_6t_5 inst_cell_71_116 (.BL(BL116),.BLN(BLN116),.WL(WL71));
sram_cell_6t_5 inst_cell_71_117 (.BL(BL117),.BLN(BLN117),.WL(WL71));
sram_cell_6t_5 inst_cell_71_118 (.BL(BL118),.BLN(BLN118),.WL(WL71));
sram_cell_6t_5 inst_cell_71_119 (.BL(BL119),.BLN(BLN119),.WL(WL71));
sram_cell_6t_5 inst_cell_71_120 (.BL(BL120),.BLN(BLN120),.WL(WL71));
sram_cell_6t_5 inst_cell_71_121 (.BL(BL121),.BLN(BLN121),.WL(WL71));
sram_cell_6t_5 inst_cell_71_122 (.BL(BL122),.BLN(BLN122),.WL(WL71));
sram_cell_6t_5 inst_cell_71_123 (.BL(BL123),.BLN(BLN123),.WL(WL71));
sram_cell_6t_5 inst_cell_71_124 (.BL(BL124),.BLN(BLN124),.WL(WL71));
sram_cell_6t_5 inst_cell_71_125 (.BL(BL125),.BLN(BLN125),.WL(WL71));
sram_cell_6t_5 inst_cell_71_126 (.BL(BL126),.BLN(BLN126),.WL(WL71));
sram_cell_6t_5 inst_cell_71_127 (.BL(BL127),.BLN(BLN127),.WL(WL71));
sram_cell_6t_5 inst_cell_72_0 (.BL(BL0),.BLN(BLN0),.WL(WL72));
sram_cell_6t_5 inst_cell_72_1 (.BL(BL1),.BLN(BLN1),.WL(WL72));
sram_cell_6t_5 inst_cell_72_2 (.BL(BL2),.BLN(BLN2),.WL(WL72));
sram_cell_6t_5 inst_cell_72_3 (.BL(BL3),.BLN(BLN3),.WL(WL72));
sram_cell_6t_5 inst_cell_72_4 (.BL(BL4),.BLN(BLN4),.WL(WL72));
sram_cell_6t_5 inst_cell_72_5 (.BL(BL5),.BLN(BLN5),.WL(WL72));
sram_cell_6t_5 inst_cell_72_6 (.BL(BL6),.BLN(BLN6),.WL(WL72));
sram_cell_6t_5 inst_cell_72_7 (.BL(BL7),.BLN(BLN7),.WL(WL72));
sram_cell_6t_5 inst_cell_72_8 (.BL(BL8),.BLN(BLN8),.WL(WL72));
sram_cell_6t_5 inst_cell_72_9 (.BL(BL9),.BLN(BLN9),.WL(WL72));
sram_cell_6t_5 inst_cell_72_10 (.BL(BL10),.BLN(BLN10),.WL(WL72));
sram_cell_6t_5 inst_cell_72_11 (.BL(BL11),.BLN(BLN11),.WL(WL72));
sram_cell_6t_5 inst_cell_72_12 (.BL(BL12),.BLN(BLN12),.WL(WL72));
sram_cell_6t_5 inst_cell_72_13 (.BL(BL13),.BLN(BLN13),.WL(WL72));
sram_cell_6t_5 inst_cell_72_14 (.BL(BL14),.BLN(BLN14),.WL(WL72));
sram_cell_6t_5 inst_cell_72_15 (.BL(BL15),.BLN(BLN15),.WL(WL72));
sram_cell_6t_5 inst_cell_72_16 (.BL(BL16),.BLN(BLN16),.WL(WL72));
sram_cell_6t_5 inst_cell_72_17 (.BL(BL17),.BLN(BLN17),.WL(WL72));
sram_cell_6t_5 inst_cell_72_18 (.BL(BL18),.BLN(BLN18),.WL(WL72));
sram_cell_6t_5 inst_cell_72_19 (.BL(BL19),.BLN(BLN19),.WL(WL72));
sram_cell_6t_5 inst_cell_72_20 (.BL(BL20),.BLN(BLN20),.WL(WL72));
sram_cell_6t_5 inst_cell_72_21 (.BL(BL21),.BLN(BLN21),.WL(WL72));
sram_cell_6t_5 inst_cell_72_22 (.BL(BL22),.BLN(BLN22),.WL(WL72));
sram_cell_6t_5 inst_cell_72_23 (.BL(BL23),.BLN(BLN23),.WL(WL72));
sram_cell_6t_5 inst_cell_72_24 (.BL(BL24),.BLN(BLN24),.WL(WL72));
sram_cell_6t_5 inst_cell_72_25 (.BL(BL25),.BLN(BLN25),.WL(WL72));
sram_cell_6t_5 inst_cell_72_26 (.BL(BL26),.BLN(BLN26),.WL(WL72));
sram_cell_6t_5 inst_cell_72_27 (.BL(BL27),.BLN(BLN27),.WL(WL72));
sram_cell_6t_5 inst_cell_72_28 (.BL(BL28),.BLN(BLN28),.WL(WL72));
sram_cell_6t_5 inst_cell_72_29 (.BL(BL29),.BLN(BLN29),.WL(WL72));
sram_cell_6t_5 inst_cell_72_30 (.BL(BL30),.BLN(BLN30),.WL(WL72));
sram_cell_6t_5 inst_cell_72_31 (.BL(BL31),.BLN(BLN31),.WL(WL72));
sram_cell_6t_5 inst_cell_72_32 (.BL(BL32),.BLN(BLN32),.WL(WL72));
sram_cell_6t_5 inst_cell_72_33 (.BL(BL33),.BLN(BLN33),.WL(WL72));
sram_cell_6t_5 inst_cell_72_34 (.BL(BL34),.BLN(BLN34),.WL(WL72));
sram_cell_6t_5 inst_cell_72_35 (.BL(BL35),.BLN(BLN35),.WL(WL72));
sram_cell_6t_5 inst_cell_72_36 (.BL(BL36),.BLN(BLN36),.WL(WL72));
sram_cell_6t_5 inst_cell_72_37 (.BL(BL37),.BLN(BLN37),.WL(WL72));
sram_cell_6t_5 inst_cell_72_38 (.BL(BL38),.BLN(BLN38),.WL(WL72));
sram_cell_6t_5 inst_cell_72_39 (.BL(BL39),.BLN(BLN39),.WL(WL72));
sram_cell_6t_5 inst_cell_72_40 (.BL(BL40),.BLN(BLN40),.WL(WL72));
sram_cell_6t_5 inst_cell_72_41 (.BL(BL41),.BLN(BLN41),.WL(WL72));
sram_cell_6t_5 inst_cell_72_42 (.BL(BL42),.BLN(BLN42),.WL(WL72));
sram_cell_6t_5 inst_cell_72_43 (.BL(BL43),.BLN(BLN43),.WL(WL72));
sram_cell_6t_5 inst_cell_72_44 (.BL(BL44),.BLN(BLN44),.WL(WL72));
sram_cell_6t_5 inst_cell_72_45 (.BL(BL45),.BLN(BLN45),.WL(WL72));
sram_cell_6t_5 inst_cell_72_46 (.BL(BL46),.BLN(BLN46),.WL(WL72));
sram_cell_6t_5 inst_cell_72_47 (.BL(BL47),.BLN(BLN47),.WL(WL72));
sram_cell_6t_5 inst_cell_72_48 (.BL(BL48),.BLN(BLN48),.WL(WL72));
sram_cell_6t_5 inst_cell_72_49 (.BL(BL49),.BLN(BLN49),.WL(WL72));
sram_cell_6t_5 inst_cell_72_50 (.BL(BL50),.BLN(BLN50),.WL(WL72));
sram_cell_6t_5 inst_cell_72_51 (.BL(BL51),.BLN(BLN51),.WL(WL72));
sram_cell_6t_5 inst_cell_72_52 (.BL(BL52),.BLN(BLN52),.WL(WL72));
sram_cell_6t_5 inst_cell_72_53 (.BL(BL53),.BLN(BLN53),.WL(WL72));
sram_cell_6t_5 inst_cell_72_54 (.BL(BL54),.BLN(BLN54),.WL(WL72));
sram_cell_6t_5 inst_cell_72_55 (.BL(BL55),.BLN(BLN55),.WL(WL72));
sram_cell_6t_5 inst_cell_72_56 (.BL(BL56),.BLN(BLN56),.WL(WL72));
sram_cell_6t_5 inst_cell_72_57 (.BL(BL57),.BLN(BLN57),.WL(WL72));
sram_cell_6t_5 inst_cell_72_58 (.BL(BL58),.BLN(BLN58),.WL(WL72));
sram_cell_6t_5 inst_cell_72_59 (.BL(BL59),.BLN(BLN59),.WL(WL72));
sram_cell_6t_5 inst_cell_72_60 (.BL(BL60),.BLN(BLN60),.WL(WL72));
sram_cell_6t_5 inst_cell_72_61 (.BL(BL61),.BLN(BLN61),.WL(WL72));
sram_cell_6t_5 inst_cell_72_62 (.BL(BL62),.BLN(BLN62),.WL(WL72));
sram_cell_6t_5 inst_cell_72_63 (.BL(BL63),.BLN(BLN63),.WL(WL72));
sram_cell_6t_5 inst_cell_72_64 (.BL(BL64),.BLN(BLN64),.WL(WL72));
sram_cell_6t_5 inst_cell_72_65 (.BL(BL65),.BLN(BLN65),.WL(WL72));
sram_cell_6t_5 inst_cell_72_66 (.BL(BL66),.BLN(BLN66),.WL(WL72));
sram_cell_6t_5 inst_cell_72_67 (.BL(BL67),.BLN(BLN67),.WL(WL72));
sram_cell_6t_5 inst_cell_72_68 (.BL(BL68),.BLN(BLN68),.WL(WL72));
sram_cell_6t_5 inst_cell_72_69 (.BL(BL69),.BLN(BLN69),.WL(WL72));
sram_cell_6t_5 inst_cell_72_70 (.BL(BL70),.BLN(BLN70),.WL(WL72));
sram_cell_6t_5 inst_cell_72_71 (.BL(BL71),.BLN(BLN71),.WL(WL72));
sram_cell_6t_5 inst_cell_72_72 (.BL(BL72),.BLN(BLN72),.WL(WL72));
sram_cell_6t_5 inst_cell_72_73 (.BL(BL73),.BLN(BLN73),.WL(WL72));
sram_cell_6t_5 inst_cell_72_74 (.BL(BL74),.BLN(BLN74),.WL(WL72));
sram_cell_6t_5 inst_cell_72_75 (.BL(BL75),.BLN(BLN75),.WL(WL72));
sram_cell_6t_5 inst_cell_72_76 (.BL(BL76),.BLN(BLN76),.WL(WL72));
sram_cell_6t_5 inst_cell_72_77 (.BL(BL77),.BLN(BLN77),.WL(WL72));
sram_cell_6t_5 inst_cell_72_78 (.BL(BL78),.BLN(BLN78),.WL(WL72));
sram_cell_6t_5 inst_cell_72_79 (.BL(BL79),.BLN(BLN79),.WL(WL72));
sram_cell_6t_5 inst_cell_72_80 (.BL(BL80),.BLN(BLN80),.WL(WL72));
sram_cell_6t_5 inst_cell_72_81 (.BL(BL81),.BLN(BLN81),.WL(WL72));
sram_cell_6t_5 inst_cell_72_82 (.BL(BL82),.BLN(BLN82),.WL(WL72));
sram_cell_6t_5 inst_cell_72_83 (.BL(BL83),.BLN(BLN83),.WL(WL72));
sram_cell_6t_5 inst_cell_72_84 (.BL(BL84),.BLN(BLN84),.WL(WL72));
sram_cell_6t_5 inst_cell_72_85 (.BL(BL85),.BLN(BLN85),.WL(WL72));
sram_cell_6t_5 inst_cell_72_86 (.BL(BL86),.BLN(BLN86),.WL(WL72));
sram_cell_6t_5 inst_cell_72_87 (.BL(BL87),.BLN(BLN87),.WL(WL72));
sram_cell_6t_5 inst_cell_72_88 (.BL(BL88),.BLN(BLN88),.WL(WL72));
sram_cell_6t_5 inst_cell_72_89 (.BL(BL89),.BLN(BLN89),.WL(WL72));
sram_cell_6t_5 inst_cell_72_90 (.BL(BL90),.BLN(BLN90),.WL(WL72));
sram_cell_6t_5 inst_cell_72_91 (.BL(BL91),.BLN(BLN91),.WL(WL72));
sram_cell_6t_5 inst_cell_72_92 (.BL(BL92),.BLN(BLN92),.WL(WL72));
sram_cell_6t_5 inst_cell_72_93 (.BL(BL93),.BLN(BLN93),.WL(WL72));
sram_cell_6t_5 inst_cell_72_94 (.BL(BL94),.BLN(BLN94),.WL(WL72));
sram_cell_6t_5 inst_cell_72_95 (.BL(BL95),.BLN(BLN95),.WL(WL72));
sram_cell_6t_5 inst_cell_72_96 (.BL(BL96),.BLN(BLN96),.WL(WL72));
sram_cell_6t_5 inst_cell_72_97 (.BL(BL97),.BLN(BLN97),.WL(WL72));
sram_cell_6t_5 inst_cell_72_98 (.BL(BL98),.BLN(BLN98),.WL(WL72));
sram_cell_6t_5 inst_cell_72_99 (.BL(BL99),.BLN(BLN99),.WL(WL72));
sram_cell_6t_5 inst_cell_72_100 (.BL(BL100),.BLN(BLN100),.WL(WL72));
sram_cell_6t_5 inst_cell_72_101 (.BL(BL101),.BLN(BLN101),.WL(WL72));
sram_cell_6t_5 inst_cell_72_102 (.BL(BL102),.BLN(BLN102),.WL(WL72));
sram_cell_6t_5 inst_cell_72_103 (.BL(BL103),.BLN(BLN103),.WL(WL72));
sram_cell_6t_5 inst_cell_72_104 (.BL(BL104),.BLN(BLN104),.WL(WL72));
sram_cell_6t_5 inst_cell_72_105 (.BL(BL105),.BLN(BLN105),.WL(WL72));
sram_cell_6t_5 inst_cell_72_106 (.BL(BL106),.BLN(BLN106),.WL(WL72));
sram_cell_6t_5 inst_cell_72_107 (.BL(BL107),.BLN(BLN107),.WL(WL72));
sram_cell_6t_5 inst_cell_72_108 (.BL(BL108),.BLN(BLN108),.WL(WL72));
sram_cell_6t_5 inst_cell_72_109 (.BL(BL109),.BLN(BLN109),.WL(WL72));
sram_cell_6t_5 inst_cell_72_110 (.BL(BL110),.BLN(BLN110),.WL(WL72));
sram_cell_6t_5 inst_cell_72_111 (.BL(BL111),.BLN(BLN111),.WL(WL72));
sram_cell_6t_5 inst_cell_72_112 (.BL(BL112),.BLN(BLN112),.WL(WL72));
sram_cell_6t_5 inst_cell_72_113 (.BL(BL113),.BLN(BLN113),.WL(WL72));
sram_cell_6t_5 inst_cell_72_114 (.BL(BL114),.BLN(BLN114),.WL(WL72));
sram_cell_6t_5 inst_cell_72_115 (.BL(BL115),.BLN(BLN115),.WL(WL72));
sram_cell_6t_5 inst_cell_72_116 (.BL(BL116),.BLN(BLN116),.WL(WL72));
sram_cell_6t_5 inst_cell_72_117 (.BL(BL117),.BLN(BLN117),.WL(WL72));
sram_cell_6t_5 inst_cell_72_118 (.BL(BL118),.BLN(BLN118),.WL(WL72));
sram_cell_6t_5 inst_cell_72_119 (.BL(BL119),.BLN(BLN119),.WL(WL72));
sram_cell_6t_5 inst_cell_72_120 (.BL(BL120),.BLN(BLN120),.WL(WL72));
sram_cell_6t_5 inst_cell_72_121 (.BL(BL121),.BLN(BLN121),.WL(WL72));
sram_cell_6t_5 inst_cell_72_122 (.BL(BL122),.BLN(BLN122),.WL(WL72));
sram_cell_6t_5 inst_cell_72_123 (.BL(BL123),.BLN(BLN123),.WL(WL72));
sram_cell_6t_5 inst_cell_72_124 (.BL(BL124),.BLN(BLN124),.WL(WL72));
sram_cell_6t_5 inst_cell_72_125 (.BL(BL125),.BLN(BLN125),.WL(WL72));
sram_cell_6t_5 inst_cell_72_126 (.BL(BL126),.BLN(BLN126),.WL(WL72));
sram_cell_6t_5 inst_cell_72_127 (.BL(BL127),.BLN(BLN127),.WL(WL72));
sram_cell_6t_5 inst_cell_73_0 (.BL(BL0),.BLN(BLN0),.WL(WL73));
sram_cell_6t_5 inst_cell_73_1 (.BL(BL1),.BLN(BLN1),.WL(WL73));
sram_cell_6t_5 inst_cell_73_2 (.BL(BL2),.BLN(BLN2),.WL(WL73));
sram_cell_6t_5 inst_cell_73_3 (.BL(BL3),.BLN(BLN3),.WL(WL73));
sram_cell_6t_5 inst_cell_73_4 (.BL(BL4),.BLN(BLN4),.WL(WL73));
sram_cell_6t_5 inst_cell_73_5 (.BL(BL5),.BLN(BLN5),.WL(WL73));
sram_cell_6t_5 inst_cell_73_6 (.BL(BL6),.BLN(BLN6),.WL(WL73));
sram_cell_6t_5 inst_cell_73_7 (.BL(BL7),.BLN(BLN7),.WL(WL73));
sram_cell_6t_5 inst_cell_73_8 (.BL(BL8),.BLN(BLN8),.WL(WL73));
sram_cell_6t_5 inst_cell_73_9 (.BL(BL9),.BLN(BLN9),.WL(WL73));
sram_cell_6t_5 inst_cell_73_10 (.BL(BL10),.BLN(BLN10),.WL(WL73));
sram_cell_6t_5 inst_cell_73_11 (.BL(BL11),.BLN(BLN11),.WL(WL73));
sram_cell_6t_5 inst_cell_73_12 (.BL(BL12),.BLN(BLN12),.WL(WL73));
sram_cell_6t_5 inst_cell_73_13 (.BL(BL13),.BLN(BLN13),.WL(WL73));
sram_cell_6t_5 inst_cell_73_14 (.BL(BL14),.BLN(BLN14),.WL(WL73));
sram_cell_6t_5 inst_cell_73_15 (.BL(BL15),.BLN(BLN15),.WL(WL73));
sram_cell_6t_5 inst_cell_73_16 (.BL(BL16),.BLN(BLN16),.WL(WL73));
sram_cell_6t_5 inst_cell_73_17 (.BL(BL17),.BLN(BLN17),.WL(WL73));
sram_cell_6t_5 inst_cell_73_18 (.BL(BL18),.BLN(BLN18),.WL(WL73));
sram_cell_6t_5 inst_cell_73_19 (.BL(BL19),.BLN(BLN19),.WL(WL73));
sram_cell_6t_5 inst_cell_73_20 (.BL(BL20),.BLN(BLN20),.WL(WL73));
sram_cell_6t_5 inst_cell_73_21 (.BL(BL21),.BLN(BLN21),.WL(WL73));
sram_cell_6t_5 inst_cell_73_22 (.BL(BL22),.BLN(BLN22),.WL(WL73));
sram_cell_6t_5 inst_cell_73_23 (.BL(BL23),.BLN(BLN23),.WL(WL73));
sram_cell_6t_5 inst_cell_73_24 (.BL(BL24),.BLN(BLN24),.WL(WL73));
sram_cell_6t_5 inst_cell_73_25 (.BL(BL25),.BLN(BLN25),.WL(WL73));
sram_cell_6t_5 inst_cell_73_26 (.BL(BL26),.BLN(BLN26),.WL(WL73));
sram_cell_6t_5 inst_cell_73_27 (.BL(BL27),.BLN(BLN27),.WL(WL73));
sram_cell_6t_5 inst_cell_73_28 (.BL(BL28),.BLN(BLN28),.WL(WL73));
sram_cell_6t_5 inst_cell_73_29 (.BL(BL29),.BLN(BLN29),.WL(WL73));
sram_cell_6t_5 inst_cell_73_30 (.BL(BL30),.BLN(BLN30),.WL(WL73));
sram_cell_6t_5 inst_cell_73_31 (.BL(BL31),.BLN(BLN31),.WL(WL73));
sram_cell_6t_5 inst_cell_73_32 (.BL(BL32),.BLN(BLN32),.WL(WL73));
sram_cell_6t_5 inst_cell_73_33 (.BL(BL33),.BLN(BLN33),.WL(WL73));
sram_cell_6t_5 inst_cell_73_34 (.BL(BL34),.BLN(BLN34),.WL(WL73));
sram_cell_6t_5 inst_cell_73_35 (.BL(BL35),.BLN(BLN35),.WL(WL73));
sram_cell_6t_5 inst_cell_73_36 (.BL(BL36),.BLN(BLN36),.WL(WL73));
sram_cell_6t_5 inst_cell_73_37 (.BL(BL37),.BLN(BLN37),.WL(WL73));
sram_cell_6t_5 inst_cell_73_38 (.BL(BL38),.BLN(BLN38),.WL(WL73));
sram_cell_6t_5 inst_cell_73_39 (.BL(BL39),.BLN(BLN39),.WL(WL73));
sram_cell_6t_5 inst_cell_73_40 (.BL(BL40),.BLN(BLN40),.WL(WL73));
sram_cell_6t_5 inst_cell_73_41 (.BL(BL41),.BLN(BLN41),.WL(WL73));
sram_cell_6t_5 inst_cell_73_42 (.BL(BL42),.BLN(BLN42),.WL(WL73));
sram_cell_6t_5 inst_cell_73_43 (.BL(BL43),.BLN(BLN43),.WL(WL73));
sram_cell_6t_5 inst_cell_73_44 (.BL(BL44),.BLN(BLN44),.WL(WL73));
sram_cell_6t_5 inst_cell_73_45 (.BL(BL45),.BLN(BLN45),.WL(WL73));
sram_cell_6t_5 inst_cell_73_46 (.BL(BL46),.BLN(BLN46),.WL(WL73));
sram_cell_6t_5 inst_cell_73_47 (.BL(BL47),.BLN(BLN47),.WL(WL73));
sram_cell_6t_5 inst_cell_73_48 (.BL(BL48),.BLN(BLN48),.WL(WL73));
sram_cell_6t_5 inst_cell_73_49 (.BL(BL49),.BLN(BLN49),.WL(WL73));
sram_cell_6t_5 inst_cell_73_50 (.BL(BL50),.BLN(BLN50),.WL(WL73));
sram_cell_6t_5 inst_cell_73_51 (.BL(BL51),.BLN(BLN51),.WL(WL73));
sram_cell_6t_5 inst_cell_73_52 (.BL(BL52),.BLN(BLN52),.WL(WL73));
sram_cell_6t_5 inst_cell_73_53 (.BL(BL53),.BLN(BLN53),.WL(WL73));
sram_cell_6t_5 inst_cell_73_54 (.BL(BL54),.BLN(BLN54),.WL(WL73));
sram_cell_6t_5 inst_cell_73_55 (.BL(BL55),.BLN(BLN55),.WL(WL73));
sram_cell_6t_5 inst_cell_73_56 (.BL(BL56),.BLN(BLN56),.WL(WL73));
sram_cell_6t_5 inst_cell_73_57 (.BL(BL57),.BLN(BLN57),.WL(WL73));
sram_cell_6t_5 inst_cell_73_58 (.BL(BL58),.BLN(BLN58),.WL(WL73));
sram_cell_6t_5 inst_cell_73_59 (.BL(BL59),.BLN(BLN59),.WL(WL73));
sram_cell_6t_5 inst_cell_73_60 (.BL(BL60),.BLN(BLN60),.WL(WL73));
sram_cell_6t_5 inst_cell_73_61 (.BL(BL61),.BLN(BLN61),.WL(WL73));
sram_cell_6t_5 inst_cell_73_62 (.BL(BL62),.BLN(BLN62),.WL(WL73));
sram_cell_6t_5 inst_cell_73_63 (.BL(BL63),.BLN(BLN63),.WL(WL73));
sram_cell_6t_5 inst_cell_73_64 (.BL(BL64),.BLN(BLN64),.WL(WL73));
sram_cell_6t_5 inst_cell_73_65 (.BL(BL65),.BLN(BLN65),.WL(WL73));
sram_cell_6t_5 inst_cell_73_66 (.BL(BL66),.BLN(BLN66),.WL(WL73));
sram_cell_6t_5 inst_cell_73_67 (.BL(BL67),.BLN(BLN67),.WL(WL73));
sram_cell_6t_5 inst_cell_73_68 (.BL(BL68),.BLN(BLN68),.WL(WL73));
sram_cell_6t_5 inst_cell_73_69 (.BL(BL69),.BLN(BLN69),.WL(WL73));
sram_cell_6t_5 inst_cell_73_70 (.BL(BL70),.BLN(BLN70),.WL(WL73));
sram_cell_6t_5 inst_cell_73_71 (.BL(BL71),.BLN(BLN71),.WL(WL73));
sram_cell_6t_5 inst_cell_73_72 (.BL(BL72),.BLN(BLN72),.WL(WL73));
sram_cell_6t_5 inst_cell_73_73 (.BL(BL73),.BLN(BLN73),.WL(WL73));
sram_cell_6t_5 inst_cell_73_74 (.BL(BL74),.BLN(BLN74),.WL(WL73));
sram_cell_6t_5 inst_cell_73_75 (.BL(BL75),.BLN(BLN75),.WL(WL73));
sram_cell_6t_5 inst_cell_73_76 (.BL(BL76),.BLN(BLN76),.WL(WL73));
sram_cell_6t_5 inst_cell_73_77 (.BL(BL77),.BLN(BLN77),.WL(WL73));
sram_cell_6t_5 inst_cell_73_78 (.BL(BL78),.BLN(BLN78),.WL(WL73));
sram_cell_6t_5 inst_cell_73_79 (.BL(BL79),.BLN(BLN79),.WL(WL73));
sram_cell_6t_5 inst_cell_73_80 (.BL(BL80),.BLN(BLN80),.WL(WL73));
sram_cell_6t_5 inst_cell_73_81 (.BL(BL81),.BLN(BLN81),.WL(WL73));
sram_cell_6t_5 inst_cell_73_82 (.BL(BL82),.BLN(BLN82),.WL(WL73));
sram_cell_6t_5 inst_cell_73_83 (.BL(BL83),.BLN(BLN83),.WL(WL73));
sram_cell_6t_5 inst_cell_73_84 (.BL(BL84),.BLN(BLN84),.WL(WL73));
sram_cell_6t_5 inst_cell_73_85 (.BL(BL85),.BLN(BLN85),.WL(WL73));
sram_cell_6t_5 inst_cell_73_86 (.BL(BL86),.BLN(BLN86),.WL(WL73));
sram_cell_6t_5 inst_cell_73_87 (.BL(BL87),.BLN(BLN87),.WL(WL73));
sram_cell_6t_5 inst_cell_73_88 (.BL(BL88),.BLN(BLN88),.WL(WL73));
sram_cell_6t_5 inst_cell_73_89 (.BL(BL89),.BLN(BLN89),.WL(WL73));
sram_cell_6t_5 inst_cell_73_90 (.BL(BL90),.BLN(BLN90),.WL(WL73));
sram_cell_6t_5 inst_cell_73_91 (.BL(BL91),.BLN(BLN91),.WL(WL73));
sram_cell_6t_5 inst_cell_73_92 (.BL(BL92),.BLN(BLN92),.WL(WL73));
sram_cell_6t_5 inst_cell_73_93 (.BL(BL93),.BLN(BLN93),.WL(WL73));
sram_cell_6t_5 inst_cell_73_94 (.BL(BL94),.BLN(BLN94),.WL(WL73));
sram_cell_6t_5 inst_cell_73_95 (.BL(BL95),.BLN(BLN95),.WL(WL73));
sram_cell_6t_5 inst_cell_73_96 (.BL(BL96),.BLN(BLN96),.WL(WL73));
sram_cell_6t_5 inst_cell_73_97 (.BL(BL97),.BLN(BLN97),.WL(WL73));
sram_cell_6t_5 inst_cell_73_98 (.BL(BL98),.BLN(BLN98),.WL(WL73));
sram_cell_6t_5 inst_cell_73_99 (.BL(BL99),.BLN(BLN99),.WL(WL73));
sram_cell_6t_5 inst_cell_73_100 (.BL(BL100),.BLN(BLN100),.WL(WL73));
sram_cell_6t_5 inst_cell_73_101 (.BL(BL101),.BLN(BLN101),.WL(WL73));
sram_cell_6t_5 inst_cell_73_102 (.BL(BL102),.BLN(BLN102),.WL(WL73));
sram_cell_6t_5 inst_cell_73_103 (.BL(BL103),.BLN(BLN103),.WL(WL73));
sram_cell_6t_5 inst_cell_73_104 (.BL(BL104),.BLN(BLN104),.WL(WL73));
sram_cell_6t_5 inst_cell_73_105 (.BL(BL105),.BLN(BLN105),.WL(WL73));
sram_cell_6t_5 inst_cell_73_106 (.BL(BL106),.BLN(BLN106),.WL(WL73));
sram_cell_6t_5 inst_cell_73_107 (.BL(BL107),.BLN(BLN107),.WL(WL73));
sram_cell_6t_5 inst_cell_73_108 (.BL(BL108),.BLN(BLN108),.WL(WL73));
sram_cell_6t_5 inst_cell_73_109 (.BL(BL109),.BLN(BLN109),.WL(WL73));
sram_cell_6t_5 inst_cell_73_110 (.BL(BL110),.BLN(BLN110),.WL(WL73));
sram_cell_6t_5 inst_cell_73_111 (.BL(BL111),.BLN(BLN111),.WL(WL73));
sram_cell_6t_5 inst_cell_73_112 (.BL(BL112),.BLN(BLN112),.WL(WL73));
sram_cell_6t_5 inst_cell_73_113 (.BL(BL113),.BLN(BLN113),.WL(WL73));
sram_cell_6t_5 inst_cell_73_114 (.BL(BL114),.BLN(BLN114),.WL(WL73));
sram_cell_6t_5 inst_cell_73_115 (.BL(BL115),.BLN(BLN115),.WL(WL73));
sram_cell_6t_5 inst_cell_73_116 (.BL(BL116),.BLN(BLN116),.WL(WL73));
sram_cell_6t_5 inst_cell_73_117 (.BL(BL117),.BLN(BLN117),.WL(WL73));
sram_cell_6t_5 inst_cell_73_118 (.BL(BL118),.BLN(BLN118),.WL(WL73));
sram_cell_6t_5 inst_cell_73_119 (.BL(BL119),.BLN(BLN119),.WL(WL73));
sram_cell_6t_5 inst_cell_73_120 (.BL(BL120),.BLN(BLN120),.WL(WL73));
sram_cell_6t_5 inst_cell_73_121 (.BL(BL121),.BLN(BLN121),.WL(WL73));
sram_cell_6t_5 inst_cell_73_122 (.BL(BL122),.BLN(BLN122),.WL(WL73));
sram_cell_6t_5 inst_cell_73_123 (.BL(BL123),.BLN(BLN123),.WL(WL73));
sram_cell_6t_5 inst_cell_73_124 (.BL(BL124),.BLN(BLN124),.WL(WL73));
sram_cell_6t_5 inst_cell_73_125 (.BL(BL125),.BLN(BLN125),.WL(WL73));
sram_cell_6t_5 inst_cell_73_126 (.BL(BL126),.BLN(BLN126),.WL(WL73));
sram_cell_6t_5 inst_cell_73_127 (.BL(BL127),.BLN(BLN127),.WL(WL73));
sram_cell_6t_5 inst_cell_74_0 (.BL(BL0),.BLN(BLN0),.WL(WL74));
sram_cell_6t_5 inst_cell_74_1 (.BL(BL1),.BLN(BLN1),.WL(WL74));
sram_cell_6t_5 inst_cell_74_2 (.BL(BL2),.BLN(BLN2),.WL(WL74));
sram_cell_6t_5 inst_cell_74_3 (.BL(BL3),.BLN(BLN3),.WL(WL74));
sram_cell_6t_5 inst_cell_74_4 (.BL(BL4),.BLN(BLN4),.WL(WL74));
sram_cell_6t_5 inst_cell_74_5 (.BL(BL5),.BLN(BLN5),.WL(WL74));
sram_cell_6t_5 inst_cell_74_6 (.BL(BL6),.BLN(BLN6),.WL(WL74));
sram_cell_6t_5 inst_cell_74_7 (.BL(BL7),.BLN(BLN7),.WL(WL74));
sram_cell_6t_5 inst_cell_74_8 (.BL(BL8),.BLN(BLN8),.WL(WL74));
sram_cell_6t_5 inst_cell_74_9 (.BL(BL9),.BLN(BLN9),.WL(WL74));
sram_cell_6t_5 inst_cell_74_10 (.BL(BL10),.BLN(BLN10),.WL(WL74));
sram_cell_6t_5 inst_cell_74_11 (.BL(BL11),.BLN(BLN11),.WL(WL74));
sram_cell_6t_5 inst_cell_74_12 (.BL(BL12),.BLN(BLN12),.WL(WL74));
sram_cell_6t_5 inst_cell_74_13 (.BL(BL13),.BLN(BLN13),.WL(WL74));
sram_cell_6t_5 inst_cell_74_14 (.BL(BL14),.BLN(BLN14),.WL(WL74));
sram_cell_6t_5 inst_cell_74_15 (.BL(BL15),.BLN(BLN15),.WL(WL74));
sram_cell_6t_5 inst_cell_74_16 (.BL(BL16),.BLN(BLN16),.WL(WL74));
sram_cell_6t_5 inst_cell_74_17 (.BL(BL17),.BLN(BLN17),.WL(WL74));
sram_cell_6t_5 inst_cell_74_18 (.BL(BL18),.BLN(BLN18),.WL(WL74));
sram_cell_6t_5 inst_cell_74_19 (.BL(BL19),.BLN(BLN19),.WL(WL74));
sram_cell_6t_5 inst_cell_74_20 (.BL(BL20),.BLN(BLN20),.WL(WL74));
sram_cell_6t_5 inst_cell_74_21 (.BL(BL21),.BLN(BLN21),.WL(WL74));
sram_cell_6t_5 inst_cell_74_22 (.BL(BL22),.BLN(BLN22),.WL(WL74));
sram_cell_6t_5 inst_cell_74_23 (.BL(BL23),.BLN(BLN23),.WL(WL74));
sram_cell_6t_5 inst_cell_74_24 (.BL(BL24),.BLN(BLN24),.WL(WL74));
sram_cell_6t_5 inst_cell_74_25 (.BL(BL25),.BLN(BLN25),.WL(WL74));
sram_cell_6t_5 inst_cell_74_26 (.BL(BL26),.BLN(BLN26),.WL(WL74));
sram_cell_6t_5 inst_cell_74_27 (.BL(BL27),.BLN(BLN27),.WL(WL74));
sram_cell_6t_5 inst_cell_74_28 (.BL(BL28),.BLN(BLN28),.WL(WL74));
sram_cell_6t_5 inst_cell_74_29 (.BL(BL29),.BLN(BLN29),.WL(WL74));
sram_cell_6t_5 inst_cell_74_30 (.BL(BL30),.BLN(BLN30),.WL(WL74));
sram_cell_6t_5 inst_cell_74_31 (.BL(BL31),.BLN(BLN31),.WL(WL74));
sram_cell_6t_5 inst_cell_74_32 (.BL(BL32),.BLN(BLN32),.WL(WL74));
sram_cell_6t_5 inst_cell_74_33 (.BL(BL33),.BLN(BLN33),.WL(WL74));
sram_cell_6t_5 inst_cell_74_34 (.BL(BL34),.BLN(BLN34),.WL(WL74));
sram_cell_6t_5 inst_cell_74_35 (.BL(BL35),.BLN(BLN35),.WL(WL74));
sram_cell_6t_5 inst_cell_74_36 (.BL(BL36),.BLN(BLN36),.WL(WL74));
sram_cell_6t_5 inst_cell_74_37 (.BL(BL37),.BLN(BLN37),.WL(WL74));
sram_cell_6t_5 inst_cell_74_38 (.BL(BL38),.BLN(BLN38),.WL(WL74));
sram_cell_6t_5 inst_cell_74_39 (.BL(BL39),.BLN(BLN39),.WL(WL74));
sram_cell_6t_5 inst_cell_74_40 (.BL(BL40),.BLN(BLN40),.WL(WL74));
sram_cell_6t_5 inst_cell_74_41 (.BL(BL41),.BLN(BLN41),.WL(WL74));
sram_cell_6t_5 inst_cell_74_42 (.BL(BL42),.BLN(BLN42),.WL(WL74));
sram_cell_6t_5 inst_cell_74_43 (.BL(BL43),.BLN(BLN43),.WL(WL74));
sram_cell_6t_5 inst_cell_74_44 (.BL(BL44),.BLN(BLN44),.WL(WL74));
sram_cell_6t_5 inst_cell_74_45 (.BL(BL45),.BLN(BLN45),.WL(WL74));
sram_cell_6t_5 inst_cell_74_46 (.BL(BL46),.BLN(BLN46),.WL(WL74));
sram_cell_6t_5 inst_cell_74_47 (.BL(BL47),.BLN(BLN47),.WL(WL74));
sram_cell_6t_5 inst_cell_74_48 (.BL(BL48),.BLN(BLN48),.WL(WL74));
sram_cell_6t_5 inst_cell_74_49 (.BL(BL49),.BLN(BLN49),.WL(WL74));
sram_cell_6t_5 inst_cell_74_50 (.BL(BL50),.BLN(BLN50),.WL(WL74));
sram_cell_6t_5 inst_cell_74_51 (.BL(BL51),.BLN(BLN51),.WL(WL74));
sram_cell_6t_5 inst_cell_74_52 (.BL(BL52),.BLN(BLN52),.WL(WL74));
sram_cell_6t_5 inst_cell_74_53 (.BL(BL53),.BLN(BLN53),.WL(WL74));
sram_cell_6t_5 inst_cell_74_54 (.BL(BL54),.BLN(BLN54),.WL(WL74));
sram_cell_6t_5 inst_cell_74_55 (.BL(BL55),.BLN(BLN55),.WL(WL74));
sram_cell_6t_5 inst_cell_74_56 (.BL(BL56),.BLN(BLN56),.WL(WL74));
sram_cell_6t_5 inst_cell_74_57 (.BL(BL57),.BLN(BLN57),.WL(WL74));
sram_cell_6t_5 inst_cell_74_58 (.BL(BL58),.BLN(BLN58),.WL(WL74));
sram_cell_6t_5 inst_cell_74_59 (.BL(BL59),.BLN(BLN59),.WL(WL74));
sram_cell_6t_5 inst_cell_74_60 (.BL(BL60),.BLN(BLN60),.WL(WL74));
sram_cell_6t_5 inst_cell_74_61 (.BL(BL61),.BLN(BLN61),.WL(WL74));
sram_cell_6t_5 inst_cell_74_62 (.BL(BL62),.BLN(BLN62),.WL(WL74));
sram_cell_6t_5 inst_cell_74_63 (.BL(BL63),.BLN(BLN63),.WL(WL74));
sram_cell_6t_5 inst_cell_74_64 (.BL(BL64),.BLN(BLN64),.WL(WL74));
sram_cell_6t_5 inst_cell_74_65 (.BL(BL65),.BLN(BLN65),.WL(WL74));
sram_cell_6t_5 inst_cell_74_66 (.BL(BL66),.BLN(BLN66),.WL(WL74));
sram_cell_6t_5 inst_cell_74_67 (.BL(BL67),.BLN(BLN67),.WL(WL74));
sram_cell_6t_5 inst_cell_74_68 (.BL(BL68),.BLN(BLN68),.WL(WL74));
sram_cell_6t_5 inst_cell_74_69 (.BL(BL69),.BLN(BLN69),.WL(WL74));
sram_cell_6t_5 inst_cell_74_70 (.BL(BL70),.BLN(BLN70),.WL(WL74));
sram_cell_6t_5 inst_cell_74_71 (.BL(BL71),.BLN(BLN71),.WL(WL74));
sram_cell_6t_5 inst_cell_74_72 (.BL(BL72),.BLN(BLN72),.WL(WL74));
sram_cell_6t_5 inst_cell_74_73 (.BL(BL73),.BLN(BLN73),.WL(WL74));
sram_cell_6t_5 inst_cell_74_74 (.BL(BL74),.BLN(BLN74),.WL(WL74));
sram_cell_6t_5 inst_cell_74_75 (.BL(BL75),.BLN(BLN75),.WL(WL74));
sram_cell_6t_5 inst_cell_74_76 (.BL(BL76),.BLN(BLN76),.WL(WL74));
sram_cell_6t_5 inst_cell_74_77 (.BL(BL77),.BLN(BLN77),.WL(WL74));
sram_cell_6t_5 inst_cell_74_78 (.BL(BL78),.BLN(BLN78),.WL(WL74));
sram_cell_6t_5 inst_cell_74_79 (.BL(BL79),.BLN(BLN79),.WL(WL74));
sram_cell_6t_5 inst_cell_74_80 (.BL(BL80),.BLN(BLN80),.WL(WL74));
sram_cell_6t_5 inst_cell_74_81 (.BL(BL81),.BLN(BLN81),.WL(WL74));
sram_cell_6t_5 inst_cell_74_82 (.BL(BL82),.BLN(BLN82),.WL(WL74));
sram_cell_6t_5 inst_cell_74_83 (.BL(BL83),.BLN(BLN83),.WL(WL74));
sram_cell_6t_5 inst_cell_74_84 (.BL(BL84),.BLN(BLN84),.WL(WL74));
sram_cell_6t_5 inst_cell_74_85 (.BL(BL85),.BLN(BLN85),.WL(WL74));
sram_cell_6t_5 inst_cell_74_86 (.BL(BL86),.BLN(BLN86),.WL(WL74));
sram_cell_6t_5 inst_cell_74_87 (.BL(BL87),.BLN(BLN87),.WL(WL74));
sram_cell_6t_5 inst_cell_74_88 (.BL(BL88),.BLN(BLN88),.WL(WL74));
sram_cell_6t_5 inst_cell_74_89 (.BL(BL89),.BLN(BLN89),.WL(WL74));
sram_cell_6t_5 inst_cell_74_90 (.BL(BL90),.BLN(BLN90),.WL(WL74));
sram_cell_6t_5 inst_cell_74_91 (.BL(BL91),.BLN(BLN91),.WL(WL74));
sram_cell_6t_5 inst_cell_74_92 (.BL(BL92),.BLN(BLN92),.WL(WL74));
sram_cell_6t_5 inst_cell_74_93 (.BL(BL93),.BLN(BLN93),.WL(WL74));
sram_cell_6t_5 inst_cell_74_94 (.BL(BL94),.BLN(BLN94),.WL(WL74));
sram_cell_6t_5 inst_cell_74_95 (.BL(BL95),.BLN(BLN95),.WL(WL74));
sram_cell_6t_5 inst_cell_74_96 (.BL(BL96),.BLN(BLN96),.WL(WL74));
sram_cell_6t_5 inst_cell_74_97 (.BL(BL97),.BLN(BLN97),.WL(WL74));
sram_cell_6t_5 inst_cell_74_98 (.BL(BL98),.BLN(BLN98),.WL(WL74));
sram_cell_6t_5 inst_cell_74_99 (.BL(BL99),.BLN(BLN99),.WL(WL74));
sram_cell_6t_5 inst_cell_74_100 (.BL(BL100),.BLN(BLN100),.WL(WL74));
sram_cell_6t_5 inst_cell_74_101 (.BL(BL101),.BLN(BLN101),.WL(WL74));
sram_cell_6t_5 inst_cell_74_102 (.BL(BL102),.BLN(BLN102),.WL(WL74));
sram_cell_6t_5 inst_cell_74_103 (.BL(BL103),.BLN(BLN103),.WL(WL74));
sram_cell_6t_5 inst_cell_74_104 (.BL(BL104),.BLN(BLN104),.WL(WL74));
sram_cell_6t_5 inst_cell_74_105 (.BL(BL105),.BLN(BLN105),.WL(WL74));
sram_cell_6t_5 inst_cell_74_106 (.BL(BL106),.BLN(BLN106),.WL(WL74));
sram_cell_6t_5 inst_cell_74_107 (.BL(BL107),.BLN(BLN107),.WL(WL74));
sram_cell_6t_5 inst_cell_74_108 (.BL(BL108),.BLN(BLN108),.WL(WL74));
sram_cell_6t_5 inst_cell_74_109 (.BL(BL109),.BLN(BLN109),.WL(WL74));
sram_cell_6t_5 inst_cell_74_110 (.BL(BL110),.BLN(BLN110),.WL(WL74));
sram_cell_6t_5 inst_cell_74_111 (.BL(BL111),.BLN(BLN111),.WL(WL74));
sram_cell_6t_5 inst_cell_74_112 (.BL(BL112),.BLN(BLN112),.WL(WL74));
sram_cell_6t_5 inst_cell_74_113 (.BL(BL113),.BLN(BLN113),.WL(WL74));
sram_cell_6t_5 inst_cell_74_114 (.BL(BL114),.BLN(BLN114),.WL(WL74));
sram_cell_6t_5 inst_cell_74_115 (.BL(BL115),.BLN(BLN115),.WL(WL74));
sram_cell_6t_5 inst_cell_74_116 (.BL(BL116),.BLN(BLN116),.WL(WL74));
sram_cell_6t_5 inst_cell_74_117 (.BL(BL117),.BLN(BLN117),.WL(WL74));
sram_cell_6t_5 inst_cell_74_118 (.BL(BL118),.BLN(BLN118),.WL(WL74));
sram_cell_6t_5 inst_cell_74_119 (.BL(BL119),.BLN(BLN119),.WL(WL74));
sram_cell_6t_5 inst_cell_74_120 (.BL(BL120),.BLN(BLN120),.WL(WL74));
sram_cell_6t_5 inst_cell_74_121 (.BL(BL121),.BLN(BLN121),.WL(WL74));
sram_cell_6t_5 inst_cell_74_122 (.BL(BL122),.BLN(BLN122),.WL(WL74));
sram_cell_6t_5 inst_cell_74_123 (.BL(BL123),.BLN(BLN123),.WL(WL74));
sram_cell_6t_5 inst_cell_74_124 (.BL(BL124),.BLN(BLN124),.WL(WL74));
sram_cell_6t_5 inst_cell_74_125 (.BL(BL125),.BLN(BLN125),.WL(WL74));
sram_cell_6t_5 inst_cell_74_126 (.BL(BL126),.BLN(BLN126),.WL(WL74));
sram_cell_6t_5 inst_cell_74_127 (.BL(BL127),.BLN(BLN127),.WL(WL74));
sram_cell_6t_5 inst_cell_75_0 (.BL(BL0),.BLN(BLN0),.WL(WL75));
sram_cell_6t_5 inst_cell_75_1 (.BL(BL1),.BLN(BLN1),.WL(WL75));
sram_cell_6t_5 inst_cell_75_2 (.BL(BL2),.BLN(BLN2),.WL(WL75));
sram_cell_6t_5 inst_cell_75_3 (.BL(BL3),.BLN(BLN3),.WL(WL75));
sram_cell_6t_5 inst_cell_75_4 (.BL(BL4),.BLN(BLN4),.WL(WL75));
sram_cell_6t_5 inst_cell_75_5 (.BL(BL5),.BLN(BLN5),.WL(WL75));
sram_cell_6t_5 inst_cell_75_6 (.BL(BL6),.BLN(BLN6),.WL(WL75));
sram_cell_6t_5 inst_cell_75_7 (.BL(BL7),.BLN(BLN7),.WL(WL75));
sram_cell_6t_5 inst_cell_75_8 (.BL(BL8),.BLN(BLN8),.WL(WL75));
sram_cell_6t_5 inst_cell_75_9 (.BL(BL9),.BLN(BLN9),.WL(WL75));
sram_cell_6t_5 inst_cell_75_10 (.BL(BL10),.BLN(BLN10),.WL(WL75));
sram_cell_6t_5 inst_cell_75_11 (.BL(BL11),.BLN(BLN11),.WL(WL75));
sram_cell_6t_5 inst_cell_75_12 (.BL(BL12),.BLN(BLN12),.WL(WL75));
sram_cell_6t_5 inst_cell_75_13 (.BL(BL13),.BLN(BLN13),.WL(WL75));
sram_cell_6t_5 inst_cell_75_14 (.BL(BL14),.BLN(BLN14),.WL(WL75));
sram_cell_6t_5 inst_cell_75_15 (.BL(BL15),.BLN(BLN15),.WL(WL75));
sram_cell_6t_5 inst_cell_75_16 (.BL(BL16),.BLN(BLN16),.WL(WL75));
sram_cell_6t_5 inst_cell_75_17 (.BL(BL17),.BLN(BLN17),.WL(WL75));
sram_cell_6t_5 inst_cell_75_18 (.BL(BL18),.BLN(BLN18),.WL(WL75));
sram_cell_6t_5 inst_cell_75_19 (.BL(BL19),.BLN(BLN19),.WL(WL75));
sram_cell_6t_5 inst_cell_75_20 (.BL(BL20),.BLN(BLN20),.WL(WL75));
sram_cell_6t_5 inst_cell_75_21 (.BL(BL21),.BLN(BLN21),.WL(WL75));
sram_cell_6t_5 inst_cell_75_22 (.BL(BL22),.BLN(BLN22),.WL(WL75));
sram_cell_6t_5 inst_cell_75_23 (.BL(BL23),.BLN(BLN23),.WL(WL75));
sram_cell_6t_5 inst_cell_75_24 (.BL(BL24),.BLN(BLN24),.WL(WL75));
sram_cell_6t_5 inst_cell_75_25 (.BL(BL25),.BLN(BLN25),.WL(WL75));
sram_cell_6t_5 inst_cell_75_26 (.BL(BL26),.BLN(BLN26),.WL(WL75));
sram_cell_6t_5 inst_cell_75_27 (.BL(BL27),.BLN(BLN27),.WL(WL75));
sram_cell_6t_5 inst_cell_75_28 (.BL(BL28),.BLN(BLN28),.WL(WL75));
sram_cell_6t_5 inst_cell_75_29 (.BL(BL29),.BLN(BLN29),.WL(WL75));
sram_cell_6t_5 inst_cell_75_30 (.BL(BL30),.BLN(BLN30),.WL(WL75));
sram_cell_6t_5 inst_cell_75_31 (.BL(BL31),.BLN(BLN31),.WL(WL75));
sram_cell_6t_5 inst_cell_75_32 (.BL(BL32),.BLN(BLN32),.WL(WL75));
sram_cell_6t_5 inst_cell_75_33 (.BL(BL33),.BLN(BLN33),.WL(WL75));
sram_cell_6t_5 inst_cell_75_34 (.BL(BL34),.BLN(BLN34),.WL(WL75));
sram_cell_6t_5 inst_cell_75_35 (.BL(BL35),.BLN(BLN35),.WL(WL75));
sram_cell_6t_5 inst_cell_75_36 (.BL(BL36),.BLN(BLN36),.WL(WL75));
sram_cell_6t_5 inst_cell_75_37 (.BL(BL37),.BLN(BLN37),.WL(WL75));
sram_cell_6t_5 inst_cell_75_38 (.BL(BL38),.BLN(BLN38),.WL(WL75));
sram_cell_6t_5 inst_cell_75_39 (.BL(BL39),.BLN(BLN39),.WL(WL75));
sram_cell_6t_5 inst_cell_75_40 (.BL(BL40),.BLN(BLN40),.WL(WL75));
sram_cell_6t_5 inst_cell_75_41 (.BL(BL41),.BLN(BLN41),.WL(WL75));
sram_cell_6t_5 inst_cell_75_42 (.BL(BL42),.BLN(BLN42),.WL(WL75));
sram_cell_6t_5 inst_cell_75_43 (.BL(BL43),.BLN(BLN43),.WL(WL75));
sram_cell_6t_5 inst_cell_75_44 (.BL(BL44),.BLN(BLN44),.WL(WL75));
sram_cell_6t_5 inst_cell_75_45 (.BL(BL45),.BLN(BLN45),.WL(WL75));
sram_cell_6t_5 inst_cell_75_46 (.BL(BL46),.BLN(BLN46),.WL(WL75));
sram_cell_6t_5 inst_cell_75_47 (.BL(BL47),.BLN(BLN47),.WL(WL75));
sram_cell_6t_5 inst_cell_75_48 (.BL(BL48),.BLN(BLN48),.WL(WL75));
sram_cell_6t_5 inst_cell_75_49 (.BL(BL49),.BLN(BLN49),.WL(WL75));
sram_cell_6t_5 inst_cell_75_50 (.BL(BL50),.BLN(BLN50),.WL(WL75));
sram_cell_6t_5 inst_cell_75_51 (.BL(BL51),.BLN(BLN51),.WL(WL75));
sram_cell_6t_5 inst_cell_75_52 (.BL(BL52),.BLN(BLN52),.WL(WL75));
sram_cell_6t_5 inst_cell_75_53 (.BL(BL53),.BLN(BLN53),.WL(WL75));
sram_cell_6t_5 inst_cell_75_54 (.BL(BL54),.BLN(BLN54),.WL(WL75));
sram_cell_6t_5 inst_cell_75_55 (.BL(BL55),.BLN(BLN55),.WL(WL75));
sram_cell_6t_5 inst_cell_75_56 (.BL(BL56),.BLN(BLN56),.WL(WL75));
sram_cell_6t_5 inst_cell_75_57 (.BL(BL57),.BLN(BLN57),.WL(WL75));
sram_cell_6t_5 inst_cell_75_58 (.BL(BL58),.BLN(BLN58),.WL(WL75));
sram_cell_6t_5 inst_cell_75_59 (.BL(BL59),.BLN(BLN59),.WL(WL75));
sram_cell_6t_5 inst_cell_75_60 (.BL(BL60),.BLN(BLN60),.WL(WL75));
sram_cell_6t_5 inst_cell_75_61 (.BL(BL61),.BLN(BLN61),.WL(WL75));
sram_cell_6t_5 inst_cell_75_62 (.BL(BL62),.BLN(BLN62),.WL(WL75));
sram_cell_6t_5 inst_cell_75_63 (.BL(BL63),.BLN(BLN63),.WL(WL75));
sram_cell_6t_5 inst_cell_75_64 (.BL(BL64),.BLN(BLN64),.WL(WL75));
sram_cell_6t_5 inst_cell_75_65 (.BL(BL65),.BLN(BLN65),.WL(WL75));
sram_cell_6t_5 inst_cell_75_66 (.BL(BL66),.BLN(BLN66),.WL(WL75));
sram_cell_6t_5 inst_cell_75_67 (.BL(BL67),.BLN(BLN67),.WL(WL75));
sram_cell_6t_5 inst_cell_75_68 (.BL(BL68),.BLN(BLN68),.WL(WL75));
sram_cell_6t_5 inst_cell_75_69 (.BL(BL69),.BLN(BLN69),.WL(WL75));
sram_cell_6t_5 inst_cell_75_70 (.BL(BL70),.BLN(BLN70),.WL(WL75));
sram_cell_6t_5 inst_cell_75_71 (.BL(BL71),.BLN(BLN71),.WL(WL75));
sram_cell_6t_5 inst_cell_75_72 (.BL(BL72),.BLN(BLN72),.WL(WL75));
sram_cell_6t_5 inst_cell_75_73 (.BL(BL73),.BLN(BLN73),.WL(WL75));
sram_cell_6t_5 inst_cell_75_74 (.BL(BL74),.BLN(BLN74),.WL(WL75));
sram_cell_6t_5 inst_cell_75_75 (.BL(BL75),.BLN(BLN75),.WL(WL75));
sram_cell_6t_5 inst_cell_75_76 (.BL(BL76),.BLN(BLN76),.WL(WL75));
sram_cell_6t_5 inst_cell_75_77 (.BL(BL77),.BLN(BLN77),.WL(WL75));
sram_cell_6t_5 inst_cell_75_78 (.BL(BL78),.BLN(BLN78),.WL(WL75));
sram_cell_6t_5 inst_cell_75_79 (.BL(BL79),.BLN(BLN79),.WL(WL75));
sram_cell_6t_5 inst_cell_75_80 (.BL(BL80),.BLN(BLN80),.WL(WL75));
sram_cell_6t_5 inst_cell_75_81 (.BL(BL81),.BLN(BLN81),.WL(WL75));
sram_cell_6t_5 inst_cell_75_82 (.BL(BL82),.BLN(BLN82),.WL(WL75));
sram_cell_6t_5 inst_cell_75_83 (.BL(BL83),.BLN(BLN83),.WL(WL75));
sram_cell_6t_5 inst_cell_75_84 (.BL(BL84),.BLN(BLN84),.WL(WL75));
sram_cell_6t_5 inst_cell_75_85 (.BL(BL85),.BLN(BLN85),.WL(WL75));
sram_cell_6t_5 inst_cell_75_86 (.BL(BL86),.BLN(BLN86),.WL(WL75));
sram_cell_6t_5 inst_cell_75_87 (.BL(BL87),.BLN(BLN87),.WL(WL75));
sram_cell_6t_5 inst_cell_75_88 (.BL(BL88),.BLN(BLN88),.WL(WL75));
sram_cell_6t_5 inst_cell_75_89 (.BL(BL89),.BLN(BLN89),.WL(WL75));
sram_cell_6t_5 inst_cell_75_90 (.BL(BL90),.BLN(BLN90),.WL(WL75));
sram_cell_6t_5 inst_cell_75_91 (.BL(BL91),.BLN(BLN91),.WL(WL75));
sram_cell_6t_5 inst_cell_75_92 (.BL(BL92),.BLN(BLN92),.WL(WL75));
sram_cell_6t_5 inst_cell_75_93 (.BL(BL93),.BLN(BLN93),.WL(WL75));
sram_cell_6t_5 inst_cell_75_94 (.BL(BL94),.BLN(BLN94),.WL(WL75));
sram_cell_6t_5 inst_cell_75_95 (.BL(BL95),.BLN(BLN95),.WL(WL75));
sram_cell_6t_5 inst_cell_75_96 (.BL(BL96),.BLN(BLN96),.WL(WL75));
sram_cell_6t_5 inst_cell_75_97 (.BL(BL97),.BLN(BLN97),.WL(WL75));
sram_cell_6t_5 inst_cell_75_98 (.BL(BL98),.BLN(BLN98),.WL(WL75));
sram_cell_6t_5 inst_cell_75_99 (.BL(BL99),.BLN(BLN99),.WL(WL75));
sram_cell_6t_5 inst_cell_75_100 (.BL(BL100),.BLN(BLN100),.WL(WL75));
sram_cell_6t_5 inst_cell_75_101 (.BL(BL101),.BLN(BLN101),.WL(WL75));
sram_cell_6t_5 inst_cell_75_102 (.BL(BL102),.BLN(BLN102),.WL(WL75));
sram_cell_6t_5 inst_cell_75_103 (.BL(BL103),.BLN(BLN103),.WL(WL75));
sram_cell_6t_5 inst_cell_75_104 (.BL(BL104),.BLN(BLN104),.WL(WL75));
sram_cell_6t_5 inst_cell_75_105 (.BL(BL105),.BLN(BLN105),.WL(WL75));
sram_cell_6t_5 inst_cell_75_106 (.BL(BL106),.BLN(BLN106),.WL(WL75));
sram_cell_6t_5 inst_cell_75_107 (.BL(BL107),.BLN(BLN107),.WL(WL75));
sram_cell_6t_5 inst_cell_75_108 (.BL(BL108),.BLN(BLN108),.WL(WL75));
sram_cell_6t_5 inst_cell_75_109 (.BL(BL109),.BLN(BLN109),.WL(WL75));
sram_cell_6t_5 inst_cell_75_110 (.BL(BL110),.BLN(BLN110),.WL(WL75));
sram_cell_6t_5 inst_cell_75_111 (.BL(BL111),.BLN(BLN111),.WL(WL75));
sram_cell_6t_5 inst_cell_75_112 (.BL(BL112),.BLN(BLN112),.WL(WL75));
sram_cell_6t_5 inst_cell_75_113 (.BL(BL113),.BLN(BLN113),.WL(WL75));
sram_cell_6t_5 inst_cell_75_114 (.BL(BL114),.BLN(BLN114),.WL(WL75));
sram_cell_6t_5 inst_cell_75_115 (.BL(BL115),.BLN(BLN115),.WL(WL75));
sram_cell_6t_5 inst_cell_75_116 (.BL(BL116),.BLN(BLN116),.WL(WL75));
sram_cell_6t_5 inst_cell_75_117 (.BL(BL117),.BLN(BLN117),.WL(WL75));
sram_cell_6t_5 inst_cell_75_118 (.BL(BL118),.BLN(BLN118),.WL(WL75));
sram_cell_6t_5 inst_cell_75_119 (.BL(BL119),.BLN(BLN119),.WL(WL75));
sram_cell_6t_5 inst_cell_75_120 (.BL(BL120),.BLN(BLN120),.WL(WL75));
sram_cell_6t_5 inst_cell_75_121 (.BL(BL121),.BLN(BLN121),.WL(WL75));
sram_cell_6t_5 inst_cell_75_122 (.BL(BL122),.BLN(BLN122),.WL(WL75));
sram_cell_6t_5 inst_cell_75_123 (.BL(BL123),.BLN(BLN123),.WL(WL75));
sram_cell_6t_5 inst_cell_75_124 (.BL(BL124),.BLN(BLN124),.WL(WL75));
sram_cell_6t_5 inst_cell_75_125 (.BL(BL125),.BLN(BLN125),.WL(WL75));
sram_cell_6t_5 inst_cell_75_126 (.BL(BL126),.BLN(BLN126),.WL(WL75));
sram_cell_6t_5 inst_cell_75_127 (.BL(BL127),.BLN(BLN127),.WL(WL75));
sram_cell_6t_5 inst_cell_76_0 (.BL(BL0),.BLN(BLN0),.WL(WL76));
sram_cell_6t_5 inst_cell_76_1 (.BL(BL1),.BLN(BLN1),.WL(WL76));
sram_cell_6t_5 inst_cell_76_2 (.BL(BL2),.BLN(BLN2),.WL(WL76));
sram_cell_6t_5 inst_cell_76_3 (.BL(BL3),.BLN(BLN3),.WL(WL76));
sram_cell_6t_5 inst_cell_76_4 (.BL(BL4),.BLN(BLN4),.WL(WL76));
sram_cell_6t_5 inst_cell_76_5 (.BL(BL5),.BLN(BLN5),.WL(WL76));
sram_cell_6t_5 inst_cell_76_6 (.BL(BL6),.BLN(BLN6),.WL(WL76));
sram_cell_6t_5 inst_cell_76_7 (.BL(BL7),.BLN(BLN7),.WL(WL76));
sram_cell_6t_5 inst_cell_76_8 (.BL(BL8),.BLN(BLN8),.WL(WL76));
sram_cell_6t_5 inst_cell_76_9 (.BL(BL9),.BLN(BLN9),.WL(WL76));
sram_cell_6t_5 inst_cell_76_10 (.BL(BL10),.BLN(BLN10),.WL(WL76));
sram_cell_6t_5 inst_cell_76_11 (.BL(BL11),.BLN(BLN11),.WL(WL76));
sram_cell_6t_5 inst_cell_76_12 (.BL(BL12),.BLN(BLN12),.WL(WL76));
sram_cell_6t_5 inst_cell_76_13 (.BL(BL13),.BLN(BLN13),.WL(WL76));
sram_cell_6t_5 inst_cell_76_14 (.BL(BL14),.BLN(BLN14),.WL(WL76));
sram_cell_6t_5 inst_cell_76_15 (.BL(BL15),.BLN(BLN15),.WL(WL76));
sram_cell_6t_5 inst_cell_76_16 (.BL(BL16),.BLN(BLN16),.WL(WL76));
sram_cell_6t_5 inst_cell_76_17 (.BL(BL17),.BLN(BLN17),.WL(WL76));
sram_cell_6t_5 inst_cell_76_18 (.BL(BL18),.BLN(BLN18),.WL(WL76));
sram_cell_6t_5 inst_cell_76_19 (.BL(BL19),.BLN(BLN19),.WL(WL76));
sram_cell_6t_5 inst_cell_76_20 (.BL(BL20),.BLN(BLN20),.WL(WL76));
sram_cell_6t_5 inst_cell_76_21 (.BL(BL21),.BLN(BLN21),.WL(WL76));
sram_cell_6t_5 inst_cell_76_22 (.BL(BL22),.BLN(BLN22),.WL(WL76));
sram_cell_6t_5 inst_cell_76_23 (.BL(BL23),.BLN(BLN23),.WL(WL76));
sram_cell_6t_5 inst_cell_76_24 (.BL(BL24),.BLN(BLN24),.WL(WL76));
sram_cell_6t_5 inst_cell_76_25 (.BL(BL25),.BLN(BLN25),.WL(WL76));
sram_cell_6t_5 inst_cell_76_26 (.BL(BL26),.BLN(BLN26),.WL(WL76));
sram_cell_6t_5 inst_cell_76_27 (.BL(BL27),.BLN(BLN27),.WL(WL76));
sram_cell_6t_5 inst_cell_76_28 (.BL(BL28),.BLN(BLN28),.WL(WL76));
sram_cell_6t_5 inst_cell_76_29 (.BL(BL29),.BLN(BLN29),.WL(WL76));
sram_cell_6t_5 inst_cell_76_30 (.BL(BL30),.BLN(BLN30),.WL(WL76));
sram_cell_6t_5 inst_cell_76_31 (.BL(BL31),.BLN(BLN31),.WL(WL76));
sram_cell_6t_5 inst_cell_76_32 (.BL(BL32),.BLN(BLN32),.WL(WL76));
sram_cell_6t_5 inst_cell_76_33 (.BL(BL33),.BLN(BLN33),.WL(WL76));
sram_cell_6t_5 inst_cell_76_34 (.BL(BL34),.BLN(BLN34),.WL(WL76));
sram_cell_6t_5 inst_cell_76_35 (.BL(BL35),.BLN(BLN35),.WL(WL76));
sram_cell_6t_5 inst_cell_76_36 (.BL(BL36),.BLN(BLN36),.WL(WL76));
sram_cell_6t_5 inst_cell_76_37 (.BL(BL37),.BLN(BLN37),.WL(WL76));
sram_cell_6t_5 inst_cell_76_38 (.BL(BL38),.BLN(BLN38),.WL(WL76));
sram_cell_6t_5 inst_cell_76_39 (.BL(BL39),.BLN(BLN39),.WL(WL76));
sram_cell_6t_5 inst_cell_76_40 (.BL(BL40),.BLN(BLN40),.WL(WL76));
sram_cell_6t_5 inst_cell_76_41 (.BL(BL41),.BLN(BLN41),.WL(WL76));
sram_cell_6t_5 inst_cell_76_42 (.BL(BL42),.BLN(BLN42),.WL(WL76));
sram_cell_6t_5 inst_cell_76_43 (.BL(BL43),.BLN(BLN43),.WL(WL76));
sram_cell_6t_5 inst_cell_76_44 (.BL(BL44),.BLN(BLN44),.WL(WL76));
sram_cell_6t_5 inst_cell_76_45 (.BL(BL45),.BLN(BLN45),.WL(WL76));
sram_cell_6t_5 inst_cell_76_46 (.BL(BL46),.BLN(BLN46),.WL(WL76));
sram_cell_6t_5 inst_cell_76_47 (.BL(BL47),.BLN(BLN47),.WL(WL76));
sram_cell_6t_5 inst_cell_76_48 (.BL(BL48),.BLN(BLN48),.WL(WL76));
sram_cell_6t_5 inst_cell_76_49 (.BL(BL49),.BLN(BLN49),.WL(WL76));
sram_cell_6t_5 inst_cell_76_50 (.BL(BL50),.BLN(BLN50),.WL(WL76));
sram_cell_6t_5 inst_cell_76_51 (.BL(BL51),.BLN(BLN51),.WL(WL76));
sram_cell_6t_5 inst_cell_76_52 (.BL(BL52),.BLN(BLN52),.WL(WL76));
sram_cell_6t_5 inst_cell_76_53 (.BL(BL53),.BLN(BLN53),.WL(WL76));
sram_cell_6t_5 inst_cell_76_54 (.BL(BL54),.BLN(BLN54),.WL(WL76));
sram_cell_6t_5 inst_cell_76_55 (.BL(BL55),.BLN(BLN55),.WL(WL76));
sram_cell_6t_5 inst_cell_76_56 (.BL(BL56),.BLN(BLN56),.WL(WL76));
sram_cell_6t_5 inst_cell_76_57 (.BL(BL57),.BLN(BLN57),.WL(WL76));
sram_cell_6t_5 inst_cell_76_58 (.BL(BL58),.BLN(BLN58),.WL(WL76));
sram_cell_6t_5 inst_cell_76_59 (.BL(BL59),.BLN(BLN59),.WL(WL76));
sram_cell_6t_5 inst_cell_76_60 (.BL(BL60),.BLN(BLN60),.WL(WL76));
sram_cell_6t_5 inst_cell_76_61 (.BL(BL61),.BLN(BLN61),.WL(WL76));
sram_cell_6t_5 inst_cell_76_62 (.BL(BL62),.BLN(BLN62),.WL(WL76));
sram_cell_6t_5 inst_cell_76_63 (.BL(BL63),.BLN(BLN63),.WL(WL76));
sram_cell_6t_5 inst_cell_76_64 (.BL(BL64),.BLN(BLN64),.WL(WL76));
sram_cell_6t_5 inst_cell_76_65 (.BL(BL65),.BLN(BLN65),.WL(WL76));
sram_cell_6t_5 inst_cell_76_66 (.BL(BL66),.BLN(BLN66),.WL(WL76));
sram_cell_6t_5 inst_cell_76_67 (.BL(BL67),.BLN(BLN67),.WL(WL76));
sram_cell_6t_5 inst_cell_76_68 (.BL(BL68),.BLN(BLN68),.WL(WL76));
sram_cell_6t_5 inst_cell_76_69 (.BL(BL69),.BLN(BLN69),.WL(WL76));
sram_cell_6t_5 inst_cell_76_70 (.BL(BL70),.BLN(BLN70),.WL(WL76));
sram_cell_6t_5 inst_cell_76_71 (.BL(BL71),.BLN(BLN71),.WL(WL76));
sram_cell_6t_5 inst_cell_76_72 (.BL(BL72),.BLN(BLN72),.WL(WL76));
sram_cell_6t_5 inst_cell_76_73 (.BL(BL73),.BLN(BLN73),.WL(WL76));
sram_cell_6t_5 inst_cell_76_74 (.BL(BL74),.BLN(BLN74),.WL(WL76));
sram_cell_6t_5 inst_cell_76_75 (.BL(BL75),.BLN(BLN75),.WL(WL76));
sram_cell_6t_5 inst_cell_76_76 (.BL(BL76),.BLN(BLN76),.WL(WL76));
sram_cell_6t_5 inst_cell_76_77 (.BL(BL77),.BLN(BLN77),.WL(WL76));
sram_cell_6t_5 inst_cell_76_78 (.BL(BL78),.BLN(BLN78),.WL(WL76));
sram_cell_6t_5 inst_cell_76_79 (.BL(BL79),.BLN(BLN79),.WL(WL76));
sram_cell_6t_5 inst_cell_76_80 (.BL(BL80),.BLN(BLN80),.WL(WL76));
sram_cell_6t_5 inst_cell_76_81 (.BL(BL81),.BLN(BLN81),.WL(WL76));
sram_cell_6t_5 inst_cell_76_82 (.BL(BL82),.BLN(BLN82),.WL(WL76));
sram_cell_6t_5 inst_cell_76_83 (.BL(BL83),.BLN(BLN83),.WL(WL76));
sram_cell_6t_5 inst_cell_76_84 (.BL(BL84),.BLN(BLN84),.WL(WL76));
sram_cell_6t_5 inst_cell_76_85 (.BL(BL85),.BLN(BLN85),.WL(WL76));
sram_cell_6t_5 inst_cell_76_86 (.BL(BL86),.BLN(BLN86),.WL(WL76));
sram_cell_6t_5 inst_cell_76_87 (.BL(BL87),.BLN(BLN87),.WL(WL76));
sram_cell_6t_5 inst_cell_76_88 (.BL(BL88),.BLN(BLN88),.WL(WL76));
sram_cell_6t_5 inst_cell_76_89 (.BL(BL89),.BLN(BLN89),.WL(WL76));
sram_cell_6t_5 inst_cell_76_90 (.BL(BL90),.BLN(BLN90),.WL(WL76));
sram_cell_6t_5 inst_cell_76_91 (.BL(BL91),.BLN(BLN91),.WL(WL76));
sram_cell_6t_5 inst_cell_76_92 (.BL(BL92),.BLN(BLN92),.WL(WL76));
sram_cell_6t_5 inst_cell_76_93 (.BL(BL93),.BLN(BLN93),.WL(WL76));
sram_cell_6t_5 inst_cell_76_94 (.BL(BL94),.BLN(BLN94),.WL(WL76));
sram_cell_6t_5 inst_cell_76_95 (.BL(BL95),.BLN(BLN95),.WL(WL76));
sram_cell_6t_5 inst_cell_76_96 (.BL(BL96),.BLN(BLN96),.WL(WL76));
sram_cell_6t_5 inst_cell_76_97 (.BL(BL97),.BLN(BLN97),.WL(WL76));
sram_cell_6t_5 inst_cell_76_98 (.BL(BL98),.BLN(BLN98),.WL(WL76));
sram_cell_6t_5 inst_cell_76_99 (.BL(BL99),.BLN(BLN99),.WL(WL76));
sram_cell_6t_5 inst_cell_76_100 (.BL(BL100),.BLN(BLN100),.WL(WL76));
sram_cell_6t_5 inst_cell_76_101 (.BL(BL101),.BLN(BLN101),.WL(WL76));
sram_cell_6t_5 inst_cell_76_102 (.BL(BL102),.BLN(BLN102),.WL(WL76));
sram_cell_6t_5 inst_cell_76_103 (.BL(BL103),.BLN(BLN103),.WL(WL76));
sram_cell_6t_5 inst_cell_76_104 (.BL(BL104),.BLN(BLN104),.WL(WL76));
sram_cell_6t_5 inst_cell_76_105 (.BL(BL105),.BLN(BLN105),.WL(WL76));
sram_cell_6t_5 inst_cell_76_106 (.BL(BL106),.BLN(BLN106),.WL(WL76));
sram_cell_6t_5 inst_cell_76_107 (.BL(BL107),.BLN(BLN107),.WL(WL76));
sram_cell_6t_5 inst_cell_76_108 (.BL(BL108),.BLN(BLN108),.WL(WL76));
sram_cell_6t_5 inst_cell_76_109 (.BL(BL109),.BLN(BLN109),.WL(WL76));
sram_cell_6t_5 inst_cell_76_110 (.BL(BL110),.BLN(BLN110),.WL(WL76));
sram_cell_6t_5 inst_cell_76_111 (.BL(BL111),.BLN(BLN111),.WL(WL76));
sram_cell_6t_5 inst_cell_76_112 (.BL(BL112),.BLN(BLN112),.WL(WL76));
sram_cell_6t_5 inst_cell_76_113 (.BL(BL113),.BLN(BLN113),.WL(WL76));
sram_cell_6t_5 inst_cell_76_114 (.BL(BL114),.BLN(BLN114),.WL(WL76));
sram_cell_6t_5 inst_cell_76_115 (.BL(BL115),.BLN(BLN115),.WL(WL76));
sram_cell_6t_5 inst_cell_76_116 (.BL(BL116),.BLN(BLN116),.WL(WL76));
sram_cell_6t_5 inst_cell_76_117 (.BL(BL117),.BLN(BLN117),.WL(WL76));
sram_cell_6t_5 inst_cell_76_118 (.BL(BL118),.BLN(BLN118),.WL(WL76));
sram_cell_6t_5 inst_cell_76_119 (.BL(BL119),.BLN(BLN119),.WL(WL76));
sram_cell_6t_5 inst_cell_76_120 (.BL(BL120),.BLN(BLN120),.WL(WL76));
sram_cell_6t_5 inst_cell_76_121 (.BL(BL121),.BLN(BLN121),.WL(WL76));
sram_cell_6t_5 inst_cell_76_122 (.BL(BL122),.BLN(BLN122),.WL(WL76));
sram_cell_6t_5 inst_cell_76_123 (.BL(BL123),.BLN(BLN123),.WL(WL76));
sram_cell_6t_5 inst_cell_76_124 (.BL(BL124),.BLN(BLN124),.WL(WL76));
sram_cell_6t_5 inst_cell_76_125 (.BL(BL125),.BLN(BLN125),.WL(WL76));
sram_cell_6t_5 inst_cell_76_126 (.BL(BL126),.BLN(BLN126),.WL(WL76));
sram_cell_6t_5 inst_cell_76_127 (.BL(BL127),.BLN(BLN127),.WL(WL76));
sram_cell_6t_5 inst_cell_77_0 (.BL(BL0),.BLN(BLN0),.WL(WL77));
sram_cell_6t_5 inst_cell_77_1 (.BL(BL1),.BLN(BLN1),.WL(WL77));
sram_cell_6t_5 inst_cell_77_2 (.BL(BL2),.BLN(BLN2),.WL(WL77));
sram_cell_6t_5 inst_cell_77_3 (.BL(BL3),.BLN(BLN3),.WL(WL77));
sram_cell_6t_5 inst_cell_77_4 (.BL(BL4),.BLN(BLN4),.WL(WL77));
sram_cell_6t_5 inst_cell_77_5 (.BL(BL5),.BLN(BLN5),.WL(WL77));
sram_cell_6t_5 inst_cell_77_6 (.BL(BL6),.BLN(BLN6),.WL(WL77));
sram_cell_6t_5 inst_cell_77_7 (.BL(BL7),.BLN(BLN7),.WL(WL77));
sram_cell_6t_5 inst_cell_77_8 (.BL(BL8),.BLN(BLN8),.WL(WL77));
sram_cell_6t_5 inst_cell_77_9 (.BL(BL9),.BLN(BLN9),.WL(WL77));
sram_cell_6t_5 inst_cell_77_10 (.BL(BL10),.BLN(BLN10),.WL(WL77));
sram_cell_6t_5 inst_cell_77_11 (.BL(BL11),.BLN(BLN11),.WL(WL77));
sram_cell_6t_5 inst_cell_77_12 (.BL(BL12),.BLN(BLN12),.WL(WL77));
sram_cell_6t_5 inst_cell_77_13 (.BL(BL13),.BLN(BLN13),.WL(WL77));
sram_cell_6t_5 inst_cell_77_14 (.BL(BL14),.BLN(BLN14),.WL(WL77));
sram_cell_6t_5 inst_cell_77_15 (.BL(BL15),.BLN(BLN15),.WL(WL77));
sram_cell_6t_5 inst_cell_77_16 (.BL(BL16),.BLN(BLN16),.WL(WL77));
sram_cell_6t_5 inst_cell_77_17 (.BL(BL17),.BLN(BLN17),.WL(WL77));
sram_cell_6t_5 inst_cell_77_18 (.BL(BL18),.BLN(BLN18),.WL(WL77));
sram_cell_6t_5 inst_cell_77_19 (.BL(BL19),.BLN(BLN19),.WL(WL77));
sram_cell_6t_5 inst_cell_77_20 (.BL(BL20),.BLN(BLN20),.WL(WL77));
sram_cell_6t_5 inst_cell_77_21 (.BL(BL21),.BLN(BLN21),.WL(WL77));
sram_cell_6t_5 inst_cell_77_22 (.BL(BL22),.BLN(BLN22),.WL(WL77));
sram_cell_6t_5 inst_cell_77_23 (.BL(BL23),.BLN(BLN23),.WL(WL77));
sram_cell_6t_5 inst_cell_77_24 (.BL(BL24),.BLN(BLN24),.WL(WL77));
sram_cell_6t_5 inst_cell_77_25 (.BL(BL25),.BLN(BLN25),.WL(WL77));
sram_cell_6t_5 inst_cell_77_26 (.BL(BL26),.BLN(BLN26),.WL(WL77));
sram_cell_6t_5 inst_cell_77_27 (.BL(BL27),.BLN(BLN27),.WL(WL77));
sram_cell_6t_5 inst_cell_77_28 (.BL(BL28),.BLN(BLN28),.WL(WL77));
sram_cell_6t_5 inst_cell_77_29 (.BL(BL29),.BLN(BLN29),.WL(WL77));
sram_cell_6t_5 inst_cell_77_30 (.BL(BL30),.BLN(BLN30),.WL(WL77));
sram_cell_6t_5 inst_cell_77_31 (.BL(BL31),.BLN(BLN31),.WL(WL77));
sram_cell_6t_5 inst_cell_77_32 (.BL(BL32),.BLN(BLN32),.WL(WL77));
sram_cell_6t_5 inst_cell_77_33 (.BL(BL33),.BLN(BLN33),.WL(WL77));
sram_cell_6t_5 inst_cell_77_34 (.BL(BL34),.BLN(BLN34),.WL(WL77));
sram_cell_6t_5 inst_cell_77_35 (.BL(BL35),.BLN(BLN35),.WL(WL77));
sram_cell_6t_5 inst_cell_77_36 (.BL(BL36),.BLN(BLN36),.WL(WL77));
sram_cell_6t_5 inst_cell_77_37 (.BL(BL37),.BLN(BLN37),.WL(WL77));
sram_cell_6t_5 inst_cell_77_38 (.BL(BL38),.BLN(BLN38),.WL(WL77));
sram_cell_6t_5 inst_cell_77_39 (.BL(BL39),.BLN(BLN39),.WL(WL77));
sram_cell_6t_5 inst_cell_77_40 (.BL(BL40),.BLN(BLN40),.WL(WL77));
sram_cell_6t_5 inst_cell_77_41 (.BL(BL41),.BLN(BLN41),.WL(WL77));
sram_cell_6t_5 inst_cell_77_42 (.BL(BL42),.BLN(BLN42),.WL(WL77));
sram_cell_6t_5 inst_cell_77_43 (.BL(BL43),.BLN(BLN43),.WL(WL77));
sram_cell_6t_5 inst_cell_77_44 (.BL(BL44),.BLN(BLN44),.WL(WL77));
sram_cell_6t_5 inst_cell_77_45 (.BL(BL45),.BLN(BLN45),.WL(WL77));
sram_cell_6t_5 inst_cell_77_46 (.BL(BL46),.BLN(BLN46),.WL(WL77));
sram_cell_6t_5 inst_cell_77_47 (.BL(BL47),.BLN(BLN47),.WL(WL77));
sram_cell_6t_5 inst_cell_77_48 (.BL(BL48),.BLN(BLN48),.WL(WL77));
sram_cell_6t_5 inst_cell_77_49 (.BL(BL49),.BLN(BLN49),.WL(WL77));
sram_cell_6t_5 inst_cell_77_50 (.BL(BL50),.BLN(BLN50),.WL(WL77));
sram_cell_6t_5 inst_cell_77_51 (.BL(BL51),.BLN(BLN51),.WL(WL77));
sram_cell_6t_5 inst_cell_77_52 (.BL(BL52),.BLN(BLN52),.WL(WL77));
sram_cell_6t_5 inst_cell_77_53 (.BL(BL53),.BLN(BLN53),.WL(WL77));
sram_cell_6t_5 inst_cell_77_54 (.BL(BL54),.BLN(BLN54),.WL(WL77));
sram_cell_6t_5 inst_cell_77_55 (.BL(BL55),.BLN(BLN55),.WL(WL77));
sram_cell_6t_5 inst_cell_77_56 (.BL(BL56),.BLN(BLN56),.WL(WL77));
sram_cell_6t_5 inst_cell_77_57 (.BL(BL57),.BLN(BLN57),.WL(WL77));
sram_cell_6t_5 inst_cell_77_58 (.BL(BL58),.BLN(BLN58),.WL(WL77));
sram_cell_6t_5 inst_cell_77_59 (.BL(BL59),.BLN(BLN59),.WL(WL77));
sram_cell_6t_5 inst_cell_77_60 (.BL(BL60),.BLN(BLN60),.WL(WL77));
sram_cell_6t_5 inst_cell_77_61 (.BL(BL61),.BLN(BLN61),.WL(WL77));
sram_cell_6t_5 inst_cell_77_62 (.BL(BL62),.BLN(BLN62),.WL(WL77));
sram_cell_6t_5 inst_cell_77_63 (.BL(BL63),.BLN(BLN63),.WL(WL77));
sram_cell_6t_5 inst_cell_77_64 (.BL(BL64),.BLN(BLN64),.WL(WL77));
sram_cell_6t_5 inst_cell_77_65 (.BL(BL65),.BLN(BLN65),.WL(WL77));
sram_cell_6t_5 inst_cell_77_66 (.BL(BL66),.BLN(BLN66),.WL(WL77));
sram_cell_6t_5 inst_cell_77_67 (.BL(BL67),.BLN(BLN67),.WL(WL77));
sram_cell_6t_5 inst_cell_77_68 (.BL(BL68),.BLN(BLN68),.WL(WL77));
sram_cell_6t_5 inst_cell_77_69 (.BL(BL69),.BLN(BLN69),.WL(WL77));
sram_cell_6t_5 inst_cell_77_70 (.BL(BL70),.BLN(BLN70),.WL(WL77));
sram_cell_6t_5 inst_cell_77_71 (.BL(BL71),.BLN(BLN71),.WL(WL77));
sram_cell_6t_5 inst_cell_77_72 (.BL(BL72),.BLN(BLN72),.WL(WL77));
sram_cell_6t_5 inst_cell_77_73 (.BL(BL73),.BLN(BLN73),.WL(WL77));
sram_cell_6t_5 inst_cell_77_74 (.BL(BL74),.BLN(BLN74),.WL(WL77));
sram_cell_6t_5 inst_cell_77_75 (.BL(BL75),.BLN(BLN75),.WL(WL77));
sram_cell_6t_5 inst_cell_77_76 (.BL(BL76),.BLN(BLN76),.WL(WL77));
sram_cell_6t_5 inst_cell_77_77 (.BL(BL77),.BLN(BLN77),.WL(WL77));
sram_cell_6t_5 inst_cell_77_78 (.BL(BL78),.BLN(BLN78),.WL(WL77));
sram_cell_6t_5 inst_cell_77_79 (.BL(BL79),.BLN(BLN79),.WL(WL77));
sram_cell_6t_5 inst_cell_77_80 (.BL(BL80),.BLN(BLN80),.WL(WL77));
sram_cell_6t_5 inst_cell_77_81 (.BL(BL81),.BLN(BLN81),.WL(WL77));
sram_cell_6t_5 inst_cell_77_82 (.BL(BL82),.BLN(BLN82),.WL(WL77));
sram_cell_6t_5 inst_cell_77_83 (.BL(BL83),.BLN(BLN83),.WL(WL77));
sram_cell_6t_5 inst_cell_77_84 (.BL(BL84),.BLN(BLN84),.WL(WL77));
sram_cell_6t_5 inst_cell_77_85 (.BL(BL85),.BLN(BLN85),.WL(WL77));
sram_cell_6t_5 inst_cell_77_86 (.BL(BL86),.BLN(BLN86),.WL(WL77));
sram_cell_6t_5 inst_cell_77_87 (.BL(BL87),.BLN(BLN87),.WL(WL77));
sram_cell_6t_5 inst_cell_77_88 (.BL(BL88),.BLN(BLN88),.WL(WL77));
sram_cell_6t_5 inst_cell_77_89 (.BL(BL89),.BLN(BLN89),.WL(WL77));
sram_cell_6t_5 inst_cell_77_90 (.BL(BL90),.BLN(BLN90),.WL(WL77));
sram_cell_6t_5 inst_cell_77_91 (.BL(BL91),.BLN(BLN91),.WL(WL77));
sram_cell_6t_5 inst_cell_77_92 (.BL(BL92),.BLN(BLN92),.WL(WL77));
sram_cell_6t_5 inst_cell_77_93 (.BL(BL93),.BLN(BLN93),.WL(WL77));
sram_cell_6t_5 inst_cell_77_94 (.BL(BL94),.BLN(BLN94),.WL(WL77));
sram_cell_6t_5 inst_cell_77_95 (.BL(BL95),.BLN(BLN95),.WL(WL77));
sram_cell_6t_5 inst_cell_77_96 (.BL(BL96),.BLN(BLN96),.WL(WL77));
sram_cell_6t_5 inst_cell_77_97 (.BL(BL97),.BLN(BLN97),.WL(WL77));
sram_cell_6t_5 inst_cell_77_98 (.BL(BL98),.BLN(BLN98),.WL(WL77));
sram_cell_6t_5 inst_cell_77_99 (.BL(BL99),.BLN(BLN99),.WL(WL77));
sram_cell_6t_5 inst_cell_77_100 (.BL(BL100),.BLN(BLN100),.WL(WL77));
sram_cell_6t_5 inst_cell_77_101 (.BL(BL101),.BLN(BLN101),.WL(WL77));
sram_cell_6t_5 inst_cell_77_102 (.BL(BL102),.BLN(BLN102),.WL(WL77));
sram_cell_6t_5 inst_cell_77_103 (.BL(BL103),.BLN(BLN103),.WL(WL77));
sram_cell_6t_5 inst_cell_77_104 (.BL(BL104),.BLN(BLN104),.WL(WL77));
sram_cell_6t_5 inst_cell_77_105 (.BL(BL105),.BLN(BLN105),.WL(WL77));
sram_cell_6t_5 inst_cell_77_106 (.BL(BL106),.BLN(BLN106),.WL(WL77));
sram_cell_6t_5 inst_cell_77_107 (.BL(BL107),.BLN(BLN107),.WL(WL77));
sram_cell_6t_5 inst_cell_77_108 (.BL(BL108),.BLN(BLN108),.WL(WL77));
sram_cell_6t_5 inst_cell_77_109 (.BL(BL109),.BLN(BLN109),.WL(WL77));
sram_cell_6t_5 inst_cell_77_110 (.BL(BL110),.BLN(BLN110),.WL(WL77));
sram_cell_6t_5 inst_cell_77_111 (.BL(BL111),.BLN(BLN111),.WL(WL77));
sram_cell_6t_5 inst_cell_77_112 (.BL(BL112),.BLN(BLN112),.WL(WL77));
sram_cell_6t_5 inst_cell_77_113 (.BL(BL113),.BLN(BLN113),.WL(WL77));
sram_cell_6t_5 inst_cell_77_114 (.BL(BL114),.BLN(BLN114),.WL(WL77));
sram_cell_6t_5 inst_cell_77_115 (.BL(BL115),.BLN(BLN115),.WL(WL77));
sram_cell_6t_5 inst_cell_77_116 (.BL(BL116),.BLN(BLN116),.WL(WL77));
sram_cell_6t_5 inst_cell_77_117 (.BL(BL117),.BLN(BLN117),.WL(WL77));
sram_cell_6t_5 inst_cell_77_118 (.BL(BL118),.BLN(BLN118),.WL(WL77));
sram_cell_6t_5 inst_cell_77_119 (.BL(BL119),.BLN(BLN119),.WL(WL77));
sram_cell_6t_5 inst_cell_77_120 (.BL(BL120),.BLN(BLN120),.WL(WL77));
sram_cell_6t_5 inst_cell_77_121 (.BL(BL121),.BLN(BLN121),.WL(WL77));
sram_cell_6t_5 inst_cell_77_122 (.BL(BL122),.BLN(BLN122),.WL(WL77));
sram_cell_6t_5 inst_cell_77_123 (.BL(BL123),.BLN(BLN123),.WL(WL77));
sram_cell_6t_5 inst_cell_77_124 (.BL(BL124),.BLN(BLN124),.WL(WL77));
sram_cell_6t_5 inst_cell_77_125 (.BL(BL125),.BLN(BLN125),.WL(WL77));
sram_cell_6t_5 inst_cell_77_126 (.BL(BL126),.BLN(BLN126),.WL(WL77));
sram_cell_6t_5 inst_cell_77_127 (.BL(BL127),.BLN(BLN127),.WL(WL77));
sram_cell_6t_5 inst_cell_78_0 (.BL(BL0),.BLN(BLN0),.WL(WL78));
sram_cell_6t_5 inst_cell_78_1 (.BL(BL1),.BLN(BLN1),.WL(WL78));
sram_cell_6t_5 inst_cell_78_2 (.BL(BL2),.BLN(BLN2),.WL(WL78));
sram_cell_6t_5 inst_cell_78_3 (.BL(BL3),.BLN(BLN3),.WL(WL78));
sram_cell_6t_5 inst_cell_78_4 (.BL(BL4),.BLN(BLN4),.WL(WL78));
sram_cell_6t_5 inst_cell_78_5 (.BL(BL5),.BLN(BLN5),.WL(WL78));
sram_cell_6t_5 inst_cell_78_6 (.BL(BL6),.BLN(BLN6),.WL(WL78));
sram_cell_6t_5 inst_cell_78_7 (.BL(BL7),.BLN(BLN7),.WL(WL78));
sram_cell_6t_5 inst_cell_78_8 (.BL(BL8),.BLN(BLN8),.WL(WL78));
sram_cell_6t_5 inst_cell_78_9 (.BL(BL9),.BLN(BLN9),.WL(WL78));
sram_cell_6t_5 inst_cell_78_10 (.BL(BL10),.BLN(BLN10),.WL(WL78));
sram_cell_6t_5 inst_cell_78_11 (.BL(BL11),.BLN(BLN11),.WL(WL78));
sram_cell_6t_5 inst_cell_78_12 (.BL(BL12),.BLN(BLN12),.WL(WL78));
sram_cell_6t_5 inst_cell_78_13 (.BL(BL13),.BLN(BLN13),.WL(WL78));
sram_cell_6t_5 inst_cell_78_14 (.BL(BL14),.BLN(BLN14),.WL(WL78));
sram_cell_6t_5 inst_cell_78_15 (.BL(BL15),.BLN(BLN15),.WL(WL78));
sram_cell_6t_5 inst_cell_78_16 (.BL(BL16),.BLN(BLN16),.WL(WL78));
sram_cell_6t_5 inst_cell_78_17 (.BL(BL17),.BLN(BLN17),.WL(WL78));
sram_cell_6t_5 inst_cell_78_18 (.BL(BL18),.BLN(BLN18),.WL(WL78));
sram_cell_6t_5 inst_cell_78_19 (.BL(BL19),.BLN(BLN19),.WL(WL78));
sram_cell_6t_5 inst_cell_78_20 (.BL(BL20),.BLN(BLN20),.WL(WL78));
sram_cell_6t_5 inst_cell_78_21 (.BL(BL21),.BLN(BLN21),.WL(WL78));
sram_cell_6t_5 inst_cell_78_22 (.BL(BL22),.BLN(BLN22),.WL(WL78));
sram_cell_6t_5 inst_cell_78_23 (.BL(BL23),.BLN(BLN23),.WL(WL78));
sram_cell_6t_5 inst_cell_78_24 (.BL(BL24),.BLN(BLN24),.WL(WL78));
sram_cell_6t_5 inst_cell_78_25 (.BL(BL25),.BLN(BLN25),.WL(WL78));
sram_cell_6t_5 inst_cell_78_26 (.BL(BL26),.BLN(BLN26),.WL(WL78));
sram_cell_6t_5 inst_cell_78_27 (.BL(BL27),.BLN(BLN27),.WL(WL78));
sram_cell_6t_5 inst_cell_78_28 (.BL(BL28),.BLN(BLN28),.WL(WL78));
sram_cell_6t_5 inst_cell_78_29 (.BL(BL29),.BLN(BLN29),.WL(WL78));
sram_cell_6t_5 inst_cell_78_30 (.BL(BL30),.BLN(BLN30),.WL(WL78));
sram_cell_6t_5 inst_cell_78_31 (.BL(BL31),.BLN(BLN31),.WL(WL78));
sram_cell_6t_5 inst_cell_78_32 (.BL(BL32),.BLN(BLN32),.WL(WL78));
sram_cell_6t_5 inst_cell_78_33 (.BL(BL33),.BLN(BLN33),.WL(WL78));
sram_cell_6t_5 inst_cell_78_34 (.BL(BL34),.BLN(BLN34),.WL(WL78));
sram_cell_6t_5 inst_cell_78_35 (.BL(BL35),.BLN(BLN35),.WL(WL78));
sram_cell_6t_5 inst_cell_78_36 (.BL(BL36),.BLN(BLN36),.WL(WL78));
sram_cell_6t_5 inst_cell_78_37 (.BL(BL37),.BLN(BLN37),.WL(WL78));
sram_cell_6t_5 inst_cell_78_38 (.BL(BL38),.BLN(BLN38),.WL(WL78));
sram_cell_6t_5 inst_cell_78_39 (.BL(BL39),.BLN(BLN39),.WL(WL78));
sram_cell_6t_5 inst_cell_78_40 (.BL(BL40),.BLN(BLN40),.WL(WL78));
sram_cell_6t_5 inst_cell_78_41 (.BL(BL41),.BLN(BLN41),.WL(WL78));
sram_cell_6t_5 inst_cell_78_42 (.BL(BL42),.BLN(BLN42),.WL(WL78));
sram_cell_6t_5 inst_cell_78_43 (.BL(BL43),.BLN(BLN43),.WL(WL78));
sram_cell_6t_5 inst_cell_78_44 (.BL(BL44),.BLN(BLN44),.WL(WL78));
sram_cell_6t_5 inst_cell_78_45 (.BL(BL45),.BLN(BLN45),.WL(WL78));
sram_cell_6t_5 inst_cell_78_46 (.BL(BL46),.BLN(BLN46),.WL(WL78));
sram_cell_6t_5 inst_cell_78_47 (.BL(BL47),.BLN(BLN47),.WL(WL78));
sram_cell_6t_5 inst_cell_78_48 (.BL(BL48),.BLN(BLN48),.WL(WL78));
sram_cell_6t_5 inst_cell_78_49 (.BL(BL49),.BLN(BLN49),.WL(WL78));
sram_cell_6t_5 inst_cell_78_50 (.BL(BL50),.BLN(BLN50),.WL(WL78));
sram_cell_6t_5 inst_cell_78_51 (.BL(BL51),.BLN(BLN51),.WL(WL78));
sram_cell_6t_5 inst_cell_78_52 (.BL(BL52),.BLN(BLN52),.WL(WL78));
sram_cell_6t_5 inst_cell_78_53 (.BL(BL53),.BLN(BLN53),.WL(WL78));
sram_cell_6t_5 inst_cell_78_54 (.BL(BL54),.BLN(BLN54),.WL(WL78));
sram_cell_6t_5 inst_cell_78_55 (.BL(BL55),.BLN(BLN55),.WL(WL78));
sram_cell_6t_5 inst_cell_78_56 (.BL(BL56),.BLN(BLN56),.WL(WL78));
sram_cell_6t_5 inst_cell_78_57 (.BL(BL57),.BLN(BLN57),.WL(WL78));
sram_cell_6t_5 inst_cell_78_58 (.BL(BL58),.BLN(BLN58),.WL(WL78));
sram_cell_6t_5 inst_cell_78_59 (.BL(BL59),.BLN(BLN59),.WL(WL78));
sram_cell_6t_5 inst_cell_78_60 (.BL(BL60),.BLN(BLN60),.WL(WL78));
sram_cell_6t_5 inst_cell_78_61 (.BL(BL61),.BLN(BLN61),.WL(WL78));
sram_cell_6t_5 inst_cell_78_62 (.BL(BL62),.BLN(BLN62),.WL(WL78));
sram_cell_6t_5 inst_cell_78_63 (.BL(BL63),.BLN(BLN63),.WL(WL78));
sram_cell_6t_5 inst_cell_78_64 (.BL(BL64),.BLN(BLN64),.WL(WL78));
sram_cell_6t_5 inst_cell_78_65 (.BL(BL65),.BLN(BLN65),.WL(WL78));
sram_cell_6t_5 inst_cell_78_66 (.BL(BL66),.BLN(BLN66),.WL(WL78));
sram_cell_6t_5 inst_cell_78_67 (.BL(BL67),.BLN(BLN67),.WL(WL78));
sram_cell_6t_5 inst_cell_78_68 (.BL(BL68),.BLN(BLN68),.WL(WL78));
sram_cell_6t_5 inst_cell_78_69 (.BL(BL69),.BLN(BLN69),.WL(WL78));
sram_cell_6t_5 inst_cell_78_70 (.BL(BL70),.BLN(BLN70),.WL(WL78));
sram_cell_6t_5 inst_cell_78_71 (.BL(BL71),.BLN(BLN71),.WL(WL78));
sram_cell_6t_5 inst_cell_78_72 (.BL(BL72),.BLN(BLN72),.WL(WL78));
sram_cell_6t_5 inst_cell_78_73 (.BL(BL73),.BLN(BLN73),.WL(WL78));
sram_cell_6t_5 inst_cell_78_74 (.BL(BL74),.BLN(BLN74),.WL(WL78));
sram_cell_6t_5 inst_cell_78_75 (.BL(BL75),.BLN(BLN75),.WL(WL78));
sram_cell_6t_5 inst_cell_78_76 (.BL(BL76),.BLN(BLN76),.WL(WL78));
sram_cell_6t_5 inst_cell_78_77 (.BL(BL77),.BLN(BLN77),.WL(WL78));
sram_cell_6t_5 inst_cell_78_78 (.BL(BL78),.BLN(BLN78),.WL(WL78));
sram_cell_6t_5 inst_cell_78_79 (.BL(BL79),.BLN(BLN79),.WL(WL78));
sram_cell_6t_5 inst_cell_78_80 (.BL(BL80),.BLN(BLN80),.WL(WL78));
sram_cell_6t_5 inst_cell_78_81 (.BL(BL81),.BLN(BLN81),.WL(WL78));
sram_cell_6t_5 inst_cell_78_82 (.BL(BL82),.BLN(BLN82),.WL(WL78));
sram_cell_6t_5 inst_cell_78_83 (.BL(BL83),.BLN(BLN83),.WL(WL78));
sram_cell_6t_5 inst_cell_78_84 (.BL(BL84),.BLN(BLN84),.WL(WL78));
sram_cell_6t_5 inst_cell_78_85 (.BL(BL85),.BLN(BLN85),.WL(WL78));
sram_cell_6t_5 inst_cell_78_86 (.BL(BL86),.BLN(BLN86),.WL(WL78));
sram_cell_6t_5 inst_cell_78_87 (.BL(BL87),.BLN(BLN87),.WL(WL78));
sram_cell_6t_5 inst_cell_78_88 (.BL(BL88),.BLN(BLN88),.WL(WL78));
sram_cell_6t_5 inst_cell_78_89 (.BL(BL89),.BLN(BLN89),.WL(WL78));
sram_cell_6t_5 inst_cell_78_90 (.BL(BL90),.BLN(BLN90),.WL(WL78));
sram_cell_6t_5 inst_cell_78_91 (.BL(BL91),.BLN(BLN91),.WL(WL78));
sram_cell_6t_5 inst_cell_78_92 (.BL(BL92),.BLN(BLN92),.WL(WL78));
sram_cell_6t_5 inst_cell_78_93 (.BL(BL93),.BLN(BLN93),.WL(WL78));
sram_cell_6t_5 inst_cell_78_94 (.BL(BL94),.BLN(BLN94),.WL(WL78));
sram_cell_6t_5 inst_cell_78_95 (.BL(BL95),.BLN(BLN95),.WL(WL78));
sram_cell_6t_5 inst_cell_78_96 (.BL(BL96),.BLN(BLN96),.WL(WL78));
sram_cell_6t_5 inst_cell_78_97 (.BL(BL97),.BLN(BLN97),.WL(WL78));
sram_cell_6t_5 inst_cell_78_98 (.BL(BL98),.BLN(BLN98),.WL(WL78));
sram_cell_6t_5 inst_cell_78_99 (.BL(BL99),.BLN(BLN99),.WL(WL78));
sram_cell_6t_5 inst_cell_78_100 (.BL(BL100),.BLN(BLN100),.WL(WL78));
sram_cell_6t_5 inst_cell_78_101 (.BL(BL101),.BLN(BLN101),.WL(WL78));
sram_cell_6t_5 inst_cell_78_102 (.BL(BL102),.BLN(BLN102),.WL(WL78));
sram_cell_6t_5 inst_cell_78_103 (.BL(BL103),.BLN(BLN103),.WL(WL78));
sram_cell_6t_5 inst_cell_78_104 (.BL(BL104),.BLN(BLN104),.WL(WL78));
sram_cell_6t_5 inst_cell_78_105 (.BL(BL105),.BLN(BLN105),.WL(WL78));
sram_cell_6t_5 inst_cell_78_106 (.BL(BL106),.BLN(BLN106),.WL(WL78));
sram_cell_6t_5 inst_cell_78_107 (.BL(BL107),.BLN(BLN107),.WL(WL78));
sram_cell_6t_5 inst_cell_78_108 (.BL(BL108),.BLN(BLN108),.WL(WL78));
sram_cell_6t_5 inst_cell_78_109 (.BL(BL109),.BLN(BLN109),.WL(WL78));
sram_cell_6t_5 inst_cell_78_110 (.BL(BL110),.BLN(BLN110),.WL(WL78));
sram_cell_6t_5 inst_cell_78_111 (.BL(BL111),.BLN(BLN111),.WL(WL78));
sram_cell_6t_5 inst_cell_78_112 (.BL(BL112),.BLN(BLN112),.WL(WL78));
sram_cell_6t_5 inst_cell_78_113 (.BL(BL113),.BLN(BLN113),.WL(WL78));
sram_cell_6t_5 inst_cell_78_114 (.BL(BL114),.BLN(BLN114),.WL(WL78));
sram_cell_6t_5 inst_cell_78_115 (.BL(BL115),.BLN(BLN115),.WL(WL78));
sram_cell_6t_5 inst_cell_78_116 (.BL(BL116),.BLN(BLN116),.WL(WL78));
sram_cell_6t_5 inst_cell_78_117 (.BL(BL117),.BLN(BLN117),.WL(WL78));
sram_cell_6t_5 inst_cell_78_118 (.BL(BL118),.BLN(BLN118),.WL(WL78));
sram_cell_6t_5 inst_cell_78_119 (.BL(BL119),.BLN(BLN119),.WL(WL78));
sram_cell_6t_5 inst_cell_78_120 (.BL(BL120),.BLN(BLN120),.WL(WL78));
sram_cell_6t_5 inst_cell_78_121 (.BL(BL121),.BLN(BLN121),.WL(WL78));
sram_cell_6t_5 inst_cell_78_122 (.BL(BL122),.BLN(BLN122),.WL(WL78));
sram_cell_6t_5 inst_cell_78_123 (.BL(BL123),.BLN(BLN123),.WL(WL78));
sram_cell_6t_5 inst_cell_78_124 (.BL(BL124),.BLN(BLN124),.WL(WL78));
sram_cell_6t_5 inst_cell_78_125 (.BL(BL125),.BLN(BLN125),.WL(WL78));
sram_cell_6t_5 inst_cell_78_126 (.BL(BL126),.BLN(BLN126),.WL(WL78));
sram_cell_6t_5 inst_cell_78_127 (.BL(BL127),.BLN(BLN127),.WL(WL78));
sram_cell_6t_5 inst_cell_79_0 (.BL(BL0),.BLN(BLN0),.WL(WL79));
sram_cell_6t_5 inst_cell_79_1 (.BL(BL1),.BLN(BLN1),.WL(WL79));
sram_cell_6t_5 inst_cell_79_2 (.BL(BL2),.BLN(BLN2),.WL(WL79));
sram_cell_6t_5 inst_cell_79_3 (.BL(BL3),.BLN(BLN3),.WL(WL79));
sram_cell_6t_5 inst_cell_79_4 (.BL(BL4),.BLN(BLN4),.WL(WL79));
sram_cell_6t_5 inst_cell_79_5 (.BL(BL5),.BLN(BLN5),.WL(WL79));
sram_cell_6t_5 inst_cell_79_6 (.BL(BL6),.BLN(BLN6),.WL(WL79));
sram_cell_6t_5 inst_cell_79_7 (.BL(BL7),.BLN(BLN7),.WL(WL79));
sram_cell_6t_5 inst_cell_79_8 (.BL(BL8),.BLN(BLN8),.WL(WL79));
sram_cell_6t_5 inst_cell_79_9 (.BL(BL9),.BLN(BLN9),.WL(WL79));
sram_cell_6t_5 inst_cell_79_10 (.BL(BL10),.BLN(BLN10),.WL(WL79));
sram_cell_6t_5 inst_cell_79_11 (.BL(BL11),.BLN(BLN11),.WL(WL79));
sram_cell_6t_5 inst_cell_79_12 (.BL(BL12),.BLN(BLN12),.WL(WL79));
sram_cell_6t_5 inst_cell_79_13 (.BL(BL13),.BLN(BLN13),.WL(WL79));
sram_cell_6t_5 inst_cell_79_14 (.BL(BL14),.BLN(BLN14),.WL(WL79));
sram_cell_6t_5 inst_cell_79_15 (.BL(BL15),.BLN(BLN15),.WL(WL79));
sram_cell_6t_5 inst_cell_79_16 (.BL(BL16),.BLN(BLN16),.WL(WL79));
sram_cell_6t_5 inst_cell_79_17 (.BL(BL17),.BLN(BLN17),.WL(WL79));
sram_cell_6t_5 inst_cell_79_18 (.BL(BL18),.BLN(BLN18),.WL(WL79));
sram_cell_6t_5 inst_cell_79_19 (.BL(BL19),.BLN(BLN19),.WL(WL79));
sram_cell_6t_5 inst_cell_79_20 (.BL(BL20),.BLN(BLN20),.WL(WL79));
sram_cell_6t_5 inst_cell_79_21 (.BL(BL21),.BLN(BLN21),.WL(WL79));
sram_cell_6t_5 inst_cell_79_22 (.BL(BL22),.BLN(BLN22),.WL(WL79));
sram_cell_6t_5 inst_cell_79_23 (.BL(BL23),.BLN(BLN23),.WL(WL79));
sram_cell_6t_5 inst_cell_79_24 (.BL(BL24),.BLN(BLN24),.WL(WL79));
sram_cell_6t_5 inst_cell_79_25 (.BL(BL25),.BLN(BLN25),.WL(WL79));
sram_cell_6t_5 inst_cell_79_26 (.BL(BL26),.BLN(BLN26),.WL(WL79));
sram_cell_6t_5 inst_cell_79_27 (.BL(BL27),.BLN(BLN27),.WL(WL79));
sram_cell_6t_5 inst_cell_79_28 (.BL(BL28),.BLN(BLN28),.WL(WL79));
sram_cell_6t_5 inst_cell_79_29 (.BL(BL29),.BLN(BLN29),.WL(WL79));
sram_cell_6t_5 inst_cell_79_30 (.BL(BL30),.BLN(BLN30),.WL(WL79));
sram_cell_6t_5 inst_cell_79_31 (.BL(BL31),.BLN(BLN31),.WL(WL79));
sram_cell_6t_5 inst_cell_79_32 (.BL(BL32),.BLN(BLN32),.WL(WL79));
sram_cell_6t_5 inst_cell_79_33 (.BL(BL33),.BLN(BLN33),.WL(WL79));
sram_cell_6t_5 inst_cell_79_34 (.BL(BL34),.BLN(BLN34),.WL(WL79));
sram_cell_6t_5 inst_cell_79_35 (.BL(BL35),.BLN(BLN35),.WL(WL79));
sram_cell_6t_5 inst_cell_79_36 (.BL(BL36),.BLN(BLN36),.WL(WL79));
sram_cell_6t_5 inst_cell_79_37 (.BL(BL37),.BLN(BLN37),.WL(WL79));
sram_cell_6t_5 inst_cell_79_38 (.BL(BL38),.BLN(BLN38),.WL(WL79));
sram_cell_6t_5 inst_cell_79_39 (.BL(BL39),.BLN(BLN39),.WL(WL79));
sram_cell_6t_5 inst_cell_79_40 (.BL(BL40),.BLN(BLN40),.WL(WL79));
sram_cell_6t_5 inst_cell_79_41 (.BL(BL41),.BLN(BLN41),.WL(WL79));
sram_cell_6t_5 inst_cell_79_42 (.BL(BL42),.BLN(BLN42),.WL(WL79));
sram_cell_6t_5 inst_cell_79_43 (.BL(BL43),.BLN(BLN43),.WL(WL79));
sram_cell_6t_5 inst_cell_79_44 (.BL(BL44),.BLN(BLN44),.WL(WL79));
sram_cell_6t_5 inst_cell_79_45 (.BL(BL45),.BLN(BLN45),.WL(WL79));
sram_cell_6t_5 inst_cell_79_46 (.BL(BL46),.BLN(BLN46),.WL(WL79));
sram_cell_6t_5 inst_cell_79_47 (.BL(BL47),.BLN(BLN47),.WL(WL79));
sram_cell_6t_5 inst_cell_79_48 (.BL(BL48),.BLN(BLN48),.WL(WL79));
sram_cell_6t_5 inst_cell_79_49 (.BL(BL49),.BLN(BLN49),.WL(WL79));
sram_cell_6t_5 inst_cell_79_50 (.BL(BL50),.BLN(BLN50),.WL(WL79));
sram_cell_6t_5 inst_cell_79_51 (.BL(BL51),.BLN(BLN51),.WL(WL79));
sram_cell_6t_5 inst_cell_79_52 (.BL(BL52),.BLN(BLN52),.WL(WL79));
sram_cell_6t_5 inst_cell_79_53 (.BL(BL53),.BLN(BLN53),.WL(WL79));
sram_cell_6t_5 inst_cell_79_54 (.BL(BL54),.BLN(BLN54),.WL(WL79));
sram_cell_6t_5 inst_cell_79_55 (.BL(BL55),.BLN(BLN55),.WL(WL79));
sram_cell_6t_5 inst_cell_79_56 (.BL(BL56),.BLN(BLN56),.WL(WL79));
sram_cell_6t_5 inst_cell_79_57 (.BL(BL57),.BLN(BLN57),.WL(WL79));
sram_cell_6t_5 inst_cell_79_58 (.BL(BL58),.BLN(BLN58),.WL(WL79));
sram_cell_6t_5 inst_cell_79_59 (.BL(BL59),.BLN(BLN59),.WL(WL79));
sram_cell_6t_5 inst_cell_79_60 (.BL(BL60),.BLN(BLN60),.WL(WL79));
sram_cell_6t_5 inst_cell_79_61 (.BL(BL61),.BLN(BLN61),.WL(WL79));
sram_cell_6t_5 inst_cell_79_62 (.BL(BL62),.BLN(BLN62),.WL(WL79));
sram_cell_6t_5 inst_cell_79_63 (.BL(BL63),.BLN(BLN63),.WL(WL79));
sram_cell_6t_5 inst_cell_79_64 (.BL(BL64),.BLN(BLN64),.WL(WL79));
sram_cell_6t_5 inst_cell_79_65 (.BL(BL65),.BLN(BLN65),.WL(WL79));
sram_cell_6t_5 inst_cell_79_66 (.BL(BL66),.BLN(BLN66),.WL(WL79));
sram_cell_6t_5 inst_cell_79_67 (.BL(BL67),.BLN(BLN67),.WL(WL79));
sram_cell_6t_5 inst_cell_79_68 (.BL(BL68),.BLN(BLN68),.WL(WL79));
sram_cell_6t_5 inst_cell_79_69 (.BL(BL69),.BLN(BLN69),.WL(WL79));
sram_cell_6t_5 inst_cell_79_70 (.BL(BL70),.BLN(BLN70),.WL(WL79));
sram_cell_6t_5 inst_cell_79_71 (.BL(BL71),.BLN(BLN71),.WL(WL79));
sram_cell_6t_5 inst_cell_79_72 (.BL(BL72),.BLN(BLN72),.WL(WL79));
sram_cell_6t_5 inst_cell_79_73 (.BL(BL73),.BLN(BLN73),.WL(WL79));
sram_cell_6t_5 inst_cell_79_74 (.BL(BL74),.BLN(BLN74),.WL(WL79));
sram_cell_6t_5 inst_cell_79_75 (.BL(BL75),.BLN(BLN75),.WL(WL79));
sram_cell_6t_5 inst_cell_79_76 (.BL(BL76),.BLN(BLN76),.WL(WL79));
sram_cell_6t_5 inst_cell_79_77 (.BL(BL77),.BLN(BLN77),.WL(WL79));
sram_cell_6t_5 inst_cell_79_78 (.BL(BL78),.BLN(BLN78),.WL(WL79));
sram_cell_6t_5 inst_cell_79_79 (.BL(BL79),.BLN(BLN79),.WL(WL79));
sram_cell_6t_5 inst_cell_79_80 (.BL(BL80),.BLN(BLN80),.WL(WL79));
sram_cell_6t_5 inst_cell_79_81 (.BL(BL81),.BLN(BLN81),.WL(WL79));
sram_cell_6t_5 inst_cell_79_82 (.BL(BL82),.BLN(BLN82),.WL(WL79));
sram_cell_6t_5 inst_cell_79_83 (.BL(BL83),.BLN(BLN83),.WL(WL79));
sram_cell_6t_5 inst_cell_79_84 (.BL(BL84),.BLN(BLN84),.WL(WL79));
sram_cell_6t_5 inst_cell_79_85 (.BL(BL85),.BLN(BLN85),.WL(WL79));
sram_cell_6t_5 inst_cell_79_86 (.BL(BL86),.BLN(BLN86),.WL(WL79));
sram_cell_6t_5 inst_cell_79_87 (.BL(BL87),.BLN(BLN87),.WL(WL79));
sram_cell_6t_5 inst_cell_79_88 (.BL(BL88),.BLN(BLN88),.WL(WL79));
sram_cell_6t_5 inst_cell_79_89 (.BL(BL89),.BLN(BLN89),.WL(WL79));
sram_cell_6t_5 inst_cell_79_90 (.BL(BL90),.BLN(BLN90),.WL(WL79));
sram_cell_6t_5 inst_cell_79_91 (.BL(BL91),.BLN(BLN91),.WL(WL79));
sram_cell_6t_5 inst_cell_79_92 (.BL(BL92),.BLN(BLN92),.WL(WL79));
sram_cell_6t_5 inst_cell_79_93 (.BL(BL93),.BLN(BLN93),.WL(WL79));
sram_cell_6t_5 inst_cell_79_94 (.BL(BL94),.BLN(BLN94),.WL(WL79));
sram_cell_6t_5 inst_cell_79_95 (.BL(BL95),.BLN(BLN95),.WL(WL79));
sram_cell_6t_5 inst_cell_79_96 (.BL(BL96),.BLN(BLN96),.WL(WL79));
sram_cell_6t_5 inst_cell_79_97 (.BL(BL97),.BLN(BLN97),.WL(WL79));
sram_cell_6t_5 inst_cell_79_98 (.BL(BL98),.BLN(BLN98),.WL(WL79));
sram_cell_6t_5 inst_cell_79_99 (.BL(BL99),.BLN(BLN99),.WL(WL79));
sram_cell_6t_5 inst_cell_79_100 (.BL(BL100),.BLN(BLN100),.WL(WL79));
sram_cell_6t_5 inst_cell_79_101 (.BL(BL101),.BLN(BLN101),.WL(WL79));
sram_cell_6t_5 inst_cell_79_102 (.BL(BL102),.BLN(BLN102),.WL(WL79));
sram_cell_6t_5 inst_cell_79_103 (.BL(BL103),.BLN(BLN103),.WL(WL79));
sram_cell_6t_5 inst_cell_79_104 (.BL(BL104),.BLN(BLN104),.WL(WL79));
sram_cell_6t_5 inst_cell_79_105 (.BL(BL105),.BLN(BLN105),.WL(WL79));
sram_cell_6t_5 inst_cell_79_106 (.BL(BL106),.BLN(BLN106),.WL(WL79));
sram_cell_6t_5 inst_cell_79_107 (.BL(BL107),.BLN(BLN107),.WL(WL79));
sram_cell_6t_5 inst_cell_79_108 (.BL(BL108),.BLN(BLN108),.WL(WL79));
sram_cell_6t_5 inst_cell_79_109 (.BL(BL109),.BLN(BLN109),.WL(WL79));
sram_cell_6t_5 inst_cell_79_110 (.BL(BL110),.BLN(BLN110),.WL(WL79));
sram_cell_6t_5 inst_cell_79_111 (.BL(BL111),.BLN(BLN111),.WL(WL79));
sram_cell_6t_5 inst_cell_79_112 (.BL(BL112),.BLN(BLN112),.WL(WL79));
sram_cell_6t_5 inst_cell_79_113 (.BL(BL113),.BLN(BLN113),.WL(WL79));
sram_cell_6t_5 inst_cell_79_114 (.BL(BL114),.BLN(BLN114),.WL(WL79));
sram_cell_6t_5 inst_cell_79_115 (.BL(BL115),.BLN(BLN115),.WL(WL79));
sram_cell_6t_5 inst_cell_79_116 (.BL(BL116),.BLN(BLN116),.WL(WL79));
sram_cell_6t_5 inst_cell_79_117 (.BL(BL117),.BLN(BLN117),.WL(WL79));
sram_cell_6t_5 inst_cell_79_118 (.BL(BL118),.BLN(BLN118),.WL(WL79));
sram_cell_6t_5 inst_cell_79_119 (.BL(BL119),.BLN(BLN119),.WL(WL79));
sram_cell_6t_5 inst_cell_79_120 (.BL(BL120),.BLN(BLN120),.WL(WL79));
sram_cell_6t_5 inst_cell_79_121 (.BL(BL121),.BLN(BLN121),.WL(WL79));
sram_cell_6t_5 inst_cell_79_122 (.BL(BL122),.BLN(BLN122),.WL(WL79));
sram_cell_6t_5 inst_cell_79_123 (.BL(BL123),.BLN(BLN123),.WL(WL79));
sram_cell_6t_5 inst_cell_79_124 (.BL(BL124),.BLN(BLN124),.WL(WL79));
sram_cell_6t_5 inst_cell_79_125 (.BL(BL125),.BLN(BLN125),.WL(WL79));
sram_cell_6t_5 inst_cell_79_126 (.BL(BL126),.BLN(BLN126),.WL(WL79));
sram_cell_6t_5 inst_cell_79_127 (.BL(BL127),.BLN(BLN127),.WL(WL79));
sram_cell_6t_5 inst_cell_80_0 (.BL(BL0),.BLN(BLN0),.WL(WL80));
sram_cell_6t_5 inst_cell_80_1 (.BL(BL1),.BLN(BLN1),.WL(WL80));
sram_cell_6t_5 inst_cell_80_2 (.BL(BL2),.BLN(BLN2),.WL(WL80));
sram_cell_6t_5 inst_cell_80_3 (.BL(BL3),.BLN(BLN3),.WL(WL80));
sram_cell_6t_5 inst_cell_80_4 (.BL(BL4),.BLN(BLN4),.WL(WL80));
sram_cell_6t_5 inst_cell_80_5 (.BL(BL5),.BLN(BLN5),.WL(WL80));
sram_cell_6t_5 inst_cell_80_6 (.BL(BL6),.BLN(BLN6),.WL(WL80));
sram_cell_6t_5 inst_cell_80_7 (.BL(BL7),.BLN(BLN7),.WL(WL80));
sram_cell_6t_5 inst_cell_80_8 (.BL(BL8),.BLN(BLN8),.WL(WL80));
sram_cell_6t_5 inst_cell_80_9 (.BL(BL9),.BLN(BLN9),.WL(WL80));
sram_cell_6t_5 inst_cell_80_10 (.BL(BL10),.BLN(BLN10),.WL(WL80));
sram_cell_6t_5 inst_cell_80_11 (.BL(BL11),.BLN(BLN11),.WL(WL80));
sram_cell_6t_5 inst_cell_80_12 (.BL(BL12),.BLN(BLN12),.WL(WL80));
sram_cell_6t_5 inst_cell_80_13 (.BL(BL13),.BLN(BLN13),.WL(WL80));
sram_cell_6t_5 inst_cell_80_14 (.BL(BL14),.BLN(BLN14),.WL(WL80));
sram_cell_6t_5 inst_cell_80_15 (.BL(BL15),.BLN(BLN15),.WL(WL80));
sram_cell_6t_5 inst_cell_80_16 (.BL(BL16),.BLN(BLN16),.WL(WL80));
sram_cell_6t_5 inst_cell_80_17 (.BL(BL17),.BLN(BLN17),.WL(WL80));
sram_cell_6t_5 inst_cell_80_18 (.BL(BL18),.BLN(BLN18),.WL(WL80));
sram_cell_6t_5 inst_cell_80_19 (.BL(BL19),.BLN(BLN19),.WL(WL80));
sram_cell_6t_5 inst_cell_80_20 (.BL(BL20),.BLN(BLN20),.WL(WL80));
sram_cell_6t_5 inst_cell_80_21 (.BL(BL21),.BLN(BLN21),.WL(WL80));
sram_cell_6t_5 inst_cell_80_22 (.BL(BL22),.BLN(BLN22),.WL(WL80));
sram_cell_6t_5 inst_cell_80_23 (.BL(BL23),.BLN(BLN23),.WL(WL80));
sram_cell_6t_5 inst_cell_80_24 (.BL(BL24),.BLN(BLN24),.WL(WL80));
sram_cell_6t_5 inst_cell_80_25 (.BL(BL25),.BLN(BLN25),.WL(WL80));
sram_cell_6t_5 inst_cell_80_26 (.BL(BL26),.BLN(BLN26),.WL(WL80));
sram_cell_6t_5 inst_cell_80_27 (.BL(BL27),.BLN(BLN27),.WL(WL80));
sram_cell_6t_5 inst_cell_80_28 (.BL(BL28),.BLN(BLN28),.WL(WL80));
sram_cell_6t_5 inst_cell_80_29 (.BL(BL29),.BLN(BLN29),.WL(WL80));
sram_cell_6t_5 inst_cell_80_30 (.BL(BL30),.BLN(BLN30),.WL(WL80));
sram_cell_6t_5 inst_cell_80_31 (.BL(BL31),.BLN(BLN31),.WL(WL80));
sram_cell_6t_5 inst_cell_80_32 (.BL(BL32),.BLN(BLN32),.WL(WL80));
sram_cell_6t_5 inst_cell_80_33 (.BL(BL33),.BLN(BLN33),.WL(WL80));
sram_cell_6t_5 inst_cell_80_34 (.BL(BL34),.BLN(BLN34),.WL(WL80));
sram_cell_6t_5 inst_cell_80_35 (.BL(BL35),.BLN(BLN35),.WL(WL80));
sram_cell_6t_5 inst_cell_80_36 (.BL(BL36),.BLN(BLN36),.WL(WL80));
sram_cell_6t_5 inst_cell_80_37 (.BL(BL37),.BLN(BLN37),.WL(WL80));
sram_cell_6t_5 inst_cell_80_38 (.BL(BL38),.BLN(BLN38),.WL(WL80));
sram_cell_6t_5 inst_cell_80_39 (.BL(BL39),.BLN(BLN39),.WL(WL80));
sram_cell_6t_5 inst_cell_80_40 (.BL(BL40),.BLN(BLN40),.WL(WL80));
sram_cell_6t_5 inst_cell_80_41 (.BL(BL41),.BLN(BLN41),.WL(WL80));
sram_cell_6t_5 inst_cell_80_42 (.BL(BL42),.BLN(BLN42),.WL(WL80));
sram_cell_6t_5 inst_cell_80_43 (.BL(BL43),.BLN(BLN43),.WL(WL80));
sram_cell_6t_5 inst_cell_80_44 (.BL(BL44),.BLN(BLN44),.WL(WL80));
sram_cell_6t_5 inst_cell_80_45 (.BL(BL45),.BLN(BLN45),.WL(WL80));
sram_cell_6t_5 inst_cell_80_46 (.BL(BL46),.BLN(BLN46),.WL(WL80));
sram_cell_6t_5 inst_cell_80_47 (.BL(BL47),.BLN(BLN47),.WL(WL80));
sram_cell_6t_5 inst_cell_80_48 (.BL(BL48),.BLN(BLN48),.WL(WL80));
sram_cell_6t_5 inst_cell_80_49 (.BL(BL49),.BLN(BLN49),.WL(WL80));
sram_cell_6t_5 inst_cell_80_50 (.BL(BL50),.BLN(BLN50),.WL(WL80));
sram_cell_6t_5 inst_cell_80_51 (.BL(BL51),.BLN(BLN51),.WL(WL80));
sram_cell_6t_5 inst_cell_80_52 (.BL(BL52),.BLN(BLN52),.WL(WL80));
sram_cell_6t_5 inst_cell_80_53 (.BL(BL53),.BLN(BLN53),.WL(WL80));
sram_cell_6t_5 inst_cell_80_54 (.BL(BL54),.BLN(BLN54),.WL(WL80));
sram_cell_6t_5 inst_cell_80_55 (.BL(BL55),.BLN(BLN55),.WL(WL80));
sram_cell_6t_5 inst_cell_80_56 (.BL(BL56),.BLN(BLN56),.WL(WL80));
sram_cell_6t_5 inst_cell_80_57 (.BL(BL57),.BLN(BLN57),.WL(WL80));
sram_cell_6t_5 inst_cell_80_58 (.BL(BL58),.BLN(BLN58),.WL(WL80));
sram_cell_6t_5 inst_cell_80_59 (.BL(BL59),.BLN(BLN59),.WL(WL80));
sram_cell_6t_5 inst_cell_80_60 (.BL(BL60),.BLN(BLN60),.WL(WL80));
sram_cell_6t_5 inst_cell_80_61 (.BL(BL61),.BLN(BLN61),.WL(WL80));
sram_cell_6t_5 inst_cell_80_62 (.BL(BL62),.BLN(BLN62),.WL(WL80));
sram_cell_6t_5 inst_cell_80_63 (.BL(BL63),.BLN(BLN63),.WL(WL80));
sram_cell_6t_5 inst_cell_80_64 (.BL(BL64),.BLN(BLN64),.WL(WL80));
sram_cell_6t_5 inst_cell_80_65 (.BL(BL65),.BLN(BLN65),.WL(WL80));
sram_cell_6t_5 inst_cell_80_66 (.BL(BL66),.BLN(BLN66),.WL(WL80));
sram_cell_6t_5 inst_cell_80_67 (.BL(BL67),.BLN(BLN67),.WL(WL80));
sram_cell_6t_5 inst_cell_80_68 (.BL(BL68),.BLN(BLN68),.WL(WL80));
sram_cell_6t_5 inst_cell_80_69 (.BL(BL69),.BLN(BLN69),.WL(WL80));
sram_cell_6t_5 inst_cell_80_70 (.BL(BL70),.BLN(BLN70),.WL(WL80));
sram_cell_6t_5 inst_cell_80_71 (.BL(BL71),.BLN(BLN71),.WL(WL80));
sram_cell_6t_5 inst_cell_80_72 (.BL(BL72),.BLN(BLN72),.WL(WL80));
sram_cell_6t_5 inst_cell_80_73 (.BL(BL73),.BLN(BLN73),.WL(WL80));
sram_cell_6t_5 inst_cell_80_74 (.BL(BL74),.BLN(BLN74),.WL(WL80));
sram_cell_6t_5 inst_cell_80_75 (.BL(BL75),.BLN(BLN75),.WL(WL80));
sram_cell_6t_5 inst_cell_80_76 (.BL(BL76),.BLN(BLN76),.WL(WL80));
sram_cell_6t_5 inst_cell_80_77 (.BL(BL77),.BLN(BLN77),.WL(WL80));
sram_cell_6t_5 inst_cell_80_78 (.BL(BL78),.BLN(BLN78),.WL(WL80));
sram_cell_6t_5 inst_cell_80_79 (.BL(BL79),.BLN(BLN79),.WL(WL80));
sram_cell_6t_5 inst_cell_80_80 (.BL(BL80),.BLN(BLN80),.WL(WL80));
sram_cell_6t_5 inst_cell_80_81 (.BL(BL81),.BLN(BLN81),.WL(WL80));
sram_cell_6t_5 inst_cell_80_82 (.BL(BL82),.BLN(BLN82),.WL(WL80));
sram_cell_6t_5 inst_cell_80_83 (.BL(BL83),.BLN(BLN83),.WL(WL80));
sram_cell_6t_5 inst_cell_80_84 (.BL(BL84),.BLN(BLN84),.WL(WL80));
sram_cell_6t_5 inst_cell_80_85 (.BL(BL85),.BLN(BLN85),.WL(WL80));
sram_cell_6t_5 inst_cell_80_86 (.BL(BL86),.BLN(BLN86),.WL(WL80));
sram_cell_6t_5 inst_cell_80_87 (.BL(BL87),.BLN(BLN87),.WL(WL80));
sram_cell_6t_5 inst_cell_80_88 (.BL(BL88),.BLN(BLN88),.WL(WL80));
sram_cell_6t_5 inst_cell_80_89 (.BL(BL89),.BLN(BLN89),.WL(WL80));
sram_cell_6t_5 inst_cell_80_90 (.BL(BL90),.BLN(BLN90),.WL(WL80));
sram_cell_6t_5 inst_cell_80_91 (.BL(BL91),.BLN(BLN91),.WL(WL80));
sram_cell_6t_5 inst_cell_80_92 (.BL(BL92),.BLN(BLN92),.WL(WL80));
sram_cell_6t_5 inst_cell_80_93 (.BL(BL93),.BLN(BLN93),.WL(WL80));
sram_cell_6t_5 inst_cell_80_94 (.BL(BL94),.BLN(BLN94),.WL(WL80));
sram_cell_6t_5 inst_cell_80_95 (.BL(BL95),.BLN(BLN95),.WL(WL80));
sram_cell_6t_5 inst_cell_80_96 (.BL(BL96),.BLN(BLN96),.WL(WL80));
sram_cell_6t_5 inst_cell_80_97 (.BL(BL97),.BLN(BLN97),.WL(WL80));
sram_cell_6t_5 inst_cell_80_98 (.BL(BL98),.BLN(BLN98),.WL(WL80));
sram_cell_6t_5 inst_cell_80_99 (.BL(BL99),.BLN(BLN99),.WL(WL80));
sram_cell_6t_5 inst_cell_80_100 (.BL(BL100),.BLN(BLN100),.WL(WL80));
sram_cell_6t_5 inst_cell_80_101 (.BL(BL101),.BLN(BLN101),.WL(WL80));
sram_cell_6t_5 inst_cell_80_102 (.BL(BL102),.BLN(BLN102),.WL(WL80));
sram_cell_6t_5 inst_cell_80_103 (.BL(BL103),.BLN(BLN103),.WL(WL80));
sram_cell_6t_5 inst_cell_80_104 (.BL(BL104),.BLN(BLN104),.WL(WL80));
sram_cell_6t_5 inst_cell_80_105 (.BL(BL105),.BLN(BLN105),.WL(WL80));
sram_cell_6t_5 inst_cell_80_106 (.BL(BL106),.BLN(BLN106),.WL(WL80));
sram_cell_6t_5 inst_cell_80_107 (.BL(BL107),.BLN(BLN107),.WL(WL80));
sram_cell_6t_5 inst_cell_80_108 (.BL(BL108),.BLN(BLN108),.WL(WL80));
sram_cell_6t_5 inst_cell_80_109 (.BL(BL109),.BLN(BLN109),.WL(WL80));
sram_cell_6t_5 inst_cell_80_110 (.BL(BL110),.BLN(BLN110),.WL(WL80));
sram_cell_6t_5 inst_cell_80_111 (.BL(BL111),.BLN(BLN111),.WL(WL80));
sram_cell_6t_5 inst_cell_80_112 (.BL(BL112),.BLN(BLN112),.WL(WL80));
sram_cell_6t_5 inst_cell_80_113 (.BL(BL113),.BLN(BLN113),.WL(WL80));
sram_cell_6t_5 inst_cell_80_114 (.BL(BL114),.BLN(BLN114),.WL(WL80));
sram_cell_6t_5 inst_cell_80_115 (.BL(BL115),.BLN(BLN115),.WL(WL80));
sram_cell_6t_5 inst_cell_80_116 (.BL(BL116),.BLN(BLN116),.WL(WL80));
sram_cell_6t_5 inst_cell_80_117 (.BL(BL117),.BLN(BLN117),.WL(WL80));
sram_cell_6t_5 inst_cell_80_118 (.BL(BL118),.BLN(BLN118),.WL(WL80));
sram_cell_6t_5 inst_cell_80_119 (.BL(BL119),.BLN(BLN119),.WL(WL80));
sram_cell_6t_5 inst_cell_80_120 (.BL(BL120),.BLN(BLN120),.WL(WL80));
sram_cell_6t_5 inst_cell_80_121 (.BL(BL121),.BLN(BLN121),.WL(WL80));
sram_cell_6t_5 inst_cell_80_122 (.BL(BL122),.BLN(BLN122),.WL(WL80));
sram_cell_6t_5 inst_cell_80_123 (.BL(BL123),.BLN(BLN123),.WL(WL80));
sram_cell_6t_5 inst_cell_80_124 (.BL(BL124),.BLN(BLN124),.WL(WL80));
sram_cell_6t_5 inst_cell_80_125 (.BL(BL125),.BLN(BLN125),.WL(WL80));
sram_cell_6t_5 inst_cell_80_126 (.BL(BL126),.BLN(BLN126),.WL(WL80));
sram_cell_6t_5 inst_cell_80_127 (.BL(BL127),.BLN(BLN127),.WL(WL80));
sram_cell_6t_5 inst_cell_81_0 (.BL(BL0),.BLN(BLN0),.WL(WL81));
sram_cell_6t_5 inst_cell_81_1 (.BL(BL1),.BLN(BLN1),.WL(WL81));
sram_cell_6t_5 inst_cell_81_2 (.BL(BL2),.BLN(BLN2),.WL(WL81));
sram_cell_6t_5 inst_cell_81_3 (.BL(BL3),.BLN(BLN3),.WL(WL81));
sram_cell_6t_5 inst_cell_81_4 (.BL(BL4),.BLN(BLN4),.WL(WL81));
sram_cell_6t_5 inst_cell_81_5 (.BL(BL5),.BLN(BLN5),.WL(WL81));
sram_cell_6t_5 inst_cell_81_6 (.BL(BL6),.BLN(BLN6),.WL(WL81));
sram_cell_6t_5 inst_cell_81_7 (.BL(BL7),.BLN(BLN7),.WL(WL81));
sram_cell_6t_5 inst_cell_81_8 (.BL(BL8),.BLN(BLN8),.WL(WL81));
sram_cell_6t_5 inst_cell_81_9 (.BL(BL9),.BLN(BLN9),.WL(WL81));
sram_cell_6t_5 inst_cell_81_10 (.BL(BL10),.BLN(BLN10),.WL(WL81));
sram_cell_6t_5 inst_cell_81_11 (.BL(BL11),.BLN(BLN11),.WL(WL81));
sram_cell_6t_5 inst_cell_81_12 (.BL(BL12),.BLN(BLN12),.WL(WL81));
sram_cell_6t_5 inst_cell_81_13 (.BL(BL13),.BLN(BLN13),.WL(WL81));
sram_cell_6t_5 inst_cell_81_14 (.BL(BL14),.BLN(BLN14),.WL(WL81));
sram_cell_6t_5 inst_cell_81_15 (.BL(BL15),.BLN(BLN15),.WL(WL81));
sram_cell_6t_5 inst_cell_81_16 (.BL(BL16),.BLN(BLN16),.WL(WL81));
sram_cell_6t_5 inst_cell_81_17 (.BL(BL17),.BLN(BLN17),.WL(WL81));
sram_cell_6t_5 inst_cell_81_18 (.BL(BL18),.BLN(BLN18),.WL(WL81));
sram_cell_6t_5 inst_cell_81_19 (.BL(BL19),.BLN(BLN19),.WL(WL81));
sram_cell_6t_5 inst_cell_81_20 (.BL(BL20),.BLN(BLN20),.WL(WL81));
sram_cell_6t_5 inst_cell_81_21 (.BL(BL21),.BLN(BLN21),.WL(WL81));
sram_cell_6t_5 inst_cell_81_22 (.BL(BL22),.BLN(BLN22),.WL(WL81));
sram_cell_6t_5 inst_cell_81_23 (.BL(BL23),.BLN(BLN23),.WL(WL81));
sram_cell_6t_5 inst_cell_81_24 (.BL(BL24),.BLN(BLN24),.WL(WL81));
sram_cell_6t_5 inst_cell_81_25 (.BL(BL25),.BLN(BLN25),.WL(WL81));
sram_cell_6t_5 inst_cell_81_26 (.BL(BL26),.BLN(BLN26),.WL(WL81));
sram_cell_6t_5 inst_cell_81_27 (.BL(BL27),.BLN(BLN27),.WL(WL81));
sram_cell_6t_5 inst_cell_81_28 (.BL(BL28),.BLN(BLN28),.WL(WL81));
sram_cell_6t_5 inst_cell_81_29 (.BL(BL29),.BLN(BLN29),.WL(WL81));
sram_cell_6t_5 inst_cell_81_30 (.BL(BL30),.BLN(BLN30),.WL(WL81));
sram_cell_6t_5 inst_cell_81_31 (.BL(BL31),.BLN(BLN31),.WL(WL81));
sram_cell_6t_5 inst_cell_81_32 (.BL(BL32),.BLN(BLN32),.WL(WL81));
sram_cell_6t_5 inst_cell_81_33 (.BL(BL33),.BLN(BLN33),.WL(WL81));
sram_cell_6t_5 inst_cell_81_34 (.BL(BL34),.BLN(BLN34),.WL(WL81));
sram_cell_6t_5 inst_cell_81_35 (.BL(BL35),.BLN(BLN35),.WL(WL81));
sram_cell_6t_5 inst_cell_81_36 (.BL(BL36),.BLN(BLN36),.WL(WL81));
sram_cell_6t_5 inst_cell_81_37 (.BL(BL37),.BLN(BLN37),.WL(WL81));
sram_cell_6t_5 inst_cell_81_38 (.BL(BL38),.BLN(BLN38),.WL(WL81));
sram_cell_6t_5 inst_cell_81_39 (.BL(BL39),.BLN(BLN39),.WL(WL81));
sram_cell_6t_5 inst_cell_81_40 (.BL(BL40),.BLN(BLN40),.WL(WL81));
sram_cell_6t_5 inst_cell_81_41 (.BL(BL41),.BLN(BLN41),.WL(WL81));
sram_cell_6t_5 inst_cell_81_42 (.BL(BL42),.BLN(BLN42),.WL(WL81));
sram_cell_6t_5 inst_cell_81_43 (.BL(BL43),.BLN(BLN43),.WL(WL81));
sram_cell_6t_5 inst_cell_81_44 (.BL(BL44),.BLN(BLN44),.WL(WL81));
sram_cell_6t_5 inst_cell_81_45 (.BL(BL45),.BLN(BLN45),.WL(WL81));
sram_cell_6t_5 inst_cell_81_46 (.BL(BL46),.BLN(BLN46),.WL(WL81));
sram_cell_6t_5 inst_cell_81_47 (.BL(BL47),.BLN(BLN47),.WL(WL81));
sram_cell_6t_5 inst_cell_81_48 (.BL(BL48),.BLN(BLN48),.WL(WL81));
sram_cell_6t_5 inst_cell_81_49 (.BL(BL49),.BLN(BLN49),.WL(WL81));
sram_cell_6t_5 inst_cell_81_50 (.BL(BL50),.BLN(BLN50),.WL(WL81));
sram_cell_6t_5 inst_cell_81_51 (.BL(BL51),.BLN(BLN51),.WL(WL81));
sram_cell_6t_5 inst_cell_81_52 (.BL(BL52),.BLN(BLN52),.WL(WL81));
sram_cell_6t_5 inst_cell_81_53 (.BL(BL53),.BLN(BLN53),.WL(WL81));
sram_cell_6t_5 inst_cell_81_54 (.BL(BL54),.BLN(BLN54),.WL(WL81));
sram_cell_6t_5 inst_cell_81_55 (.BL(BL55),.BLN(BLN55),.WL(WL81));
sram_cell_6t_5 inst_cell_81_56 (.BL(BL56),.BLN(BLN56),.WL(WL81));
sram_cell_6t_5 inst_cell_81_57 (.BL(BL57),.BLN(BLN57),.WL(WL81));
sram_cell_6t_5 inst_cell_81_58 (.BL(BL58),.BLN(BLN58),.WL(WL81));
sram_cell_6t_5 inst_cell_81_59 (.BL(BL59),.BLN(BLN59),.WL(WL81));
sram_cell_6t_5 inst_cell_81_60 (.BL(BL60),.BLN(BLN60),.WL(WL81));
sram_cell_6t_5 inst_cell_81_61 (.BL(BL61),.BLN(BLN61),.WL(WL81));
sram_cell_6t_5 inst_cell_81_62 (.BL(BL62),.BLN(BLN62),.WL(WL81));
sram_cell_6t_5 inst_cell_81_63 (.BL(BL63),.BLN(BLN63),.WL(WL81));
sram_cell_6t_5 inst_cell_81_64 (.BL(BL64),.BLN(BLN64),.WL(WL81));
sram_cell_6t_5 inst_cell_81_65 (.BL(BL65),.BLN(BLN65),.WL(WL81));
sram_cell_6t_5 inst_cell_81_66 (.BL(BL66),.BLN(BLN66),.WL(WL81));
sram_cell_6t_5 inst_cell_81_67 (.BL(BL67),.BLN(BLN67),.WL(WL81));
sram_cell_6t_5 inst_cell_81_68 (.BL(BL68),.BLN(BLN68),.WL(WL81));
sram_cell_6t_5 inst_cell_81_69 (.BL(BL69),.BLN(BLN69),.WL(WL81));
sram_cell_6t_5 inst_cell_81_70 (.BL(BL70),.BLN(BLN70),.WL(WL81));
sram_cell_6t_5 inst_cell_81_71 (.BL(BL71),.BLN(BLN71),.WL(WL81));
sram_cell_6t_5 inst_cell_81_72 (.BL(BL72),.BLN(BLN72),.WL(WL81));
sram_cell_6t_5 inst_cell_81_73 (.BL(BL73),.BLN(BLN73),.WL(WL81));
sram_cell_6t_5 inst_cell_81_74 (.BL(BL74),.BLN(BLN74),.WL(WL81));
sram_cell_6t_5 inst_cell_81_75 (.BL(BL75),.BLN(BLN75),.WL(WL81));
sram_cell_6t_5 inst_cell_81_76 (.BL(BL76),.BLN(BLN76),.WL(WL81));
sram_cell_6t_5 inst_cell_81_77 (.BL(BL77),.BLN(BLN77),.WL(WL81));
sram_cell_6t_5 inst_cell_81_78 (.BL(BL78),.BLN(BLN78),.WL(WL81));
sram_cell_6t_5 inst_cell_81_79 (.BL(BL79),.BLN(BLN79),.WL(WL81));
sram_cell_6t_5 inst_cell_81_80 (.BL(BL80),.BLN(BLN80),.WL(WL81));
sram_cell_6t_5 inst_cell_81_81 (.BL(BL81),.BLN(BLN81),.WL(WL81));
sram_cell_6t_5 inst_cell_81_82 (.BL(BL82),.BLN(BLN82),.WL(WL81));
sram_cell_6t_5 inst_cell_81_83 (.BL(BL83),.BLN(BLN83),.WL(WL81));
sram_cell_6t_5 inst_cell_81_84 (.BL(BL84),.BLN(BLN84),.WL(WL81));
sram_cell_6t_5 inst_cell_81_85 (.BL(BL85),.BLN(BLN85),.WL(WL81));
sram_cell_6t_5 inst_cell_81_86 (.BL(BL86),.BLN(BLN86),.WL(WL81));
sram_cell_6t_5 inst_cell_81_87 (.BL(BL87),.BLN(BLN87),.WL(WL81));
sram_cell_6t_5 inst_cell_81_88 (.BL(BL88),.BLN(BLN88),.WL(WL81));
sram_cell_6t_5 inst_cell_81_89 (.BL(BL89),.BLN(BLN89),.WL(WL81));
sram_cell_6t_5 inst_cell_81_90 (.BL(BL90),.BLN(BLN90),.WL(WL81));
sram_cell_6t_5 inst_cell_81_91 (.BL(BL91),.BLN(BLN91),.WL(WL81));
sram_cell_6t_5 inst_cell_81_92 (.BL(BL92),.BLN(BLN92),.WL(WL81));
sram_cell_6t_5 inst_cell_81_93 (.BL(BL93),.BLN(BLN93),.WL(WL81));
sram_cell_6t_5 inst_cell_81_94 (.BL(BL94),.BLN(BLN94),.WL(WL81));
sram_cell_6t_5 inst_cell_81_95 (.BL(BL95),.BLN(BLN95),.WL(WL81));
sram_cell_6t_5 inst_cell_81_96 (.BL(BL96),.BLN(BLN96),.WL(WL81));
sram_cell_6t_5 inst_cell_81_97 (.BL(BL97),.BLN(BLN97),.WL(WL81));
sram_cell_6t_5 inst_cell_81_98 (.BL(BL98),.BLN(BLN98),.WL(WL81));
sram_cell_6t_5 inst_cell_81_99 (.BL(BL99),.BLN(BLN99),.WL(WL81));
sram_cell_6t_5 inst_cell_81_100 (.BL(BL100),.BLN(BLN100),.WL(WL81));
sram_cell_6t_5 inst_cell_81_101 (.BL(BL101),.BLN(BLN101),.WL(WL81));
sram_cell_6t_5 inst_cell_81_102 (.BL(BL102),.BLN(BLN102),.WL(WL81));
sram_cell_6t_5 inst_cell_81_103 (.BL(BL103),.BLN(BLN103),.WL(WL81));
sram_cell_6t_5 inst_cell_81_104 (.BL(BL104),.BLN(BLN104),.WL(WL81));
sram_cell_6t_5 inst_cell_81_105 (.BL(BL105),.BLN(BLN105),.WL(WL81));
sram_cell_6t_5 inst_cell_81_106 (.BL(BL106),.BLN(BLN106),.WL(WL81));
sram_cell_6t_5 inst_cell_81_107 (.BL(BL107),.BLN(BLN107),.WL(WL81));
sram_cell_6t_5 inst_cell_81_108 (.BL(BL108),.BLN(BLN108),.WL(WL81));
sram_cell_6t_5 inst_cell_81_109 (.BL(BL109),.BLN(BLN109),.WL(WL81));
sram_cell_6t_5 inst_cell_81_110 (.BL(BL110),.BLN(BLN110),.WL(WL81));
sram_cell_6t_5 inst_cell_81_111 (.BL(BL111),.BLN(BLN111),.WL(WL81));
sram_cell_6t_5 inst_cell_81_112 (.BL(BL112),.BLN(BLN112),.WL(WL81));
sram_cell_6t_5 inst_cell_81_113 (.BL(BL113),.BLN(BLN113),.WL(WL81));
sram_cell_6t_5 inst_cell_81_114 (.BL(BL114),.BLN(BLN114),.WL(WL81));
sram_cell_6t_5 inst_cell_81_115 (.BL(BL115),.BLN(BLN115),.WL(WL81));
sram_cell_6t_5 inst_cell_81_116 (.BL(BL116),.BLN(BLN116),.WL(WL81));
sram_cell_6t_5 inst_cell_81_117 (.BL(BL117),.BLN(BLN117),.WL(WL81));
sram_cell_6t_5 inst_cell_81_118 (.BL(BL118),.BLN(BLN118),.WL(WL81));
sram_cell_6t_5 inst_cell_81_119 (.BL(BL119),.BLN(BLN119),.WL(WL81));
sram_cell_6t_5 inst_cell_81_120 (.BL(BL120),.BLN(BLN120),.WL(WL81));
sram_cell_6t_5 inst_cell_81_121 (.BL(BL121),.BLN(BLN121),.WL(WL81));
sram_cell_6t_5 inst_cell_81_122 (.BL(BL122),.BLN(BLN122),.WL(WL81));
sram_cell_6t_5 inst_cell_81_123 (.BL(BL123),.BLN(BLN123),.WL(WL81));
sram_cell_6t_5 inst_cell_81_124 (.BL(BL124),.BLN(BLN124),.WL(WL81));
sram_cell_6t_5 inst_cell_81_125 (.BL(BL125),.BLN(BLN125),.WL(WL81));
sram_cell_6t_5 inst_cell_81_126 (.BL(BL126),.BLN(BLN126),.WL(WL81));
sram_cell_6t_5 inst_cell_81_127 (.BL(BL127),.BLN(BLN127),.WL(WL81));
sram_cell_6t_5 inst_cell_82_0 (.BL(BL0),.BLN(BLN0),.WL(WL82));
sram_cell_6t_5 inst_cell_82_1 (.BL(BL1),.BLN(BLN1),.WL(WL82));
sram_cell_6t_5 inst_cell_82_2 (.BL(BL2),.BLN(BLN2),.WL(WL82));
sram_cell_6t_5 inst_cell_82_3 (.BL(BL3),.BLN(BLN3),.WL(WL82));
sram_cell_6t_5 inst_cell_82_4 (.BL(BL4),.BLN(BLN4),.WL(WL82));
sram_cell_6t_5 inst_cell_82_5 (.BL(BL5),.BLN(BLN5),.WL(WL82));
sram_cell_6t_5 inst_cell_82_6 (.BL(BL6),.BLN(BLN6),.WL(WL82));
sram_cell_6t_5 inst_cell_82_7 (.BL(BL7),.BLN(BLN7),.WL(WL82));
sram_cell_6t_5 inst_cell_82_8 (.BL(BL8),.BLN(BLN8),.WL(WL82));
sram_cell_6t_5 inst_cell_82_9 (.BL(BL9),.BLN(BLN9),.WL(WL82));
sram_cell_6t_5 inst_cell_82_10 (.BL(BL10),.BLN(BLN10),.WL(WL82));
sram_cell_6t_5 inst_cell_82_11 (.BL(BL11),.BLN(BLN11),.WL(WL82));
sram_cell_6t_5 inst_cell_82_12 (.BL(BL12),.BLN(BLN12),.WL(WL82));
sram_cell_6t_5 inst_cell_82_13 (.BL(BL13),.BLN(BLN13),.WL(WL82));
sram_cell_6t_5 inst_cell_82_14 (.BL(BL14),.BLN(BLN14),.WL(WL82));
sram_cell_6t_5 inst_cell_82_15 (.BL(BL15),.BLN(BLN15),.WL(WL82));
sram_cell_6t_5 inst_cell_82_16 (.BL(BL16),.BLN(BLN16),.WL(WL82));
sram_cell_6t_5 inst_cell_82_17 (.BL(BL17),.BLN(BLN17),.WL(WL82));
sram_cell_6t_5 inst_cell_82_18 (.BL(BL18),.BLN(BLN18),.WL(WL82));
sram_cell_6t_5 inst_cell_82_19 (.BL(BL19),.BLN(BLN19),.WL(WL82));
sram_cell_6t_5 inst_cell_82_20 (.BL(BL20),.BLN(BLN20),.WL(WL82));
sram_cell_6t_5 inst_cell_82_21 (.BL(BL21),.BLN(BLN21),.WL(WL82));
sram_cell_6t_5 inst_cell_82_22 (.BL(BL22),.BLN(BLN22),.WL(WL82));
sram_cell_6t_5 inst_cell_82_23 (.BL(BL23),.BLN(BLN23),.WL(WL82));
sram_cell_6t_5 inst_cell_82_24 (.BL(BL24),.BLN(BLN24),.WL(WL82));
sram_cell_6t_5 inst_cell_82_25 (.BL(BL25),.BLN(BLN25),.WL(WL82));
sram_cell_6t_5 inst_cell_82_26 (.BL(BL26),.BLN(BLN26),.WL(WL82));
sram_cell_6t_5 inst_cell_82_27 (.BL(BL27),.BLN(BLN27),.WL(WL82));
sram_cell_6t_5 inst_cell_82_28 (.BL(BL28),.BLN(BLN28),.WL(WL82));
sram_cell_6t_5 inst_cell_82_29 (.BL(BL29),.BLN(BLN29),.WL(WL82));
sram_cell_6t_5 inst_cell_82_30 (.BL(BL30),.BLN(BLN30),.WL(WL82));
sram_cell_6t_5 inst_cell_82_31 (.BL(BL31),.BLN(BLN31),.WL(WL82));
sram_cell_6t_5 inst_cell_82_32 (.BL(BL32),.BLN(BLN32),.WL(WL82));
sram_cell_6t_5 inst_cell_82_33 (.BL(BL33),.BLN(BLN33),.WL(WL82));
sram_cell_6t_5 inst_cell_82_34 (.BL(BL34),.BLN(BLN34),.WL(WL82));
sram_cell_6t_5 inst_cell_82_35 (.BL(BL35),.BLN(BLN35),.WL(WL82));
sram_cell_6t_5 inst_cell_82_36 (.BL(BL36),.BLN(BLN36),.WL(WL82));
sram_cell_6t_5 inst_cell_82_37 (.BL(BL37),.BLN(BLN37),.WL(WL82));
sram_cell_6t_5 inst_cell_82_38 (.BL(BL38),.BLN(BLN38),.WL(WL82));
sram_cell_6t_5 inst_cell_82_39 (.BL(BL39),.BLN(BLN39),.WL(WL82));
sram_cell_6t_5 inst_cell_82_40 (.BL(BL40),.BLN(BLN40),.WL(WL82));
sram_cell_6t_5 inst_cell_82_41 (.BL(BL41),.BLN(BLN41),.WL(WL82));
sram_cell_6t_5 inst_cell_82_42 (.BL(BL42),.BLN(BLN42),.WL(WL82));
sram_cell_6t_5 inst_cell_82_43 (.BL(BL43),.BLN(BLN43),.WL(WL82));
sram_cell_6t_5 inst_cell_82_44 (.BL(BL44),.BLN(BLN44),.WL(WL82));
sram_cell_6t_5 inst_cell_82_45 (.BL(BL45),.BLN(BLN45),.WL(WL82));
sram_cell_6t_5 inst_cell_82_46 (.BL(BL46),.BLN(BLN46),.WL(WL82));
sram_cell_6t_5 inst_cell_82_47 (.BL(BL47),.BLN(BLN47),.WL(WL82));
sram_cell_6t_5 inst_cell_82_48 (.BL(BL48),.BLN(BLN48),.WL(WL82));
sram_cell_6t_5 inst_cell_82_49 (.BL(BL49),.BLN(BLN49),.WL(WL82));
sram_cell_6t_5 inst_cell_82_50 (.BL(BL50),.BLN(BLN50),.WL(WL82));
sram_cell_6t_5 inst_cell_82_51 (.BL(BL51),.BLN(BLN51),.WL(WL82));
sram_cell_6t_5 inst_cell_82_52 (.BL(BL52),.BLN(BLN52),.WL(WL82));
sram_cell_6t_5 inst_cell_82_53 (.BL(BL53),.BLN(BLN53),.WL(WL82));
sram_cell_6t_5 inst_cell_82_54 (.BL(BL54),.BLN(BLN54),.WL(WL82));
sram_cell_6t_5 inst_cell_82_55 (.BL(BL55),.BLN(BLN55),.WL(WL82));
sram_cell_6t_5 inst_cell_82_56 (.BL(BL56),.BLN(BLN56),.WL(WL82));
sram_cell_6t_5 inst_cell_82_57 (.BL(BL57),.BLN(BLN57),.WL(WL82));
sram_cell_6t_5 inst_cell_82_58 (.BL(BL58),.BLN(BLN58),.WL(WL82));
sram_cell_6t_5 inst_cell_82_59 (.BL(BL59),.BLN(BLN59),.WL(WL82));
sram_cell_6t_5 inst_cell_82_60 (.BL(BL60),.BLN(BLN60),.WL(WL82));
sram_cell_6t_5 inst_cell_82_61 (.BL(BL61),.BLN(BLN61),.WL(WL82));
sram_cell_6t_5 inst_cell_82_62 (.BL(BL62),.BLN(BLN62),.WL(WL82));
sram_cell_6t_5 inst_cell_82_63 (.BL(BL63),.BLN(BLN63),.WL(WL82));
sram_cell_6t_5 inst_cell_82_64 (.BL(BL64),.BLN(BLN64),.WL(WL82));
sram_cell_6t_5 inst_cell_82_65 (.BL(BL65),.BLN(BLN65),.WL(WL82));
sram_cell_6t_5 inst_cell_82_66 (.BL(BL66),.BLN(BLN66),.WL(WL82));
sram_cell_6t_5 inst_cell_82_67 (.BL(BL67),.BLN(BLN67),.WL(WL82));
sram_cell_6t_5 inst_cell_82_68 (.BL(BL68),.BLN(BLN68),.WL(WL82));
sram_cell_6t_5 inst_cell_82_69 (.BL(BL69),.BLN(BLN69),.WL(WL82));
sram_cell_6t_5 inst_cell_82_70 (.BL(BL70),.BLN(BLN70),.WL(WL82));
sram_cell_6t_5 inst_cell_82_71 (.BL(BL71),.BLN(BLN71),.WL(WL82));
sram_cell_6t_5 inst_cell_82_72 (.BL(BL72),.BLN(BLN72),.WL(WL82));
sram_cell_6t_5 inst_cell_82_73 (.BL(BL73),.BLN(BLN73),.WL(WL82));
sram_cell_6t_5 inst_cell_82_74 (.BL(BL74),.BLN(BLN74),.WL(WL82));
sram_cell_6t_5 inst_cell_82_75 (.BL(BL75),.BLN(BLN75),.WL(WL82));
sram_cell_6t_5 inst_cell_82_76 (.BL(BL76),.BLN(BLN76),.WL(WL82));
sram_cell_6t_5 inst_cell_82_77 (.BL(BL77),.BLN(BLN77),.WL(WL82));
sram_cell_6t_5 inst_cell_82_78 (.BL(BL78),.BLN(BLN78),.WL(WL82));
sram_cell_6t_5 inst_cell_82_79 (.BL(BL79),.BLN(BLN79),.WL(WL82));
sram_cell_6t_5 inst_cell_82_80 (.BL(BL80),.BLN(BLN80),.WL(WL82));
sram_cell_6t_5 inst_cell_82_81 (.BL(BL81),.BLN(BLN81),.WL(WL82));
sram_cell_6t_5 inst_cell_82_82 (.BL(BL82),.BLN(BLN82),.WL(WL82));
sram_cell_6t_5 inst_cell_82_83 (.BL(BL83),.BLN(BLN83),.WL(WL82));
sram_cell_6t_5 inst_cell_82_84 (.BL(BL84),.BLN(BLN84),.WL(WL82));
sram_cell_6t_5 inst_cell_82_85 (.BL(BL85),.BLN(BLN85),.WL(WL82));
sram_cell_6t_5 inst_cell_82_86 (.BL(BL86),.BLN(BLN86),.WL(WL82));
sram_cell_6t_5 inst_cell_82_87 (.BL(BL87),.BLN(BLN87),.WL(WL82));
sram_cell_6t_5 inst_cell_82_88 (.BL(BL88),.BLN(BLN88),.WL(WL82));
sram_cell_6t_5 inst_cell_82_89 (.BL(BL89),.BLN(BLN89),.WL(WL82));
sram_cell_6t_5 inst_cell_82_90 (.BL(BL90),.BLN(BLN90),.WL(WL82));
sram_cell_6t_5 inst_cell_82_91 (.BL(BL91),.BLN(BLN91),.WL(WL82));
sram_cell_6t_5 inst_cell_82_92 (.BL(BL92),.BLN(BLN92),.WL(WL82));
sram_cell_6t_5 inst_cell_82_93 (.BL(BL93),.BLN(BLN93),.WL(WL82));
sram_cell_6t_5 inst_cell_82_94 (.BL(BL94),.BLN(BLN94),.WL(WL82));
sram_cell_6t_5 inst_cell_82_95 (.BL(BL95),.BLN(BLN95),.WL(WL82));
sram_cell_6t_5 inst_cell_82_96 (.BL(BL96),.BLN(BLN96),.WL(WL82));
sram_cell_6t_5 inst_cell_82_97 (.BL(BL97),.BLN(BLN97),.WL(WL82));
sram_cell_6t_5 inst_cell_82_98 (.BL(BL98),.BLN(BLN98),.WL(WL82));
sram_cell_6t_5 inst_cell_82_99 (.BL(BL99),.BLN(BLN99),.WL(WL82));
sram_cell_6t_5 inst_cell_82_100 (.BL(BL100),.BLN(BLN100),.WL(WL82));
sram_cell_6t_5 inst_cell_82_101 (.BL(BL101),.BLN(BLN101),.WL(WL82));
sram_cell_6t_5 inst_cell_82_102 (.BL(BL102),.BLN(BLN102),.WL(WL82));
sram_cell_6t_5 inst_cell_82_103 (.BL(BL103),.BLN(BLN103),.WL(WL82));
sram_cell_6t_5 inst_cell_82_104 (.BL(BL104),.BLN(BLN104),.WL(WL82));
sram_cell_6t_5 inst_cell_82_105 (.BL(BL105),.BLN(BLN105),.WL(WL82));
sram_cell_6t_5 inst_cell_82_106 (.BL(BL106),.BLN(BLN106),.WL(WL82));
sram_cell_6t_5 inst_cell_82_107 (.BL(BL107),.BLN(BLN107),.WL(WL82));
sram_cell_6t_5 inst_cell_82_108 (.BL(BL108),.BLN(BLN108),.WL(WL82));
sram_cell_6t_5 inst_cell_82_109 (.BL(BL109),.BLN(BLN109),.WL(WL82));
sram_cell_6t_5 inst_cell_82_110 (.BL(BL110),.BLN(BLN110),.WL(WL82));
sram_cell_6t_5 inst_cell_82_111 (.BL(BL111),.BLN(BLN111),.WL(WL82));
sram_cell_6t_5 inst_cell_82_112 (.BL(BL112),.BLN(BLN112),.WL(WL82));
sram_cell_6t_5 inst_cell_82_113 (.BL(BL113),.BLN(BLN113),.WL(WL82));
sram_cell_6t_5 inst_cell_82_114 (.BL(BL114),.BLN(BLN114),.WL(WL82));
sram_cell_6t_5 inst_cell_82_115 (.BL(BL115),.BLN(BLN115),.WL(WL82));
sram_cell_6t_5 inst_cell_82_116 (.BL(BL116),.BLN(BLN116),.WL(WL82));
sram_cell_6t_5 inst_cell_82_117 (.BL(BL117),.BLN(BLN117),.WL(WL82));
sram_cell_6t_5 inst_cell_82_118 (.BL(BL118),.BLN(BLN118),.WL(WL82));
sram_cell_6t_5 inst_cell_82_119 (.BL(BL119),.BLN(BLN119),.WL(WL82));
sram_cell_6t_5 inst_cell_82_120 (.BL(BL120),.BLN(BLN120),.WL(WL82));
sram_cell_6t_5 inst_cell_82_121 (.BL(BL121),.BLN(BLN121),.WL(WL82));
sram_cell_6t_5 inst_cell_82_122 (.BL(BL122),.BLN(BLN122),.WL(WL82));
sram_cell_6t_5 inst_cell_82_123 (.BL(BL123),.BLN(BLN123),.WL(WL82));
sram_cell_6t_5 inst_cell_82_124 (.BL(BL124),.BLN(BLN124),.WL(WL82));
sram_cell_6t_5 inst_cell_82_125 (.BL(BL125),.BLN(BLN125),.WL(WL82));
sram_cell_6t_5 inst_cell_82_126 (.BL(BL126),.BLN(BLN126),.WL(WL82));
sram_cell_6t_5 inst_cell_82_127 (.BL(BL127),.BLN(BLN127),.WL(WL82));
sram_cell_6t_5 inst_cell_83_0 (.BL(BL0),.BLN(BLN0),.WL(WL83));
sram_cell_6t_5 inst_cell_83_1 (.BL(BL1),.BLN(BLN1),.WL(WL83));
sram_cell_6t_5 inst_cell_83_2 (.BL(BL2),.BLN(BLN2),.WL(WL83));
sram_cell_6t_5 inst_cell_83_3 (.BL(BL3),.BLN(BLN3),.WL(WL83));
sram_cell_6t_5 inst_cell_83_4 (.BL(BL4),.BLN(BLN4),.WL(WL83));
sram_cell_6t_5 inst_cell_83_5 (.BL(BL5),.BLN(BLN5),.WL(WL83));
sram_cell_6t_5 inst_cell_83_6 (.BL(BL6),.BLN(BLN6),.WL(WL83));
sram_cell_6t_5 inst_cell_83_7 (.BL(BL7),.BLN(BLN7),.WL(WL83));
sram_cell_6t_5 inst_cell_83_8 (.BL(BL8),.BLN(BLN8),.WL(WL83));
sram_cell_6t_5 inst_cell_83_9 (.BL(BL9),.BLN(BLN9),.WL(WL83));
sram_cell_6t_5 inst_cell_83_10 (.BL(BL10),.BLN(BLN10),.WL(WL83));
sram_cell_6t_5 inst_cell_83_11 (.BL(BL11),.BLN(BLN11),.WL(WL83));
sram_cell_6t_5 inst_cell_83_12 (.BL(BL12),.BLN(BLN12),.WL(WL83));
sram_cell_6t_5 inst_cell_83_13 (.BL(BL13),.BLN(BLN13),.WL(WL83));
sram_cell_6t_5 inst_cell_83_14 (.BL(BL14),.BLN(BLN14),.WL(WL83));
sram_cell_6t_5 inst_cell_83_15 (.BL(BL15),.BLN(BLN15),.WL(WL83));
sram_cell_6t_5 inst_cell_83_16 (.BL(BL16),.BLN(BLN16),.WL(WL83));
sram_cell_6t_5 inst_cell_83_17 (.BL(BL17),.BLN(BLN17),.WL(WL83));
sram_cell_6t_5 inst_cell_83_18 (.BL(BL18),.BLN(BLN18),.WL(WL83));
sram_cell_6t_5 inst_cell_83_19 (.BL(BL19),.BLN(BLN19),.WL(WL83));
sram_cell_6t_5 inst_cell_83_20 (.BL(BL20),.BLN(BLN20),.WL(WL83));
sram_cell_6t_5 inst_cell_83_21 (.BL(BL21),.BLN(BLN21),.WL(WL83));
sram_cell_6t_5 inst_cell_83_22 (.BL(BL22),.BLN(BLN22),.WL(WL83));
sram_cell_6t_5 inst_cell_83_23 (.BL(BL23),.BLN(BLN23),.WL(WL83));
sram_cell_6t_5 inst_cell_83_24 (.BL(BL24),.BLN(BLN24),.WL(WL83));
sram_cell_6t_5 inst_cell_83_25 (.BL(BL25),.BLN(BLN25),.WL(WL83));
sram_cell_6t_5 inst_cell_83_26 (.BL(BL26),.BLN(BLN26),.WL(WL83));
sram_cell_6t_5 inst_cell_83_27 (.BL(BL27),.BLN(BLN27),.WL(WL83));
sram_cell_6t_5 inst_cell_83_28 (.BL(BL28),.BLN(BLN28),.WL(WL83));
sram_cell_6t_5 inst_cell_83_29 (.BL(BL29),.BLN(BLN29),.WL(WL83));
sram_cell_6t_5 inst_cell_83_30 (.BL(BL30),.BLN(BLN30),.WL(WL83));
sram_cell_6t_5 inst_cell_83_31 (.BL(BL31),.BLN(BLN31),.WL(WL83));
sram_cell_6t_5 inst_cell_83_32 (.BL(BL32),.BLN(BLN32),.WL(WL83));
sram_cell_6t_5 inst_cell_83_33 (.BL(BL33),.BLN(BLN33),.WL(WL83));
sram_cell_6t_5 inst_cell_83_34 (.BL(BL34),.BLN(BLN34),.WL(WL83));
sram_cell_6t_5 inst_cell_83_35 (.BL(BL35),.BLN(BLN35),.WL(WL83));
sram_cell_6t_5 inst_cell_83_36 (.BL(BL36),.BLN(BLN36),.WL(WL83));
sram_cell_6t_5 inst_cell_83_37 (.BL(BL37),.BLN(BLN37),.WL(WL83));
sram_cell_6t_5 inst_cell_83_38 (.BL(BL38),.BLN(BLN38),.WL(WL83));
sram_cell_6t_5 inst_cell_83_39 (.BL(BL39),.BLN(BLN39),.WL(WL83));
sram_cell_6t_5 inst_cell_83_40 (.BL(BL40),.BLN(BLN40),.WL(WL83));
sram_cell_6t_5 inst_cell_83_41 (.BL(BL41),.BLN(BLN41),.WL(WL83));
sram_cell_6t_5 inst_cell_83_42 (.BL(BL42),.BLN(BLN42),.WL(WL83));
sram_cell_6t_5 inst_cell_83_43 (.BL(BL43),.BLN(BLN43),.WL(WL83));
sram_cell_6t_5 inst_cell_83_44 (.BL(BL44),.BLN(BLN44),.WL(WL83));
sram_cell_6t_5 inst_cell_83_45 (.BL(BL45),.BLN(BLN45),.WL(WL83));
sram_cell_6t_5 inst_cell_83_46 (.BL(BL46),.BLN(BLN46),.WL(WL83));
sram_cell_6t_5 inst_cell_83_47 (.BL(BL47),.BLN(BLN47),.WL(WL83));
sram_cell_6t_5 inst_cell_83_48 (.BL(BL48),.BLN(BLN48),.WL(WL83));
sram_cell_6t_5 inst_cell_83_49 (.BL(BL49),.BLN(BLN49),.WL(WL83));
sram_cell_6t_5 inst_cell_83_50 (.BL(BL50),.BLN(BLN50),.WL(WL83));
sram_cell_6t_5 inst_cell_83_51 (.BL(BL51),.BLN(BLN51),.WL(WL83));
sram_cell_6t_5 inst_cell_83_52 (.BL(BL52),.BLN(BLN52),.WL(WL83));
sram_cell_6t_5 inst_cell_83_53 (.BL(BL53),.BLN(BLN53),.WL(WL83));
sram_cell_6t_5 inst_cell_83_54 (.BL(BL54),.BLN(BLN54),.WL(WL83));
sram_cell_6t_5 inst_cell_83_55 (.BL(BL55),.BLN(BLN55),.WL(WL83));
sram_cell_6t_5 inst_cell_83_56 (.BL(BL56),.BLN(BLN56),.WL(WL83));
sram_cell_6t_5 inst_cell_83_57 (.BL(BL57),.BLN(BLN57),.WL(WL83));
sram_cell_6t_5 inst_cell_83_58 (.BL(BL58),.BLN(BLN58),.WL(WL83));
sram_cell_6t_5 inst_cell_83_59 (.BL(BL59),.BLN(BLN59),.WL(WL83));
sram_cell_6t_5 inst_cell_83_60 (.BL(BL60),.BLN(BLN60),.WL(WL83));
sram_cell_6t_5 inst_cell_83_61 (.BL(BL61),.BLN(BLN61),.WL(WL83));
sram_cell_6t_5 inst_cell_83_62 (.BL(BL62),.BLN(BLN62),.WL(WL83));
sram_cell_6t_5 inst_cell_83_63 (.BL(BL63),.BLN(BLN63),.WL(WL83));
sram_cell_6t_5 inst_cell_83_64 (.BL(BL64),.BLN(BLN64),.WL(WL83));
sram_cell_6t_5 inst_cell_83_65 (.BL(BL65),.BLN(BLN65),.WL(WL83));
sram_cell_6t_5 inst_cell_83_66 (.BL(BL66),.BLN(BLN66),.WL(WL83));
sram_cell_6t_5 inst_cell_83_67 (.BL(BL67),.BLN(BLN67),.WL(WL83));
sram_cell_6t_5 inst_cell_83_68 (.BL(BL68),.BLN(BLN68),.WL(WL83));
sram_cell_6t_5 inst_cell_83_69 (.BL(BL69),.BLN(BLN69),.WL(WL83));
sram_cell_6t_5 inst_cell_83_70 (.BL(BL70),.BLN(BLN70),.WL(WL83));
sram_cell_6t_5 inst_cell_83_71 (.BL(BL71),.BLN(BLN71),.WL(WL83));
sram_cell_6t_5 inst_cell_83_72 (.BL(BL72),.BLN(BLN72),.WL(WL83));
sram_cell_6t_5 inst_cell_83_73 (.BL(BL73),.BLN(BLN73),.WL(WL83));
sram_cell_6t_5 inst_cell_83_74 (.BL(BL74),.BLN(BLN74),.WL(WL83));
sram_cell_6t_5 inst_cell_83_75 (.BL(BL75),.BLN(BLN75),.WL(WL83));
sram_cell_6t_5 inst_cell_83_76 (.BL(BL76),.BLN(BLN76),.WL(WL83));
sram_cell_6t_5 inst_cell_83_77 (.BL(BL77),.BLN(BLN77),.WL(WL83));
sram_cell_6t_5 inst_cell_83_78 (.BL(BL78),.BLN(BLN78),.WL(WL83));
sram_cell_6t_5 inst_cell_83_79 (.BL(BL79),.BLN(BLN79),.WL(WL83));
sram_cell_6t_5 inst_cell_83_80 (.BL(BL80),.BLN(BLN80),.WL(WL83));
sram_cell_6t_5 inst_cell_83_81 (.BL(BL81),.BLN(BLN81),.WL(WL83));
sram_cell_6t_5 inst_cell_83_82 (.BL(BL82),.BLN(BLN82),.WL(WL83));
sram_cell_6t_5 inst_cell_83_83 (.BL(BL83),.BLN(BLN83),.WL(WL83));
sram_cell_6t_5 inst_cell_83_84 (.BL(BL84),.BLN(BLN84),.WL(WL83));
sram_cell_6t_5 inst_cell_83_85 (.BL(BL85),.BLN(BLN85),.WL(WL83));
sram_cell_6t_5 inst_cell_83_86 (.BL(BL86),.BLN(BLN86),.WL(WL83));
sram_cell_6t_5 inst_cell_83_87 (.BL(BL87),.BLN(BLN87),.WL(WL83));
sram_cell_6t_5 inst_cell_83_88 (.BL(BL88),.BLN(BLN88),.WL(WL83));
sram_cell_6t_5 inst_cell_83_89 (.BL(BL89),.BLN(BLN89),.WL(WL83));
sram_cell_6t_5 inst_cell_83_90 (.BL(BL90),.BLN(BLN90),.WL(WL83));
sram_cell_6t_5 inst_cell_83_91 (.BL(BL91),.BLN(BLN91),.WL(WL83));
sram_cell_6t_5 inst_cell_83_92 (.BL(BL92),.BLN(BLN92),.WL(WL83));
sram_cell_6t_5 inst_cell_83_93 (.BL(BL93),.BLN(BLN93),.WL(WL83));
sram_cell_6t_5 inst_cell_83_94 (.BL(BL94),.BLN(BLN94),.WL(WL83));
sram_cell_6t_5 inst_cell_83_95 (.BL(BL95),.BLN(BLN95),.WL(WL83));
sram_cell_6t_5 inst_cell_83_96 (.BL(BL96),.BLN(BLN96),.WL(WL83));
sram_cell_6t_5 inst_cell_83_97 (.BL(BL97),.BLN(BLN97),.WL(WL83));
sram_cell_6t_5 inst_cell_83_98 (.BL(BL98),.BLN(BLN98),.WL(WL83));
sram_cell_6t_5 inst_cell_83_99 (.BL(BL99),.BLN(BLN99),.WL(WL83));
sram_cell_6t_5 inst_cell_83_100 (.BL(BL100),.BLN(BLN100),.WL(WL83));
sram_cell_6t_5 inst_cell_83_101 (.BL(BL101),.BLN(BLN101),.WL(WL83));
sram_cell_6t_5 inst_cell_83_102 (.BL(BL102),.BLN(BLN102),.WL(WL83));
sram_cell_6t_5 inst_cell_83_103 (.BL(BL103),.BLN(BLN103),.WL(WL83));
sram_cell_6t_5 inst_cell_83_104 (.BL(BL104),.BLN(BLN104),.WL(WL83));
sram_cell_6t_5 inst_cell_83_105 (.BL(BL105),.BLN(BLN105),.WL(WL83));
sram_cell_6t_5 inst_cell_83_106 (.BL(BL106),.BLN(BLN106),.WL(WL83));
sram_cell_6t_5 inst_cell_83_107 (.BL(BL107),.BLN(BLN107),.WL(WL83));
sram_cell_6t_5 inst_cell_83_108 (.BL(BL108),.BLN(BLN108),.WL(WL83));
sram_cell_6t_5 inst_cell_83_109 (.BL(BL109),.BLN(BLN109),.WL(WL83));
sram_cell_6t_5 inst_cell_83_110 (.BL(BL110),.BLN(BLN110),.WL(WL83));
sram_cell_6t_5 inst_cell_83_111 (.BL(BL111),.BLN(BLN111),.WL(WL83));
sram_cell_6t_5 inst_cell_83_112 (.BL(BL112),.BLN(BLN112),.WL(WL83));
sram_cell_6t_5 inst_cell_83_113 (.BL(BL113),.BLN(BLN113),.WL(WL83));
sram_cell_6t_5 inst_cell_83_114 (.BL(BL114),.BLN(BLN114),.WL(WL83));
sram_cell_6t_5 inst_cell_83_115 (.BL(BL115),.BLN(BLN115),.WL(WL83));
sram_cell_6t_5 inst_cell_83_116 (.BL(BL116),.BLN(BLN116),.WL(WL83));
sram_cell_6t_5 inst_cell_83_117 (.BL(BL117),.BLN(BLN117),.WL(WL83));
sram_cell_6t_5 inst_cell_83_118 (.BL(BL118),.BLN(BLN118),.WL(WL83));
sram_cell_6t_5 inst_cell_83_119 (.BL(BL119),.BLN(BLN119),.WL(WL83));
sram_cell_6t_5 inst_cell_83_120 (.BL(BL120),.BLN(BLN120),.WL(WL83));
sram_cell_6t_5 inst_cell_83_121 (.BL(BL121),.BLN(BLN121),.WL(WL83));
sram_cell_6t_5 inst_cell_83_122 (.BL(BL122),.BLN(BLN122),.WL(WL83));
sram_cell_6t_5 inst_cell_83_123 (.BL(BL123),.BLN(BLN123),.WL(WL83));
sram_cell_6t_5 inst_cell_83_124 (.BL(BL124),.BLN(BLN124),.WL(WL83));
sram_cell_6t_5 inst_cell_83_125 (.BL(BL125),.BLN(BLN125),.WL(WL83));
sram_cell_6t_5 inst_cell_83_126 (.BL(BL126),.BLN(BLN126),.WL(WL83));
sram_cell_6t_5 inst_cell_83_127 (.BL(BL127),.BLN(BLN127),.WL(WL83));
sram_cell_6t_5 inst_cell_84_0 (.BL(BL0),.BLN(BLN0),.WL(WL84));
sram_cell_6t_5 inst_cell_84_1 (.BL(BL1),.BLN(BLN1),.WL(WL84));
sram_cell_6t_5 inst_cell_84_2 (.BL(BL2),.BLN(BLN2),.WL(WL84));
sram_cell_6t_5 inst_cell_84_3 (.BL(BL3),.BLN(BLN3),.WL(WL84));
sram_cell_6t_5 inst_cell_84_4 (.BL(BL4),.BLN(BLN4),.WL(WL84));
sram_cell_6t_5 inst_cell_84_5 (.BL(BL5),.BLN(BLN5),.WL(WL84));
sram_cell_6t_5 inst_cell_84_6 (.BL(BL6),.BLN(BLN6),.WL(WL84));
sram_cell_6t_5 inst_cell_84_7 (.BL(BL7),.BLN(BLN7),.WL(WL84));
sram_cell_6t_5 inst_cell_84_8 (.BL(BL8),.BLN(BLN8),.WL(WL84));
sram_cell_6t_5 inst_cell_84_9 (.BL(BL9),.BLN(BLN9),.WL(WL84));
sram_cell_6t_5 inst_cell_84_10 (.BL(BL10),.BLN(BLN10),.WL(WL84));
sram_cell_6t_5 inst_cell_84_11 (.BL(BL11),.BLN(BLN11),.WL(WL84));
sram_cell_6t_5 inst_cell_84_12 (.BL(BL12),.BLN(BLN12),.WL(WL84));
sram_cell_6t_5 inst_cell_84_13 (.BL(BL13),.BLN(BLN13),.WL(WL84));
sram_cell_6t_5 inst_cell_84_14 (.BL(BL14),.BLN(BLN14),.WL(WL84));
sram_cell_6t_5 inst_cell_84_15 (.BL(BL15),.BLN(BLN15),.WL(WL84));
sram_cell_6t_5 inst_cell_84_16 (.BL(BL16),.BLN(BLN16),.WL(WL84));
sram_cell_6t_5 inst_cell_84_17 (.BL(BL17),.BLN(BLN17),.WL(WL84));
sram_cell_6t_5 inst_cell_84_18 (.BL(BL18),.BLN(BLN18),.WL(WL84));
sram_cell_6t_5 inst_cell_84_19 (.BL(BL19),.BLN(BLN19),.WL(WL84));
sram_cell_6t_5 inst_cell_84_20 (.BL(BL20),.BLN(BLN20),.WL(WL84));
sram_cell_6t_5 inst_cell_84_21 (.BL(BL21),.BLN(BLN21),.WL(WL84));
sram_cell_6t_5 inst_cell_84_22 (.BL(BL22),.BLN(BLN22),.WL(WL84));
sram_cell_6t_5 inst_cell_84_23 (.BL(BL23),.BLN(BLN23),.WL(WL84));
sram_cell_6t_5 inst_cell_84_24 (.BL(BL24),.BLN(BLN24),.WL(WL84));
sram_cell_6t_5 inst_cell_84_25 (.BL(BL25),.BLN(BLN25),.WL(WL84));
sram_cell_6t_5 inst_cell_84_26 (.BL(BL26),.BLN(BLN26),.WL(WL84));
sram_cell_6t_5 inst_cell_84_27 (.BL(BL27),.BLN(BLN27),.WL(WL84));
sram_cell_6t_5 inst_cell_84_28 (.BL(BL28),.BLN(BLN28),.WL(WL84));
sram_cell_6t_5 inst_cell_84_29 (.BL(BL29),.BLN(BLN29),.WL(WL84));
sram_cell_6t_5 inst_cell_84_30 (.BL(BL30),.BLN(BLN30),.WL(WL84));
sram_cell_6t_5 inst_cell_84_31 (.BL(BL31),.BLN(BLN31),.WL(WL84));
sram_cell_6t_5 inst_cell_84_32 (.BL(BL32),.BLN(BLN32),.WL(WL84));
sram_cell_6t_5 inst_cell_84_33 (.BL(BL33),.BLN(BLN33),.WL(WL84));
sram_cell_6t_5 inst_cell_84_34 (.BL(BL34),.BLN(BLN34),.WL(WL84));
sram_cell_6t_5 inst_cell_84_35 (.BL(BL35),.BLN(BLN35),.WL(WL84));
sram_cell_6t_5 inst_cell_84_36 (.BL(BL36),.BLN(BLN36),.WL(WL84));
sram_cell_6t_5 inst_cell_84_37 (.BL(BL37),.BLN(BLN37),.WL(WL84));
sram_cell_6t_5 inst_cell_84_38 (.BL(BL38),.BLN(BLN38),.WL(WL84));
sram_cell_6t_5 inst_cell_84_39 (.BL(BL39),.BLN(BLN39),.WL(WL84));
sram_cell_6t_5 inst_cell_84_40 (.BL(BL40),.BLN(BLN40),.WL(WL84));
sram_cell_6t_5 inst_cell_84_41 (.BL(BL41),.BLN(BLN41),.WL(WL84));
sram_cell_6t_5 inst_cell_84_42 (.BL(BL42),.BLN(BLN42),.WL(WL84));
sram_cell_6t_5 inst_cell_84_43 (.BL(BL43),.BLN(BLN43),.WL(WL84));
sram_cell_6t_5 inst_cell_84_44 (.BL(BL44),.BLN(BLN44),.WL(WL84));
sram_cell_6t_5 inst_cell_84_45 (.BL(BL45),.BLN(BLN45),.WL(WL84));
sram_cell_6t_5 inst_cell_84_46 (.BL(BL46),.BLN(BLN46),.WL(WL84));
sram_cell_6t_5 inst_cell_84_47 (.BL(BL47),.BLN(BLN47),.WL(WL84));
sram_cell_6t_5 inst_cell_84_48 (.BL(BL48),.BLN(BLN48),.WL(WL84));
sram_cell_6t_5 inst_cell_84_49 (.BL(BL49),.BLN(BLN49),.WL(WL84));
sram_cell_6t_5 inst_cell_84_50 (.BL(BL50),.BLN(BLN50),.WL(WL84));
sram_cell_6t_5 inst_cell_84_51 (.BL(BL51),.BLN(BLN51),.WL(WL84));
sram_cell_6t_5 inst_cell_84_52 (.BL(BL52),.BLN(BLN52),.WL(WL84));
sram_cell_6t_5 inst_cell_84_53 (.BL(BL53),.BLN(BLN53),.WL(WL84));
sram_cell_6t_5 inst_cell_84_54 (.BL(BL54),.BLN(BLN54),.WL(WL84));
sram_cell_6t_5 inst_cell_84_55 (.BL(BL55),.BLN(BLN55),.WL(WL84));
sram_cell_6t_5 inst_cell_84_56 (.BL(BL56),.BLN(BLN56),.WL(WL84));
sram_cell_6t_5 inst_cell_84_57 (.BL(BL57),.BLN(BLN57),.WL(WL84));
sram_cell_6t_5 inst_cell_84_58 (.BL(BL58),.BLN(BLN58),.WL(WL84));
sram_cell_6t_5 inst_cell_84_59 (.BL(BL59),.BLN(BLN59),.WL(WL84));
sram_cell_6t_5 inst_cell_84_60 (.BL(BL60),.BLN(BLN60),.WL(WL84));
sram_cell_6t_5 inst_cell_84_61 (.BL(BL61),.BLN(BLN61),.WL(WL84));
sram_cell_6t_5 inst_cell_84_62 (.BL(BL62),.BLN(BLN62),.WL(WL84));
sram_cell_6t_5 inst_cell_84_63 (.BL(BL63),.BLN(BLN63),.WL(WL84));
sram_cell_6t_5 inst_cell_84_64 (.BL(BL64),.BLN(BLN64),.WL(WL84));
sram_cell_6t_5 inst_cell_84_65 (.BL(BL65),.BLN(BLN65),.WL(WL84));
sram_cell_6t_5 inst_cell_84_66 (.BL(BL66),.BLN(BLN66),.WL(WL84));
sram_cell_6t_5 inst_cell_84_67 (.BL(BL67),.BLN(BLN67),.WL(WL84));
sram_cell_6t_5 inst_cell_84_68 (.BL(BL68),.BLN(BLN68),.WL(WL84));
sram_cell_6t_5 inst_cell_84_69 (.BL(BL69),.BLN(BLN69),.WL(WL84));
sram_cell_6t_5 inst_cell_84_70 (.BL(BL70),.BLN(BLN70),.WL(WL84));
sram_cell_6t_5 inst_cell_84_71 (.BL(BL71),.BLN(BLN71),.WL(WL84));
sram_cell_6t_5 inst_cell_84_72 (.BL(BL72),.BLN(BLN72),.WL(WL84));
sram_cell_6t_5 inst_cell_84_73 (.BL(BL73),.BLN(BLN73),.WL(WL84));
sram_cell_6t_5 inst_cell_84_74 (.BL(BL74),.BLN(BLN74),.WL(WL84));
sram_cell_6t_5 inst_cell_84_75 (.BL(BL75),.BLN(BLN75),.WL(WL84));
sram_cell_6t_5 inst_cell_84_76 (.BL(BL76),.BLN(BLN76),.WL(WL84));
sram_cell_6t_5 inst_cell_84_77 (.BL(BL77),.BLN(BLN77),.WL(WL84));
sram_cell_6t_5 inst_cell_84_78 (.BL(BL78),.BLN(BLN78),.WL(WL84));
sram_cell_6t_5 inst_cell_84_79 (.BL(BL79),.BLN(BLN79),.WL(WL84));
sram_cell_6t_5 inst_cell_84_80 (.BL(BL80),.BLN(BLN80),.WL(WL84));
sram_cell_6t_5 inst_cell_84_81 (.BL(BL81),.BLN(BLN81),.WL(WL84));
sram_cell_6t_5 inst_cell_84_82 (.BL(BL82),.BLN(BLN82),.WL(WL84));
sram_cell_6t_5 inst_cell_84_83 (.BL(BL83),.BLN(BLN83),.WL(WL84));
sram_cell_6t_5 inst_cell_84_84 (.BL(BL84),.BLN(BLN84),.WL(WL84));
sram_cell_6t_5 inst_cell_84_85 (.BL(BL85),.BLN(BLN85),.WL(WL84));
sram_cell_6t_5 inst_cell_84_86 (.BL(BL86),.BLN(BLN86),.WL(WL84));
sram_cell_6t_5 inst_cell_84_87 (.BL(BL87),.BLN(BLN87),.WL(WL84));
sram_cell_6t_5 inst_cell_84_88 (.BL(BL88),.BLN(BLN88),.WL(WL84));
sram_cell_6t_5 inst_cell_84_89 (.BL(BL89),.BLN(BLN89),.WL(WL84));
sram_cell_6t_5 inst_cell_84_90 (.BL(BL90),.BLN(BLN90),.WL(WL84));
sram_cell_6t_5 inst_cell_84_91 (.BL(BL91),.BLN(BLN91),.WL(WL84));
sram_cell_6t_5 inst_cell_84_92 (.BL(BL92),.BLN(BLN92),.WL(WL84));
sram_cell_6t_5 inst_cell_84_93 (.BL(BL93),.BLN(BLN93),.WL(WL84));
sram_cell_6t_5 inst_cell_84_94 (.BL(BL94),.BLN(BLN94),.WL(WL84));
sram_cell_6t_5 inst_cell_84_95 (.BL(BL95),.BLN(BLN95),.WL(WL84));
sram_cell_6t_5 inst_cell_84_96 (.BL(BL96),.BLN(BLN96),.WL(WL84));
sram_cell_6t_5 inst_cell_84_97 (.BL(BL97),.BLN(BLN97),.WL(WL84));
sram_cell_6t_5 inst_cell_84_98 (.BL(BL98),.BLN(BLN98),.WL(WL84));
sram_cell_6t_5 inst_cell_84_99 (.BL(BL99),.BLN(BLN99),.WL(WL84));
sram_cell_6t_5 inst_cell_84_100 (.BL(BL100),.BLN(BLN100),.WL(WL84));
sram_cell_6t_5 inst_cell_84_101 (.BL(BL101),.BLN(BLN101),.WL(WL84));
sram_cell_6t_5 inst_cell_84_102 (.BL(BL102),.BLN(BLN102),.WL(WL84));
sram_cell_6t_5 inst_cell_84_103 (.BL(BL103),.BLN(BLN103),.WL(WL84));
sram_cell_6t_5 inst_cell_84_104 (.BL(BL104),.BLN(BLN104),.WL(WL84));
sram_cell_6t_5 inst_cell_84_105 (.BL(BL105),.BLN(BLN105),.WL(WL84));
sram_cell_6t_5 inst_cell_84_106 (.BL(BL106),.BLN(BLN106),.WL(WL84));
sram_cell_6t_5 inst_cell_84_107 (.BL(BL107),.BLN(BLN107),.WL(WL84));
sram_cell_6t_5 inst_cell_84_108 (.BL(BL108),.BLN(BLN108),.WL(WL84));
sram_cell_6t_5 inst_cell_84_109 (.BL(BL109),.BLN(BLN109),.WL(WL84));
sram_cell_6t_5 inst_cell_84_110 (.BL(BL110),.BLN(BLN110),.WL(WL84));
sram_cell_6t_5 inst_cell_84_111 (.BL(BL111),.BLN(BLN111),.WL(WL84));
sram_cell_6t_5 inst_cell_84_112 (.BL(BL112),.BLN(BLN112),.WL(WL84));
sram_cell_6t_5 inst_cell_84_113 (.BL(BL113),.BLN(BLN113),.WL(WL84));
sram_cell_6t_5 inst_cell_84_114 (.BL(BL114),.BLN(BLN114),.WL(WL84));
sram_cell_6t_5 inst_cell_84_115 (.BL(BL115),.BLN(BLN115),.WL(WL84));
sram_cell_6t_5 inst_cell_84_116 (.BL(BL116),.BLN(BLN116),.WL(WL84));
sram_cell_6t_5 inst_cell_84_117 (.BL(BL117),.BLN(BLN117),.WL(WL84));
sram_cell_6t_5 inst_cell_84_118 (.BL(BL118),.BLN(BLN118),.WL(WL84));
sram_cell_6t_5 inst_cell_84_119 (.BL(BL119),.BLN(BLN119),.WL(WL84));
sram_cell_6t_5 inst_cell_84_120 (.BL(BL120),.BLN(BLN120),.WL(WL84));
sram_cell_6t_5 inst_cell_84_121 (.BL(BL121),.BLN(BLN121),.WL(WL84));
sram_cell_6t_5 inst_cell_84_122 (.BL(BL122),.BLN(BLN122),.WL(WL84));
sram_cell_6t_5 inst_cell_84_123 (.BL(BL123),.BLN(BLN123),.WL(WL84));
sram_cell_6t_5 inst_cell_84_124 (.BL(BL124),.BLN(BLN124),.WL(WL84));
sram_cell_6t_5 inst_cell_84_125 (.BL(BL125),.BLN(BLN125),.WL(WL84));
sram_cell_6t_5 inst_cell_84_126 (.BL(BL126),.BLN(BLN126),.WL(WL84));
sram_cell_6t_5 inst_cell_84_127 (.BL(BL127),.BLN(BLN127),.WL(WL84));
sram_cell_6t_5 inst_cell_85_0 (.BL(BL0),.BLN(BLN0),.WL(WL85));
sram_cell_6t_5 inst_cell_85_1 (.BL(BL1),.BLN(BLN1),.WL(WL85));
sram_cell_6t_5 inst_cell_85_2 (.BL(BL2),.BLN(BLN2),.WL(WL85));
sram_cell_6t_5 inst_cell_85_3 (.BL(BL3),.BLN(BLN3),.WL(WL85));
sram_cell_6t_5 inst_cell_85_4 (.BL(BL4),.BLN(BLN4),.WL(WL85));
sram_cell_6t_5 inst_cell_85_5 (.BL(BL5),.BLN(BLN5),.WL(WL85));
sram_cell_6t_5 inst_cell_85_6 (.BL(BL6),.BLN(BLN6),.WL(WL85));
sram_cell_6t_5 inst_cell_85_7 (.BL(BL7),.BLN(BLN7),.WL(WL85));
sram_cell_6t_5 inst_cell_85_8 (.BL(BL8),.BLN(BLN8),.WL(WL85));
sram_cell_6t_5 inst_cell_85_9 (.BL(BL9),.BLN(BLN9),.WL(WL85));
sram_cell_6t_5 inst_cell_85_10 (.BL(BL10),.BLN(BLN10),.WL(WL85));
sram_cell_6t_5 inst_cell_85_11 (.BL(BL11),.BLN(BLN11),.WL(WL85));
sram_cell_6t_5 inst_cell_85_12 (.BL(BL12),.BLN(BLN12),.WL(WL85));
sram_cell_6t_5 inst_cell_85_13 (.BL(BL13),.BLN(BLN13),.WL(WL85));
sram_cell_6t_5 inst_cell_85_14 (.BL(BL14),.BLN(BLN14),.WL(WL85));
sram_cell_6t_5 inst_cell_85_15 (.BL(BL15),.BLN(BLN15),.WL(WL85));
sram_cell_6t_5 inst_cell_85_16 (.BL(BL16),.BLN(BLN16),.WL(WL85));
sram_cell_6t_5 inst_cell_85_17 (.BL(BL17),.BLN(BLN17),.WL(WL85));
sram_cell_6t_5 inst_cell_85_18 (.BL(BL18),.BLN(BLN18),.WL(WL85));
sram_cell_6t_5 inst_cell_85_19 (.BL(BL19),.BLN(BLN19),.WL(WL85));
sram_cell_6t_5 inst_cell_85_20 (.BL(BL20),.BLN(BLN20),.WL(WL85));
sram_cell_6t_5 inst_cell_85_21 (.BL(BL21),.BLN(BLN21),.WL(WL85));
sram_cell_6t_5 inst_cell_85_22 (.BL(BL22),.BLN(BLN22),.WL(WL85));
sram_cell_6t_5 inst_cell_85_23 (.BL(BL23),.BLN(BLN23),.WL(WL85));
sram_cell_6t_5 inst_cell_85_24 (.BL(BL24),.BLN(BLN24),.WL(WL85));
sram_cell_6t_5 inst_cell_85_25 (.BL(BL25),.BLN(BLN25),.WL(WL85));
sram_cell_6t_5 inst_cell_85_26 (.BL(BL26),.BLN(BLN26),.WL(WL85));
sram_cell_6t_5 inst_cell_85_27 (.BL(BL27),.BLN(BLN27),.WL(WL85));
sram_cell_6t_5 inst_cell_85_28 (.BL(BL28),.BLN(BLN28),.WL(WL85));
sram_cell_6t_5 inst_cell_85_29 (.BL(BL29),.BLN(BLN29),.WL(WL85));
sram_cell_6t_5 inst_cell_85_30 (.BL(BL30),.BLN(BLN30),.WL(WL85));
sram_cell_6t_5 inst_cell_85_31 (.BL(BL31),.BLN(BLN31),.WL(WL85));
sram_cell_6t_5 inst_cell_85_32 (.BL(BL32),.BLN(BLN32),.WL(WL85));
sram_cell_6t_5 inst_cell_85_33 (.BL(BL33),.BLN(BLN33),.WL(WL85));
sram_cell_6t_5 inst_cell_85_34 (.BL(BL34),.BLN(BLN34),.WL(WL85));
sram_cell_6t_5 inst_cell_85_35 (.BL(BL35),.BLN(BLN35),.WL(WL85));
sram_cell_6t_5 inst_cell_85_36 (.BL(BL36),.BLN(BLN36),.WL(WL85));
sram_cell_6t_5 inst_cell_85_37 (.BL(BL37),.BLN(BLN37),.WL(WL85));
sram_cell_6t_5 inst_cell_85_38 (.BL(BL38),.BLN(BLN38),.WL(WL85));
sram_cell_6t_5 inst_cell_85_39 (.BL(BL39),.BLN(BLN39),.WL(WL85));
sram_cell_6t_5 inst_cell_85_40 (.BL(BL40),.BLN(BLN40),.WL(WL85));
sram_cell_6t_5 inst_cell_85_41 (.BL(BL41),.BLN(BLN41),.WL(WL85));
sram_cell_6t_5 inst_cell_85_42 (.BL(BL42),.BLN(BLN42),.WL(WL85));
sram_cell_6t_5 inst_cell_85_43 (.BL(BL43),.BLN(BLN43),.WL(WL85));
sram_cell_6t_5 inst_cell_85_44 (.BL(BL44),.BLN(BLN44),.WL(WL85));
sram_cell_6t_5 inst_cell_85_45 (.BL(BL45),.BLN(BLN45),.WL(WL85));
sram_cell_6t_5 inst_cell_85_46 (.BL(BL46),.BLN(BLN46),.WL(WL85));
sram_cell_6t_5 inst_cell_85_47 (.BL(BL47),.BLN(BLN47),.WL(WL85));
sram_cell_6t_5 inst_cell_85_48 (.BL(BL48),.BLN(BLN48),.WL(WL85));
sram_cell_6t_5 inst_cell_85_49 (.BL(BL49),.BLN(BLN49),.WL(WL85));
sram_cell_6t_5 inst_cell_85_50 (.BL(BL50),.BLN(BLN50),.WL(WL85));
sram_cell_6t_5 inst_cell_85_51 (.BL(BL51),.BLN(BLN51),.WL(WL85));
sram_cell_6t_5 inst_cell_85_52 (.BL(BL52),.BLN(BLN52),.WL(WL85));
sram_cell_6t_5 inst_cell_85_53 (.BL(BL53),.BLN(BLN53),.WL(WL85));
sram_cell_6t_5 inst_cell_85_54 (.BL(BL54),.BLN(BLN54),.WL(WL85));
sram_cell_6t_5 inst_cell_85_55 (.BL(BL55),.BLN(BLN55),.WL(WL85));
sram_cell_6t_5 inst_cell_85_56 (.BL(BL56),.BLN(BLN56),.WL(WL85));
sram_cell_6t_5 inst_cell_85_57 (.BL(BL57),.BLN(BLN57),.WL(WL85));
sram_cell_6t_5 inst_cell_85_58 (.BL(BL58),.BLN(BLN58),.WL(WL85));
sram_cell_6t_5 inst_cell_85_59 (.BL(BL59),.BLN(BLN59),.WL(WL85));
sram_cell_6t_5 inst_cell_85_60 (.BL(BL60),.BLN(BLN60),.WL(WL85));
sram_cell_6t_5 inst_cell_85_61 (.BL(BL61),.BLN(BLN61),.WL(WL85));
sram_cell_6t_5 inst_cell_85_62 (.BL(BL62),.BLN(BLN62),.WL(WL85));
sram_cell_6t_5 inst_cell_85_63 (.BL(BL63),.BLN(BLN63),.WL(WL85));
sram_cell_6t_5 inst_cell_85_64 (.BL(BL64),.BLN(BLN64),.WL(WL85));
sram_cell_6t_5 inst_cell_85_65 (.BL(BL65),.BLN(BLN65),.WL(WL85));
sram_cell_6t_5 inst_cell_85_66 (.BL(BL66),.BLN(BLN66),.WL(WL85));
sram_cell_6t_5 inst_cell_85_67 (.BL(BL67),.BLN(BLN67),.WL(WL85));
sram_cell_6t_5 inst_cell_85_68 (.BL(BL68),.BLN(BLN68),.WL(WL85));
sram_cell_6t_5 inst_cell_85_69 (.BL(BL69),.BLN(BLN69),.WL(WL85));
sram_cell_6t_5 inst_cell_85_70 (.BL(BL70),.BLN(BLN70),.WL(WL85));
sram_cell_6t_5 inst_cell_85_71 (.BL(BL71),.BLN(BLN71),.WL(WL85));
sram_cell_6t_5 inst_cell_85_72 (.BL(BL72),.BLN(BLN72),.WL(WL85));
sram_cell_6t_5 inst_cell_85_73 (.BL(BL73),.BLN(BLN73),.WL(WL85));
sram_cell_6t_5 inst_cell_85_74 (.BL(BL74),.BLN(BLN74),.WL(WL85));
sram_cell_6t_5 inst_cell_85_75 (.BL(BL75),.BLN(BLN75),.WL(WL85));
sram_cell_6t_5 inst_cell_85_76 (.BL(BL76),.BLN(BLN76),.WL(WL85));
sram_cell_6t_5 inst_cell_85_77 (.BL(BL77),.BLN(BLN77),.WL(WL85));
sram_cell_6t_5 inst_cell_85_78 (.BL(BL78),.BLN(BLN78),.WL(WL85));
sram_cell_6t_5 inst_cell_85_79 (.BL(BL79),.BLN(BLN79),.WL(WL85));
sram_cell_6t_5 inst_cell_85_80 (.BL(BL80),.BLN(BLN80),.WL(WL85));
sram_cell_6t_5 inst_cell_85_81 (.BL(BL81),.BLN(BLN81),.WL(WL85));
sram_cell_6t_5 inst_cell_85_82 (.BL(BL82),.BLN(BLN82),.WL(WL85));
sram_cell_6t_5 inst_cell_85_83 (.BL(BL83),.BLN(BLN83),.WL(WL85));
sram_cell_6t_5 inst_cell_85_84 (.BL(BL84),.BLN(BLN84),.WL(WL85));
sram_cell_6t_5 inst_cell_85_85 (.BL(BL85),.BLN(BLN85),.WL(WL85));
sram_cell_6t_5 inst_cell_85_86 (.BL(BL86),.BLN(BLN86),.WL(WL85));
sram_cell_6t_5 inst_cell_85_87 (.BL(BL87),.BLN(BLN87),.WL(WL85));
sram_cell_6t_5 inst_cell_85_88 (.BL(BL88),.BLN(BLN88),.WL(WL85));
sram_cell_6t_5 inst_cell_85_89 (.BL(BL89),.BLN(BLN89),.WL(WL85));
sram_cell_6t_5 inst_cell_85_90 (.BL(BL90),.BLN(BLN90),.WL(WL85));
sram_cell_6t_5 inst_cell_85_91 (.BL(BL91),.BLN(BLN91),.WL(WL85));
sram_cell_6t_5 inst_cell_85_92 (.BL(BL92),.BLN(BLN92),.WL(WL85));
sram_cell_6t_5 inst_cell_85_93 (.BL(BL93),.BLN(BLN93),.WL(WL85));
sram_cell_6t_5 inst_cell_85_94 (.BL(BL94),.BLN(BLN94),.WL(WL85));
sram_cell_6t_5 inst_cell_85_95 (.BL(BL95),.BLN(BLN95),.WL(WL85));
sram_cell_6t_5 inst_cell_85_96 (.BL(BL96),.BLN(BLN96),.WL(WL85));
sram_cell_6t_5 inst_cell_85_97 (.BL(BL97),.BLN(BLN97),.WL(WL85));
sram_cell_6t_5 inst_cell_85_98 (.BL(BL98),.BLN(BLN98),.WL(WL85));
sram_cell_6t_5 inst_cell_85_99 (.BL(BL99),.BLN(BLN99),.WL(WL85));
sram_cell_6t_5 inst_cell_85_100 (.BL(BL100),.BLN(BLN100),.WL(WL85));
sram_cell_6t_5 inst_cell_85_101 (.BL(BL101),.BLN(BLN101),.WL(WL85));
sram_cell_6t_5 inst_cell_85_102 (.BL(BL102),.BLN(BLN102),.WL(WL85));
sram_cell_6t_5 inst_cell_85_103 (.BL(BL103),.BLN(BLN103),.WL(WL85));
sram_cell_6t_5 inst_cell_85_104 (.BL(BL104),.BLN(BLN104),.WL(WL85));
sram_cell_6t_5 inst_cell_85_105 (.BL(BL105),.BLN(BLN105),.WL(WL85));
sram_cell_6t_5 inst_cell_85_106 (.BL(BL106),.BLN(BLN106),.WL(WL85));
sram_cell_6t_5 inst_cell_85_107 (.BL(BL107),.BLN(BLN107),.WL(WL85));
sram_cell_6t_5 inst_cell_85_108 (.BL(BL108),.BLN(BLN108),.WL(WL85));
sram_cell_6t_5 inst_cell_85_109 (.BL(BL109),.BLN(BLN109),.WL(WL85));
sram_cell_6t_5 inst_cell_85_110 (.BL(BL110),.BLN(BLN110),.WL(WL85));
sram_cell_6t_5 inst_cell_85_111 (.BL(BL111),.BLN(BLN111),.WL(WL85));
sram_cell_6t_5 inst_cell_85_112 (.BL(BL112),.BLN(BLN112),.WL(WL85));
sram_cell_6t_5 inst_cell_85_113 (.BL(BL113),.BLN(BLN113),.WL(WL85));
sram_cell_6t_5 inst_cell_85_114 (.BL(BL114),.BLN(BLN114),.WL(WL85));
sram_cell_6t_5 inst_cell_85_115 (.BL(BL115),.BLN(BLN115),.WL(WL85));
sram_cell_6t_5 inst_cell_85_116 (.BL(BL116),.BLN(BLN116),.WL(WL85));
sram_cell_6t_5 inst_cell_85_117 (.BL(BL117),.BLN(BLN117),.WL(WL85));
sram_cell_6t_5 inst_cell_85_118 (.BL(BL118),.BLN(BLN118),.WL(WL85));
sram_cell_6t_5 inst_cell_85_119 (.BL(BL119),.BLN(BLN119),.WL(WL85));
sram_cell_6t_5 inst_cell_85_120 (.BL(BL120),.BLN(BLN120),.WL(WL85));
sram_cell_6t_5 inst_cell_85_121 (.BL(BL121),.BLN(BLN121),.WL(WL85));
sram_cell_6t_5 inst_cell_85_122 (.BL(BL122),.BLN(BLN122),.WL(WL85));
sram_cell_6t_5 inst_cell_85_123 (.BL(BL123),.BLN(BLN123),.WL(WL85));
sram_cell_6t_5 inst_cell_85_124 (.BL(BL124),.BLN(BLN124),.WL(WL85));
sram_cell_6t_5 inst_cell_85_125 (.BL(BL125),.BLN(BLN125),.WL(WL85));
sram_cell_6t_5 inst_cell_85_126 (.BL(BL126),.BLN(BLN126),.WL(WL85));
sram_cell_6t_5 inst_cell_85_127 (.BL(BL127),.BLN(BLN127),.WL(WL85));
sram_cell_6t_5 inst_cell_86_0 (.BL(BL0),.BLN(BLN0),.WL(WL86));
sram_cell_6t_5 inst_cell_86_1 (.BL(BL1),.BLN(BLN1),.WL(WL86));
sram_cell_6t_5 inst_cell_86_2 (.BL(BL2),.BLN(BLN2),.WL(WL86));
sram_cell_6t_5 inst_cell_86_3 (.BL(BL3),.BLN(BLN3),.WL(WL86));
sram_cell_6t_5 inst_cell_86_4 (.BL(BL4),.BLN(BLN4),.WL(WL86));
sram_cell_6t_5 inst_cell_86_5 (.BL(BL5),.BLN(BLN5),.WL(WL86));
sram_cell_6t_5 inst_cell_86_6 (.BL(BL6),.BLN(BLN6),.WL(WL86));
sram_cell_6t_5 inst_cell_86_7 (.BL(BL7),.BLN(BLN7),.WL(WL86));
sram_cell_6t_5 inst_cell_86_8 (.BL(BL8),.BLN(BLN8),.WL(WL86));
sram_cell_6t_5 inst_cell_86_9 (.BL(BL9),.BLN(BLN9),.WL(WL86));
sram_cell_6t_5 inst_cell_86_10 (.BL(BL10),.BLN(BLN10),.WL(WL86));
sram_cell_6t_5 inst_cell_86_11 (.BL(BL11),.BLN(BLN11),.WL(WL86));
sram_cell_6t_5 inst_cell_86_12 (.BL(BL12),.BLN(BLN12),.WL(WL86));
sram_cell_6t_5 inst_cell_86_13 (.BL(BL13),.BLN(BLN13),.WL(WL86));
sram_cell_6t_5 inst_cell_86_14 (.BL(BL14),.BLN(BLN14),.WL(WL86));
sram_cell_6t_5 inst_cell_86_15 (.BL(BL15),.BLN(BLN15),.WL(WL86));
sram_cell_6t_5 inst_cell_86_16 (.BL(BL16),.BLN(BLN16),.WL(WL86));
sram_cell_6t_5 inst_cell_86_17 (.BL(BL17),.BLN(BLN17),.WL(WL86));
sram_cell_6t_5 inst_cell_86_18 (.BL(BL18),.BLN(BLN18),.WL(WL86));
sram_cell_6t_5 inst_cell_86_19 (.BL(BL19),.BLN(BLN19),.WL(WL86));
sram_cell_6t_5 inst_cell_86_20 (.BL(BL20),.BLN(BLN20),.WL(WL86));
sram_cell_6t_5 inst_cell_86_21 (.BL(BL21),.BLN(BLN21),.WL(WL86));
sram_cell_6t_5 inst_cell_86_22 (.BL(BL22),.BLN(BLN22),.WL(WL86));
sram_cell_6t_5 inst_cell_86_23 (.BL(BL23),.BLN(BLN23),.WL(WL86));
sram_cell_6t_5 inst_cell_86_24 (.BL(BL24),.BLN(BLN24),.WL(WL86));
sram_cell_6t_5 inst_cell_86_25 (.BL(BL25),.BLN(BLN25),.WL(WL86));
sram_cell_6t_5 inst_cell_86_26 (.BL(BL26),.BLN(BLN26),.WL(WL86));
sram_cell_6t_5 inst_cell_86_27 (.BL(BL27),.BLN(BLN27),.WL(WL86));
sram_cell_6t_5 inst_cell_86_28 (.BL(BL28),.BLN(BLN28),.WL(WL86));
sram_cell_6t_5 inst_cell_86_29 (.BL(BL29),.BLN(BLN29),.WL(WL86));
sram_cell_6t_5 inst_cell_86_30 (.BL(BL30),.BLN(BLN30),.WL(WL86));
sram_cell_6t_5 inst_cell_86_31 (.BL(BL31),.BLN(BLN31),.WL(WL86));
sram_cell_6t_5 inst_cell_86_32 (.BL(BL32),.BLN(BLN32),.WL(WL86));
sram_cell_6t_5 inst_cell_86_33 (.BL(BL33),.BLN(BLN33),.WL(WL86));
sram_cell_6t_5 inst_cell_86_34 (.BL(BL34),.BLN(BLN34),.WL(WL86));
sram_cell_6t_5 inst_cell_86_35 (.BL(BL35),.BLN(BLN35),.WL(WL86));
sram_cell_6t_5 inst_cell_86_36 (.BL(BL36),.BLN(BLN36),.WL(WL86));
sram_cell_6t_5 inst_cell_86_37 (.BL(BL37),.BLN(BLN37),.WL(WL86));
sram_cell_6t_5 inst_cell_86_38 (.BL(BL38),.BLN(BLN38),.WL(WL86));
sram_cell_6t_5 inst_cell_86_39 (.BL(BL39),.BLN(BLN39),.WL(WL86));
sram_cell_6t_5 inst_cell_86_40 (.BL(BL40),.BLN(BLN40),.WL(WL86));
sram_cell_6t_5 inst_cell_86_41 (.BL(BL41),.BLN(BLN41),.WL(WL86));
sram_cell_6t_5 inst_cell_86_42 (.BL(BL42),.BLN(BLN42),.WL(WL86));
sram_cell_6t_5 inst_cell_86_43 (.BL(BL43),.BLN(BLN43),.WL(WL86));
sram_cell_6t_5 inst_cell_86_44 (.BL(BL44),.BLN(BLN44),.WL(WL86));
sram_cell_6t_5 inst_cell_86_45 (.BL(BL45),.BLN(BLN45),.WL(WL86));
sram_cell_6t_5 inst_cell_86_46 (.BL(BL46),.BLN(BLN46),.WL(WL86));
sram_cell_6t_5 inst_cell_86_47 (.BL(BL47),.BLN(BLN47),.WL(WL86));
sram_cell_6t_5 inst_cell_86_48 (.BL(BL48),.BLN(BLN48),.WL(WL86));
sram_cell_6t_5 inst_cell_86_49 (.BL(BL49),.BLN(BLN49),.WL(WL86));
sram_cell_6t_5 inst_cell_86_50 (.BL(BL50),.BLN(BLN50),.WL(WL86));
sram_cell_6t_5 inst_cell_86_51 (.BL(BL51),.BLN(BLN51),.WL(WL86));
sram_cell_6t_5 inst_cell_86_52 (.BL(BL52),.BLN(BLN52),.WL(WL86));
sram_cell_6t_5 inst_cell_86_53 (.BL(BL53),.BLN(BLN53),.WL(WL86));
sram_cell_6t_5 inst_cell_86_54 (.BL(BL54),.BLN(BLN54),.WL(WL86));
sram_cell_6t_5 inst_cell_86_55 (.BL(BL55),.BLN(BLN55),.WL(WL86));
sram_cell_6t_5 inst_cell_86_56 (.BL(BL56),.BLN(BLN56),.WL(WL86));
sram_cell_6t_5 inst_cell_86_57 (.BL(BL57),.BLN(BLN57),.WL(WL86));
sram_cell_6t_5 inst_cell_86_58 (.BL(BL58),.BLN(BLN58),.WL(WL86));
sram_cell_6t_5 inst_cell_86_59 (.BL(BL59),.BLN(BLN59),.WL(WL86));
sram_cell_6t_5 inst_cell_86_60 (.BL(BL60),.BLN(BLN60),.WL(WL86));
sram_cell_6t_5 inst_cell_86_61 (.BL(BL61),.BLN(BLN61),.WL(WL86));
sram_cell_6t_5 inst_cell_86_62 (.BL(BL62),.BLN(BLN62),.WL(WL86));
sram_cell_6t_5 inst_cell_86_63 (.BL(BL63),.BLN(BLN63),.WL(WL86));
sram_cell_6t_5 inst_cell_86_64 (.BL(BL64),.BLN(BLN64),.WL(WL86));
sram_cell_6t_5 inst_cell_86_65 (.BL(BL65),.BLN(BLN65),.WL(WL86));
sram_cell_6t_5 inst_cell_86_66 (.BL(BL66),.BLN(BLN66),.WL(WL86));
sram_cell_6t_5 inst_cell_86_67 (.BL(BL67),.BLN(BLN67),.WL(WL86));
sram_cell_6t_5 inst_cell_86_68 (.BL(BL68),.BLN(BLN68),.WL(WL86));
sram_cell_6t_5 inst_cell_86_69 (.BL(BL69),.BLN(BLN69),.WL(WL86));
sram_cell_6t_5 inst_cell_86_70 (.BL(BL70),.BLN(BLN70),.WL(WL86));
sram_cell_6t_5 inst_cell_86_71 (.BL(BL71),.BLN(BLN71),.WL(WL86));
sram_cell_6t_5 inst_cell_86_72 (.BL(BL72),.BLN(BLN72),.WL(WL86));
sram_cell_6t_5 inst_cell_86_73 (.BL(BL73),.BLN(BLN73),.WL(WL86));
sram_cell_6t_5 inst_cell_86_74 (.BL(BL74),.BLN(BLN74),.WL(WL86));
sram_cell_6t_5 inst_cell_86_75 (.BL(BL75),.BLN(BLN75),.WL(WL86));
sram_cell_6t_5 inst_cell_86_76 (.BL(BL76),.BLN(BLN76),.WL(WL86));
sram_cell_6t_5 inst_cell_86_77 (.BL(BL77),.BLN(BLN77),.WL(WL86));
sram_cell_6t_5 inst_cell_86_78 (.BL(BL78),.BLN(BLN78),.WL(WL86));
sram_cell_6t_5 inst_cell_86_79 (.BL(BL79),.BLN(BLN79),.WL(WL86));
sram_cell_6t_5 inst_cell_86_80 (.BL(BL80),.BLN(BLN80),.WL(WL86));
sram_cell_6t_5 inst_cell_86_81 (.BL(BL81),.BLN(BLN81),.WL(WL86));
sram_cell_6t_5 inst_cell_86_82 (.BL(BL82),.BLN(BLN82),.WL(WL86));
sram_cell_6t_5 inst_cell_86_83 (.BL(BL83),.BLN(BLN83),.WL(WL86));
sram_cell_6t_5 inst_cell_86_84 (.BL(BL84),.BLN(BLN84),.WL(WL86));
sram_cell_6t_5 inst_cell_86_85 (.BL(BL85),.BLN(BLN85),.WL(WL86));
sram_cell_6t_5 inst_cell_86_86 (.BL(BL86),.BLN(BLN86),.WL(WL86));
sram_cell_6t_5 inst_cell_86_87 (.BL(BL87),.BLN(BLN87),.WL(WL86));
sram_cell_6t_5 inst_cell_86_88 (.BL(BL88),.BLN(BLN88),.WL(WL86));
sram_cell_6t_5 inst_cell_86_89 (.BL(BL89),.BLN(BLN89),.WL(WL86));
sram_cell_6t_5 inst_cell_86_90 (.BL(BL90),.BLN(BLN90),.WL(WL86));
sram_cell_6t_5 inst_cell_86_91 (.BL(BL91),.BLN(BLN91),.WL(WL86));
sram_cell_6t_5 inst_cell_86_92 (.BL(BL92),.BLN(BLN92),.WL(WL86));
sram_cell_6t_5 inst_cell_86_93 (.BL(BL93),.BLN(BLN93),.WL(WL86));
sram_cell_6t_5 inst_cell_86_94 (.BL(BL94),.BLN(BLN94),.WL(WL86));
sram_cell_6t_5 inst_cell_86_95 (.BL(BL95),.BLN(BLN95),.WL(WL86));
sram_cell_6t_5 inst_cell_86_96 (.BL(BL96),.BLN(BLN96),.WL(WL86));
sram_cell_6t_5 inst_cell_86_97 (.BL(BL97),.BLN(BLN97),.WL(WL86));
sram_cell_6t_5 inst_cell_86_98 (.BL(BL98),.BLN(BLN98),.WL(WL86));
sram_cell_6t_5 inst_cell_86_99 (.BL(BL99),.BLN(BLN99),.WL(WL86));
sram_cell_6t_5 inst_cell_86_100 (.BL(BL100),.BLN(BLN100),.WL(WL86));
sram_cell_6t_5 inst_cell_86_101 (.BL(BL101),.BLN(BLN101),.WL(WL86));
sram_cell_6t_5 inst_cell_86_102 (.BL(BL102),.BLN(BLN102),.WL(WL86));
sram_cell_6t_5 inst_cell_86_103 (.BL(BL103),.BLN(BLN103),.WL(WL86));
sram_cell_6t_5 inst_cell_86_104 (.BL(BL104),.BLN(BLN104),.WL(WL86));
sram_cell_6t_5 inst_cell_86_105 (.BL(BL105),.BLN(BLN105),.WL(WL86));
sram_cell_6t_5 inst_cell_86_106 (.BL(BL106),.BLN(BLN106),.WL(WL86));
sram_cell_6t_5 inst_cell_86_107 (.BL(BL107),.BLN(BLN107),.WL(WL86));
sram_cell_6t_5 inst_cell_86_108 (.BL(BL108),.BLN(BLN108),.WL(WL86));
sram_cell_6t_5 inst_cell_86_109 (.BL(BL109),.BLN(BLN109),.WL(WL86));
sram_cell_6t_5 inst_cell_86_110 (.BL(BL110),.BLN(BLN110),.WL(WL86));
sram_cell_6t_5 inst_cell_86_111 (.BL(BL111),.BLN(BLN111),.WL(WL86));
sram_cell_6t_5 inst_cell_86_112 (.BL(BL112),.BLN(BLN112),.WL(WL86));
sram_cell_6t_5 inst_cell_86_113 (.BL(BL113),.BLN(BLN113),.WL(WL86));
sram_cell_6t_5 inst_cell_86_114 (.BL(BL114),.BLN(BLN114),.WL(WL86));
sram_cell_6t_5 inst_cell_86_115 (.BL(BL115),.BLN(BLN115),.WL(WL86));
sram_cell_6t_5 inst_cell_86_116 (.BL(BL116),.BLN(BLN116),.WL(WL86));
sram_cell_6t_5 inst_cell_86_117 (.BL(BL117),.BLN(BLN117),.WL(WL86));
sram_cell_6t_5 inst_cell_86_118 (.BL(BL118),.BLN(BLN118),.WL(WL86));
sram_cell_6t_5 inst_cell_86_119 (.BL(BL119),.BLN(BLN119),.WL(WL86));
sram_cell_6t_5 inst_cell_86_120 (.BL(BL120),.BLN(BLN120),.WL(WL86));
sram_cell_6t_5 inst_cell_86_121 (.BL(BL121),.BLN(BLN121),.WL(WL86));
sram_cell_6t_5 inst_cell_86_122 (.BL(BL122),.BLN(BLN122),.WL(WL86));
sram_cell_6t_5 inst_cell_86_123 (.BL(BL123),.BLN(BLN123),.WL(WL86));
sram_cell_6t_5 inst_cell_86_124 (.BL(BL124),.BLN(BLN124),.WL(WL86));
sram_cell_6t_5 inst_cell_86_125 (.BL(BL125),.BLN(BLN125),.WL(WL86));
sram_cell_6t_5 inst_cell_86_126 (.BL(BL126),.BLN(BLN126),.WL(WL86));
sram_cell_6t_5 inst_cell_86_127 (.BL(BL127),.BLN(BLN127),.WL(WL86));
sram_cell_6t_5 inst_cell_87_0 (.BL(BL0),.BLN(BLN0),.WL(WL87));
sram_cell_6t_5 inst_cell_87_1 (.BL(BL1),.BLN(BLN1),.WL(WL87));
sram_cell_6t_5 inst_cell_87_2 (.BL(BL2),.BLN(BLN2),.WL(WL87));
sram_cell_6t_5 inst_cell_87_3 (.BL(BL3),.BLN(BLN3),.WL(WL87));
sram_cell_6t_5 inst_cell_87_4 (.BL(BL4),.BLN(BLN4),.WL(WL87));
sram_cell_6t_5 inst_cell_87_5 (.BL(BL5),.BLN(BLN5),.WL(WL87));
sram_cell_6t_5 inst_cell_87_6 (.BL(BL6),.BLN(BLN6),.WL(WL87));
sram_cell_6t_5 inst_cell_87_7 (.BL(BL7),.BLN(BLN7),.WL(WL87));
sram_cell_6t_5 inst_cell_87_8 (.BL(BL8),.BLN(BLN8),.WL(WL87));
sram_cell_6t_5 inst_cell_87_9 (.BL(BL9),.BLN(BLN9),.WL(WL87));
sram_cell_6t_5 inst_cell_87_10 (.BL(BL10),.BLN(BLN10),.WL(WL87));
sram_cell_6t_5 inst_cell_87_11 (.BL(BL11),.BLN(BLN11),.WL(WL87));
sram_cell_6t_5 inst_cell_87_12 (.BL(BL12),.BLN(BLN12),.WL(WL87));
sram_cell_6t_5 inst_cell_87_13 (.BL(BL13),.BLN(BLN13),.WL(WL87));
sram_cell_6t_5 inst_cell_87_14 (.BL(BL14),.BLN(BLN14),.WL(WL87));
sram_cell_6t_5 inst_cell_87_15 (.BL(BL15),.BLN(BLN15),.WL(WL87));
sram_cell_6t_5 inst_cell_87_16 (.BL(BL16),.BLN(BLN16),.WL(WL87));
sram_cell_6t_5 inst_cell_87_17 (.BL(BL17),.BLN(BLN17),.WL(WL87));
sram_cell_6t_5 inst_cell_87_18 (.BL(BL18),.BLN(BLN18),.WL(WL87));
sram_cell_6t_5 inst_cell_87_19 (.BL(BL19),.BLN(BLN19),.WL(WL87));
sram_cell_6t_5 inst_cell_87_20 (.BL(BL20),.BLN(BLN20),.WL(WL87));
sram_cell_6t_5 inst_cell_87_21 (.BL(BL21),.BLN(BLN21),.WL(WL87));
sram_cell_6t_5 inst_cell_87_22 (.BL(BL22),.BLN(BLN22),.WL(WL87));
sram_cell_6t_5 inst_cell_87_23 (.BL(BL23),.BLN(BLN23),.WL(WL87));
sram_cell_6t_5 inst_cell_87_24 (.BL(BL24),.BLN(BLN24),.WL(WL87));
sram_cell_6t_5 inst_cell_87_25 (.BL(BL25),.BLN(BLN25),.WL(WL87));
sram_cell_6t_5 inst_cell_87_26 (.BL(BL26),.BLN(BLN26),.WL(WL87));
sram_cell_6t_5 inst_cell_87_27 (.BL(BL27),.BLN(BLN27),.WL(WL87));
sram_cell_6t_5 inst_cell_87_28 (.BL(BL28),.BLN(BLN28),.WL(WL87));
sram_cell_6t_5 inst_cell_87_29 (.BL(BL29),.BLN(BLN29),.WL(WL87));
sram_cell_6t_5 inst_cell_87_30 (.BL(BL30),.BLN(BLN30),.WL(WL87));
sram_cell_6t_5 inst_cell_87_31 (.BL(BL31),.BLN(BLN31),.WL(WL87));
sram_cell_6t_5 inst_cell_87_32 (.BL(BL32),.BLN(BLN32),.WL(WL87));
sram_cell_6t_5 inst_cell_87_33 (.BL(BL33),.BLN(BLN33),.WL(WL87));
sram_cell_6t_5 inst_cell_87_34 (.BL(BL34),.BLN(BLN34),.WL(WL87));
sram_cell_6t_5 inst_cell_87_35 (.BL(BL35),.BLN(BLN35),.WL(WL87));
sram_cell_6t_5 inst_cell_87_36 (.BL(BL36),.BLN(BLN36),.WL(WL87));
sram_cell_6t_5 inst_cell_87_37 (.BL(BL37),.BLN(BLN37),.WL(WL87));
sram_cell_6t_5 inst_cell_87_38 (.BL(BL38),.BLN(BLN38),.WL(WL87));
sram_cell_6t_5 inst_cell_87_39 (.BL(BL39),.BLN(BLN39),.WL(WL87));
sram_cell_6t_5 inst_cell_87_40 (.BL(BL40),.BLN(BLN40),.WL(WL87));
sram_cell_6t_5 inst_cell_87_41 (.BL(BL41),.BLN(BLN41),.WL(WL87));
sram_cell_6t_5 inst_cell_87_42 (.BL(BL42),.BLN(BLN42),.WL(WL87));
sram_cell_6t_5 inst_cell_87_43 (.BL(BL43),.BLN(BLN43),.WL(WL87));
sram_cell_6t_5 inst_cell_87_44 (.BL(BL44),.BLN(BLN44),.WL(WL87));
sram_cell_6t_5 inst_cell_87_45 (.BL(BL45),.BLN(BLN45),.WL(WL87));
sram_cell_6t_5 inst_cell_87_46 (.BL(BL46),.BLN(BLN46),.WL(WL87));
sram_cell_6t_5 inst_cell_87_47 (.BL(BL47),.BLN(BLN47),.WL(WL87));
sram_cell_6t_5 inst_cell_87_48 (.BL(BL48),.BLN(BLN48),.WL(WL87));
sram_cell_6t_5 inst_cell_87_49 (.BL(BL49),.BLN(BLN49),.WL(WL87));
sram_cell_6t_5 inst_cell_87_50 (.BL(BL50),.BLN(BLN50),.WL(WL87));
sram_cell_6t_5 inst_cell_87_51 (.BL(BL51),.BLN(BLN51),.WL(WL87));
sram_cell_6t_5 inst_cell_87_52 (.BL(BL52),.BLN(BLN52),.WL(WL87));
sram_cell_6t_5 inst_cell_87_53 (.BL(BL53),.BLN(BLN53),.WL(WL87));
sram_cell_6t_5 inst_cell_87_54 (.BL(BL54),.BLN(BLN54),.WL(WL87));
sram_cell_6t_5 inst_cell_87_55 (.BL(BL55),.BLN(BLN55),.WL(WL87));
sram_cell_6t_5 inst_cell_87_56 (.BL(BL56),.BLN(BLN56),.WL(WL87));
sram_cell_6t_5 inst_cell_87_57 (.BL(BL57),.BLN(BLN57),.WL(WL87));
sram_cell_6t_5 inst_cell_87_58 (.BL(BL58),.BLN(BLN58),.WL(WL87));
sram_cell_6t_5 inst_cell_87_59 (.BL(BL59),.BLN(BLN59),.WL(WL87));
sram_cell_6t_5 inst_cell_87_60 (.BL(BL60),.BLN(BLN60),.WL(WL87));
sram_cell_6t_5 inst_cell_87_61 (.BL(BL61),.BLN(BLN61),.WL(WL87));
sram_cell_6t_5 inst_cell_87_62 (.BL(BL62),.BLN(BLN62),.WL(WL87));
sram_cell_6t_5 inst_cell_87_63 (.BL(BL63),.BLN(BLN63),.WL(WL87));
sram_cell_6t_5 inst_cell_87_64 (.BL(BL64),.BLN(BLN64),.WL(WL87));
sram_cell_6t_5 inst_cell_87_65 (.BL(BL65),.BLN(BLN65),.WL(WL87));
sram_cell_6t_5 inst_cell_87_66 (.BL(BL66),.BLN(BLN66),.WL(WL87));
sram_cell_6t_5 inst_cell_87_67 (.BL(BL67),.BLN(BLN67),.WL(WL87));
sram_cell_6t_5 inst_cell_87_68 (.BL(BL68),.BLN(BLN68),.WL(WL87));
sram_cell_6t_5 inst_cell_87_69 (.BL(BL69),.BLN(BLN69),.WL(WL87));
sram_cell_6t_5 inst_cell_87_70 (.BL(BL70),.BLN(BLN70),.WL(WL87));
sram_cell_6t_5 inst_cell_87_71 (.BL(BL71),.BLN(BLN71),.WL(WL87));
sram_cell_6t_5 inst_cell_87_72 (.BL(BL72),.BLN(BLN72),.WL(WL87));
sram_cell_6t_5 inst_cell_87_73 (.BL(BL73),.BLN(BLN73),.WL(WL87));
sram_cell_6t_5 inst_cell_87_74 (.BL(BL74),.BLN(BLN74),.WL(WL87));
sram_cell_6t_5 inst_cell_87_75 (.BL(BL75),.BLN(BLN75),.WL(WL87));
sram_cell_6t_5 inst_cell_87_76 (.BL(BL76),.BLN(BLN76),.WL(WL87));
sram_cell_6t_5 inst_cell_87_77 (.BL(BL77),.BLN(BLN77),.WL(WL87));
sram_cell_6t_5 inst_cell_87_78 (.BL(BL78),.BLN(BLN78),.WL(WL87));
sram_cell_6t_5 inst_cell_87_79 (.BL(BL79),.BLN(BLN79),.WL(WL87));
sram_cell_6t_5 inst_cell_87_80 (.BL(BL80),.BLN(BLN80),.WL(WL87));
sram_cell_6t_5 inst_cell_87_81 (.BL(BL81),.BLN(BLN81),.WL(WL87));
sram_cell_6t_5 inst_cell_87_82 (.BL(BL82),.BLN(BLN82),.WL(WL87));
sram_cell_6t_5 inst_cell_87_83 (.BL(BL83),.BLN(BLN83),.WL(WL87));
sram_cell_6t_5 inst_cell_87_84 (.BL(BL84),.BLN(BLN84),.WL(WL87));
sram_cell_6t_5 inst_cell_87_85 (.BL(BL85),.BLN(BLN85),.WL(WL87));
sram_cell_6t_5 inst_cell_87_86 (.BL(BL86),.BLN(BLN86),.WL(WL87));
sram_cell_6t_5 inst_cell_87_87 (.BL(BL87),.BLN(BLN87),.WL(WL87));
sram_cell_6t_5 inst_cell_87_88 (.BL(BL88),.BLN(BLN88),.WL(WL87));
sram_cell_6t_5 inst_cell_87_89 (.BL(BL89),.BLN(BLN89),.WL(WL87));
sram_cell_6t_5 inst_cell_87_90 (.BL(BL90),.BLN(BLN90),.WL(WL87));
sram_cell_6t_5 inst_cell_87_91 (.BL(BL91),.BLN(BLN91),.WL(WL87));
sram_cell_6t_5 inst_cell_87_92 (.BL(BL92),.BLN(BLN92),.WL(WL87));
sram_cell_6t_5 inst_cell_87_93 (.BL(BL93),.BLN(BLN93),.WL(WL87));
sram_cell_6t_5 inst_cell_87_94 (.BL(BL94),.BLN(BLN94),.WL(WL87));
sram_cell_6t_5 inst_cell_87_95 (.BL(BL95),.BLN(BLN95),.WL(WL87));
sram_cell_6t_5 inst_cell_87_96 (.BL(BL96),.BLN(BLN96),.WL(WL87));
sram_cell_6t_5 inst_cell_87_97 (.BL(BL97),.BLN(BLN97),.WL(WL87));
sram_cell_6t_5 inst_cell_87_98 (.BL(BL98),.BLN(BLN98),.WL(WL87));
sram_cell_6t_5 inst_cell_87_99 (.BL(BL99),.BLN(BLN99),.WL(WL87));
sram_cell_6t_5 inst_cell_87_100 (.BL(BL100),.BLN(BLN100),.WL(WL87));
sram_cell_6t_5 inst_cell_87_101 (.BL(BL101),.BLN(BLN101),.WL(WL87));
sram_cell_6t_5 inst_cell_87_102 (.BL(BL102),.BLN(BLN102),.WL(WL87));
sram_cell_6t_5 inst_cell_87_103 (.BL(BL103),.BLN(BLN103),.WL(WL87));
sram_cell_6t_5 inst_cell_87_104 (.BL(BL104),.BLN(BLN104),.WL(WL87));
sram_cell_6t_5 inst_cell_87_105 (.BL(BL105),.BLN(BLN105),.WL(WL87));
sram_cell_6t_5 inst_cell_87_106 (.BL(BL106),.BLN(BLN106),.WL(WL87));
sram_cell_6t_5 inst_cell_87_107 (.BL(BL107),.BLN(BLN107),.WL(WL87));
sram_cell_6t_5 inst_cell_87_108 (.BL(BL108),.BLN(BLN108),.WL(WL87));
sram_cell_6t_5 inst_cell_87_109 (.BL(BL109),.BLN(BLN109),.WL(WL87));
sram_cell_6t_5 inst_cell_87_110 (.BL(BL110),.BLN(BLN110),.WL(WL87));
sram_cell_6t_5 inst_cell_87_111 (.BL(BL111),.BLN(BLN111),.WL(WL87));
sram_cell_6t_5 inst_cell_87_112 (.BL(BL112),.BLN(BLN112),.WL(WL87));
sram_cell_6t_5 inst_cell_87_113 (.BL(BL113),.BLN(BLN113),.WL(WL87));
sram_cell_6t_5 inst_cell_87_114 (.BL(BL114),.BLN(BLN114),.WL(WL87));
sram_cell_6t_5 inst_cell_87_115 (.BL(BL115),.BLN(BLN115),.WL(WL87));
sram_cell_6t_5 inst_cell_87_116 (.BL(BL116),.BLN(BLN116),.WL(WL87));
sram_cell_6t_5 inst_cell_87_117 (.BL(BL117),.BLN(BLN117),.WL(WL87));
sram_cell_6t_5 inst_cell_87_118 (.BL(BL118),.BLN(BLN118),.WL(WL87));
sram_cell_6t_5 inst_cell_87_119 (.BL(BL119),.BLN(BLN119),.WL(WL87));
sram_cell_6t_5 inst_cell_87_120 (.BL(BL120),.BLN(BLN120),.WL(WL87));
sram_cell_6t_5 inst_cell_87_121 (.BL(BL121),.BLN(BLN121),.WL(WL87));
sram_cell_6t_5 inst_cell_87_122 (.BL(BL122),.BLN(BLN122),.WL(WL87));
sram_cell_6t_5 inst_cell_87_123 (.BL(BL123),.BLN(BLN123),.WL(WL87));
sram_cell_6t_5 inst_cell_87_124 (.BL(BL124),.BLN(BLN124),.WL(WL87));
sram_cell_6t_5 inst_cell_87_125 (.BL(BL125),.BLN(BLN125),.WL(WL87));
sram_cell_6t_5 inst_cell_87_126 (.BL(BL126),.BLN(BLN126),.WL(WL87));
sram_cell_6t_5 inst_cell_87_127 (.BL(BL127),.BLN(BLN127),.WL(WL87));
sram_cell_6t_5 inst_cell_88_0 (.BL(BL0),.BLN(BLN0),.WL(WL88));
sram_cell_6t_5 inst_cell_88_1 (.BL(BL1),.BLN(BLN1),.WL(WL88));
sram_cell_6t_5 inst_cell_88_2 (.BL(BL2),.BLN(BLN2),.WL(WL88));
sram_cell_6t_5 inst_cell_88_3 (.BL(BL3),.BLN(BLN3),.WL(WL88));
sram_cell_6t_5 inst_cell_88_4 (.BL(BL4),.BLN(BLN4),.WL(WL88));
sram_cell_6t_5 inst_cell_88_5 (.BL(BL5),.BLN(BLN5),.WL(WL88));
sram_cell_6t_5 inst_cell_88_6 (.BL(BL6),.BLN(BLN6),.WL(WL88));
sram_cell_6t_5 inst_cell_88_7 (.BL(BL7),.BLN(BLN7),.WL(WL88));
sram_cell_6t_5 inst_cell_88_8 (.BL(BL8),.BLN(BLN8),.WL(WL88));
sram_cell_6t_5 inst_cell_88_9 (.BL(BL9),.BLN(BLN9),.WL(WL88));
sram_cell_6t_5 inst_cell_88_10 (.BL(BL10),.BLN(BLN10),.WL(WL88));
sram_cell_6t_5 inst_cell_88_11 (.BL(BL11),.BLN(BLN11),.WL(WL88));
sram_cell_6t_5 inst_cell_88_12 (.BL(BL12),.BLN(BLN12),.WL(WL88));
sram_cell_6t_5 inst_cell_88_13 (.BL(BL13),.BLN(BLN13),.WL(WL88));
sram_cell_6t_5 inst_cell_88_14 (.BL(BL14),.BLN(BLN14),.WL(WL88));
sram_cell_6t_5 inst_cell_88_15 (.BL(BL15),.BLN(BLN15),.WL(WL88));
sram_cell_6t_5 inst_cell_88_16 (.BL(BL16),.BLN(BLN16),.WL(WL88));
sram_cell_6t_5 inst_cell_88_17 (.BL(BL17),.BLN(BLN17),.WL(WL88));
sram_cell_6t_5 inst_cell_88_18 (.BL(BL18),.BLN(BLN18),.WL(WL88));
sram_cell_6t_5 inst_cell_88_19 (.BL(BL19),.BLN(BLN19),.WL(WL88));
sram_cell_6t_5 inst_cell_88_20 (.BL(BL20),.BLN(BLN20),.WL(WL88));
sram_cell_6t_5 inst_cell_88_21 (.BL(BL21),.BLN(BLN21),.WL(WL88));
sram_cell_6t_5 inst_cell_88_22 (.BL(BL22),.BLN(BLN22),.WL(WL88));
sram_cell_6t_5 inst_cell_88_23 (.BL(BL23),.BLN(BLN23),.WL(WL88));
sram_cell_6t_5 inst_cell_88_24 (.BL(BL24),.BLN(BLN24),.WL(WL88));
sram_cell_6t_5 inst_cell_88_25 (.BL(BL25),.BLN(BLN25),.WL(WL88));
sram_cell_6t_5 inst_cell_88_26 (.BL(BL26),.BLN(BLN26),.WL(WL88));
sram_cell_6t_5 inst_cell_88_27 (.BL(BL27),.BLN(BLN27),.WL(WL88));
sram_cell_6t_5 inst_cell_88_28 (.BL(BL28),.BLN(BLN28),.WL(WL88));
sram_cell_6t_5 inst_cell_88_29 (.BL(BL29),.BLN(BLN29),.WL(WL88));
sram_cell_6t_5 inst_cell_88_30 (.BL(BL30),.BLN(BLN30),.WL(WL88));
sram_cell_6t_5 inst_cell_88_31 (.BL(BL31),.BLN(BLN31),.WL(WL88));
sram_cell_6t_5 inst_cell_88_32 (.BL(BL32),.BLN(BLN32),.WL(WL88));
sram_cell_6t_5 inst_cell_88_33 (.BL(BL33),.BLN(BLN33),.WL(WL88));
sram_cell_6t_5 inst_cell_88_34 (.BL(BL34),.BLN(BLN34),.WL(WL88));
sram_cell_6t_5 inst_cell_88_35 (.BL(BL35),.BLN(BLN35),.WL(WL88));
sram_cell_6t_5 inst_cell_88_36 (.BL(BL36),.BLN(BLN36),.WL(WL88));
sram_cell_6t_5 inst_cell_88_37 (.BL(BL37),.BLN(BLN37),.WL(WL88));
sram_cell_6t_5 inst_cell_88_38 (.BL(BL38),.BLN(BLN38),.WL(WL88));
sram_cell_6t_5 inst_cell_88_39 (.BL(BL39),.BLN(BLN39),.WL(WL88));
sram_cell_6t_5 inst_cell_88_40 (.BL(BL40),.BLN(BLN40),.WL(WL88));
sram_cell_6t_5 inst_cell_88_41 (.BL(BL41),.BLN(BLN41),.WL(WL88));
sram_cell_6t_5 inst_cell_88_42 (.BL(BL42),.BLN(BLN42),.WL(WL88));
sram_cell_6t_5 inst_cell_88_43 (.BL(BL43),.BLN(BLN43),.WL(WL88));
sram_cell_6t_5 inst_cell_88_44 (.BL(BL44),.BLN(BLN44),.WL(WL88));
sram_cell_6t_5 inst_cell_88_45 (.BL(BL45),.BLN(BLN45),.WL(WL88));
sram_cell_6t_5 inst_cell_88_46 (.BL(BL46),.BLN(BLN46),.WL(WL88));
sram_cell_6t_5 inst_cell_88_47 (.BL(BL47),.BLN(BLN47),.WL(WL88));
sram_cell_6t_5 inst_cell_88_48 (.BL(BL48),.BLN(BLN48),.WL(WL88));
sram_cell_6t_5 inst_cell_88_49 (.BL(BL49),.BLN(BLN49),.WL(WL88));
sram_cell_6t_5 inst_cell_88_50 (.BL(BL50),.BLN(BLN50),.WL(WL88));
sram_cell_6t_5 inst_cell_88_51 (.BL(BL51),.BLN(BLN51),.WL(WL88));
sram_cell_6t_5 inst_cell_88_52 (.BL(BL52),.BLN(BLN52),.WL(WL88));
sram_cell_6t_5 inst_cell_88_53 (.BL(BL53),.BLN(BLN53),.WL(WL88));
sram_cell_6t_5 inst_cell_88_54 (.BL(BL54),.BLN(BLN54),.WL(WL88));
sram_cell_6t_5 inst_cell_88_55 (.BL(BL55),.BLN(BLN55),.WL(WL88));
sram_cell_6t_5 inst_cell_88_56 (.BL(BL56),.BLN(BLN56),.WL(WL88));
sram_cell_6t_5 inst_cell_88_57 (.BL(BL57),.BLN(BLN57),.WL(WL88));
sram_cell_6t_5 inst_cell_88_58 (.BL(BL58),.BLN(BLN58),.WL(WL88));
sram_cell_6t_5 inst_cell_88_59 (.BL(BL59),.BLN(BLN59),.WL(WL88));
sram_cell_6t_5 inst_cell_88_60 (.BL(BL60),.BLN(BLN60),.WL(WL88));
sram_cell_6t_5 inst_cell_88_61 (.BL(BL61),.BLN(BLN61),.WL(WL88));
sram_cell_6t_5 inst_cell_88_62 (.BL(BL62),.BLN(BLN62),.WL(WL88));
sram_cell_6t_5 inst_cell_88_63 (.BL(BL63),.BLN(BLN63),.WL(WL88));
sram_cell_6t_5 inst_cell_88_64 (.BL(BL64),.BLN(BLN64),.WL(WL88));
sram_cell_6t_5 inst_cell_88_65 (.BL(BL65),.BLN(BLN65),.WL(WL88));
sram_cell_6t_5 inst_cell_88_66 (.BL(BL66),.BLN(BLN66),.WL(WL88));
sram_cell_6t_5 inst_cell_88_67 (.BL(BL67),.BLN(BLN67),.WL(WL88));
sram_cell_6t_5 inst_cell_88_68 (.BL(BL68),.BLN(BLN68),.WL(WL88));
sram_cell_6t_5 inst_cell_88_69 (.BL(BL69),.BLN(BLN69),.WL(WL88));
sram_cell_6t_5 inst_cell_88_70 (.BL(BL70),.BLN(BLN70),.WL(WL88));
sram_cell_6t_5 inst_cell_88_71 (.BL(BL71),.BLN(BLN71),.WL(WL88));
sram_cell_6t_5 inst_cell_88_72 (.BL(BL72),.BLN(BLN72),.WL(WL88));
sram_cell_6t_5 inst_cell_88_73 (.BL(BL73),.BLN(BLN73),.WL(WL88));
sram_cell_6t_5 inst_cell_88_74 (.BL(BL74),.BLN(BLN74),.WL(WL88));
sram_cell_6t_5 inst_cell_88_75 (.BL(BL75),.BLN(BLN75),.WL(WL88));
sram_cell_6t_5 inst_cell_88_76 (.BL(BL76),.BLN(BLN76),.WL(WL88));
sram_cell_6t_5 inst_cell_88_77 (.BL(BL77),.BLN(BLN77),.WL(WL88));
sram_cell_6t_5 inst_cell_88_78 (.BL(BL78),.BLN(BLN78),.WL(WL88));
sram_cell_6t_5 inst_cell_88_79 (.BL(BL79),.BLN(BLN79),.WL(WL88));
sram_cell_6t_5 inst_cell_88_80 (.BL(BL80),.BLN(BLN80),.WL(WL88));
sram_cell_6t_5 inst_cell_88_81 (.BL(BL81),.BLN(BLN81),.WL(WL88));
sram_cell_6t_5 inst_cell_88_82 (.BL(BL82),.BLN(BLN82),.WL(WL88));
sram_cell_6t_5 inst_cell_88_83 (.BL(BL83),.BLN(BLN83),.WL(WL88));
sram_cell_6t_5 inst_cell_88_84 (.BL(BL84),.BLN(BLN84),.WL(WL88));
sram_cell_6t_5 inst_cell_88_85 (.BL(BL85),.BLN(BLN85),.WL(WL88));
sram_cell_6t_5 inst_cell_88_86 (.BL(BL86),.BLN(BLN86),.WL(WL88));
sram_cell_6t_5 inst_cell_88_87 (.BL(BL87),.BLN(BLN87),.WL(WL88));
sram_cell_6t_5 inst_cell_88_88 (.BL(BL88),.BLN(BLN88),.WL(WL88));
sram_cell_6t_5 inst_cell_88_89 (.BL(BL89),.BLN(BLN89),.WL(WL88));
sram_cell_6t_5 inst_cell_88_90 (.BL(BL90),.BLN(BLN90),.WL(WL88));
sram_cell_6t_5 inst_cell_88_91 (.BL(BL91),.BLN(BLN91),.WL(WL88));
sram_cell_6t_5 inst_cell_88_92 (.BL(BL92),.BLN(BLN92),.WL(WL88));
sram_cell_6t_5 inst_cell_88_93 (.BL(BL93),.BLN(BLN93),.WL(WL88));
sram_cell_6t_5 inst_cell_88_94 (.BL(BL94),.BLN(BLN94),.WL(WL88));
sram_cell_6t_5 inst_cell_88_95 (.BL(BL95),.BLN(BLN95),.WL(WL88));
sram_cell_6t_5 inst_cell_88_96 (.BL(BL96),.BLN(BLN96),.WL(WL88));
sram_cell_6t_5 inst_cell_88_97 (.BL(BL97),.BLN(BLN97),.WL(WL88));
sram_cell_6t_5 inst_cell_88_98 (.BL(BL98),.BLN(BLN98),.WL(WL88));
sram_cell_6t_5 inst_cell_88_99 (.BL(BL99),.BLN(BLN99),.WL(WL88));
sram_cell_6t_5 inst_cell_88_100 (.BL(BL100),.BLN(BLN100),.WL(WL88));
sram_cell_6t_5 inst_cell_88_101 (.BL(BL101),.BLN(BLN101),.WL(WL88));
sram_cell_6t_5 inst_cell_88_102 (.BL(BL102),.BLN(BLN102),.WL(WL88));
sram_cell_6t_5 inst_cell_88_103 (.BL(BL103),.BLN(BLN103),.WL(WL88));
sram_cell_6t_5 inst_cell_88_104 (.BL(BL104),.BLN(BLN104),.WL(WL88));
sram_cell_6t_5 inst_cell_88_105 (.BL(BL105),.BLN(BLN105),.WL(WL88));
sram_cell_6t_5 inst_cell_88_106 (.BL(BL106),.BLN(BLN106),.WL(WL88));
sram_cell_6t_5 inst_cell_88_107 (.BL(BL107),.BLN(BLN107),.WL(WL88));
sram_cell_6t_5 inst_cell_88_108 (.BL(BL108),.BLN(BLN108),.WL(WL88));
sram_cell_6t_5 inst_cell_88_109 (.BL(BL109),.BLN(BLN109),.WL(WL88));
sram_cell_6t_5 inst_cell_88_110 (.BL(BL110),.BLN(BLN110),.WL(WL88));
sram_cell_6t_5 inst_cell_88_111 (.BL(BL111),.BLN(BLN111),.WL(WL88));
sram_cell_6t_5 inst_cell_88_112 (.BL(BL112),.BLN(BLN112),.WL(WL88));
sram_cell_6t_5 inst_cell_88_113 (.BL(BL113),.BLN(BLN113),.WL(WL88));
sram_cell_6t_5 inst_cell_88_114 (.BL(BL114),.BLN(BLN114),.WL(WL88));
sram_cell_6t_5 inst_cell_88_115 (.BL(BL115),.BLN(BLN115),.WL(WL88));
sram_cell_6t_5 inst_cell_88_116 (.BL(BL116),.BLN(BLN116),.WL(WL88));
sram_cell_6t_5 inst_cell_88_117 (.BL(BL117),.BLN(BLN117),.WL(WL88));
sram_cell_6t_5 inst_cell_88_118 (.BL(BL118),.BLN(BLN118),.WL(WL88));
sram_cell_6t_5 inst_cell_88_119 (.BL(BL119),.BLN(BLN119),.WL(WL88));
sram_cell_6t_5 inst_cell_88_120 (.BL(BL120),.BLN(BLN120),.WL(WL88));
sram_cell_6t_5 inst_cell_88_121 (.BL(BL121),.BLN(BLN121),.WL(WL88));
sram_cell_6t_5 inst_cell_88_122 (.BL(BL122),.BLN(BLN122),.WL(WL88));
sram_cell_6t_5 inst_cell_88_123 (.BL(BL123),.BLN(BLN123),.WL(WL88));
sram_cell_6t_5 inst_cell_88_124 (.BL(BL124),.BLN(BLN124),.WL(WL88));
sram_cell_6t_5 inst_cell_88_125 (.BL(BL125),.BLN(BLN125),.WL(WL88));
sram_cell_6t_5 inst_cell_88_126 (.BL(BL126),.BLN(BLN126),.WL(WL88));
sram_cell_6t_5 inst_cell_88_127 (.BL(BL127),.BLN(BLN127),.WL(WL88));
sram_cell_6t_5 inst_cell_89_0 (.BL(BL0),.BLN(BLN0),.WL(WL89));
sram_cell_6t_5 inst_cell_89_1 (.BL(BL1),.BLN(BLN1),.WL(WL89));
sram_cell_6t_5 inst_cell_89_2 (.BL(BL2),.BLN(BLN2),.WL(WL89));
sram_cell_6t_5 inst_cell_89_3 (.BL(BL3),.BLN(BLN3),.WL(WL89));
sram_cell_6t_5 inst_cell_89_4 (.BL(BL4),.BLN(BLN4),.WL(WL89));
sram_cell_6t_5 inst_cell_89_5 (.BL(BL5),.BLN(BLN5),.WL(WL89));
sram_cell_6t_5 inst_cell_89_6 (.BL(BL6),.BLN(BLN6),.WL(WL89));
sram_cell_6t_5 inst_cell_89_7 (.BL(BL7),.BLN(BLN7),.WL(WL89));
sram_cell_6t_5 inst_cell_89_8 (.BL(BL8),.BLN(BLN8),.WL(WL89));
sram_cell_6t_5 inst_cell_89_9 (.BL(BL9),.BLN(BLN9),.WL(WL89));
sram_cell_6t_5 inst_cell_89_10 (.BL(BL10),.BLN(BLN10),.WL(WL89));
sram_cell_6t_5 inst_cell_89_11 (.BL(BL11),.BLN(BLN11),.WL(WL89));
sram_cell_6t_5 inst_cell_89_12 (.BL(BL12),.BLN(BLN12),.WL(WL89));
sram_cell_6t_5 inst_cell_89_13 (.BL(BL13),.BLN(BLN13),.WL(WL89));
sram_cell_6t_5 inst_cell_89_14 (.BL(BL14),.BLN(BLN14),.WL(WL89));
sram_cell_6t_5 inst_cell_89_15 (.BL(BL15),.BLN(BLN15),.WL(WL89));
sram_cell_6t_5 inst_cell_89_16 (.BL(BL16),.BLN(BLN16),.WL(WL89));
sram_cell_6t_5 inst_cell_89_17 (.BL(BL17),.BLN(BLN17),.WL(WL89));
sram_cell_6t_5 inst_cell_89_18 (.BL(BL18),.BLN(BLN18),.WL(WL89));
sram_cell_6t_5 inst_cell_89_19 (.BL(BL19),.BLN(BLN19),.WL(WL89));
sram_cell_6t_5 inst_cell_89_20 (.BL(BL20),.BLN(BLN20),.WL(WL89));
sram_cell_6t_5 inst_cell_89_21 (.BL(BL21),.BLN(BLN21),.WL(WL89));
sram_cell_6t_5 inst_cell_89_22 (.BL(BL22),.BLN(BLN22),.WL(WL89));
sram_cell_6t_5 inst_cell_89_23 (.BL(BL23),.BLN(BLN23),.WL(WL89));
sram_cell_6t_5 inst_cell_89_24 (.BL(BL24),.BLN(BLN24),.WL(WL89));
sram_cell_6t_5 inst_cell_89_25 (.BL(BL25),.BLN(BLN25),.WL(WL89));
sram_cell_6t_5 inst_cell_89_26 (.BL(BL26),.BLN(BLN26),.WL(WL89));
sram_cell_6t_5 inst_cell_89_27 (.BL(BL27),.BLN(BLN27),.WL(WL89));
sram_cell_6t_5 inst_cell_89_28 (.BL(BL28),.BLN(BLN28),.WL(WL89));
sram_cell_6t_5 inst_cell_89_29 (.BL(BL29),.BLN(BLN29),.WL(WL89));
sram_cell_6t_5 inst_cell_89_30 (.BL(BL30),.BLN(BLN30),.WL(WL89));
sram_cell_6t_5 inst_cell_89_31 (.BL(BL31),.BLN(BLN31),.WL(WL89));
sram_cell_6t_5 inst_cell_89_32 (.BL(BL32),.BLN(BLN32),.WL(WL89));
sram_cell_6t_5 inst_cell_89_33 (.BL(BL33),.BLN(BLN33),.WL(WL89));
sram_cell_6t_5 inst_cell_89_34 (.BL(BL34),.BLN(BLN34),.WL(WL89));
sram_cell_6t_5 inst_cell_89_35 (.BL(BL35),.BLN(BLN35),.WL(WL89));
sram_cell_6t_5 inst_cell_89_36 (.BL(BL36),.BLN(BLN36),.WL(WL89));
sram_cell_6t_5 inst_cell_89_37 (.BL(BL37),.BLN(BLN37),.WL(WL89));
sram_cell_6t_5 inst_cell_89_38 (.BL(BL38),.BLN(BLN38),.WL(WL89));
sram_cell_6t_5 inst_cell_89_39 (.BL(BL39),.BLN(BLN39),.WL(WL89));
sram_cell_6t_5 inst_cell_89_40 (.BL(BL40),.BLN(BLN40),.WL(WL89));
sram_cell_6t_5 inst_cell_89_41 (.BL(BL41),.BLN(BLN41),.WL(WL89));
sram_cell_6t_5 inst_cell_89_42 (.BL(BL42),.BLN(BLN42),.WL(WL89));
sram_cell_6t_5 inst_cell_89_43 (.BL(BL43),.BLN(BLN43),.WL(WL89));
sram_cell_6t_5 inst_cell_89_44 (.BL(BL44),.BLN(BLN44),.WL(WL89));
sram_cell_6t_5 inst_cell_89_45 (.BL(BL45),.BLN(BLN45),.WL(WL89));
sram_cell_6t_5 inst_cell_89_46 (.BL(BL46),.BLN(BLN46),.WL(WL89));
sram_cell_6t_5 inst_cell_89_47 (.BL(BL47),.BLN(BLN47),.WL(WL89));
sram_cell_6t_5 inst_cell_89_48 (.BL(BL48),.BLN(BLN48),.WL(WL89));
sram_cell_6t_5 inst_cell_89_49 (.BL(BL49),.BLN(BLN49),.WL(WL89));
sram_cell_6t_5 inst_cell_89_50 (.BL(BL50),.BLN(BLN50),.WL(WL89));
sram_cell_6t_5 inst_cell_89_51 (.BL(BL51),.BLN(BLN51),.WL(WL89));
sram_cell_6t_5 inst_cell_89_52 (.BL(BL52),.BLN(BLN52),.WL(WL89));
sram_cell_6t_5 inst_cell_89_53 (.BL(BL53),.BLN(BLN53),.WL(WL89));
sram_cell_6t_5 inst_cell_89_54 (.BL(BL54),.BLN(BLN54),.WL(WL89));
sram_cell_6t_5 inst_cell_89_55 (.BL(BL55),.BLN(BLN55),.WL(WL89));
sram_cell_6t_5 inst_cell_89_56 (.BL(BL56),.BLN(BLN56),.WL(WL89));
sram_cell_6t_5 inst_cell_89_57 (.BL(BL57),.BLN(BLN57),.WL(WL89));
sram_cell_6t_5 inst_cell_89_58 (.BL(BL58),.BLN(BLN58),.WL(WL89));
sram_cell_6t_5 inst_cell_89_59 (.BL(BL59),.BLN(BLN59),.WL(WL89));
sram_cell_6t_5 inst_cell_89_60 (.BL(BL60),.BLN(BLN60),.WL(WL89));
sram_cell_6t_5 inst_cell_89_61 (.BL(BL61),.BLN(BLN61),.WL(WL89));
sram_cell_6t_5 inst_cell_89_62 (.BL(BL62),.BLN(BLN62),.WL(WL89));
sram_cell_6t_5 inst_cell_89_63 (.BL(BL63),.BLN(BLN63),.WL(WL89));
sram_cell_6t_5 inst_cell_89_64 (.BL(BL64),.BLN(BLN64),.WL(WL89));
sram_cell_6t_5 inst_cell_89_65 (.BL(BL65),.BLN(BLN65),.WL(WL89));
sram_cell_6t_5 inst_cell_89_66 (.BL(BL66),.BLN(BLN66),.WL(WL89));
sram_cell_6t_5 inst_cell_89_67 (.BL(BL67),.BLN(BLN67),.WL(WL89));
sram_cell_6t_5 inst_cell_89_68 (.BL(BL68),.BLN(BLN68),.WL(WL89));
sram_cell_6t_5 inst_cell_89_69 (.BL(BL69),.BLN(BLN69),.WL(WL89));
sram_cell_6t_5 inst_cell_89_70 (.BL(BL70),.BLN(BLN70),.WL(WL89));
sram_cell_6t_5 inst_cell_89_71 (.BL(BL71),.BLN(BLN71),.WL(WL89));
sram_cell_6t_5 inst_cell_89_72 (.BL(BL72),.BLN(BLN72),.WL(WL89));
sram_cell_6t_5 inst_cell_89_73 (.BL(BL73),.BLN(BLN73),.WL(WL89));
sram_cell_6t_5 inst_cell_89_74 (.BL(BL74),.BLN(BLN74),.WL(WL89));
sram_cell_6t_5 inst_cell_89_75 (.BL(BL75),.BLN(BLN75),.WL(WL89));
sram_cell_6t_5 inst_cell_89_76 (.BL(BL76),.BLN(BLN76),.WL(WL89));
sram_cell_6t_5 inst_cell_89_77 (.BL(BL77),.BLN(BLN77),.WL(WL89));
sram_cell_6t_5 inst_cell_89_78 (.BL(BL78),.BLN(BLN78),.WL(WL89));
sram_cell_6t_5 inst_cell_89_79 (.BL(BL79),.BLN(BLN79),.WL(WL89));
sram_cell_6t_5 inst_cell_89_80 (.BL(BL80),.BLN(BLN80),.WL(WL89));
sram_cell_6t_5 inst_cell_89_81 (.BL(BL81),.BLN(BLN81),.WL(WL89));
sram_cell_6t_5 inst_cell_89_82 (.BL(BL82),.BLN(BLN82),.WL(WL89));
sram_cell_6t_5 inst_cell_89_83 (.BL(BL83),.BLN(BLN83),.WL(WL89));
sram_cell_6t_5 inst_cell_89_84 (.BL(BL84),.BLN(BLN84),.WL(WL89));
sram_cell_6t_5 inst_cell_89_85 (.BL(BL85),.BLN(BLN85),.WL(WL89));
sram_cell_6t_5 inst_cell_89_86 (.BL(BL86),.BLN(BLN86),.WL(WL89));
sram_cell_6t_5 inst_cell_89_87 (.BL(BL87),.BLN(BLN87),.WL(WL89));
sram_cell_6t_5 inst_cell_89_88 (.BL(BL88),.BLN(BLN88),.WL(WL89));
sram_cell_6t_5 inst_cell_89_89 (.BL(BL89),.BLN(BLN89),.WL(WL89));
sram_cell_6t_5 inst_cell_89_90 (.BL(BL90),.BLN(BLN90),.WL(WL89));
sram_cell_6t_5 inst_cell_89_91 (.BL(BL91),.BLN(BLN91),.WL(WL89));
sram_cell_6t_5 inst_cell_89_92 (.BL(BL92),.BLN(BLN92),.WL(WL89));
sram_cell_6t_5 inst_cell_89_93 (.BL(BL93),.BLN(BLN93),.WL(WL89));
sram_cell_6t_5 inst_cell_89_94 (.BL(BL94),.BLN(BLN94),.WL(WL89));
sram_cell_6t_5 inst_cell_89_95 (.BL(BL95),.BLN(BLN95),.WL(WL89));
sram_cell_6t_5 inst_cell_89_96 (.BL(BL96),.BLN(BLN96),.WL(WL89));
sram_cell_6t_5 inst_cell_89_97 (.BL(BL97),.BLN(BLN97),.WL(WL89));
sram_cell_6t_5 inst_cell_89_98 (.BL(BL98),.BLN(BLN98),.WL(WL89));
sram_cell_6t_5 inst_cell_89_99 (.BL(BL99),.BLN(BLN99),.WL(WL89));
sram_cell_6t_5 inst_cell_89_100 (.BL(BL100),.BLN(BLN100),.WL(WL89));
sram_cell_6t_5 inst_cell_89_101 (.BL(BL101),.BLN(BLN101),.WL(WL89));
sram_cell_6t_5 inst_cell_89_102 (.BL(BL102),.BLN(BLN102),.WL(WL89));
sram_cell_6t_5 inst_cell_89_103 (.BL(BL103),.BLN(BLN103),.WL(WL89));
sram_cell_6t_5 inst_cell_89_104 (.BL(BL104),.BLN(BLN104),.WL(WL89));
sram_cell_6t_5 inst_cell_89_105 (.BL(BL105),.BLN(BLN105),.WL(WL89));
sram_cell_6t_5 inst_cell_89_106 (.BL(BL106),.BLN(BLN106),.WL(WL89));
sram_cell_6t_5 inst_cell_89_107 (.BL(BL107),.BLN(BLN107),.WL(WL89));
sram_cell_6t_5 inst_cell_89_108 (.BL(BL108),.BLN(BLN108),.WL(WL89));
sram_cell_6t_5 inst_cell_89_109 (.BL(BL109),.BLN(BLN109),.WL(WL89));
sram_cell_6t_5 inst_cell_89_110 (.BL(BL110),.BLN(BLN110),.WL(WL89));
sram_cell_6t_5 inst_cell_89_111 (.BL(BL111),.BLN(BLN111),.WL(WL89));
sram_cell_6t_5 inst_cell_89_112 (.BL(BL112),.BLN(BLN112),.WL(WL89));
sram_cell_6t_5 inst_cell_89_113 (.BL(BL113),.BLN(BLN113),.WL(WL89));
sram_cell_6t_5 inst_cell_89_114 (.BL(BL114),.BLN(BLN114),.WL(WL89));
sram_cell_6t_5 inst_cell_89_115 (.BL(BL115),.BLN(BLN115),.WL(WL89));
sram_cell_6t_5 inst_cell_89_116 (.BL(BL116),.BLN(BLN116),.WL(WL89));
sram_cell_6t_5 inst_cell_89_117 (.BL(BL117),.BLN(BLN117),.WL(WL89));
sram_cell_6t_5 inst_cell_89_118 (.BL(BL118),.BLN(BLN118),.WL(WL89));
sram_cell_6t_5 inst_cell_89_119 (.BL(BL119),.BLN(BLN119),.WL(WL89));
sram_cell_6t_5 inst_cell_89_120 (.BL(BL120),.BLN(BLN120),.WL(WL89));
sram_cell_6t_5 inst_cell_89_121 (.BL(BL121),.BLN(BLN121),.WL(WL89));
sram_cell_6t_5 inst_cell_89_122 (.BL(BL122),.BLN(BLN122),.WL(WL89));
sram_cell_6t_5 inst_cell_89_123 (.BL(BL123),.BLN(BLN123),.WL(WL89));
sram_cell_6t_5 inst_cell_89_124 (.BL(BL124),.BLN(BLN124),.WL(WL89));
sram_cell_6t_5 inst_cell_89_125 (.BL(BL125),.BLN(BLN125),.WL(WL89));
sram_cell_6t_5 inst_cell_89_126 (.BL(BL126),.BLN(BLN126),.WL(WL89));
sram_cell_6t_5 inst_cell_89_127 (.BL(BL127),.BLN(BLN127),.WL(WL89));
sram_cell_6t_5 inst_cell_90_0 (.BL(BL0),.BLN(BLN0),.WL(WL90));
sram_cell_6t_5 inst_cell_90_1 (.BL(BL1),.BLN(BLN1),.WL(WL90));
sram_cell_6t_5 inst_cell_90_2 (.BL(BL2),.BLN(BLN2),.WL(WL90));
sram_cell_6t_5 inst_cell_90_3 (.BL(BL3),.BLN(BLN3),.WL(WL90));
sram_cell_6t_5 inst_cell_90_4 (.BL(BL4),.BLN(BLN4),.WL(WL90));
sram_cell_6t_5 inst_cell_90_5 (.BL(BL5),.BLN(BLN5),.WL(WL90));
sram_cell_6t_5 inst_cell_90_6 (.BL(BL6),.BLN(BLN6),.WL(WL90));
sram_cell_6t_5 inst_cell_90_7 (.BL(BL7),.BLN(BLN7),.WL(WL90));
sram_cell_6t_5 inst_cell_90_8 (.BL(BL8),.BLN(BLN8),.WL(WL90));
sram_cell_6t_5 inst_cell_90_9 (.BL(BL9),.BLN(BLN9),.WL(WL90));
sram_cell_6t_5 inst_cell_90_10 (.BL(BL10),.BLN(BLN10),.WL(WL90));
sram_cell_6t_5 inst_cell_90_11 (.BL(BL11),.BLN(BLN11),.WL(WL90));
sram_cell_6t_5 inst_cell_90_12 (.BL(BL12),.BLN(BLN12),.WL(WL90));
sram_cell_6t_5 inst_cell_90_13 (.BL(BL13),.BLN(BLN13),.WL(WL90));
sram_cell_6t_5 inst_cell_90_14 (.BL(BL14),.BLN(BLN14),.WL(WL90));
sram_cell_6t_5 inst_cell_90_15 (.BL(BL15),.BLN(BLN15),.WL(WL90));
sram_cell_6t_5 inst_cell_90_16 (.BL(BL16),.BLN(BLN16),.WL(WL90));
sram_cell_6t_5 inst_cell_90_17 (.BL(BL17),.BLN(BLN17),.WL(WL90));
sram_cell_6t_5 inst_cell_90_18 (.BL(BL18),.BLN(BLN18),.WL(WL90));
sram_cell_6t_5 inst_cell_90_19 (.BL(BL19),.BLN(BLN19),.WL(WL90));
sram_cell_6t_5 inst_cell_90_20 (.BL(BL20),.BLN(BLN20),.WL(WL90));
sram_cell_6t_5 inst_cell_90_21 (.BL(BL21),.BLN(BLN21),.WL(WL90));
sram_cell_6t_5 inst_cell_90_22 (.BL(BL22),.BLN(BLN22),.WL(WL90));
sram_cell_6t_5 inst_cell_90_23 (.BL(BL23),.BLN(BLN23),.WL(WL90));
sram_cell_6t_5 inst_cell_90_24 (.BL(BL24),.BLN(BLN24),.WL(WL90));
sram_cell_6t_5 inst_cell_90_25 (.BL(BL25),.BLN(BLN25),.WL(WL90));
sram_cell_6t_5 inst_cell_90_26 (.BL(BL26),.BLN(BLN26),.WL(WL90));
sram_cell_6t_5 inst_cell_90_27 (.BL(BL27),.BLN(BLN27),.WL(WL90));
sram_cell_6t_5 inst_cell_90_28 (.BL(BL28),.BLN(BLN28),.WL(WL90));
sram_cell_6t_5 inst_cell_90_29 (.BL(BL29),.BLN(BLN29),.WL(WL90));
sram_cell_6t_5 inst_cell_90_30 (.BL(BL30),.BLN(BLN30),.WL(WL90));
sram_cell_6t_5 inst_cell_90_31 (.BL(BL31),.BLN(BLN31),.WL(WL90));
sram_cell_6t_5 inst_cell_90_32 (.BL(BL32),.BLN(BLN32),.WL(WL90));
sram_cell_6t_5 inst_cell_90_33 (.BL(BL33),.BLN(BLN33),.WL(WL90));
sram_cell_6t_5 inst_cell_90_34 (.BL(BL34),.BLN(BLN34),.WL(WL90));
sram_cell_6t_5 inst_cell_90_35 (.BL(BL35),.BLN(BLN35),.WL(WL90));
sram_cell_6t_5 inst_cell_90_36 (.BL(BL36),.BLN(BLN36),.WL(WL90));
sram_cell_6t_5 inst_cell_90_37 (.BL(BL37),.BLN(BLN37),.WL(WL90));
sram_cell_6t_5 inst_cell_90_38 (.BL(BL38),.BLN(BLN38),.WL(WL90));
sram_cell_6t_5 inst_cell_90_39 (.BL(BL39),.BLN(BLN39),.WL(WL90));
sram_cell_6t_5 inst_cell_90_40 (.BL(BL40),.BLN(BLN40),.WL(WL90));
sram_cell_6t_5 inst_cell_90_41 (.BL(BL41),.BLN(BLN41),.WL(WL90));
sram_cell_6t_5 inst_cell_90_42 (.BL(BL42),.BLN(BLN42),.WL(WL90));
sram_cell_6t_5 inst_cell_90_43 (.BL(BL43),.BLN(BLN43),.WL(WL90));
sram_cell_6t_5 inst_cell_90_44 (.BL(BL44),.BLN(BLN44),.WL(WL90));
sram_cell_6t_5 inst_cell_90_45 (.BL(BL45),.BLN(BLN45),.WL(WL90));
sram_cell_6t_5 inst_cell_90_46 (.BL(BL46),.BLN(BLN46),.WL(WL90));
sram_cell_6t_5 inst_cell_90_47 (.BL(BL47),.BLN(BLN47),.WL(WL90));
sram_cell_6t_5 inst_cell_90_48 (.BL(BL48),.BLN(BLN48),.WL(WL90));
sram_cell_6t_5 inst_cell_90_49 (.BL(BL49),.BLN(BLN49),.WL(WL90));
sram_cell_6t_5 inst_cell_90_50 (.BL(BL50),.BLN(BLN50),.WL(WL90));
sram_cell_6t_5 inst_cell_90_51 (.BL(BL51),.BLN(BLN51),.WL(WL90));
sram_cell_6t_5 inst_cell_90_52 (.BL(BL52),.BLN(BLN52),.WL(WL90));
sram_cell_6t_5 inst_cell_90_53 (.BL(BL53),.BLN(BLN53),.WL(WL90));
sram_cell_6t_5 inst_cell_90_54 (.BL(BL54),.BLN(BLN54),.WL(WL90));
sram_cell_6t_5 inst_cell_90_55 (.BL(BL55),.BLN(BLN55),.WL(WL90));
sram_cell_6t_5 inst_cell_90_56 (.BL(BL56),.BLN(BLN56),.WL(WL90));
sram_cell_6t_5 inst_cell_90_57 (.BL(BL57),.BLN(BLN57),.WL(WL90));
sram_cell_6t_5 inst_cell_90_58 (.BL(BL58),.BLN(BLN58),.WL(WL90));
sram_cell_6t_5 inst_cell_90_59 (.BL(BL59),.BLN(BLN59),.WL(WL90));
sram_cell_6t_5 inst_cell_90_60 (.BL(BL60),.BLN(BLN60),.WL(WL90));
sram_cell_6t_5 inst_cell_90_61 (.BL(BL61),.BLN(BLN61),.WL(WL90));
sram_cell_6t_5 inst_cell_90_62 (.BL(BL62),.BLN(BLN62),.WL(WL90));
sram_cell_6t_5 inst_cell_90_63 (.BL(BL63),.BLN(BLN63),.WL(WL90));
sram_cell_6t_5 inst_cell_90_64 (.BL(BL64),.BLN(BLN64),.WL(WL90));
sram_cell_6t_5 inst_cell_90_65 (.BL(BL65),.BLN(BLN65),.WL(WL90));
sram_cell_6t_5 inst_cell_90_66 (.BL(BL66),.BLN(BLN66),.WL(WL90));
sram_cell_6t_5 inst_cell_90_67 (.BL(BL67),.BLN(BLN67),.WL(WL90));
sram_cell_6t_5 inst_cell_90_68 (.BL(BL68),.BLN(BLN68),.WL(WL90));
sram_cell_6t_5 inst_cell_90_69 (.BL(BL69),.BLN(BLN69),.WL(WL90));
sram_cell_6t_5 inst_cell_90_70 (.BL(BL70),.BLN(BLN70),.WL(WL90));
sram_cell_6t_5 inst_cell_90_71 (.BL(BL71),.BLN(BLN71),.WL(WL90));
sram_cell_6t_5 inst_cell_90_72 (.BL(BL72),.BLN(BLN72),.WL(WL90));
sram_cell_6t_5 inst_cell_90_73 (.BL(BL73),.BLN(BLN73),.WL(WL90));
sram_cell_6t_5 inst_cell_90_74 (.BL(BL74),.BLN(BLN74),.WL(WL90));
sram_cell_6t_5 inst_cell_90_75 (.BL(BL75),.BLN(BLN75),.WL(WL90));
sram_cell_6t_5 inst_cell_90_76 (.BL(BL76),.BLN(BLN76),.WL(WL90));
sram_cell_6t_5 inst_cell_90_77 (.BL(BL77),.BLN(BLN77),.WL(WL90));
sram_cell_6t_5 inst_cell_90_78 (.BL(BL78),.BLN(BLN78),.WL(WL90));
sram_cell_6t_5 inst_cell_90_79 (.BL(BL79),.BLN(BLN79),.WL(WL90));
sram_cell_6t_5 inst_cell_90_80 (.BL(BL80),.BLN(BLN80),.WL(WL90));
sram_cell_6t_5 inst_cell_90_81 (.BL(BL81),.BLN(BLN81),.WL(WL90));
sram_cell_6t_5 inst_cell_90_82 (.BL(BL82),.BLN(BLN82),.WL(WL90));
sram_cell_6t_5 inst_cell_90_83 (.BL(BL83),.BLN(BLN83),.WL(WL90));
sram_cell_6t_5 inst_cell_90_84 (.BL(BL84),.BLN(BLN84),.WL(WL90));
sram_cell_6t_5 inst_cell_90_85 (.BL(BL85),.BLN(BLN85),.WL(WL90));
sram_cell_6t_5 inst_cell_90_86 (.BL(BL86),.BLN(BLN86),.WL(WL90));
sram_cell_6t_5 inst_cell_90_87 (.BL(BL87),.BLN(BLN87),.WL(WL90));
sram_cell_6t_5 inst_cell_90_88 (.BL(BL88),.BLN(BLN88),.WL(WL90));
sram_cell_6t_5 inst_cell_90_89 (.BL(BL89),.BLN(BLN89),.WL(WL90));
sram_cell_6t_5 inst_cell_90_90 (.BL(BL90),.BLN(BLN90),.WL(WL90));
sram_cell_6t_5 inst_cell_90_91 (.BL(BL91),.BLN(BLN91),.WL(WL90));
sram_cell_6t_5 inst_cell_90_92 (.BL(BL92),.BLN(BLN92),.WL(WL90));
sram_cell_6t_5 inst_cell_90_93 (.BL(BL93),.BLN(BLN93),.WL(WL90));
sram_cell_6t_5 inst_cell_90_94 (.BL(BL94),.BLN(BLN94),.WL(WL90));
sram_cell_6t_5 inst_cell_90_95 (.BL(BL95),.BLN(BLN95),.WL(WL90));
sram_cell_6t_5 inst_cell_90_96 (.BL(BL96),.BLN(BLN96),.WL(WL90));
sram_cell_6t_5 inst_cell_90_97 (.BL(BL97),.BLN(BLN97),.WL(WL90));
sram_cell_6t_5 inst_cell_90_98 (.BL(BL98),.BLN(BLN98),.WL(WL90));
sram_cell_6t_5 inst_cell_90_99 (.BL(BL99),.BLN(BLN99),.WL(WL90));
sram_cell_6t_5 inst_cell_90_100 (.BL(BL100),.BLN(BLN100),.WL(WL90));
sram_cell_6t_5 inst_cell_90_101 (.BL(BL101),.BLN(BLN101),.WL(WL90));
sram_cell_6t_5 inst_cell_90_102 (.BL(BL102),.BLN(BLN102),.WL(WL90));
sram_cell_6t_5 inst_cell_90_103 (.BL(BL103),.BLN(BLN103),.WL(WL90));
sram_cell_6t_5 inst_cell_90_104 (.BL(BL104),.BLN(BLN104),.WL(WL90));
sram_cell_6t_5 inst_cell_90_105 (.BL(BL105),.BLN(BLN105),.WL(WL90));
sram_cell_6t_5 inst_cell_90_106 (.BL(BL106),.BLN(BLN106),.WL(WL90));
sram_cell_6t_5 inst_cell_90_107 (.BL(BL107),.BLN(BLN107),.WL(WL90));
sram_cell_6t_5 inst_cell_90_108 (.BL(BL108),.BLN(BLN108),.WL(WL90));
sram_cell_6t_5 inst_cell_90_109 (.BL(BL109),.BLN(BLN109),.WL(WL90));
sram_cell_6t_5 inst_cell_90_110 (.BL(BL110),.BLN(BLN110),.WL(WL90));
sram_cell_6t_5 inst_cell_90_111 (.BL(BL111),.BLN(BLN111),.WL(WL90));
sram_cell_6t_5 inst_cell_90_112 (.BL(BL112),.BLN(BLN112),.WL(WL90));
sram_cell_6t_5 inst_cell_90_113 (.BL(BL113),.BLN(BLN113),.WL(WL90));
sram_cell_6t_5 inst_cell_90_114 (.BL(BL114),.BLN(BLN114),.WL(WL90));
sram_cell_6t_5 inst_cell_90_115 (.BL(BL115),.BLN(BLN115),.WL(WL90));
sram_cell_6t_5 inst_cell_90_116 (.BL(BL116),.BLN(BLN116),.WL(WL90));
sram_cell_6t_5 inst_cell_90_117 (.BL(BL117),.BLN(BLN117),.WL(WL90));
sram_cell_6t_5 inst_cell_90_118 (.BL(BL118),.BLN(BLN118),.WL(WL90));
sram_cell_6t_5 inst_cell_90_119 (.BL(BL119),.BLN(BLN119),.WL(WL90));
sram_cell_6t_5 inst_cell_90_120 (.BL(BL120),.BLN(BLN120),.WL(WL90));
sram_cell_6t_5 inst_cell_90_121 (.BL(BL121),.BLN(BLN121),.WL(WL90));
sram_cell_6t_5 inst_cell_90_122 (.BL(BL122),.BLN(BLN122),.WL(WL90));
sram_cell_6t_5 inst_cell_90_123 (.BL(BL123),.BLN(BLN123),.WL(WL90));
sram_cell_6t_5 inst_cell_90_124 (.BL(BL124),.BLN(BLN124),.WL(WL90));
sram_cell_6t_5 inst_cell_90_125 (.BL(BL125),.BLN(BLN125),.WL(WL90));
sram_cell_6t_5 inst_cell_90_126 (.BL(BL126),.BLN(BLN126),.WL(WL90));
sram_cell_6t_5 inst_cell_90_127 (.BL(BL127),.BLN(BLN127),.WL(WL90));
sram_cell_6t_5 inst_cell_91_0 (.BL(BL0),.BLN(BLN0),.WL(WL91));
sram_cell_6t_5 inst_cell_91_1 (.BL(BL1),.BLN(BLN1),.WL(WL91));
sram_cell_6t_5 inst_cell_91_2 (.BL(BL2),.BLN(BLN2),.WL(WL91));
sram_cell_6t_5 inst_cell_91_3 (.BL(BL3),.BLN(BLN3),.WL(WL91));
sram_cell_6t_5 inst_cell_91_4 (.BL(BL4),.BLN(BLN4),.WL(WL91));
sram_cell_6t_5 inst_cell_91_5 (.BL(BL5),.BLN(BLN5),.WL(WL91));
sram_cell_6t_5 inst_cell_91_6 (.BL(BL6),.BLN(BLN6),.WL(WL91));
sram_cell_6t_5 inst_cell_91_7 (.BL(BL7),.BLN(BLN7),.WL(WL91));
sram_cell_6t_5 inst_cell_91_8 (.BL(BL8),.BLN(BLN8),.WL(WL91));
sram_cell_6t_5 inst_cell_91_9 (.BL(BL9),.BLN(BLN9),.WL(WL91));
sram_cell_6t_5 inst_cell_91_10 (.BL(BL10),.BLN(BLN10),.WL(WL91));
sram_cell_6t_5 inst_cell_91_11 (.BL(BL11),.BLN(BLN11),.WL(WL91));
sram_cell_6t_5 inst_cell_91_12 (.BL(BL12),.BLN(BLN12),.WL(WL91));
sram_cell_6t_5 inst_cell_91_13 (.BL(BL13),.BLN(BLN13),.WL(WL91));
sram_cell_6t_5 inst_cell_91_14 (.BL(BL14),.BLN(BLN14),.WL(WL91));
sram_cell_6t_5 inst_cell_91_15 (.BL(BL15),.BLN(BLN15),.WL(WL91));
sram_cell_6t_5 inst_cell_91_16 (.BL(BL16),.BLN(BLN16),.WL(WL91));
sram_cell_6t_5 inst_cell_91_17 (.BL(BL17),.BLN(BLN17),.WL(WL91));
sram_cell_6t_5 inst_cell_91_18 (.BL(BL18),.BLN(BLN18),.WL(WL91));
sram_cell_6t_5 inst_cell_91_19 (.BL(BL19),.BLN(BLN19),.WL(WL91));
sram_cell_6t_5 inst_cell_91_20 (.BL(BL20),.BLN(BLN20),.WL(WL91));
sram_cell_6t_5 inst_cell_91_21 (.BL(BL21),.BLN(BLN21),.WL(WL91));
sram_cell_6t_5 inst_cell_91_22 (.BL(BL22),.BLN(BLN22),.WL(WL91));
sram_cell_6t_5 inst_cell_91_23 (.BL(BL23),.BLN(BLN23),.WL(WL91));
sram_cell_6t_5 inst_cell_91_24 (.BL(BL24),.BLN(BLN24),.WL(WL91));
sram_cell_6t_5 inst_cell_91_25 (.BL(BL25),.BLN(BLN25),.WL(WL91));
sram_cell_6t_5 inst_cell_91_26 (.BL(BL26),.BLN(BLN26),.WL(WL91));
sram_cell_6t_5 inst_cell_91_27 (.BL(BL27),.BLN(BLN27),.WL(WL91));
sram_cell_6t_5 inst_cell_91_28 (.BL(BL28),.BLN(BLN28),.WL(WL91));
sram_cell_6t_5 inst_cell_91_29 (.BL(BL29),.BLN(BLN29),.WL(WL91));
sram_cell_6t_5 inst_cell_91_30 (.BL(BL30),.BLN(BLN30),.WL(WL91));
sram_cell_6t_5 inst_cell_91_31 (.BL(BL31),.BLN(BLN31),.WL(WL91));
sram_cell_6t_5 inst_cell_91_32 (.BL(BL32),.BLN(BLN32),.WL(WL91));
sram_cell_6t_5 inst_cell_91_33 (.BL(BL33),.BLN(BLN33),.WL(WL91));
sram_cell_6t_5 inst_cell_91_34 (.BL(BL34),.BLN(BLN34),.WL(WL91));
sram_cell_6t_5 inst_cell_91_35 (.BL(BL35),.BLN(BLN35),.WL(WL91));
sram_cell_6t_5 inst_cell_91_36 (.BL(BL36),.BLN(BLN36),.WL(WL91));
sram_cell_6t_5 inst_cell_91_37 (.BL(BL37),.BLN(BLN37),.WL(WL91));
sram_cell_6t_5 inst_cell_91_38 (.BL(BL38),.BLN(BLN38),.WL(WL91));
sram_cell_6t_5 inst_cell_91_39 (.BL(BL39),.BLN(BLN39),.WL(WL91));
sram_cell_6t_5 inst_cell_91_40 (.BL(BL40),.BLN(BLN40),.WL(WL91));
sram_cell_6t_5 inst_cell_91_41 (.BL(BL41),.BLN(BLN41),.WL(WL91));
sram_cell_6t_5 inst_cell_91_42 (.BL(BL42),.BLN(BLN42),.WL(WL91));
sram_cell_6t_5 inst_cell_91_43 (.BL(BL43),.BLN(BLN43),.WL(WL91));
sram_cell_6t_5 inst_cell_91_44 (.BL(BL44),.BLN(BLN44),.WL(WL91));
sram_cell_6t_5 inst_cell_91_45 (.BL(BL45),.BLN(BLN45),.WL(WL91));
sram_cell_6t_5 inst_cell_91_46 (.BL(BL46),.BLN(BLN46),.WL(WL91));
sram_cell_6t_5 inst_cell_91_47 (.BL(BL47),.BLN(BLN47),.WL(WL91));
sram_cell_6t_5 inst_cell_91_48 (.BL(BL48),.BLN(BLN48),.WL(WL91));
sram_cell_6t_5 inst_cell_91_49 (.BL(BL49),.BLN(BLN49),.WL(WL91));
sram_cell_6t_5 inst_cell_91_50 (.BL(BL50),.BLN(BLN50),.WL(WL91));
sram_cell_6t_5 inst_cell_91_51 (.BL(BL51),.BLN(BLN51),.WL(WL91));
sram_cell_6t_5 inst_cell_91_52 (.BL(BL52),.BLN(BLN52),.WL(WL91));
sram_cell_6t_5 inst_cell_91_53 (.BL(BL53),.BLN(BLN53),.WL(WL91));
sram_cell_6t_5 inst_cell_91_54 (.BL(BL54),.BLN(BLN54),.WL(WL91));
sram_cell_6t_5 inst_cell_91_55 (.BL(BL55),.BLN(BLN55),.WL(WL91));
sram_cell_6t_5 inst_cell_91_56 (.BL(BL56),.BLN(BLN56),.WL(WL91));
sram_cell_6t_5 inst_cell_91_57 (.BL(BL57),.BLN(BLN57),.WL(WL91));
sram_cell_6t_5 inst_cell_91_58 (.BL(BL58),.BLN(BLN58),.WL(WL91));
sram_cell_6t_5 inst_cell_91_59 (.BL(BL59),.BLN(BLN59),.WL(WL91));
sram_cell_6t_5 inst_cell_91_60 (.BL(BL60),.BLN(BLN60),.WL(WL91));
sram_cell_6t_5 inst_cell_91_61 (.BL(BL61),.BLN(BLN61),.WL(WL91));
sram_cell_6t_5 inst_cell_91_62 (.BL(BL62),.BLN(BLN62),.WL(WL91));
sram_cell_6t_5 inst_cell_91_63 (.BL(BL63),.BLN(BLN63),.WL(WL91));
sram_cell_6t_5 inst_cell_91_64 (.BL(BL64),.BLN(BLN64),.WL(WL91));
sram_cell_6t_5 inst_cell_91_65 (.BL(BL65),.BLN(BLN65),.WL(WL91));
sram_cell_6t_5 inst_cell_91_66 (.BL(BL66),.BLN(BLN66),.WL(WL91));
sram_cell_6t_5 inst_cell_91_67 (.BL(BL67),.BLN(BLN67),.WL(WL91));
sram_cell_6t_5 inst_cell_91_68 (.BL(BL68),.BLN(BLN68),.WL(WL91));
sram_cell_6t_5 inst_cell_91_69 (.BL(BL69),.BLN(BLN69),.WL(WL91));
sram_cell_6t_5 inst_cell_91_70 (.BL(BL70),.BLN(BLN70),.WL(WL91));
sram_cell_6t_5 inst_cell_91_71 (.BL(BL71),.BLN(BLN71),.WL(WL91));
sram_cell_6t_5 inst_cell_91_72 (.BL(BL72),.BLN(BLN72),.WL(WL91));
sram_cell_6t_5 inst_cell_91_73 (.BL(BL73),.BLN(BLN73),.WL(WL91));
sram_cell_6t_5 inst_cell_91_74 (.BL(BL74),.BLN(BLN74),.WL(WL91));
sram_cell_6t_5 inst_cell_91_75 (.BL(BL75),.BLN(BLN75),.WL(WL91));
sram_cell_6t_5 inst_cell_91_76 (.BL(BL76),.BLN(BLN76),.WL(WL91));
sram_cell_6t_5 inst_cell_91_77 (.BL(BL77),.BLN(BLN77),.WL(WL91));
sram_cell_6t_5 inst_cell_91_78 (.BL(BL78),.BLN(BLN78),.WL(WL91));
sram_cell_6t_5 inst_cell_91_79 (.BL(BL79),.BLN(BLN79),.WL(WL91));
sram_cell_6t_5 inst_cell_91_80 (.BL(BL80),.BLN(BLN80),.WL(WL91));
sram_cell_6t_5 inst_cell_91_81 (.BL(BL81),.BLN(BLN81),.WL(WL91));
sram_cell_6t_5 inst_cell_91_82 (.BL(BL82),.BLN(BLN82),.WL(WL91));
sram_cell_6t_5 inst_cell_91_83 (.BL(BL83),.BLN(BLN83),.WL(WL91));
sram_cell_6t_5 inst_cell_91_84 (.BL(BL84),.BLN(BLN84),.WL(WL91));
sram_cell_6t_5 inst_cell_91_85 (.BL(BL85),.BLN(BLN85),.WL(WL91));
sram_cell_6t_5 inst_cell_91_86 (.BL(BL86),.BLN(BLN86),.WL(WL91));
sram_cell_6t_5 inst_cell_91_87 (.BL(BL87),.BLN(BLN87),.WL(WL91));
sram_cell_6t_5 inst_cell_91_88 (.BL(BL88),.BLN(BLN88),.WL(WL91));
sram_cell_6t_5 inst_cell_91_89 (.BL(BL89),.BLN(BLN89),.WL(WL91));
sram_cell_6t_5 inst_cell_91_90 (.BL(BL90),.BLN(BLN90),.WL(WL91));
sram_cell_6t_5 inst_cell_91_91 (.BL(BL91),.BLN(BLN91),.WL(WL91));
sram_cell_6t_5 inst_cell_91_92 (.BL(BL92),.BLN(BLN92),.WL(WL91));
sram_cell_6t_5 inst_cell_91_93 (.BL(BL93),.BLN(BLN93),.WL(WL91));
sram_cell_6t_5 inst_cell_91_94 (.BL(BL94),.BLN(BLN94),.WL(WL91));
sram_cell_6t_5 inst_cell_91_95 (.BL(BL95),.BLN(BLN95),.WL(WL91));
sram_cell_6t_5 inst_cell_91_96 (.BL(BL96),.BLN(BLN96),.WL(WL91));
sram_cell_6t_5 inst_cell_91_97 (.BL(BL97),.BLN(BLN97),.WL(WL91));
sram_cell_6t_5 inst_cell_91_98 (.BL(BL98),.BLN(BLN98),.WL(WL91));
sram_cell_6t_5 inst_cell_91_99 (.BL(BL99),.BLN(BLN99),.WL(WL91));
sram_cell_6t_5 inst_cell_91_100 (.BL(BL100),.BLN(BLN100),.WL(WL91));
sram_cell_6t_5 inst_cell_91_101 (.BL(BL101),.BLN(BLN101),.WL(WL91));
sram_cell_6t_5 inst_cell_91_102 (.BL(BL102),.BLN(BLN102),.WL(WL91));
sram_cell_6t_5 inst_cell_91_103 (.BL(BL103),.BLN(BLN103),.WL(WL91));
sram_cell_6t_5 inst_cell_91_104 (.BL(BL104),.BLN(BLN104),.WL(WL91));
sram_cell_6t_5 inst_cell_91_105 (.BL(BL105),.BLN(BLN105),.WL(WL91));
sram_cell_6t_5 inst_cell_91_106 (.BL(BL106),.BLN(BLN106),.WL(WL91));
sram_cell_6t_5 inst_cell_91_107 (.BL(BL107),.BLN(BLN107),.WL(WL91));
sram_cell_6t_5 inst_cell_91_108 (.BL(BL108),.BLN(BLN108),.WL(WL91));
sram_cell_6t_5 inst_cell_91_109 (.BL(BL109),.BLN(BLN109),.WL(WL91));
sram_cell_6t_5 inst_cell_91_110 (.BL(BL110),.BLN(BLN110),.WL(WL91));
sram_cell_6t_5 inst_cell_91_111 (.BL(BL111),.BLN(BLN111),.WL(WL91));
sram_cell_6t_5 inst_cell_91_112 (.BL(BL112),.BLN(BLN112),.WL(WL91));
sram_cell_6t_5 inst_cell_91_113 (.BL(BL113),.BLN(BLN113),.WL(WL91));
sram_cell_6t_5 inst_cell_91_114 (.BL(BL114),.BLN(BLN114),.WL(WL91));
sram_cell_6t_5 inst_cell_91_115 (.BL(BL115),.BLN(BLN115),.WL(WL91));
sram_cell_6t_5 inst_cell_91_116 (.BL(BL116),.BLN(BLN116),.WL(WL91));
sram_cell_6t_5 inst_cell_91_117 (.BL(BL117),.BLN(BLN117),.WL(WL91));
sram_cell_6t_5 inst_cell_91_118 (.BL(BL118),.BLN(BLN118),.WL(WL91));
sram_cell_6t_5 inst_cell_91_119 (.BL(BL119),.BLN(BLN119),.WL(WL91));
sram_cell_6t_5 inst_cell_91_120 (.BL(BL120),.BLN(BLN120),.WL(WL91));
sram_cell_6t_5 inst_cell_91_121 (.BL(BL121),.BLN(BLN121),.WL(WL91));
sram_cell_6t_5 inst_cell_91_122 (.BL(BL122),.BLN(BLN122),.WL(WL91));
sram_cell_6t_5 inst_cell_91_123 (.BL(BL123),.BLN(BLN123),.WL(WL91));
sram_cell_6t_5 inst_cell_91_124 (.BL(BL124),.BLN(BLN124),.WL(WL91));
sram_cell_6t_5 inst_cell_91_125 (.BL(BL125),.BLN(BLN125),.WL(WL91));
sram_cell_6t_5 inst_cell_91_126 (.BL(BL126),.BLN(BLN126),.WL(WL91));
sram_cell_6t_5 inst_cell_91_127 (.BL(BL127),.BLN(BLN127),.WL(WL91));
sram_cell_6t_5 inst_cell_92_0 (.BL(BL0),.BLN(BLN0),.WL(WL92));
sram_cell_6t_5 inst_cell_92_1 (.BL(BL1),.BLN(BLN1),.WL(WL92));
sram_cell_6t_5 inst_cell_92_2 (.BL(BL2),.BLN(BLN2),.WL(WL92));
sram_cell_6t_5 inst_cell_92_3 (.BL(BL3),.BLN(BLN3),.WL(WL92));
sram_cell_6t_5 inst_cell_92_4 (.BL(BL4),.BLN(BLN4),.WL(WL92));
sram_cell_6t_5 inst_cell_92_5 (.BL(BL5),.BLN(BLN5),.WL(WL92));
sram_cell_6t_5 inst_cell_92_6 (.BL(BL6),.BLN(BLN6),.WL(WL92));
sram_cell_6t_5 inst_cell_92_7 (.BL(BL7),.BLN(BLN7),.WL(WL92));
sram_cell_6t_5 inst_cell_92_8 (.BL(BL8),.BLN(BLN8),.WL(WL92));
sram_cell_6t_5 inst_cell_92_9 (.BL(BL9),.BLN(BLN9),.WL(WL92));
sram_cell_6t_5 inst_cell_92_10 (.BL(BL10),.BLN(BLN10),.WL(WL92));
sram_cell_6t_5 inst_cell_92_11 (.BL(BL11),.BLN(BLN11),.WL(WL92));
sram_cell_6t_5 inst_cell_92_12 (.BL(BL12),.BLN(BLN12),.WL(WL92));
sram_cell_6t_5 inst_cell_92_13 (.BL(BL13),.BLN(BLN13),.WL(WL92));
sram_cell_6t_5 inst_cell_92_14 (.BL(BL14),.BLN(BLN14),.WL(WL92));
sram_cell_6t_5 inst_cell_92_15 (.BL(BL15),.BLN(BLN15),.WL(WL92));
sram_cell_6t_5 inst_cell_92_16 (.BL(BL16),.BLN(BLN16),.WL(WL92));
sram_cell_6t_5 inst_cell_92_17 (.BL(BL17),.BLN(BLN17),.WL(WL92));
sram_cell_6t_5 inst_cell_92_18 (.BL(BL18),.BLN(BLN18),.WL(WL92));
sram_cell_6t_5 inst_cell_92_19 (.BL(BL19),.BLN(BLN19),.WL(WL92));
sram_cell_6t_5 inst_cell_92_20 (.BL(BL20),.BLN(BLN20),.WL(WL92));
sram_cell_6t_5 inst_cell_92_21 (.BL(BL21),.BLN(BLN21),.WL(WL92));
sram_cell_6t_5 inst_cell_92_22 (.BL(BL22),.BLN(BLN22),.WL(WL92));
sram_cell_6t_5 inst_cell_92_23 (.BL(BL23),.BLN(BLN23),.WL(WL92));
sram_cell_6t_5 inst_cell_92_24 (.BL(BL24),.BLN(BLN24),.WL(WL92));
sram_cell_6t_5 inst_cell_92_25 (.BL(BL25),.BLN(BLN25),.WL(WL92));
sram_cell_6t_5 inst_cell_92_26 (.BL(BL26),.BLN(BLN26),.WL(WL92));
sram_cell_6t_5 inst_cell_92_27 (.BL(BL27),.BLN(BLN27),.WL(WL92));
sram_cell_6t_5 inst_cell_92_28 (.BL(BL28),.BLN(BLN28),.WL(WL92));
sram_cell_6t_5 inst_cell_92_29 (.BL(BL29),.BLN(BLN29),.WL(WL92));
sram_cell_6t_5 inst_cell_92_30 (.BL(BL30),.BLN(BLN30),.WL(WL92));
sram_cell_6t_5 inst_cell_92_31 (.BL(BL31),.BLN(BLN31),.WL(WL92));
sram_cell_6t_5 inst_cell_92_32 (.BL(BL32),.BLN(BLN32),.WL(WL92));
sram_cell_6t_5 inst_cell_92_33 (.BL(BL33),.BLN(BLN33),.WL(WL92));
sram_cell_6t_5 inst_cell_92_34 (.BL(BL34),.BLN(BLN34),.WL(WL92));
sram_cell_6t_5 inst_cell_92_35 (.BL(BL35),.BLN(BLN35),.WL(WL92));
sram_cell_6t_5 inst_cell_92_36 (.BL(BL36),.BLN(BLN36),.WL(WL92));
sram_cell_6t_5 inst_cell_92_37 (.BL(BL37),.BLN(BLN37),.WL(WL92));
sram_cell_6t_5 inst_cell_92_38 (.BL(BL38),.BLN(BLN38),.WL(WL92));
sram_cell_6t_5 inst_cell_92_39 (.BL(BL39),.BLN(BLN39),.WL(WL92));
sram_cell_6t_5 inst_cell_92_40 (.BL(BL40),.BLN(BLN40),.WL(WL92));
sram_cell_6t_5 inst_cell_92_41 (.BL(BL41),.BLN(BLN41),.WL(WL92));
sram_cell_6t_5 inst_cell_92_42 (.BL(BL42),.BLN(BLN42),.WL(WL92));
sram_cell_6t_5 inst_cell_92_43 (.BL(BL43),.BLN(BLN43),.WL(WL92));
sram_cell_6t_5 inst_cell_92_44 (.BL(BL44),.BLN(BLN44),.WL(WL92));
sram_cell_6t_5 inst_cell_92_45 (.BL(BL45),.BLN(BLN45),.WL(WL92));
sram_cell_6t_5 inst_cell_92_46 (.BL(BL46),.BLN(BLN46),.WL(WL92));
sram_cell_6t_5 inst_cell_92_47 (.BL(BL47),.BLN(BLN47),.WL(WL92));
sram_cell_6t_5 inst_cell_92_48 (.BL(BL48),.BLN(BLN48),.WL(WL92));
sram_cell_6t_5 inst_cell_92_49 (.BL(BL49),.BLN(BLN49),.WL(WL92));
sram_cell_6t_5 inst_cell_92_50 (.BL(BL50),.BLN(BLN50),.WL(WL92));
sram_cell_6t_5 inst_cell_92_51 (.BL(BL51),.BLN(BLN51),.WL(WL92));
sram_cell_6t_5 inst_cell_92_52 (.BL(BL52),.BLN(BLN52),.WL(WL92));
sram_cell_6t_5 inst_cell_92_53 (.BL(BL53),.BLN(BLN53),.WL(WL92));
sram_cell_6t_5 inst_cell_92_54 (.BL(BL54),.BLN(BLN54),.WL(WL92));
sram_cell_6t_5 inst_cell_92_55 (.BL(BL55),.BLN(BLN55),.WL(WL92));
sram_cell_6t_5 inst_cell_92_56 (.BL(BL56),.BLN(BLN56),.WL(WL92));
sram_cell_6t_5 inst_cell_92_57 (.BL(BL57),.BLN(BLN57),.WL(WL92));
sram_cell_6t_5 inst_cell_92_58 (.BL(BL58),.BLN(BLN58),.WL(WL92));
sram_cell_6t_5 inst_cell_92_59 (.BL(BL59),.BLN(BLN59),.WL(WL92));
sram_cell_6t_5 inst_cell_92_60 (.BL(BL60),.BLN(BLN60),.WL(WL92));
sram_cell_6t_5 inst_cell_92_61 (.BL(BL61),.BLN(BLN61),.WL(WL92));
sram_cell_6t_5 inst_cell_92_62 (.BL(BL62),.BLN(BLN62),.WL(WL92));
sram_cell_6t_5 inst_cell_92_63 (.BL(BL63),.BLN(BLN63),.WL(WL92));
sram_cell_6t_5 inst_cell_92_64 (.BL(BL64),.BLN(BLN64),.WL(WL92));
sram_cell_6t_5 inst_cell_92_65 (.BL(BL65),.BLN(BLN65),.WL(WL92));
sram_cell_6t_5 inst_cell_92_66 (.BL(BL66),.BLN(BLN66),.WL(WL92));
sram_cell_6t_5 inst_cell_92_67 (.BL(BL67),.BLN(BLN67),.WL(WL92));
sram_cell_6t_5 inst_cell_92_68 (.BL(BL68),.BLN(BLN68),.WL(WL92));
sram_cell_6t_5 inst_cell_92_69 (.BL(BL69),.BLN(BLN69),.WL(WL92));
sram_cell_6t_5 inst_cell_92_70 (.BL(BL70),.BLN(BLN70),.WL(WL92));
sram_cell_6t_5 inst_cell_92_71 (.BL(BL71),.BLN(BLN71),.WL(WL92));
sram_cell_6t_5 inst_cell_92_72 (.BL(BL72),.BLN(BLN72),.WL(WL92));
sram_cell_6t_5 inst_cell_92_73 (.BL(BL73),.BLN(BLN73),.WL(WL92));
sram_cell_6t_5 inst_cell_92_74 (.BL(BL74),.BLN(BLN74),.WL(WL92));
sram_cell_6t_5 inst_cell_92_75 (.BL(BL75),.BLN(BLN75),.WL(WL92));
sram_cell_6t_5 inst_cell_92_76 (.BL(BL76),.BLN(BLN76),.WL(WL92));
sram_cell_6t_5 inst_cell_92_77 (.BL(BL77),.BLN(BLN77),.WL(WL92));
sram_cell_6t_5 inst_cell_92_78 (.BL(BL78),.BLN(BLN78),.WL(WL92));
sram_cell_6t_5 inst_cell_92_79 (.BL(BL79),.BLN(BLN79),.WL(WL92));
sram_cell_6t_5 inst_cell_92_80 (.BL(BL80),.BLN(BLN80),.WL(WL92));
sram_cell_6t_5 inst_cell_92_81 (.BL(BL81),.BLN(BLN81),.WL(WL92));
sram_cell_6t_5 inst_cell_92_82 (.BL(BL82),.BLN(BLN82),.WL(WL92));
sram_cell_6t_5 inst_cell_92_83 (.BL(BL83),.BLN(BLN83),.WL(WL92));
sram_cell_6t_5 inst_cell_92_84 (.BL(BL84),.BLN(BLN84),.WL(WL92));
sram_cell_6t_5 inst_cell_92_85 (.BL(BL85),.BLN(BLN85),.WL(WL92));
sram_cell_6t_5 inst_cell_92_86 (.BL(BL86),.BLN(BLN86),.WL(WL92));
sram_cell_6t_5 inst_cell_92_87 (.BL(BL87),.BLN(BLN87),.WL(WL92));
sram_cell_6t_5 inst_cell_92_88 (.BL(BL88),.BLN(BLN88),.WL(WL92));
sram_cell_6t_5 inst_cell_92_89 (.BL(BL89),.BLN(BLN89),.WL(WL92));
sram_cell_6t_5 inst_cell_92_90 (.BL(BL90),.BLN(BLN90),.WL(WL92));
sram_cell_6t_5 inst_cell_92_91 (.BL(BL91),.BLN(BLN91),.WL(WL92));
sram_cell_6t_5 inst_cell_92_92 (.BL(BL92),.BLN(BLN92),.WL(WL92));
sram_cell_6t_5 inst_cell_92_93 (.BL(BL93),.BLN(BLN93),.WL(WL92));
sram_cell_6t_5 inst_cell_92_94 (.BL(BL94),.BLN(BLN94),.WL(WL92));
sram_cell_6t_5 inst_cell_92_95 (.BL(BL95),.BLN(BLN95),.WL(WL92));
sram_cell_6t_5 inst_cell_92_96 (.BL(BL96),.BLN(BLN96),.WL(WL92));
sram_cell_6t_5 inst_cell_92_97 (.BL(BL97),.BLN(BLN97),.WL(WL92));
sram_cell_6t_5 inst_cell_92_98 (.BL(BL98),.BLN(BLN98),.WL(WL92));
sram_cell_6t_5 inst_cell_92_99 (.BL(BL99),.BLN(BLN99),.WL(WL92));
sram_cell_6t_5 inst_cell_92_100 (.BL(BL100),.BLN(BLN100),.WL(WL92));
sram_cell_6t_5 inst_cell_92_101 (.BL(BL101),.BLN(BLN101),.WL(WL92));
sram_cell_6t_5 inst_cell_92_102 (.BL(BL102),.BLN(BLN102),.WL(WL92));
sram_cell_6t_5 inst_cell_92_103 (.BL(BL103),.BLN(BLN103),.WL(WL92));
sram_cell_6t_5 inst_cell_92_104 (.BL(BL104),.BLN(BLN104),.WL(WL92));
sram_cell_6t_5 inst_cell_92_105 (.BL(BL105),.BLN(BLN105),.WL(WL92));
sram_cell_6t_5 inst_cell_92_106 (.BL(BL106),.BLN(BLN106),.WL(WL92));
sram_cell_6t_5 inst_cell_92_107 (.BL(BL107),.BLN(BLN107),.WL(WL92));
sram_cell_6t_5 inst_cell_92_108 (.BL(BL108),.BLN(BLN108),.WL(WL92));
sram_cell_6t_5 inst_cell_92_109 (.BL(BL109),.BLN(BLN109),.WL(WL92));
sram_cell_6t_5 inst_cell_92_110 (.BL(BL110),.BLN(BLN110),.WL(WL92));
sram_cell_6t_5 inst_cell_92_111 (.BL(BL111),.BLN(BLN111),.WL(WL92));
sram_cell_6t_5 inst_cell_92_112 (.BL(BL112),.BLN(BLN112),.WL(WL92));
sram_cell_6t_5 inst_cell_92_113 (.BL(BL113),.BLN(BLN113),.WL(WL92));
sram_cell_6t_5 inst_cell_92_114 (.BL(BL114),.BLN(BLN114),.WL(WL92));
sram_cell_6t_5 inst_cell_92_115 (.BL(BL115),.BLN(BLN115),.WL(WL92));
sram_cell_6t_5 inst_cell_92_116 (.BL(BL116),.BLN(BLN116),.WL(WL92));
sram_cell_6t_5 inst_cell_92_117 (.BL(BL117),.BLN(BLN117),.WL(WL92));
sram_cell_6t_5 inst_cell_92_118 (.BL(BL118),.BLN(BLN118),.WL(WL92));
sram_cell_6t_5 inst_cell_92_119 (.BL(BL119),.BLN(BLN119),.WL(WL92));
sram_cell_6t_5 inst_cell_92_120 (.BL(BL120),.BLN(BLN120),.WL(WL92));
sram_cell_6t_5 inst_cell_92_121 (.BL(BL121),.BLN(BLN121),.WL(WL92));
sram_cell_6t_5 inst_cell_92_122 (.BL(BL122),.BLN(BLN122),.WL(WL92));
sram_cell_6t_5 inst_cell_92_123 (.BL(BL123),.BLN(BLN123),.WL(WL92));
sram_cell_6t_5 inst_cell_92_124 (.BL(BL124),.BLN(BLN124),.WL(WL92));
sram_cell_6t_5 inst_cell_92_125 (.BL(BL125),.BLN(BLN125),.WL(WL92));
sram_cell_6t_5 inst_cell_92_126 (.BL(BL126),.BLN(BLN126),.WL(WL92));
sram_cell_6t_5 inst_cell_92_127 (.BL(BL127),.BLN(BLN127),.WL(WL92));
sram_cell_6t_5 inst_cell_93_0 (.BL(BL0),.BLN(BLN0),.WL(WL93));
sram_cell_6t_5 inst_cell_93_1 (.BL(BL1),.BLN(BLN1),.WL(WL93));
sram_cell_6t_5 inst_cell_93_2 (.BL(BL2),.BLN(BLN2),.WL(WL93));
sram_cell_6t_5 inst_cell_93_3 (.BL(BL3),.BLN(BLN3),.WL(WL93));
sram_cell_6t_5 inst_cell_93_4 (.BL(BL4),.BLN(BLN4),.WL(WL93));
sram_cell_6t_5 inst_cell_93_5 (.BL(BL5),.BLN(BLN5),.WL(WL93));
sram_cell_6t_5 inst_cell_93_6 (.BL(BL6),.BLN(BLN6),.WL(WL93));
sram_cell_6t_5 inst_cell_93_7 (.BL(BL7),.BLN(BLN7),.WL(WL93));
sram_cell_6t_5 inst_cell_93_8 (.BL(BL8),.BLN(BLN8),.WL(WL93));
sram_cell_6t_5 inst_cell_93_9 (.BL(BL9),.BLN(BLN9),.WL(WL93));
sram_cell_6t_5 inst_cell_93_10 (.BL(BL10),.BLN(BLN10),.WL(WL93));
sram_cell_6t_5 inst_cell_93_11 (.BL(BL11),.BLN(BLN11),.WL(WL93));
sram_cell_6t_5 inst_cell_93_12 (.BL(BL12),.BLN(BLN12),.WL(WL93));
sram_cell_6t_5 inst_cell_93_13 (.BL(BL13),.BLN(BLN13),.WL(WL93));
sram_cell_6t_5 inst_cell_93_14 (.BL(BL14),.BLN(BLN14),.WL(WL93));
sram_cell_6t_5 inst_cell_93_15 (.BL(BL15),.BLN(BLN15),.WL(WL93));
sram_cell_6t_5 inst_cell_93_16 (.BL(BL16),.BLN(BLN16),.WL(WL93));
sram_cell_6t_5 inst_cell_93_17 (.BL(BL17),.BLN(BLN17),.WL(WL93));
sram_cell_6t_5 inst_cell_93_18 (.BL(BL18),.BLN(BLN18),.WL(WL93));
sram_cell_6t_5 inst_cell_93_19 (.BL(BL19),.BLN(BLN19),.WL(WL93));
sram_cell_6t_5 inst_cell_93_20 (.BL(BL20),.BLN(BLN20),.WL(WL93));
sram_cell_6t_5 inst_cell_93_21 (.BL(BL21),.BLN(BLN21),.WL(WL93));
sram_cell_6t_5 inst_cell_93_22 (.BL(BL22),.BLN(BLN22),.WL(WL93));
sram_cell_6t_5 inst_cell_93_23 (.BL(BL23),.BLN(BLN23),.WL(WL93));
sram_cell_6t_5 inst_cell_93_24 (.BL(BL24),.BLN(BLN24),.WL(WL93));
sram_cell_6t_5 inst_cell_93_25 (.BL(BL25),.BLN(BLN25),.WL(WL93));
sram_cell_6t_5 inst_cell_93_26 (.BL(BL26),.BLN(BLN26),.WL(WL93));
sram_cell_6t_5 inst_cell_93_27 (.BL(BL27),.BLN(BLN27),.WL(WL93));
sram_cell_6t_5 inst_cell_93_28 (.BL(BL28),.BLN(BLN28),.WL(WL93));
sram_cell_6t_5 inst_cell_93_29 (.BL(BL29),.BLN(BLN29),.WL(WL93));
sram_cell_6t_5 inst_cell_93_30 (.BL(BL30),.BLN(BLN30),.WL(WL93));
sram_cell_6t_5 inst_cell_93_31 (.BL(BL31),.BLN(BLN31),.WL(WL93));
sram_cell_6t_5 inst_cell_93_32 (.BL(BL32),.BLN(BLN32),.WL(WL93));
sram_cell_6t_5 inst_cell_93_33 (.BL(BL33),.BLN(BLN33),.WL(WL93));
sram_cell_6t_5 inst_cell_93_34 (.BL(BL34),.BLN(BLN34),.WL(WL93));
sram_cell_6t_5 inst_cell_93_35 (.BL(BL35),.BLN(BLN35),.WL(WL93));
sram_cell_6t_5 inst_cell_93_36 (.BL(BL36),.BLN(BLN36),.WL(WL93));
sram_cell_6t_5 inst_cell_93_37 (.BL(BL37),.BLN(BLN37),.WL(WL93));
sram_cell_6t_5 inst_cell_93_38 (.BL(BL38),.BLN(BLN38),.WL(WL93));
sram_cell_6t_5 inst_cell_93_39 (.BL(BL39),.BLN(BLN39),.WL(WL93));
sram_cell_6t_5 inst_cell_93_40 (.BL(BL40),.BLN(BLN40),.WL(WL93));
sram_cell_6t_5 inst_cell_93_41 (.BL(BL41),.BLN(BLN41),.WL(WL93));
sram_cell_6t_5 inst_cell_93_42 (.BL(BL42),.BLN(BLN42),.WL(WL93));
sram_cell_6t_5 inst_cell_93_43 (.BL(BL43),.BLN(BLN43),.WL(WL93));
sram_cell_6t_5 inst_cell_93_44 (.BL(BL44),.BLN(BLN44),.WL(WL93));
sram_cell_6t_5 inst_cell_93_45 (.BL(BL45),.BLN(BLN45),.WL(WL93));
sram_cell_6t_5 inst_cell_93_46 (.BL(BL46),.BLN(BLN46),.WL(WL93));
sram_cell_6t_5 inst_cell_93_47 (.BL(BL47),.BLN(BLN47),.WL(WL93));
sram_cell_6t_5 inst_cell_93_48 (.BL(BL48),.BLN(BLN48),.WL(WL93));
sram_cell_6t_5 inst_cell_93_49 (.BL(BL49),.BLN(BLN49),.WL(WL93));
sram_cell_6t_5 inst_cell_93_50 (.BL(BL50),.BLN(BLN50),.WL(WL93));
sram_cell_6t_5 inst_cell_93_51 (.BL(BL51),.BLN(BLN51),.WL(WL93));
sram_cell_6t_5 inst_cell_93_52 (.BL(BL52),.BLN(BLN52),.WL(WL93));
sram_cell_6t_5 inst_cell_93_53 (.BL(BL53),.BLN(BLN53),.WL(WL93));
sram_cell_6t_5 inst_cell_93_54 (.BL(BL54),.BLN(BLN54),.WL(WL93));
sram_cell_6t_5 inst_cell_93_55 (.BL(BL55),.BLN(BLN55),.WL(WL93));
sram_cell_6t_5 inst_cell_93_56 (.BL(BL56),.BLN(BLN56),.WL(WL93));
sram_cell_6t_5 inst_cell_93_57 (.BL(BL57),.BLN(BLN57),.WL(WL93));
sram_cell_6t_5 inst_cell_93_58 (.BL(BL58),.BLN(BLN58),.WL(WL93));
sram_cell_6t_5 inst_cell_93_59 (.BL(BL59),.BLN(BLN59),.WL(WL93));
sram_cell_6t_5 inst_cell_93_60 (.BL(BL60),.BLN(BLN60),.WL(WL93));
sram_cell_6t_5 inst_cell_93_61 (.BL(BL61),.BLN(BLN61),.WL(WL93));
sram_cell_6t_5 inst_cell_93_62 (.BL(BL62),.BLN(BLN62),.WL(WL93));
sram_cell_6t_5 inst_cell_93_63 (.BL(BL63),.BLN(BLN63),.WL(WL93));
sram_cell_6t_5 inst_cell_93_64 (.BL(BL64),.BLN(BLN64),.WL(WL93));
sram_cell_6t_5 inst_cell_93_65 (.BL(BL65),.BLN(BLN65),.WL(WL93));
sram_cell_6t_5 inst_cell_93_66 (.BL(BL66),.BLN(BLN66),.WL(WL93));
sram_cell_6t_5 inst_cell_93_67 (.BL(BL67),.BLN(BLN67),.WL(WL93));
sram_cell_6t_5 inst_cell_93_68 (.BL(BL68),.BLN(BLN68),.WL(WL93));
sram_cell_6t_5 inst_cell_93_69 (.BL(BL69),.BLN(BLN69),.WL(WL93));
sram_cell_6t_5 inst_cell_93_70 (.BL(BL70),.BLN(BLN70),.WL(WL93));
sram_cell_6t_5 inst_cell_93_71 (.BL(BL71),.BLN(BLN71),.WL(WL93));
sram_cell_6t_5 inst_cell_93_72 (.BL(BL72),.BLN(BLN72),.WL(WL93));
sram_cell_6t_5 inst_cell_93_73 (.BL(BL73),.BLN(BLN73),.WL(WL93));
sram_cell_6t_5 inst_cell_93_74 (.BL(BL74),.BLN(BLN74),.WL(WL93));
sram_cell_6t_5 inst_cell_93_75 (.BL(BL75),.BLN(BLN75),.WL(WL93));
sram_cell_6t_5 inst_cell_93_76 (.BL(BL76),.BLN(BLN76),.WL(WL93));
sram_cell_6t_5 inst_cell_93_77 (.BL(BL77),.BLN(BLN77),.WL(WL93));
sram_cell_6t_5 inst_cell_93_78 (.BL(BL78),.BLN(BLN78),.WL(WL93));
sram_cell_6t_5 inst_cell_93_79 (.BL(BL79),.BLN(BLN79),.WL(WL93));
sram_cell_6t_5 inst_cell_93_80 (.BL(BL80),.BLN(BLN80),.WL(WL93));
sram_cell_6t_5 inst_cell_93_81 (.BL(BL81),.BLN(BLN81),.WL(WL93));
sram_cell_6t_5 inst_cell_93_82 (.BL(BL82),.BLN(BLN82),.WL(WL93));
sram_cell_6t_5 inst_cell_93_83 (.BL(BL83),.BLN(BLN83),.WL(WL93));
sram_cell_6t_5 inst_cell_93_84 (.BL(BL84),.BLN(BLN84),.WL(WL93));
sram_cell_6t_5 inst_cell_93_85 (.BL(BL85),.BLN(BLN85),.WL(WL93));
sram_cell_6t_5 inst_cell_93_86 (.BL(BL86),.BLN(BLN86),.WL(WL93));
sram_cell_6t_5 inst_cell_93_87 (.BL(BL87),.BLN(BLN87),.WL(WL93));
sram_cell_6t_5 inst_cell_93_88 (.BL(BL88),.BLN(BLN88),.WL(WL93));
sram_cell_6t_5 inst_cell_93_89 (.BL(BL89),.BLN(BLN89),.WL(WL93));
sram_cell_6t_5 inst_cell_93_90 (.BL(BL90),.BLN(BLN90),.WL(WL93));
sram_cell_6t_5 inst_cell_93_91 (.BL(BL91),.BLN(BLN91),.WL(WL93));
sram_cell_6t_5 inst_cell_93_92 (.BL(BL92),.BLN(BLN92),.WL(WL93));
sram_cell_6t_5 inst_cell_93_93 (.BL(BL93),.BLN(BLN93),.WL(WL93));
sram_cell_6t_5 inst_cell_93_94 (.BL(BL94),.BLN(BLN94),.WL(WL93));
sram_cell_6t_5 inst_cell_93_95 (.BL(BL95),.BLN(BLN95),.WL(WL93));
sram_cell_6t_5 inst_cell_93_96 (.BL(BL96),.BLN(BLN96),.WL(WL93));
sram_cell_6t_5 inst_cell_93_97 (.BL(BL97),.BLN(BLN97),.WL(WL93));
sram_cell_6t_5 inst_cell_93_98 (.BL(BL98),.BLN(BLN98),.WL(WL93));
sram_cell_6t_5 inst_cell_93_99 (.BL(BL99),.BLN(BLN99),.WL(WL93));
sram_cell_6t_5 inst_cell_93_100 (.BL(BL100),.BLN(BLN100),.WL(WL93));
sram_cell_6t_5 inst_cell_93_101 (.BL(BL101),.BLN(BLN101),.WL(WL93));
sram_cell_6t_5 inst_cell_93_102 (.BL(BL102),.BLN(BLN102),.WL(WL93));
sram_cell_6t_5 inst_cell_93_103 (.BL(BL103),.BLN(BLN103),.WL(WL93));
sram_cell_6t_5 inst_cell_93_104 (.BL(BL104),.BLN(BLN104),.WL(WL93));
sram_cell_6t_5 inst_cell_93_105 (.BL(BL105),.BLN(BLN105),.WL(WL93));
sram_cell_6t_5 inst_cell_93_106 (.BL(BL106),.BLN(BLN106),.WL(WL93));
sram_cell_6t_5 inst_cell_93_107 (.BL(BL107),.BLN(BLN107),.WL(WL93));
sram_cell_6t_5 inst_cell_93_108 (.BL(BL108),.BLN(BLN108),.WL(WL93));
sram_cell_6t_5 inst_cell_93_109 (.BL(BL109),.BLN(BLN109),.WL(WL93));
sram_cell_6t_5 inst_cell_93_110 (.BL(BL110),.BLN(BLN110),.WL(WL93));
sram_cell_6t_5 inst_cell_93_111 (.BL(BL111),.BLN(BLN111),.WL(WL93));
sram_cell_6t_5 inst_cell_93_112 (.BL(BL112),.BLN(BLN112),.WL(WL93));
sram_cell_6t_5 inst_cell_93_113 (.BL(BL113),.BLN(BLN113),.WL(WL93));
sram_cell_6t_5 inst_cell_93_114 (.BL(BL114),.BLN(BLN114),.WL(WL93));
sram_cell_6t_5 inst_cell_93_115 (.BL(BL115),.BLN(BLN115),.WL(WL93));
sram_cell_6t_5 inst_cell_93_116 (.BL(BL116),.BLN(BLN116),.WL(WL93));
sram_cell_6t_5 inst_cell_93_117 (.BL(BL117),.BLN(BLN117),.WL(WL93));
sram_cell_6t_5 inst_cell_93_118 (.BL(BL118),.BLN(BLN118),.WL(WL93));
sram_cell_6t_5 inst_cell_93_119 (.BL(BL119),.BLN(BLN119),.WL(WL93));
sram_cell_6t_5 inst_cell_93_120 (.BL(BL120),.BLN(BLN120),.WL(WL93));
sram_cell_6t_5 inst_cell_93_121 (.BL(BL121),.BLN(BLN121),.WL(WL93));
sram_cell_6t_5 inst_cell_93_122 (.BL(BL122),.BLN(BLN122),.WL(WL93));
sram_cell_6t_5 inst_cell_93_123 (.BL(BL123),.BLN(BLN123),.WL(WL93));
sram_cell_6t_5 inst_cell_93_124 (.BL(BL124),.BLN(BLN124),.WL(WL93));
sram_cell_6t_5 inst_cell_93_125 (.BL(BL125),.BLN(BLN125),.WL(WL93));
sram_cell_6t_5 inst_cell_93_126 (.BL(BL126),.BLN(BLN126),.WL(WL93));
sram_cell_6t_5 inst_cell_93_127 (.BL(BL127),.BLN(BLN127),.WL(WL93));
sram_cell_6t_5 inst_cell_94_0 (.BL(BL0),.BLN(BLN0),.WL(WL94));
sram_cell_6t_5 inst_cell_94_1 (.BL(BL1),.BLN(BLN1),.WL(WL94));
sram_cell_6t_5 inst_cell_94_2 (.BL(BL2),.BLN(BLN2),.WL(WL94));
sram_cell_6t_5 inst_cell_94_3 (.BL(BL3),.BLN(BLN3),.WL(WL94));
sram_cell_6t_5 inst_cell_94_4 (.BL(BL4),.BLN(BLN4),.WL(WL94));
sram_cell_6t_5 inst_cell_94_5 (.BL(BL5),.BLN(BLN5),.WL(WL94));
sram_cell_6t_5 inst_cell_94_6 (.BL(BL6),.BLN(BLN6),.WL(WL94));
sram_cell_6t_5 inst_cell_94_7 (.BL(BL7),.BLN(BLN7),.WL(WL94));
sram_cell_6t_5 inst_cell_94_8 (.BL(BL8),.BLN(BLN8),.WL(WL94));
sram_cell_6t_5 inst_cell_94_9 (.BL(BL9),.BLN(BLN9),.WL(WL94));
sram_cell_6t_5 inst_cell_94_10 (.BL(BL10),.BLN(BLN10),.WL(WL94));
sram_cell_6t_5 inst_cell_94_11 (.BL(BL11),.BLN(BLN11),.WL(WL94));
sram_cell_6t_5 inst_cell_94_12 (.BL(BL12),.BLN(BLN12),.WL(WL94));
sram_cell_6t_5 inst_cell_94_13 (.BL(BL13),.BLN(BLN13),.WL(WL94));
sram_cell_6t_5 inst_cell_94_14 (.BL(BL14),.BLN(BLN14),.WL(WL94));
sram_cell_6t_5 inst_cell_94_15 (.BL(BL15),.BLN(BLN15),.WL(WL94));
sram_cell_6t_5 inst_cell_94_16 (.BL(BL16),.BLN(BLN16),.WL(WL94));
sram_cell_6t_5 inst_cell_94_17 (.BL(BL17),.BLN(BLN17),.WL(WL94));
sram_cell_6t_5 inst_cell_94_18 (.BL(BL18),.BLN(BLN18),.WL(WL94));
sram_cell_6t_5 inst_cell_94_19 (.BL(BL19),.BLN(BLN19),.WL(WL94));
sram_cell_6t_5 inst_cell_94_20 (.BL(BL20),.BLN(BLN20),.WL(WL94));
sram_cell_6t_5 inst_cell_94_21 (.BL(BL21),.BLN(BLN21),.WL(WL94));
sram_cell_6t_5 inst_cell_94_22 (.BL(BL22),.BLN(BLN22),.WL(WL94));
sram_cell_6t_5 inst_cell_94_23 (.BL(BL23),.BLN(BLN23),.WL(WL94));
sram_cell_6t_5 inst_cell_94_24 (.BL(BL24),.BLN(BLN24),.WL(WL94));
sram_cell_6t_5 inst_cell_94_25 (.BL(BL25),.BLN(BLN25),.WL(WL94));
sram_cell_6t_5 inst_cell_94_26 (.BL(BL26),.BLN(BLN26),.WL(WL94));
sram_cell_6t_5 inst_cell_94_27 (.BL(BL27),.BLN(BLN27),.WL(WL94));
sram_cell_6t_5 inst_cell_94_28 (.BL(BL28),.BLN(BLN28),.WL(WL94));
sram_cell_6t_5 inst_cell_94_29 (.BL(BL29),.BLN(BLN29),.WL(WL94));
sram_cell_6t_5 inst_cell_94_30 (.BL(BL30),.BLN(BLN30),.WL(WL94));
sram_cell_6t_5 inst_cell_94_31 (.BL(BL31),.BLN(BLN31),.WL(WL94));
sram_cell_6t_5 inst_cell_94_32 (.BL(BL32),.BLN(BLN32),.WL(WL94));
sram_cell_6t_5 inst_cell_94_33 (.BL(BL33),.BLN(BLN33),.WL(WL94));
sram_cell_6t_5 inst_cell_94_34 (.BL(BL34),.BLN(BLN34),.WL(WL94));
sram_cell_6t_5 inst_cell_94_35 (.BL(BL35),.BLN(BLN35),.WL(WL94));
sram_cell_6t_5 inst_cell_94_36 (.BL(BL36),.BLN(BLN36),.WL(WL94));
sram_cell_6t_5 inst_cell_94_37 (.BL(BL37),.BLN(BLN37),.WL(WL94));
sram_cell_6t_5 inst_cell_94_38 (.BL(BL38),.BLN(BLN38),.WL(WL94));
sram_cell_6t_5 inst_cell_94_39 (.BL(BL39),.BLN(BLN39),.WL(WL94));
sram_cell_6t_5 inst_cell_94_40 (.BL(BL40),.BLN(BLN40),.WL(WL94));
sram_cell_6t_5 inst_cell_94_41 (.BL(BL41),.BLN(BLN41),.WL(WL94));
sram_cell_6t_5 inst_cell_94_42 (.BL(BL42),.BLN(BLN42),.WL(WL94));
sram_cell_6t_5 inst_cell_94_43 (.BL(BL43),.BLN(BLN43),.WL(WL94));
sram_cell_6t_5 inst_cell_94_44 (.BL(BL44),.BLN(BLN44),.WL(WL94));
sram_cell_6t_5 inst_cell_94_45 (.BL(BL45),.BLN(BLN45),.WL(WL94));
sram_cell_6t_5 inst_cell_94_46 (.BL(BL46),.BLN(BLN46),.WL(WL94));
sram_cell_6t_5 inst_cell_94_47 (.BL(BL47),.BLN(BLN47),.WL(WL94));
sram_cell_6t_5 inst_cell_94_48 (.BL(BL48),.BLN(BLN48),.WL(WL94));
sram_cell_6t_5 inst_cell_94_49 (.BL(BL49),.BLN(BLN49),.WL(WL94));
sram_cell_6t_5 inst_cell_94_50 (.BL(BL50),.BLN(BLN50),.WL(WL94));
sram_cell_6t_5 inst_cell_94_51 (.BL(BL51),.BLN(BLN51),.WL(WL94));
sram_cell_6t_5 inst_cell_94_52 (.BL(BL52),.BLN(BLN52),.WL(WL94));
sram_cell_6t_5 inst_cell_94_53 (.BL(BL53),.BLN(BLN53),.WL(WL94));
sram_cell_6t_5 inst_cell_94_54 (.BL(BL54),.BLN(BLN54),.WL(WL94));
sram_cell_6t_5 inst_cell_94_55 (.BL(BL55),.BLN(BLN55),.WL(WL94));
sram_cell_6t_5 inst_cell_94_56 (.BL(BL56),.BLN(BLN56),.WL(WL94));
sram_cell_6t_5 inst_cell_94_57 (.BL(BL57),.BLN(BLN57),.WL(WL94));
sram_cell_6t_5 inst_cell_94_58 (.BL(BL58),.BLN(BLN58),.WL(WL94));
sram_cell_6t_5 inst_cell_94_59 (.BL(BL59),.BLN(BLN59),.WL(WL94));
sram_cell_6t_5 inst_cell_94_60 (.BL(BL60),.BLN(BLN60),.WL(WL94));
sram_cell_6t_5 inst_cell_94_61 (.BL(BL61),.BLN(BLN61),.WL(WL94));
sram_cell_6t_5 inst_cell_94_62 (.BL(BL62),.BLN(BLN62),.WL(WL94));
sram_cell_6t_5 inst_cell_94_63 (.BL(BL63),.BLN(BLN63),.WL(WL94));
sram_cell_6t_5 inst_cell_94_64 (.BL(BL64),.BLN(BLN64),.WL(WL94));
sram_cell_6t_5 inst_cell_94_65 (.BL(BL65),.BLN(BLN65),.WL(WL94));
sram_cell_6t_5 inst_cell_94_66 (.BL(BL66),.BLN(BLN66),.WL(WL94));
sram_cell_6t_5 inst_cell_94_67 (.BL(BL67),.BLN(BLN67),.WL(WL94));
sram_cell_6t_5 inst_cell_94_68 (.BL(BL68),.BLN(BLN68),.WL(WL94));
sram_cell_6t_5 inst_cell_94_69 (.BL(BL69),.BLN(BLN69),.WL(WL94));
sram_cell_6t_5 inst_cell_94_70 (.BL(BL70),.BLN(BLN70),.WL(WL94));
sram_cell_6t_5 inst_cell_94_71 (.BL(BL71),.BLN(BLN71),.WL(WL94));
sram_cell_6t_5 inst_cell_94_72 (.BL(BL72),.BLN(BLN72),.WL(WL94));
sram_cell_6t_5 inst_cell_94_73 (.BL(BL73),.BLN(BLN73),.WL(WL94));
sram_cell_6t_5 inst_cell_94_74 (.BL(BL74),.BLN(BLN74),.WL(WL94));
sram_cell_6t_5 inst_cell_94_75 (.BL(BL75),.BLN(BLN75),.WL(WL94));
sram_cell_6t_5 inst_cell_94_76 (.BL(BL76),.BLN(BLN76),.WL(WL94));
sram_cell_6t_5 inst_cell_94_77 (.BL(BL77),.BLN(BLN77),.WL(WL94));
sram_cell_6t_5 inst_cell_94_78 (.BL(BL78),.BLN(BLN78),.WL(WL94));
sram_cell_6t_5 inst_cell_94_79 (.BL(BL79),.BLN(BLN79),.WL(WL94));
sram_cell_6t_5 inst_cell_94_80 (.BL(BL80),.BLN(BLN80),.WL(WL94));
sram_cell_6t_5 inst_cell_94_81 (.BL(BL81),.BLN(BLN81),.WL(WL94));
sram_cell_6t_5 inst_cell_94_82 (.BL(BL82),.BLN(BLN82),.WL(WL94));
sram_cell_6t_5 inst_cell_94_83 (.BL(BL83),.BLN(BLN83),.WL(WL94));
sram_cell_6t_5 inst_cell_94_84 (.BL(BL84),.BLN(BLN84),.WL(WL94));
sram_cell_6t_5 inst_cell_94_85 (.BL(BL85),.BLN(BLN85),.WL(WL94));
sram_cell_6t_5 inst_cell_94_86 (.BL(BL86),.BLN(BLN86),.WL(WL94));
sram_cell_6t_5 inst_cell_94_87 (.BL(BL87),.BLN(BLN87),.WL(WL94));
sram_cell_6t_5 inst_cell_94_88 (.BL(BL88),.BLN(BLN88),.WL(WL94));
sram_cell_6t_5 inst_cell_94_89 (.BL(BL89),.BLN(BLN89),.WL(WL94));
sram_cell_6t_5 inst_cell_94_90 (.BL(BL90),.BLN(BLN90),.WL(WL94));
sram_cell_6t_5 inst_cell_94_91 (.BL(BL91),.BLN(BLN91),.WL(WL94));
sram_cell_6t_5 inst_cell_94_92 (.BL(BL92),.BLN(BLN92),.WL(WL94));
sram_cell_6t_5 inst_cell_94_93 (.BL(BL93),.BLN(BLN93),.WL(WL94));
sram_cell_6t_5 inst_cell_94_94 (.BL(BL94),.BLN(BLN94),.WL(WL94));
sram_cell_6t_5 inst_cell_94_95 (.BL(BL95),.BLN(BLN95),.WL(WL94));
sram_cell_6t_5 inst_cell_94_96 (.BL(BL96),.BLN(BLN96),.WL(WL94));
sram_cell_6t_5 inst_cell_94_97 (.BL(BL97),.BLN(BLN97),.WL(WL94));
sram_cell_6t_5 inst_cell_94_98 (.BL(BL98),.BLN(BLN98),.WL(WL94));
sram_cell_6t_5 inst_cell_94_99 (.BL(BL99),.BLN(BLN99),.WL(WL94));
sram_cell_6t_5 inst_cell_94_100 (.BL(BL100),.BLN(BLN100),.WL(WL94));
sram_cell_6t_5 inst_cell_94_101 (.BL(BL101),.BLN(BLN101),.WL(WL94));
sram_cell_6t_5 inst_cell_94_102 (.BL(BL102),.BLN(BLN102),.WL(WL94));
sram_cell_6t_5 inst_cell_94_103 (.BL(BL103),.BLN(BLN103),.WL(WL94));
sram_cell_6t_5 inst_cell_94_104 (.BL(BL104),.BLN(BLN104),.WL(WL94));
sram_cell_6t_5 inst_cell_94_105 (.BL(BL105),.BLN(BLN105),.WL(WL94));
sram_cell_6t_5 inst_cell_94_106 (.BL(BL106),.BLN(BLN106),.WL(WL94));
sram_cell_6t_5 inst_cell_94_107 (.BL(BL107),.BLN(BLN107),.WL(WL94));
sram_cell_6t_5 inst_cell_94_108 (.BL(BL108),.BLN(BLN108),.WL(WL94));
sram_cell_6t_5 inst_cell_94_109 (.BL(BL109),.BLN(BLN109),.WL(WL94));
sram_cell_6t_5 inst_cell_94_110 (.BL(BL110),.BLN(BLN110),.WL(WL94));
sram_cell_6t_5 inst_cell_94_111 (.BL(BL111),.BLN(BLN111),.WL(WL94));
sram_cell_6t_5 inst_cell_94_112 (.BL(BL112),.BLN(BLN112),.WL(WL94));
sram_cell_6t_5 inst_cell_94_113 (.BL(BL113),.BLN(BLN113),.WL(WL94));
sram_cell_6t_5 inst_cell_94_114 (.BL(BL114),.BLN(BLN114),.WL(WL94));
sram_cell_6t_5 inst_cell_94_115 (.BL(BL115),.BLN(BLN115),.WL(WL94));
sram_cell_6t_5 inst_cell_94_116 (.BL(BL116),.BLN(BLN116),.WL(WL94));
sram_cell_6t_5 inst_cell_94_117 (.BL(BL117),.BLN(BLN117),.WL(WL94));
sram_cell_6t_5 inst_cell_94_118 (.BL(BL118),.BLN(BLN118),.WL(WL94));
sram_cell_6t_5 inst_cell_94_119 (.BL(BL119),.BLN(BLN119),.WL(WL94));
sram_cell_6t_5 inst_cell_94_120 (.BL(BL120),.BLN(BLN120),.WL(WL94));
sram_cell_6t_5 inst_cell_94_121 (.BL(BL121),.BLN(BLN121),.WL(WL94));
sram_cell_6t_5 inst_cell_94_122 (.BL(BL122),.BLN(BLN122),.WL(WL94));
sram_cell_6t_5 inst_cell_94_123 (.BL(BL123),.BLN(BLN123),.WL(WL94));
sram_cell_6t_5 inst_cell_94_124 (.BL(BL124),.BLN(BLN124),.WL(WL94));
sram_cell_6t_5 inst_cell_94_125 (.BL(BL125),.BLN(BLN125),.WL(WL94));
sram_cell_6t_5 inst_cell_94_126 (.BL(BL126),.BLN(BLN126),.WL(WL94));
sram_cell_6t_5 inst_cell_94_127 (.BL(BL127),.BLN(BLN127),.WL(WL94));
sram_cell_6t_5 inst_cell_95_0 (.BL(BL0),.BLN(BLN0),.WL(WL95));
sram_cell_6t_5 inst_cell_95_1 (.BL(BL1),.BLN(BLN1),.WL(WL95));
sram_cell_6t_5 inst_cell_95_2 (.BL(BL2),.BLN(BLN2),.WL(WL95));
sram_cell_6t_5 inst_cell_95_3 (.BL(BL3),.BLN(BLN3),.WL(WL95));
sram_cell_6t_5 inst_cell_95_4 (.BL(BL4),.BLN(BLN4),.WL(WL95));
sram_cell_6t_5 inst_cell_95_5 (.BL(BL5),.BLN(BLN5),.WL(WL95));
sram_cell_6t_5 inst_cell_95_6 (.BL(BL6),.BLN(BLN6),.WL(WL95));
sram_cell_6t_5 inst_cell_95_7 (.BL(BL7),.BLN(BLN7),.WL(WL95));
sram_cell_6t_5 inst_cell_95_8 (.BL(BL8),.BLN(BLN8),.WL(WL95));
sram_cell_6t_5 inst_cell_95_9 (.BL(BL9),.BLN(BLN9),.WL(WL95));
sram_cell_6t_5 inst_cell_95_10 (.BL(BL10),.BLN(BLN10),.WL(WL95));
sram_cell_6t_5 inst_cell_95_11 (.BL(BL11),.BLN(BLN11),.WL(WL95));
sram_cell_6t_5 inst_cell_95_12 (.BL(BL12),.BLN(BLN12),.WL(WL95));
sram_cell_6t_5 inst_cell_95_13 (.BL(BL13),.BLN(BLN13),.WL(WL95));
sram_cell_6t_5 inst_cell_95_14 (.BL(BL14),.BLN(BLN14),.WL(WL95));
sram_cell_6t_5 inst_cell_95_15 (.BL(BL15),.BLN(BLN15),.WL(WL95));
sram_cell_6t_5 inst_cell_95_16 (.BL(BL16),.BLN(BLN16),.WL(WL95));
sram_cell_6t_5 inst_cell_95_17 (.BL(BL17),.BLN(BLN17),.WL(WL95));
sram_cell_6t_5 inst_cell_95_18 (.BL(BL18),.BLN(BLN18),.WL(WL95));
sram_cell_6t_5 inst_cell_95_19 (.BL(BL19),.BLN(BLN19),.WL(WL95));
sram_cell_6t_5 inst_cell_95_20 (.BL(BL20),.BLN(BLN20),.WL(WL95));
sram_cell_6t_5 inst_cell_95_21 (.BL(BL21),.BLN(BLN21),.WL(WL95));
sram_cell_6t_5 inst_cell_95_22 (.BL(BL22),.BLN(BLN22),.WL(WL95));
sram_cell_6t_5 inst_cell_95_23 (.BL(BL23),.BLN(BLN23),.WL(WL95));
sram_cell_6t_5 inst_cell_95_24 (.BL(BL24),.BLN(BLN24),.WL(WL95));
sram_cell_6t_5 inst_cell_95_25 (.BL(BL25),.BLN(BLN25),.WL(WL95));
sram_cell_6t_5 inst_cell_95_26 (.BL(BL26),.BLN(BLN26),.WL(WL95));
sram_cell_6t_5 inst_cell_95_27 (.BL(BL27),.BLN(BLN27),.WL(WL95));
sram_cell_6t_5 inst_cell_95_28 (.BL(BL28),.BLN(BLN28),.WL(WL95));
sram_cell_6t_5 inst_cell_95_29 (.BL(BL29),.BLN(BLN29),.WL(WL95));
sram_cell_6t_5 inst_cell_95_30 (.BL(BL30),.BLN(BLN30),.WL(WL95));
sram_cell_6t_5 inst_cell_95_31 (.BL(BL31),.BLN(BLN31),.WL(WL95));
sram_cell_6t_5 inst_cell_95_32 (.BL(BL32),.BLN(BLN32),.WL(WL95));
sram_cell_6t_5 inst_cell_95_33 (.BL(BL33),.BLN(BLN33),.WL(WL95));
sram_cell_6t_5 inst_cell_95_34 (.BL(BL34),.BLN(BLN34),.WL(WL95));
sram_cell_6t_5 inst_cell_95_35 (.BL(BL35),.BLN(BLN35),.WL(WL95));
sram_cell_6t_5 inst_cell_95_36 (.BL(BL36),.BLN(BLN36),.WL(WL95));
sram_cell_6t_5 inst_cell_95_37 (.BL(BL37),.BLN(BLN37),.WL(WL95));
sram_cell_6t_5 inst_cell_95_38 (.BL(BL38),.BLN(BLN38),.WL(WL95));
sram_cell_6t_5 inst_cell_95_39 (.BL(BL39),.BLN(BLN39),.WL(WL95));
sram_cell_6t_5 inst_cell_95_40 (.BL(BL40),.BLN(BLN40),.WL(WL95));
sram_cell_6t_5 inst_cell_95_41 (.BL(BL41),.BLN(BLN41),.WL(WL95));
sram_cell_6t_5 inst_cell_95_42 (.BL(BL42),.BLN(BLN42),.WL(WL95));
sram_cell_6t_5 inst_cell_95_43 (.BL(BL43),.BLN(BLN43),.WL(WL95));
sram_cell_6t_5 inst_cell_95_44 (.BL(BL44),.BLN(BLN44),.WL(WL95));
sram_cell_6t_5 inst_cell_95_45 (.BL(BL45),.BLN(BLN45),.WL(WL95));
sram_cell_6t_5 inst_cell_95_46 (.BL(BL46),.BLN(BLN46),.WL(WL95));
sram_cell_6t_5 inst_cell_95_47 (.BL(BL47),.BLN(BLN47),.WL(WL95));
sram_cell_6t_5 inst_cell_95_48 (.BL(BL48),.BLN(BLN48),.WL(WL95));
sram_cell_6t_5 inst_cell_95_49 (.BL(BL49),.BLN(BLN49),.WL(WL95));
sram_cell_6t_5 inst_cell_95_50 (.BL(BL50),.BLN(BLN50),.WL(WL95));
sram_cell_6t_5 inst_cell_95_51 (.BL(BL51),.BLN(BLN51),.WL(WL95));
sram_cell_6t_5 inst_cell_95_52 (.BL(BL52),.BLN(BLN52),.WL(WL95));
sram_cell_6t_5 inst_cell_95_53 (.BL(BL53),.BLN(BLN53),.WL(WL95));
sram_cell_6t_5 inst_cell_95_54 (.BL(BL54),.BLN(BLN54),.WL(WL95));
sram_cell_6t_5 inst_cell_95_55 (.BL(BL55),.BLN(BLN55),.WL(WL95));
sram_cell_6t_5 inst_cell_95_56 (.BL(BL56),.BLN(BLN56),.WL(WL95));
sram_cell_6t_5 inst_cell_95_57 (.BL(BL57),.BLN(BLN57),.WL(WL95));
sram_cell_6t_5 inst_cell_95_58 (.BL(BL58),.BLN(BLN58),.WL(WL95));
sram_cell_6t_5 inst_cell_95_59 (.BL(BL59),.BLN(BLN59),.WL(WL95));
sram_cell_6t_5 inst_cell_95_60 (.BL(BL60),.BLN(BLN60),.WL(WL95));
sram_cell_6t_5 inst_cell_95_61 (.BL(BL61),.BLN(BLN61),.WL(WL95));
sram_cell_6t_5 inst_cell_95_62 (.BL(BL62),.BLN(BLN62),.WL(WL95));
sram_cell_6t_5 inst_cell_95_63 (.BL(BL63),.BLN(BLN63),.WL(WL95));
sram_cell_6t_5 inst_cell_95_64 (.BL(BL64),.BLN(BLN64),.WL(WL95));
sram_cell_6t_5 inst_cell_95_65 (.BL(BL65),.BLN(BLN65),.WL(WL95));
sram_cell_6t_5 inst_cell_95_66 (.BL(BL66),.BLN(BLN66),.WL(WL95));
sram_cell_6t_5 inst_cell_95_67 (.BL(BL67),.BLN(BLN67),.WL(WL95));
sram_cell_6t_5 inst_cell_95_68 (.BL(BL68),.BLN(BLN68),.WL(WL95));
sram_cell_6t_5 inst_cell_95_69 (.BL(BL69),.BLN(BLN69),.WL(WL95));
sram_cell_6t_5 inst_cell_95_70 (.BL(BL70),.BLN(BLN70),.WL(WL95));
sram_cell_6t_5 inst_cell_95_71 (.BL(BL71),.BLN(BLN71),.WL(WL95));
sram_cell_6t_5 inst_cell_95_72 (.BL(BL72),.BLN(BLN72),.WL(WL95));
sram_cell_6t_5 inst_cell_95_73 (.BL(BL73),.BLN(BLN73),.WL(WL95));
sram_cell_6t_5 inst_cell_95_74 (.BL(BL74),.BLN(BLN74),.WL(WL95));
sram_cell_6t_5 inst_cell_95_75 (.BL(BL75),.BLN(BLN75),.WL(WL95));
sram_cell_6t_5 inst_cell_95_76 (.BL(BL76),.BLN(BLN76),.WL(WL95));
sram_cell_6t_5 inst_cell_95_77 (.BL(BL77),.BLN(BLN77),.WL(WL95));
sram_cell_6t_5 inst_cell_95_78 (.BL(BL78),.BLN(BLN78),.WL(WL95));
sram_cell_6t_5 inst_cell_95_79 (.BL(BL79),.BLN(BLN79),.WL(WL95));
sram_cell_6t_5 inst_cell_95_80 (.BL(BL80),.BLN(BLN80),.WL(WL95));
sram_cell_6t_5 inst_cell_95_81 (.BL(BL81),.BLN(BLN81),.WL(WL95));
sram_cell_6t_5 inst_cell_95_82 (.BL(BL82),.BLN(BLN82),.WL(WL95));
sram_cell_6t_5 inst_cell_95_83 (.BL(BL83),.BLN(BLN83),.WL(WL95));
sram_cell_6t_5 inst_cell_95_84 (.BL(BL84),.BLN(BLN84),.WL(WL95));
sram_cell_6t_5 inst_cell_95_85 (.BL(BL85),.BLN(BLN85),.WL(WL95));
sram_cell_6t_5 inst_cell_95_86 (.BL(BL86),.BLN(BLN86),.WL(WL95));
sram_cell_6t_5 inst_cell_95_87 (.BL(BL87),.BLN(BLN87),.WL(WL95));
sram_cell_6t_5 inst_cell_95_88 (.BL(BL88),.BLN(BLN88),.WL(WL95));
sram_cell_6t_5 inst_cell_95_89 (.BL(BL89),.BLN(BLN89),.WL(WL95));
sram_cell_6t_5 inst_cell_95_90 (.BL(BL90),.BLN(BLN90),.WL(WL95));
sram_cell_6t_5 inst_cell_95_91 (.BL(BL91),.BLN(BLN91),.WL(WL95));
sram_cell_6t_5 inst_cell_95_92 (.BL(BL92),.BLN(BLN92),.WL(WL95));
sram_cell_6t_5 inst_cell_95_93 (.BL(BL93),.BLN(BLN93),.WL(WL95));
sram_cell_6t_5 inst_cell_95_94 (.BL(BL94),.BLN(BLN94),.WL(WL95));
sram_cell_6t_5 inst_cell_95_95 (.BL(BL95),.BLN(BLN95),.WL(WL95));
sram_cell_6t_5 inst_cell_95_96 (.BL(BL96),.BLN(BLN96),.WL(WL95));
sram_cell_6t_5 inst_cell_95_97 (.BL(BL97),.BLN(BLN97),.WL(WL95));
sram_cell_6t_5 inst_cell_95_98 (.BL(BL98),.BLN(BLN98),.WL(WL95));
sram_cell_6t_5 inst_cell_95_99 (.BL(BL99),.BLN(BLN99),.WL(WL95));
sram_cell_6t_5 inst_cell_95_100 (.BL(BL100),.BLN(BLN100),.WL(WL95));
sram_cell_6t_5 inst_cell_95_101 (.BL(BL101),.BLN(BLN101),.WL(WL95));
sram_cell_6t_5 inst_cell_95_102 (.BL(BL102),.BLN(BLN102),.WL(WL95));
sram_cell_6t_5 inst_cell_95_103 (.BL(BL103),.BLN(BLN103),.WL(WL95));
sram_cell_6t_5 inst_cell_95_104 (.BL(BL104),.BLN(BLN104),.WL(WL95));
sram_cell_6t_5 inst_cell_95_105 (.BL(BL105),.BLN(BLN105),.WL(WL95));
sram_cell_6t_5 inst_cell_95_106 (.BL(BL106),.BLN(BLN106),.WL(WL95));
sram_cell_6t_5 inst_cell_95_107 (.BL(BL107),.BLN(BLN107),.WL(WL95));
sram_cell_6t_5 inst_cell_95_108 (.BL(BL108),.BLN(BLN108),.WL(WL95));
sram_cell_6t_5 inst_cell_95_109 (.BL(BL109),.BLN(BLN109),.WL(WL95));
sram_cell_6t_5 inst_cell_95_110 (.BL(BL110),.BLN(BLN110),.WL(WL95));
sram_cell_6t_5 inst_cell_95_111 (.BL(BL111),.BLN(BLN111),.WL(WL95));
sram_cell_6t_5 inst_cell_95_112 (.BL(BL112),.BLN(BLN112),.WL(WL95));
sram_cell_6t_5 inst_cell_95_113 (.BL(BL113),.BLN(BLN113),.WL(WL95));
sram_cell_6t_5 inst_cell_95_114 (.BL(BL114),.BLN(BLN114),.WL(WL95));
sram_cell_6t_5 inst_cell_95_115 (.BL(BL115),.BLN(BLN115),.WL(WL95));
sram_cell_6t_5 inst_cell_95_116 (.BL(BL116),.BLN(BLN116),.WL(WL95));
sram_cell_6t_5 inst_cell_95_117 (.BL(BL117),.BLN(BLN117),.WL(WL95));
sram_cell_6t_5 inst_cell_95_118 (.BL(BL118),.BLN(BLN118),.WL(WL95));
sram_cell_6t_5 inst_cell_95_119 (.BL(BL119),.BLN(BLN119),.WL(WL95));
sram_cell_6t_5 inst_cell_95_120 (.BL(BL120),.BLN(BLN120),.WL(WL95));
sram_cell_6t_5 inst_cell_95_121 (.BL(BL121),.BLN(BLN121),.WL(WL95));
sram_cell_6t_5 inst_cell_95_122 (.BL(BL122),.BLN(BLN122),.WL(WL95));
sram_cell_6t_5 inst_cell_95_123 (.BL(BL123),.BLN(BLN123),.WL(WL95));
sram_cell_6t_5 inst_cell_95_124 (.BL(BL124),.BLN(BLN124),.WL(WL95));
sram_cell_6t_5 inst_cell_95_125 (.BL(BL125),.BLN(BLN125),.WL(WL95));
sram_cell_6t_5 inst_cell_95_126 (.BL(BL126),.BLN(BLN126),.WL(WL95));
sram_cell_6t_5 inst_cell_95_127 (.BL(BL127),.BLN(BLN127),.WL(WL95));
sram_cell_6t_5 inst_cell_96_0 (.BL(BL0),.BLN(BLN0),.WL(WL96));
sram_cell_6t_5 inst_cell_96_1 (.BL(BL1),.BLN(BLN1),.WL(WL96));
sram_cell_6t_5 inst_cell_96_2 (.BL(BL2),.BLN(BLN2),.WL(WL96));
sram_cell_6t_5 inst_cell_96_3 (.BL(BL3),.BLN(BLN3),.WL(WL96));
sram_cell_6t_5 inst_cell_96_4 (.BL(BL4),.BLN(BLN4),.WL(WL96));
sram_cell_6t_5 inst_cell_96_5 (.BL(BL5),.BLN(BLN5),.WL(WL96));
sram_cell_6t_5 inst_cell_96_6 (.BL(BL6),.BLN(BLN6),.WL(WL96));
sram_cell_6t_5 inst_cell_96_7 (.BL(BL7),.BLN(BLN7),.WL(WL96));
sram_cell_6t_5 inst_cell_96_8 (.BL(BL8),.BLN(BLN8),.WL(WL96));
sram_cell_6t_5 inst_cell_96_9 (.BL(BL9),.BLN(BLN9),.WL(WL96));
sram_cell_6t_5 inst_cell_96_10 (.BL(BL10),.BLN(BLN10),.WL(WL96));
sram_cell_6t_5 inst_cell_96_11 (.BL(BL11),.BLN(BLN11),.WL(WL96));
sram_cell_6t_5 inst_cell_96_12 (.BL(BL12),.BLN(BLN12),.WL(WL96));
sram_cell_6t_5 inst_cell_96_13 (.BL(BL13),.BLN(BLN13),.WL(WL96));
sram_cell_6t_5 inst_cell_96_14 (.BL(BL14),.BLN(BLN14),.WL(WL96));
sram_cell_6t_5 inst_cell_96_15 (.BL(BL15),.BLN(BLN15),.WL(WL96));
sram_cell_6t_5 inst_cell_96_16 (.BL(BL16),.BLN(BLN16),.WL(WL96));
sram_cell_6t_5 inst_cell_96_17 (.BL(BL17),.BLN(BLN17),.WL(WL96));
sram_cell_6t_5 inst_cell_96_18 (.BL(BL18),.BLN(BLN18),.WL(WL96));
sram_cell_6t_5 inst_cell_96_19 (.BL(BL19),.BLN(BLN19),.WL(WL96));
sram_cell_6t_5 inst_cell_96_20 (.BL(BL20),.BLN(BLN20),.WL(WL96));
sram_cell_6t_5 inst_cell_96_21 (.BL(BL21),.BLN(BLN21),.WL(WL96));
sram_cell_6t_5 inst_cell_96_22 (.BL(BL22),.BLN(BLN22),.WL(WL96));
sram_cell_6t_5 inst_cell_96_23 (.BL(BL23),.BLN(BLN23),.WL(WL96));
sram_cell_6t_5 inst_cell_96_24 (.BL(BL24),.BLN(BLN24),.WL(WL96));
sram_cell_6t_5 inst_cell_96_25 (.BL(BL25),.BLN(BLN25),.WL(WL96));
sram_cell_6t_5 inst_cell_96_26 (.BL(BL26),.BLN(BLN26),.WL(WL96));
sram_cell_6t_5 inst_cell_96_27 (.BL(BL27),.BLN(BLN27),.WL(WL96));
sram_cell_6t_5 inst_cell_96_28 (.BL(BL28),.BLN(BLN28),.WL(WL96));
sram_cell_6t_5 inst_cell_96_29 (.BL(BL29),.BLN(BLN29),.WL(WL96));
sram_cell_6t_5 inst_cell_96_30 (.BL(BL30),.BLN(BLN30),.WL(WL96));
sram_cell_6t_5 inst_cell_96_31 (.BL(BL31),.BLN(BLN31),.WL(WL96));
sram_cell_6t_5 inst_cell_96_32 (.BL(BL32),.BLN(BLN32),.WL(WL96));
sram_cell_6t_5 inst_cell_96_33 (.BL(BL33),.BLN(BLN33),.WL(WL96));
sram_cell_6t_5 inst_cell_96_34 (.BL(BL34),.BLN(BLN34),.WL(WL96));
sram_cell_6t_5 inst_cell_96_35 (.BL(BL35),.BLN(BLN35),.WL(WL96));
sram_cell_6t_5 inst_cell_96_36 (.BL(BL36),.BLN(BLN36),.WL(WL96));
sram_cell_6t_5 inst_cell_96_37 (.BL(BL37),.BLN(BLN37),.WL(WL96));
sram_cell_6t_5 inst_cell_96_38 (.BL(BL38),.BLN(BLN38),.WL(WL96));
sram_cell_6t_5 inst_cell_96_39 (.BL(BL39),.BLN(BLN39),.WL(WL96));
sram_cell_6t_5 inst_cell_96_40 (.BL(BL40),.BLN(BLN40),.WL(WL96));
sram_cell_6t_5 inst_cell_96_41 (.BL(BL41),.BLN(BLN41),.WL(WL96));
sram_cell_6t_5 inst_cell_96_42 (.BL(BL42),.BLN(BLN42),.WL(WL96));
sram_cell_6t_5 inst_cell_96_43 (.BL(BL43),.BLN(BLN43),.WL(WL96));
sram_cell_6t_5 inst_cell_96_44 (.BL(BL44),.BLN(BLN44),.WL(WL96));
sram_cell_6t_5 inst_cell_96_45 (.BL(BL45),.BLN(BLN45),.WL(WL96));
sram_cell_6t_5 inst_cell_96_46 (.BL(BL46),.BLN(BLN46),.WL(WL96));
sram_cell_6t_5 inst_cell_96_47 (.BL(BL47),.BLN(BLN47),.WL(WL96));
sram_cell_6t_5 inst_cell_96_48 (.BL(BL48),.BLN(BLN48),.WL(WL96));
sram_cell_6t_5 inst_cell_96_49 (.BL(BL49),.BLN(BLN49),.WL(WL96));
sram_cell_6t_5 inst_cell_96_50 (.BL(BL50),.BLN(BLN50),.WL(WL96));
sram_cell_6t_5 inst_cell_96_51 (.BL(BL51),.BLN(BLN51),.WL(WL96));
sram_cell_6t_5 inst_cell_96_52 (.BL(BL52),.BLN(BLN52),.WL(WL96));
sram_cell_6t_5 inst_cell_96_53 (.BL(BL53),.BLN(BLN53),.WL(WL96));
sram_cell_6t_5 inst_cell_96_54 (.BL(BL54),.BLN(BLN54),.WL(WL96));
sram_cell_6t_5 inst_cell_96_55 (.BL(BL55),.BLN(BLN55),.WL(WL96));
sram_cell_6t_5 inst_cell_96_56 (.BL(BL56),.BLN(BLN56),.WL(WL96));
sram_cell_6t_5 inst_cell_96_57 (.BL(BL57),.BLN(BLN57),.WL(WL96));
sram_cell_6t_5 inst_cell_96_58 (.BL(BL58),.BLN(BLN58),.WL(WL96));
sram_cell_6t_5 inst_cell_96_59 (.BL(BL59),.BLN(BLN59),.WL(WL96));
sram_cell_6t_5 inst_cell_96_60 (.BL(BL60),.BLN(BLN60),.WL(WL96));
sram_cell_6t_5 inst_cell_96_61 (.BL(BL61),.BLN(BLN61),.WL(WL96));
sram_cell_6t_5 inst_cell_96_62 (.BL(BL62),.BLN(BLN62),.WL(WL96));
sram_cell_6t_5 inst_cell_96_63 (.BL(BL63),.BLN(BLN63),.WL(WL96));
sram_cell_6t_5 inst_cell_96_64 (.BL(BL64),.BLN(BLN64),.WL(WL96));
sram_cell_6t_5 inst_cell_96_65 (.BL(BL65),.BLN(BLN65),.WL(WL96));
sram_cell_6t_5 inst_cell_96_66 (.BL(BL66),.BLN(BLN66),.WL(WL96));
sram_cell_6t_5 inst_cell_96_67 (.BL(BL67),.BLN(BLN67),.WL(WL96));
sram_cell_6t_5 inst_cell_96_68 (.BL(BL68),.BLN(BLN68),.WL(WL96));
sram_cell_6t_5 inst_cell_96_69 (.BL(BL69),.BLN(BLN69),.WL(WL96));
sram_cell_6t_5 inst_cell_96_70 (.BL(BL70),.BLN(BLN70),.WL(WL96));
sram_cell_6t_5 inst_cell_96_71 (.BL(BL71),.BLN(BLN71),.WL(WL96));
sram_cell_6t_5 inst_cell_96_72 (.BL(BL72),.BLN(BLN72),.WL(WL96));
sram_cell_6t_5 inst_cell_96_73 (.BL(BL73),.BLN(BLN73),.WL(WL96));
sram_cell_6t_5 inst_cell_96_74 (.BL(BL74),.BLN(BLN74),.WL(WL96));
sram_cell_6t_5 inst_cell_96_75 (.BL(BL75),.BLN(BLN75),.WL(WL96));
sram_cell_6t_5 inst_cell_96_76 (.BL(BL76),.BLN(BLN76),.WL(WL96));
sram_cell_6t_5 inst_cell_96_77 (.BL(BL77),.BLN(BLN77),.WL(WL96));
sram_cell_6t_5 inst_cell_96_78 (.BL(BL78),.BLN(BLN78),.WL(WL96));
sram_cell_6t_5 inst_cell_96_79 (.BL(BL79),.BLN(BLN79),.WL(WL96));
sram_cell_6t_5 inst_cell_96_80 (.BL(BL80),.BLN(BLN80),.WL(WL96));
sram_cell_6t_5 inst_cell_96_81 (.BL(BL81),.BLN(BLN81),.WL(WL96));
sram_cell_6t_5 inst_cell_96_82 (.BL(BL82),.BLN(BLN82),.WL(WL96));
sram_cell_6t_5 inst_cell_96_83 (.BL(BL83),.BLN(BLN83),.WL(WL96));
sram_cell_6t_5 inst_cell_96_84 (.BL(BL84),.BLN(BLN84),.WL(WL96));
sram_cell_6t_5 inst_cell_96_85 (.BL(BL85),.BLN(BLN85),.WL(WL96));
sram_cell_6t_5 inst_cell_96_86 (.BL(BL86),.BLN(BLN86),.WL(WL96));
sram_cell_6t_5 inst_cell_96_87 (.BL(BL87),.BLN(BLN87),.WL(WL96));
sram_cell_6t_5 inst_cell_96_88 (.BL(BL88),.BLN(BLN88),.WL(WL96));
sram_cell_6t_5 inst_cell_96_89 (.BL(BL89),.BLN(BLN89),.WL(WL96));
sram_cell_6t_5 inst_cell_96_90 (.BL(BL90),.BLN(BLN90),.WL(WL96));
sram_cell_6t_5 inst_cell_96_91 (.BL(BL91),.BLN(BLN91),.WL(WL96));
sram_cell_6t_5 inst_cell_96_92 (.BL(BL92),.BLN(BLN92),.WL(WL96));
sram_cell_6t_5 inst_cell_96_93 (.BL(BL93),.BLN(BLN93),.WL(WL96));
sram_cell_6t_5 inst_cell_96_94 (.BL(BL94),.BLN(BLN94),.WL(WL96));
sram_cell_6t_5 inst_cell_96_95 (.BL(BL95),.BLN(BLN95),.WL(WL96));
sram_cell_6t_5 inst_cell_96_96 (.BL(BL96),.BLN(BLN96),.WL(WL96));
sram_cell_6t_5 inst_cell_96_97 (.BL(BL97),.BLN(BLN97),.WL(WL96));
sram_cell_6t_5 inst_cell_96_98 (.BL(BL98),.BLN(BLN98),.WL(WL96));
sram_cell_6t_5 inst_cell_96_99 (.BL(BL99),.BLN(BLN99),.WL(WL96));
sram_cell_6t_5 inst_cell_96_100 (.BL(BL100),.BLN(BLN100),.WL(WL96));
sram_cell_6t_5 inst_cell_96_101 (.BL(BL101),.BLN(BLN101),.WL(WL96));
sram_cell_6t_5 inst_cell_96_102 (.BL(BL102),.BLN(BLN102),.WL(WL96));
sram_cell_6t_5 inst_cell_96_103 (.BL(BL103),.BLN(BLN103),.WL(WL96));
sram_cell_6t_5 inst_cell_96_104 (.BL(BL104),.BLN(BLN104),.WL(WL96));
sram_cell_6t_5 inst_cell_96_105 (.BL(BL105),.BLN(BLN105),.WL(WL96));
sram_cell_6t_5 inst_cell_96_106 (.BL(BL106),.BLN(BLN106),.WL(WL96));
sram_cell_6t_5 inst_cell_96_107 (.BL(BL107),.BLN(BLN107),.WL(WL96));
sram_cell_6t_5 inst_cell_96_108 (.BL(BL108),.BLN(BLN108),.WL(WL96));
sram_cell_6t_5 inst_cell_96_109 (.BL(BL109),.BLN(BLN109),.WL(WL96));
sram_cell_6t_5 inst_cell_96_110 (.BL(BL110),.BLN(BLN110),.WL(WL96));
sram_cell_6t_5 inst_cell_96_111 (.BL(BL111),.BLN(BLN111),.WL(WL96));
sram_cell_6t_5 inst_cell_96_112 (.BL(BL112),.BLN(BLN112),.WL(WL96));
sram_cell_6t_5 inst_cell_96_113 (.BL(BL113),.BLN(BLN113),.WL(WL96));
sram_cell_6t_5 inst_cell_96_114 (.BL(BL114),.BLN(BLN114),.WL(WL96));
sram_cell_6t_5 inst_cell_96_115 (.BL(BL115),.BLN(BLN115),.WL(WL96));
sram_cell_6t_5 inst_cell_96_116 (.BL(BL116),.BLN(BLN116),.WL(WL96));
sram_cell_6t_5 inst_cell_96_117 (.BL(BL117),.BLN(BLN117),.WL(WL96));
sram_cell_6t_5 inst_cell_96_118 (.BL(BL118),.BLN(BLN118),.WL(WL96));
sram_cell_6t_5 inst_cell_96_119 (.BL(BL119),.BLN(BLN119),.WL(WL96));
sram_cell_6t_5 inst_cell_96_120 (.BL(BL120),.BLN(BLN120),.WL(WL96));
sram_cell_6t_5 inst_cell_96_121 (.BL(BL121),.BLN(BLN121),.WL(WL96));
sram_cell_6t_5 inst_cell_96_122 (.BL(BL122),.BLN(BLN122),.WL(WL96));
sram_cell_6t_5 inst_cell_96_123 (.BL(BL123),.BLN(BLN123),.WL(WL96));
sram_cell_6t_5 inst_cell_96_124 (.BL(BL124),.BLN(BLN124),.WL(WL96));
sram_cell_6t_5 inst_cell_96_125 (.BL(BL125),.BLN(BLN125),.WL(WL96));
sram_cell_6t_5 inst_cell_96_126 (.BL(BL126),.BLN(BLN126),.WL(WL96));
sram_cell_6t_5 inst_cell_96_127 (.BL(BL127),.BLN(BLN127),.WL(WL96));
sram_cell_6t_5 inst_cell_97_0 (.BL(BL0),.BLN(BLN0),.WL(WL97));
sram_cell_6t_5 inst_cell_97_1 (.BL(BL1),.BLN(BLN1),.WL(WL97));
sram_cell_6t_5 inst_cell_97_2 (.BL(BL2),.BLN(BLN2),.WL(WL97));
sram_cell_6t_5 inst_cell_97_3 (.BL(BL3),.BLN(BLN3),.WL(WL97));
sram_cell_6t_5 inst_cell_97_4 (.BL(BL4),.BLN(BLN4),.WL(WL97));
sram_cell_6t_5 inst_cell_97_5 (.BL(BL5),.BLN(BLN5),.WL(WL97));
sram_cell_6t_5 inst_cell_97_6 (.BL(BL6),.BLN(BLN6),.WL(WL97));
sram_cell_6t_5 inst_cell_97_7 (.BL(BL7),.BLN(BLN7),.WL(WL97));
sram_cell_6t_5 inst_cell_97_8 (.BL(BL8),.BLN(BLN8),.WL(WL97));
sram_cell_6t_5 inst_cell_97_9 (.BL(BL9),.BLN(BLN9),.WL(WL97));
sram_cell_6t_5 inst_cell_97_10 (.BL(BL10),.BLN(BLN10),.WL(WL97));
sram_cell_6t_5 inst_cell_97_11 (.BL(BL11),.BLN(BLN11),.WL(WL97));
sram_cell_6t_5 inst_cell_97_12 (.BL(BL12),.BLN(BLN12),.WL(WL97));
sram_cell_6t_5 inst_cell_97_13 (.BL(BL13),.BLN(BLN13),.WL(WL97));
sram_cell_6t_5 inst_cell_97_14 (.BL(BL14),.BLN(BLN14),.WL(WL97));
sram_cell_6t_5 inst_cell_97_15 (.BL(BL15),.BLN(BLN15),.WL(WL97));
sram_cell_6t_5 inst_cell_97_16 (.BL(BL16),.BLN(BLN16),.WL(WL97));
sram_cell_6t_5 inst_cell_97_17 (.BL(BL17),.BLN(BLN17),.WL(WL97));
sram_cell_6t_5 inst_cell_97_18 (.BL(BL18),.BLN(BLN18),.WL(WL97));
sram_cell_6t_5 inst_cell_97_19 (.BL(BL19),.BLN(BLN19),.WL(WL97));
sram_cell_6t_5 inst_cell_97_20 (.BL(BL20),.BLN(BLN20),.WL(WL97));
sram_cell_6t_5 inst_cell_97_21 (.BL(BL21),.BLN(BLN21),.WL(WL97));
sram_cell_6t_5 inst_cell_97_22 (.BL(BL22),.BLN(BLN22),.WL(WL97));
sram_cell_6t_5 inst_cell_97_23 (.BL(BL23),.BLN(BLN23),.WL(WL97));
sram_cell_6t_5 inst_cell_97_24 (.BL(BL24),.BLN(BLN24),.WL(WL97));
sram_cell_6t_5 inst_cell_97_25 (.BL(BL25),.BLN(BLN25),.WL(WL97));
sram_cell_6t_5 inst_cell_97_26 (.BL(BL26),.BLN(BLN26),.WL(WL97));
sram_cell_6t_5 inst_cell_97_27 (.BL(BL27),.BLN(BLN27),.WL(WL97));
sram_cell_6t_5 inst_cell_97_28 (.BL(BL28),.BLN(BLN28),.WL(WL97));
sram_cell_6t_5 inst_cell_97_29 (.BL(BL29),.BLN(BLN29),.WL(WL97));
sram_cell_6t_5 inst_cell_97_30 (.BL(BL30),.BLN(BLN30),.WL(WL97));
sram_cell_6t_5 inst_cell_97_31 (.BL(BL31),.BLN(BLN31),.WL(WL97));
sram_cell_6t_5 inst_cell_97_32 (.BL(BL32),.BLN(BLN32),.WL(WL97));
sram_cell_6t_5 inst_cell_97_33 (.BL(BL33),.BLN(BLN33),.WL(WL97));
sram_cell_6t_5 inst_cell_97_34 (.BL(BL34),.BLN(BLN34),.WL(WL97));
sram_cell_6t_5 inst_cell_97_35 (.BL(BL35),.BLN(BLN35),.WL(WL97));
sram_cell_6t_5 inst_cell_97_36 (.BL(BL36),.BLN(BLN36),.WL(WL97));
sram_cell_6t_5 inst_cell_97_37 (.BL(BL37),.BLN(BLN37),.WL(WL97));
sram_cell_6t_5 inst_cell_97_38 (.BL(BL38),.BLN(BLN38),.WL(WL97));
sram_cell_6t_5 inst_cell_97_39 (.BL(BL39),.BLN(BLN39),.WL(WL97));
sram_cell_6t_5 inst_cell_97_40 (.BL(BL40),.BLN(BLN40),.WL(WL97));
sram_cell_6t_5 inst_cell_97_41 (.BL(BL41),.BLN(BLN41),.WL(WL97));
sram_cell_6t_5 inst_cell_97_42 (.BL(BL42),.BLN(BLN42),.WL(WL97));
sram_cell_6t_5 inst_cell_97_43 (.BL(BL43),.BLN(BLN43),.WL(WL97));
sram_cell_6t_5 inst_cell_97_44 (.BL(BL44),.BLN(BLN44),.WL(WL97));
sram_cell_6t_5 inst_cell_97_45 (.BL(BL45),.BLN(BLN45),.WL(WL97));
sram_cell_6t_5 inst_cell_97_46 (.BL(BL46),.BLN(BLN46),.WL(WL97));
sram_cell_6t_5 inst_cell_97_47 (.BL(BL47),.BLN(BLN47),.WL(WL97));
sram_cell_6t_5 inst_cell_97_48 (.BL(BL48),.BLN(BLN48),.WL(WL97));
sram_cell_6t_5 inst_cell_97_49 (.BL(BL49),.BLN(BLN49),.WL(WL97));
sram_cell_6t_5 inst_cell_97_50 (.BL(BL50),.BLN(BLN50),.WL(WL97));
sram_cell_6t_5 inst_cell_97_51 (.BL(BL51),.BLN(BLN51),.WL(WL97));
sram_cell_6t_5 inst_cell_97_52 (.BL(BL52),.BLN(BLN52),.WL(WL97));
sram_cell_6t_5 inst_cell_97_53 (.BL(BL53),.BLN(BLN53),.WL(WL97));
sram_cell_6t_5 inst_cell_97_54 (.BL(BL54),.BLN(BLN54),.WL(WL97));
sram_cell_6t_5 inst_cell_97_55 (.BL(BL55),.BLN(BLN55),.WL(WL97));
sram_cell_6t_5 inst_cell_97_56 (.BL(BL56),.BLN(BLN56),.WL(WL97));
sram_cell_6t_5 inst_cell_97_57 (.BL(BL57),.BLN(BLN57),.WL(WL97));
sram_cell_6t_5 inst_cell_97_58 (.BL(BL58),.BLN(BLN58),.WL(WL97));
sram_cell_6t_5 inst_cell_97_59 (.BL(BL59),.BLN(BLN59),.WL(WL97));
sram_cell_6t_5 inst_cell_97_60 (.BL(BL60),.BLN(BLN60),.WL(WL97));
sram_cell_6t_5 inst_cell_97_61 (.BL(BL61),.BLN(BLN61),.WL(WL97));
sram_cell_6t_5 inst_cell_97_62 (.BL(BL62),.BLN(BLN62),.WL(WL97));
sram_cell_6t_5 inst_cell_97_63 (.BL(BL63),.BLN(BLN63),.WL(WL97));
sram_cell_6t_5 inst_cell_97_64 (.BL(BL64),.BLN(BLN64),.WL(WL97));
sram_cell_6t_5 inst_cell_97_65 (.BL(BL65),.BLN(BLN65),.WL(WL97));
sram_cell_6t_5 inst_cell_97_66 (.BL(BL66),.BLN(BLN66),.WL(WL97));
sram_cell_6t_5 inst_cell_97_67 (.BL(BL67),.BLN(BLN67),.WL(WL97));
sram_cell_6t_5 inst_cell_97_68 (.BL(BL68),.BLN(BLN68),.WL(WL97));
sram_cell_6t_5 inst_cell_97_69 (.BL(BL69),.BLN(BLN69),.WL(WL97));
sram_cell_6t_5 inst_cell_97_70 (.BL(BL70),.BLN(BLN70),.WL(WL97));
sram_cell_6t_5 inst_cell_97_71 (.BL(BL71),.BLN(BLN71),.WL(WL97));
sram_cell_6t_5 inst_cell_97_72 (.BL(BL72),.BLN(BLN72),.WL(WL97));
sram_cell_6t_5 inst_cell_97_73 (.BL(BL73),.BLN(BLN73),.WL(WL97));
sram_cell_6t_5 inst_cell_97_74 (.BL(BL74),.BLN(BLN74),.WL(WL97));
sram_cell_6t_5 inst_cell_97_75 (.BL(BL75),.BLN(BLN75),.WL(WL97));
sram_cell_6t_5 inst_cell_97_76 (.BL(BL76),.BLN(BLN76),.WL(WL97));
sram_cell_6t_5 inst_cell_97_77 (.BL(BL77),.BLN(BLN77),.WL(WL97));
sram_cell_6t_5 inst_cell_97_78 (.BL(BL78),.BLN(BLN78),.WL(WL97));
sram_cell_6t_5 inst_cell_97_79 (.BL(BL79),.BLN(BLN79),.WL(WL97));
sram_cell_6t_5 inst_cell_97_80 (.BL(BL80),.BLN(BLN80),.WL(WL97));
sram_cell_6t_5 inst_cell_97_81 (.BL(BL81),.BLN(BLN81),.WL(WL97));
sram_cell_6t_5 inst_cell_97_82 (.BL(BL82),.BLN(BLN82),.WL(WL97));
sram_cell_6t_5 inst_cell_97_83 (.BL(BL83),.BLN(BLN83),.WL(WL97));
sram_cell_6t_5 inst_cell_97_84 (.BL(BL84),.BLN(BLN84),.WL(WL97));
sram_cell_6t_5 inst_cell_97_85 (.BL(BL85),.BLN(BLN85),.WL(WL97));
sram_cell_6t_5 inst_cell_97_86 (.BL(BL86),.BLN(BLN86),.WL(WL97));
sram_cell_6t_5 inst_cell_97_87 (.BL(BL87),.BLN(BLN87),.WL(WL97));
sram_cell_6t_5 inst_cell_97_88 (.BL(BL88),.BLN(BLN88),.WL(WL97));
sram_cell_6t_5 inst_cell_97_89 (.BL(BL89),.BLN(BLN89),.WL(WL97));
sram_cell_6t_5 inst_cell_97_90 (.BL(BL90),.BLN(BLN90),.WL(WL97));
sram_cell_6t_5 inst_cell_97_91 (.BL(BL91),.BLN(BLN91),.WL(WL97));
sram_cell_6t_5 inst_cell_97_92 (.BL(BL92),.BLN(BLN92),.WL(WL97));
sram_cell_6t_5 inst_cell_97_93 (.BL(BL93),.BLN(BLN93),.WL(WL97));
sram_cell_6t_5 inst_cell_97_94 (.BL(BL94),.BLN(BLN94),.WL(WL97));
sram_cell_6t_5 inst_cell_97_95 (.BL(BL95),.BLN(BLN95),.WL(WL97));
sram_cell_6t_5 inst_cell_97_96 (.BL(BL96),.BLN(BLN96),.WL(WL97));
sram_cell_6t_5 inst_cell_97_97 (.BL(BL97),.BLN(BLN97),.WL(WL97));
sram_cell_6t_5 inst_cell_97_98 (.BL(BL98),.BLN(BLN98),.WL(WL97));
sram_cell_6t_5 inst_cell_97_99 (.BL(BL99),.BLN(BLN99),.WL(WL97));
sram_cell_6t_5 inst_cell_97_100 (.BL(BL100),.BLN(BLN100),.WL(WL97));
sram_cell_6t_5 inst_cell_97_101 (.BL(BL101),.BLN(BLN101),.WL(WL97));
sram_cell_6t_5 inst_cell_97_102 (.BL(BL102),.BLN(BLN102),.WL(WL97));
sram_cell_6t_5 inst_cell_97_103 (.BL(BL103),.BLN(BLN103),.WL(WL97));
sram_cell_6t_5 inst_cell_97_104 (.BL(BL104),.BLN(BLN104),.WL(WL97));
sram_cell_6t_5 inst_cell_97_105 (.BL(BL105),.BLN(BLN105),.WL(WL97));
sram_cell_6t_5 inst_cell_97_106 (.BL(BL106),.BLN(BLN106),.WL(WL97));
sram_cell_6t_5 inst_cell_97_107 (.BL(BL107),.BLN(BLN107),.WL(WL97));
sram_cell_6t_5 inst_cell_97_108 (.BL(BL108),.BLN(BLN108),.WL(WL97));
sram_cell_6t_5 inst_cell_97_109 (.BL(BL109),.BLN(BLN109),.WL(WL97));
sram_cell_6t_5 inst_cell_97_110 (.BL(BL110),.BLN(BLN110),.WL(WL97));
sram_cell_6t_5 inst_cell_97_111 (.BL(BL111),.BLN(BLN111),.WL(WL97));
sram_cell_6t_5 inst_cell_97_112 (.BL(BL112),.BLN(BLN112),.WL(WL97));
sram_cell_6t_5 inst_cell_97_113 (.BL(BL113),.BLN(BLN113),.WL(WL97));
sram_cell_6t_5 inst_cell_97_114 (.BL(BL114),.BLN(BLN114),.WL(WL97));
sram_cell_6t_5 inst_cell_97_115 (.BL(BL115),.BLN(BLN115),.WL(WL97));
sram_cell_6t_5 inst_cell_97_116 (.BL(BL116),.BLN(BLN116),.WL(WL97));
sram_cell_6t_5 inst_cell_97_117 (.BL(BL117),.BLN(BLN117),.WL(WL97));
sram_cell_6t_5 inst_cell_97_118 (.BL(BL118),.BLN(BLN118),.WL(WL97));
sram_cell_6t_5 inst_cell_97_119 (.BL(BL119),.BLN(BLN119),.WL(WL97));
sram_cell_6t_5 inst_cell_97_120 (.BL(BL120),.BLN(BLN120),.WL(WL97));
sram_cell_6t_5 inst_cell_97_121 (.BL(BL121),.BLN(BLN121),.WL(WL97));
sram_cell_6t_5 inst_cell_97_122 (.BL(BL122),.BLN(BLN122),.WL(WL97));
sram_cell_6t_5 inst_cell_97_123 (.BL(BL123),.BLN(BLN123),.WL(WL97));
sram_cell_6t_5 inst_cell_97_124 (.BL(BL124),.BLN(BLN124),.WL(WL97));
sram_cell_6t_5 inst_cell_97_125 (.BL(BL125),.BLN(BLN125),.WL(WL97));
sram_cell_6t_5 inst_cell_97_126 (.BL(BL126),.BLN(BLN126),.WL(WL97));
sram_cell_6t_5 inst_cell_97_127 (.BL(BL127),.BLN(BLN127),.WL(WL97));
sram_cell_6t_5 inst_cell_98_0 (.BL(BL0),.BLN(BLN0),.WL(WL98));
sram_cell_6t_5 inst_cell_98_1 (.BL(BL1),.BLN(BLN1),.WL(WL98));
sram_cell_6t_5 inst_cell_98_2 (.BL(BL2),.BLN(BLN2),.WL(WL98));
sram_cell_6t_5 inst_cell_98_3 (.BL(BL3),.BLN(BLN3),.WL(WL98));
sram_cell_6t_5 inst_cell_98_4 (.BL(BL4),.BLN(BLN4),.WL(WL98));
sram_cell_6t_5 inst_cell_98_5 (.BL(BL5),.BLN(BLN5),.WL(WL98));
sram_cell_6t_5 inst_cell_98_6 (.BL(BL6),.BLN(BLN6),.WL(WL98));
sram_cell_6t_5 inst_cell_98_7 (.BL(BL7),.BLN(BLN7),.WL(WL98));
sram_cell_6t_5 inst_cell_98_8 (.BL(BL8),.BLN(BLN8),.WL(WL98));
sram_cell_6t_5 inst_cell_98_9 (.BL(BL9),.BLN(BLN9),.WL(WL98));
sram_cell_6t_5 inst_cell_98_10 (.BL(BL10),.BLN(BLN10),.WL(WL98));
sram_cell_6t_5 inst_cell_98_11 (.BL(BL11),.BLN(BLN11),.WL(WL98));
sram_cell_6t_5 inst_cell_98_12 (.BL(BL12),.BLN(BLN12),.WL(WL98));
sram_cell_6t_5 inst_cell_98_13 (.BL(BL13),.BLN(BLN13),.WL(WL98));
sram_cell_6t_5 inst_cell_98_14 (.BL(BL14),.BLN(BLN14),.WL(WL98));
sram_cell_6t_5 inst_cell_98_15 (.BL(BL15),.BLN(BLN15),.WL(WL98));
sram_cell_6t_5 inst_cell_98_16 (.BL(BL16),.BLN(BLN16),.WL(WL98));
sram_cell_6t_5 inst_cell_98_17 (.BL(BL17),.BLN(BLN17),.WL(WL98));
sram_cell_6t_5 inst_cell_98_18 (.BL(BL18),.BLN(BLN18),.WL(WL98));
sram_cell_6t_5 inst_cell_98_19 (.BL(BL19),.BLN(BLN19),.WL(WL98));
sram_cell_6t_5 inst_cell_98_20 (.BL(BL20),.BLN(BLN20),.WL(WL98));
sram_cell_6t_5 inst_cell_98_21 (.BL(BL21),.BLN(BLN21),.WL(WL98));
sram_cell_6t_5 inst_cell_98_22 (.BL(BL22),.BLN(BLN22),.WL(WL98));
sram_cell_6t_5 inst_cell_98_23 (.BL(BL23),.BLN(BLN23),.WL(WL98));
sram_cell_6t_5 inst_cell_98_24 (.BL(BL24),.BLN(BLN24),.WL(WL98));
sram_cell_6t_5 inst_cell_98_25 (.BL(BL25),.BLN(BLN25),.WL(WL98));
sram_cell_6t_5 inst_cell_98_26 (.BL(BL26),.BLN(BLN26),.WL(WL98));
sram_cell_6t_5 inst_cell_98_27 (.BL(BL27),.BLN(BLN27),.WL(WL98));
sram_cell_6t_5 inst_cell_98_28 (.BL(BL28),.BLN(BLN28),.WL(WL98));
sram_cell_6t_5 inst_cell_98_29 (.BL(BL29),.BLN(BLN29),.WL(WL98));
sram_cell_6t_5 inst_cell_98_30 (.BL(BL30),.BLN(BLN30),.WL(WL98));
sram_cell_6t_5 inst_cell_98_31 (.BL(BL31),.BLN(BLN31),.WL(WL98));
sram_cell_6t_5 inst_cell_98_32 (.BL(BL32),.BLN(BLN32),.WL(WL98));
sram_cell_6t_5 inst_cell_98_33 (.BL(BL33),.BLN(BLN33),.WL(WL98));
sram_cell_6t_5 inst_cell_98_34 (.BL(BL34),.BLN(BLN34),.WL(WL98));
sram_cell_6t_5 inst_cell_98_35 (.BL(BL35),.BLN(BLN35),.WL(WL98));
sram_cell_6t_5 inst_cell_98_36 (.BL(BL36),.BLN(BLN36),.WL(WL98));
sram_cell_6t_5 inst_cell_98_37 (.BL(BL37),.BLN(BLN37),.WL(WL98));
sram_cell_6t_5 inst_cell_98_38 (.BL(BL38),.BLN(BLN38),.WL(WL98));
sram_cell_6t_5 inst_cell_98_39 (.BL(BL39),.BLN(BLN39),.WL(WL98));
sram_cell_6t_5 inst_cell_98_40 (.BL(BL40),.BLN(BLN40),.WL(WL98));
sram_cell_6t_5 inst_cell_98_41 (.BL(BL41),.BLN(BLN41),.WL(WL98));
sram_cell_6t_5 inst_cell_98_42 (.BL(BL42),.BLN(BLN42),.WL(WL98));
sram_cell_6t_5 inst_cell_98_43 (.BL(BL43),.BLN(BLN43),.WL(WL98));
sram_cell_6t_5 inst_cell_98_44 (.BL(BL44),.BLN(BLN44),.WL(WL98));
sram_cell_6t_5 inst_cell_98_45 (.BL(BL45),.BLN(BLN45),.WL(WL98));
sram_cell_6t_5 inst_cell_98_46 (.BL(BL46),.BLN(BLN46),.WL(WL98));
sram_cell_6t_5 inst_cell_98_47 (.BL(BL47),.BLN(BLN47),.WL(WL98));
sram_cell_6t_5 inst_cell_98_48 (.BL(BL48),.BLN(BLN48),.WL(WL98));
sram_cell_6t_5 inst_cell_98_49 (.BL(BL49),.BLN(BLN49),.WL(WL98));
sram_cell_6t_5 inst_cell_98_50 (.BL(BL50),.BLN(BLN50),.WL(WL98));
sram_cell_6t_5 inst_cell_98_51 (.BL(BL51),.BLN(BLN51),.WL(WL98));
sram_cell_6t_5 inst_cell_98_52 (.BL(BL52),.BLN(BLN52),.WL(WL98));
sram_cell_6t_5 inst_cell_98_53 (.BL(BL53),.BLN(BLN53),.WL(WL98));
sram_cell_6t_5 inst_cell_98_54 (.BL(BL54),.BLN(BLN54),.WL(WL98));
sram_cell_6t_5 inst_cell_98_55 (.BL(BL55),.BLN(BLN55),.WL(WL98));
sram_cell_6t_5 inst_cell_98_56 (.BL(BL56),.BLN(BLN56),.WL(WL98));
sram_cell_6t_5 inst_cell_98_57 (.BL(BL57),.BLN(BLN57),.WL(WL98));
sram_cell_6t_5 inst_cell_98_58 (.BL(BL58),.BLN(BLN58),.WL(WL98));
sram_cell_6t_5 inst_cell_98_59 (.BL(BL59),.BLN(BLN59),.WL(WL98));
sram_cell_6t_5 inst_cell_98_60 (.BL(BL60),.BLN(BLN60),.WL(WL98));
sram_cell_6t_5 inst_cell_98_61 (.BL(BL61),.BLN(BLN61),.WL(WL98));
sram_cell_6t_5 inst_cell_98_62 (.BL(BL62),.BLN(BLN62),.WL(WL98));
sram_cell_6t_5 inst_cell_98_63 (.BL(BL63),.BLN(BLN63),.WL(WL98));
sram_cell_6t_5 inst_cell_98_64 (.BL(BL64),.BLN(BLN64),.WL(WL98));
sram_cell_6t_5 inst_cell_98_65 (.BL(BL65),.BLN(BLN65),.WL(WL98));
sram_cell_6t_5 inst_cell_98_66 (.BL(BL66),.BLN(BLN66),.WL(WL98));
sram_cell_6t_5 inst_cell_98_67 (.BL(BL67),.BLN(BLN67),.WL(WL98));
sram_cell_6t_5 inst_cell_98_68 (.BL(BL68),.BLN(BLN68),.WL(WL98));
sram_cell_6t_5 inst_cell_98_69 (.BL(BL69),.BLN(BLN69),.WL(WL98));
sram_cell_6t_5 inst_cell_98_70 (.BL(BL70),.BLN(BLN70),.WL(WL98));
sram_cell_6t_5 inst_cell_98_71 (.BL(BL71),.BLN(BLN71),.WL(WL98));
sram_cell_6t_5 inst_cell_98_72 (.BL(BL72),.BLN(BLN72),.WL(WL98));
sram_cell_6t_5 inst_cell_98_73 (.BL(BL73),.BLN(BLN73),.WL(WL98));
sram_cell_6t_5 inst_cell_98_74 (.BL(BL74),.BLN(BLN74),.WL(WL98));
sram_cell_6t_5 inst_cell_98_75 (.BL(BL75),.BLN(BLN75),.WL(WL98));
sram_cell_6t_5 inst_cell_98_76 (.BL(BL76),.BLN(BLN76),.WL(WL98));
sram_cell_6t_5 inst_cell_98_77 (.BL(BL77),.BLN(BLN77),.WL(WL98));
sram_cell_6t_5 inst_cell_98_78 (.BL(BL78),.BLN(BLN78),.WL(WL98));
sram_cell_6t_5 inst_cell_98_79 (.BL(BL79),.BLN(BLN79),.WL(WL98));
sram_cell_6t_5 inst_cell_98_80 (.BL(BL80),.BLN(BLN80),.WL(WL98));
sram_cell_6t_5 inst_cell_98_81 (.BL(BL81),.BLN(BLN81),.WL(WL98));
sram_cell_6t_5 inst_cell_98_82 (.BL(BL82),.BLN(BLN82),.WL(WL98));
sram_cell_6t_5 inst_cell_98_83 (.BL(BL83),.BLN(BLN83),.WL(WL98));
sram_cell_6t_5 inst_cell_98_84 (.BL(BL84),.BLN(BLN84),.WL(WL98));
sram_cell_6t_5 inst_cell_98_85 (.BL(BL85),.BLN(BLN85),.WL(WL98));
sram_cell_6t_5 inst_cell_98_86 (.BL(BL86),.BLN(BLN86),.WL(WL98));
sram_cell_6t_5 inst_cell_98_87 (.BL(BL87),.BLN(BLN87),.WL(WL98));
sram_cell_6t_5 inst_cell_98_88 (.BL(BL88),.BLN(BLN88),.WL(WL98));
sram_cell_6t_5 inst_cell_98_89 (.BL(BL89),.BLN(BLN89),.WL(WL98));
sram_cell_6t_5 inst_cell_98_90 (.BL(BL90),.BLN(BLN90),.WL(WL98));
sram_cell_6t_5 inst_cell_98_91 (.BL(BL91),.BLN(BLN91),.WL(WL98));
sram_cell_6t_5 inst_cell_98_92 (.BL(BL92),.BLN(BLN92),.WL(WL98));
sram_cell_6t_5 inst_cell_98_93 (.BL(BL93),.BLN(BLN93),.WL(WL98));
sram_cell_6t_5 inst_cell_98_94 (.BL(BL94),.BLN(BLN94),.WL(WL98));
sram_cell_6t_5 inst_cell_98_95 (.BL(BL95),.BLN(BLN95),.WL(WL98));
sram_cell_6t_5 inst_cell_98_96 (.BL(BL96),.BLN(BLN96),.WL(WL98));
sram_cell_6t_5 inst_cell_98_97 (.BL(BL97),.BLN(BLN97),.WL(WL98));
sram_cell_6t_5 inst_cell_98_98 (.BL(BL98),.BLN(BLN98),.WL(WL98));
sram_cell_6t_5 inst_cell_98_99 (.BL(BL99),.BLN(BLN99),.WL(WL98));
sram_cell_6t_5 inst_cell_98_100 (.BL(BL100),.BLN(BLN100),.WL(WL98));
sram_cell_6t_5 inst_cell_98_101 (.BL(BL101),.BLN(BLN101),.WL(WL98));
sram_cell_6t_5 inst_cell_98_102 (.BL(BL102),.BLN(BLN102),.WL(WL98));
sram_cell_6t_5 inst_cell_98_103 (.BL(BL103),.BLN(BLN103),.WL(WL98));
sram_cell_6t_5 inst_cell_98_104 (.BL(BL104),.BLN(BLN104),.WL(WL98));
sram_cell_6t_5 inst_cell_98_105 (.BL(BL105),.BLN(BLN105),.WL(WL98));
sram_cell_6t_5 inst_cell_98_106 (.BL(BL106),.BLN(BLN106),.WL(WL98));
sram_cell_6t_5 inst_cell_98_107 (.BL(BL107),.BLN(BLN107),.WL(WL98));
sram_cell_6t_5 inst_cell_98_108 (.BL(BL108),.BLN(BLN108),.WL(WL98));
sram_cell_6t_5 inst_cell_98_109 (.BL(BL109),.BLN(BLN109),.WL(WL98));
sram_cell_6t_5 inst_cell_98_110 (.BL(BL110),.BLN(BLN110),.WL(WL98));
sram_cell_6t_5 inst_cell_98_111 (.BL(BL111),.BLN(BLN111),.WL(WL98));
sram_cell_6t_5 inst_cell_98_112 (.BL(BL112),.BLN(BLN112),.WL(WL98));
sram_cell_6t_5 inst_cell_98_113 (.BL(BL113),.BLN(BLN113),.WL(WL98));
sram_cell_6t_5 inst_cell_98_114 (.BL(BL114),.BLN(BLN114),.WL(WL98));
sram_cell_6t_5 inst_cell_98_115 (.BL(BL115),.BLN(BLN115),.WL(WL98));
sram_cell_6t_5 inst_cell_98_116 (.BL(BL116),.BLN(BLN116),.WL(WL98));
sram_cell_6t_5 inst_cell_98_117 (.BL(BL117),.BLN(BLN117),.WL(WL98));
sram_cell_6t_5 inst_cell_98_118 (.BL(BL118),.BLN(BLN118),.WL(WL98));
sram_cell_6t_5 inst_cell_98_119 (.BL(BL119),.BLN(BLN119),.WL(WL98));
sram_cell_6t_5 inst_cell_98_120 (.BL(BL120),.BLN(BLN120),.WL(WL98));
sram_cell_6t_5 inst_cell_98_121 (.BL(BL121),.BLN(BLN121),.WL(WL98));
sram_cell_6t_5 inst_cell_98_122 (.BL(BL122),.BLN(BLN122),.WL(WL98));
sram_cell_6t_5 inst_cell_98_123 (.BL(BL123),.BLN(BLN123),.WL(WL98));
sram_cell_6t_5 inst_cell_98_124 (.BL(BL124),.BLN(BLN124),.WL(WL98));
sram_cell_6t_5 inst_cell_98_125 (.BL(BL125),.BLN(BLN125),.WL(WL98));
sram_cell_6t_5 inst_cell_98_126 (.BL(BL126),.BLN(BLN126),.WL(WL98));
sram_cell_6t_5 inst_cell_98_127 (.BL(BL127),.BLN(BLN127),.WL(WL98));
sram_cell_6t_5 inst_cell_99_0 (.BL(BL0),.BLN(BLN0),.WL(WL99));
sram_cell_6t_5 inst_cell_99_1 (.BL(BL1),.BLN(BLN1),.WL(WL99));
sram_cell_6t_5 inst_cell_99_2 (.BL(BL2),.BLN(BLN2),.WL(WL99));
sram_cell_6t_5 inst_cell_99_3 (.BL(BL3),.BLN(BLN3),.WL(WL99));
sram_cell_6t_5 inst_cell_99_4 (.BL(BL4),.BLN(BLN4),.WL(WL99));
sram_cell_6t_5 inst_cell_99_5 (.BL(BL5),.BLN(BLN5),.WL(WL99));
sram_cell_6t_5 inst_cell_99_6 (.BL(BL6),.BLN(BLN6),.WL(WL99));
sram_cell_6t_5 inst_cell_99_7 (.BL(BL7),.BLN(BLN7),.WL(WL99));
sram_cell_6t_5 inst_cell_99_8 (.BL(BL8),.BLN(BLN8),.WL(WL99));
sram_cell_6t_5 inst_cell_99_9 (.BL(BL9),.BLN(BLN9),.WL(WL99));
sram_cell_6t_5 inst_cell_99_10 (.BL(BL10),.BLN(BLN10),.WL(WL99));
sram_cell_6t_5 inst_cell_99_11 (.BL(BL11),.BLN(BLN11),.WL(WL99));
sram_cell_6t_5 inst_cell_99_12 (.BL(BL12),.BLN(BLN12),.WL(WL99));
sram_cell_6t_5 inst_cell_99_13 (.BL(BL13),.BLN(BLN13),.WL(WL99));
sram_cell_6t_5 inst_cell_99_14 (.BL(BL14),.BLN(BLN14),.WL(WL99));
sram_cell_6t_5 inst_cell_99_15 (.BL(BL15),.BLN(BLN15),.WL(WL99));
sram_cell_6t_5 inst_cell_99_16 (.BL(BL16),.BLN(BLN16),.WL(WL99));
sram_cell_6t_5 inst_cell_99_17 (.BL(BL17),.BLN(BLN17),.WL(WL99));
sram_cell_6t_5 inst_cell_99_18 (.BL(BL18),.BLN(BLN18),.WL(WL99));
sram_cell_6t_5 inst_cell_99_19 (.BL(BL19),.BLN(BLN19),.WL(WL99));
sram_cell_6t_5 inst_cell_99_20 (.BL(BL20),.BLN(BLN20),.WL(WL99));
sram_cell_6t_5 inst_cell_99_21 (.BL(BL21),.BLN(BLN21),.WL(WL99));
sram_cell_6t_5 inst_cell_99_22 (.BL(BL22),.BLN(BLN22),.WL(WL99));
sram_cell_6t_5 inst_cell_99_23 (.BL(BL23),.BLN(BLN23),.WL(WL99));
sram_cell_6t_5 inst_cell_99_24 (.BL(BL24),.BLN(BLN24),.WL(WL99));
sram_cell_6t_5 inst_cell_99_25 (.BL(BL25),.BLN(BLN25),.WL(WL99));
sram_cell_6t_5 inst_cell_99_26 (.BL(BL26),.BLN(BLN26),.WL(WL99));
sram_cell_6t_5 inst_cell_99_27 (.BL(BL27),.BLN(BLN27),.WL(WL99));
sram_cell_6t_5 inst_cell_99_28 (.BL(BL28),.BLN(BLN28),.WL(WL99));
sram_cell_6t_5 inst_cell_99_29 (.BL(BL29),.BLN(BLN29),.WL(WL99));
sram_cell_6t_5 inst_cell_99_30 (.BL(BL30),.BLN(BLN30),.WL(WL99));
sram_cell_6t_5 inst_cell_99_31 (.BL(BL31),.BLN(BLN31),.WL(WL99));
sram_cell_6t_5 inst_cell_99_32 (.BL(BL32),.BLN(BLN32),.WL(WL99));
sram_cell_6t_5 inst_cell_99_33 (.BL(BL33),.BLN(BLN33),.WL(WL99));
sram_cell_6t_5 inst_cell_99_34 (.BL(BL34),.BLN(BLN34),.WL(WL99));
sram_cell_6t_5 inst_cell_99_35 (.BL(BL35),.BLN(BLN35),.WL(WL99));
sram_cell_6t_5 inst_cell_99_36 (.BL(BL36),.BLN(BLN36),.WL(WL99));
sram_cell_6t_5 inst_cell_99_37 (.BL(BL37),.BLN(BLN37),.WL(WL99));
sram_cell_6t_5 inst_cell_99_38 (.BL(BL38),.BLN(BLN38),.WL(WL99));
sram_cell_6t_5 inst_cell_99_39 (.BL(BL39),.BLN(BLN39),.WL(WL99));
sram_cell_6t_5 inst_cell_99_40 (.BL(BL40),.BLN(BLN40),.WL(WL99));
sram_cell_6t_5 inst_cell_99_41 (.BL(BL41),.BLN(BLN41),.WL(WL99));
sram_cell_6t_5 inst_cell_99_42 (.BL(BL42),.BLN(BLN42),.WL(WL99));
sram_cell_6t_5 inst_cell_99_43 (.BL(BL43),.BLN(BLN43),.WL(WL99));
sram_cell_6t_5 inst_cell_99_44 (.BL(BL44),.BLN(BLN44),.WL(WL99));
sram_cell_6t_5 inst_cell_99_45 (.BL(BL45),.BLN(BLN45),.WL(WL99));
sram_cell_6t_5 inst_cell_99_46 (.BL(BL46),.BLN(BLN46),.WL(WL99));
sram_cell_6t_5 inst_cell_99_47 (.BL(BL47),.BLN(BLN47),.WL(WL99));
sram_cell_6t_5 inst_cell_99_48 (.BL(BL48),.BLN(BLN48),.WL(WL99));
sram_cell_6t_5 inst_cell_99_49 (.BL(BL49),.BLN(BLN49),.WL(WL99));
sram_cell_6t_5 inst_cell_99_50 (.BL(BL50),.BLN(BLN50),.WL(WL99));
sram_cell_6t_5 inst_cell_99_51 (.BL(BL51),.BLN(BLN51),.WL(WL99));
sram_cell_6t_5 inst_cell_99_52 (.BL(BL52),.BLN(BLN52),.WL(WL99));
sram_cell_6t_5 inst_cell_99_53 (.BL(BL53),.BLN(BLN53),.WL(WL99));
sram_cell_6t_5 inst_cell_99_54 (.BL(BL54),.BLN(BLN54),.WL(WL99));
sram_cell_6t_5 inst_cell_99_55 (.BL(BL55),.BLN(BLN55),.WL(WL99));
sram_cell_6t_5 inst_cell_99_56 (.BL(BL56),.BLN(BLN56),.WL(WL99));
sram_cell_6t_5 inst_cell_99_57 (.BL(BL57),.BLN(BLN57),.WL(WL99));
sram_cell_6t_5 inst_cell_99_58 (.BL(BL58),.BLN(BLN58),.WL(WL99));
sram_cell_6t_5 inst_cell_99_59 (.BL(BL59),.BLN(BLN59),.WL(WL99));
sram_cell_6t_5 inst_cell_99_60 (.BL(BL60),.BLN(BLN60),.WL(WL99));
sram_cell_6t_5 inst_cell_99_61 (.BL(BL61),.BLN(BLN61),.WL(WL99));
sram_cell_6t_5 inst_cell_99_62 (.BL(BL62),.BLN(BLN62),.WL(WL99));
sram_cell_6t_5 inst_cell_99_63 (.BL(BL63),.BLN(BLN63),.WL(WL99));
sram_cell_6t_5 inst_cell_99_64 (.BL(BL64),.BLN(BLN64),.WL(WL99));
sram_cell_6t_5 inst_cell_99_65 (.BL(BL65),.BLN(BLN65),.WL(WL99));
sram_cell_6t_5 inst_cell_99_66 (.BL(BL66),.BLN(BLN66),.WL(WL99));
sram_cell_6t_5 inst_cell_99_67 (.BL(BL67),.BLN(BLN67),.WL(WL99));
sram_cell_6t_5 inst_cell_99_68 (.BL(BL68),.BLN(BLN68),.WL(WL99));
sram_cell_6t_5 inst_cell_99_69 (.BL(BL69),.BLN(BLN69),.WL(WL99));
sram_cell_6t_5 inst_cell_99_70 (.BL(BL70),.BLN(BLN70),.WL(WL99));
sram_cell_6t_5 inst_cell_99_71 (.BL(BL71),.BLN(BLN71),.WL(WL99));
sram_cell_6t_5 inst_cell_99_72 (.BL(BL72),.BLN(BLN72),.WL(WL99));
sram_cell_6t_5 inst_cell_99_73 (.BL(BL73),.BLN(BLN73),.WL(WL99));
sram_cell_6t_5 inst_cell_99_74 (.BL(BL74),.BLN(BLN74),.WL(WL99));
sram_cell_6t_5 inst_cell_99_75 (.BL(BL75),.BLN(BLN75),.WL(WL99));
sram_cell_6t_5 inst_cell_99_76 (.BL(BL76),.BLN(BLN76),.WL(WL99));
sram_cell_6t_5 inst_cell_99_77 (.BL(BL77),.BLN(BLN77),.WL(WL99));
sram_cell_6t_5 inst_cell_99_78 (.BL(BL78),.BLN(BLN78),.WL(WL99));
sram_cell_6t_5 inst_cell_99_79 (.BL(BL79),.BLN(BLN79),.WL(WL99));
sram_cell_6t_5 inst_cell_99_80 (.BL(BL80),.BLN(BLN80),.WL(WL99));
sram_cell_6t_5 inst_cell_99_81 (.BL(BL81),.BLN(BLN81),.WL(WL99));
sram_cell_6t_5 inst_cell_99_82 (.BL(BL82),.BLN(BLN82),.WL(WL99));
sram_cell_6t_5 inst_cell_99_83 (.BL(BL83),.BLN(BLN83),.WL(WL99));
sram_cell_6t_5 inst_cell_99_84 (.BL(BL84),.BLN(BLN84),.WL(WL99));
sram_cell_6t_5 inst_cell_99_85 (.BL(BL85),.BLN(BLN85),.WL(WL99));
sram_cell_6t_5 inst_cell_99_86 (.BL(BL86),.BLN(BLN86),.WL(WL99));
sram_cell_6t_5 inst_cell_99_87 (.BL(BL87),.BLN(BLN87),.WL(WL99));
sram_cell_6t_5 inst_cell_99_88 (.BL(BL88),.BLN(BLN88),.WL(WL99));
sram_cell_6t_5 inst_cell_99_89 (.BL(BL89),.BLN(BLN89),.WL(WL99));
sram_cell_6t_5 inst_cell_99_90 (.BL(BL90),.BLN(BLN90),.WL(WL99));
sram_cell_6t_5 inst_cell_99_91 (.BL(BL91),.BLN(BLN91),.WL(WL99));
sram_cell_6t_5 inst_cell_99_92 (.BL(BL92),.BLN(BLN92),.WL(WL99));
sram_cell_6t_5 inst_cell_99_93 (.BL(BL93),.BLN(BLN93),.WL(WL99));
sram_cell_6t_5 inst_cell_99_94 (.BL(BL94),.BLN(BLN94),.WL(WL99));
sram_cell_6t_5 inst_cell_99_95 (.BL(BL95),.BLN(BLN95),.WL(WL99));
sram_cell_6t_5 inst_cell_99_96 (.BL(BL96),.BLN(BLN96),.WL(WL99));
sram_cell_6t_5 inst_cell_99_97 (.BL(BL97),.BLN(BLN97),.WL(WL99));
sram_cell_6t_5 inst_cell_99_98 (.BL(BL98),.BLN(BLN98),.WL(WL99));
sram_cell_6t_5 inst_cell_99_99 (.BL(BL99),.BLN(BLN99),.WL(WL99));
sram_cell_6t_5 inst_cell_99_100 (.BL(BL100),.BLN(BLN100),.WL(WL99));
sram_cell_6t_5 inst_cell_99_101 (.BL(BL101),.BLN(BLN101),.WL(WL99));
sram_cell_6t_5 inst_cell_99_102 (.BL(BL102),.BLN(BLN102),.WL(WL99));
sram_cell_6t_5 inst_cell_99_103 (.BL(BL103),.BLN(BLN103),.WL(WL99));
sram_cell_6t_5 inst_cell_99_104 (.BL(BL104),.BLN(BLN104),.WL(WL99));
sram_cell_6t_5 inst_cell_99_105 (.BL(BL105),.BLN(BLN105),.WL(WL99));
sram_cell_6t_5 inst_cell_99_106 (.BL(BL106),.BLN(BLN106),.WL(WL99));
sram_cell_6t_5 inst_cell_99_107 (.BL(BL107),.BLN(BLN107),.WL(WL99));
sram_cell_6t_5 inst_cell_99_108 (.BL(BL108),.BLN(BLN108),.WL(WL99));
sram_cell_6t_5 inst_cell_99_109 (.BL(BL109),.BLN(BLN109),.WL(WL99));
sram_cell_6t_5 inst_cell_99_110 (.BL(BL110),.BLN(BLN110),.WL(WL99));
sram_cell_6t_5 inst_cell_99_111 (.BL(BL111),.BLN(BLN111),.WL(WL99));
sram_cell_6t_5 inst_cell_99_112 (.BL(BL112),.BLN(BLN112),.WL(WL99));
sram_cell_6t_5 inst_cell_99_113 (.BL(BL113),.BLN(BLN113),.WL(WL99));
sram_cell_6t_5 inst_cell_99_114 (.BL(BL114),.BLN(BLN114),.WL(WL99));
sram_cell_6t_5 inst_cell_99_115 (.BL(BL115),.BLN(BLN115),.WL(WL99));
sram_cell_6t_5 inst_cell_99_116 (.BL(BL116),.BLN(BLN116),.WL(WL99));
sram_cell_6t_5 inst_cell_99_117 (.BL(BL117),.BLN(BLN117),.WL(WL99));
sram_cell_6t_5 inst_cell_99_118 (.BL(BL118),.BLN(BLN118),.WL(WL99));
sram_cell_6t_5 inst_cell_99_119 (.BL(BL119),.BLN(BLN119),.WL(WL99));
sram_cell_6t_5 inst_cell_99_120 (.BL(BL120),.BLN(BLN120),.WL(WL99));
sram_cell_6t_5 inst_cell_99_121 (.BL(BL121),.BLN(BLN121),.WL(WL99));
sram_cell_6t_5 inst_cell_99_122 (.BL(BL122),.BLN(BLN122),.WL(WL99));
sram_cell_6t_5 inst_cell_99_123 (.BL(BL123),.BLN(BLN123),.WL(WL99));
sram_cell_6t_5 inst_cell_99_124 (.BL(BL124),.BLN(BLN124),.WL(WL99));
sram_cell_6t_5 inst_cell_99_125 (.BL(BL125),.BLN(BLN125),.WL(WL99));
sram_cell_6t_5 inst_cell_99_126 (.BL(BL126),.BLN(BLN126),.WL(WL99));
sram_cell_6t_5 inst_cell_99_127 (.BL(BL127),.BLN(BLN127),.WL(WL99));
sram_cell_6t_5 inst_cell_100_0 (.BL(BL0),.BLN(BLN0),.WL(WL100));
sram_cell_6t_5 inst_cell_100_1 (.BL(BL1),.BLN(BLN1),.WL(WL100));
sram_cell_6t_5 inst_cell_100_2 (.BL(BL2),.BLN(BLN2),.WL(WL100));
sram_cell_6t_5 inst_cell_100_3 (.BL(BL3),.BLN(BLN3),.WL(WL100));
sram_cell_6t_5 inst_cell_100_4 (.BL(BL4),.BLN(BLN4),.WL(WL100));
sram_cell_6t_5 inst_cell_100_5 (.BL(BL5),.BLN(BLN5),.WL(WL100));
sram_cell_6t_5 inst_cell_100_6 (.BL(BL6),.BLN(BLN6),.WL(WL100));
sram_cell_6t_5 inst_cell_100_7 (.BL(BL7),.BLN(BLN7),.WL(WL100));
sram_cell_6t_5 inst_cell_100_8 (.BL(BL8),.BLN(BLN8),.WL(WL100));
sram_cell_6t_5 inst_cell_100_9 (.BL(BL9),.BLN(BLN9),.WL(WL100));
sram_cell_6t_5 inst_cell_100_10 (.BL(BL10),.BLN(BLN10),.WL(WL100));
sram_cell_6t_5 inst_cell_100_11 (.BL(BL11),.BLN(BLN11),.WL(WL100));
sram_cell_6t_5 inst_cell_100_12 (.BL(BL12),.BLN(BLN12),.WL(WL100));
sram_cell_6t_5 inst_cell_100_13 (.BL(BL13),.BLN(BLN13),.WL(WL100));
sram_cell_6t_5 inst_cell_100_14 (.BL(BL14),.BLN(BLN14),.WL(WL100));
sram_cell_6t_5 inst_cell_100_15 (.BL(BL15),.BLN(BLN15),.WL(WL100));
sram_cell_6t_5 inst_cell_100_16 (.BL(BL16),.BLN(BLN16),.WL(WL100));
sram_cell_6t_5 inst_cell_100_17 (.BL(BL17),.BLN(BLN17),.WL(WL100));
sram_cell_6t_5 inst_cell_100_18 (.BL(BL18),.BLN(BLN18),.WL(WL100));
sram_cell_6t_5 inst_cell_100_19 (.BL(BL19),.BLN(BLN19),.WL(WL100));
sram_cell_6t_5 inst_cell_100_20 (.BL(BL20),.BLN(BLN20),.WL(WL100));
sram_cell_6t_5 inst_cell_100_21 (.BL(BL21),.BLN(BLN21),.WL(WL100));
sram_cell_6t_5 inst_cell_100_22 (.BL(BL22),.BLN(BLN22),.WL(WL100));
sram_cell_6t_5 inst_cell_100_23 (.BL(BL23),.BLN(BLN23),.WL(WL100));
sram_cell_6t_5 inst_cell_100_24 (.BL(BL24),.BLN(BLN24),.WL(WL100));
sram_cell_6t_5 inst_cell_100_25 (.BL(BL25),.BLN(BLN25),.WL(WL100));
sram_cell_6t_5 inst_cell_100_26 (.BL(BL26),.BLN(BLN26),.WL(WL100));
sram_cell_6t_5 inst_cell_100_27 (.BL(BL27),.BLN(BLN27),.WL(WL100));
sram_cell_6t_5 inst_cell_100_28 (.BL(BL28),.BLN(BLN28),.WL(WL100));
sram_cell_6t_5 inst_cell_100_29 (.BL(BL29),.BLN(BLN29),.WL(WL100));
sram_cell_6t_5 inst_cell_100_30 (.BL(BL30),.BLN(BLN30),.WL(WL100));
sram_cell_6t_5 inst_cell_100_31 (.BL(BL31),.BLN(BLN31),.WL(WL100));
sram_cell_6t_5 inst_cell_100_32 (.BL(BL32),.BLN(BLN32),.WL(WL100));
sram_cell_6t_5 inst_cell_100_33 (.BL(BL33),.BLN(BLN33),.WL(WL100));
sram_cell_6t_5 inst_cell_100_34 (.BL(BL34),.BLN(BLN34),.WL(WL100));
sram_cell_6t_5 inst_cell_100_35 (.BL(BL35),.BLN(BLN35),.WL(WL100));
sram_cell_6t_5 inst_cell_100_36 (.BL(BL36),.BLN(BLN36),.WL(WL100));
sram_cell_6t_5 inst_cell_100_37 (.BL(BL37),.BLN(BLN37),.WL(WL100));
sram_cell_6t_5 inst_cell_100_38 (.BL(BL38),.BLN(BLN38),.WL(WL100));
sram_cell_6t_5 inst_cell_100_39 (.BL(BL39),.BLN(BLN39),.WL(WL100));
sram_cell_6t_5 inst_cell_100_40 (.BL(BL40),.BLN(BLN40),.WL(WL100));
sram_cell_6t_5 inst_cell_100_41 (.BL(BL41),.BLN(BLN41),.WL(WL100));
sram_cell_6t_5 inst_cell_100_42 (.BL(BL42),.BLN(BLN42),.WL(WL100));
sram_cell_6t_5 inst_cell_100_43 (.BL(BL43),.BLN(BLN43),.WL(WL100));
sram_cell_6t_5 inst_cell_100_44 (.BL(BL44),.BLN(BLN44),.WL(WL100));
sram_cell_6t_5 inst_cell_100_45 (.BL(BL45),.BLN(BLN45),.WL(WL100));
sram_cell_6t_5 inst_cell_100_46 (.BL(BL46),.BLN(BLN46),.WL(WL100));
sram_cell_6t_5 inst_cell_100_47 (.BL(BL47),.BLN(BLN47),.WL(WL100));
sram_cell_6t_5 inst_cell_100_48 (.BL(BL48),.BLN(BLN48),.WL(WL100));
sram_cell_6t_5 inst_cell_100_49 (.BL(BL49),.BLN(BLN49),.WL(WL100));
sram_cell_6t_5 inst_cell_100_50 (.BL(BL50),.BLN(BLN50),.WL(WL100));
sram_cell_6t_5 inst_cell_100_51 (.BL(BL51),.BLN(BLN51),.WL(WL100));
sram_cell_6t_5 inst_cell_100_52 (.BL(BL52),.BLN(BLN52),.WL(WL100));
sram_cell_6t_5 inst_cell_100_53 (.BL(BL53),.BLN(BLN53),.WL(WL100));
sram_cell_6t_5 inst_cell_100_54 (.BL(BL54),.BLN(BLN54),.WL(WL100));
sram_cell_6t_5 inst_cell_100_55 (.BL(BL55),.BLN(BLN55),.WL(WL100));
sram_cell_6t_5 inst_cell_100_56 (.BL(BL56),.BLN(BLN56),.WL(WL100));
sram_cell_6t_5 inst_cell_100_57 (.BL(BL57),.BLN(BLN57),.WL(WL100));
sram_cell_6t_5 inst_cell_100_58 (.BL(BL58),.BLN(BLN58),.WL(WL100));
sram_cell_6t_5 inst_cell_100_59 (.BL(BL59),.BLN(BLN59),.WL(WL100));
sram_cell_6t_5 inst_cell_100_60 (.BL(BL60),.BLN(BLN60),.WL(WL100));
sram_cell_6t_5 inst_cell_100_61 (.BL(BL61),.BLN(BLN61),.WL(WL100));
sram_cell_6t_5 inst_cell_100_62 (.BL(BL62),.BLN(BLN62),.WL(WL100));
sram_cell_6t_5 inst_cell_100_63 (.BL(BL63),.BLN(BLN63),.WL(WL100));
sram_cell_6t_5 inst_cell_100_64 (.BL(BL64),.BLN(BLN64),.WL(WL100));
sram_cell_6t_5 inst_cell_100_65 (.BL(BL65),.BLN(BLN65),.WL(WL100));
sram_cell_6t_5 inst_cell_100_66 (.BL(BL66),.BLN(BLN66),.WL(WL100));
sram_cell_6t_5 inst_cell_100_67 (.BL(BL67),.BLN(BLN67),.WL(WL100));
sram_cell_6t_5 inst_cell_100_68 (.BL(BL68),.BLN(BLN68),.WL(WL100));
sram_cell_6t_5 inst_cell_100_69 (.BL(BL69),.BLN(BLN69),.WL(WL100));
sram_cell_6t_5 inst_cell_100_70 (.BL(BL70),.BLN(BLN70),.WL(WL100));
sram_cell_6t_5 inst_cell_100_71 (.BL(BL71),.BLN(BLN71),.WL(WL100));
sram_cell_6t_5 inst_cell_100_72 (.BL(BL72),.BLN(BLN72),.WL(WL100));
sram_cell_6t_5 inst_cell_100_73 (.BL(BL73),.BLN(BLN73),.WL(WL100));
sram_cell_6t_5 inst_cell_100_74 (.BL(BL74),.BLN(BLN74),.WL(WL100));
sram_cell_6t_5 inst_cell_100_75 (.BL(BL75),.BLN(BLN75),.WL(WL100));
sram_cell_6t_5 inst_cell_100_76 (.BL(BL76),.BLN(BLN76),.WL(WL100));
sram_cell_6t_5 inst_cell_100_77 (.BL(BL77),.BLN(BLN77),.WL(WL100));
sram_cell_6t_5 inst_cell_100_78 (.BL(BL78),.BLN(BLN78),.WL(WL100));
sram_cell_6t_5 inst_cell_100_79 (.BL(BL79),.BLN(BLN79),.WL(WL100));
sram_cell_6t_5 inst_cell_100_80 (.BL(BL80),.BLN(BLN80),.WL(WL100));
sram_cell_6t_5 inst_cell_100_81 (.BL(BL81),.BLN(BLN81),.WL(WL100));
sram_cell_6t_5 inst_cell_100_82 (.BL(BL82),.BLN(BLN82),.WL(WL100));
sram_cell_6t_5 inst_cell_100_83 (.BL(BL83),.BLN(BLN83),.WL(WL100));
sram_cell_6t_5 inst_cell_100_84 (.BL(BL84),.BLN(BLN84),.WL(WL100));
sram_cell_6t_5 inst_cell_100_85 (.BL(BL85),.BLN(BLN85),.WL(WL100));
sram_cell_6t_5 inst_cell_100_86 (.BL(BL86),.BLN(BLN86),.WL(WL100));
sram_cell_6t_5 inst_cell_100_87 (.BL(BL87),.BLN(BLN87),.WL(WL100));
sram_cell_6t_5 inst_cell_100_88 (.BL(BL88),.BLN(BLN88),.WL(WL100));
sram_cell_6t_5 inst_cell_100_89 (.BL(BL89),.BLN(BLN89),.WL(WL100));
sram_cell_6t_5 inst_cell_100_90 (.BL(BL90),.BLN(BLN90),.WL(WL100));
sram_cell_6t_5 inst_cell_100_91 (.BL(BL91),.BLN(BLN91),.WL(WL100));
sram_cell_6t_5 inst_cell_100_92 (.BL(BL92),.BLN(BLN92),.WL(WL100));
sram_cell_6t_5 inst_cell_100_93 (.BL(BL93),.BLN(BLN93),.WL(WL100));
sram_cell_6t_5 inst_cell_100_94 (.BL(BL94),.BLN(BLN94),.WL(WL100));
sram_cell_6t_5 inst_cell_100_95 (.BL(BL95),.BLN(BLN95),.WL(WL100));
sram_cell_6t_5 inst_cell_100_96 (.BL(BL96),.BLN(BLN96),.WL(WL100));
sram_cell_6t_5 inst_cell_100_97 (.BL(BL97),.BLN(BLN97),.WL(WL100));
sram_cell_6t_5 inst_cell_100_98 (.BL(BL98),.BLN(BLN98),.WL(WL100));
sram_cell_6t_5 inst_cell_100_99 (.BL(BL99),.BLN(BLN99),.WL(WL100));
sram_cell_6t_5 inst_cell_100_100 (.BL(BL100),.BLN(BLN100),.WL(WL100));
sram_cell_6t_5 inst_cell_100_101 (.BL(BL101),.BLN(BLN101),.WL(WL100));
sram_cell_6t_5 inst_cell_100_102 (.BL(BL102),.BLN(BLN102),.WL(WL100));
sram_cell_6t_5 inst_cell_100_103 (.BL(BL103),.BLN(BLN103),.WL(WL100));
sram_cell_6t_5 inst_cell_100_104 (.BL(BL104),.BLN(BLN104),.WL(WL100));
sram_cell_6t_5 inst_cell_100_105 (.BL(BL105),.BLN(BLN105),.WL(WL100));
sram_cell_6t_5 inst_cell_100_106 (.BL(BL106),.BLN(BLN106),.WL(WL100));
sram_cell_6t_5 inst_cell_100_107 (.BL(BL107),.BLN(BLN107),.WL(WL100));
sram_cell_6t_5 inst_cell_100_108 (.BL(BL108),.BLN(BLN108),.WL(WL100));
sram_cell_6t_5 inst_cell_100_109 (.BL(BL109),.BLN(BLN109),.WL(WL100));
sram_cell_6t_5 inst_cell_100_110 (.BL(BL110),.BLN(BLN110),.WL(WL100));
sram_cell_6t_5 inst_cell_100_111 (.BL(BL111),.BLN(BLN111),.WL(WL100));
sram_cell_6t_5 inst_cell_100_112 (.BL(BL112),.BLN(BLN112),.WL(WL100));
sram_cell_6t_5 inst_cell_100_113 (.BL(BL113),.BLN(BLN113),.WL(WL100));
sram_cell_6t_5 inst_cell_100_114 (.BL(BL114),.BLN(BLN114),.WL(WL100));
sram_cell_6t_5 inst_cell_100_115 (.BL(BL115),.BLN(BLN115),.WL(WL100));
sram_cell_6t_5 inst_cell_100_116 (.BL(BL116),.BLN(BLN116),.WL(WL100));
sram_cell_6t_5 inst_cell_100_117 (.BL(BL117),.BLN(BLN117),.WL(WL100));
sram_cell_6t_5 inst_cell_100_118 (.BL(BL118),.BLN(BLN118),.WL(WL100));
sram_cell_6t_5 inst_cell_100_119 (.BL(BL119),.BLN(BLN119),.WL(WL100));
sram_cell_6t_5 inst_cell_100_120 (.BL(BL120),.BLN(BLN120),.WL(WL100));
sram_cell_6t_5 inst_cell_100_121 (.BL(BL121),.BLN(BLN121),.WL(WL100));
sram_cell_6t_5 inst_cell_100_122 (.BL(BL122),.BLN(BLN122),.WL(WL100));
sram_cell_6t_5 inst_cell_100_123 (.BL(BL123),.BLN(BLN123),.WL(WL100));
sram_cell_6t_5 inst_cell_100_124 (.BL(BL124),.BLN(BLN124),.WL(WL100));
sram_cell_6t_5 inst_cell_100_125 (.BL(BL125),.BLN(BLN125),.WL(WL100));
sram_cell_6t_5 inst_cell_100_126 (.BL(BL126),.BLN(BLN126),.WL(WL100));
sram_cell_6t_5 inst_cell_100_127 (.BL(BL127),.BLN(BLN127),.WL(WL100));
sram_cell_6t_5 inst_cell_101_0 (.BL(BL0),.BLN(BLN0),.WL(WL101));
sram_cell_6t_5 inst_cell_101_1 (.BL(BL1),.BLN(BLN1),.WL(WL101));
sram_cell_6t_5 inst_cell_101_2 (.BL(BL2),.BLN(BLN2),.WL(WL101));
sram_cell_6t_5 inst_cell_101_3 (.BL(BL3),.BLN(BLN3),.WL(WL101));
sram_cell_6t_5 inst_cell_101_4 (.BL(BL4),.BLN(BLN4),.WL(WL101));
sram_cell_6t_5 inst_cell_101_5 (.BL(BL5),.BLN(BLN5),.WL(WL101));
sram_cell_6t_5 inst_cell_101_6 (.BL(BL6),.BLN(BLN6),.WL(WL101));
sram_cell_6t_5 inst_cell_101_7 (.BL(BL7),.BLN(BLN7),.WL(WL101));
sram_cell_6t_5 inst_cell_101_8 (.BL(BL8),.BLN(BLN8),.WL(WL101));
sram_cell_6t_5 inst_cell_101_9 (.BL(BL9),.BLN(BLN9),.WL(WL101));
sram_cell_6t_5 inst_cell_101_10 (.BL(BL10),.BLN(BLN10),.WL(WL101));
sram_cell_6t_5 inst_cell_101_11 (.BL(BL11),.BLN(BLN11),.WL(WL101));
sram_cell_6t_5 inst_cell_101_12 (.BL(BL12),.BLN(BLN12),.WL(WL101));
sram_cell_6t_5 inst_cell_101_13 (.BL(BL13),.BLN(BLN13),.WL(WL101));
sram_cell_6t_5 inst_cell_101_14 (.BL(BL14),.BLN(BLN14),.WL(WL101));
sram_cell_6t_5 inst_cell_101_15 (.BL(BL15),.BLN(BLN15),.WL(WL101));
sram_cell_6t_5 inst_cell_101_16 (.BL(BL16),.BLN(BLN16),.WL(WL101));
sram_cell_6t_5 inst_cell_101_17 (.BL(BL17),.BLN(BLN17),.WL(WL101));
sram_cell_6t_5 inst_cell_101_18 (.BL(BL18),.BLN(BLN18),.WL(WL101));
sram_cell_6t_5 inst_cell_101_19 (.BL(BL19),.BLN(BLN19),.WL(WL101));
sram_cell_6t_5 inst_cell_101_20 (.BL(BL20),.BLN(BLN20),.WL(WL101));
sram_cell_6t_5 inst_cell_101_21 (.BL(BL21),.BLN(BLN21),.WL(WL101));
sram_cell_6t_5 inst_cell_101_22 (.BL(BL22),.BLN(BLN22),.WL(WL101));
sram_cell_6t_5 inst_cell_101_23 (.BL(BL23),.BLN(BLN23),.WL(WL101));
sram_cell_6t_5 inst_cell_101_24 (.BL(BL24),.BLN(BLN24),.WL(WL101));
sram_cell_6t_5 inst_cell_101_25 (.BL(BL25),.BLN(BLN25),.WL(WL101));
sram_cell_6t_5 inst_cell_101_26 (.BL(BL26),.BLN(BLN26),.WL(WL101));
sram_cell_6t_5 inst_cell_101_27 (.BL(BL27),.BLN(BLN27),.WL(WL101));
sram_cell_6t_5 inst_cell_101_28 (.BL(BL28),.BLN(BLN28),.WL(WL101));
sram_cell_6t_5 inst_cell_101_29 (.BL(BL29),.BLN(BLN29),.WL(WL101));
sram_cell_6t_5 inst_cell_101_30 (.BL(BL30),.BLN(BLN30),.WL(WL101));
sram_cell_6t_5 inst_cell_101_31 (.BL(BL31),.BLN(BLN31),.WL(WL101));
sram_cell_6t_5 inst_cell_101_32 (.BL(BL32),.BLN(BLN32),.WL(WL101));
sram_cell_6t_5 inst_cell_101_33 (.BL(BL33),.BLN(BLN33),.WL(WL101));
sram_cell_6t_5 inst_cell_101_34 (.BL(BL34),.BLN(BLN34),.WL(WL101));
sram_cell_6t_5 inst_cell_101_35 (.BL(BL35),.BLN(BLN35),.WL(WL101));
sram_cell_6t_5 inst_cell_101_36 (.BL(BL36),.BLN(BLN36),.WL(WL101));
sram_cell_6t_5 inst_cell_101_37 (.BL(BL37),.BLN(BLN37),.WL(WL101));
sram_cell_6t_5 inst_cell_101_38 (.BL(BL38),.BLN(BLN38),.WL(WL101));
sram_cell_6t_5 inst_cell_101_39 (.BL(BL39),.BLN(BLN39),.WL(WL101));
sram_cell_6t_5 inst_cell_101_40 (.BL(BL40),.BLN(BLN40),.WL(WL101));
sram_cell_6t_5 inst_cell_101_41 (.BL(BL41),.BLN(BLN41),.WL(WL101));
sram_cell_6t_5 inst_cell_101_42 (.BL(BL42),.BLN(BLN42),.WL(WL101));
sram_cell_6t_5 inst_cell_101_43 (.BL(BL43),.BLN(BLN43),.WL(WL101));
sram_cell_6t_5 inst_cell_101_44 (.BL(BL44),.BLN(BLN44),.WL(WL101));
sram_cell_6t_5 inst_cell_101_45 (.BL(BL45),.BLN(BLN45),.WL(WL101));
sram_cell_6t_5 inst_cell_101_46 (.BL(BL46),.BLN(BLN46),.WL(WL101));
sram_cell_6t_5 inst_cell_101_47 (.BL(BL47),.BLN(BLN47),.WL(WL101));
sram_cell_6t_5 inst_cell_101_48 (.BL(BL48),.BLN(BLN48),.WL(WL101));
sram_cell_6t_5 inst_cell_101_49 (.BL(BL49),.BLN(BLN49),.WL(WL101));
sram_cell_6t_5 inst_cell_101_50 (.BL(BL50),.BLN(BLN50),.WL(WL101));
sram_cell_6t_5 inst_cell_101_51 (.BL(BL51),.BLN(BLN51),.WL(WL101));
sram_cell_6t_5 inst_cell_101_52 (.BL(BL52),.BLN(BLN52),.WL(WL101));
sram_cell_6t_5 inst_cell_101_53 (.BL(BL53),.BLN(BLN53),.WL(WL101));
sram_cell_6t_5 inst_cell_101_54 (.BL(BL54),.BLN(BLN54),.WL(WL101));
sram_cell_6t_5 inst_cell_101_55 (.BL(BL55),.BLN(BLN55),.WL(WL101));
sram_cell_6t_5 inst_cell_101_56 (.BL(BL56),.BLN(BLN56),.WL(WL101));
sram_cell_6t_5 inst_cell_101_57 (.BL(BL57),.BLN(BLN57),.WL(WL101));
sram_cell_6t_5 inst_cell_101_58 (.BL(BL58),.BLN(BLN58),.WL(WL101));
sram_cell_6t_5 inst_cell_101_59 (.BL(BL59),.BLN(BLN59),.WL(WL101));
sram_cell_6t_5 inst_cell_101_60 (.BL(BL60),.BLN(BLN60),.WL(WL101));
sram_cell_6t_5 inst_cell_101_61 (.BL(BL61),.BLN(BLN61),.WL(WL101));
sram_cell_6t_5 inst_cell_101_62 (.BL(BL62),.BLN(BLN62),.WL(WL101));
sram_cell_6t_5 inst_cell_101_63 (.BL(BL63),.BLN(BLN63),.WL(WL101));
sram_cell_6t_5 inst_cell_101_64 (.BL(BL64),.BLN(BLN64),.WL(WL101));
sram_cell_6t_5 inst_cell_101_65 (.BL(BL65),.BLN(BLN65),.WL(WL101));
sram_cell_6t_5 inst_cell_101_66 (.BL(BL66),.BLN(BLN66),.WL(WL101));
sram_cell_6t_5 inst_cell_101_67 (.BL(BL67),.BLN(BLN67),.WL(WL101));
sram_cell_6t_5 inst_cell_101_68 (.BL(BL68),.BLN(BLN68),.WL(WL101));
sram_cell_6t_5 inst_cell_101_69 (.BL(BL69),.BLN(BLN69),.WL(WL101));
sram_cell_6t_5 inst_cell_101_70 (.BL(BL70),.BLN(BLN70),.WL(WL101));
sram_cell_6t_5 inst_cell_101_71 (.BL(BL71),.BLN(BLN71),.WL(WL101));
sram_cell_6t_5 inst_cell_101_72 (.BL(BL72),.BLN(BLN72),.WL(WL101));
sram_cell_6t_5 inst_cell_101_73 (.BL(BL73),.BLN(BLN73),.WL(WL101));
sram_cell_6t_5 inst_cell_101_74 (.BL(BL74),.BLN(BLN74),.WL(WL101));
sram_cell_6t_5 inst_cell_101_75 (.BL(BL75),.BLN(BLN75),.WL(WL101));
sram_cell_6t_5 inst_cell_101_76 (.BL(BL76),.BLN(BLN76),.WL(WL101));
sram_cell_6t_5 inst_cell_101_77 (.BL(BL77),.BLN(BLN77),.WL(WL101));
sram_cell_6t_5 inst_cell_101_78 (.BL(BL78),.BLN(BLN78),.WL(WL101));
sram_cell_6t_5 inst_cell_101_79 (.BL(BL79),.BLN(BLN79),.WL(WL101));
sram_cell_6t_5 inst_cell_101_80 (.BL(BL80),.BLN(BLN80),.WL(WL101));
sram_cell_6t_5 inst_cell_101_81 (.BL(BL81),.BLN(BLN81),.WL(WL101));
sram_cell_6t_5 inst_cell_101_82 (.BL(BL82),.BLN(BLN82),.WL(WL101));
sram_cell_6t_5 inst_cell_101_83 (.BL(BL83),.BLN(BLN83),.WL(WL101));
sram_cell_6t_5 inst_cell_101_84 (.BL(BL84),.BLN(BLN84),.WL(WL101));
sram_cell_6t_5 inst_cell_101_85 (.BL(BL85),.BLN(BLN85),.WL(WL101));
sram_cell_6t_5 inst_cell_101_86 (.BL(BL86),.BLN(BLN86),.WL(WL101));
sram_cell_6t_5 inst_cell_101_87 (.BL(BL87),.BLN(BLN87),.WL(WL101));
sram_cell_6t_5 inst_cell_101_88 (.BL(BL88),.BLN(BLN88),.WL(WL101));
sram_cell_6t_5 inst_cell_101_89 (.BL(BL89),.BLN(BLN89),.WL(WL101));
sram_cell_6t_5 inst_cell_101_90 (.BL(BL90),.BLN(BLN90),.WL(WL101));
sram_cell_6t_5 inst_cell_101_91 (.BL(BL91),.BLN(BLN91),.WL(WL101));
sram_cell_6t_5 inst_cell_101_92 (.BL(BL92),.BLN(BLN92),.WL(WL101));
sram_cell_6t_5 inst_cell_101_93 (.BL(BL93),.BLN(BLN93),.WL(WL101));
sram_cell_6t_5 inst_cell_101_94 (.BL(BL94),.BLN(BLN94),.WL(WL101));
sram_cell_6t_5 inst_cell_101_95 (.BL(BL95),.BLN(BLN95),.WL(WL101));
sram_cell_6t_5 inst_cell_101_96 (.BL(BL96),.BLN(BLN96),.WL(WL101));
sram_cell_6t_5 inst_cell_101_97 (.BL(BL97),.BLN(BLN97),.WL(WL101));
sram_cell_6t_5 inst_cell_101_98 (.BL(BL98),.BLN(BLN98),.WL(WL101));
sram_cell_6t_5 inst_cell_101_99 (.BL(BL99),.BLN(BLN99),.WL(WL101));
sram_cell_6t_5 inst_cell_101_100 (.BL(BL100),.BLN(BLN100),.WL(WL101));
sram_cell_6t_5 inst_cell_101_101 (.BL(BL101),.BLN(BLN101),.WL(WL101));
sram_cell_6t_5 inst_cell_101_102 (.BL(BL102),.BLN(BLN102),.WL(WL101));
sram_cell_6t_5 inst_cell_101_103 (.BL(BL103),.BLN(BLN103),.WL(WL101));
sram_cell_6t_5 inst_cell_101_104 (.BL(BL104),.BLN(BLN104),.WL(WL101));
sram_cell_6t_5 inst_cell_101_105 (.BL(BL105),.BLN(BLN105),.WL(WL101));
sram_cell_6t_5 inst_cell_101_106 (.BL(BL106),.BLN(BLN106),.WL(WL101));
sram_cell_6t_5 inst_cell_101_107 (.BL(BL107),.BLN(BLN107),.WL(WL101));
sram_cell_6t_5 inst_cell_101_108 (.BL(BL108),.BLN(BLN108),.WL(WL101));
sram_cell_6t_5 inst_cell_101_109 (.BL(BL109),.BLN(BLN109),.WL(WL101));
sram_cell_6t_5 inst_cell_101_110 (.BL(BL110),.BLN(BLN110),.WL(WL101));
sram_cell_6t_5 inst_cell_101_111 (.BL(BL111),.BLN(BLN111),.WL(WL101));
sram_cell_6t_5 inst_cell_101_112 (.BL(BL112),.BLN(BLN112),.WL(WL101));
sram_cell_6t_5 inst_cell_101_113 (.BL(BL113),.BLN(BLN113),.WL(WL101));
sram_cell_6t_5 inst_cell_101_114 (.BL(BL114),.BLN(BLN114),.WL(WL101));
sram_cell_6t_5 inst_cell_101_115 (.BL(BL115),.BLN(BLN115),.WL(WL101));
sram_cell_6t_5 inst_cell_101_116 (.BL(BL116),.BLN(BLN116),.WL(WL101));
sram_cell_6t_5 inst_cell_101_117 (.BL(BL117),.BLN(BLN117),.WL(WL101));
sram_cell_6t_5 inst_cell_101_118 (.BL(BL118),.BLN(BLN118),.WL(WL101));
sram_cell_6t_5 inst_cell_101_119 (.BL(BL119),.BLN(BLN119),.WL(WL101));
sram_cell_6t_5 inst_cell_101_120 (.BL(BL120),.BLN(BLN120),.WL(WL101));
sram_cell_6t_5 inst_cell_101_121 (.BL(BL121),.BLN(BLN121),.WL(WL101));
sram_cell_6t_5 inst_cell_101_122 (.BL(BL122),.BLN(BLN122),.WL(WL101));
sram_cell_6t_5 inst_cell_101_123 (.BL(BL123),.BLN(BLN123),.WL(WL101));
sram_cell_6t_5 inst_cell_101_124 (.BL(BL124),.BLN(BLN124),.WL(WL101));
sram_cell_6t_5 inst_cell_101_125 (.BL(BL125),.BLN(BLN125),.WL(WL101));
sram_cell_6t_5 inst_cell_101_126 (.BL(BL126),.BLN(BLN126),.WL(WL101));
sram_cell_6t_5 inst_cell_101_127 (.BL(BL127),.BLN(BLN127),.WL(WL101));
sram_cell_6t_5 inst_cell_102_0 (.BL(BL0),.BLN(BLN0),.WL(WL102));
sram_cell_6t_5 inst_cell_102_1 (.BL(BL1),.BLN(BLN1),.WL(WL102));
sram_cell_6t_5 inst_cell_102_2 (.BL(BL2),.BLN(BLN2),.WL(WL102));
sram_cell_6t_5 inst_cell_102_3 (.BL(BL3),.BLN(BLN3),.WL(WL102));
sram_cell_6t_5 inst_cell_102_4 (.BL(BL4),.BLN(BLN4),.WL(WL102));
sram_cell_6t_5 inst_cell_102_5 (.BL(BL5),.BLN(BLN5),.WL(WL102));
sram_cell_6t_5 inst_cell_102_6 (.BL(BL6),.BLN(BLN6),.WL(WL102));
sram_cell_6t_5 inst_cell_102_7 (.BL(BL7),.BLN(BLN7),.WL(WL102));
sram_cell_6t_5 inst_cell_102_8 (.BL(BL8),.BLN(BLN8),.WL(WL102));
sram_cell_6t_5 inst_cell_102_9 (.BL(BL9),.BLN(BLN9),.WL(WL102));
sram_cell_6t_5 inst_cell_102_10 (.BL(BL10),.BLN(BLN10),.WL(WL102));
sram_cell_6t_5 inst_cell_102_11 (.BL(BL11),.BLN(BLN11),.WL(WL102));
sram_cell_6t_5 inst_cell_102_12 (.BL(BL12),.BLN(BLN12),.WL(WL102));
sram_cell_6t_5 inst_cell_102_13 (.BL(BL13),.BLN(BLN13),.WL(WL102));
sram_cell_6t_5 inst_cell_102_14 (.BL(BL14),.BLN(BLN14),.WL(WL102));
sram_cell_6t_5 inst_cell_102_15 (.BL(BL15),.BLN(BLN15),.WL(WL102));
sram_cell_6t_5 inst_cell_102_16 (.BL(BL16),.BLN(BLN16),.WL(WL102));
sram_cell_6t_5 inst_cell_102_17 (.BL(BL17),.BLN(BLN17),.WL(WL102));
sram_cell_6t_5 inst_cell_102_18 (.BL(BL18),.BLN(BLN18),.WL(WL102));
sram_cell_6t_5 inst_cell_102_19 (.BL(BL19),.BLN(BLN19),.WL(WL102));
sram_cell_6t_5 inst_cell_102_20 (.BL(BL20),.BLN(BLN20),.WL(WL102));
sram_cell_6t_5 inst_cell_102_21 (.BL(BL21),.BLN(BLN21),.WL(WL102));
sram_cell_6t_5 inst_cell_102_22 (.BL(BL22),.BLN(BLN22),.WL(WL102));
sram_cell_6t_5 inst_cell_102_23 (.BL(BL23),.BLN(BLN23),.WL(WL102));
sram_cell_6t_5 inst_cell_102_24 (.BL(BL24),.BLN(BLN24),.WL(WL102));
sram_cell_6t_5 inst_cell_102_25 (.BL(BL25),.BLN(BLN25),.WL(WL102));
sram_cell_6t_5 inst_cell_102_26 (.BL(BL26),.BLN(BLN26),.WL(WL102));
sram_cell_6t_5 inst_cell_102_27 (.BL(BL27),.BLN(BLN27),.WL(WL102));
sram_cell_6t_5 inst_cell_102_28 (.BL(BL28),.BLN(BLN28),.WL(WL102));
sram_cell_6t_5 inst_cell_102_29 (.BL(BL29),.BLN(BLN29),.WL(WL102));
sram_cell_6t_5 inst_cell_102_30 (.BL(BL30),.BLN(BLN30),.WL(WL102));
sram_cell_6t_5 inst_cell_102_31 (.BL(BL31),.BLN(BLN31),.WL(WL102));
sram_cell_6t_5 inst_cell_102_32 (.BL(BL32),.BLN(BLN32),.WL(WL102));
sram_cell_6t_5 inst_cell_102_33 (.BL(BL33),.BLN(BLN33),.WL(WL102));
sram_cell_6t_5 inst_cell_102_34 (.BL(BL34),.BLN(BLN34),.WL(WL102));
sram_cell_6t_5 inst_cell_102_35 (.BL(BL35),.BLN(BLN35),.WL(WL102));
sram_cell_6t_5 inst_cell_102_36 (.BL(BL36),.BLN(BLN36),.WL(WL102));
sram_cell_6t_5 inst_cell_102_37 (.BL(BL37),.BLN(BLN37),.WL(WL102));
sram_cell_6t_5 inst_cell_102_38 (.BL(BL38),.BLN(BLN38),.WL(WL102));
sram_cell_6t_5 inst_cell_102_39 (.BL(BL39),.BLN(BLN39),.WL(WL102));
sram_cell_6t_5 inst_cell_102_40 (.BL(BL40),.BLN(BLN40),.WL(WL102));
sram_cell_6t_5 inst_cell_102_41 (.BL(BL41),.BLN(BLN41),.WL(WL102));
sram_cell_6t_5 inst_cell_102_42 (.BL(BL42),.BLN(BLN42),.WL(WL102));
sram_cell_6t_5 inst_cell_102_43 (.BL(BL43),.BLN(BLN43),.WL(WL102));
sram_cell_6t_5 inst_cell_102_44 (.BL(BL44),.BLN(BLN44),.WL(WL102));
sram_cell_6t_5 inst_cell_102_45 (.BL(BL45),.BLN(BLN45),.WL(WL102));
sram_cell_6t_5 inst_cell_102_46 (.BL(BL46),.BLN(BLN46),.WL(WL102));
sram_cell_6t_5 inst_cell_102_47 (.BL(BL47),.BLN(BLN47),.WL(WL102));
sram_cell_6t_5 inst_cell_102_48 (.BL(BL48),.BLN(BLN48),.WL(WL102));
sram_cell_6t_5 inst_cell_102_49 (.BL(BL49),.BLN(BLN49),.WL(WL102));
sram_cell_6t_5 inst_cell_102_50 (.BL(BL50),.BLN(BLN50),.WL(WL102));
sram_cell_6t_5 inst_cell_102_51 (.BL(BL51),.BLN(BLN51),.WL(WL102));
sram_cell_6t_5 inst_cell_102_52 (.BL(BL52),.BLN(BLN52),.WL(WL102));
sram_cell_6t_5 inst_cell_102_53 (.BL(BL53),.BLN(BLN53),.WL(WL102));
sram_cell_6t_5 inst_cell_102_54 (.BL(BL54),.BLN(BLN54),.WL(WL102));
sram_cell_6t_5 inst_cell_102_55 (.BL(BL55),.BLN(BLN55),.WL(WL102));
sram_cell_6t_5 inst_cell_102_56 (.BL(BL56),.BLN(BLN56),.WL(WL102));
sram_cell_6t_5 inst_cell_102_57 (.BL(BL57),.BLN(BLN57),.WL(WL102));
sram_cell_6t_5 inst_cell_102_58 (.BL(BL58),.BLN(BLN58),.WL(WL102));
sram_cell_6t_5 inst_cell_102_59 (.BL(BL59),.BLN(BLN59),.WL(WL102));
sram_cell_6t_5 inst_cell_102_60 (.BL(BL60),.BLN(BLN60),.WL(WL102));
sram_cell_6t_5 inst_cell_102_61 (.BL(BL61),.BLN(BLN61),.WL(WL102));
sram_cell_6t_5 inst_cell_102_62 (.BL(BL62),.BLN(BLN62),.WL(WL102));
sram_cell_6t_5 inst_cell_102_63 (.BL(BL63),.BLN(BLN63),.WL(WL102));
sram_cell_6t_5 inst_cell_102_64 (.BL(BL64),.BLN(BLN64),.WL(WL102));
sram_cell_6t_5 inst_cell_102_65 (.BL(BL65),.BLN(BLN65),.WL(WL102));
sram_cell_6t_5 inst_cell_102_66 (.BL(BL66),.BLN(BLN66),.WL(WL102));
sram_cell_6t_5 inst_cell_102_67 (.BL(BL67),.BLN(BLN67),.WL(WL102));
sram_cell_6t_5 inst_cell_102_68 (.BL(BL68),.BLN(BLN68),.WL(WL102));
sram_cell_6t_5 inst_cell_102_69 (.BL(BL69),.BLN(BLN69),.WL(WL102));
sram_cell_6t_5 inst_cell_102_70 (.BL(BL70),.BLN(BLN70),.WL(WL102));
sram_cell_6t_5 inst_cell_102_71 (.BL(BL71),.BLN(BLN71),.WL(WL102));
sram_cell_6t_5 inst_cell_102_72 (.BL(BL72),.BLN(BLN72),.WL(WL102));
sram_cell_6t_5 inst_cell_102_73 (.BL(BL73),.BLN(BLN73),.WL(WL102));
sram_cell_6t_5 inst_cell_102_74 (.BL(BL74),.BLN(BLN74),.WL(WL102));
sram_cell_6t_5 inst_cell_102_75 (.BL(BL75),.BLN(BLN75),.WL(WL102));
sram_cell_6t_5 inst_cell_102_76 (.BL(BL76),.BLN(BLN76),.WL(WL102));
sram_cell_6t_5 inst_cell_102_77 (.BL(BL77),.BLN(BLN77),.WL(WL102));
sram_cell_6t_5 inst_cell_102_78 (.BL(BL78),.BLN(BLN78),.WL(WL102));
sram_cell_6t_5 inst_cell_102_79 (.BL(BL79),.BLN(BLN79),.WL(WL102));
sram_cell_6t_5 inst_cell_102_80 (.BL(BL80),.BLN(BLN80),.WL(WL102));
sram_cell_6t_5 inst_cell_102_81 (.BL(BL81),.BLN(BLN81),.WL(WL102));
sram_cell_6t_5 inst_cell_102_82 (.BL(BL82),.BLN(BLN82),.WL(WL102));
sram_cell_6t_5 inst_cell_102_83 (.BL(BL83),.BLN(BLN83),.WL(WL102));
sram_cell_6t_5 inst_cell_102_84 (.BL(BL84),.BLN(BLN84),.WL(WL102));
sram_cell_6t_5 inst_cell_102_85 (.BL(BL85),.BLN(BLN85),.WL(WL102));
sram_cell_6t_5 inst_cell_102_86 (.BL(BL86),.BLN(BLN86),.WL(WL102));
sram_cell_6t_5 inst_cell_102_87 (.BL(BL87),.BLN(BLN87),.WL(WL102));
sram_cell_6t_5 inst_cell_102_88 (.BL(BL88),.BLN(BLN88),.WL(WL102));
sram_cell_6t_5 inst_cell_102_89 (.BL(BL89),.BLN(BLN89),.WL(WL102));
sram_cell_6t_5 inst_cell_102_90 (.BL(BL90),.BLN(BLN90),.WL(WL102));
sram_cell_6t_5 inst_cell_102_91 (.BL(BL91),.BLN(BLN91),.WL(WL102));
sram_cell_6t_5 inst_cell_102_92 (.BL(BL92),.BLN(BLN92),.WL(WL102));
sram_cell_6t_5 inst_cell_102_93 (.BL(BL93),.BLN(BLN93),.WL(WL102));
sram_cell_6t_5 inst_cell_102_94 (.BL(BL94),.BLN(BLN94),.WL(WL102));
sram_cell_6t_5 inst_cell_102_95 (.BL(BL95),.BLN(BLN95),.WL(WL102));
sram_cell_6t_5 inst_cell_102_96 (.BL(BL96),.BLN(BLN96),.WL(WL102));
sram_cell_6t_5 inst_cell_102_97 (.BL(BL97),.BLN(BLN97),.WL(WL102));
sram_cell_6t_5 inst_cell_102_98 (.BL(BL98),.BLN(BLN98),.WL(WL102));
sram_cell_6t_5 inst_cell_102_99 (.BL(BL99),.BLN(BLN99),.WL(WL102));
sram_cell_6t_5 inst_cell_102_100 (.BL(BL100),.BLN(BLN100),.WL(WL102));
sram_cell_6t_5 inst_cell_102_101 (.BL(BL101),.BLN(BLN101),.WL(WL102));
sram_cell_6t_5 inst_cell_102_102 (.BL(BL102),.BLN(BLN102),.WL(WL102));
sram_cell_6t_5 inst_cell_102_103 (.BL(BL103),.BLN(BLN103),.WL(WL102));
sram_cell_6t_5 inst_cell_102_104 (.BL(BL104),.BLN(BLN104),.WL(WL102));
sram_cell_6t_5 inst_cell_102_105 (.BL(BL105),.BLN(BLN105),.WL(WL102));
sram_cell_6t_5 inst_cell_102_106 (.BL(BL106),.BLN(BLN106),.WL(WL102));
sram_cell_6t_5 inst_cell_102_107 (.BL(BL107),.BLN(BLN107),.WL(WL102));
sram_cell_6t_5 inst_cell_102_108 (.BL(BL108),.BLN(BLN108),.WL(WL102));
sram_cell_6t_5 inst_cell_102_109 (.BL(BL109),.BLN(BLN109),.WL(WL102));
sram_cell_6t_5 inst_cell_102_110 (.BL(BL110),.BLN(BLN110),.WL(WL102));
sram_cell_6t_5 inst_cell_102_111 (.BL(BL111),.BLN(BLN111),.WL(WL102));
sram_cell_6t_5 inst_cell_102_112 (.BL(BL112),.BLN(BLN112),.WL(WL102));
sram_cell_6t_5 inst_cell_102_113 (.BL(BL113),.BLN(BLN113),.WL(WL102));
sram_cell_6t_5 inst_cell_102_114 (.BL(BL114),.BLN(BLN114),.WL(WL102));
sram_cell_6t_5 inst_cell_102_115 (.BL(BL115),.BLN(BLN115),.WL(WL102));
sram_cell_6t_5 inst_cell_102_116 (.BL(BL116),.BLN(BLN116),.WL(WL102));
sram_cell_6t_5 inst_cell_102_117 (.BL(BL117),.BLN(BLN117),.WL(WL102));
sram_cell_6t_5 inst_cell_102_118 (.BL(BL118),.BLN(BLN118),.WL(WL102));
sram_cell_6t_5 inst_cell_102_119 (.BL(BL119),.BLN(BLN119),.WL(WL102));
sram_cell_6t_5 inst_cell_102_120 (.BL(BL120),.BLN(BLN120),.WL(WL102));
sram_cell_6t_5 inst_cell_102_121 (.BL(BL121),.BLN(BLN121),.WL(WL102));
sram_cell_6t_5 inst_cell_102_122 (.BL(BL122),.BLN(BLN122),.WL(WL102));
sram_cell_6t_5 inst_cell_102_123 (.BL(BL123),.BLN(BLN123),.WL(WL102));
sram_cell_6t_5 inst_cell_102_124 (.BL(BL124),.BLN(BLN124),.WL(WL102));
sram_cell_6t_5 inst_cell_102_125 (.BL(BL125),.BLN(BLN125),.WL(WL102));
sram_cell_6t_5 inst_cell_102_126 (.BL(BL126),.BLN(BLN126),.WL(WL102));
sram_cell_6t_5 inst_cell_102_127 (.BL(BL127),.BLN(BLN127),.WL(WL102));
sram_cell_6t_5 inst_cell_103_0 (.BL(BL0),.BLN(BLN0),.WL(WL103));
sram_cell_6t_5 inst_cell_103_1 (.BL(BL1),.BLN(BLN1),.WL(WL103));
sram_cell_6t_5 inst_cell_103_2 (.BL(BL2),.BLN(BLN2),.WL(WL103));
sram_cell_6t_5 inst_cell_103_3 (.BL(BL3),.BLN(BLN3),.WL(WL103));
sram_cell_6t_5 inst_cell_103_4 (.BL(BL4),.BLN(BLN4),.WL(WL103));
sram_cell_6t_5 inst_cell_103_5 (.BL(BL5),.BLN(BLN5),.WL(WL103));
sram_cell_6t_5 inst_cell_103_6 (.BL(BL6),.BLN(BLN6),.WL(WL103));
sram_cell_6t_5 inst_cell_103_7 (.BL(BL7),.BLN(BLN7),.WL(WL103));
sram_cell_6t_5 inst_cell_103_8 (.BL(BL8),.BLN(BLN8),.WL(WL103));
sram_cell_6t_5 inst_cell_103_9 (.BL(BL9),.BLN(BLN9),.WL(WL103));
sram_cell_6t_5 inst_cell_103_10 (.BL(BL10),.BLN(BLN10),.WL(WL103));
sram_cell_6t_5 inst_cell_103_11 (.BL(BL11),.BLN(BLN11),.WL(WL103));
sram_cell_6t_5 inst_cell_103_12 (.BL(BL12),.BLN(BLN12),.WL(WL103));
sram_cell_6t_5 inst_cell_103_13 (.BL(BL13),.BLN(BLN13),.WL(WL103));
sram_cell_6t_5 inst_cell_103_14 (.BL(BL14),.BLN(BLN14),.WL(WL103));
sram_cell_6t_5 inst_cell_103_15 (.BL(BL15),.BLN(BLN15),.WL(WL103));
sram_cell_6t_5 inst_cell_103_16 (.BL(BL16),.BLN(BLN16),.WL(WL103));
sram_cell_6t_5 inst_cell_103_17 (.BL(BL17),.BLN(BLN17),.WL(WL103));
sram_cell_6t_5 inst_cell_103_18 (.BL(BL18),.BLN(BLN18),.WL(WL103));
sram_cell_6t_5 inst_cell_103_19 (.BL(BL19),.BLN(BLN19),.WL(WL103));
sram_cell_6t_5 inst_cell_103_20 (.BL(BL20),.BLN(BLN20),.WL(WL103));
sram_cell_6t_5 inst_cell_103_21 (.BL(BL21),.BLN(BLN21),.WL(WL103));
sram_cell_6t_5 inst_cell_103_22 (.BL(BL22),.BLN(BLN22),.WL(WL103));
sram_cell_6t_5 inst_cell_103_23 (.BL(BL23),.BLN(BLN23),.WL(WL103));
sram_cell_6t_5 inst_cell_103_24 (.BL(BL24),.BLN(BLN24),.WL(WL103));
sram_cell_6t_5 inst_cell_103_25 (.BL(BL25),.BLN(BLN25),.WL(WL103));
sram_cell_6t_5 inst_cell_103_26 (.BL(BL26),.BLN(BLN26),.WL(WL103));
sram_cell_6t_5 inst_cell_103_27 (.BL(BL27),.BLN(BLN27),.WL(WL103));
sram_cell_6t_5 inst_cell_103_28 (.BL(BL28),.BLN(BLN28),.WL(WL103));
sram_cell_6t_5 inst_cell_103_29 (.BL(BL29),.BLN(BLN29),.WL(WL103));
sram_cell_6t_5 inst_cell_103_30 (.BL(BL30),.BLN(BLN30),.WL(WL103));
sram_cell_6t_5 inst_cell_103_31 (.BL(BL31),.BLN(BLN31),.WL(WL103));
sram_cell_6t_5 inst_cell_103_32 (.BL(BL32),.BLN(BLN32),.WL(WL103));
sram_cell_6t_5 inst_cell_103_33 (.BL(BL33),.BLN(BLN33),.WL(WL103));
sram_cell_6t_5 inst_cell_103_34 (.BL(BL34),.BLN(BLN34),.WL(WL103));
sram_cell_6t_5 inst_cell_103_35 (.BL(BL35),.BLN(BLN35),.WL(WL103));
sram_cell_6t_5 inst_cell_103_36 (.BL(BL36),.BLN(BLN36),.WL(WL103));
sram_cell_6t_5 inst_cell_103_37 (.BL(BL37),.BLN(BLN37),.WL(WL103));
sram_cell_6t_5 inst_cell_103_38 (.BL(BL38),.BLN(BLN38),.WL(WL103));
sram_cell_6t_5 inst_cell_103_39 (.BL(BL39),.BLN(BLN39),.WL(WL103));
sram_cell_6t_5 inst_cell_103_40 (.BL(BL40),.BLN(BLN40),.WL(WL103));
sram_cell_6t_5 inst_cell_103_41 (.BL(BL41),.BLN(BLN41),.WL(WL103));
sram_cell_6t_5 inst_cell_103_42 (.BL(BL42),.BLN(BLN42),.WL(WL103));
sram_cell_6t_5 inst_cell_103_43 (.BL(BL43),.BLN(BLN43),.WL(WL103));
sram_cell_6t_5 inst_cell_103_44 (.BL(BL44),.BLN(BLN44),.WL(WL103));
sram_cell_6t_5 inst_cell_103_45 (.BL(BL45),.BLN(BLN45),.WL(WL103));
sram_cell_6t_5 inst_cell_103_46 (.BL(BL46),.BLN(BLN46),.WL(WL103));
sram_cell_6t_5 inst_cell_103_47 (.BL(BL47),.BLN(BLN47),.WL(WL103));
sram_cell_6t_5 inst_cell_103_48 (.BL(BL48),.BLN(BLN48),.WL(WL103));
sram_cell_6t_5 inst_cell_103_49 (.BL(BL49),.BLN(BLN49),.WL(WL103));
sram_cell_6t_5 inst_cell_103_50 (.BL(BL50),.BLN(BLN50),.WL(WL103));
sram_cell_6t_5 inst_cell_103_51 (.BL(BL51),.BLN(BLN51),.WL(WL103));
sram_cell_6t_5 inst_cell_103_52 (.BL(BL52),.BLN(BLN52),.WL(WL103));
sram_cell_6t_5 inst_cell_103_53 (.BL(BL53),.BLN(BLN53),.WL(WL103));
sram_cell_6t_5 inst_cell_103_54 (.BL(BL54),.BLN(BLN54),.WL(WL103));
sram_cell_6t_5 inst_cell_103_55 (.BL(BL55),.BLN(BLN55),.WL(WL103));
sram_cell_6t_5 inst_cell_103_56 (.BL(BL56),.BLN(BLN56),.WL(WL103));
sram_cell_6t_5 inst_cell_103_57 (.BL(BL57),.BLN(BLN57),.WL(WL103));
sram_cell_6t_5 inst_cell_103_58 (.BL(BL58),.BLN(BLN58),.WL(WL103));
sram_cell_6t_5 inst_cell_103_59 (.BL(BL59),.BLN(BLN59),.WL(WL103));
sram_cell_6t_5 inst_cell_103_60 (.BL(BL60),.BLN(BLN60),.WL(WL103));
sram_cell_6t_5 inst_cell_103_61 (.BL(BL61),.BLN(BLN61),.WL(WL103));
sram_cell_6t_5 inst_cell_103_62 (.BL(BL62),.BLN(BLN62),.WL(WL103));
sram_cell_6t_5 inst_cell_103_63 (.BL(BL63),.BLN(BLN63),.WL(WL103));
sram_cell_6t_5 inst_cell_103_64 (.BL(BL64),.BLN(BLN64),.WL(WL103));
sram_cell_6t_5 inst_cell_103_65 (.BL(BL65),.BLN(BLN65),.WL(WL103));
sram_cell_6t_5 inst_cell_103_66 (.BL(BL66),.BLN(BLN66),.WL(WL103));
sram_cell_6t_5 inst_cell_103_67 (.BL(BL67),.BLN(BLN67),.WL(WL103));
sram_cell_6t_5 inst_cell_103_68 (.BL(BL68),.BLN(BLN68),.WL(WL103));
sram_cell_6t_5 inst_cell_103_69 (.BL(BL69),.BLN(BLN69),.WL(WL103));
sram_cell_6t_5 inst_cell_103_70 (.BL(BL70),.BLN(BLN70),.WL(WL103));
sram_cell_6t_5 inst_cell_103_71 (.BL(BL71),.BLN(BLN71),.WL(WL103));
sram_cell_6t_5 inst_cell_103_72 (.BL(BL72),.BLN(BLN72),.WL(WL103));
sram_cell_6t_5 inst_cell_103_73 (.BL(BL73),.BLN(BLN73),.WL(WL103));
sram_cell_6t_5 inst_cell_103_74 (.BL(BL74),.BLN(BLN74),.WL(WL103));
sram_cell_6t_5 inst_cell_103_75 (.BL(BL75),.BLN(BLN75),.WL(WL103));
sram_cell_6t_5 inst_cell_103_76 (.BL(BL76),.BLN(BLN76),.WL(WL103));
sram_cell_6t_5 inst_cell_103_77 (.BL(BL77),.BLN(BLN77),.WL(WL103));
sram_cell_6t_5 inst_cell_103_78 (.BL(BL78),.BLN(BLN78),.WL(WL103));
sram_cell_6t_5 inst_cell_103_79 (.BL(BL79),.BLN(BLN79),.WL(WL103));
sram_cell_6t_5 inst_cell_103_80 (.BL(BL80),.BLN(BLN80),.WL(WL103));
sram_cell_6t_5 inst_cell_103_81 (.BL(BL81),.BLN(BLN81),.WL(WL103));
sram_cell_6t_5 inst_cell_103_82 (.BL(BL82),.BLN(BLN82),.WL(WL103));
sram_cell_6t_5 inst_cell_103_83 (.BL(BL83),.BLN(BLN83),.WL(WL103));
sram_cell_6t_5 inst_cell_103_84 (.BL(BL84),.BLN(BLN84),.WL(WL103));
sram_cell_6t_5 inst_cell_103_85 (.BL(BL85),.BLN(BLN85),.WL(WL103));
sram_cell_6t_5 inst_cell_103_86 (.BL(BL86),.BLN(BLN86),.WL(WL103));
sram_cell_6t_5 inst_cell_103_87 (.BL(BL87),.BLN(BLN87),.WL(WL103));
sram_cell_6t_5 inst_cell_103_88 (.BL(BL88),.BLN(BLN88),.WL(WL103));
sram_cell_6t_5 inst_cell_103_89 (.BL(BL89),.BLN(BLN89),.WL(WL103));
sram_cell_6t_5 inst_cell_103_90 (.BL(BL90),.BLN(BLN90),.WL(WL103));
sram_cell_6t_5 inst_cell_103_91 (.BL(BL91),.BLN(BLN91),.WL(WL103));
sram_cell_6t_5 inst_cell_103_92 (.BL(BL92),.BLN(BLN92),.WL(WL103));
sram_cell_6t_5 inst_cell_103_93 (.BL(BL93),.BLN(BLN93),.WL(WL103));
sram_cell_6t_5 inst_cell_103_94 (.BL(BL94),.BLN(BLN94),.WL(WL103));
sram_cell_6t_5 inst_cell_103_95 (.BL(BL95),.BLN(BLN95),.WL(WL103));
sram_cell_6t_5 inst_cell_103_96 (.BL(BL96),.BLN(BLN96),.WL(WL103));
sram_cell_6t_5 inst_cell_103_97 (.BL(BL97),.BLN(BLN97),.WL(WL103));
sram_cell_6t_5 inst_cell_103_98 (.BL(BL98),.BLN(BLN98),.WL(WL103));
sram_cell_6t_5 inst_cell_103_99 (.BL(BL99),.BLN(BLN99),.WL(WL103));
sram_cell_6t_5 inst_cell_103_100 (.BL(BL100),.BLN(BLN100),.WL(WL103));
sram_cell_6t_5 inst_cell_103_101 (.BL(BL101),.BLN(BLN101),.WL(WL103));
sram_cell_6t_5 inst_cell_103_102 (.BL(BL102),.BLN(BLN102),.WL(WL103));
sram_cell_6t_5 inst_cell_103_103 (.BL(BL103),.BLN(BLN103),.WL(WL103));
sram_cell_6t_5 inst_cell_103_104 (.BL(BL104),.BLN(BLN104),.WL(WL103));
sram_cell_6t_5 inst_cell_103_105 (.BL(BL105),.BLN(BLN105),.WL(WL103));
sram_cell_6t_5 inst_cell_103_106 (.BL(BL106),.BLN(BLN106),.WL(WL103));
sram_cell_6t_5 inst_cell_103_107 (.BL(BL107),.BLN(BLN107),.WL(WL103));
sram_cell_6t_5 inst_cell_103_108 (.BL(BL108),.BLN(BLN108),.WL(WL103));
sram_cell_6t_5 inst_cell_103_109 (.BL(BL109),.BLN(BLN109),.WL(WL103));
sram_cell_6t_5 inst_cell_103_110 (.BL(BL110),.BLN(BLN110),.WL(WL103));
sram_cell_6t_5 inst_cell_103_111 (.BL(BL111),.BLN(BLN111),.WL(WL103));
sram_cell_6t_5 inst_cell_103_112 (.BL(BL112),.BLN(BLN112),.WL(WL103));
sram_cell_6t_5 inst_cell_103_113 (.BL(BL113),.BLN(BLN113),.WL(WL103));
sram_cell_6t_5 inst_cell_103_114 (.BL(BL114),.BLN(BLN114),.WL(WL103));
sram_cell_6t_5 inst_cell_103_115 (.BL(BL115),.BLN(BLN115),.WL(WL103));
sram_cell_6t_5 inst_cell_103_116 (.BL(BL116),.BLN(BLN116),.WL(WL103));
sram_cell_6t_5 inst_cell_103_117 (.BL(BL117),.BLN(BLN117),.WL(WL103));
sram_cell_6t_5 inst_cell_103_118 (.BL(BL118),.BLN(BLN118),.WL(WL103));
sram_cell_6t_5 inst_cell_103_119 (.BL(BL119),.BLN(BLN119),.WL(WL103));
sram_cell_6t_5 inst_cell_103_120 (.BL(BL120),.BLN(BLN120),.WL(WL103));
sram_cell_6t_5 inst_cell_103_121 (.BL(BL121),.BLN(BLN121),.WL(WL103));
sram_cell_6t_5 inst_cell_103_122 (.BL(BL122),.BLN(BLN122),.WL(WL103));
sram_cell_6t_5 inst_cell_103_123 (.BL(BL123),.BLN(BLN123),.WL(WL103));
sram_cell_6t_5 inst_cell_103_124 (.BL(BL124),.BLN(BLN124),.WL(WL103));
sram_cell_6t_5 inst_cell_103_125 (.BL(BL125),.BLN(BLN125),.WL(WL103));
sram_cell_6t_5 inst_cell_103_126 (.BL(BL126),.BLN(BLN126),.WL(WL103));
sram_cell_6t_5 inst_cell_103_127 (.BL(BL127),.BLN(BLN127),.WL(WL103));
sram_cell_6t_5 inst_cell_104_0 (.BL(BL0),.BLN(BLN0),.WL(WL104));
sram_cell_6t_5 inst_cell_104_1 (.BL(BL1),.BLN(BLN1),.WL(WL104));
sram_cell_6t_5 inst_cell_104_2 (.BL(BL2),.BLN(BLN2),.WL(WL104));
sram_cell_6t_5 inst_cell_104_3 (.BL(BL3),.BLN(BLN3),.WL(WL104));
sram_cell_6t_5 inst_cell_104_4 (.BL(BL4),.BLN(BLN4),.WL(WL104));
sram_cell_6t_5 inst_cell_104_5 (.BL(BL5),.BLN(BLN5),.WL(WL104));
sram_cell_6t_5 inst_cell_104_6 (.BL(BL6),.BLN(BLN6),.WL(WL104));
sram_cell_6t_5 inst_cell_104_7 (.BL(BL7),.BLN(BLN7),.WL(WL104));
sram_cell_6t_5 inst_cell_104_8 (.BL(BL8),.BLN(BLN8),.WL(WL104));
sram_cell_6t_5 inst_cell_104_9 (.BL(BL9),.BLN(BLN9),.WL(WL104));
sram_cell_6t_5 inst_cell_104_10 (.BL(BL10),.BLN(BLN10),.WL(WL104));
sram_cell_6t_5 inst_cell_104_11 (.BL(BL11),.BLN(BLN11),.WL(WL104));
sram_cell_6t_5 inst_cell_104_12 (.BL(BL12),.BLN(BLN12),.WL(WL104));
sram_cell_6t_5 inst_cell_104_13 (.BL(BL13),.BLN(BLN13),.WL(WL104));
sram_cell_6t_5 inst_cell_104_14 (.BL(BL14),.BLN(BLN14),.WL(WL104));
sram_cell_6t_5 inst_cell_104_15 (.BL(BL15),.BLN(BLN15),.WL(WL104));
sram_cell_6t_5 inst_cell_104_16 (.BL(BL16),.BLN(BLN16),.WL(WL104));
sram_cell_6t_5 inst_cell_104_17 (.BL(BL17),.BLN(BLN17),.WL(WL104));
sram_cell_6t_5 inst_cell_104_18 (.BL(BL18),.BLN(BLN18),.WL(WL104));
sram_cell_6t_5 inst_cell_104_19 (.BL(BL19),.BLN(BLN19),.WL(WL104));
sram_cell_6t_5 inst_cell_104_20 (.BL(BL20),.BLN(BLN20),.WL(WL104));
sram_cell_6t_5 inst_cell_104_21 (.BL(BL21),.BLN(BLN21),.WL(WL104));
sram_cell_6t_5 inst_cell_104_22 (.BL(BL22),.BLN(BLN22),.WL(WL104));
sram_cell_6t_5 inst_cell_104_23 (.BL(BL23),.BLN(BLN23),.WL(WL104));
sram_cell_6t_5 inst_cell_104_24 (.BL(BL24),.BLN(BLN24),.WL(WL104));
sram_cell_6t_5 inst_cell_104_25 (.BL(BL25),.BLN(BLN25),.WL(WL104));
sram_cell_6t_5 inst_cell_104_26 (.BL(BL26),.BLN(BLN26),.WL(WL104));
sram_cell_6t_5 inst_cell_104_27 (.BL(BL27),.BLN(BLN27),.WL(WL104));
sram_cell_6t_5 inst_cell_104_28 (.BL(BL28),.BLN(BLN28),.WL(WL104));
sram_cell_6t_5 inst_cell_104_29 (.BL(BL29),.BLN(BLN29),.WL(WL104));
sram_cell_6t_5 inst_cell_104_30 (.BL(BL30),.BLN(BLN30),.WL(WL104));
sram_cell_6t_5 inst_cell_104_31 (.BL(BL31),.BLN(BLN31),.WL(WL104));
sram_cell_6t_5 inst_cell_104_32 (.BL(BL32),.BLN(BLN32),.WL(WL104));
sram_cell_6t_5 inst_cell_104_33 (.BL(BL33),.BLN(BLN33),.WL(WL104));
sram_cell_6t_5 inst_cell_104_34 (.BL(BL34),.BLN(BLN34),.WL(WL104));
sram_cell_6t_5 inst_cell_104_35 (.BL(BL35),.BLN(BLN35),.WL(WL104));
sram_cell_6t_5 inst_cell_104_36 (.BL(BL36),.BLN(BLN36),.WL(WL104));
sram_cell_6t_5 inst_cell_104_37 (.BL(BL37),.BLN(BLN37),.WL(WL104));
sram_cell_6t_5 inst_cell_104_38 (.BL(BL38),.BLN(BLN38),.WL(WL104));
sram_cell_6t_5 inst_cell_104_39 (.BL(BL39),.BLN(BLN39),.WL(WL104));
sram_cell_6t_5 inst_cell_104_40 (.BL(BL40),.BLN(BLN40),.WL(WL104));
sram_cell_6t_5 inst_cell_104_41 (.BL(BL41),.BLN(BLN41),.WL(WL104));
sram_cell_6t_5 inst_cell_104_42 (.BL(BL42),.BLN(BLN42),.WL(WL104));
sram_cell_6t_5 inst_cell_104_43 (.BL(BL43),.BLN(BLN43),.WL(WL104));
sram_cell_6t_5 inst_cell_104_44 (.BL(BL44),.BLN(BLN44),.WL(WL104));
sram_cell_6t_5 inst_cell_104_45 (.BL(BL45),.BLN(BLN45),.WL(WL104));
sram_cell_6t_5 inst_cell_104_46 (.BL(BL46),.BLN(BLN46),.WL(WL104));
sram_cell_6t_5 inst_cell_104_47 (.BL(BL47),.BLN(BLN47),.WL(WL104));
sram_cell_6t_5 inst_cell_104_48 (.BL(BL48),.BLN(BLN48),.WL(WL104));
sram_cell_6t_5 inst_cell_104_49 (.BL(BL49),.BLN(BLN49),.WL(WL104));
sram_cell_6t_5 inst_cell_104_50 (.BL(BL50),.BLN(BLN50),.WL(WL104));
sram_cell_6t_5 inst_cell_104_51 (.BL(BL51),.BLN(BLN51),.WL(WL104));
sram_cell_6t_5 inst_cell_104_52 (.BL(BL52),.BLN(BLN52),.WL(WL104));
sram_cell_6t_5 inst_cell_104_53 (.BL(BL53),.BLN(BLN53),.WL(WL104));
sram_cell_6t_5 inst_cell_104_54 (.BL(BL54),.BLN(BLN54),.WL(WL104));
sram_cell_6t_5 inst_cell_104_55 (.BL(BL55),.BLN(BLN55),.WL(WL104));
sram_cell_6t_5 inst_cell_104_56 (.BL(BL56),.BLN(BLN56),.WL(WL104));
sram_cell_6t_5 inst_cell_104_57 (.BL(BL57),.BLN(BLN57),.WL(WL104));
sram_cell_6t_5 inst_cell_104_58 (.BL(BL58),.BLN(BLN58),.WL(WL104));
sram_cell_6t_5 inst_cell_104_59 (.BL(BL59),.BLN(BLN59),.WL(WL104));
sram_cell_6t_5 inst_cell_104_60 (.BL(BL60),.BLN(BLN60),.WL(WL104));
sram_cell_6t_5 inst_cell_104_61 (.BL(BL61),.BLN(BLN61),.WL(WL104));
sram_cell_6t_5 inst_cell_104_62 (.BL(BL62),.BLN(BLN62),.WL(WL104));
sram_cell_6t_5 inst_cell_104_63 (.BL(BL63),.BLN(BLN63),.WL(WL104));
sram_cell_6t_5 inst_cell_104_64 (.BL(BL64),.BLN(BLN64),.WL(WL104));
sram_cell_6t_5 inst_cell_104_65 (.BL(BL65),.BLN(BLN65),.WL(WL104));
sram_cell_6t_5 inst_cell_104_66 (.BL(BL66),.BLN(BLN66),.WL(WL104));
sram_cell_6t_5 inst_cell_104_67 (.BL(BL67),.BLN(BLN67),.WL(WL104));
sram_cell_6t_5 inst_cell_104_68 (.BL(BL68),.BLN(BLN68),.WL(WL104));
sram_cell_6t_5 inst_cell_104_69 (.BL(BL69),.BLN(BLN69),.WL(WL104));
sram_cell_6t_5 inst_cell_104_70 (.BL(BL70),.BLN(BLN70),.WL(WL104));
sram_cell_6t_5 inst_cell_104_71 (.BL(BL71),.BLN(BLN71),.WL(WL104));
sram_cell_6t_5 inst_cell_104_72 (.BL(BL72),.BLN(BLN72),.WL(WL104));
sram_cell_6t_5 inst_cell_104_73 (.BL(BL73),.BLN(BLN73),.WL(WL104));
sram_cell_6t_5 inst_cell_104_74 (.BL(BL74),.BLN(BLN74),.WL(WL104));
sram_cell_6t_5 inst_cell_104_75 (.BL(BL75),.BLN(BLN75),.WL(WL104));
sram_cell_6t_5 inst_cell_104_76 (.BL(BL76),.BLN(BLN76),.WL(WL104));
sram_cell_6t_5 inst_cell_104_77 (.BL(BL77),.BLN(BLN77),.WL(WL104));
sram_cell_6t_5 inst_cell_104_78 (.BL(BL78),.BLN(BLN78),.WL(WL104));
sram_cell_6t_5 inst_cell_104_79 (.BL(BL79),.BLN(BLN79),.WL(WL104));
sram_cell_6t_5 inst_cell_104_80 (.BL(BL80),.BLN(BLN80),.WL(WL104));
sram_cell_6t_5 inst_cell_104_81 (.BL(BL81),.BLN(BLN81),.WL(WL104));
sram_cell_6t_5 inst_cell_104_82 (.BL(BL82),.BLN(BLN82),.WL(WL104));
sram_cell_6t_5 inst_cell_104_83 (.BL(BL83),.BLN(BLN83),.WL(WL104));
sram_cell_6t_5 inst_cell_104_84 (.BL(BL84),.BLN(BLN84),.WL(WL104));
sram_cell_6t_5 inst_cell_104_85 (.BL(BL85),.BLN(BLN85),.WL(WL104));
sram_cell_6t_5 inst_cell_104_86 (.BL(BL86),.BLN(BLN86),.WL(WL104));
sram_cell_6t_5 inst_cell_104_87 (.BL(BL87),.BLN(BLN87),.WL(WL104));
sram_cell_6t_5 inst_cell_104_88 (.BL(BL88),.BLN(BLN88),.WL(WL104));
sram_cell_6t_5 inst_cell_104_89 (.BL(BL89),.BLN(BLN89),.WL(WL104));
sram_cell_6t_5 inst_cell_104_90 (.BL(BL90),.BLN(BLN90),.WL(WL104));
sram_cell_6t_5 inst_cell_104_91 (.BL(BL91),.BLN(BLN91),.WL(WL104));
sram_cell_6t_5 inst_cell_104_92 (.BL(BL92),.BLN(BLN92),.WL(WL104));
sram_cell_6t_5 inst_cell_104_93 (.BL(BL93),.BLN(BLN93),.WL(WL104));
sram_cell_6t_5 inst_cell_104_94 (.BL(BL94),.BLN(BLN94),.WL(WL104));
sram_cell_6t_5 inst_cell_104_95 (.BL(BL95),.BLN(BLN95),.WL(WL104));
sram_cell_6t_5 inst_cell_104_96 (.BL(BL96),.BLN(BLN96),.WL(WL104));
sram_cell_6t_5 inst_cell_104_97 (.BL(BL97),.BLN(BLN97),.WL(WL104));
sram_cell_6t_5 inst_cell_104_98 (.BL(BL98),.BLN(BLN98),.WL(WL104));
sram_cell_6t_5 inst_cell_104_99 (.BL(BL99),.BLN(BLN99),.WL(WL104));
sram_cell_6t_5 inst_cell_104_100 (.BL(BL100),.BLN(BLN100),.WL(WL104));
sram_cell_6t_5 inst_cell_104_101 (.BL(BL101),.BLN(BLN101),.WL(WL104));
sram_cell_6t_5 inst_cell_104_102 (.BL(BL102),.BLN(BLN102),.WL(WL104));
sram_cell_6t_5 inst_cell_104_103 (.BL(BL103),.BLN(BLN103),.WL(WL104));
sram_cell_6t_5 inst_cell_104_104 (.BL(BL104),.BLN(BLN104),.WL(WL104));
sram_cell_6t_5 inst_cell_104_105 (.BL(BL105),.BLN(BLN105),.WL(WL104));
sram_cell_6t_5 inst_cell_104_106 (.BL(BL106),.BLN(BLN106),.WL(WL104));
sram_cell_6t_5 inst_cell_104_107 (.BL(BL107),.BLN(BLN107),.WL(WL104));
sram_cell_6t_5 inst_cell_104_108 (.BL(BL108),.BLN(BLN108),.WL(WL104));
sram_cell_6t_5 inst_cell_104_109 (.BL(BL109),.BLN(BLN109),.WL(WL104));
sram_cell_6t_5 inst_cell_104_110 (.BL(BL110),.BLN(BLN110),.WL(WL104));
sram_cell_6t_5 inst_cell_104_111 (.BL(BL111),.BLN(BLN111),.WL(WL104));
sram_cell_6t_5 inst_cell_104_112 (.BL(BL112),.BLN(BLN112),.WL(WL104));
sram_cell_6t_5 inst_cell_104_113 (.BL(BL113),.BLN(BLN113),.WL(WL104));
sram_cell_6t_5 inst_cell_104_114 (.BL(BL114),.BLN(BLN114),.WL(WL104));
sram_cell_6t_5 inst_cell_104_115 (.BL(BL115),.BLN(BLN115),.WL(WL104));
sram_cell_6t_5 inst_cell_104_116 (.BL(BL116),.BLN(BLN116),.WL(WL104));
sram_cell_6t_5 inst_cell_104_117 (.BL(BL117),.BLN(BLN117),.WL(WL104));
sram_cell_6t_5 inst_cell_104_118 (.BL(BL118),.BLN(BLN118),.WL(WL104));
sram_cell_6t_5 inst_cell_104_119 (.BL(BL119),.BLN(BLN119),.WL(WL104));
sram_cell_6t_5 inst_cell_104_120 (.BL(BL120),.BLN(BLN120),.WL(WL104));
sram_cell_6t_5 inst_cell_104_121 (.BL(BL121),.BLN(BLN121),.WL(WL104));
sram_cell_6t_5 inst_cell_104_122 (.BL(BL122),.BLN(BLN122),.WL(WL104));
sram_cell_6t_5 inst_cell_104_123 (.BL(BL123),.BLN(BLN123),.WL(WL104));
sram_cell_6t_5 inst_cell_104_124 (.BL(BL124),.BLN(BLN124),.WL(WL104));
sram_cell_6t_5 inst_cell_104_125 (.BL(BL125),.BLN(BLN125),.WL(WL104));
sram_cell_6t_5 inst_cell_104_126 (.BL(BL126),.BLN(BLN126),.WL(WL104));
sram_cell_6t_5 inst_cell_104_127 (.BL(BL127),.BLN(BLN127),.WL(WL104));
sram_cell_6t_5 inst_cell_105_0 (.BL(BL0),.BLN(BLN0),.WL(WL105));
sram_cell_6t_5 inst_cell_105_1 (.BL(BL1),.BLN(BLN1),.WL(WL105));
sram_cell_6t_5 inst_cell_105_2 (.BL(BL2),.BLN(BLN2),.WL(WL105));
sram_cell_6t_5 inst_cell_105_3 (.BL(BL3),.BLN(BLN3),.WL(WL105));
sram_cell_6t_5 inst_cell_105_4 (.BL(BL4),.BLN(BLN4),.WL(WL105));
sram_cell_6t_5 inst_cell_105_5 (.BL(BL5),.BLN(BLN5),.WL(WL105));
sram_cell_6t_5 inst_cell_105_6 (.BL(BL6),.BLN(BLN6),.WL(WL105));
sram_cell_6t_5 inst_cell_105_7 (.BL(BL7),.BLN(BLN7),.WL(WL105));
sram_cell_6t_5 inst_cell_105_8 (.BL(BL8),.BLN(BLN8),.WL(WL105));
sram_cell_6t_5 inst_cell_105_9 (.BL(BL9),.BLN(BLN9),.WL(WL105));
sram_cell_6t_5 inst_cell_105_10 (.BL(BL10),.BLN(BLN10),.WL(WL105));
sram_cell_6t_5 inst_cell_105_11 (.BL(BL11),.BLN(BLN11),.WL(WL105));
sram_cell_6t_5 inst_cell_105_12 (.BL(BL12),.BLN(BLN12),.WL(WL105));
sram_cell_6t_5 inst_cell_105_13 (.BL(BL13),.BLN(BLN13),.WL(WL105));
sram_cell_6t_5 inst_cell_105_14 (.BL(BL14),.BLN(BLN14),.WL(WL105));
sram_cell_6t_5 inst_cell_105_15 (.BL(BL15),.BLN(BLN15),.WL(WL105));
sram_cell_6t_5 inst_cell_105_16 (.BL(BL16),.BLN(BLN16),.WL(WL105));
sram_cell_6t_5 inst_cell_105_17 (.BL(BL17),.BLN(BLN17),.WL(WL105));
sram_cell_6t_5 inst_cell_105_18 (.BL(BL18),.BLN(BLN18),.WL(WL105));
sram_cell_6t_5 inst_cell_105_19 (.BL(BL19),.BLN(BLN19),.WL(WL105));
sram_cell_6t_5 inst_cell_105_20 (.BL(BL20),.BLN(BLN20),.WL(WL105));
sram_cell_6t_5 inst_cell_105_21 (.BL(BL21),.BLN(BLN21),.WL(WL105));
sram_cell_6t_5 inst_cell_105_22 (.BL(BL22),.BLN(BLN22),.WL(WL105));
sram_cell_6t_5 inst_cell_105_23 (.BL(BL23),.BLN(BLN23),.WL(WL105));
sram_cell_6t_5 inst_cell_105_24 (.BL(BL24),.BLN(BLN24),.WL(WL105));
sram_cell_6t_5 inst_cell_105_25 (.BL(BL25),.BLN(BLN25),.WL(WL105));
sram_cell_6t_5 inst_cell_105_26 (.BL(BL26),.BLN(BLN26),.WL(WL105));
sram_cell_6t_5 inst_cell_105_27 (.BL(BL27),.BLN(BLN27),.WL(WL105));
sram_cell_6t_5 inst_cell_105_28 (.BL(BL28),.BLN(BLN28),.WL(WL105));
sram_cell_6t_5 inst_cell_105_29 (.BL(BL29),.BLN(BLN29),.WL(WL105));
sram_cell_6t_5 inst_cell_105_30 (.BL(BL30),.BLN(BLN30),.WL(WL105));
sram_cell_6t_5 inst_cell_105_31 (.BL(BL31),.BLN(BLN31),.WL(WL105));
sram_cell_6t_5 inst_cell_105_32 (.BL(BL32),.BLN(BLN32),.WL(WL105));
sram_cell_6t_5 inst_cell_105_33 (.BL(BL33),.BLN(BLN33),.WL(WL105));
sram_cell_6t_5 inst_cell_105_34 (.BL(BL34),.BLN(BLN34),.WL(WL105));
sram_cell_6t_5 inst_cell_105_35 (.BL(BL35),.BLN(BLN35),.WL(WL105));
sram_cell_6t_5 inst_cell_105_36 (.BL(BL36),.BLN(BLN36),.WL(WL105));
sram_cell_6t_5 inst_cell_105_37 (.BL(BL37),.BLN(BLN37),.WL(WL105));
sram_cell_6t_5 inst_cell_105_38 (.BL(BL38),.BLN(BLN38),.WL(WL105));
sram_cell_6t_5 inst_cell_105_39 (.BL(BL39),.BLN(BLN39),.WL(WL105));
sram_cell_6t_5 inst_cell_105_40 (.BL(BL40),.BLN(BLN40),.WL(WL105));
sram_cell_6t_5 inst_cell_105_41 (.BL(BL41),.BLN(BLN41),.WL(WL105));
sram_cell_6t_5 inst_cell_105_42 (.BL(BL42),.BLN(BLN42),.WL(WL105));
sram_cell_6t_5 inst_cell_105_43 (.BL(BL43),.BLN(BLN43),.WL(WL105));
sram_cell_6t_5 inst_cell_105_44 (.BL(BL44),.BLN(BLN44),.WL(WL105));
sram_cell_6t_5 inst_cell_105_45 (.BL(BL45),.BLN(BLN45),.WL(WL105));
sram_cell_6t_5 inst_cell_105_46 (.BL(BL46),.BLN(BLN46),.WL(WL105));
sram_cell_6t_5 inst_cell_105_47 (.BL(BL47),.BLN(BLN47),.WL(WL105));
sram_cell_6t_5 inst_cell_105_48 (.BL(BL48),.BLN(BLN48),.WL(WL105));
sram_cell_6t_5 inst_cell_105_49 (.BL(BL49),.BLN(BLN49),.WL(WL105));
sram_cell_6t_5 inst_cell_105_50 (.BL(BL50),.BLN(BLN50),.WL(WL105));
sram_cell_6t_5 inst_cell_105_51 (.BL(BL51),.BLN(BLN51),.WL(WL105));
sram_cell_6t_5 inst_cell_105_52 (.BL(BL52),.BLN(BLN52),.WL(WL105));
sram_cell_6t_5 inst_cell_105_53 (.BL(BL53),.BLN(BLN53),.WL(WL105));
sram_cell_6t_5 inst_cell_105_54 (.BL(BL54),.BLN(BLN54),.WL(WL105));
sram_cell_6t_5 inst_cell_105_55 (.BL(BL55),.BLN(BLN55),.WL(WL105));
sram_cell_6t_5 inst_cell_105_56 (.BL(BL56),.BLN(BLN56),.WL(WL105));
sram_cell_6t_5 inst_cell_105_57 (.BL(BL57),.BLN(BLN57),.WL(WL105));
sram_cell_6t_5 inst_cell_105_58 (.BL(BL58),.BLN(BLN58),.WL(WL105));
sram_cell_6t_5 inst_cell_105_59 (.BL(BL59),.BLN(BLN59),.WL(WL105));
sram_cell_6t_5 inst_cell_105_60 (.BL(BL60),.BLN(BLN60),.WL(WL105));
sram_cell_6t_5 inst_cell_105_61 (.BL(BL61),.BLN(BLN61),.WL(WL105));
sram_cell_6t_5 inst_cell_105_62 (.BL(BL62),.BLN(BLN62),.WL(WL105));
sram_cell_6t_5 inst_cell_105_63 (.BL(BL63),.BLN(BLN63),.WL(WL105));
sram_cell_6t_5 inst_cell_105_64 (.BL(BL64),.BLN(BLN64),.WL(WL105));
sram_cell_6t_5 inst_cell_105_65 (.BL(BL65),.BLN(BLN65),.WL(WL105));
sram_cell_6t_5 inst_cell_105_66 (.BL(BL66),.BLN(BLN66),.WL(WL105));
sram_cell_6t_5 inst_cell_105_67 (.BL(BL67),.BLN(BLN67),.WL(WL105));
sram_cell_6t_5 inst_cell_105_68 (.BL(BL68),.BLN(BLN68),.WL(WL105));
sram_cell_6t_5 inst_cell_105_69 (.BL(BL69),.BLN(BLN69),.WL(WL105));
sram_cell_6t_5 inst_cell_105_70 (.BL(BL70),.BLN(BLN70),.WL(WL105));
sram_cell_6t_5 inst_cell_105_71 (.BL(BL71),.BLN(BLN71),.WL(WL105));
sram_cell_6t_5 inst_cell_105_72 (.BL(BL72),.BLN(BLN72),.WL(WL105));
sram_cell_6t_5 inst_cell_105_73 (.BL(BL73),.BLN(BLN73),.WL(WL105));
sram_cell_6t_5 inst_cell_105_74 (.BL(BL74),.BLN(BLN74),.WL(WL105));
sram_cell_6t_5 inst_cell_105_75 (.BL(BL75),.BLN(BLN75),.WL(WL105));
sram_cell_6t_5 inst_cell_105_76 (.BL(BL76),.BLN(BLN76),.WL(WL105));
sram_cell_6t_5 inst_cell_105_77 (.BL(BL77),.BLN(BLN77),.WL(WL105));
sram_cell_6t_5 inst_cell_105_78 (.BL(BL78),.BLN(BLN78),.WL(WL105));
sram_cell_6t_5 inst_cell_105_79 (.BL(BL79),.BLN(BLN79),.WL(WL105));
sram_cell_6t_5 inst_cell_105_80 (.BL(BL80),.BLN(BLN80),.WL(WL105));
sram_cell_6t_5 inst_cell_105_81 (.BL(BL81),.BLN(BLN81),.WL(WL105));
sram_cell_6t_5 inst_cell_105_82 (.BL(BL82),.BLN(BLN82),.WL(WL105));
sram_cell_6t_5 inst_cell_105_83 (.BL(BL83),.BLN(BLN83),.WL(WL105));
sram_cell_6t_5 inst_cell_105_84 (.BL(BL84),.BLN(BLN84),.WL(WL105));
sram_cell_6t_5 inst_cell_105_85 (.BL(BL85),.BLN(BLN85),.WL(WL105));
sram_cell_6t_5 inst_cell_105_86 (.BL(BL86),.BLN(BLN86),.WL(WL105));
sram_cell_6t_5 inst_cell_105_87 (.BL(BL87),.BLN(BLN87),.WL(WL105));
sram_cell_6t_5 inst_cell_105_88 (.BL(BL88),.BLN(BLN88),.WL(WL105));
sram_cell_6t_5 inst_cell_105_89 (.BL(BL89),.BLN(BLN89),.WL(WL105));
sram_cell_6t_5 inst_cell_105_90 (.BL(BL90),.BLN(BLN90),.WL(WL105));
sram_cell_6t_5 inst_cell_105_91 (.BL(BL91),.BLN(BLN91),.WL(WL105));
sram_cell_6t_5 inst_cell_105_92 (.BL(BL92),.BLN(BLN92),.WL(WL105));
sram_cell_6t_5 inst_cell_105_93 (.BL(BL93),.BLN(BLN93),.WL(WL105));
sram_cell_6t_5 inst_cell_105_94 (.BL(BL94),.BLN(BLN94),.WL(WL105));
sram_cell_6t_5 inst_cell_105_95 (.BL(BL95),.BLN(BLN95),.WL(WL105));
sram_cell_6t_5 inst_cell_105_96 (.BL(BL96),.BLN(BLN96),.WL(WL105));
sram_cell_6t_5 inst_cell_105_97 (.BL(BL97),.BLN(BLN97),.WL(WL105));
sram_cell_6t_5 inst_cell_105_98 (.BL(BL98),.BLN(BLN98),.WL(WL105));
sram_cell_6t_5 inst_cell_105_99 (.BL(BL99),.BLN(BLN99),.WL(WL105));
sram_cell_6t_5 inst_cell_105_100 (.BL(BL100),.BLN(BLN100),.WL(WL105));
sram_cell_6t_5 inst_cell_105_101 (.BL(BL101),.BLN(BLN101),.WL(WL105));
sram_cell_6t_5 inst_cell_105_102 (.BL(BL102),.BLN(BLN102),.WL(WL105));
sram_cell_6t_5 inst_cell_105_103 (.BL(BL103),.BLN(BLN103),.WL(WL105));
sram_cell_6t_5 inst_cell_105_104 (.BL(BL104),.BLN(BLN104),.WL(WL105));
sram_cell_6t_5 inst_cell_105_105 (.BL(BL105),.BLN(BLN105),.WL(WL105));
sram_cell_6t_5 inst_cell_105_106 (.BL(BL106),.BLN(BLN106),.WL(WL105));
sram_cell_6t_5 inst_cell_105_107 (.BL(BL107),.BLN(BLN107),.WL(WL105));
sram_cell_6t_5 inst_cell_105_108 (.BL(BL108),.BLN(BLN108),.WL(WL105));
sram_cell_6t_5 inst_cell_105_109 (.BL(BL109),.BLN(BLN109),.WL(WL105));
sram_cell_6t_5 inst_cell_105_110 (.BL(BL110),.BLN(BLN110),.WL(WL105));
sram_cell_6t_5 inst_cell_105_111 (.BL(BL111),.BLN(BLN111),.WL(WL105));
sram_cell_6t_5 inst_cell_105_112 (.BL(BL112),.BLN(BLN112),.WL(WL105));
sram_cell_6t_5 inst_cell_105_113 (.BL(BL113),.BLN(BLN113),.WL(WL105));
sram_cell_6t_5 inst_cell_105_114 (.BL(BL114),.BLN(BLN114),.WL(WL105));
sram_cell_6t_5 inst_cell_105_115 (.BL(BL115),.BLN(BLN115),.WL(WL105));
sram_cell_6t_5 inst_cell_105_116 (.BL(BL116),.BLN(BLN116),.WL(WL105));
sram_cell_6t_5 inst_cell_105_117 (.BL(BL117),.BLN(BLN117),.WL(WL105));
sram_cell_6t_5 inst_cell_105_118 (.BL(BL118),.BLN(BLN118),.WL(WL105));
sram_cell_6t_5 inst_cell_105_119 (.BL(BL119),.BLN(BLN119),.WL(WL105));
sram_cell_6t_5 inst_cell_105_120 (.BL(BL120),.BLN(BLN120),.WL(WL105));
sram_cell_6t_5 inst_cell_105_121 (.BL(BL121),.BLN(BLN121),.WL(WL105));
sram_cell_6t_5 inst_cell_105_122 (.BL(BL122),.BLN(BLN122),.WL(WL105));
sram_cell_6t_5 inst_cell_105_123 (.BL(BL123),.BLN(BLN123),.WL(WL105));
sram_cell_6t_5 inst_cell_105_124 (.BL(BL124),.BLN(BLN124),.WL(WL105));
sram_cell_6t_5 inst_cell_105_125 (.BL(BL125),.BLN(BLN125),.WL(WL105));
sram_cell_6t_5 inst_cell_105_126 (.BL(BL126),.BLN(BLN126),.WL(WL105));
sram_cell_6t_5 inst_cell_105_127 (.BL(BL127),.BLN(BLN127),.WL(WL105));
sram_cell_6t_5 inst_cell_106_0 (.BL(BL0),.BLN(BLN0),.WL(WL106));
sram_cell_6t_5 inst_cell_106_1 (.BL(BL1),.BLN(BLN1),.WL(WL106));
sram_cell_6t_5 inst_cell_106_2 (.BL(BL2),.BLN(BLN2),.WL(WL106));
sram_cell_6t_5 inst_cell_106_3 (.BL(BL3),.BLN(BLN3),.WL(WL106));
sram_cell_6t_5 inst_cell_106_4 (.BL(BL4),.BLN(BLN4),.WL(WL106));
sram_cell_6t_5 inst_cell_106_5 (.BL(BL5),.BLN(BLN5),.WL(WL106));
sram_cell_6t_5 inst_cell_106_6 (.BL(BL6),.BLN(BLN6),.WL(WL106));
sram_cell_6t_5 inst_cell_106_7 (.BL(BL7),.BLN(BLN7),.WL(WL106));
sram_cell_6t_5 inst_cell_106_8 (.BL(BL8),.BLN(BLN8),.WL(WL106));
sram_cell_6t_5 inst_cell_106_9 (.BL(BL9),.BLN(BLN9),.WL(WL106));
sram_cell_6t_5 inst_cell_106_10 (.BL(BL10),.BLN(BLN10),.WL(WL106));
sram_cell_6t_5 inst_cell_106_11 (.BL(BL11),.BLN(BLN11),.WL(WL106));
sram_cell_6t_5 inst_cell_106_12 (.BL(BL12),.BLN(BLN12),.WL(WL106));
sram_cell_6t_5 inst_cell_106_13 (.BL(BL13),.BLN(BLN13),.WL(WL106));
sram_cell_6t_5 inst_cell_106_14 (.BL(BL14),.BLN(BLN14),.WL(WL106));
sram_cell_6t_5 inst_cell_106_15 (.BL(BL15),.BLN(BLN15),.WL(WL106));
sram_cell_6t_5 inst_cell_106_16 (.BL(BL16),.BLN(BLN16),.WL(WL106));
sram_cell_6t_5 inst_cell_106_17 (.BL(BL17),.BLN(BLN17),.WL(WL106));
sram_cell_6t_5 inst_cell_106_18 (.BL(BL18),.BLN(BLN18),.WL(WL106));
sram_cell_6t_5 inst_cell_106_19 (.BL(BL19),.BLN(BLN19),.WL(WL106));
sram_cell_6t_5 inst_cell_106_20 (.BL(BL20),.BLN(BLN20),.WL(WL106));
sram_cell_6t_5 inst_cell_106_21 (.BL(BL21),.BLN(BLN21),.WL(WL106));
sram_cell_6t_5 inst_cell_106_22 (.BL(BL22),.BLN(BLN22),.WL(WL106));
sram_cell_6t_5 inst_cell_106_23 (.BL(BL23),.BLN(BLN23),.WL(WL106));
sram_cell_6t_5 inst_cell_106_24 (.BL(BL24),.BLN(BLN24),.WL(WL106));
sram_cell_6t_5 inst_cell_106_25 (.BL(BL25),.BLN(BLN25),.WL(WL106));
sram_cell_6t_5 inst_cell_106_26 (.BL(BL26),.BLN(BLN26),.WL(WL106));
sram_cell_6t_5 inst_cell_106_27 (.BL(BL27),.BLN(BLN27),.WL(WL106));
sram_cell_6t_5 inst_cell_106_28 (.BL(BL28),.BLN(BLN28),.WL(WL106));
sram_cell_6t_5 inst_cell_106_29 (.BL(BL29),.BLN(BLN29),.WL(WL106));
sram_cell_6t_5 inst_cell_106_30 (.BL(BL30),.BLN(BLN30),.WL(WL106));
sram_cell_6t_5 inst_cell_106_31 (.BL(BL31),.BLN(BLN31),.WL(WL106));
sram_cell_6t_5 inst_cell_106_32 (.BL(BL32),.BLN(BLN32),.WL(WL106));
sram_cell_6t_5 inst_cell_106_33 (.BL(BL33),.BLN(BLN33),.WL(WL106));
sram_cell_6t_5 inst_cell_106_34 (.BL(BL34),.BLN(BLN34),.WL(WL106));
sram_cell_6t_5 inst_cell_106_35 (.BL(BL35),.BLN(BLN35),.WL(WL106));
sram_cell_6t_5 inst_cell_106_36 (.BL(BL36),.BLN(BLN36),.WL(WL106));
sram_cell_6t_5 inst_cell_106_37 (.BL(BL37),.BLN(BLN37),.WL(WL106));
sram_cell_6t_5 inst_cell_106_38 (.BL(BL38),.BLN(BLN38),.WL(WL106));
sram_cell_6t_5 inst_cell_106_39 (.BL(BL39),.BLN(BLN39),.WL(WL106));
sram_cell_6t_5 inst_cell_106_40 (.BL(BL40),.BLN(BLN40),.WL(WL106));
sram_cell_6t_5 inst_cell_106_41 (.BL(BL41),.BLN(BLN41),.WL(WL106));
sram_cell_6t_5 inst_cell_106_42 (.BL(BL42),.BLN(BLN42),.WL(WL106));
sram_cell_6t_5 inst_cell_106_43 (.BL(BL43),.BLN(BLN43),.WL(WL106));
sram_cell_6t_5 inst_cell_106_44 (.BL(BL44),.BLN(BLN44),.WL(WL106));
sram_cell_6t_5 inst_cell_106_45 (.BL(BL45),.BLN(BLN45),.WL(WL106));
sram_cell_6t_5 inst_cell_106_46 (.BL(BL46),.BLN(BLN46),.WL(WL106));
sram_cell_6t_5 inst_cell_106_47 (.BL(BL47),.BLN(BLN47),.WL(WL106));
sram_cell_6t_5 inst_cell_106_48 (.BL(BL48),.BLN(BLN48),.WL(WL106));
sram_cell_6t_5 inst_cell_106_49 (.BL(BL49),.BLN(BLN49),.WL(WL106));
sram_cell_6t_5 inst_cell_106_50 (.BL(BL50),.BLN(BLN50),.WL(WL106));
sram_cell_6t_5 inst_cell_106_51 (.BL(BL51),.BLN(BLN51),.WL(WL106));
sram_cell_6t_5 inst_cell_106_52 (.BL(BL52),.BLN(BLN52),.WL(WL106));
sram_cell_6t_5 inst_cell_106_53 (.BL(BL53),.BLN(BLN53),.WL(WL106));
sram_cell_6t_5 inst_cell_106_54 (.BL(BL54),.BLN(BLN54),.WL(WL106));
sram_cell_6t_5 inst_cell_106_55 (.BL(BL55),.BLN(BLN55),.WL(WL106));
sram_cell_6t_5 inst_cell_106_56 (.BL(BL56),.BLN(BLN56),.WL(WL106));
sram_cell_6t_5 inst_cell_106_57 (.BL(BL57),.BLN(BLN57),.WL(WL106));
sram_cell_6t_5 inst_cell_106_58 (.BL(BL58),.BLN(BLN58),.WL(WL106));
sram_cell_6t_5 inst_cell_106_59 (.BL(BL59),.BLN(BLN59),.WL(WL106));
sram_cell_6t_5 inst_cell_106_60 (.BL(BL60),.BLN(BLN60),.WL(WL106));
sram_cell_6t_5 inst_cell_106_61 (.BL(BL61),.BLN(BLN61),.WL(WL106));
sram_cell_6t_5 inst_cell_106_62 (.BL(BL62),.BLN(BLN62),.WL(WL106));
sram_cell_6t_5 inst_cell_106_63 (.BL(BL63),.BLN(BLN63),.WL(WL106));
sram_cell_6t_5 inst_cell_106_64 (.BL(BL64),.BLN(BLN64),.WL(WL106));
sram_cell_6t_5 inst_cell_106_65 (.BL(BL65),.BLN(BLN65),.WL(WL106));
sram_cell_6t_5 inst_cell_106_66 (.BL(BL66),.BLN(BLN66),.WL(WL106));
sram_cell_6t_5 inst_cell_106_67 (.BL(BL67),.BLN(BLN67),.WL(WL106));
sram_cell_6t_5 inst_cell_106_68 (.BL(BL68),.BLN(BLN68),.WL(WL106));
sram_cell_6t_5 inst_cell_106_69 (.BL(BL69),.BLN(BLN69),.WL(WL106));
sram_cell_6t_5 inst_cell_106_70 (.BL(BL70),.BLN(BLN70),.WL(WL106));
sram_cell_6t_5 inst_cell_106_71 (.BL(BL71),.BLN(BLN71),.WL(WL106));
sram_cell_6t_5 inst_cell_106_72 (.BL(BL72),.BLN(BLN72),.WL(WL106));
sram_cell_6t_5 inst_cell_106_73 (.BL(BL73),.BLN(BLN73),.WL(WL106));
sram_cell_6t_5 inst_cell_106_74 (.BL(BL74),.BLN(BLN74),.WL(WL106));
sram_cell_6t_5 inst_cell_106_75 (.BL(BL75),.BLN(BLN75),.WL(WL106));
sram_cell_6t_5 inst_cell_106_76 (.BL(BL76),.BLN(BLN76),.WL(WL106));
sram_cell_6t_5 inst_cell_106_77 (.BL(BL77),.BLN(BLN77),.WL(WL106));
sram_cell_6t_5 inst_cell_106_78 (.BL(BL78),.BLN(BLN78),.WL(WL106));
sram_cell_6t_5 inst_cell_106_79 (.BL(BL79),.BLN(BLN79),.WL(WL106));
sram_cell_6t_5 inst_cell_106_80 (.BL(BL80),.BLN(BLN80),.WL(WL106));
sram_cell_6t_5 inst_cell_106_81 (.BL(BL81),.BLN(BLN81),.WL(WL106));
sram_cell_6t_5 inst_cell_106_82 (.BL(BL82),.BLN(BLN82),.WL(WL106));
sram_cell_6t_5 inst_cell_106_83 (.BL(BL83),.BLN(BLN83),.WL(WL106));
sram_cell_6t_5 inst_cell_106_84 (.BL(BL84),.BLN(BLN84),.WL(WL106));
sram_cell_6t_5 inst_cell_106_85 (.BL(BL85),.BLN(BLN85),.WL(WL106));
sram_cell_6t_5 inst_cell_106_86 (.BL(BL86),.BLN(BLN86),.WL(WL106));
sram_cell_6t_5 inst_cell_106_87 (.BL(BL87),.BLN(BLN87),.WL(WL106));
sram_cell_6t_5 inst_cell_106_88 (.BL(BL88),.BLN(BLN88),.WL(WL106));
sram_cell_6t_5 inst_cell_106_89 (.BL(BL89),.BLN(BLN89),.WL(WL106));
sram_cell_6t_5 inst_cell_106_90 (.BL(BL90),.BLN(BLN90),.WL(WL106));
sram_cell_6t_5 inst_cell_106_91 (.BL(BL91),.BLN(BLN91),.WL(WL106));
sram_cell_6t_5 inst_cell_106_92 (.BL(BL92),.BLN(BLN92),.WL(WL106));
sram_cell_6t_5 inst_cell_106_93 (.BL(BL93),.BLN(BLN93),.WL(WL106));
sram_cell_6t_5 inst_cell_106_94 (.BL(BL94),.BLN(BLN94),.WL(WL106));
sram_cell_6t_5 inst_cell_106_95 (.BL(BL95),.BLN(BLN95),.WL(WL106));
sram_cell_6t_5 inst_cell_106_96 (.BL(BL96),.BLN(BLN96),.WL(WL106));
sram_cell_6t_5 inst_cell_106_97 (.BL(BL97),.BLN(BLN97),.WL(WL106));
sram_cell_6t_5 inst_cell_106_98 (.BL(BL98),.BLN(BLN98),.WL(WL106));
sram_cell_6t_5 inst_cell_106_99 (.BL(BL99),.BLN(BLN99),.WL(WL106));
sram_cell_6t_5 inst_cell_106_100 (.BL(BL100),.BLN(BLN100),.WL(WL106));
sram_cell_6t_5 inst_cell_106_101 (.BL(BL101),.BLN(BLN101),.WL(WL106));
sram_cell_6t_5 inst_cell_106_102 (.BL(BL102),.BLN(BLN102),.WL(WL106));
sram_cell_6t_5 inst_cell_106_103 (.BL(BL103),.BLN(BLN103),.WL(WL106));
sram_cell_6t_5 inst_cell_106_104 (.BL(BL104),.BLN(BLN104),.WL(WL106));
sram_cell_6t_5 inst_cell_106_105 (.BL(BL105),.BLN(BLN105),.WL(WL106));
sram_cell_6t_5 inst_cell_106_106 (.BL(BL106),.BLN(BLN106),.WL(WL106));
sram_cell_6t_5 inst_cell_106_107 (.BL(BL107),.BLN(BLN107),.WL(WL106));
sram_cell_6t_5 inst_cell_106_108 (.BL(BL108),.BLN(BLN108),.WL(WL106));
sram_cell_6t_5 inst_cell_106_109 (.BL(BL109),.BLN(BLN109),.WL(WL106));
sram_cell_6t_5 inst_cell_106_110 (.BL(BL110),.BLN(BLN110),.WL(WL106));
sram_cell_6t_5 inst_cell_106_111 (.BL(BL111),.BLN(BLN111),.WL(WL106));
sram_cell_6t_5 inst_cell_106_112 (.BL(BL112),.BLN(BLN112),.WL(WL106));
sram_cell_6t_5 inst_cell_106_113 (.BL(BL113),.BLN(BLN113),.WL(WL106));
sram_cell_6t_5 inst_cell_106_114 (.BL(BL114),.BLN(BLN114),.WL(WL106));
sram_cell_6t_5 inst_cell_106_115 (.BL(BL115),.BLN(BLN115),.WL(WL106));
sram_cell_6t_5 inst_cell_106_116 (.BL(BL116),.BLN(BLN116),.WL(WL106));
sram_cell_6t_5 inst_cell_106_117 (.BL(BL117),.BLN(BLN117),.WL(WL106));
sram_cell_6t_5 inst_cell_106_118 (.BL(BL118),.BLN(BLN118),.WL(WL106));
sram_cell_6t_5 inst_cell_106_119 (.BL(BL119),.BLN(BLN119),.WL(WL106));
sram_cell_6t_5 inst_cell_106_120 (.BL(BL120),.BLN(BLN120),.WL(WL106));
sram_cell_6t_5 inst_cell_106_121 (.BL(BL121),.BLN(BLN121),.WL(WL106));
sram_cell_6t_5 inst_cell_106_122 (.BL(BL122),.BLN(BLN122),.WL(WL106));
sram_cell_6t_5 inst_cell_106_123 (.BL(BL123),.BLN(BLN123),.WL(WL106));
sram_cell_6t_5 inst_cell_106_124 (.BL(BL124),.BLN(BLN124),.WL(WL106));
sram_cell_6t_5 inst_cell_106_125 (.BL(BL125),.BLN(BLN125),.WL(WL106));
sram_cell_6t_5 inst_cell_106_126 (.BL(BL126),.BLN(BLN126),.WL(WL106));
sram_cell_6t_5 inst_cell_106_127 (.BL(BL127),.BLN(BLN127),.WL(WL106));
sram_cell_6t_5 inst_cell_107_0 (.BL(BL0),.BLN(BLN0),.WL(WL107));
sram_cell_6t_5 inst_cell_107_1 (.BL(BL1),.BLN(BLN1),.WL(WL107));
sram_cell_6t_5 inst_cell_107_2 (.BL(BL2),.BLN(BLN2),.WL(WL107));
sram_cell_6t_5 inst_cell_107_3 (.BL(BL3),.BLN(BLN3),.WL(WL107));
sram_cell_6t_5 inst_cell_107_4 (.BL(BL4),.BLN(BLN4),.WL(WL107));
sram_cell_6t_5 inst_cell_107_5 (.BL(BL5),.BLN(BLN5),.WL(WL107));
sram_cell_6t_5 inst_cell_107_6 (.BL(BL6),.BLN(BLN6),.WL(WL107));
sram_cell_6t_5 inst_cell_107_7 (.BL(BL7),.BLN(BLN7),.WL(WL107));
sram_cell_6t_5 inst_cell_107_8 (.BL(BL8),.BLN(BLN8),.WL(WL107));
sram_cell_6t_5 inst_cell_107_9 (.BL(BL9),.BLN(BLN9),.WL(WL107));
sram_cell_6t_5 inst_cell_107_10 (.BL(BL10),.BLN(BLN10),.WL(WL107));
sram_cell_6t_5 inst_cell_107_11 (.BL(BL11),.BLN(BLN11),.WL(WL107));
sram_cell_6t_5 inst_cell_107_12 (.BL(BL12),.BLN(BLN12),.WL(WL107));
sram_cell_6t_5 inst_cell_107_13 (.BL(BL13),.BLN(BLN13),.WL(WL107));
sram_cell_6t_5 inst_cell_107_14 (.BL(BL14),.BLN(BLN14),.WL(WL107));
sram_cell_6t_5 inst_cell_107_15 (.BL(BL15),.BLN(BLN15),.WL(WL107));
sram_cell_6t_5 inst_cell_107_16 (.BL(BL16),.BLN(BLN16),.WL(WL107));
sram_cell_6t_5 inst_cell_107_17 (.BL(BL17),.BLN(BLN17),.WL(WL107));
sram_cell_6t_5 inst_cell_107_18 (.BL(BL18),.BLN(BLN18),.WL(WL107));
sram_cell_6t_5 inst_cell_107_19 (.BL(BL19),.BLN(BLN19),.WL(WL107));
sram_cell_6t_5 inst_cell_107_20 (.BL(BL20),.BLN(BLN20),.WL(WL107));
sram_cell_6t_5 inst_cell_107_21 (.BL(BL21),.BLN(BLN21),.WL(WL107));
sram_cell_6t_5 inst_cell_107_22 (.BL(BL22),.BLN(BLN22),.WL(WL107));
sram_cell_6t_5 inst_cell_107_23 (.BL(BL23),.BLN(BLN23),.WL(WL107));
sram_cell_6t_5 inst_cell_107_24 (.BL(BL24),.BLN(BLN24),.WL(WL107));
sram_cell_6t_5 inst_cell_107_25 (.BL(BL25),.BLN(BLN25),.WL(WL107));
sram_cell_6t_5 inst_cell_107_26 (.BL(BL26),.BLN(BLN26),.WL(WL107));
sram_cell_6t_5 inst_cell_107_27 (.BL(BL27),.BLN(BLN27),.WL(WL107));
sram_cell_6t_5 inst_cell_107_28 (.BL(BL28),.BLN(BLN28),.WL(WL107));
sram_cell_6t_5 inst_cell_107_29 (.BL(BL29),.BLN(BLN29),.WL(WL107));
sram_cell_6t_5 inst_cell_107_30 (.BL(BL30),.BLN(BLN30),.WL(WL107));
sram_cell_6t_5 inst_cell_107_31 (.BL(BL31),.BLN(BLN31),.WL(WL107));
sram_cell_6t_5 inst_cell_107_32 (.BL(BL32),.BLN(BLN32),.WL(WL107));
sram_cell_6t_5 inst_cell_107_33 (.BL(BL33),.BLN(BLN33),.WL(WL107));
sram_cell_6t_5 inst_cell_107_34 (.BL(BL34),.BLN(BLN34),.WL(WL107));
sram_cell_6t_5 inst_cell_107_35 (.BL(BL35),.BLN(BLN35),.WL(WL107));
sram_cell_6t_5 inst_cell_107_36 (.BL(BL36),.BLN(BLN36),.WL(WL107));
sram_cell_6t_5 inst_cell_107_37 (.BL(BL37),.BLN(BLN37),.WL(WL107));
sram_cell_6t_5 inst_cell_107_38 (.BL(BL38),.BLN(BLN38),.WL(WL107));
sram_cell_6t_5 inst_cell_107_39 (.BL(BL39),.BLN(BLN39),.WL(WL107));
sram_cell_6t_5 inst_cell_107_40 (.BL(BL40),.BLN(BLN40),.WL(WL107));
sram_cell_6t_5 inst_cell_107_41 (.BL(BL41),.BLN(BLN41),.WL(WL107));
sram_cell_6t_5 inst_cell_107_42 (.BL(BL42),.BLN(BLN42),.WL(WL107));
sram_cell_6t_5 inst_cell_107_43 (.BL(BL43),.BLN(BLN43),.WL(WL107));
sram_cell_6t_5 inst_cell_107_44 (.BL(BL44),.BLN(BLN44),.WL(WL107));
sram_cell_6t_5 inst_cell_107_45 (.BL(BL45),.BLN(BLN45),.WL(WL107));
sram_cell_6t_5 inst_cell_107_46 (.BL(BL46),.BLN(BLN46),.WL(WL107));
sram_cell_6t_5 inst_cell_107_47 (.BL(BL47),.BLN(BLN47),.WL(WL107));
sram_cell_6t_5 inst_cell_107_48 (.BL(BL48),.BLN(BLN48),.WL(WL107));
sram_cell_6t_5 inst_cell_107_49 (.BL(BL49),.BLN(BLN49),.WL(WL107));
sram_cell_6t_5 inst_cell_107_50 (.BL(BL50),.BLN(BLN50),.WL(WL107));
sram_cell_6t_5 inst_cell_107_51 (.BL(BL51),.BLN(BLN51),.WL(WL107));
sram_cell_6t_5 inst_cell_107_52 (.BL(BL52),.BLN(BLN52),.WL(WL107));
sram_cell_6t_5 inst_cell_107_53 (.BL(BL53),.BLN(BLN53),.WL(WL107));
sram_cell_6t_5 inst_cell_107_54 (.BL(BL54),.BLN(BLN54),.WL(WL107));
sram_cell_6t_5 inst_cell_107_55 (.BL(BL55),.BLN(BLN55),.WL(WL107));
sram_cell_6t_5 inst_cell_107_56 (.BL(BL56),.BLN(BLN56),.WL(WL107));
sram_cell_6t_5 inst_cell_107_57 (.BL(BL57),.BLN(BLN57),.WL(WL107));
sram_cell_6t_5 inst_cell_107_58 (.BL(BL58),.BLN(BLN58),.WL(WL107));
sram_cell_6t_5 inst_cell_107_59 (.BL(BL59),.BLN(BLN59),.WL(WL107));
sram_cell_6t_5 inst_cell_107_60 (.BL(BL60),.BLN(BLN60),.WL(WL107));
sram_cell_6t_5 inst_cell_107_61 (.BL(BL61),.BLN(BLN61),.WL(WL107));
sram_cell_6t_5 inst_cell_107_62 (.BL(BL62),.BLN(BLN62),.WL(WL107));
sram_cell_6t_5 inst_cell_107_63 (.BL(BL63),.BLN(BLN63),.WL(WL107));
sram_cell_6t_5 inst_cell_107_64 (.BL(BL64),.BLN(BLN64),.WL(WL107));
sram_cell_6t_5 inst_cell_107_65 (.BL(BL65),.BLN(BLN65),.WL(WL107));
sram_cell_6t_5 inst_cell_107_66 (.BL(BL66),.BLN(BLN66),.WL(WL107));
sram_cell_6t_5 inst_cell_107_67 (.BL(BL67),.BLN(BLN67),.WL(WL107));
sram_cell_6t_5 inst_cell_107_68 (.BL(BL68),.BLN(BLN68),.WL(WL107));
sram_cell_6t_5 inst_cell_107_69 (.BL(BL69),.BLN(BLN69),.WL(WL107));
sram_cell_6t_5 inst_cell_107_70 (.BL(BL70),.BLN(BLN70),.WL(WL107));
sram_cell_6t_5 inst_cell_107_71 (.BL(BL71),.BLN(BLN71),.WL(WL107));
sram_cell_6t_5 inst_cell_107_72 (.BL(BL72),.BLN(BLN72),.WL(WL107));
sram_cell_6t_5 inst_cell_107_73 (.BL(BL73),.BLN(BLN73),.WL(WL107));
sram_cell_6t_5 inst_cell_107_74 (.BL(BL74),.BLN(BLN74),.WL(WL107));
sram_cell_6t_5 inst_cell_107_75 (.BL(BL75),.BLN(BLN75),.WL(WL107));
sram_cell_6t_5 inst_cell_107_76 (.BL(BL76),.BLN(BLN76),.WL(WL107));
sram_cell_6t_5 inst_cell_107_77 (.BL(BL77),.BLN(BLN77),.WL(WL107));
sram_cell_6t_5 inst_cell_107_78 (.BL(BL78),.BLN(BLN78),.WL(WL107));
sram_cell_6t_5 inst_cell_107_79 (.BL(BL79),.BLN(BLN79),.WL(WL107));
sram_cell_6t_5 inst_cell_107_80 (.BL(BL80),.BLN(BLN80),.WL(WL107));
sram_cell_6t_5 inst_cell_107_81 (.BL(BL81),.BLN(BLN81),.WL(WL107));
sram_cell_6t_5 inst_cell_107_82 (.BL(BL82),.BLN(BLN82),.WL(WL107));
sram_cell_6t_5 inst_cell_107_83 (.BL(BL83),.BLN(BLN83),.WL(WL107));
sram_cell_6t_5 inst_cell_107_84 (.BL(BL84),.BLN(BLN84),.WL(WL107));
sram_cell_6t_5 inst_cell_107_85 (.BL(BL85),.BLN(BLN85),.WL(WL107));
sram_cell_6t_5 inst_cell_107_86 (.BL(BL86),.BLN(BLN86),.WL(WL107));
sram_cell_6t_5 inst_cell_107_87 (.BL(BL87),.BLN(BLN87),.WL(WL107));
sram_cell_6t_5 inst_cell_107_88 (.BL(BL88),.BLN(BLN88),.WL(WL107));
sram_cell_6t_5 inst_cell_107_89 (.BL(BL89),.BLN(BLN89),.WL(WL107));
sram_cell_6t_5 inst_cell_107_90 (.BL(BL90),.BLN(BLN90),.WL(WL107));
sram_cell_6t_5 inst_cell_107_91 (.BL(BL91),.BLN(BLN91),.WL(WL107));
sram_cell_6t_5 inst_cell_107_92 (.BL(BL92),.BLN(BLN92),.WL(WL107));
sram_cell_6t_5 inst_cell_107_93 (.BL(BL93),.BLN(BLN93),.WL(WL107));
sram_cell_6t_5 inst_cell_107_94 (.BL(BL94),.BLN(BLN94),.WL(WL107));
sram_cell_6t_5 inst_cell_107_95 (.BL(BL95),.BLN(BLN95),.WL(WL107));
sram_cell_6t_5 inst_cell_107_96 (.BL(BL96),.BLN(BLN96),.WL(WL107));
sram_cell_6t_5 inst_cell_107_97 (.BL(BL97),.BLN(BLN97),.WL(WL107));
sram_cell_6t_5 inst_cell_107_98 (.BL(BL98),.BLN(BLN98),.WL(WL107));
sram_cell_6t_5 inst_cell_107_99 (.BL(BL99),.BLN(BLN99),.WL(WL107));
sram_cell_6t_5 inst_cell_107_100 (.BL(BL100),.BLN(BLN100),.WL(WL107));
sram_cell_6t_5 inst_cell_107_101 (.BL(BL101),.BLN(BLN101),.WL(WL107));
sram_cell_6t_5 inst_cell_107_102 (.BL(BL102),.BLN(BLN102),.WL(WL107));
sram_cell_6t_5 inst_cell_107_103 (.BL(BL103),.BLN(BLN103),.WL(WL107));
sram_cell_6t_5 inst_cell_107_104 (.BL(BL104),.BLN(BLN104),.WL(WL107));
sram_cell_6t_5 inst_cell_107_105 (.BL(BL105),.BLN(BLN105),.WL(WL107));
sram_cell_6t_5 inst_cell_107_106 (.BL(BL106),.BLN(BLN106),.WL(WL107));
sram_cell_6t_5 inst_cell_107_107 (.BL(BL107),.BLN(BLN107),.WL(WL107));
sram_cell_6t_5 inst_cell_107_108 (.BL(BL108),.BLN(BLN108),.WL(WL107));
sram_cell_6t_5 inst_cell_107_109 (.BL(BL109),.BLN(BLN109),.WL(WL107));
sram_cell_6t_5 inst_cell_107_110 (.BL(BL110),.BLN(BLN110),.WL(WL107));
sram_cell_6t_5 inst_cell_107_111 (.BL(BL111),.BLN(BLN111),.WL(WL107));
sram_cell_6t_5 inst_cell_107_112 (.BL(BL112),.BLN(BLN112),.WL(WL107));
sram_cell_6t_5 inst_cell_107_113 (.BL(BL113),.BLN(BLN113),.WL(WL107));
sram_cell_6t_5 inst_cell_107_114 (.BL(BL114),.BLN(BLN114),.WL(WL107));
sram_cell_6t_5 inst_cell_107_115 (.BL(BL115),.BLN(BLN115),.WL(WL107));
sram_cell_6t_5 inst_cell_107_116 (.BL(BL116),.BLN(BLN116),.WL(WL107));
sram_cell_6t_5 inst_cell_107_117 (.BL(BL117),.BLN(BLN117),.WL(WL107));
sram_cell_6t_5 inst_cell_107_118 (.BL(BL118),.BLN(BLN118),.WL(WL107));
sram_cell_6t_5 inst_cell_107_119 (.BL(BL119),.BLN(BLN119),.WL(WL107));
sram_cell_6t_5 inst_cell_107_120 (.BL(BL120),.BLN(BLN120),.WL(WL107));
sram_cell_6t_5 inst_cell_107_121 (.BL(BL121),.BLN(BLN121),.WL(WL107));
sram_cell_6t_5 inst_cell_107_122 (.BL(BL122),.BLN(BLN122),.WL(WL107));
sram_cell_6t_5 inst_cell_107_123 (.BL(BL123),.BLN(BLN123),.WL(WL107));
sram_cell_6t_5 inst_cell_107_124 (.BL(BL124),.BLN(BLN124),.WL(WL107));
sram_cell_6t_5 inst_cell_107_125 (.BL(BL125),.BLN(BLN125),.WL(WL107));
sram_cell_6t_5 inst_cell_107_126 (.BL(BL126),.BLN(BLN126),.WL(WL107));
sram_cell_6t_5 inst_cell_107_127 (.BL(BL127),.BLN(BLN127),.WL(WL107));
sram_cell_6t_5 inst_cell_108_0 (.BL(BL0),.BLN(BLN0),.WL(WL108));
sram_cell_6t_5 inst_cell_108_1 (.BL(BL1),.BLN(BLN1),.WL(WL108));
sram_cell_6t_5 inst_cell_108_2 (.BL(BL2),.BLN(BLN2),.WL(WL108));
sram_cell_6t_5 inst_cell_108_3 (.BL(BL3),.BLN(BLN3),.WL(WL108));
sram_cell_6t_5 inst_cell_108_4 (.BL(BL4),.BLN(BLN4),.WL(WL108));
sram_cell_6t_5 inst_cell_108_5 (.BL(BL5),.BLN(BLN5),.WL(WL108));
sram_cell_6t_5 inst_cell_108_6 (.BL(BL6),.BLN(BLN6),.WL(WL108));
sram_cell_6t_5 inst_cell_108_7 (.BL(BL7),.BLN(BLN7),.WL(WL108));
sram_cell_6t_5 inst_cell_108_8 (.BL(BL8),.BLN(BLN8),.WL(WL108));
sram_cell_6t_5 inst_cell_108_9 (.BL(BL9),.BLN(BLN9),.WL(WL108));
sram_cell_6t_5 inst_cell_108_10 (.BL(BL10),.BLN(BLN10),.WL(WL108));
sram_cell_6t_5 inst_cell_108_11 (.BL(BL11),.BLN(BLN11),.WL(WL108));
sram_cell_6t_5 inst_cell_108_12 (.BL(BL12),.BLN(BLN12),.WL(WL108));
sram_cell_6t_5 inst_cell_108_13 (.BL(BL13),.BLN(BLN13),.WL(WL108));
sram_cell_6t_5 inst_cell_108_14 (.BL(BL14),.BLN(BLN14),.WL(WL108));
sram_cell_6t_5 inst_cell_108_15 (.BL(BL15),.BLN(BLN15),.WL(WL108));
sram_cell_6t_5 inst_cell_108_16 (.BL(BL16),.BLN(BLN16),.WL(WL108));
sram_cell_6t_5 inst_cell_108_17 (.BL(BL17),.BLN(BLN17),.WL(WL108));
sram_cell_6t_5 inst_cell_108_18 (.BL(BL18),.BLN(BLN18),.WL(WL108));
sram_cell_6t_5 inst_cell_108_19 (.BL(BL19),.BLN(BLN19),.WL(WL108));
sram_cell_6t_5 inst_cell_108_20 (.BL(BL20),.BLN(BLN20),.WL(WL108));
sram_cell_6t_5 inst_cell_108_21 (.BL(BL21),.BLN(BLN21),.WL(WL108));
sram_cell_6t_5 inst_cell_108_22 (.BL(BL22),.BLN(BLN22),.WL(WL108));
sram_cell_6t_5 inst_cell_108_23 (.BL(BL23),.BLN(BLN23),.WL(WL108));
sram_cell_6t_5 inst_cell_108_24 (.BL(BL24),.BLN(BLN24),.WL(WL108));
sram_cell_6t_5 inst_cell_108_25 (.BL(BL25),.BLN(BLN25),.WL(WL108));
sram_cell_6t_5 inst_cell_108_26 (.BL(BL26),.BLN(BLN26),.WL(WL108));
sram_cell_6t_5 inst_cell_108_27 (.BL(BL27),.BLN(BLN27),.WL(WL108));
sram_cell_6t_5 inst_cell_108_28 (.BL(BL28),.BLN(BLN28),.WL(WL108));
sram_cell_6t_5 inst_cell_108_29 (.BL(BL29),.BLN(BLN29),.WL(WL108));
sram_cell_6t_5 inst_cell_108_30 (.BL(BL30),.BLN(BLN30),.WL(WL108));
sram_cell_6t_5 inst_cell_108_31 (.BL(BL31),.BLN(BLN31),.WL(WL108));
sram_cell_6t_5 inst_cell_108_32 (.BL(BL32),.BLN(BLN32),.WL(WL108));
sram_cell_6t_5 inst_cell_108_33 (.BL(BL33),.BLN(BLN33),.WL(WL108));
sram_cell_6t_5 inst_cell_108_34 (.BL(BL34),.BLN(BLN34),.WL(WL108));
sram_cell_6t_5 inst_cell_108_35 (.BL(BL35),.BLN(BLN35),.WL(WL108));
sram_cell_6t_5 inst_cell_108_36 (.BL(BL36),.BLN(BLN36),.WL(WL108));
sram_cell_6t_5 inst_cell_108_37 (.BL(BL37),.BLN(BLN37),.WL(WL108));
sram_cell_6t_5 inst_cell_108_38 (.BL(BL38),.BLN(BLN38),.WL(WL108));
sram_cell_6t_5 inst_cell_108_39 (.BL(BL39),.BLN(BLN39),.WL(WL108));
sram_cell_6t_5 inst_cell_108_40 (.BL(BL40),.BLN(BLN40),.WL(WL108));
sram_cell_6t_5 inst_cell_108_41 (.BL(BL41),.BLN(BLN41),.WL(WL108));
sram_cell_6t_5 inst_cell_108_42 (.BL(BL42),.BLN(BLN42),.WL(WL108));
sram_cell_6t_5 inst_cell_108_43 (.BL(BL43),.BLN(BLN43),.WL(WL108));
sram_cell_6t_5 inst_cell_108_44 (.BL(BL44),.BLN(BLN44),.WL(WL108));
sram_cell_6t_5 inst_cell_108_45 (.BL(BL45),.BLN(BLN45),.WL(WL108));
sram_cell_6t_5 inst_cell_108_46 (.BL(BL46),.BLN(BLN46),.WL(WL108));
sram_cell_6t_5 inst_cell_108_47 (.BL(BL47),.BLN(BLN47),.WL(WL108));
sram_cell_6t_5 inst_cell_108_48 (.BL(BL48),.BLN(BLN48),.WL(WL108));
sram_cell_6t_5 inst_cell_108_49 (.BL(BL49),.BLN(BLN49),.WL(WL108));
sram_cell_6t_5 inst_cell_108_50 (.BL(BL50),.BLN(BLN50),.WL(WL108));
sram_cell_6t_5 inst_cell_108_51 (.BL(BL51),.BLN(BLN51),.WL(WL108));
sram_cell_6t_5 inst_cell_108_52 (.BL(BL52),.BLN(BLN52),.WL(WL108));
sram_cell_6t_5 inst_cell_108_53 (.BL(BL53),.BLN(BLN53),.WL(WL108));
sram_cell_6t_5 inst_cell_108_54 (.BL(BL54),.BLN(BLN54),.WL(WL108));
sram_cell_6t_5 inst_cell_108_55 (.BL(BL55),.BLN(BLN55),.WL(WL108));
sram_cell_6t_5 inst_cell_108_56 (.BL(BL56),.BLN(BLN56),.WL(WL108));
sram_cell_6t_5 inst_cell_108_57 (.BL(BL57),.BLN(BLN57),.WL(WL108));
sram_cell_6t_5 inst_cell_108_58 (.BL(BL58),.BLN(BLN58),.WL(WL108));
sram_cell_6t_5 inst_cell_108_59 (.BL(BL59),.BLN(BLN59),.WL(WL108));
sram_cell_6t_5 inst_cell_108_60 (.BL(BL60),.BLN(BLN60),.WL(WL108));
sram_cell_6t_5 inst_cell_108_61 (.BL(BL61),.BLN(BLN61),.WL(WL108));
sram_cell_6t_5 inst_cell_108_62 (.BL(BL62),.BLN(BLN62),.WL(WL108));
sram_cell_6t_5 inst_cell_108_63 (.BL(BL63),.BLN(BLN63),.WL(WL108));
sram_cell_6t_5 inst_cell_108_64 (.BL(BL64),.BLN(BLN64),.WL(WL108));
sram_cell_6t_5 inst_cell_108_65 (.BL(BL65),.BLN(BLN65),.WL(WL108));
sram_cell_6t_5 inst_cell_108_66 (.BL(BL66),.BLN(BLN66),.WL(WL108));
sram_cell_6t_5 inst_cell_108_67 (.BL(BL67),.BLN(BLN67),.WL(WL108));
sram_cell_6t_5 inst_cell_108_68 (.BL(BL68),.BLN(BLN68),.WL(WL108));
sram_cell_6t_5 inst_cell_108_69 (.BL(BL69),.BLN(BLN69),.WL(WL108));
sram_cell_6t_5 inst_cell_108_70 (.BL(BL70),.BLN(BLN70),.WL(WL108));
sram_cell_6t_5 inst_cell_108_71 (.BL(BL71),.BLN(BLN71),.WL(WL108));
sram_cell_6t_5 inst_cell_108_72 (.BL(BL72),.BLN(BLN72),.WL(WL108));
sram_cell_6t_5 inst_cell_108_73 (.BL(BL73),.BLN(BLN73),.WL(WL108));
sram_cell_6t_5 inst_cell_108_74 (.BL(BL74),.BLN(BLN74),.WL(WL108));
sram_cell_6t_5 inst_cell_108_75 (.BL(BL75),.BLN(BLN75),.WL(WL108));
sram_cell_6t_5 inst_cell_108_76 (.BL(BL76),.BLN(BLN76),.WL(WL108));
sram_cell_6t_5 inst_cell_108_77 (.BL(BL77),.BLN(BLN77),.WL(WL108));
sram_cell_6t_5 inst_cell_108_78 (.BL(BL78),.BLN(BLN78),.WL(WL108));
sram_cell_6t_5 inst_cell_108_79 (.BL(BL79),.BLN(BLN79),.WL(WL108));
sram_cell_6t_5 inst_cell_108_80 (.BL(BL80),.BLN(BLN80),.WL(WL108));
sram_cell_6t_5 inst_cell_108_81 (.BL(BL81),.BLN(BLN81),.WL(WL108));
sram_cell_6t_5 inst_cell_108_82 (.BL(BL82),.BLN(BLN82),.WL(WL108));
sram_cell_6t_5 inst_cell_108_83 (.BL(BL83),.BLN(BLN83),.WL(WL108));
sram_cell_6t_5 inst_cell_108_84 (.BL(BL84),.BLN(BLN84),.WL(WL108));
sram_cell_6t_5 inst_cell_108_85 (.BL(BL85),.BLN(BLN85),.WL(WL108));
sram_cell_6t_5 inst_cell_108_86 (.BL(BL86),.BLN(BLN86),.WL(WL108));
sram_cell_6t_5 inst_cell_108_87 (.BL(BL87),.BLN(BLN87),.WL(WL108));
sram_cell_6t_5 inst_cell_108_88 (.BL(BL88),.BLN(BLN88),.WL(WL108));
sram_cell_6t_5 inst_cell_108_89 (.BL(BL89),.BLN(BLN89),.WL(WL108));
sram_cell_6t_5 inst_cell_108_90 (.BL(BL90),.BLN(BLN90),.WL(WL108));
sram_cell_6t_5 inst_cell_108_91 (.BL(BL91),.BLN(BLN91),.WL(WL108));
sram_cell_6t_5 inst_cell_108_92 (.BL(BL92),.BLN(BLN92),.WL(WL108));
sram_cell_6t_5 inst_cell_108_93 (.BL(BL93),.BLN(BLN93),.WL(WL108));
sram_cell_6t_5 inst_cell_108_94 (.BL(BL94),.BLN(BLN94),.WL(WL108));
sram_cell_6t_5 inst_cell_108_95 (.BL(BL95),.BLN(BLN95),.WL(WL108));
sram_cell_6t_5 inst_cell_108_96 (.BL(BL96),.BLN(BLN96),.WL(WL108));
sram_cell_6t_5 inst_cell_108_97 (.BL(BL97),.BLN(BLN97),.WL(WL108));
sram_cell_6t_5 inst_cell_108_98 (.BL(BL98),.BLN(BLN98),.WL(WL108));
sram_cell_6t_5 inst_cell_108_99 (.BL(BL99),.BLN(BLN99),.WL(WL108));
sram_cell_6t_5 inst_cell_108_100 (.BL(BL100),.BLN(BLN100),.WL(WL108));
sram_cell_6t_5 inst_cell_108_101 (.BL(BL101),.BLN(BLN101),.WL(WL108));
sram_cell_6t_5 inst_cell_108_102 (.BL(BL102),.BLN(BLN102),.WL(WL108));
sram_cell_6t_5 inst_cell_108_103 (.BL(BL103),.BLN(BLN103),.WL(WL108));
sram_cell_6t_5 inst_cell_108_104 (.BL(BL104),.BLN(BLN104),.WL(WL108));
sram_cell_6t_5 inst_cell_108_105 (.BL(BL105),.BLN(BLN105),.WL(WL108));
sram_cell_6t_5 inst_cell_108_106 (.BL(BL106),.BLN(BLN106),.WL(WL108));
sram_cell_6t_5 inst_cell_108_107 (.BL(BL107),.BLN(BLN107),.WL(WL108));
sram_cell_6t_5 inst_cell_108_108 (.BL(BL108),.BLN(BLN108),.WL(WL108));
sram_cell_6t_5 inst_cell_108_109 (.BL(BL109),.BLN(BLN109),.WL(WL108));
sram_cell_6t_5 inst_cell_108_110 (.BL(BL110),.BLN(BLN110),.WL(WL108));
sram_cell_6t_5 inst_cell_108_111 (.BL(BL111),.BLN(BLN111),.WL(WL108));
sram_cell_6t_5 inst_cell_108_112 (.BL(BL112),.BLN(BLN112),.WL(WL108));
sram_cell_6t_5 inst_cell_108_113 (.BL(BL113),.BLN(BLN113),.WL(WL108));
sram_cell_6t_5 inst_cell_108_114 (.BL(BL114),.BLN(BLN114),.WL(WL108));
sram_cell_6t_5 inst_cell_108_115 (.BL(BL115),.BLN(BLN115),.WL(WL108));
sram_cell_6t_5 inst_cell_108_116 (.BL(BL116),.BLN(BLN116),.WL(WL108));
sram_cell_6t_5 inst_cell_108_117 (.BL(BL117),.BLN(BLN117),.WL(WL108));
sram_cell_6t_5 inst_cell_108_118 (.BL(BL118),.BLN(BLN118),.WL(WL108));
sram_cell_6t_5 inst_cell_108_119 (.BL(BL119),.BLN(BLN119),.WL(WL108));
sram_cell_6t_5 inst_cell_108_120 (.BL(BL120),.BLN(BLN120),.WL(WL108));
sram_cell_6t_5 inst_cell_108_121 (.BL(BL121),.BLN(BLN121),.WL(WL108));
sram_cell_6t_5 inst_cell_108_122 (.BL(BL122),.BLN(BLN122),.WL(WL108));
sram_cell_6t_5 inst_cell_108_123 (.BL(BL123),.BLN(BLN123),.WL(WL108));
sram_cell_6t_5 inst_cell_108_124 (.BL(BL124),.BLN(BLN124),.WL(WL108));
sram_cell_6t_5 inst_cell_108_125 (.BL(BL125),.BLN(BLN125),.WL(WL108));
sram_cell_6t_5 inst_cell_108_126 (.BL(BL126),.BLN(BLN126),.WL(WL108));
sram_cell_6t_5 inst_cell_108_127 (.BL(BL127),.BLN(BLN127),.WL(WL108));
sram_cell_6t_5 inst_cell_109_0 (.BL(BL0),.BLN(BLN0),.WL(WL109));
sram_cell_6t_5 inst_cell_109_1 (.BL(BL1),.BLN(BLN1),.WL(WL109));
sram_cell_6t_5 inst_cell_109_2 (.BL(BL2),.BLN(BLN2),.WL(WL109));
sram_cell_6t_5 inst_cell_109_3 (.BL(BL3),.BLN(BLN3),.WL(WL109));
sram_cell_6t_5 inst_cell_109_4 (.BL(BL4),.BLN(BLN4),.WL(WL109));
sram_cell_6t_5 inst_cell_109_5 (.BL(BL5),.BLN(BLN5),.WL(WL109));
sram_cell_6t_5 inst_cell_109_6 (.BL(BL6),.BLN(BLN6),.WL(WL109));
sram_cell_6t_5 inst_cell_109_7 (.BL(BL7),.BLN(BLN7),.WL(WL109));
sram_cell_6t_5 inst_cell_109_8 (.BL(BL8),.BLN(BLN8),.WL(WL109));
sram_cell_6t_5 inst_cell_109_9 (.BL(BL9),.BLN(BLN9),.WL(WL109));
sram_cell_6t_5 inst_cell_109_10 (.BL(BL10),.BLN(BLN10),.WL(WL109));
sram_cell_6t_5 inst_cell_109_11 (.BL(BL11),.BLN(BLN11),.WL(WL109));
sram_cell_6t_5 inst_cell_109_12 (.BL(BL12),.BLN(BLN12),.WL(WL109));
sram_cell_6t_5 inst_cell_109_13 (.BL(BL13),.BLN(BLN13),.WL(WL109));
sram_cell_6t_5 inst_cell_109_14 (.BL(BL14),.BLN(BLN14),.WL(WL109));
sram_cell_6t_5 inst_cell_109_15 (.BL(BL15),.BLN(BLN15),.WL(WL109));
sram_cell_6t_5 inst_cell_109_16 (.BL(BL16),.BLN(BLN16),.WL(WL109));
sram_cell_6t_5 inst_cell_109_17 (.BL(BL17),.BLN(BLN17),.WL(WL109));
sram_cell_6t_5 inst_cell_109_18 (.BL(BL18),.BLN(BLN18),.WL(WL109));
sram_cell_6t_5 inst_cell_109_19 (.BL(BL19),.BLN(BLN19),.WL(WL109));
sram_cell_6t_5 inst_cell_109_20 (.BL(BL20),.BLN(BLN20),.WL(WL109));
sram_cell_6t_5 inst_cell_109_21 (.BL(BL21),.BLN(BLN21),.WL(WL109));
sram_cell_6t_5 inst_cell_109_22 (.BL(BL22),.BLN(BLN22),.WL(WL109));
sram_cell_6t_5 inst_cell_109_23 (.BL(BL23),.BLN(BLN23),.WL(WL109));
sram_cell_6t_5 inst_cell_109_24 (.BL(BL24),.BLN(BLN24),.WL(WL109));
sram_cell_6t_5 inst_cell_109_25 (.BL(BL25),.BLN(BLN25),.WL(WL109));
sram_cell_6t_5 inst_cell_109_26 (.BL(BL26),.BLN(BLN26),.WL(WL109));
sram_cell_6t_5 inst_cell_109_27 (.BL(BL27),.BLN(BLN27),.WL(WL109));
sram_cell_6t_5 inst_cell_109_28 (.BL(BL28),.BLN(BLN28),.WL(WL109));
sram_cell_6t_5 inst_cell_109_29 (.BL(BL29),.BLN(BLN29),.WL(WL109));
sram_cell_6t_5 inst_cell_109_30 (.BL(BL30),.BLN(BLN30),.WL(WL109));
sram_cell_6t_5 inst_cell_109_31 (.BL(BL31),.BLN(BLN31),.WL(WL109));
sram_cell_6t_5 inst_cell_109_32 (.BL(BL32),.BLN(BLN32),.WL(WL109));
sram_cell_6t_5 inst_cell_109_33 (.BL(BL33),.BLN(BLN33),.WL(WL109));
sram_cell_6t_5 inst_cell_109_34 (.BL(BL34),.BLN(BLN34),.WL(WL109));
sram_cell_6t_5 inst_cell_109_35 (.BL(BL35),.BLN(BLN35),.WL(WL109));
sram_cell_6t_5 inst_cell_109_36 (.BL(BL36),.BLN(BLN36),.WL(WL109));
sram_cell_6t_5 inst_cell_109_37 (.BL(BL37),.BLN(BLN37),.WL(WL109));
sram_cell_6t_5 inst_cell_109_38 (.BL(BL38),.BLN(BLN38),.WL(WL109));
sram_cell_6t_5 inst_cell_109_39 (.BL(BL39),.BLN(BLN39),.WL(WL109));
sram_cell_6t_5 inst_cell_109_40 (.BL(BL40),.BLN(BLN40),.WL(WL109));
sram_cell_6t_5 inst_cell_109_41 (.BL(BL41),.BLN(BLN41),.WL(WL109));
sram_cell_6t_5 inst_cell_109_42 (.BL(BL42),.BLN(BLN42),.WL(WL109));
sram_cell_6t_5 inst_cell_109_43 (.BL(BL43),.BLN(BLN43),.WL(WL109));
sram_cell_6t_5 inst_cell_109_44 (.BL(BL44),.BLN(BLN44),.WL(WL109));
sram_cell_6t_5 inst_cell_109_45 (.BL(BL45),.BLN(BLN45),.WL(WL109));
sram_cell_6t_5 inst_cell_109_46 (.BL(BL46),.BLN(BLN46),.WL(WL109));
sram_cell_6t_5 inst_cell_109_47 (.BL(BL47),.BLN(BLN47),.WL(WL109));
sram_cell_6t_5 inst_cell_109_48 (.BL(BL48),.BLN(BLN48),.WL(WL109));
sram_cell_6t_5 inst_cell_109_49 (.BL(BL49),.BLN(BLN49),.WL(WL109));
sram_cell_6t_5 inst_cell_109_50 (.BL(BL50),.BLN(BLN50),.WL(WL109));
sram_cell_6t_5 inst_cell_109_51 (.BL(BL51),.BLN(BLN51),.WL(WL109));
sram_cell_6t_5 inst_cell_109_52 (.BL(BL52),.BLN(BLN52),.WL(WL109));
sram_cell_6t_5 inst_cell_109_53 (.BL(BL53),.BLN(BLN53),.WL(WL109));
sram_cell_6t_5 inst_cell_109_54 (.BL(BL54),.BLN(BLN54),.WL(WL109));
sram_cell_6t_5 inst_cell_109_55 (.BL(BL55),.BLN(BLN55),.WL(WL109));
sram_cell_6t_5 inst_cell_109_56 (.BL(BL56),.BLN(BLN56),.WL(WL109));
sram_cell_6t_5 inst_cell_109_57 (.BL(BL57),.BLN(BLN57),.WL(WL109));
sram_cell_6t_5 inst_cell_109_58 (.BL(BL58),.BLN(BLN58),.WL(WL109));
sram_cell_6t_5 inst_cell_109_59 (.BL(BL59),.BLN(BLN59),.WL(WL109));
sram_cell_6t_5 inst_cell_109_60 (.BL(BL60),.BLN(BLN60),.WL(WL109));
sram_cell_6t_5 inst_cell_109_61 (.BL(BL61),.BLN(BLN61),.WL(WL109));
sram_cell_6t_5 inst_cell_109_62 (.BL(BL62),.BLN(BLN62),.WL(WL109));
sram_cell_6t_5 inst_cell_109_63 (.BL(BL63),.BLN(BLN63),.WL(WL109));
sram_cell_6t_5 inst_cell_109_64 (.BL(BL64),.BLN(BLN64),.WL(WL109));
sram_cell_6t_5 inst_cell_109_65 (.BL(BL65),.BLN(BLN65),.WL(WL109));
sram_cell_6t_5 inst_cell_109_66 (.BL(BL66),.BLN(BLN66),.WL(WL109));
sram_cell_6t_5 inst_cell_109_67 (.BL(BL67),.BLN(BLN67),.WL(WL109));
sram_cell_6t_5 inst_cell_109_68 (.BL(BL68),.BLN(BLN68),.WL(WL109));
sram_cell_6t_5 inst_cell_109_69 (.BL(BL69),.BLN(BLN69),.WL(WL109));
sram_cell_6t_5 inst_cell_109_70 (.BL(BL70),.BLN(BLN70),.WL(WL109));
sram_cell_6t_5 inst_cell_109_71 (.BL(BL71),.BLN(BLN71),.WL(WL109));
sram_cell_6t_5 inst_cell_109_72 (.BL(BL72),.BLN(BLN72),.WL(WL109));
sram_cell_6t_5 inst_cell_109_73 (.BL(BL73),.BLN(BLN73),.WL(WL109));
sram_cell_6t_5 inst_cell_109_74 (.BL(BL74),.BLN(BLN74),.WL(WL109));
sram_cell_6t_5 inst_cell_109_75 (.BL(BL75),.BLN(BLN75),.WL(WL109));
sram_cell_6t_5 inst_cell_109_76 (.BL(BL76),.BLN(BLN76),.WL(WL109));
sram_cell_6t_5 inst_cell_109_77 (.BL(BL77),.BLN(BLN77),.WL(WL109));
sram_cell_6t_5 inst_cell_109_78 (.BL(BL78),.BLN(BLN78),.WL(WL109));
sram_cell_6t_5 inst_cell_109_79 (.BL(BL79),.BLN(BLN79),.WL(WL109));
sram_cell_6t_5 inst_cell_109_80 (.BL(BL80),.BLN(BLN80),.WL(WL109));
sram_cell_6t_5 inst_cell_109_81 (.BL(BL81),.BLN(BLN81),.WL(WL109));
sram_cell_6t_5 inst_cell_109_82 (.BL(BL82),.BLN(BLN82),.WL(WL109));
sram_cell_6t_5 inst_cell_109_83 (.BL(BL83),.BLN(BLN83),.WL(WL109));
sram_cell_6t_5 inst_cell_109_84 (.BL(BL84),.BLN(BLN84),.WL(WL109));
sram_cell_6t_5 inst_cell_109_85 (.BL(BL85),.BLN(BLN85),.WL(WL109));
sram_cell_6t_5 inst_cell_109_86 (.BL(BL86),.BLN(BLN86),.WL(WL109));
sram_cell_6t_5 inst_cell_109_87 (.BL(BL87),.BLN(BLN87),.WL(WL109));
sram_cell_6t_5 inst_cell_109_88 (.BL(BL88),.BLN(BLN88),.WL(WL109));
sram_cell_6t_5 inst_cell_109_89 (.BL(BL89),.BLN(BLN89),.WL(WL109));
sram_cell_6t_5 inst_cell_109_90 (.BL(BL90),.BLN(BLN90),.WL(WL109));
sram_cell_6t_5 inst_cell_109_91 (.BL(BL91),.BLN(BLN91),.WL(WL109));
sram_cell_6t_5 inst_cell_109_92 (.BL(BL92),.BLN(BLN92),.WL(WL109));
sram_cell_6t_5 inst_cell_109_93 (.BL(BL93),.BLN(BLN93),.WL(WL109));
sram_cell_6t_5 inst_cell_109_94 (.BL(BL94),.BLN(BLN94),.WL(WL109));
sram_cell_6t_5 inst_cell_109_95 (.BL(BL95),.BLN(BLN95),.WL(WL109));
sram_cell_6t_5 inst_cell_109_96 (.BL(BL96),.BLN(BLN96),.WL(WL109));
sram_cell_6t_5 inst_cell_109_97 (.BL(BL97),.BLN(BLN97),.WL(WL109));
sram_cell_6t_5 inst_cell_109_98 (.BL(BL98),.BLN(BLN98),.WL(WL109));
sram_cell_6t_5 inst_cell_109_99 (.BL(BL99),.BLN(BLN99),.WL(WL109));
sram_cell_6t_5 inst_cell_109_100 (.BL(BL100),.BLN(BLN100),.WL(WL109));
sram_cell_6t_5 inst_cell_109_101 (.BL(BL101),.BLN(BLN101),.WL(WL109));
sram_cell_6t_5 inst_cell_109_102 (.BL(BL102),.BLN(BLN102),.WL(WL109));
sram_cell_6t_5 inst_cell_109_103 (.BL(BL103),.BLN(BLN103),.WL(WL109));
sram_cell_6t_5 inst_cell_109_104 (.BL(BL104),.BLN(BLN104),.WL(WL109));
sram_cell_6t_5 inst_cell_109_105 (.BL(BL105),.BLN(BLN105),.WL(WL109));
sram_cell_6t_5 inst_cell_109_106 (.BL(BL106),.BLN(BLN106),.WL(WL109));
sram_cell_6t_5 inst_cell_109_107 (.BL(BL107),.BLN(BLN107),.WL(WL109));
sram_cell_6t_5 inst_cell_109_108 (.BL(BL108),.BLN(BLN108),.WL(WL109));
sram_cell_6t_5 inst_cell_109_109 (.BL(BL109),.BLN(BLN109),.WL(WL109));
sram_cell_6t_5 inst_cell_109_110 (.BL(BL110),.BLN(BLN110),.WL(WL109));
sram_cell_6t_5 inst_cell_109_111 (.BL(BL111),.BLN(BLN111),.WL(WL109));
sram_cell_6t_5 inst_cell_109_112 (.BL(BL112),.BLN(BLN112),.WL(WL109));
sram_cell_6t_5 inst_cell_109_113 (.BL(BL113),.BLN(BLN113),.WL(WL109));
sram_cell_6t_5 inst_cell_109_114 (.BL(BL114),.BLN(BLN114),.WL(WL109));
sram_cell_6t_5 inst_cell_109_115 (.BL(BL115),.BLN(BLN115),.WL(WL109));
sram_cell_6t_5 inst_cell_109_116 (.BL(BL116),.BLN(BLN116),.WL(WL109));
sram_cell_6t_5 inst_cell_109_117 (.BL(BL117),.BLN(BLN117),.WL(WL109));
sram_cell_6t_5 inst_cell_109_118 (.BL(BL118),.BLN(BLN118),.WL(WL109));
sram_cell_6t_5 inst_cell_109_119 (.BL(BL119),.BLN(BLN119),.WL(WL109));
sram_cell_6t_5 inst_cell_109_120 (.BL(BL120),.BLN(BLN120),.WL(WL109));
sram_cell_6t_5 inst_cell_109_121 (.BL(BL121),.BLN(BLN121),.WL(WL109));
sram_cell_6t_5 inst_cell_109_122 (.BL(BL122),.BLN(BLN122),.WL(WL109));
sram_cell_6t_5 inst_cell_109_123 (.BL(BL123),.BLN(BLN123),.WL(WL109));
sram_cell_6t_5 inst_cell_109_124 (.BL(BL124),.BLN(BLN124),.WL(WL109));
sram_cell_6t_5 inst_cell_109_125 (.BL(BL125),.BLN(BLN125),.WL(WL109));
sram_cell_6t_5 inst_cell_109_126 (.BL(BL126),.BLN(BLN126),.WL(WL109));
sram_cell_6t_5 inst_cell_109_127 (.BL(BL127),.BLN(BLN127),.WL(WL109));
sram_cell_6t_5 inst_cell_110_0 (.BL(BL0),.BLN(BLN0),.WL(WL110));
sram_cell_6t_5 inst_cell_110_1 (.BL(BL1),.BLN(BLN1),.WL(WL110));
sram_cell_6t_5 inst_cell_110_2 (.BL(BL2),.BLN(BLN2),.WL(WL110));
sram_cell_6t_5 inst_cell_110_3 (.BL(BL3),.BLN(BLN3),.WL(WL110));
sram_cell_6t_5 inst_cell_110_4 (.BL(BL4),.BLN(BLN4),.WL(WL110));
sram_cell_6t_5 inst_cell_110_5 (.BL(BL5),.BLN(BLN5),.WL(WL110));
sram_cell_6t_5 inst_cell_110_6 (.BL(BL6),.BLN(BLN6),.WL(WL110));
sram_cell_6t_5 inst_cell_110_7 (.BL(BL7),.BLN(BLN7),.WL(WL110));
sram_cell_6t_5 inst_cell_110_8 (.BL(BL8),.BLN(BLN8),.WL(WL110));
sram_cell_6t_5 inst_cell_110_9 (.BL(BL9),.BLN(BLN9),.WL(WL110));
sram_cell_6t_5 inst_cell_110_10 (.BL(BL10),.BLN(BLN10),.WL(WL110));
sram_cell_6t_5 inst_cell_110_11 (.BL(BL11),.BLN(BLN11),.WL(WL110));
sram_cell_6t_5 inst_cell_110_12 (.BL(BL12),.BLN(BLN12),.WL(WL110));
sram_cell_6t_5 inst_cell_110_13 (.BL(BL13),.BLN(BLN13),.WL(WL110));
sram_cell_6t_5 inst_cell_110_14 (.BL(BL14),.BLN(BLN14),.WL(WL110));
sram_cell_6t_5 inst_cell_110_15 (.BL(BL15),.BLN(BLN15),.WL(WL110));
sram_cell_6t_5 inst_cell_110_16 (.BL(BL16),.BLN(BLN16),.WL(WL110));
sram_cell_6t_5 inst_cell_110_17 (.BL(BL17),.BLN(BLN17),.WL(WL110));
sram_cell_6t_5 inst_cell_110_18 (.BL(BL18),.BLN(BLN18),.WL(WL110));
sram_cell_6t_5 inst_cell_110_19 (.BL(BL19),.BLN(BLN19),.WL(WL110));
sram_cell_6t_5 inst_cell_110_20 (.BL(BL20),.BLN(BLN20),.WL(WL110));
sram_cell_6t_5 inst_cell_110_21 (.BL(BL21),.BLN(BLN21),.WL(WL110));
sram_cell_6t_5 inst_cell_110_22 (.BL(BL22),.BLN(BLN22),.WL(WL110));
sram_cell_6t_5 inst_cell_110_23 (.BL(BL23),.BLN(BLN23),.WL(WL110));
sram_cell_6t_5 inst_cell_110_24 (.BL(BL24),.BLN(BLN24),.WL(WL110));
sram_cell_6t_5 inst_cell_110_25 (.BL(BL25),.BLN(BLN25),.WL(WL110));
sram_cell_6t_5 inst_cell_110_26 (.BL(BL26),.BLN(BLN26),.WL(WL110));
sram_cell_6t_5 inst_cell_110_27 (.BL(BL27),.BLN(BLN27),.WL(WL110));
sram_cell_6t_5 inst_cell_110_28 (.BL(BL28),.BLN(BLN28),.WL(WL110));
sram_cell_6t_5 inst_cell_110_29 (.BL(BL29),.BLN(BLN29),.WL(WL110));
sram_cell_6t_5 inst_cell_110_30 (.BL(BL30),.BLN(BLN30),.WL(WL110));
sram_cell_6t_5 inst_cell_110_31 (.BL(BL31),.BLN(BLN31),.WL(WL110));
sram_cell_6t_5 inst_cell_110_32 (.BL(BL32),.BLN(BLN32),.WL(WL110));
sram_cell_6t_5 inst_cell_110_33 (.BL(BL33),.BLN(BLN33),.WL(WL110));
sram_cell_6t_5 inst_cell_110_34 (.BL(BL34),.BLN(BLN34),.WL(WL110));
sram_cell_6t_5 inst_cell_110_35 (.BL(BL35),.BLN(BLN35),.WL(WL110));
sram_cell_6t_5 inst_cell_110_36 (.BL(BL36),.BLN(BLN36),.WL(WL110));
sram_cell_6t_5 inst_cell_110_37 (.BL(BL37),.BLN(BLN37),.WL(WL110));
sram_cell_6t_5 inst_cell_110_38 (.BL(BL38),.BLN(BLN38),.WL(WL110));
sram_cell_6t_5 inst_cell_110_39 (.BL(BL39),.BLN(BLN39),.WL(WL110));
sram_cell_6t_5 inst_cell_110_40 (.BL(BL40),.BLN(BLN40),.WL(WL110));
sram_cell_6t_5 inst_cell_110_41 (.BL(BL41),.BLN(BLN41),.WL(WL110));
sram_cell_6t_5 inst_cell_110_42 (.BL(BL42),.BLN(BLN42),.WL(WL110));
sram_cell_6t_5 inst_cell_110_43 (.BL(BL43),.BLN(BLN43),.WL(WL110));
sram_cell_6t_5 inst_cell_110_44 (.BL(BL44),.BLN(BLN44),.WL(WL110));
sram_cell_6t_5 inst_cell_110_45 (.BL(BL45),.BLN(BLN45),.WL(WL110));
sram_cell_6t_5 inst_cell_110_46 (.BL(BL46),.BLN(BLN46),.WL(WL110));
sram_cell_6t_5 inst_cell_110_47 (.BL(BL47),.BLN(BLN47),.WL(WL110));
sram_cell_6t_5 inst_cell_110_48 (.BL(BL48),.BLN(BLN48),.WL(WL110));
sram_cell_6t_5 inst_cell_110_49 (.BL(BL49),.BLN(BLN49),.WL(WL110));
sram_cell_6t_5 inst_cell_110_50 (.BL(BL50),.BLN(BLN50),.WL(WL110));
sram_cell_6t_5 inst_cell_110_51 (.BL(BL51),.BLN(BLN51),.WL(WL110));
sram_cell_6t_5 inst_cell_110_52 (.BL(BL52),.BLN(BLN52),.WL(WL110));
sram_cell_6t_5 inst_cell_110_53 (.BL(BL53),.BLN(BLN53),.WL(WL110));
sram_cell_6t_5 inst_cell_110_54 (.BL(BL54),.BLN(BLN54),.WL(WL110));
sram_cell_6t_5 inst_cell_110_55 (.BL(BL55),.BLN(BLN55),.WL(WL110));
sram_cell_6t_5 inst_cell_110_56 (.BL(BL56),.BLN(BLN56),.WL(WL110));
sram_cell_6t_5 inst_cell_110_57 (.BL(BL57),.BLN(BLN57),.WL(WL110));
sram_cell_6t_5 inst_cell_110_58 (.BL(BL58),.BLN(BLN58),.WL(WL110));
sram_cell_6t_5 inst_cell_110_59 (.BL(BL59),.BLN(BLN59),.WL(WL110));
sram_cell_6t_5 inst_cell_110_60 (.BL(BL60),.BLN(BLN60),.WL(WL110));
sram_cell_6t_5 inst_cell_110_61 (.BL(BL61),.BLN(BLN61),.WL(WL110));
sram_cell_6t_5 inst_cell_110_62 (.BL(BL62),.BLN(BLN62),.WL(WL110));
sram_cell_6t_5 inst_cell_110_63 (.BL(BL63),.BLN(BLN63),.WL(WL110));
sram_cell_6t_5 inst_cell_110_64 (.BL(BL64),.BLN(BLN64),.WL(WL110));
sram_cell_6t_5 inst_cell_110_65 (.BL(BL65),.BLN(BLN65),.WL(WL110));
sram_cell_6t_5 inst_cell_110_66 (.BL(BL66),.BLN(BLN66),.WL(WL110));
sram_cell_6t_5 inst_cell_110_67 (.BL(BL67),.BLN(BLN67),.WL(WL110));
sram_cell_6t_5 inst_cell_110_68 (.BL(BL68),.BLN(BLN68),.WL(WL110));
sram_cell_6t_5 inst_cell_110_69 (.BL(BL69),.BLN(BLN69),.WL(WL110));
sram_cell_6t_5 inst_cell_110_70 (.BL(BL70),.BLN(BLN70),.WL(WL110));
sram_cell_6t_5 inst_cell_110_71 (.BL(BL71),.BLN(BLN71),.WL(WL110));
sram_cell_6t_5 inst_cell_110_72 (.BL(BL72),.BLN(BLN72),.WL(WL110));
sram_cell_6t_5 inst_cell_110_73 (.BL(BL73),.BLN(BLN73),.WL(WL110));
sram_cell_6t_5 inst_cell_110_74 (.BL(BL74),.BLN(BLN74),.WL(WL110));
sram_cell_6t_5 inst_cell_110_75 (.BL(BL75),.BLN(BLN75),.WL(WL110));
sram_cell_6t_5 inst_cell_110_76 (.BL(BL76),.BLN(BLN76),.WL(WL110));
sram_cell_6t_5 inst_cell_110_77 (.BL(BL77),.BLN(BLN77),.WL(WL110));
sram_cell_6t_5 inst_cell_110_78 (.BL(BL78),.BLN(BLN78),.WL(WL110));
sram_cell_6t_5 inst_cell_110_79 (.BL(BL79),.BLN(BLN79),.WL(WL110));
sram_cell_6t_5 inst_cell_110_80 (.BL(BL80),.BLN(BLN80),.WL(WL110));
sram_cell_6t_5 inst_cell_110_81 (.BL(BL81),.BLN(BLN81),.WL(WL110));
sram_cell_6t_5 inst_cell_110_82 (.BL(BL82),.BLN(BLN82),.WL(WL110));
sram_cell_6t_5 inst_cell_110_83 (.BL(BL83),.BLN(BLN83),.WL(WL110));
sram_cell_6t_5 inst_cell_110_84 (.BL(BL84),.BLN(BLN84),.WL(WL110));
sram_cell_6t_5 inst_cell_110_85 (.BL(BL85),.BLN(BLN85),.WL(WL110));
sram_cell_6t_5 inst_cell_110_86 (.BL(BL86),.BLN(BLN86),.WL(WL110));
sram_cell_6t_5 inst_cell_110_87 (.BL(BL87),.BLN(BLN87),.WL(WL110));
sram_cell_6t_5 inst_cell_110_88 (.BL(BL88),.BLN(BLN88),.WL(WL110));
sram_cell_6t_5 inst_cell_110_89 (.BL(BL89),.BLN(BLN89),.WL(WL110));
sram_cell_6t_5 inst_cell_110_90 (.BL(BL90),.BLN(BLN90),.WL(WL110));
sram_cell_6t_5 inst_cell_110_91 (.BL(BL91),.BLN(BLN91),.WL(WL110));
sram_cell_6t_5 inst_cell_110_92 (.BL(BL92),.BLN(BLN92),.WL(WL110));
sram_cell_6t_5 inst_cell_110_93 (.BL(BL93),.BLN(BLN93),.WL(WL110));
sram_cell_6t_5 inst_cell_110_94 (.BL(BL94),.BLN(BLN94),.WL(WL110));
sram_cell_6t_5 inst_cell_110_95 (.BL(BL95),.BLN(BLN95),.WL(WL110));
sram_cell_6t_5 inst_cell_110_96 (.BL(BL96),.BLN(BLN96),.WL(WL110));
sram_cell_6t_5 inst_cell_110_97 (.BL(BL97),.BLN(BLN97),.WL(WL110));
sram_cell_6t_5 inst_cell_110_98 (.BL(BL98),.BLN(BLN98),.WL(WL110));
sram_cell_6t_5 inst_cell_110_99 (.BL(BL99),.BLN(BLN99),.WL(WL110));
sram_cell_6t_5 inst_cell_110_100 (.BL(BL100),.BLN(BLN100),.WL(WL110));
sram_cell_6t_5 inst_cell_110_101 (.BL(BL101),.BLN(BLN101),.WL(WL110));
sram_cell_6t_5 inst_cell_110_102 (.BL(BL102),.BLN(BLN102),.WL(WL110));
sram_cell_6t_5 inst_cell_110_103 (.BL(BL103),.BLN(BLN103),.WL(WL110));
sram_cell_6t_5 inst_cell_110_104 (.BL(BL104),.BLN(BLN104),.WL(WL110));
sram_cell_6t_5 inst_cell_110_105 (.BL(BL105),.BLN(BLN105),.WL(WL110));
sram_cell_6t_5 inst_cell_110_106 (.BL(BL106),.BLN(BLN106),.WL(WL110));
sram_cell_6t_5 inst_cell_110_107 (.BL(BL107),.BLN(BLN107),.WL(WL110));
sram_cell_6t_5 inst_cell_110_108 (.BL(BL108),.BLN(BLN108),.WL(WL110));
sram_cell_6t_5 inst_cell_110_109 (.BL(BL109),.BLN(BLN109),.WL(WL110));
sram_cell_6t_5 inst_cell_110_110 (.BL(BL110),.BLN(BLN110),.WL(WL110));
sram_cell_6t_5 inst_cell_110_111 (.BL(BL111),.BLN(BLN111),.WL(WL110));
sram_cell_6t_5 inst_cell_110_112 (.BL(BL112),.BLN(BLN112),.WL(WL110));
sram_cell_6t_5 inst_cell_110_113 (.BL(BL113),.BLN(BLN113),.WL(WL110));
sram_cell_6t_5 inst_cell_110_114 (.BL(BL114),.BLN(BLN114),.WL(WL110));
sram_cell_6t_5 inst_cell_110_115 (.BL(BL115),.BLN(BLN115),.WL(WL110));
sram_cell_6t_5 inst_cell_110_116 (.BL(BL116),.BLN(BLN116),.WL(WL110));
sram_cell_6t_5 inst_cell_110_117 (.BL(BL117),.BLN(BLN117),.WL(WL110));
sram_cell_6t_5 inst_cell_110_118 (.BL(BL118),.BLN(BLN118),.WL(WL110));
sram_cell_6t_5 inst_cell_110_119 (.BL(BL119),.BLN(BLN119),.WL(WL110));
sram_cell_6t_5 inst_cell_110_120 (.BL(BL120),.BLN(BLN120),.WL(WL110));
sram_cell_6t_5 inst_cell_110_121 (.BL(BL121),.BLN(BLN121),.WL(WL110));
sram_cell_6t_5 inst_cell_110_122 (.BL(BL122),.BLN(BLN122),.WL(WL110));
sram_cell_6t_5 inst_cell_110_123 (.BL(BL123),.BLN(BLN123),.WL(WL110));
sram_cell_6t_5 inst_cell_110_124 (.BL(BL124),.BLN(BLN124),.WL(WL110));
sram_cell_6t_5 inst_cell_110_125 (.BL(BL125),.BLN(BLN125),.WL(WL110));
sram_cell_6t_5 inst_cell_110_126 (.BL(BL126),.BLN(BLN126),.WL(WL110));
sram_cell_6t_5 inst_cell_110_127 (.BL(BL127),.BLN(BLN127),.WL(WL110));
sram_cell_6t_5 inst_cell_111_0 (.BL(BL0),.BLN(BLN0),.WL(WL111));
sram_cell_6t_5 inst_cell_111_1 (.BL(BL1),.BLN(BLN1),.WL(WL111));
sram_cell_6t_5 inst_cell_111_2 (.BL(BL2),.BLN(BLN2),.WL(WL111));
sram_cell_6t_5 inst_cell_111_3 (.BL(BL3),.BLN(BLN3),.WL(WL111));
sram_cell_6t_5 inst_cell_111_4 (.BL(BL4),.BLN(BLN4),.WL(WL111));
sram_cell_6t_5 inst_cell_111_5 (.BL(BL5),.BLN(BLN5),.WL(WL111));
sram_cell_6t_5 inst_cell_111_6 (.BL(BL6),.BLN(BLN6),.WL(WL111));
sram_cell_6t_5 inst_cell_111_7 (.BL(BL7),.BLN(BLN7),.WL(WL111));
sram_cell_6t_5 inst_cell_111_8 (.BL(BL8),.BLN(BLN8),.WL(WL111));
sram_cell_6t_5 inst_cell_111_9 (.BL(BL9),.BLN(BLN9),.WL(WL111));
sram_cell_6t_5 inst_cell_111_10 (.BL(BL10),.BLN(BLN10),.WL(WL111));
sram_cell_6t_5 inst_cell_111_11 (.BL(BL11),.BLN(BLN11),.WL(WL111));
sram_cell_6t_5 inst_cell_111_12 (.BL(BL12),.BLN(BLN12),.WL(WL111));
sram_cell_6t_5 inst_cell_111_13 (.BL(BL13),.BLN(BLN13),.WL(WL111));
sram_cell_6t_5 inst_cell_111_14 (.BL(BL14),.BLN(BLN14),.WL(WL111));
sram_cell_6t_5 inst_cell_111_15 (.BL(BL15),.BLN(BLN15),.WL(WL111));
sram_cell_6t_5 inst_cell_111_16 (.BL(BL16),.BLN(BLN16),.WL(WL111));
sram_cell_6t_5 inst_cell_111_17 (.BL(BL17),.BLN(BLN17),.WL(WL111));
sram_cell_6t_5 inst_cell_111_18 (.BL(BL18),.BLN(BLN18),.WL(WL111));
sram_cell_6t_5 inst_cell_111_19 (.BL(BL19),.BLN(BLN19),.WL(WL111));
sram_cell_6t_5 inst_cell_111_20 (.BL(BL20),.BLN(BLN20),.WL(WL111));
sram_cell_6t_5 inst_cell_111_21 (.BL(BL21),.BLN(BLN21),.WL(WL111));
sram_cell_6t_5 inst_cell_111_22 (.BL(BL22),.BLN(BLN22),.WL(WL111));
sram_cell_6t_5 inst_cell_111_23 (.BL(BL23),.BLN(BLN23),.WL(WL111));
sram_cell_6t_5 inst_cell_111_24 (.BL(BL24),.BLN(BLN24),.WL(WL111));
sram_cell_6t_5 inst_cell_111_25 (.BL(BL25),.BLN(BLN25),.WL(WL111));
sram_cell_6t_5 inst_cell_111_26 (.BL(BL26),.BLN(BLN26),.WL(WL111));
sram_cell_6t_5 inst_cell_111_27 (.BL(BL27),.BLN(BLN27),.WL(WL111));
sram_cell_6t_5 inst_cell_111_28 (.BL(BL28),.BLN(BLN28),.WL(WL111));
sram_cell_6t_5 inst_cell_111_29 (.BL(BL29),.BLN(BLN29),.WL(WL111));
sram_cell_6t_5 inst_cell_111_30 (.BL(BL30),.BLN(BLN30),.WL(WL111));
sram_cell_6t_5 inst_cell_111_31 (.BL(BL31),.BLN(BLN31),.WL(WL111));
sram_cell_6t_5 inst_cell_111_32 (.BL(BL32),.BLN(BLN32),.WL(WL111));
sram_cell_6t_5 inst_cell_111_33 (.BL(BL33),.BLN(BLN33),.WL(WL111));
sram_cell_6t_5 inst_cell_111_34 (.BL(BL34),.BLN(BLN34),.WL(WL111));
sram_cell_6t_5 inst_cell_111_35 (.BL(BL35),.BLN(BLN35),.WL(WL111));
sram_cell_6t_5 inst_cell_111_36 (.BL(BL36),.BLN(BLN36),.WL(WL111));
sram_cell_6t_5 inst_cell_111_37 (.BL(BL37),.BLN(BLN37),.WL(WL111));
sram_cell_6t_5 inst_cell_111_38 (.BL(BL38),.BLN(BLN38),.WL(WL111));
sram_cell_6t_5 inst_cell_111_39 (.BL(BL39),.BLN(BLN39),.WL(WL111));
sram_cell_6t_5 inst_cell_111_40 (.BL(BL40),.BLN(BLN40),.WL(WL111));
sram_cell_6t_5 inst_cell_111_41 (.BL(BL41),.BLN(BLN41),.WL(WL111));
sram_cell_6t_5 inst_cell_111_42 (.BL(BL42),.BLN(BLN42),.WL(WL111));
sram_cell_6t_5 inst_cell_111_43 (.BL(BL43),.BLN(BLN43),.WL(WL111));
sram_cell_6t_5 inst_cell_111_44 (.BL(BL44),.BLN(BLN44),.WL(WL111));
sram_cell_6t_5 inst_cell_111_45 (.BL(BL45),.BLN(BLN45),.WL(WL111));
sram_cell_6t_5 inst_cell_111_46 (.BL(BL46),.BLN(BLN46),.WL(WL111));
sram_cell_6t_5 inst_cell_111_47 (.BL(BL47),.BLN(BLN47),.WL(WL111));
sram_cell_6t_5 inst_cell_111_48 (.BL(BL48),.BLN(BLN48),.WL(WL111));
sram_cell_6t_5 inst_cell_111_49 (.BL(BL49),.BLN(BLN49),.WL(WL111));
sram_cell_6t_5 inst_cell_111_50 (.BL(BL50),.BLN(BLN50),.WL(WL111));
sram_cell_6t_5 inst_cell_111_51 (.BL(BL51),.BLN(BLN51),.WL(WL111));
sram_cell_6t_5 inst_cell_111_52 (.BL(BL52),.BLN(BLN52),.WL(WL111));
sram_cell_6t_5 inst_cell_111_53 (.BL(BL53),.BLN(BLN53),.WL(WL111));
sram_cell_6t_5 inst_cell_111_54 (.BL(BL54),.BLN(BLN54),.WL(WL111));
sram_cell_6t_5 inst_cell_111_55 (.BL(BL55),.BLN(BLN55),.WL(WL111));
sram_cell_6t_5 inst_cell_111_56 (.BL(BL56),.BLN(BLN56),.WL(WL111));
sram_cell_6t_5 inst_cell_111_57 (.BL(BL57),.BLN(BLN57),.WL(WL111));
sram_cell_6t_5 inst_cell_111_58 (.BL(BL58),.BLN(BLN58),.WL(WL111));
sram_cell_6t_5 inst_cell_111_59 (.BL(BL59),.BLN(BLN59),.WL(WL111));
sram_cell_6t_5 inst_cell_111_60 (.BL(BL60),.BLN(BLN60),.WL(WL111));
sram_cell_6t_5 inst_cell_111_61 (.BL(BL61),.BLN(BLN61),.WL(WL111));
sram_cell_6t_5 inst_cell_111_62 (.BL(BL62),.BLN(BLN62),.WL(WL111));
sram_cell_6t_5 inst_cell_111_63 (.BL(BL63),.BLN(BLN63),.WL(WL111));
sram_cell_6t_5 inst_cell_111_64 (.BL(BL64),.BLN(BLN64),.WL(WL111));
sram_cell_6t_5 inst_cell_111_65 (.BL(BL65),.BLN(BLN65),.WL(WL111));
sram_cell_6t_5 inst_cell_111_66 (.BL(BL66),.BLN(BLN66),.WL(WL111));
sram_cell_6t_5 inst_cell_111_67 (.BL(BL67),.BLN(BLN67),.WL(WL111));
sram_cell_6t_5 inst_cell_111_68 (.BL(BL68),.BLN(BLN68),.WL(WL111));
sram_cell_6t_5 inst_cell_111_69 (.BL(BL69),.BLN(BLN69),.WL(WL111));
sram_cell_6t_5 inst_cell_111_70 (.BL(BL70),.BLN(BLN70),.WL(WL111));
sram_cell_6t_5 inst_cell_111_71 (.BL(BL71),.BLN(BLN71),.WL(WL111));
sram_cell_6t_5 inst_cell_111_72 (.BL(BL72),.BLN(BLN72),.WL(WL111));
sram_cell_6t_5 inst_cell_111_73 (.BL(BL73),.BLN(BLN73),.WL(WL111));
sram_cell_6t_5 inst_cell_111_74 (.BL(BL74),.BLN(BLN74),.WL(WL111));
sram_cell_6t_5 inst_cell_111_75 (.BL(BL75),.BLN(BLN75),.WL(WL111));
sram_cell_6t_5 inst_cell_111_76 (.BL(BL76),.BLN(BLN76),.WL(WL111));
sram_cell_6t_5 inst_cell_111_77 (.BL(BL77),.BLN(BLN77),.WL(WL111));
sram_cell_6t_5 inst_cell_111_78 (.BL(BL78),.BLN(BLN78),.WL(WL111));
sram_cell_6t_5 inst_cell_111_79 (.BL(BL79),.BLN(BLN79),.WL(WL111));
sram_cell_6t_5 inst_cell_111_80 (.BL(BL80),.BLN(BLN80),.WL(WL111));
sram_cell_6t_5 inst_cell_111_81 (.BL(BL81),.BLN(BLN81),.WL(WL111));
sram_cell_6t_5 inst_cell_111_82 (.BL(BL82),.BLN(BLN82),.WL(WL111));
sram_cell_6t_5 inst_cell_111_83 (.BL(BL83),.BLN(BLN83),.WL(WL111));
sram_cell_6t_5 inst_cell_111_84 (.BL(BL84),.BLN(BLN84),.WL(WL111));
sram_cell_6t_5 inst_cell_111_85 (.BL(BL85),.BLN(BLN85),.WL(WL111));
sram_cell_6t_5 inst_cell_111_86 (.BL(BL86),.BLN(BLN86),.WL(WL111));
sram_cell_6t_5 inst_cell_111_87 (.BL(BL87),.BLN(BLN87),.WL(WL111));
sram_cell_6t_5 inst_cell_111_88 (.BL(BL88),.BLN(BLN88),.WL(WL111));
sram_cell_6t_5 inst_cell_111_89 (.BL(BL89),.BLN(BLN89),.WL(WL111));
sram_cell_6t_5 inst_cell_111_90 (.BL(BL90),.BLN(BLN90),.WL(WL111));
sram_cell_6t_5 inst_cell_111_91 (.BL(BL91),.BLN(BLN91),.WL(WL111));
sram_cell_6t_5 inst_cell_111_92 (.BL(BL92),.BLN(BLN92),.WL(WL111));
sram_cell_6t_5 inst_cell_111_93 (.BL(BL93),.BLN(BLN93),.WL(WL111));
sram_cell_6t_5 inst_cell_111_94 (.BL(BL94),.BLN(BLN94),.WL(WL111));
sram_cell_6t_5 inst_cell_111_95 (.BL(BL95),.BLN(BLN95),.WL(WL111));
sram_cell_6t_5 inst_cell_111_96 (.BL(BL96),.BLN(BLN96),.WL(WL111));
sram_cell_6t_5 inst_cell_111_97 (.BL(BL97),.BLN(BLN97),.WL(WL111));
sram_cell_6t_5 inst_cell_111_98 (.BL(BL98),.BLN(BLN98),.WL(WL111));
sram_cell_6t_5 inst_cell_111_99 (.BL(BL99),.BLN(BLN99),.WL(WL111));
sram_cell_6t_5 inst_cell_111_100 (.BL(BL100),.BLN(BLN100),.WL(WL111));
sram_cell_6t_5 inst_cell_111_101 (.BL(BL101),.BLN(BLN101),.WL(WL111));
sram_cell_6t_5 inst_cell_111_102 (.BL(BL102),.BLN(BLN102),.WL(WL111));
sram_cell_6t_5 inst_cell_111_103 (.BL(BL103),.BLN(BLN103),.WL(WL111));
sram_cell_6t_5 inst_cell_111_104 (.BL(BL104),.BLN(BLN104),.WL(WL111));
sram_cell_6t_5 inst_cell_111_105 (.BL(BL105),.BLN(BLN105),.WL(WL111));
sram_cell_6t_5 inst_cell_111_106 (.BL(BL106),.BLN(BLN106),.WL(WL111));
sram_cell_6t_5 inst_cell_111_107 (.BL(BL107),.BLN(BLN107),.WL(WL111));
sram_cell_6t_5 inst_cell_111_108 (.BL(BL108),.BLN(BLN108),.WL(WL111));
sram_cell_6t_5 inst_cell_111_109 (.BL(BL109),.BLN(BLN109),.WL(WL111));
sram_cell_6t_5 inst_cell_111_110 (.BL(BL110),.BLN(BLN110),.WL(WL111));
sram_cell_6t_5 inst_cell_111_111 (.BL(BL111),.BLN(BLN111),.WL(WL111));
sram_cell_6t_5 inst_cell_111_112 (.BL(BL112),.BLN(BLN112),.WL(WL111));
sram_cell_6t_5 inst_cell_111_113 (.BL(BL113),.BLN(BLN113),.WL(WL111));
sram_cell_6t_5 inst_cell_111_114 (.BL(BL114),.BLN(BLN114),.WL(WL111));
sram_cell_6t_5 inst_cell_111_115 (.BL(BL115),.BLN(BLN115),.WL(WL111));
sram_cell_6t_5 inst_cell_111_116 (.BL(BL116),.BLN(BLN116),.WL(WL111));
sram_cell_6t_5 inst_cell_111_117 (.BL(BL117),.BLN(BLN117),.WL(WL111));
sram_cell_6t_5 inst_cell_111_118 (.BL(BL118),.BLN(BLN118),.WL(WL111));
sram_cell_6t_5 inst_cell_111_119 (.BL(BL119),.BLN(BLN119),.WL(WL111));
sram_cell_6t_5 inst_cell_111_120 (.BL(BL120),.BLN(BLN120),.WL(WL111));
sram_cell_6t_5 inst_cell_111_121 (.BL(BL121),.BLN(BLN121),.WL(WL111));
sram_cell_6t_5 inst_cell_111_122 (.BL(BL122),.BLN(BLN122),.WL(WL111));
sram_cell_6t_5 inst_cell_111_123 (.BL(BL123),.BLN(BLN123),.WL(WL111));
sram_cell_6t_5 inst_cell_111_124 (.BL(BL124),.BLN(BLN124),.WL(WL111));
sram_cell_6t_5 inst_cell_111_125 (.BL(BL125),.BLN(BLN125),.WL(WL111));
sram_cell_6t_5 inst_cell_111_126 (.BL(BL126),.BLN(BLN126),.WL(WL111));
sram_cell_6t_5 inst_cell_111_127 (.BL(BL127),.BLN(BLN127),.WL(WL111));
sram_cell_6t_5 inst_cell_112_0 (.BL(BL0),.BLN(BLN0),.WL(WL112));
sram_cell_6t_5 inst_cell_112_1 (.BL(BL1),.BLN(BLN1),.WL(WL112));
sram_cell_6t_5 inst_cell_112_2 (.BL(BL2),.BLN(BLN2),.WL(WL112));
sram_cell_6t_5 inst_cell_112_3 (.BL(BL3),.BLN(BLN3),.WL(WL112));
sram_cell_6t_5 inst_cell_112_4 (.BL(BL4),.BLN(BLN4),.WL(WL112));
sram_cell_6t_5 inst_cell_112_5 (.BL(BL5),.BLN(BLN5),.WL(WL112));
sram_cell_6t_5 inst_cell_112_6 (.BL(BL6),.BLN(BLN6),.WL(WL112));
sram_cell_6t_5 inst_cell_112_7 (.BL(BL7),.BLN(BLN7),.WL(WL112));
sram_cell_6t_5 inst_cell_112_8 (.BL(BL8),.BLN(BLN8),.WL(WL112));
sram_cell_6t_5 inst_cell_112_9 (.BL(BL9),.BLN(BLN9),.WL(WL112));
sram_cell_6t_5 inst_cell_112_10 (.BL(BL10),.BLN(BLN10),.WL(WL112));
sram_cell_6t_5 inst_cell_112_11 (.BL(BL11),.BLN(BLN11),.WL(WL112));
sram_cell_6t_5 inst_cell_112_12 (.BL(BL12),.BLN(BLN12),.WL(WL112));
sram_cell_6t_5 inst_cell_112_13 (.BL(BL13),.BLN(BLN13),.WL(WL112));
sram_cell_6t_5 inst_cell_112_14 (.BL(BL14),.BLN(BLN14),.WL(WL112));
sram_cell_6t_5 inst_cell_112_15 (.BL(BL15),.BLN(BLN15),.WL(WL112));
sram_cell_6t_5 inst_cell_112_16 (.BL(BL16),.BLN(BLN16),.WL(WL112));
sram_cell_6t_5 inst_cell_112_17 (.BL(BL17),.BLN(BLN17),.WL(WL112));
sram_cell_6t_5 inst_cell_112_18 (.BL(BL18),.BLN(BLN18),.WL(WL112));
sram_cell_6t_5 inst_cell_112_19 (.BL(BL19),.BLN(BLN19),.WL(WL112));
sram_cell_6t_5 inst_cell_112_20 (.BL(BL20),.BLN(BLN20),.WL(WL112));
sram_cell_6t_5 inst_cell_112_21 (.BL(BL21),.BLN(BLN21),.WL(WL112));
sram_cell_6t_5 inst_cell_112_22 (.BL(BL22),.BLN(BLN22),.WL(WL112));
sram_cell_6t_5 inst_cell_112_23 (.BL(BL23),.BLN(BLN23),.WL(WL112));
sram_cell_6t_5 inst_cell_112_24 (.BL(BL24),.BLN(BLN24),.WL(WL112));
sram_cell_6t_5 inst_cell_112_25 (.BL(BL25),.BLN(BLN25),.WL(WL112));
sram_cell_6t_5 inst_cell_112_26 (.BL(BL26),.BLN(BLN26),.WL(WL112));
sram_cell_6t_5 inst_cell_112_27 (.BL(BL27),.BLN(BLN27),.WL(WL112));
sram_cell_6t_5 inst_cell_112_28 (.BL(BL28),.BLN(BLN28),.WL(WL112));
sram_cell_6t_5 inst_cell_112_29 (.BL(BL29),.BLN(BLN29),.WL(WL112));
sram_cell_6t_5 inst_cell_112_30 (.BL(BL30),.BLN(BLN30),.WL(WL112));
sram_cell_6t_5 inst_cell_112_31 (.BL(BL31),.BLN(BLN31),.WL(WL112));
sram_cell_6t_5 inst_cell_112_32 (.BL(BL32),.BLN(BLN32),.WL(WL112));
sram_cell_6t_5 inst_cell_112_33 (.BL(BL33),.BLN(BLN33),.WL(WL112));
sram_cell_6t_5 inst_cell_112_34 (.BL(BL34),.BLN(BLN34),.WL(WL112));
sram_cell_6t_5 inst_cell_112_35 (.BL(BL35),.BLN(BLN35),.WL(WL112));
sram_cell_6t_5 inst_cell_112_36 (.BL(BL36),.BLN(BLN36),.WL(WL112));
sram_cell_6t_5 inst_cell_112_37 (.BL(BL37),.BLN(BLN37),.WL(WL112));
sram_cell_6t_5 inst_cell_112_38 (.BL(BL38),.BLN(BLN38),.WL(WL112));
sram_cell_6t_5 inst_cell_112_39 (.BL(BL39),.BLN(BLN39),.WL(WL112));
sram_cell_6t_5 inst_cell_112_40 (.BL(BL40),.BLN(BLN40),.WL(WL112));
sram_cell_6t_5 inst_cell_112_41 (.BL(BL41),.BLN(BLN41),.WL(WL112));
sram_cell_6t_5 inst_cell_112_42 (.BL(BL42),.BLN(BLN42),.WL(WL112));
sram_cell_6t_5 inst_cell_112_43 (.BL(BL43),.BLN(BLN43),.WL(WL112));
sram_cell_6t_5 inst_cell_112_44 (.BL(BL44),.BLN(BLN44),.WL(WL112));
sram_cell_6t_5 inst_cell_112_45 (.BL(BL45),.BLN(BLN45),.WL(WL112));
sram_cell_6t_5 inst_cell_112_46 (.BL(BL46),.BLN(BLN46),.WL(WL112));
sram_cell_6t_5 inst_cell_112_47 (.BL(BL47),.BLN(BLN47),.WL(WL112));
sram_cell_6t_5 inst_cell_112_48 (.BL(BL48),.BLN(BLN48),.WL(WL112));
sram_cell_6t_5 inst_cell_112_49 (.BL(BL49),.BLN(BLN49),.WL(WL112));
sram_cell_6t_5 inst_cell_112_50 (.BL(BL50),.BLN(BLN50),.WL(WL112));
sram_cell_6t_5 inst_cell_112_51 (.BL(BL51),.BLN(BLN51),.WL(WL112));
sram_cell_6t_5 inst_cell_112_52 (.BL(BL52),.BLN(BLN52),.WL(WL112));
sram_cell_6t_5 inst_cell_112_53 (.BL(BL53),.BLN(BLN53),.WL(WL112));
sram_cell_6t_5 inst_cell_112_54 (.BL(BL54),.BLN(BLN54),.WL(WL112));
sram_cell_6t_5 inst_cell_112_55 (.BL(BL55),.BLN(BLN55),.WL(WL112));
sram_cell_6t_5 inst_cell_112_56 (.BL(BL56),.BLN(BLN56),.WL(WL112));
sram_cell_6t_5 inst_cell_112_57 (.BL(BL57),.BLN(BLN57),.WL(WL112));
sram_cell_6t_5 inst_cell_112_58 (.BL(BL58),.BLN(BLN58),.WL(WL112));
sram_cell_6t_5 inst_cell_112_59 (.BL(BL59),.BLN(BLN59),.WL(WL112));
sram_cell_6t_5 inst_cell_112_60 (.BL(BL60),.BLN(BLN60),.WL(WL112));
sram_cell_6t_5 inst_cell_112_61 (.BL(BL61),.BLN(BLN61),.WL(WL112));
sram_cell_6t_5 inst_cell_112_62 (.BL(BL62),.BLN(BLN62),.WL(WL112));
sram_cell_6t_5 inst_cell_112_63 (.BL(BL63),.BLN(BLN63),.WL(WL112));
sram_cell_6t_5 inst_cell_112_64 (.BL(BL64),.BLN(BLN64),.WL(WL112));
sram_cell_6t_5 inst_cell_112_65 (.BL(BL65),.BLN(BLN65),.WL(WL112));
sram_cell_6t_5 inst_cell_112_66 (.BL(BL66),.BLN(BLN66),.WL(WL112));
sram_cell_6t_5 inst_cell_112_67 (.BL(BL67),.BLN(BLN67),.WL(WL112));
sram_cell_6t_5 inst_cell_112_68 (.BL(BL68),.BLN(BLN68),.WL(WL112));
sram_cell_6t_5 inst_cell_112_69 (.BL(BL69),.BLN(BLN69),.WL(WL112));
sram_cell_6t_5 inst_cell_112_70 (.BL(BL70),.BLN(BLN70),.WL(WL112));
sram_cell_6t_5 inst_cell_112_71 (.BL(BL71),.BLN(BLN71),.WL(WL112));
sram_cell_6t_5 inst_cell_112_72 (.BL(BL72),.BLN(BLN72),.WL(WL112));
sram_cell_6t_5 inst_cell_112_73 (.BL(BL73),.BLN(BLN73),.WL(WL112));
sram_cell_6t_5 inst_cell_112_74 (.BL(BL74),.BLN(BLN74),.WL(WL112));
sram_cell_6t_5 inst_cell_112_75 (.BL(BL75),.BLN(BLN75),.WL(WL112));
sram_cell_6t_5 inst_cell_112_76 (.BL(BL76),.BLN(BLN76),.WL(WL112));
sram_cell_6t_5 inst_cell_112_77 (.BL(BL77),.BLN(BLN77),.WL(WL112));
sram_cell_6t_5 inst_cell_112_78 (.BL(BL78),.BLN(BLN78),.WL(WL112));
sram_cell_6t_5 inst_cell_112_79 (.BL(BL79),.BLN(BLN79),.WL(WL112));
sram_cell_6t_5 inst_cell_112_80 (.BL(BL80),.BLN(BLN80),.WL(WL112));
sram_cell_6t_5 inst_cell_112_81 (.BL(BL81),.BLN(BLN81),.WL(WL112));
sram_cell_6t_5 inst_cell_112_82 (.BL(BL82),.BLN(BLN82),.WL(WL112));
sram_cell_6t_5 inst_cell_112_83 (.BL(BL83),.BLN(BLN83),.WL(WL112));
sram_cell_6t_5 inst_cell_112_84 (.BL(BL84),.BLN(BLN84),.WL(WL112));
sram_cell_6t_5 inst_cell_112_85 (.BL(BL85),.BLN(BLN85),.WL(WL112));
sram_cell_6t_5 inst_cell_112_86 (.BL(BL86),.BLN(BLN86),.WL(WL112));
sram_cell_6t_5 inst_cell_112_87 (.BL(BL87),.BLN(BLN87),.WL(WL112));
sram_cell_6t_5 inst_cell_112_88 (.BL(BL88),.BLN(BLN88),.WL(WL112));
sram_cell_6t_5 inst_cell_112_89 (.BL(BL89),.BLN(BLN89),.WL(WL112));
sram_cell_6t_5 inst_cell_112_90 (.BL(BL90),.BLN(BLN90),.WL(WL112));
sram_cell_6t_5 inst_cell_112_91 (.BL(BL91),.BLN(BLN91),.WL(WL112));
sram_cell_6t_5 inst_cell_112_92 (.BL(BL92),.BLN(BLN92),.WL(WL112));
sram_cell_6t_5 inst_cell_112_93 (.BL(BL93),.BLN(BLN93),.WL(WL112));
sram_cell_6t_5 inst_cell_112_94 (.BL(BL94),.BLN(BLN94),.WL(WL112));
sram_cell_6t_5 inst_cell_112_95 (.BL(BL95),.BLN(BLN95),.WL(WL112));
sram_cell_6t_5 inst_cell_112_96 (.BL(BL96),.BLN(BLN96),.WL(WL112));
sram_cell_6t_5 inst_cell_112_97 (.BL(BL97),.BLN(BLN97),.WL(WL112));
sram_cell_6t_5 inst_cell_112_98 (.BL(BL98),.BLN(BLN98),.WL(WL112));
sram_cell_6t_5 inst_cell_112_99 (.BL(BL99),.BLN(BLN99),.WL(WL112));
sram_cell_6t_5 inst_cell_112_100 (.BL(BL100),.BLN(BLN100),.WL(WL112));
sram_cell_6t_5 inst_cell_112_101 (.BL(BL101),.BLN(BLN101),.WL(WL112));
sram_cell_6t_5 inst_cell_112_102 (.BL(BL102),.BLN(BLN102),.WL(WL112));
sram_cell_6t_5 inst_cell_112_103 (.BL(BL103),.BLN(BLN103),.WL(WL112));
sram_cell_6t_5 inst_cell_112_104 (.BL(BL104),.BLN(BLN104),.WL(WL112));
sram_cell_6t_5 inst_cell_112_105 (.BL(BL105),.BLN(BLN105),.WL(WL112));
sram_cell_6t_5 inst_cell_112_106 (.BL(BL106),.BLN(BLN106),.WL(WL112));
sram_cell_6t_5 inst_cell_112_107 (.BL(BL107),.BLN(BLN107),.WL(WL112));
sram_cell_6t_5 inst_cell_112_108 (.BL(BL108),.BLN(BLN108),.WL(WL112));
sram_cell_6t_5 inst_cell_112_109 (.BL(BL109),.BLN(BLN109),.WL(WL112));
sram_cell_6t_5 inst_cell_112_110 (.BL(BL110),.BLN(BLN110),.WL(WL112));
sram_cell_6t_5 inst_cell_112_111 (.BL(BL111),.BLN(BLN111),.WL(WL112));
sram_cell_6t_5 inst_cell_112_112 (.BL(BL112),.BLN(BLN112),.WL(WL112));
sram_cell_6t_5 inst_cell_112_113 (.BL(BL113),.BLN(BLN113),.WL(WL112));
sram_cell_6t_5 inst_cell_112_114 (.BL(BL114),.BLN(BLN114),.WL(WL112));
sram_cell_6t_5 inst_cell_112_115 (.BL(BL115),.BLN(BLN115),.WL(WL112));
sram_cell_6t_5 inst_cell_112_116 (.BL(BL116),.BLN(BLN116),.WL(WL112));
sram_cell_6t_5 inst_cell_112_117 (.BL(BL117),.BLN(BLN117),.WL(WL112));
sram_cell_6t_5 inst_cell_112_118 (.BL(BL118),.BLN(BLN118),.WL(WL112));
sram_cell_6t_5 inst_cell_112_119 (.BL(BL119),.BLN(BLN119),.WL(WL112));
sram_cell_6t_5 inst_cell_112_120 (.BL(BL120),.BLN(BLN120),.WL(WL112));
sram_cell_6t_5 inst_cell_112_121 (.BL(BL121),.BLN(BLN121),.WL(WL112));
sram_cell_6t_5 inst_cell_112_122 (.BL(BL122),.BLN(BLN122),.WL(WL112));
sram_cell_6t_5 inst_cell_112_123 (.BL(BL123),.BLN(BLN123),.WL(WL112));
sram_cell_6t_5 inst_cell_112_124 (.BL(BL124),.BLN(BLN124),.WL(WL112));
sram_cell_6t_5 inst_cell_112_125 (.BL(BL125),.BLN(BLN125),.WL(WL112));
sram_cell_6t_5 inst_cell_112_126 (.BL(BL126),.BLN(BLN126),.WL(WL112));
sram_cell_6t_5 inst_cell_112_127 (.BL(BL127),.BLN(BLN127),.WL(WL112));
sram_cell_6t_5 inst_cell_113_0 (.BL(BL0),.BLN(BLN0),.WL(WL113));
sram_cell_6t_5 inst_cell_113_1 (.BL(BL1),.BLN(BLN1),.WL(WL113));
sram_cell_6t_5 inst_cell_113_2 (.BL(BL2),.BLN(BLN2),.WL(WL113));
sram_cell_6t_5 inst_cell_113_3 (.BL(BL3),.BLN(BLN3),.WL(WL113));
sram_cell_6t_5 inst_cell_113_4 (.BL(BL4),.BLN(BLN4),.WL(WL113));
sram_cell_6t_5 inst_cell_113_5 (.BL(BL5),.BLN(BLN5),.WL(WL113));
sram_cell_6t_5 inst_cell_113_6 (.BL(BL6),.BLN(BLN6),.WL(WL113));
sram_cell_6t_5 inst_cell_113_7 (.BL(BL7),.BLN(BLN7),.WL(WL113));
sram_cell_6t_5 inst_cell_113_8 (.BL(BL8),.BLN(BLN8),.WL(WL113));
sram_cell_6t_5 inst_cell_113_9 (.BL(BL9),.BLN(BLN9),.WL(WL113));
sram_cell_6t_5 inst_cell_113_10 (.BL(BL10),.BLN(BLN10),.WL(WL113));
sram_cell_6t_5 inst_cell_113_11 (.BL(BL11),.BLN(BLN11),.WL(WL113));
sram_cell_6t_5 inst_cell_113_12 (.BL(BL12),.BLN(BLN12),.WL(WL113));
sram_cell_6t_5 inst_cell_113_13 (.BL(BL13),.BLN(BLN13),.WL(WL113));
sram_cell_6t_5 inst_cell_113_14 (.BL(BL14),.BLN(BLN14),.WL(WL113));
sram_cell_6t_5 inst_cell_113_15 (.BL(BL15),.BLN(BLN15),.WL(WL113));
sram_cell_6t_5 inst_cell_113_16 (.BL(BL16),.BLN(BLN16),.WL(WL113));
sram_cell_6t_5 inst_cell_113_17 (.BL(BL17),.BLN(BLN17),.WL(WL113));
sram_cell_6t_5 inst_cell_113_18 (.BL(BL18),.BLN(BLN18),.WL(WL113));
sram_cell_6t_5 inst_cell_113_19 (.BL(BL19),.BLN(BLN19),.WL(WL113));
sram_cell_6t_5 inst_cell_113_20 (.BL(BL20),.BLN(BLN20),.WL(WL113));
sram_cell_6t_5 inst_cell_113_21 (.BL(BL21),.BLN(BLN21),.WL(WL113));
sram_cell_6t_5 inst_cell_113_22 (.BL(BL22),.BLN(BLN22),.WL(WL113));
sram_cell_6t_5 inst_cell_113_23 (.BL(BL23),.BLN(BLN23),.WL(WL113));
sram_cell_6t_5 inst_cell_113_24 (.BL(BL24),.BLN(BLN24),.WL(WL113));
sram_cell_6t_5 inst_cell_113_25 (.BL(BL25),.BLN(BLN25),.WL(WL113));
sram_cell_6t_5 inst_cell_113_26 (.BL(BL26),.BLN(BLN26),.WL(WL113));
sram_cell_6t_5 inst_cell_113_27 (.BL(BL27),.BLN(BLN27),.WL(WL113));
sram_cell_6t_5 inst_cell_113_28 (.BL(BL28),.BLN(BLN28),.WL(WL113));
sram_cell_6t_5 inst_cell_113_29 (.BL(BL29),.BLN(BLN29),.WL(WL113));
sram_cell_6t_5 inst_cell_113_30 (.BL(BL30),.BLN(BLN30),.WL(WL113));
sram_cell_6t_5 inst_cell_113_31 (.BL(BL31),.BLN(BLN31),.WL(WL113));
sram_cell_6t_5 inst_cell_113_32 (.BL(BL32),.BLN(BLN32),.WL(WL113));
sram_cell_6t_5 inst_cell_113_33 (.BL(BL33),.BLN(BLN33),.WL(WL113));
sram_cell_6t_5 inst_cell_113_34 (.BL(BL34),.BLN(BLN34),.WL(WL113));
sram_cell_6t_5 inst_cell_113_35 (.BL(BL35),.BLN(BLN35),.WL(WL113));
sram_cell_6t_5 inst_cell_113_36 (.BL(BL36),.BLN(BLN36),.WL(WL113));
sram_cell_6t_5 inst_cell_113_37 (.BL(BL37),.BLN(BLN37),.WL(WL113));
sram_cell_6t_5 inst_cell_113_38 (.BL(BL38),.BLN(BLN38),.WL(WL113));
sram_cell_6t_5 inst_cell_113_39 (.BL(BL39),.BLN(BLN39),.WL(WL113));
sram_cell_6t_5 inst_cell_113_40 (.BL(BL40),.BLN(BLN40),.WL(WL113));
sram_cell_6t_5 inst_cell_113_41 (.BL(BL41),.BLN(BLN41),.WL(WL113));
sram_cell_6t_5 inst_cell_113_42 (.BL(BL42),.BLN(BLN42),.WL(WL113));
sram_cell_6t_5 inst_cell_113_43 (.BL(BL43),.BLN(BLN43),.WL(WL113));
sram_cell_6t_5 inst_cell_113_44 (.BL(BL44),.BLN(BLN44),.WL(WL113));
sram_cell_6t_5 inst_cell_113_45 (.BL(BL45),.BLN(BLN45),.WL(WL113));
sram_cell_6t_5 inst_cell_113_46 (.BL(BL46),.BLN(BLN46),.WL(WL113));
sram_cell_6t_5 inst_cell_113_47 (.BL(BL47),.BLN(BLN47),.WL(WL113));
sram_cell_6t_5 inst_cell_113_48 (.BL(BL48),.BLN(BLN48),.WL(WL113));
sram_cell_6t_5 inst_cell_113_49 (.BL(BL49),.BLN(BLN49),.WL(WL113));
sram_cell_6t_5 inst_cell_113_50 (.BL(BL50),.BLN(BLN50),.WL(WL113));
sram_cell_6t_5 inst_cell_113_51 (.BL(BL51),.BLN(BLN51),.WL(WL113));
sram_cell_6t_5 inst_cell_113_52 (.BL(BL52),.BLN(BLN52),.WL(WL113));
sram_cell_6t_5 inst_cell_113_53 (.BL(BL53),.BLN(BLN53),.WL(WL113));
sram_cell_6t_5 inst_cell_113_54 (.BL(BL54),.BLN(BLN54),.WL(WL113));
sram_cell_6t_5 inst_cell_113_55 (.BL(BL55),.BLN(BLN55),.WL(WL113));
sram_cell_6t_5 inst_cell_113_56 (.BL(BL56),.BLN(BLN56),.WL(WL113));
sram_cell_6t_5 inst_cell_113_57 (.BL(BL57),.BLN(BLN57),.WL(WL113));
sram_cell_6t_5 inst_cell_113_58 (.BL(BL58),.BLN(BLN58),.WL(WL113));
sram_cell_6t_5 inst_cell_113_59 (.BL(BL59),.BLN(BLN59),.WL(WL113));
sram_cell_6t_5 inst_cell_113_60 (.BL(BL60),.BLN(BLN60),.WL(WL113));
sram_cell_6t_5 inst_cell_113_61 (.BL(BL61),.BLN(BLN61),.WL(WL113));
sram_cell_6t_5 inst_cell_113_62 (.BL(BL62),.BLN(BLN62),.WL(WL113));
sram_cell_6t_5 inst_cell_113_63 (.BL(BL63),.BLN(BLN63),.WL(WL113));
sram_cell_6t_5 inst_cell_113_64 (.BL(BL64),.BLN(BLN64),.WL(WL113));
sram_cell_6t_5 inst_cell_113_65 (.BL(BL65),.BLN(BLN65),.WL(WL113));
sram_cell_6t_5 inst_cell_113_66 (.BL(BL66),.BLN(BLN66),.WL(WL113));
sram_cell_6t_5 inst_cell_113_67 (.BL(BL67),.BLN(BLN67),.WL(WL113));
sram_cell_6t_5 inst_cell_113_68 (.BL(BL68),.BLN(BLN68),.WL(WL113));
sram_cell_6t_5 inst_cell_113_69 (.BL(BL69),.BLN(BLN69),.WL(WL113));
sram_cell_6t_5 inst_cell_113_70 (.BL(BL70),.BLN(BLN70),.WL(WL113));
sram_cell_6t_5 inst_cell_113_71 (.BL(BL71),.BLN(BLN71),.WL(WL113));
sram_cell_6t_5 inst_cell_113_72 (.BL(BL72),.BLN(BLN72),.WL(WL113));
sram_cell_6t_5 inst_cell_113_73 (.BL(BL73),.BLN(BLN73),.WL(WL113));
sram_cell_6t_5 inst_cell_113_74 (.BL(BL74),.BLN(BLN74),.WL(WL113));
sram_cell_6t_5 inst_cell_113_75 (.BL(BL75),.BLN(BLN75),.WL(WL113));
sram_cell_6t_5 inst_cell_113_76 (.BL(BL76),.BLN(BLN76),.WL(WL113));
sram_cell_6t_5 inst_cell_113_77 (.BL(BL77),.BLN(BLN77),.WL(WL113));
sram_cell_6t_5 inst_cell_113_78 (.BL(BL78),.BLN(BLN78),.WL(WL113));
sram_cell_6t_5 inst_cell_113_79 (.BL(BL79),.BLN(BLN79),.WL(WL113));
sram_cell_6t_5 inst_cell_113_80 (.BL(BL80),.BLN(BLN80),.WL(WL113));
sram_cell_6t_5 inst_cell_113_81 (.BL(BL81),.BLN(BLN81),.WL(WL113));
sram_cell_6t_5 inst_cell_113_82 (.BL(BL82),.BLN(BLN82),.WL(WL113));
sram_cell_6t_5 inst_cell_113_83 (.BL(BL83),.BLN(BLN83),.WL(WL113));
sram_cell_6t_5 inst_cell_113_84 (.BL(BL84),.BLN(BLN84),.WL(WL113));
sram_cell_6t_5 inst_cell_113_85 (.BL(BL85),.BLN(BLN85),.WL(WL113));
sram_cell_6t_5 inst_cell_113_86 (.BL(BL86),.BLN(BLN86),.WL(WL113));
sram_cell_6t_5 inst_cell_113_87 (.BL(BL87),.BLN(BLN87),.WL(WL113));
sram_cell_6t_5 inst_cell_113_88 (.BL(BL88),.BLN(BLN88),.WL(WL113));
sram_cell_6t_5 inst_cell_113_89 (.BL(BL89),.BLN(BLN89),.WL(WL113));
sram_cell_6t_5 inst_cell_113_90 (.BL(BL90),.BLN(BLN90),.WL(WL113));
sram_cell_6t_5 inst_cell_113_91 (.BL(BL91),.BLN(BLN91),.WL(WL113));
sram_cell_6t_5 inst_cell_113_92 (.BL(BL92),.BLN(BLN92),.WL(WL113));
sram_cell_6t_5 inst_cell_113_93 (.BL(BL93),.BLN(BLN93),.WL(WL113));
sram_cell_6t_5 inst_cell_113_94 (.BL(BL94),.BLN(BLN94),.WL(WL113));
sram_cell_6t_5 inst_cell_113_95 (.BL(BL95),.BLN(BLN95),.WL(WL113));
sram_cell_6t_5 inst_cell_113_96 (.BL(BL96),.BLN(BLN96),.WL(WL113));
sram_cell_6t_5 inst_cell_113_97 (.BL(BL97),.BLN(BLN97),.WL(WL113));
sram_cell_6t_5 inst_cell_113_98 (.BL(BL98),.BLN(BLN98),.WL(WL113));
sram_cell_6t_5 inst_cell_113_99 (.BL(BL99),.BLN(BLN99),.WL(WL113));
sram_cell_6t_5 inst_cell_113_100 (.BL(BL100),.BLN(BLN100),.WL(WL113));
sram_cell_6t_5 inst_cell_113_101 (.BL(BL101),.BLN(BLN101),.WL(WL113));
sram_cell_6t_5 inst_cell_113_102 (.BL(BL102),.BLN(BLN102),.WL(WL113));
sram_cell_6t_5 inst_cell_113_103 (.BL(BL103),.BLN(BLN103),.WL(WL113));
sram_cell_6t_5 inst_cell_113_104 (.BL(BL104),.BLN(BLN104),.WL(WL113));
sram_cell_6t_5 inst_cell_113_105 (.BL(BL105),.BLN(BLN105),.WL(WL113));
sram_cell_6t_5 inst_cell_113_106 (.BL(BL106),.BLN(BLN106),.WL(WL113));
sram_cell_6t_5 inst_cell_113_107 (.BL(BL107),.BLN(BLN107),.WL(WL113));
sram_cell_6t_5 inst_cell_113_108 (.BL(BL108),.BLN(BLN108),.WL(WL113));
sram_cell_6t_5 inst_cell_113_109 (.BL(BL109),.BLN(BLN109),.WL(WL113));
sram_cell_6t_5 inst_cell_113_110 (.BL(BL110),.BLN(BLN110),.WL(WL113));
sram_cell_6t_5 inst_cell_113_111 (.BL(BL111),.BLN(BLN111),.WL(WL113));
sram_cell_6t_5 inst_cell_113_112 (.BL(BL112),.BLN(BLN112),.WL(WL113));
sram_cell_6t_5 inst_cell_113_113 (.BL(BL113),.BLN(BLN113),.WL(WL113));
sram_cell_6t_5 inst_cell_113_114 (.BL(BL114),.BLN(BLN114),.WL(WL113));
sram_cell_6t_5 inst_cell_113_115 (.BL(BL115),.BLN(BLN115),.WL(WL113));
sram_cell_6t_5 inst_cell_113_116 (.BL(BL116),.BLN(BLN116),.WL(WL113));
sram_cell_6t_5 inst_cell_113_117 (.BL(BL117),.BLN(BLN117),.WL(WL113));
sram_cell_6t_5 inst_cell_113_118 (.BL(BL118),.BLN(BLN118),.WL(WL113));
sram_cell_6t_5 inst_cell_113_119 (.BL(BL119),.BLN(BLN119),.WL(WL113));
sram_cell_6t_5 inst_cell_113_120 (.BL(BL120),.BLN(BLN120),.WL(WL113));
sram_cell_6t_5 inst_cell_113_121 (.BL(BL121),.BLN(BLN121),.WL(WL113));
sram_cell_6t_5 inst_cell_113_122 (.BL(BL122),.BLN(BLN122),.WL(WL113));
sram_cell_6t_5 inst_cell_113_123 (.BL(BL123),.BLN(BLN123),.WL(WL113));
sram_cell_6t_5 inst_cell_113_124 (.BL(BL124),.BLN(BLN124),.WL(WL113));
sram_cell_6t_5 inst_cell_113_125 (.BL(BL125),.BLN(BLN125),.WL(WL113));
sram_cell_6t_5 inst_cell_113_126 (.BL(BL126),.BLN(BLN126),.WL(WL113));
sram_cell_6t_5 inst_cell_113_127 (.BL(BL127),.BLN(BLN127),.WL(WL113));
sram_cell_6t_5 inst_cell_114_0 (.BL(BL0),.BLN(BLN0),.WL(WL114));
sram_cell_6t_5 inst_cell_114_1 (.BL(BL1),.BLN(BLN1),.WL(WL114));
sram_cell_6t_5 inst_cell_114_2 (.BL(BL2),.BLN(BLN2),.WL(WL114));
sram_cell_6t_5 inst_cell_114_3 (.BL(BL3),.BLN(BLN3),.WL(WL114));
sram_cell_6t_5 inst_cell_114_4 (.BL(BL4),.BLN(BLN4),.WL(WL114));
sram_cell_6t_5 inst_cell_114_5 (.BL(BL5),.BLN(BLN5),.WL(WL114));
sram_cell_6t_5 inst_cell_114_6 (.BL(BL6),.BLN(BLN6),.WL(WL114));
sram_cell_6t_5 inst_cell_114_7 (.BL(BL7),.BLN(BLN7),.WL(WL114));
sram_cell_6t_5 inst_cell_114_8 (.BL(BL8),.BLN(BLN8),.WL(WL114));
sram_cell_6t_5 inst_cell_114_9 (.BL(BL9),.BLN(BLN9),.WL(WL114));
sram_cell_6t_5 inst_cell_114_10 (.BL(BL10),.BLN(BLN10),.WL(WL114));
sram_cell_6t_5 inst_cell_114_11 (.BL(BL11),.BLN(BLN11),.WL(WL114));
sram_cell_6t_5 inst_cell_114_12 (.BL(BL12),.BLN(BLN12),.WL(WL114));
sram_cell_6t_5 inst_cell_114_13 (.BL(BL13),.BLN(BLN13),.WL(WL114));
sram_cell_6t_5 inst_cell_114_14 (.BL(BL14),.BLN(BLN14),.WL(WL114));
sram_cell_6t_5 inst_cell_114_15 (.BL(BL15),.BLN(BLN15),.WL(WL114));
sram_cell_6t_5 inst_cell_114_16 (.BL(BL16),.BLN(BLN16),.WL(WL114));
sram_cell_6t_5 inst_cell_114_17 (.BL(BL17),.BLN(BLN17),.WL(WL114));
sram_cell_6t_5 inst_cell_114_18 (.BL(BL18),.BLN(BLN18),.WL(WL114));
sram_cell_6t_5 inst_cell_114_19 (.BL(BL19),.BLN(BLN19),.WL(WL114));
sram_cell_6t_5 inst_cell_114_20 (.BL(BL20),.BLN(BLN20),.WL(WL114));
sram_cell_6t_5 inst_cell_114_21 (.BL(BL21),.BLN(BLN21),.WL(WL114));
sram_cell_6t_5 inst_cell_114_22 (.BL(BL22),.BLN(BLN22),.WL(WL114));
sram_cell_6t_5 inst_cell_114_23 (.BL(BL23),.BLN(BLN23),.WL(WL114));
sram_cell_6t_5 inst_cell_114_24 (.BL(BL24),.BLN(BLN24),.WL(WL114));
sram_cell_6t_5 inst_cell_114_25 (.BL(BL25),.BLN(BLN25),.WL(WL114));
sram_cell_6t_5 inst_cell_114_26 (.BL(BL26),.BLN(BLN26),.WL(WL114));
sram_cell_6t_5 inst_cell_114_27 (.BL(BL27),.BLN(BLN27),.WL(WL114));
sram_cell_6t_5 inst_cell_114_28 (.BL(BL28),.BLN(BLN28),.WL(WL114));
sram_cell_6t_5 inst_cell_114_29 (.BL(BL29),.BLN(BLN29),.WL(WL114));
sram_cell_6t_5 inst_cell_114_30 (.BL(BL30),.BLN(BLN30),.WL(WL114));
sram_cell_6t_5 inst_cell_114_31 (.BL(BL31),.BLN(BLN31),.WL(WL114));
sram_cell_6t_5 inst_cell_114_32 (.BL(BL32),.BLN(BLN32),.WL(WL114));
sram_cell_6t_5 inst_cell_114_33 (.BL(BL33),.BLN(BLN33),.WL(WL114));
sram_cell_6t_5 inst_cell_114_34 (.BL(BL34),.BLN(BLN34),.WL(WL114));
sram_cell_6t_5 inst_cell_114_35 (.BL(BL35),.BLN(BLN35),.WL(WL114));
sram_cell_6t_5 inst_cell_114_36 (.BL(BL36),.BLN(BLN36),.WL(WL114));
sram_cell_6t_5 inst_cell_114_37 (.BL(BL37),.BLN(BLN37),.WL(WL114));
sram_cell_6t_5 inst_cell_114_38 (.BL(BL38),.BLN(BLN38),.WL(WL114));
sram_cell_6t_5 inst_cell_114_39 (.BL(BL39),.BLN(BLN39),.WL(WL114));
sram_cell_6t_5 inst_cell_114_40 (.BL(BL40),.BLN(BLN40),.WL(WL114));
sram_cell_6t_5 inst_cell_114_41 (.BL(BL41),.BLN(BLN41),.WL(WL114));
sram_cell_6t_5 inst_cell_114_42 (.BL(BL42),.BLN(BLN42),.WL(WL114));
sram_cell_6t_5 inst_cell_114_43 (.BL(BL43),.BLN(BLN43),.WL(WL114));
sram_cell_6t_5 inst_cell_114_44 (.BL(BL44),.BLN(BLN44),.WL(WL114));
sram_cell_6t_5 inst_cell_114_45 (.BL(BL45),.BLN(BLN45),.WL(WL114));
sram_cell_6t_5 inst_cell_114_46 (.BL(BL46),.BLN(BLN46),.WL(WL114));
sram_cell_6t_5 inst_cell_114_47 (.BL(BL47),.BLN(BLN47),.WL(WL114));
sram_cell_6t_5 inst_cell_114_48 (.BL(BL48),.BLN(BLN48),.WL(WL114));
sram_cell_6t_5 inst_cell_114_49 (.BL(BL49),.BLN(BLN49),.WL(WL114));
sram_cell_6t_5 inst_cell_114_50 (.BL(BL50),.BLN(BLN50),.WL(WL114));
sram_cell_6t_5 inst_cell_114_51 (.BL(BL51),.BLN(BLN51),.WL(WL114));
sram_cell_6t_5 inst_cell_114_52 (.BL(BL52),.BLN(BLN52),.WL(WL114));
sram_cell_6t_5 inst_cell_114_53 (.BL(BL53),.BLN(BLN53),.WL(WL114));
sram_cell_6t_5 inst_cell_114_54 (.BL(BL54),.BLN(BLN54),.WL(WL114));
sram_cell_6t_5 inst_cell_114_55 (.BL(BL55),.BLN(BLN55),.WL(WL114));
sram_cell_6t_5 inst_cell_114_56 (.BL(BL56),.BLN(BLN56),.WL(WL114));
sram_cell_6t_5 inst_cell_114_57 (.BL(BL57),.BLN(BLN57),.WL(WL114));
sram_cell_6t_5 inst_cell_114_58 (.BL(BL58),.BLN(BLN58),.WL(WL114));
sram_cell_6t_5 inst_cell_114_59 (.BL(BL59),.BLN(BLN59),.WL(WL114));
sram_cell_6t_5 inst_cell_114_60 (.BL(BL60),.BLN(BLN60),.WL(WL114));
sram_cell_6t_5 inst_cell_114_61 (.BL(BL61),.BLN(BLN61),.WL(WL114));
sram_cell_6t_5 inst_cell_114_62 (.BL(BL62),.BLN(BLN62),.WL(WL114));
sram_cell_6t_5 inst_cell_114_63 (.BL(BL63),.BLN(BLN63),.WL(WL114));
sram_cell_6t_5 inst_cell_114_64 (.BL(BL64),.BLN(BLN64),.WL(WL114));
sram_cell_6t_5 inst_cell_114_65 (.BL(BL65),.BLN(BLN65),.WL(WL114));
sram_cell_6t_5 inst_cell_114_66 (.BL(BL66),.BLN(BLN66),.WL(WL114));
sram_cell_6t_5 inst_cell_114_67 (.BL(BL67),.BLN(BLN67),.WL(WL114));
sram_cell_6t_5 inst_cell_114_68 (.BL(BL68),.BLN(BLN68),.WL(WL114));
sram_cell_6t_5 inst_cell_114_69 (.BL(BL69),.BLN(BLN69),.WL(WL114));
sram_cell_6t_5 inst_cell_114_70 (.BL(BL70),.BLN(BLN70),.WL(WL114));
sram_cell_6t_5 inst_cell_114_71 (.BL(BL71),.BLN(BLN71),.WL(WL114));
sram_cell_6t_5 inst_cell_114_72 (.BL(BL72),.BLN(BLN72),.WL(WL114));
sram_cell_6t_5 inst_cell_114_73 (.BL(BL73),.BLN(BLN73),.WL(WL114));
sram_cell_6t_5 inst_cell_114_74 (.BL(BL74),.BLN(BLN74),.WL(WL114));
sram_cell_6t_5 inst_cell_114_75 (.BL(BL75),.BLN(BLN75),.WL(WL114));
sram_cell_6t_5 inst_cell_114_76 (.BL(BL76),.BLN(BLN76),.WL(WL114));
sram_cell_6t_5 inst_cell_114_77 (.BL(BL77),.BLN(BLN77),.WL(WL114));
sram_cell_6t_5 inst_cell_114_78 (.BL(BL78),.BLN(BLN78),.WL(WL114));
sram_cell_6t_5 inst_cell_114_79 (.BL(BL79),.BLN(BLN79),.WL(WL114));
sram_cell_6t_5 inst_cell_114_80 (.BL(BL80),.BLN(BLN80),.WL(WL114));
sram_cell_6t_5 inst_cell_114_81 (.BL(BL81),.BLN(BLN81),.WL(WL114));
sram_cell_6t_5 inst_cell_114_82 (.BL(BL82),.BLN(BLN82),.WL(WL114));
sram_cell_6t_5 inst_cell_114_83 (.BL(BL83),.BLN(BLN83),.WL(WL114));
sram_cell_6t_5 inst_cell_114_84 (.BL(BL84),.BLN(BLN84),.WL(WL114));
sram_cell_6t_5 inst_cell_114_85 (.BL(BL85),.BLN(BLN85),.WL(WL114));
sram_cell_6t_5 inst_cell_114_86 (.BL(BL86),.BLN(BLN86),.WL(WL114));
sram_cell_6t_5 inst_cell_114_87 (.BL(BL87),.BLN(BLN87),.WL(WL114));
sram_cell_6t_5 inst_cell_114_88 (.BL(BL88),.BLN(BLN88),.WL(WL114));
sram_cell_6t_5 inst_cell_114_89 (.BL(BL89),.BLN(BLN89),.WL(WL114));
sram_cell_6t_5 inst_cell_114_90 (.BL(BL90),.BLN(BLN90),.WL(WL114));
sram_cell_6t_5 inst_cell_114_91 (.BL(BL91),.BLN(BLN91),.WL(WL114));
sram_cell_6t_5 inst_cell_114_92 (.BL(BL92),.BLN(BLN92),.WL(WL114));
sram_cell_6t_5 inst_cell_114_93 (.BL(BL93),.BLN(BLN93),.WL(WL114));
sram_cell_6t_5 inst_cell_114_94 (.BL(BL94),.BLN(BLN94),.WL(WL114));
sram_cell_6t_5 inst_cell_114_95 (.BL(BL95),.BLN(BLN95),.WL(WL114));
sram_cell_6t_5 inst_cell_114_96 (.BL(BL96),.BLN(BLN96),.WL(WL114));
sram_cell_6t_5 inst_cell_114_97 (.BL(BL97),.BLN(BLN97),.WL(WL114));
sram_cell_6t_5 inst_cell_114_98 (.BL(BL98),.BLN(BLN98),.WL(WL114));
sram_cell_6t_5 inst_cell_114_99 (.BL(BL99),.BLN(BLN99),.WL(WL114));
sram_cell_6t_5 inst_cell_114_100 (.BL(BL100),.BLN(BLN100),.WL(WL114));
sram_cell_6t_5 inst_cell_114_101 (.BL(BL101),.BLN(BLN101),.WL(WL114));
sram_cell_6t_5 inst_cell_114_102 (.BL(BL102),.BLN(BLN102),.WL(WL114));
sram_cell_6t_5 inst_cell_114_103 (.BL(BL103),.BLN(BLN103),.WL(WL114));
sram_cell_6t_5 inst_cell_114_104 (.BL(BL104),.BLN(BLN104),.WL(WL114));
sram_cell_6t_5 inst_cell_114_105 (.BL(BL105),.BLN(BLN105),.WL(WL114));
sram_cell_6t_5 inst_cell_114_106 (.BL(BL106),.BLN(BLN106),.WL(WL114));
sram_cell_6t_5 inst_cell_114_107 (.BL(BL107),.BLN(BLN107),.WL(WL114));
sram_cell_6t_5 inst_cell_114_108 (.BL(BL108),.BLN(BLN108),.WL(WL114));
sram_cell_6t_5 inst_cell_114_109 (.BL(BL109),.BLN(BLN109),.WL(WL114));
sram_cell_6t_5 inst_cell_114_110 (.BL(BL110),.BLN(BLN110),.WL(WL114));
sram_cell_6t_5 inst_cell_114_111 (.BL(BL111),.BLN(BLN111),.WL(WL114));
sram_cell_6t_5 inst_cell_114_112 (.BL(BL112),.BLN(BLN112),.WL(WL114));
sram_cell_6t_5 inst_cell_114_113 (.BL(BL113),.BLN(BLN113),.WL(WL114));
sram_cell_6t_5 inst_cell_114_114 (.BL(BL114),.BLN(BLN114),.WL(WL114));
sram_cell_6t_5 inst_cell_114_115 (.BL(BL115),.BLN(BLN115),.WL(WL114));
sram_cell_6t_5 inst_cell_114_116 (.BL(BL116),.BLN(BLN116),.WL(WL114));
sram_cell_6t_5 inst_cell_114_117 (.BL(BL117),.BLN(BLN117),.WL(WL114));
sram_cell_6t_5 inst_cell_114_118 (.BL(BL118),.BLN(BLN118),.WL(WL114));
sram_cell_6t_5 inst_cell_114_119 (.BL(BL119),.BLN(BLN119),.WL(WL114));
sram_cell_6t_5 inst_cell_114_120 (.BL(BL120),.BLN(BLN120),.WL(WL114));
sram_cell_6t_5 inst_cell_114_121 (.BL(BL121),.BLN(BLN121),.WL(WL114));
sram_cell_6t_5 inst_cell_114_122 (.BL(BL122),.BLN(BLN122),.WL(WL114));
sram_cell_6t_5 inst_cell_114_123 (.BL(BL123),.BLN(BLN123),.WL(WL114));
sram_cell_6t_5 inst_cell_114_124 (.BL(BL124),.BLN(BLN124),.WL(WL114));
sram_cell_6t_5 inst_cell_114_125 (.BL(BL125),.BLN(BLN125),.WL(WL114));
sram_cell_6t_5 inst_cell_114_126 (.BL(BL126),.BLN(BLN126),.WL(WL114));
sram_cell_6t_5 inst_cell_114_127 (.BL(BL127),.BLN(BLN127),.WL(WL114));
sram_cell_6t_5 inst_cell_115_0 (.BL(BL0),.BLN(BLN0),.WL(WL115));
sram_cell_6t_5 inst_cell_115_1 (.BL(BL1),.BLN(BLN1),.WL(WL115));
sram_cell_6t_5 inst_cell_115_2 (.BL(BL2),.BLN(BLN2),.WL(WL115));
sram_cell_6t_5 inst_cell_115_3 (.BL(BL3),.BLN(BLN3),.WL(WL115));
sram_cell_6t_5 inst_cell_115_4 (.BL(BL4),.BLN(BLN4),.WL(WL115));
sram_cell_6t_5 inst_cell_115_5 (.BL(BL5),.BLN(BLN5),.WL(WL115));
sram_cell_6t_5 inst_cell_115_6 (.BL(BL6),.BLN(BLN6),.WL(WL115));
sram_cell_6t_5 inst_cell_115_7 (.BL(BL7),.BLN(BLN7),.WL(WL115));
sram_cell_6t_5 inst_cell_115_8 (.BL(BL8),.BLN(BLN8),.WL(WL115));
sram_cell_6t_5 inst_cell_115_9 (.BL(BL9),.BLN(BLN9),.WL(WL115));
sram_cell_6t_5 inst_cell_115_10 (.BL(BL10),.BLN(BLN10),.WL(WL115));
sram_cell_6t_5 inst_cell_115_11 (.BL(BL11),.BLN(BLN11),.WL(WL115));
sram_cell_6t_5 inst_cell_115_12 (.BL(BL12),.BLN(BLN12),.WL(WL115));
sram_cell_6t_5 inst_cell_115_13 (.BL(BL13),.BLN(BLN13),.WL(WL115));
sram_cell_6t_5 inst_cell_115_14 (.BL(BL14),.BLN(BLN14),.WL(WL115));
sram_cell_6t_5 inst_cell_115_15 (.BL(BL15),.BLN(BLN15),.WL(WL115));
sram_cell_6t_5 inst_cell_115_16 (.BL(BL16),.BLN(BLN16),.WL(WL115));
sram_cell_6t_5 inst_cell_115_17 (.BL(BL17),.BLN(BLN17),.WL(WL115));
sram_cell_6t_5 inst_cell_115_18 (.BL(BL18),.BLN(BLN18),.WL(WL115));
sram_cell_6t_5 inst_cell_115_19 (.BL(BL19),.BLN(BLN19),.WL(WL115));
sram_cell_6t_5 inst_cell_115_20 (.BL(BL20),.BLN(BLN20),.WL(WL115));
sram_cell_6t_5 inst_cell_115_21 (.BL(BL21),.BLN(BLN21),.WL(WL115));
sram_cell_6t_5 inst_cell_115_22 (.BL(BL22),.BLN(BLN22),.WL(WL115));
sram_cell_6t_5 inst_cell_115_23 (.BL(BL23),.BLN(BLN23),.WL(WL115));
sram_cell_6t_5 inst_cell_115_24 (.BL(BL24),.BLN(BLN24),.WL(WL115));
sram_cell_6t_5 inst_cell_115_25 (.BL(BL25),.BLN(BLN25),.WL(WL115));
sram_cell_6t_5 inst_cell_115_26 (.BL(BL26),.BLN(BLN26),.WL(WL115));
sram_cell_6t_5 inst_cell_115_27 (.BL(BL27),.BLN(BLN27),.WL(WL115));
sram_cell_6t_5 inst_cell_115_28 (.BL(BL28),.BLN(BLN28),.WL(WL115));
sram_cell_6t_5 inst_cell_115_29 (.BL(BL29),.BLN(BLN29),.WL(WL115));
sram_cell_6t_5 inst_cell_115_30 (.BL(BL30),.BLN(BLN30),.WL(WL115));
sram_cell_6t_5 inst_cell_115_31 (.BL(BL31),.BLN(BLN31),.WL(WL115));
sram_cell_6t_5 inst_cell_115_32 (.BL(BL32),.BLN(BLN32),.WL(WL115));
sram_cell_6t_5 inst_cell_115_33 (.BL(BL33),.BLN(BLN33),.WL(WL115));
sram_cell_6t_5 inst_cell_115_34 (.BL(BL34),.BLN(BLN34),.WL(WL115));
sram_cell_6t_5 inst_cell_115_35 (.BL(BL35),.BLN(BLN35),.WL(WL115));
sram_cell_6t_5 inst_cell_115_36 (.BL(BL36),.BLN(BLN36),.WL(WL115));
sram_cell_6t_5 inst_cell_115_37 (.BL(BL37),.BLN(BLN37),.WL(WL115));
sram_cell_6t_5 inst_cell_115_38 (.BL(BL38),.BLN(BLN38),.WL(WL115));
sram_cell_6t_5 inst_cell_115_39 (.BL(BL39),.BLN(BLN39),.WL(WL115));
sram_cell_6t_5 inst_cell_115_40 (.BL(BL40),.BLN(BLN40),.WL(WL115));
sram_cell_6t_5 inst_cell_115_41 (.BL(BL41),.BLN(BLN41),.WL(WL115));
sram_cell_6t_5 inst_cell_115_42 (.BL(BL42),.BLN(BLN42),.WL(WL115));
sram_cell_6t_5 inst_cell_115_43 (.BL(BL43),.BLN(BLN43),.WL(WL115));
sram_cell_6t_5 inst_cell_115_44 (.BL(BL44),.BLN(BLN44),.WL(WL115));
sram_cell_6t_5 inst_cell_115_45 (.BL(BL45),.BLN(BLN45),.WL(WL115));
sram_cell_6t_5 inst_cell_115_46 (.BL(BL46),.BLN(BLN46),.WL(WL115));
sram_cell_6t_5 inst_cell_115_47 (.BL(BL47),.BLN(BLN47),.WL(WL115));
sram_cell_6t_5 inst_cell_115_48 (.BL(BL48),.BLN(BLN48),.WL(WL115));
sram_cell_6t_5 inst_cell_115_49 (.BL(BL49),.BLN(BLN49),.WL(WL115));
sram_cell_6t_5 inst_cell_115_50 (.BL(BL50),.BLN(BLN50),.WL(WL115));
sram_cell_6t_5 inst_cell_115_51 (.BL(BL51),.BLN(BLN51),.WL(WL115));
sram_cell_6t_5 inst_cell_115_52 (.BL(BL52),.BLN(BLN52),.WL(WL115));
sram_cell_6t_5 inst_cell_115_53 (.BL(BL53),.BLN(BLN53),.WL(WL115));
sram_cell_6t_5 inst_cell_115_54 (.BL(BL54),.BLN(BLN54),.WL(WL115));
sram_cell_6t_5 inst_cell_115_55 (.BL(BL55),.BLN(BLN55),.WL(WL115));
sram_cell_6t_5 inst_cell_115_56 (.BL(BL56),.BLN(BLN56),.WL(WL115));
sram_cell_6t_5 inst_cell_115_57 (.BL(BL57),.BLN(BLN57),.WL(WL115));
sram_cell_6t_5 inst_cell_115_58 (.BL(BL58),.BLN(BLN58),.WL(WL115));
sram_cell_6t_5 inst_cell_115_59 (.BL(BL59),.BLN(BLN59),.WL(WL115));
sram_cell_6t_5 inst_cell_115_60 (.BL(BL60),.BLN(BLN60),.WL(WL115));
sram_cell_6t_5 inst_cell_115_61 (.BL(BL61),.BLN(BLN61),.WL(WL115));
sram_cell_6t_5 inst_cell_115_62 (.BL(BL62),.BLN(BLN62),.WL(WL115));
sram_cell_6t_5 inst_cell_115_63 (.BL(BL63),.BLN(BLN63),.WL(WL115));
sram_cell_6t_5 inst_cell_115_64 (.BL(BL64),.BLN(BLN64),.WL(WL115));
sram_cell_6t_5 inst_cell_115_65 (.BL(BL65),.BLN(BLN65),.WL(WL115));
sram_cell_6t_5 inst_cell_115_66 (.BL(BL66),.BLN(BLN66),.WL(WL115));
sram_cell_6t_5 inst_cell_115_67 (.BL(BL67),.BLN(BLN67),.WL(WL115));
sram_cell_6t_5 inst_cell_115_68 (.BL(BL68),.BLN(BLN68),.WL(WL115));
sram_cell_6t_5 inst_cell_115_69 (.BL(BL69),.BLN(BLN69),.WL(WL115));
sram_cell_6t_5 inst_cell_115_70 (.BL(BL70),.BLN(BLN70),.WL(WL115));
sram_cell_6t_5 inst_cell_115_71 (.BL(BL71),.BLN(BLN71),.WL(WL115));
sram_cell_6t_5 inst_cell_115_72 (.BL(BL72),.BLN(BLN72),.WL(WL115));
sram_cell_6t_5 inst_cell_115_73 (.BL(BL73),.BLN(BLN73),.WL(WL115));
sram_cell_6t_5 inst_cell_115_74 (.BL(BL74),.BLN(BLN74),.WL(WL115));
sram_cell_6t_5 inst_cell_115_75 (.BL(BL75),.BLN(BLN75),.WL(WL115));
sram_cell_6t_5 inst_cell_115_76 (.BL(BL76),.BLN(BLN76),.WL(WL115));
sram_cell_6t_5 inst_cell_115_77 (.BL(BL77),.BLN(BLN77),.WL(WL115));
sram_cell_6t_5 inst_cell_115_78 (.BL(BL78),.BLN(BLN78),.WL(WL115));
sram_cell_6t_5 inst_cell_115_79 (.BL(BL79),.BLN(BLN79),.WL(WL115));
sram_cell_6t_5 inst_cell_115_80 (.BL(BL80),.BLN(BLN80),.WL(WL115));
sram_cell_6t_5 inst_cell_115_81 (.BL(BL81),.BLN(BLN81),.WL(WL115));
sram_cell_6t_5 inst_cell_115_82 (.BL(BL82),.BLN(BLN82),.WL(WL115));
sram_cell_6t_5 inst_cell_115_83 (.BL(BL83),.BLN(BLN83),.WL(WL115));
sram_cell_6t_5 inst_cell_115_84 (.BL(BL84),.BLN(BLN84),.WL(WL115));
sram_cell_6t_5 inst_cell_115_85 (.BL(BL85),.BLN(BLN85),.WL(WL115));
sram_cell_6t_5 inst_cell_115_86 (.BL(BL86),.BLN(BLN86),.WL(WL115));
sram_cell_6t_5 inst_cell_115_87 (.BL(BL87),.BLN(BLN87),.WL(WL115));
sram_cell_6t_5 inst_cell_115_88 (.BL(BL88),.BLN(BLN88),.WL(WL115));
sram_cell_6t_5 inst_cell_115_89 (.BL(BL89),.BLN(BLN89),.WL(WL115));
sram_cell_6t_5 inst_cell_115_90 (.BL(BL90),.BLN(BLN90),.WL(WL115));
sram_cell_6t_5 inst_cell_115_91 (.BL(BL91),.BLN(BLN91),.WL(WL115));
sram_cell_6t_5 inst_cell_115_92 (.BL(BL92),.BLN(BLN92),.WL(WL115));
sram_cell_6t_5 inst_cell_115_93 (.BL(BL93),.BLN(BLN93),.WL(WL115));
sram_cell_6t_5 inst_cell_115_94 (.BL(BL94),.BLN(BLN94),.WL(WL115));
sram_cell_6t_5 inst_cell_115_95 (.BL(BL95),.BLN(BLN95),.WL(WL115));
sram_cell_6t_5 inst_cell_115_96 (.BL(BL96),.BLN(BLN96),.WL(WL115));
sram_cell_6t_5 inst_cell_115_97 (.BL(BL97),.BLN(BLN97),.WL(WL115));
sram_cell_6t_5 inst_cell_115_98 (.BL(BL98),.BLN(BLN98),.WL(WL115));
sram_cell_6t_5 inst_cell_115_99 (.BL(BL99),.BLN(BLN99),.WL(WL115));
sram_cell_6t_5 inst_cell_115_100 (.BL(BL100),.BLN(BLN100),.WL(WL115));
sram_cell_6t_5 inst_cell_115_101 (.BL(BL101),.BLN(BLN101),.WL(WL115));
sram_cell_6t_5 inst_cell_115_102 (.BL(BL102),.BLN(BLN102),.WL(WL115));
sram_cell_6t_5 inst_cell_115_103 (.BL(BL103),.BLN(BLN103),.WL(WL115));
sram_cell_6t_5 inst_cell_115_104 (.BL(BL104),.BLN(BLN104),.WL(WL115));
sram_cell_6t_5 inst_cell_115_105 (.BL(BL105),.BLN(BLN105),.WL(WL115));
sram_cell_6t_5 inst_cell_115_106 (.BL(BL106),.BLN(BLN106),.WL(WL115));
sram_cell_6t_5 inst_cell_115_107 (.BL(BL107),.BLN(BLN107),.WL(WL115));
sram_cell_6t_5 inst_cell_115_108 (.BL(BL108),.BLN(BLN108),.WL(WL115));
sram_cell_6t_5 inst_cell_115_109 (.BL(BL109),.BLN(BLN109),.WL(WL115));
sram_cell_6t_5 inst_cell_115_110 (.BL(BL110),.BLN(BLN110),.WL(WL115));
sram_cell_6t_5 inst_cell_115_111 (.BL(BL111),.BLN(BLN111),.WL(WL115));
sram_cell_6t_5 inst_cell_115_112 (.BL(BL112),.BLN(BLN112),.WL(WL115));
sram_cell_6t_5 inst_cell_115_113 (.BL(BL113),.BLN(BLN113),.WL(WL115));
sram_cell_6t_5 inst_cell_115_114 (.BL(BL114),.BLN(BLN114),.WL(WL115));
sram_cell_6t_5 inst_cell_115_115 (.BL(BL115),.BLN(BLN115),.WL(WL115));
sram_cell_6t_5 inst_cell_115_116 (.BL(BL116),.BLN(BLN116),.WL(WL115));
sram_cell_6t_5 inst_cell_115_117 (.BL(BL117),.BLN(BLN117),.WL(WL115));
sram_cell_6t_5 inst_cell_115_118 (.BL(BL118),.BLN(BLN118),.WL(WL115));
sram_cell_6t_5 inst_cell_115_119 (.BL(BL119),.BLN(BLN119),.WL(WL115));
sram_cell_6t_5 inst_cell_115_120 (.BL(BL120),.BLN(BLN120),.WL(WL115));
sram_cell_6t_5 inst_cell_115_121 (.BL(BL121),.BLN(BLN121),.WL(WL115));
sram_cell_6t_5 inst_cell_115_122 (.BL(BL122),.BLN(BLN122),.WL(WL115));
sram_cell_6t_5 inst_cell_115_123 (.BL(BL123),.BLN(BLN123),.WL(WL115));
sram_cell_6t_5 inst_cell_115_124 (.BL(BL124),.BLN(BLN124),.WL(WL115));
sram_cell_6t_5 inst_cell_115_125 (.BL(BL125),.BLN(BLN125),.WL(WL115));
sram_cell_6t_5 inst_cell_115_126 (.BL(BL126),.BLN(BLN126),.WL(WL115));
sram_cell_6t_5 inst_cell_115_127 (.BL(BL127),.BLN(BLN127),.WL(WL115));
sram_cell_6t_5 inst_cell_116_0 (.BL(BL0),.BLN(BLN0),.WL(WL116));
sram_cell_6t_5 inst_cell_116_1 (.BL(BL1),.BLN(BLN1),.WL(WL116));
sram_cell_6t_5 inst_cell_116_2 (.BL(BL2),.BLN(BLN2),.WL(WL116));
sram_cell_6t_5 inst_cell_116_3 (.BL(BL3),.BLN(BLN3),.WL(WL116));
sram_cell_6t_5 inst_cell_116_4 (.BL(BL4),.BLN(BLN4),.WL(WL116));
sram_cell_6t_5 inst_cell_116_5 (.BL(BL5),.BLN(BLN5),.WL(WL116));
sram_cell_6t_5 inst_cell_116_6 (.BL(BL6),.BLN(BLN6),.WL(WL116));
sram_cell_6t_5 inst_cell_116_7 (.BL(BL7),.BLN(BLN7),.WL(WL116));
sram_cell_6t_5 inst_cell_116_8 (.BL(BL8),.BLN(BLN8),.WL(WL116));
sram_cell_6t_5 inst_cell_116_9 (.BL(BL9),.BLN(BLN9),.WL(WL116));
sram_cell_6t_5 inst_cell_116_10 (.BL(BL10),.BLN(BLN10),.WL(WL116));
sram_cell_6t_5 inst_cell_116_11 (.BL(BL11),.BLN(BLN11),.WL(WL116));
sram_cell_6t_5 inst_cell_116_12 (.BL(BL12),.BLN(BLN12),.WL(WL116));
sram_cell_6t_5 inst_cell_116_13 (.BL(BL13),.BLN(BLN13),.WL(WL116));
sram_cell_6t_5 inst_cell_116_14 (.BL(BL14),.BLN(BLN14),.WL(WL116));
sram_cell_6t_5 inst_cell_116_15 (.BL(BL15),.BLN(BLN15),.WL(WL116));
sram_cell_6t_5 inst_cell_116_16 (.BL(BL16),.BLN(BLN16),.WL(WL116));
sram_cell_6t_5 inst_cell_116_17 (.BL(BL17),.BLN(BLN17),.WL(WL116));
sram_cell_6t_5 inst_cell_116_18 (.BL(BL18),.BLN(BLN18),.WL(WL116));
sram_cell_6t_5 inst_cell_116_19 (.BL(BL19),.BLN(BLN19),.WL(WL116));
sram_cell_6t_5 inst_cell_116_20 (.BL(BL20),.BLN(BLN20),.WL(WL116));
sram_cell_6t_5 inst_cell_116_21 (.BL(BL21),.BLN(BLN21),.WL(WL116));
sram_cell_6t_5 inst_cell_116_22 (.BL(BL22),.BLN(BLN22),.WL(WL116));
sram_cell_6t_5 inst_cell_116_23 (.BL(BL23),.BLN(BLN23),.WL(WL116));
sram_cell_6t_5 inst_cell_116_24 (.BL(BL24),.BLN(BLN24),.WL(WL116));
sram_cell_6t_5 inst_cell_116_25 (.BL(BL25),.BLN(BLN25),.WL(WL116));
sram_cell_6t_5 inst_cell_116_26 (.BL(BL26),.BLN(BLN26),.WL(WL116));
sram_cell_6t_5 inst_cell_116_27 (.BL(BL27),.BLN(BLN27),.WL(WL116));
sram_cell_6t_5 inst_cell_116_28 (.BL(BL28),.BLN(BLN28),.WL(WL116));
sram_cell_6t_5 inst_cell_116_29 (.BL(BL29),.BLN(BLN29),.WL(WL116));
sram_cell_6t_5 inst_cell_116_30 (.BL(BL30),.BLN(BLN30),.WL(WL116));
sram_cell_6t_5 inst_cell_116_31 (.BL(BL31),.BLN(BLN31),.WL(WL116));
sram_cell_6t_5 inst_cell_116_32 (.BL(BL32),.BLN(BLN32),.WL(WL116));
sram_cell_6t_5 inst_cell_116_33 (.BL(BL33),.BLN(BLN33),.WL(WL116));
sram_cell_6t_5 inst_cell_116_34 (.BL(BL34),.BLN(BLN34),.WL(WL116));
sram_cell_6t_5 inst_cell_116_35 (.BL(BL35),.BLN(BLN35),.WL(WL116));
sram_cell_6t_5 inst_cell_116_36 (.BL(BL36),.BLN(BLN36),.WL(WL116));
sram_cell_6t_5 inst_cell_116_37 (.BL(BL37),.BLN(BLN37),.WL(WL116));
sram_cell_6t_5 inst_cell_116_38 (.BL(BL38),.BLN(BLN38),.WL(WL116));
sram_cell_6t_5 inst_cell_116_39 (.BL(BL39),.BLN(BLN39),.WL(WL116));
sram_cell_6t_5 inst_cell_116_40 (.BL(BL40),.BLN(BLN40),.WL(WL116));
sram_cell_6t_5 inst_cell_116_41 (.BL(BL41),.BLN(BLN41),.WL(WL116));
sram_cell_6t_5 inst_cell_116_42 (.BL(BL42),.BLN(BLN42),.WL(WL116));
sram_cell_6t_5 inst_cell_116_43 (.BL(BL43),.BLN(BLN43),.WL(WL116));
sram_cell_6t_5 inst_cell_116_44 (.BL(BL44),.BLN(BLN44),.WL(WL116));
sram_cell_6t_5 inst_cell_116_45 (.BL(BL45),.BLN(BLN45),.WL(WL116));
sram_cell_6t_5 inst_cell_116_46 (.BL(BL46),.BLN(BLN46),.WL(WL116));
sram_cell_6t_5 inst_cell_116_47 (.BL(BL47),.BLN(BLN47),.WL(WL116));
sram_cell_6t_5 inst_cell_116_48 (.BL(BL48),.BLN(BLN48),.WL(WL116));
sram_cell_6t_5 inst_cell_116_49 (.BL(BL49),.BLN(BLN49),.WL(WL116));
sram_cell_6t_5 inst_cell_116_50 (.BL(BL50),.BLN(BLN50),.WL(WL116));
sram_cell_6t_5 inst_cell_116_51 (.BL(BL51),.BLN(BLN51),.WL(WL116));
sram_cell_6t_5 inst_cell_116_52 (.BL(BL52),.BLN(BLN52),.WL(WL116));
sram_cell_6t_5 inst_cell_116_53 (.BL(BL53),.BLN(BLN53),.WL(WL116));
sram_cell_6t_5 inst_cell_116_54 (.BL(BL54),.BLN(BLN54),.WL(WL116));
sram_cell_6t_5 inst_cell_116_55 (.BL(BL55),.BLN(BLN55),.WL(WL116));
sram_cell_6t_5 inst_cell_116_56 (.BL(BL56),.BLN(BLN56),.WL(WL116));
sram_cell_6t_5 inst_cell_116_57 (.BL(BL57),.BLN(BLN57),.WL(WL116));
sram_cell_6t_5 inst_cell_116_58 (.BL(BL58),.BLN(BLN58),.WL(WL116));
sram_cell_6t_5 inst_cell_116_59 (.BL(BL59),.BLN(BLN59),.WL(WL116));
sram_cell_6t_5 inst_cell_116_60 (.BL(BL60),.BLN(BLN60),.WL(WL116));
sram_cell_6t_5 inst_cell_116_61 (.BL(BL61),.BLN(BLN61),.WL(WL116));
sram_cell_6t_5 inst_cell_116_62 (.BL(BL62),.BLN(BLN62),.WL(WL116));
sram_cell_6t_5 inst_cell_116_63 (.BL(BL63),.BLN(BLN63),.WL(WL116));
sram_cell_6t_5 inst_cell_116_64 (.BL(BL64),.BLN(BLN64),.WL(WL116));
sram_cell_6t_5 inst_cell_116_65 (.BL(BL65),.BLN(BLN65),.WL(WL116));
sram_cell_6t_5 inst_cell_116_66 (.BL(BL66),.BLN(BLN66),.WL(WL116));
sram_cell_6t_5 inst_cell_116_67 (.BL(BL67),.BLN(BLN67),.WL(WL116));
sram_cell_6t_5 inst_cell_116_68 (.BL(BL68),.BLN(BLN68),.WL(WL116));
sram_cell_6t_5 inst_cell_116_69 (.BL(BL69),.BLN(BLN69),.WL(WL116));
sram_cell_6t_5 inst_cell_116_70 (.BL(BL70),.BLN(BLN70),.WL(WL116));
sram_cell_6t_5 inst_cell_116_71 (.BL(BL71),.BLN(BLN71),.WL(WL116));
sram_cell_6t_5 inst_cell_116_72 (.BL(BL72),.BLN(BLN72),.WL(WL116));
sram_cell_6t_5 inst_cell_116_73 (.BL(BL73),.BLN(BLN73),.WL(WL116));
sram_cell_6t_5 inst_cell_116_74 (.BL(BL74),.BLN(BLN74),.WL(WL116));
sram_cell_6t_5 inst_cell_116_75 (.BL(BL75),.BLN(BLN75),.WL(WL116));
sram_cell_6t_5 inst_cell_116_76 (.BL(BL76),.BLN(BLN76),.WL(WL116));
sram_cell_6t_5 inst_cell_116_77 (.BL(BL77),.BLN(BLN77),.WL(WL116));
sram_cell_6t_5 inst_cell_116_78 (.BL(BL78),.BLN(BLN78),.WL(WL116));
sram_cell_6t_5 inst_cell_116_79 (.BL(BL79),.BLN(BLN79),.WL(WL116));
sram_cell_6t_5 inst_cell_116_80 (.BL(BL80),.BLN(BLN80),.WL(WL116));
sram_cell_6t_5 inst_cell_116_81 (.BL(BL81),.BLN(BLN81),.WL(WL116));
sram_cell_6t_5 inst_cell_116_82 (.BL(BL82),.BLN(BLN82),.WL(WL116));
sram_cell_6t_5 inst_cell_116_83 (.BL(BL83),.BLN(BLN83),.WL(WL116));
sram_cell_6t_5 inst_cell_116_84 (.BL(BL84),.BLN(BLN84),.WL(WL116));
sram_cell_6t_5 inst_cell_116_85 (.BL(BL85),.BLN(BLN85),.WL(WL116));
sram_cell_6t_5 inst_cell_116_86 (.BL(BL86),.BLN(BLN86),.WL(WL116));
sram_cell_6t_5 inst_cell_116_87 (.BL(BL87),.BLN(BLN87),.WL(WL116));
sram_cell_6t_5 inst_cell_116_88 (.BL(BL88),.BLN(BLN88),.WL(WL116));
sram_cell_6t_5 inst_cell_116_89 (.BL(BL89),.BLN(BLN89),.WL(WL116));
sram_cell_6t_5 inst_cell_116_90 (.BL(BL90),.BLN(BLN90),.WL(WL116));
sram_cell_6t_5 inst_cell_116_91 (.BL(BL91),.BLN(BLN91),.WL(WL116));
sram_cell_6t_5 inst_cell_116_92 (.BL(BL92),.BLN(BLN92),.WL(WL116));
sram_cell_6t_5 inst_cell_116_93 (.BL(BL93),.BLN(BLN93),.WL(WL116));
sram_cell_6t_5 inst_cell_116_94 (.BL(BL94),.BLN(BLN94),.WL(WL116));
sram_cell_6t_5 inst_cell_116_95 (.BL(BL95),.BLN(BLN95),.WL(WL116));
sram_cell_6t_5 inst_cell_116_96 (.BL(BL96),.BLN(BLN96),.WL(WL116));
sram_cell_6t_5 inst_cell_116_97 (.BL(BL97),.BLN(BLN97),.WL(WL116));
sram_cell_6t_5 inst_cell_116_98 (.BL(BL98),.BLN(BLN98),.WL(WL116));
sram_cell_6t_5 inst_cell_116_99 (.BL(BL99),.BLN(BLN99),.WL(WL116));
sram_cell_6t_5 inst_cell_116_100 (.BL(BL100),.BLN(BLN100),.WL(WL116));
sram_cell_6t_5 inst_cell_116_101 (.BL(BL101),.BLN(BLN101),.WL(WL116));
sram_cell_6t_5 inst_cell_116_102 (.BL(BL102),.BLN(BLN102),.WL(WL116));
sram_cell_6t_5 inst_cell_116_103 (.BL(BL103),.BLN(BLN103),.WL(WL116));
sram_cell_6t_5 inst_cell_116_104 (.BL(BL104),.BLN(BLN104),.WL(WL116));
sram_cell_6t_5 inst_cell_116_105 (.BL(BL105),.BLN(BLN105),.WL(WL116));
sram_cell_6t_5 inst_cell_116_106 (.BL(BL106),.BLN(BLN106),.WL(WL116));
sram_cell_6t_5 inst_cell_116_107 (.BL(BL107),.BLN(BLN107),.WL(WL116));
sram_cell_6t_5 inst_cell_116_108 (.BL(BL108),.BLN(BLN108),.WL(WL116));
sram_cell_6t_5 inst_cell_116_109 (.BL(BL109),.BLN(BLN109),.WL(WL116));
sram_cell_6t_5 inst_cell_116_110 (.BL(BL110),.BLN(BLN110),.WL(WL116));
sram_cell_6t_5 inst_cell_116_111 (.BL(BL111),.BLN(BLN111),.WL(WL116));
sram_cell_6t_5 inst_cell_116_112 (.BL(BL112),.BLN(BLN112),.WL(WL116));
sram_cell_6t_5 inst_cell_116_113 (.BL(BL113),.BLN(BLN113),.WL(WL116));
sram_cell_6t_5 inst_cell_116_114 (.BL(BL114),.BLN(BLN114),.WL(WL116));
sram_cell_6t_5 inst_cell_116_115 (.BL(BL115),.BLN(BLN115),.WL(WL116));
sram_cell_6t_5 inst_cell_116_116 (.BL(BL116),.BLN(BLN116),.WL(WL116));
sram_cell_6t_5 inst_cell_116_117 (.BL(BL117),.BLN(BLN117),.WL(WL116));
sram_cell_6t_5 inst_cell_116_118 (.BL(BL118),.BLN(BLN118),.WL(WL116));
sram_cell_6t_5 inst_cell_116_119 (.BL(BL119),.BLN(BLN119),.WL(WL116));
sram_cell_6t_5 inst_cell_116_120 (.BL(BL120),.BLN(BLN120),.WL(WL116));
sram_cell_6t_5 inst_cell_116_121 (.BL(BL121),.BLN(BLN121),.WL(WL116));
sram_cell_6t_5 inst_cell_116_122 (.BL(BL122),.BLN(BLN122),.WL(WL116));
sram_cell_6t_5 inst_cell_116_123 (.BL(BL123),.BLN(BLN123),.WL(WL116));
sram_cell_6t_5 inst_cell_116_124 (.BL(BL124),.BLN(BLN124),.WL(WL116));
sram_cell_6t_5 inst_cell_116_125 (.BL(BL125),.BLN(BLN125),.WL(WL116));
sram_cell_6t_5 inst_cell_116_126 (.BL(BL126),.BLN(BLN126),.WL(WL116));
sram_cell_6t_5 inst_cell_116_127 (.BL(BL127),.BLN(BLN127),.WL(WL116));
sram_cell_6t_5 inst_cell_117_0 (.BL(BL0),.BLN(BLN0),.WL(WL117));
sram_cell_6t_5 inst_cell_117_1 (.BL(BL1),.BLN(BLN1),.WL(WL117));
sram_cell_6t_5 inst_cell_117_2 (.BL(BL2),.BLN(BLN2),.WL(WL117));
sram_cell_6t_5 inst_cell_117_3 (.BL(BL3),.BLN(BLN3),.WL(WL117));
sram_cell_6t_5 inst_cell_117_4 (.BL(BL4),.BLN(BLN4),.WL(WL117));
sram_cell_6t_5 inst_cell_117_5 (.BL(BL5),.BLN(BLN5),.WL(WL117));
sram_cell_6t_5 inst_cell_117_6 (.BL(BL6),.BLN(BLN6),.WL(WL117));
sram_cell_6t_5 inst_cell_117_7 (.BL(BL7),.BLN(BLN7),.WL(WL117));
sram_cell_6t_5 inst_cell_117_8 (.BL(BL8),.BLN(BLN8),.WL(WL117));
sram_cell_6t_5 inst_cell_117_9 (.BL(BL9),.BLN(BLN9),.WL(WL117));
sram_cell_6t_5 inst_cell_117_10 (.BL(BL10),.BLN(BLN10),.WL(WL117));
sram_cell_6t_5 inst_cell_117_11 (.BL(BL11),.BLN(BLN11),.WL(WL117));
sram_cell_6t_5 inst_cell_117_12 (.BL(BL12),.BLN(BLN12),.WL(WL117));
sram_cell_6t_5 inst_cell_117_13 (.BL(BL13),.BLN(BLN13),.WL(WL117));
sram_cell_6t_5 inst_cell_117_14 (.BL(BL14),.BLN(BLN14),.WL(WL117));
sram_cell_6t_5 inst_cell_117_15 (.BL(BL15),.BLN(BLN15),.WL(WL117));
sram_cell_6t_5 inst_cell_117_16 (.BL(BL16),.BLN(BLN16),.WL(WL117));
sram_cell_6t_5 inst_cell_117_17 (.BL(BL17),.BLN(BLN17),.WL(WL117));
sram_cell_6t_5 inst_cell_117_18 (.BL(BL18),.BLN(BLN18),.WL(WL117));
sram_cell_6t_5 inst_cell_117_19 (.BL(BL19),.BLN(BLN19),.WL(WL117));
sram_cell_6t_5 inst_cell_117_20 (.BL(BL20),.BLN(BLN20),.WL(WL117));
sram_cell_6t_5 inst_cell_117_21 (.BL(BL21),.BLN(BLN21),.WL(WL117));
sram_cell_6t_5 inst_cell_117_22 (.BL(BL22),.BLN(BLN22),.WL(WL117));
sram_cell_6t_5 inst_cell_117_23 (.BL(BL23),.BLN(BLN23),.WL(WL117));
sram_cell_6t_5 inst_cell_117_24 (.BL(BL24),.BLN(BLN24),.WL(WL117));
sram_cell_6t_5 inst_cell_117_25 (.BL(BL25),.BLN(BLN25),.WL(WL117));
sram_cell_6t_5 inst_cell_117_26 (.BL(BL26),.BLN(BLN26),.WL(WL117));
sram_cell_6t_5 inst_cell_117_27 (.BL(BL27),.BLN(BLN27),.WL(WL117));
sram_cell_6t_5 inst_cell_117_28 (.BL(BL28),.BLN(BLN28),.WL(WL117));
sram_cell_6t_5 inst_cell_117_29 (.BL(BL29),.BLN(BLN29),.WL(WL117));
sram_cell_6t_5 inst_cell_117_30 (.BL(BL30),.BLN(BLN30),.WL(WL117));
sram_cell_6t_5 inst_cell_117_31 (.BL(BL31),.BLN(BLN31),.WL(WL117));
sram_cell_6t_5 inst_cell_117_32 (.BL(BL32),.BLN(BLN32),.WL(WL117));
sram_cell_6t_5 inst_cell_117_33 (.BL(BL33),.BLN(BLN33),.WL(WL117));
sram_cell_6t_5 inst_cell_117_34 (.BL(BL34),.BLN(BLN34),.WL(WL117));
sram_cell_6t_5 inst_cell_117_35 (.BL(BL35),.BLN(BLN35),.WL(WL117));
sram_cell_6t_5 inst_cell_117_36 (.BL(BL36),.BLN(BLN36),.WL(WL117));
sram_cell_6t_5 inst_cell_117_37 (.BL(BL37),.BLN(BLN37),.WL(WL117));
sram_cell_6t_5 inst_cell_117_38 (.BL(BL38),.BLN(BLN38),.WL(WL117));
sram_cell_6t_5 inst_cell_117_39 (.BL(BL39),.BLN(BLN39),.WL(WL117));
sram_cell_6t_5 inst_cell_117_40 (.BL(BL40),.BLN(BLN40),.WL(WL117));
sram_cell_6t_5 inst_cell_117_41 (.BL(BL41),.BLN(BLN41),.WL(WL117));
sram_cell_6t_5 inst_cell_117_42 (.BL(BL42),.BLN(BLN42),.WL(WL117));
sram_cell_6t_5 inst_cell_117_43 (.BL(BL43),.BLN(BLN43),.WL(WL117));
sram_cell_6t_5 inst_cell_117_44 (.BL(BL44),.BLN(BLN44),.WL(WL117));
sram_cell_6t_5 inst_cell_117_45 (.BL(BL45),.BLN(BLN45),.WL(WL117));
sram_cell_6t_5 inst_cell_117_46 (.BL(BL46),.BLN(BLN46),.WL(WL117));
sram_cell_6t_5 inst_cell_117_47 (.BL(BL47),.BLN(BLN47),.WL(WL117));
sram_cell_6t_5 inst_cell_117_48 (.BL(BL48),.BLN(BLN48),.WL(WL117));
sram_cell_6t_5 inst_cell_117_49 (.BL(BL49),.BLN(BLN49),.WL(WL117));
sram_cell_6t_5 inst_cell_117_50 (.BL(BL50),.BLN(BLN50),.WL(WL117));
sram_cell_6t_5 inst_cell_117_51 (.BL(BL51),.BLN(BLN51),.WL(WL117));
sram_cell_6t_5 inst_cell_117_52 (.BL(BL52),.BLN(BLN52),.WL(WL117));
sram_cell_6t_5 inst_cell_117_53 (.BL(BL53),.BLN(BLN53),.WL(WL117));
sram_cell_6t_5 inst_cell_117_54 (.BL(BL54),.BLN(BLN54),.WL(WL117));
sram_cell_6t_5 inst_cell_117_55 (.BL(BL55),.BLN(BLN55),.WL(WL117));
sram_cell_6t_5 inst_cell_117_56 (.BL(BL56),.BLN(BLN56),.WL(WL117));
sram_cell_6t_5 inst_cell_117_57 (.BL(BL57),.BLN(BLN57),.WL(WL117));
sram_cell_6t_5 inst_cell_117_58 (.BL(BL58),.BLN(BLN58),.WL(WL117));
sram_cell_6t_5 inst_cell_117_59 (.BL(BL59),.BLN(BLN59),.WL(WL117));
sram_cell_6t_5 inst_cell_117_60 (.BL(BL60),.BLN(BLN60),.WL(WL117));
sram_cell_6t_5 inst_cell_117_61 (.BL(BL61),.BLN(BLN61),.WL(WL117));
sram_cell_6t_5 inst_cell_117_62 (.BL(BL62),.BLN(BLN62),.WL(WL117));
sram_cell_6t_5 inst_cell_117_63 (.BL(BL63),.BLN(BLN63),.WL(WL117));
sram_cell_6t_5 inst_cell_117_64 (.BL(BL64),.BLN(BLN64),.WL(WL117));
sram_cell_6t_5 inst_cell_117_65 (.BL(BL65),.BLN(BLN65),.WL(WL117));
sram_cell_6t_5 inst_cell_117_66 (.BL(BL66),.BLN(BLN66),.WL(WL117));
sram_cell_6t_5 inst_cell_117_67 (.BL(BL67),.BLN(BLN67),.WL(WL117));
sram_cell_6t_5 inst_cell_117_68 (.BL(BL68),.BLN(BLN68),.WL(WL117));
sram_cell_6t_5 inst_cell_117_69 (.BL(BL69),.BLN(BLN69),.WL(WL117));
sram_cell_6t_5 inst_cell_117_70 (.BL(BL70),.BLN(BLN70),.WL(WL117));
sram_cell_6t_5 inst_cell_117_71 (.BL(BL71),.BLN(BLN71),.WL(WL117));
sram_cell_6t_5 inst_cell_117_72 (.BL(BL72),.BLN(BLN72),.WL(WL117));
sram_cell_6t_5 inst_cell_117_73 (.BL(BL73),.BLN(BLN73),.WL(WL117));
sram_cell_6t_5 inst_cell_117_74 (.BL(BL74),.BLN(BLN74),.WL(WL117));
sram_cell_6t_5 inst_cell_117_75 (.BL(BL75),.BLN(BLN75),.WL(WL117));
sram_cell_6t_5 inst_cell_117_76 (.BL(BL76),.BLN(BLN76),.WL(WL117));
sram_cell_6t_5 inst_cell_117_77 (.BL(BL77),.BLN(BLN77),.WL(WL117));
sram_cell_6t_5 inst_cell_117_78 (.BL(BL78),.BLN(BLN78),.WL(WL117));
sram_cell_6t_5 inst_cell_117_79 (.BL(BL79),.BLN(BLN79),.WL(WL117));
sram_cell_6t_5 inst_cell_117_80 (.BL(BL80),.BLN(BLN80),.WL(WL117));
sram_cell_6t_5 inst_cell_117_81 (.BL(BL81),.BLN(BLN81),.WL(WL117));
sram_cell_6t_5 inst_cell_117_82 (.BL(BL82),.BLN(BLN82),.WL(WL117));
sram_cell_6t_5 inst_cell_117_83 (.BL(BL83),.BLN(BLN83),.WL(WL117));
sram_cell_6t_5 inst_cell_117_84 (.BL(BL84),.BLN(BLN84),.WL(WL117));
sram_cell_6t_5 inst_cell_117_85 (.BL(BL85),.BLN(BLN85),.WL(WL117));
sram_cell_6t_5 inst_cell_117_86 (.BL(BL86),.BLN(BLN86),.WL(WL117));
sram_cell_6t_5 inst_cell_117_87 (.BL(BL87),.BLN(BLN87),.WL(WL117));
sram_cell_6t_5 inst_cell_117_88 (.BL(BL88),.BLN(BLN88),.WL(WL117));
sram_cell_6t_5 inst_cell_117_89 (.BL(BL89),.BLN(BLN89),.WL(WL117));
sram_cell_6t_5 inst_cell_117_90 (.BL(BL90),.BLN(BLN90),.WL(WL117));
sram_cell_6t_5 inst_cell_117_91 (.BL(BL91),.BLN(BLN91),.WL(WL117));
sram_cell_6t_5 inst_cell_117_92 (.BL(BL92),.BLN(BLN92),.WL(WL117));
sram_cell_6t_5 inst_cell_117_93 (.BL(BL93),.BLN(BLN93),.WL(WL117));
sram_cell_6t_5 inst_cell_117_94 (.BL(BL94),.BLN(BLN94),.WL(WL117));
sram_cell_6t_5 inst_cell_117_95 (.BL(BL95),.BLN(BLN95),.WL(WL117));
sram_cell_6t_5 inst_cell_117_96 (.BL(BL96),.BLN(BLN96),.WL(WL117));
sram_cell_6t_5 inst_cell_117_97 (.BL(BL97),.BLN(BLN97),.WL(WL117));
sram_cell_6t_5 inst_cell_117_98 (.BL(BL98),.BLN(BLN98),.WL(WL117));
sram_cell_6t_5 inst_cell_117_99 (.BL(BL99),.BLN(BLN99),.WL(WL117));
sram_cell_6t_5 inst_cell_117_100 (.BL(BL100),.BLN(BLN100),.WL(WL117));
sram_cell_6t_5 inst_cell_117_101 (.BL(BL101),.BLN(BLN101),.WL(WL117));
sram_cell_6t_5 inst_cell_117_102 (.BL(BL102),.BLN(BLN102),.WL(WL117));
sram_cell_6t_5 inst_cell_117_103 (.BL(BL103),.BLN(BLN103),.WL(WL117));
sram_cell_6t_5 inst_cell_117_104 (.BL(BL104),.BLN(BLN104),.WL(WL117));
sram_cell_6t_5 inst_cell_117_105 (.BL(BL105),.BLN(BLN105),.WL(WL117));
sram_cell_6t_5 inst_cell_117_106 (.BL(BL106),.BLN(BLN106),.WL(WL117));
sram_cell_6t_5 inst_cell_117_107 (.BL(BL107),.BLN(BLN107),.WL(WL117));
sram_cell_6t_5 inst_cell_117_108 (.BL(BL108),.BLN(BLN108),.WL(WL117));
sram_cell_6t_5 inst_cell_117_109 (.BL(BL109),.BLN(BLN109),.WL(WL117));
sram_cell_6t_5 inst_cell_117_110 (.BL(BL110),.BLN(BLN110),.WL(WL117));
sram_cell_6t_5 inst_cell_117_111 (.BL(BL111),.BLN(BLN111),.WL(WL117));
sram_cell_6t_5 inst_cell_117_112 (.BL(BL112),.BLN(BLN112),.WL(WL117));
sram_cell_6t_5 inst_cell_117_113 (.BL(BL113),.BLN(BLN113),.WL(WL117));
sram_cell_6t_5 inst_cell_117_114 (.BL(BL114),.BLN(BLN114),.WL(WL117));
sram_cell_6t_5 inst_cell_117_115 (.BL(BL115),.BLN(BLN115),.WL(WL117));
sram_cell_6t_5 inst_cell_117_116 (.BL(BL116),.BLN(BLN116),.WL(WL117));
sram_cell_6t_5 inst_cell_117_117 (.BL(BL117),.BLN(BLN117),.WL(WL117));
sram_cell_6t_5 inst_cell_117_118 (.BL(BL118),.BLN(BLN118),.WL(WL117));
sram_cell_6t_5 inst_cell_117_119 (.BL(BL119),.BLN(BLN119),.WL(WL117));
sram_cell_6t_5 inst_cell_117_120 (.BL(BL120),.BLN(BLN120),.WL(WL117));
sram_cell_6t_5 inst_cell_117_121 (.BL(BL121),.BLN(BLN121),.WL(WL117));
sram_cell_6t_5 inst_cell_117_122 (.BL(BL122),.BLN(BLN122),.WL(WL117));
sram_cell_6t_5 inst_cell_117_123 (.BL(BL123),.BLN(BLN123),.WL(WL117));
sram_cell_6t_5 inst_cell_117_124 (.BL(BL124),.BLN(BLN124),.WL(WL117));
sram_cell_6t_5 inst_cell_117_125 (.BL(BL125),.BLN(BLN125),.WL(WL117));
sram_cell_6t_5 inst_cell_117_126 (.BL(BL126),.BLN(BLN126),.WL(WL117));
sram_cell_6t_5 inst_cell_117_127 (.BL(BL127),.BLN(BLN127),.WL(WL117));
sram_cell_6t_5 inst_cell_118_0 (.BL(BL0),.BLN(BLN0),.WL(WL118));
sram_cell_6t_5 inst_cell_118_1 (.BL(BL1),.BLN(BLN1),.WL(WL118));
sram_cell_6t_5 inst_cell_118_2 (.BL(BL2),.BLN(BLN2),.WL(WL118));
sram_cell_6t_5 inst_cell_118_3 (.BL(BL3),.BLN(BLN3),.WL(WL118));
sram_cell_6t_5 inst_cell_118_4 (.BL(BL4),.BLN(BLN4),.WL(WL118));
sram_cell_6t_5 inst_cell_118_5 (.BL(BL5),.BLN(BLN5),.WL(WL118));
sram_cell_6t_5 inst_cell_118_6 (.BL(BL6),.BLN(BLN6),.WL(WL118));
sram_cell_6t_5 inst_cell_118_7 (.BL(BL7),.BLN(BLN7),.WL(WL118));
sram_cell_6t_5 inst_cell_118_8 (.BL(BL8),.BLN(BLN8),.WL(WL118));
sram_cell_6t_5 inst_cell_118_9 (.BL(BL9),.BLN(BLN9),.WL(WL118));
sram_cell_6t_5 inst_cell_118_10 (.BL(BL10),.BLN(BLN10),.WL(WL118));
sram_cell_6t_5 inst_cell_118_11 (.BL(BL11),.BLN(BLN11),.WL(WL118));
sram_cell_6t_5 inst_cell_118_12 (.BL(BL12),.BLN(BLN12),.WL(WL118));
sram_cell_6t_5 inst_cell_118_13 (.BL(BL13),.BLN(BLN13),.WL(WL118));
sram_cell_6t_5 inst_cell_118_14 (.BL(BL14),.BLN(BLN14),.WL(WL118));
sram_cell_6t_5 inst_cell_118_15 (.BL(BL15),.BLN(BLN15),.WL(WL118));
sram_cell_6t_5 inst_cell_118_16 (.BL(BL16),.BLN(BLN16),.WL(WL118));
sram_cell_6t_5 inst_cell_118_17 (.BL(BL17),.BLN(BLN17),.WL(WL118));
sram_cell_6t_5 inst_cell_118_18 (.BL(BL18),.BLN(BLN18),.WL(WL118));
sram_cell_6t_5 inst_cell_118_19 (.BL(BL19),.BLN(BLN19),.WL(WL118));
sram_cell_6t_5 inst_cell_118_20 (.BL(BL20),.BLN(BLN20),.WL(WL118));
sram_cell_6t_5 inst_cell_118_21 (.BL(BL21),.BLN(BLN21),.WL(WL118));
sram_cell_6t_5 inst_cell_118_22 (.BL(BL22),.BLN(BLN22),.WL(WL118));
sram_cell_6t_5 inst_cell_118_23 (.BL(BL23),.BLN(BLN23),.WL(WL118));
sram_cell_6t_5 inst_cell_118_24 (.BL(BL24),.BLN(BLN24),.WL(WL118));
sram_cell_6t_5 inst_cell_118_25 (.BL(BL25),.BLN(BLN25),.WL(WL118));
sram_cell_6t_5 inst_cell_118_26 (.BL(BL26),.BLN(BLN26),.WL(WL118));
sram_cell_6t_5 inst_cell_118_27 (.BL(BL27),.BLN(BLN27),.WL(WL118));
sram_cell_6t_5 inst_cell_118_28 (.BL(BL28),.BLN(BLN28),.WL(WL118));
sram_cell_6t_5 inst_cell_118_29 (.BL(BL29),.BLN(BLN29),.WL(WL118));
sram_cell_6t_5 inst_cell_118_30 (.BL(BL30),.BLN(BLN30),.WL(WL118));
sram_cell_6t_5 inst_cell_118_31 (.BL(BL31),.BLN(BLN31),.WL(WL118));
sram_cell_6t_5 inst_cell_118_32 (.BL(BL32),.BLN(BLN32),.WL(WL118));
sram_cell_6t_5 inst_cell_118_33 (.BL(BL33),.BLN(BLN33),.WL(WL118));
sram_cell_6t_5 inst_cell_118_34 (.BL(BL34),.BLN(BLN34),.WL(WL118));
sram_cell_6t_5 inst_cell_118_35 (.BL(BL35),.BLN(BLN35),.WL(WL118));
sram_cell_6t_5 inst_cell_118_36 (.BL(BL36),.BLN(BLN36),.WL(WL118));
sram_cell_6t_5 inst_cell_118_37 (.BL(BL37),.BLN(BLN37),.WL(WL118));
sram_cell_6t_5 inst_cell_118_38 (.BL(BL38),.BLN(BLN38),.WL(WL118));
sram_cell_6t_5 inst_cell_118_39 (.BL(BL39),.BLN(BLN39),.WL(WL118));
sram_cell_6t_5 inst_cell_118_40 (.BL(BL40),.BLN(BLN40),.WL(WL118));
sram_cell_6t_5 inst_cell_118_41 (.BL(BL41),.BLN(BLN41),.WL(WL118));
sram_cell_6t_5 inst_cell_118_42 (.BL(BL42),.BLN(BLN42),.WL(WL118));
sram_cell_6t_5 inst_cell_118_43 (.BL(BL43),.BLN(BLN43),.WL(WL118));
sram_cell_6t_5 inst_cell_118_44 (.BL(BL44),.BLN(BLN44),.WL(WL118));
sram_cell_6t_5 inst_cell_118_45 (.BL(BL45),.BLN(BLN45),.WL(WL118));
sram_cell_6t_5 inst_cell_118_46 (.BL(BL46),.BLN(BLN46),.WL(WL118));
sram_cell_6t_5 inst_cell_118_47 (.BL(BL47),.BLN(BLN47),.WL(WL118));
sram_cell_6t_5 inst_cell_118_48 (.BL(BL48),.BLN(BLN48),.WL(WL118));
sram_cell_6t_5 inst_cell_118_49 (.BL(BL49),.BLN(BLN49),.WL(WL118));
sram_cell_6t_5 inst_cell_118_50 (.BL(BL50),.BLN(BLN50),.WL(WL118));
sram_cell_6t_5 inst_cell_118_51 (.BL(BL51),.BLN(BLN51),.WL(WL118));
sram_cell_6t_5 inst_cell_118_52 (.BL(BL52),.BLN(BLN52),.WL(WL118));
sram_cell_6t_5 inst_cell_118_53 (.BL(BL53),.BLN(BLN53),.WL(WL118));
sram_cell_6t_5 inst_cell_118_54 (.BL(BL54),.BLN(BLN54),.WL(WL118));
sram_cell_6t_5 inst_cell_118_55 (.BL(BL55),.BLN(BLN55),.WL(WL118));
sram_cell_6t_5 inst_cell_118_56 (.BL(BL56),.BLN(BLN56),.WL(WL118));
sram_cell_6t_5 inst_cell_118_57 (.BL(BL57),.BLN(BLN57),.WL(WL118));
sram_cell_6t_5 inst_cell_118_58 (.BL(BL58),.BLN(BLN58),.WL(WL118));
sram_cell_6t_5 inst_cell_118_59 (.BL(BL59),.BLN(BLN59),.WL(WL118));
sram_cell_6t_5 inst_cell_118_60 (.BL(BL60),.BLN(BLN60),.WL(WL118));
sram_cell_6t_5 inst_cell_118_61 (.BL(BL61),.BLN(BLN61),.WL(WL118));
sram_cell_6t_5 inst_cell_118_62 (.BL(BL62),.BLN(BLN62),.WL(WL118));
sram_cell_6t_5 inst_cell_118_63 (.BL(BL63),.BLN(BLN63),.WL(WL118));
sram_cell_6t_5 inst_cell_118_64 (.BL(BL64),.BLN(BLN64),.WL(WL118));
sram_cell_6t_5 inst_cell_118_65 (.BL(BL65),.BLN(BLN65),.WL(WL118));
sram_cell_6t_5 inst_cell_118_66 (.BL(BL66),.BLN(BLN66),.WL(WL118));
sram_cell_6t_5 inst_cell_118_67 (.BL(BL67),.BLN(BLN67),.WL(WL118));
sram_cell_6t_5 inst_cell_118_68 (.BL(BL68),.BLN(BLN68),.WL(WL118));
sram_cell_6t_5 inst_cell_118_69 (.BL(BL69),.BLN(BLN69),.WL(WL118));
sram_cell_6t_5 inst_cell_118_70 (.BL(BL70),.BLN(BLN70),.WL(WL118));
sram_cell_6t_5 inst_cell_118_71 (.BL(BL71),.BLN(BLN71),.WL(WL118));
sram_cell_6t_5 inst_cell_118_72 (.BL(BL72),.BLN(BLN72),.WL(WL118));
sram_cell_6t_5 inst_cell_118_73 (.BL(BL73),.BLN(BLN73),.WL(WL118));
sram_cell_6t_5 inst_cell_118_74 (.BL(BL74),.BLN(BLN74),.WL(WL118));
sram_cell_6t_5 inst_cell_118_75 (.BL(BL75),.BLN(BLN75),.WL(WL118));
sram_cell_6t_5 inst_cell_118_76 (.BL(BL76),.BLN(BLN76),.WL(WL118));
sram_cell_6t_5 inst_cell_118_77 (.BL(BL77),.BLN(BLN77),.WL(WL118));
sram_cell_6t_5 inst_cell_118_78 (.BL(BL78),.BLN(BLN78),.WL(WL118));
sram_cell_6t_5 inst_cell_118_79 (.BL(BL79),.BLN(BLN79),.WL(WL118));
sram_cell_6t_5 inst_cell_118_80 (.BL(BL80),.BLN(BLN80),.WL(WL118));
sram_cell_6t_5 inst_cell_118_81 (.BL(BL81),.BLN(BLN81),.WL(WL118));
sram_cell_6t_5 inst_cell_118_82 (.BL(BL82),.BLN(BLN82),.WL(WL118));
sram_cell_6t_5 inst_cell_118_83 (.BL(BL83),.BLN(BLN83),.WL(WL118));
sram_cell_6t_5 inst_cell_118_84 (.BL(BL84),.BLN(BLN84),.WL(WL118));
sram_cell_6t_5 inst_cell_118_85 (.BL(BL85),.BLN(BLN85),.WL(WL118));
sram_cell_6t_5 inst_cell_118_86 (.BL(BL86),.BLN(BLN86),.WL(WL118));
sram_cell_6t_5 inst_cell_118_87 (.BL(BL87),.BLN(BLN87),.WL(WL118));
sram_cell_6t_5 inst_cell_118_88 (.BL(BL88),.BLN(BLN88),.WL(WL118));
sram_cell_6t_5 inst_cell_118_89 (.BL(BL89),.BLN(BLN89),.WL(WL118));
sram_cell_6t_5 inst_cell_118_90 (.BL(BL90),.BLN(BLN90),.WL(WL118));
sram_cell_6t_5 inst_cell_118_91 (.BL(BL91),.BLN(BLN91),.WL(WL118));
sram_cell_6t_5 inst_cell_118_92 (.BL(BL92),.BLN(BLN92),.WL(WL118));
sram_cell_6t_5 inst_cell_118_93 (.BL(BL93),.BLN(BLN93),.WL(WL118));
sram_cell_6t_5 inst_cell_118_94 (.BL(BL94),.BLN(BLN94),.WL(WL118));
sram_cell_6t_5 inst_cell_118_95 (.BL(BL95),.BLN(BLN95),.WL(WL118));
sram_cell_6t_5 inst_cell_118_96 (.BL(BL96),.BLN(BLN96),.WL(WL118));
sram_cell_6t_5 inst_cell_118_97 (.BL(BL97),.BLN(BLN97),.WL(WL118));
sram_cell_6t_5 inst_cell_118_98 (.BL(BL98),.BLN(BLN98),.WL(WL118));
sram_cell_6t_5 inst_cell_118_99 (.BL(BL99),.BLN(BLN99),.WL(WL118));
sram_cell_6t_5 inst_cell_118_100 (.BL(BL100),.BLN(BLN100),.WL(WL118));
sram_cell_6t_5 inst_cell_118_101 (.BL(BL101),.BLN(BLN101),.WL(WL118));
sram_cell_6t_5 inst_cell_118_102 (.BL(BL102),.BLN(BLN102),.WL(WL118));
sram_cell_6t_5 inst_cell_118_103 (.BL(BL103),.BLN(BLN103),.WL(WL118));
sram_cell_6t_5 inst_cell_118_104 (.BL(BL104),.BLN(BLN104),.WL(WL118));
sram_cell_6t_5 inst_cell_118_105 (.BL(BL105),.BLN(BLN105),.WL(WL118));
sram_cell_6t_5 inst_cell_118_106 (.BL(BL106),.BLN(BLN106),.WL(WL118));
sram_cell_6t_5 inst_cell_118_107 (.BL(BL107),.BLN(BLN107),.WL(WL118));
sram_cell_6t_5 inst_cell_118_108 (.BL(BL108),.BLN(BLN108),.WL(WL118));
sram_cell_6t_5 inst_cell_118_109 (.BL(BL109),.BLN(BLN109),.WL(WL118));
sram_cell_6t_5 inst_cell_118_110 (.BL(BL110),.BLN(BLN110),.WL(WL118));
sram_cell_6t_5 inst_cell_118_111 (.BL(BL111),.BLN(BLN111),.WL(WL118));
sram_cell_6t_5 inst_cell_118_112 (.BL(BL112),.BLN(BLN112),.WL(WL118));
sram_cell_6t_5 inst_cell_118_113 (.BL(BL113),.BLN(BLN113),.WL(WL118));
sram_cell_6t_5 inst_cell_118_114 (.BL(BL114),.BLN(BLN114),.WL(WL118));
sram_cell_6t_5 inst_cell_118_115 (.BL(BL115),.BLN(BLN115),.WL(WL118));
sram_cell_6t_5 inst_cell_118_116 (.BL(BL116),.BLN(BLN116),.WL(WL118));
sram_cell_6t_5 inst_cell_118_117 (.BL(BL117),.BLN(BLN117),.WL(WL118));
sram_cell_6t_5 inst_cell_118_118 (.BL(BL118),.BLN(BLN118),.WL(WL118));
sram_cell_6t_5 inst_cell_118_119 (.BL(BL119),.BLN(BLN119),.WL(WL118));
sram_cell_6t_5 inst_cell_118_120 (.BL(BL120),.BLN(BLN120),.WL(WL118));
sram_cell_6t_5 inst_cell_118_121 (.BL(BL121),.BLN(BLN121),.WL(WL118));
sram_cell_6t_5 inst_cell_118_122 (.BL(BL122),.BLN(BLN122),.WL(WL118));
sram_cell_6t_5 inst_cell_118_123 (.BL(BL123),.BLN(BLN123),.WL(WL118));
sram_cell_6t_5 inst_cell_118_124 (.BL(BL124),.BLN(BLN124),.WL(WL118));
sram_cell_6t_5 inst_cell_118_125 (.BL(BL125),.BLN(BLN125),.WL(WL118));
sram_cell_6t_5 inst_cell_118_126 (.BL(BL126),.BLN(BLN126),.WL(WL118));
sram_cell_6t_5 inst_cell_118_127 (.BL(BL127),.BLN(BLN127),.WL(WL118));
sram_cell_6t_5 inst_cell_119_0 (.BL(BL0),.BLN(BLN0),.WL(WL119));
sram_cell_6t_5 inst_cell_119_1 (.BL(BL1),.BLN(BLN1),.WL(WL119));
sram_cell_6t_5 inst_cell_119_2 (.BL(BL2),.BLN(BLN2),.WL(WL119));
sram_cell_6t_5 inst_cell_119_3 (.BL(BL3),.BLN(BLN3),.WL(WL119));
sram_cell_6t_5 inst_cell_119_4 (.BL(BL4),.BLN(BLN4),.WL(WL119));
sram_cell_6t_5 inst_cell_119_5 (.BL(BL5),.BLN(BLN5),.WL(WL119));
sram_cell_6t_5 inst_cell_119_6 (.BL(BL6),.BLN(BLN6),.WL(WL119));
sram_cell_6t_5 inst_cell_119_7 (.BL(BL7),.BLN(BLN7),.WL(WL119));
sram_cell_6t_5 inst_cell_119_8 (.BL(BL8),.BLN(BLN8),.WL(WL119));
sram_cell_6t_5 inst_cell_119_9 (.BL(BL9),.BLN(BLN9),.WL(WL119));
sram_cell_6t_5 inst_cell_119_10 (.BL(BL10),.BLN(BLN10),.WL(WL119));
sram_cell_6t_5 inst_cell_119_11 (.BL(BL11),.BLN(BLN11),.WL(WL119));
sram_cell_6t_5 inst_cell_119_12 (.BL(BL12),.BLN(BLN12),.WL(WL119));
sram_cell_6t_5 inst_cell_119_13 (.BL(BL13),.BLN(BLN13),.WL(WL119));
sram_cell_6t_5 inst_cell_119_14 (.BL(BL14),.BLN(BLN14),.WL(WL119));
sram_cell_6t_5 inst_cell_119_15 (.BL(BL15),.BLN(BLN15),.WL(WL119));
sram_cell_6t_5 inst_cell_119_16 (.BL(BL16),.BLN(BLN16),.WL(WL119));
sram_cell_6t_5 inst_cell_119_17 (.BL(BL17),.BLN(BLN17),.WL(WL119));
sram_cell_6t_5 inst_cell_119_18 (.BL(BL18),.BLN(BLN18),.WL(WL119));
sram_cell_6t_5 inst_cell_119_19 (.BL(BL19),.BLN(BLN19),.WL(WL119));
sram_cell_6t_5 inst_cell_119_20 (.BL(BL20),.BLN(BLN20),.WL(WL119));
sram_cell_6t_5 inst_cell_119_21 (.BL(BL21),.BLN(BLN21),.WL(WL119));
sram_cell_6t_5 inst_cell_119_22 (.BL(BL22),.BLN(BLN22),.WL(WL119));
sram_cell_6t_5 inst_cell_119_23 (.BL(BL23),.BLN(BLN23),.WL(WL119));
sram_cell_6t_5 inst_cell_119_24 (.BL(BL24),.BLN(BLN24),.WL(WL119));
sram_cell_6t_5 inst_cell_119_25 (.BL(BL25),.BLN(BLN25),.WL(WL119));
sram_cell_6t_5 inst_cell_119_26 (.BL(BL26),.BLN(BLN26),.WL(WL119));
sram_cell_6t_5 inst_cell_119_27 (.BL(BL27),.BLN(BLN27),.WL(WL119));
sram_cell_6t_5 inst_cell_119_28 (.BL(BL28),.BLN(BLN28),.WL(WL119));
sram_cell_6t_5 inst_cell_119_29 (.BL(BL29),.BLN(BLN29),.WL(WL119));
sram_cell_6t_5 inst_cell_119_30 (.BL(BL30),.BLN(BLN30),.WL(WL119));
sram_cell_6t_5 inst_cell_119_31 (.BL(BL31),.BLN(BLN31),.WL(WL119));
sram_cell_6t_5 inst_cell_119_32 (.BL(BL32),.BLN(BLN32),.WL(WL119));
sram_cell_6t_5 inst_cell_119_33 (.BL(BL33),.BLN(BLN33),.WL(WL119));
sram_cell_6t_5 inst_cell_119_34 (.BL(BL34),.BLN(BLN34),.WL(WL119));
sram_cell_6t_5 inst_cell_119_35 (.BL(BL35),.BLN(BLN35),.WL(WL119));
sram_cell_6t_5 inst_cell_119_36 (.BL(BL36),.BLN(BLN36),.WL(WL119));
sram_cell_6t_5 inst_cell_119_37 (.BL(BL37),.BLN(BLN37),.WL(WL119));
sram_cell_6t_5 inst_cell_119_38 (.BL(BL38),.BLN(BLN38),.WL(WL119));
sram_cell_6t_5 inst_cell_119_39 (.BL(BL39),.BLN(BLN39),.WL(WL119));
sram_cell_6t_5 inst_cell_119_40 (.BL(BL40),.BLN(BLN40),.WL(WL119));
sram_cell_6t_5 inst_cell_119_41 (.BL(BL41),.BLN(BLN41),.WL(WL119));
sram_cell_6t_5 inst_cell_119_42 (.BL(BL42),.BLN(BLN42),.WL(WL119));
sram_cell_6t_5 inst_cell_119_43 (.BL(BL43),.BLN(BLN43),.WL(WL119));
sram_cell_6t_5 inst_cell_119_44 (.BL(BL44),.BLN(BLN44),.WL(WL119));
sram_cell_6t_5 inst_cell_119_45 (.BL(BL45),.BLN(BLN45),.WL(WL119));
sram_cell_6t_5 inst_cell_119_46 (.BL(BL46),.BLN(BLN46),.WL(WL119));
sram_cell_6t_5 inst_cell_119_47 (.BL(BL47),.BLN(BLN47),.WL(WL119));
sram_cell_6t_5 inst_cell_119_48 (.BL(BL48),.BLN(BLN48),.WL(WL119));
sram_cell_6t_5 inst_cell_119_49 (.BL(BL49),.BLN(BLN49),.WL(WL119));
sram_cell_6t_5 inst_cell_119_50 (.BL(BL50),.BLN(BLN50),.WL(WL119));
sram_cell_6t_5 inst_cell_119_51 (.BL(BL51),.BLN(BLN51),.WL(WL119));
sram_cell_6t_5 inst_cell_119_52 (.BL(BL52),.BLN(BLN52),.WL(WL119));
sram_cell_6t_5 inst_cell_119_53 (.BL(BL53),.BLN(BLN53),.WL(WL119));
sram_cell_6t_5 inst_cell_119_54 (.BL(BL54),.BLN(BLN54),.WL(WL119));
sram_cell_6t_5 inst_cell_119_55 (.BL(BL55),.BLN(BLN55),.WL(WL119));
sram_cell_6t_5 inst_cell_119_56 (.BL(BL56),.BLN(BLN56),.WL(WL119));
sram_cell_6t_5 inst_cell_119_57 (.BL(BL57),.BLN(BLN57),.WL(WL119));
sram_cell_6t_5 inst_cell_119_58 (.BL(BL58),.BLN(BLN58),.WL(WL119));
sram_cell_6t_5 inst_cell_119_59 (.BL(BL59),.BLN(BLN59),.WL(WL119));
sram_cell_6t_5 inst_cell_119_60 (.BL(BL60),.BLN(BLN60),.WL(WL119));
sram_cell_6t_5 inst_cell_119_61 (.BL(BL61),.BLN(BLN61),.WL(WL119));
sram_cell_6t_5 inst_cell_119_62 (.BL(BL62),.BLN(BLN62),.WL(WL119));
sram_cell_6t_5 inst_cell_119_63 (.BL(BL63),.BLN(BLN63),.WL(WL119));
sram_cell_6t_5 inst_cell_119_64 (.BL(BL64),.BLN(BLN64),.WL(WL119));
sram_cell_6t_5 inst_cell_119_65 (.BL(BL65),.BLN(BLN65),.WL(WL119));
sram_cell_6t_5 inst_cell_119_66 (.BL(BL66),.BLN(BLN66),.WL(WL119));
sram_cell_6t_5 inst_cell_119_67 (.BL(BL67),.BLN(BLN67),.WL(WL119));
sram_cell_6t_5 inst_cell_119_68 (.BL(BL68),.BLN(BLN68),.WL(WL119));
sram_cell_6t_5 inst_cell_119_69 (.BL(BL69),.BLN(BLN69),.WL(WL119));
sram_cell_6t_5 inst_cell_119_70 (.BL(BL70),.BLN(BLN70),.WL(WL119));
sram_cell_6t_5 inst_cell_119_71 (.BL(BL71),.BLN(BLN71),.WL(WL119));
sram_cell_6t_5 inst_cell_119_72 (.BL(BL72),.BLN(BLN72),.WL(WL119));
sram_cell_6t_5 inst_cell_119_73 (.BL(BL73),.BLN(BLN73),.WL(WL119));
sram_cell_6t_5 inst_cell_119_74 (.BL(BL74),.BLN(BLN74),.WL(WL119));
sram_cell_6t_5 inst_cell_119_75 (.BL(BL75),.BLN(BLN75),.WL(WL119));
sram_cell_6t_5 inst_cell_119_76 (.BL(BL76),.BLN(BLN76),.WL(WL119));
sram_cell_6t_5 inst_cell_119_77 (.BL(BL77),.BLN(BLN77),.WL(WL119));
sram_cell_6t_5 inst_cell_119_78 (.BL(BL78),.BLN(BLN78),.WL(WL119));
sram_cell_6t_5 inst_cell_119_79 (.BL(BL79),.BLN(BLN79),.WL(WL119));
sram_cell_6t_5 inst_cell_119_80 (.BL(BL80),.BLN(BLN80),.WL(WL119));
sram_cell_6t_5 inst_cell_119_81 (.BL(BL81),.BLN(BLN81),.WL(WL119));
sram_cell_6t_5 inst_cell_119_82 (.BL(BL82),.BLN(BLN82),.WL(WL119));
sram_cell_6t_5 inst_cell_119_83 (.BL(BL83),.BLN(BLN83),.WL(WL119));
sram_cell_6t_5 inst_cell_119_84 (.BL(BL84),.BLN(BLN84),.WL(WL119));
sram_cell_6t_5 inst_cell_119_85 (.BL(BL85),.BLN(BLN85),.WL(WL119));
sram_cell_6t_5 inst_cell_119_86 (.BL(BL86),.BLN(BLN86),.WL(WL119));
sram_cell_6t_5 inst_cell_119_87 (.BL(BL87),.BLN(BLN87),.WL(WL119));
sram_cell_6t_5 inst_cell_119_88 (.BL(BL88),.BLN(BLN88),.WL(WL119));
sram_cell_6t_5 inst_cell_119_89 (.BL(BL89),.BLN(BLN89),.WL(WL119));
sram_cell_6t_5 inst_cell_119_90 (.BL(BL90),.BLN(BLN90),.WL(WL119));
sram_cell_6t_5 inst_cell_119_91 (.BL(BL91),.BLN(BLN91),.WL(WL119));
sram_cell_6t_5 inst_cell_119_92 (.BL(BL92),.BLN(BLN92),.WL(WL119));
sram_cell_6t_5 inst_cell_119_93 (.BL(BL93),.BLN(BLN93),.WL(WL119));
sram_cell_6t_5 inst_cell_119_94 (.BL(BL94),.BLN(BLN94),.WL(WL119));
sram_cell_6t_5 inst_cell_119_95 (.BL(BL95),.BLN(BLN95),.WL(WL119));
sram_cell_6t_5 inst_cell_119_96 (.BL(BL96),.BLN(BLN96),.WL(WL119));
sram_cell_6t_5 inst_cell_119_97 (.BL(BL97),.BLN(BLN97),.WL(WL119));
sram_cell_6t_5 inst_cell_119_98 (.BL(BL98),.BLN(BLN98),.WL(WL119));
sram_cell_6t_5 inst_cell_119_99 (.BL(BL99),.BLN(BLN99),.WL(WL119));
sram_cell_6t_5 inst_cell_119_100 (.BL(BL100),.BLN(BLN100),.WL(WL119));
sram_cell_6t_5 inst_cell_119_101 (.BL(BL101),.BLN(BLN101),.WL(WL119));
sram_cell_6t_5 inst_cell_119_102 (.BL(BL102),.BLN(BLN102),.WL(WL119));
sram_cell_6t_5 inst_cell_119_103 (.BL(BL103),.BLN(BLN103),.WL(WL119));
sram_cell_6t_5 inst_cell_119_104 (.BL(BL104),.BLN(BLN104),.WL(WL119));
sram_cell_6t_5 inst_cell_119_105 (.BL(BL105),.BLN(BLN105),.WL(WL119));
sram_cell_6t_5 inst_cell_119_106 (.BL(BL106),.BLN(BLN106),.WL(WL119));
sram_cell_6t_5 inst_cell_119_107 (.BL(BL107),.BLN(BLN107),.WL(WL119));
sram_cell_6t_5 inst_cell_119_108 (.BL(BL108),.BLN(BLN108),.WL(WL119));
sram_cell_6t_5 inst_cell_119_109 (.BL(BL109),.BLN(BLN109),.WL(WL119));
sram_cell_6t_5 inst_cell_119_110 (.BL(BL110),.BLN(BLN110),.WL(WL119));
sram_cell_6t_5 inst_cell_119_111 (.BL(BL111),.BLN(BLN111),.WL(WL119));
sram_cell_6t_5 inst_cell_119_112 (.BL(BL112),.BLN(BLN112),.WL(WL119));
sram_cell_6t_5 inst_cell_119_113 (.BL(BL113),.BLN(BLN113),.WL(WL119));
sram_cell_6t_5 inst_cell_119_114 (.BL(BL114),.BLN(BLN114),.WL(WL119));
sram_cell_6t_5 inst_cell_119_115 (.BL(BL115),.BLN(BLN115),.WL(WL119));
sram_cell_6t_5 inst_cell_119_116 (.BL(BL116),.BLN(BLN116),.WL(WL119));
sram_cell_6t_5 inst_cell_119_117 (.BL(BL117),.BLN(BLN117),.WL(WL119));
sram_cell_6t_5 inst_cell_119_118 (.BL(BL118),.BLN(BLN118),.WL(WL119));
sram_cell_6t_5 inst_cell_119_119 (.BL(BL119),.BLN(BLN119),.WL(WL119));
sram_cell_6t_5 inst_cell_119_120 (.BL(BL120),.BLN(BLN120),.WL(WL119));
sram_cell_6t_5 inst_cell_119_121 (.BL(BL121),.BLN(BLN121),.WL(WL119));
sram_cell_6t_5 inst_cell_119_122 (.BL(BL122),.BLN(BLN122),.WL(WL119));
sram_cell_6t_5 inst_cell_119_123 (.BL(BL123),.BLN(BLN123),.WL(WL119));
sram_cell_6t_5 inst_cell_119_124 (.BL(BL124),.BLN(BLN124),.WL(WL119));
sram_cell_6t_5 inst_cell_119_125 (.BL(BL125),.BLN(BLN125),.WL(WL119));
sram_cell_6t_5 inst_cell_119_126 (.BL(BL126),.BLN(BLN126),.WL(WL119));
sram_cell_6t_5 inst_cell_119_127 (.BL(BL127),.BLN(BLN127),.WL(WL119));
sram_cell_6t_5 inst_cell_120_0 (.BL(BL0),.BLN(BLN0),.WL(WL120));
sram_cell_6t_5 inst_cell_120_1 (.BL(BL1),.BLN(BLN1),.WL(WL120));
sram_cell_6t_5 inst_cell_120_2 (.BL(BL2),.BLN(BLN2),.WL(WL120));
sram_cell_6t_5 inst_cell_120_3 (.BL(BL3),.BLN(BLN3),.WL(WL120));
sram_cell_6t_5 inst_cell_120_4 (.BL(BL4),.BLN(BLN4),.WL(WL120));
sram_cell_6t_5 inst_cell_120_5 (.BL(BL5),.BLN(BLN5),.WL(WL120));
sram_cell_6t_5 inst_cell_120_6 (.BL(BL6),.BLN(BLN6),.WL(WL120));
sram_cell_6t_5 inst_cell_120_7 (.BL(BL7),.BLN(BLN7),.WL(WL120));
sram_cell_6t_5 inst_cell_120_8 (.BL(BL8),.BLN(BLN8),.WL(WL120));
sram_cell_6t_5 inst_cell_120_9 (.BL(BL9),.BLN(BLN9),.WL(WL120));
sram_cell_6t_5 inst_cell_120_10 (.BL(BL10),.BLN(BLN10),.WL(WL120));
sram_cell_6t_5 inst_cell_120_11 (.BL(BL11),.BLN(BLN11),.WL(WL120));
sram_cell_6t_5 inst_cell_120_12 (.BL(BL12),.BLN(BLN12),.WL(WL120));
sram_cell_6t_5 inst_cell_120_13 (.BL(BL13),.BLN(BLN13),.WL(WL120));
sram_cell_6t_5 inst_cell_120_14 (.BL(BL14),.BLN(BLN14),.WL(WL120));
sram_cell_6t_5 inst_cell_120_15 (.BL(BL15),.BLN(BLN15),.WL(WL120));
sram_cell_6t_5 inst_cell_120_16 (.BL(BL16),.BLN(BLN16),.WL(WL120));
sram_cell_6t_5 inst_cell_120_17 (.BL(BL17),.BLN(BLN17),.WL(WL120));
sram_cell_6t_5 inst_cell_120_18 (.BL(BL18),.BLN(BLN18),.WL(WL120));
sram_cell_6t_5 inst_cell_120_19 (.BL(BL19),.BLN(BLN19),.WL(WL120));
sram_cell_6t_5 inst_cell_120_20 (.BL(BL20),.BLN(BLN20),.WL(WL120));
sram_cell_6t_5 inst_cell_120_21 (.BL(BL21),.BLN(BLN21),.WL(WL120));
sram_cell_6t_5 inst_cell_120_22 (.BL(BL22),.BLN(BLN22),.WL(WL120));
sram_cell_6t_5 inst_cell_120_23 (.BL(BL23),.BLN(BLN23),.WL(WL120));
sram_cell_6t_5 inst_cell_120_24 (.BL(BL24),.BLN(BLN24),.WL(WL120));
sram_cell_6t_5 inst_cell_120_25 (.BL(BL25),.BLN(BLN25),.WL(WL120));
sram_cell_6t_5 inst_cell_120_26 (.BL(BL26),.BLN(BLN26),.WL(WL120));
sram_cell_6t_5 inst_cell_120_27 (.BL(BL27),.BLN(BLN27),.WL(WL120));
sram_cell_6t_5 inst_cell_120_28 (.BL(BL28),.BLN(BLN28),.WL(WL120));
sram_cell_6t_5 inst_cell_120_29 (.BL(BL29),.BLN(BLN29),.WL(WL120));
sram_cell_6t_5 inst_cell_120_30 (.BL(BL30),.BLN(BLN30),.WL(WL120));
sram_cell_6t_5 inst_cell_120_31 (.BL(BL31),.BLN(BLN31),.WL(WL120));
sram_cell_6t_5 inst_cell_120_32 (.BL(BL32),.BLN(BLN32),.WL(WL120));
sram_cell_6t_5 inst_cell_120_33 (.BL(BL33),.BLN(BLN33),.WL(WL120));
sram_cell_6t_5 inst_cell_120_34 (.BL(BL34),.BLN(BLN34),.WL(WL120));
sram_cell_6t_5 inst_cell_120_35 (.BL(BL35),.BLN(BLN35),.WL(WL120));
sram_cell_6t_5 inst_cell_120_36 (.BL(BL36),.BLN(BLN36),.WL(WL120));
sram_cell_6t_5 inst_cell_120_37 (.BL(BL37),.BLN(BLN37),.WL(WL120));
sram_cell_6t_5 inst_cell_120_38 (.BL(BL38),.BLN(BLN38),.WL(WL120));
sram_cell_6t_5 inst_cell_120_39 (.BL(BL39),.BLN(BLN39),.WL(WL120));
sram_cell_6t_5 inst_cell_120_40 (.BL(BL40),.BLN(BLN40),.WL(WL120));
sram_cell_6t_5 inst_cell_120_41 (.BL(BL41),.BLN(BLN41),.WL(WL120));
sram_cell_6t_5 inst_cell_120_42 (.BL(BL42),.BLN(BLN42),.WL(WL120));
sram_cell_6t_5 inst_cell_120_43 (.BL(BL43),.BLN(BLN43),.WL(WL120));
sram_cell_6t_5 inst_cell_120_44 (.BL(BL44),.BLN(BLN44),.WL(WL120));
sram_cell_6t_5 inst_cell_120_45 (.BL(BL45),.BLN(BLN45),.WL(WL120));
sram_cell_6t_5 inst_cell_120_46 (.BL(BL46),.BLN(BLN46),.WL(WL120));
sram_cell_6t_5 inst_cell_120_47 (.BL(BL47),.BLN(BLN47),.WL(WL120));
sram_cell_6t_5 inst_cell_120_48 (.BL(BL48),.BLN(BLN48),.WL(WL120));
sram_cell_6t_5 inst_cell_120_49 (.BL(BL49),.BLN(BLN49),.WL(WL120));
sram_cell_6t_5 inst_cell_120_50 (.BL(BL50),.BLN(BLN50),.WL(WL120));
sram_cell_6t_5 inst_cell_120_51 (.BL(BL51),.BLN(BLN51),.WL(WL120));
sram_cell_6t_5 inst_cell_120_52 (.BL(BL52),.BLN(BLN52),.WL(WL120));
sram_cell_6t_5 inst_cell_120_53 (.BL(BL53),.BLN(BLN53),.WL(WL120));
sram_cell_6t_5 inst_cell_120_54 (.BL(BL54),.BLN(BLN54),.WL(WL120));
sram_cell_6t_5 inst_cell_120_55 (.BL(BL55),.BLN(BLN55),.WL(WL120));
sram_cell_6t_5 inst_cell_120_56 (.BL(BL56),.BLN(BLN56),.WL(WL120));
sram_cell_6t_5 inst_cell_120_57 (.BL(BL57),.BLN(BLN57),.WL(WL120));
sram_cell_6t_5 inst_cell_120_58 (.BL(BL58),.BLN(BLN58),.WL(WL120));
sram_cell_6t_5 inst_cell_120_59 (.BL(BL59),.BLN(BLN59),.WL(WL120));
sram_cell_6t_5 inst_cell_120_60 (.BL(BL60),.BLN(BLN60),.WL(WL120));
sram_cell_6t_5 inst_cell_120_61 (.BL(BL61),.BLN(BLN61),.WL(WL120));
sram_cell_6t_5 inst_cell_120_62 (.BL(BL62),.BLN(BLN62),.WL(WL120));
sram_cell_6t_5 inst_cell_120_63 (.BL(BL63),.BLN(BLN63),.WL(WL120));
sram_cell_6t_5 inst_cell_120_64 (.BL(BL64),.BLN(BLN64),.WL(WL120));
sram_cell_6t_5 inst_cell_120_65 (.BL(BL65),.BLN(BLN65),.WL(WL120));
sram_cell_6t_5 inst_cell_120_66 (.BL(BL66),.BLN(BLN66),.WL(WL120));
sram_cell_6t_5 inst_cell_120_67 (.BL(BL67),.BLN(BLN67),.WL(WL120));
sram_cell_6t_5 inst_cell_120_68 (.BL(BL68),.BLN(BLN68),.WL(WL120));
sram_cell_6t_5 inst_cell_120_69 (.BL(BL69),.BLN(BLN69),.WL(WL120));
sram_cell_6t_5 inst_cell_120_70 (.BL(BL70),.BLN(BLN70),.WL(WL120));
sram_cell_6t_5 inst_cell_120_71 (.BL(BL71),.BLN(BLN71),.WL(WL120));
sram_cell_6t_5 inst_cell_120_72 (.BL(BL72),.BLN(BLN72),.WL(WL120));
sram_cell_6t_5 inst_cell_120_73 (.BL(BL73),.BLN(BLN73),.WL(WL120));
sram_cell_6t_5 inst_cell_120_74 (.BL(BL74),.BLN(BLN74),.WL(WL120));
sram_cell_6t_5 inst_cell_120_75 (.BL(BL75),.BLN(BLN75),.WL(WL120));
sram_cell_6t_5 inst_cell_120_76 (.BL(BL76),.BLN(BLN76),.WL(WL120));
sram_cell_6t_5 inst_cell_120_77 (.BL(BL77),.BLN(BLN77),.WL(WL120));
sram_cell_6t_5 inst_cell_120_78 (.BL(BL78),.BLN(BLN78),.WL(WL120));
sram_cell_6t_5 inst_cell_120_79 (.BL(BL79),.BLN(BLN79),.WL(WL120));
sram_cell_6t_5 inst_cell_120_80 (.BL(BL80),.BLN(BLN80),.WL(WL120));
sram_cell_6t_5 inst_cell_120_81 (.BL(BL81),.BLN(BLN81),.WL(WL120));
sram_cell_6t_5 inst_cell_120_82 (.BL(BL82),.BLN(BLN82),.WL(WL120));
sram_cell_6t_5 inst_cell_120_83 (.BL(BL83),.BLN(BLN83),.WL(WL120));
sram_cell_6t_5 inst_cell_120_84 (.BL(BL84),.BLN(BLN84),.WL(WL120));
sram_cell_6t_5 inst_cell_120_85 (.BL(BL85),.BLN(BLN85),.WL(WL120));
sram_cell_6t_5 inst_cell_120_86 (.BL(BL86),.BLN(BLN86),.WL(WL120));
sram_cell_6t_5 inst_cell_120_87 (.BL(BL87),.BLN(BLN87),.WL(WL120));
sram_cell_6t_5 inst_cell_120_88 (.BL(BL88),.BLN(BLN88),.WL(WL120));
sram_cell_6t_5 inst_cell_120_89 (.BL(BL89),.BLN(BLN89),.WL(WL120));
sram_cell_6t_5 inst_cell_120_90 (.BL(BL90),.BLN(BLN90),.WL(WL120));
sram_cell_6t_5 inst_cell_120_91 (.BL(BL91),.BLN(BLN91),.WL(WL120));
sram_cell_6t_5 inst_cell_120_92 (.BL(BL92),.BLN(BLN92),.WL(WL120));
sram_cell_6t_5 inst_cell_120_93 (.BL(BL93),.BLN(BLN93),.WL(WL120));
sram_cell_6t_5 inst_cell_120_94 (.BL(BL94),.BLN(BLN94),.WL(WL120));
sram_cell_6t_5 inst_cell_120_95 (.BL(BL95),.BLN(BLN95),.WL(WL120));
sram_cell_6t_5 inst_cell_120_96 (.BL(BL96),.BLN(BLN96),.WL(WL120));
sram_cell_6t_5 inst_cell_120_97 (.BL(BL97),.BLN(BLN97),.WL(WL120));
sram_cell_6t_5 inst_cell_120_98 (.BL(BL98),.BLN(BLN98),.WL(WL120));
sram_cell_6t_5 inst_cell_120_99 (.BL(BL99),.BLN(BLN99),.WL(WL120));
sram_cell_6t_5 inst_cell_120_100 (.BL(BL100),.BLN(BLN100),.WL(WL120));
sram_cell_6t_5 inst_cell_120_101 (.BL(BL101),.BLN(BLN101),.WL(WL120));
sram_cell_6t_5 inst_cell_120_102 (.BL(BL102),.BLN(BLN102),.WL(WL120));
sram_cell_6t_5 inst_cell_120_103 (.BL(BL103),.BLN(BLN103),.WL(WL120));
sram_cell_6t_5 inst_cell_120_104 (.BL(BL104),.BLN(BLN104),.WL(WL120));
sram_cell_6t_5 inst_cell_120_105 (.BL(BL105),.BLN(BLN105),.WL(WL120));
sram_cell_6t_5 inst_cell_120_106 (.BL(BL106),.BLN(BLN106),.WL(WL120));
sram_cell_6t_5 inst_cell_120_107 (.BL(BL107),.BLN(BLN107),.WL(WL120));
sram_cell_6t_5 inst_cell_120_108 (.BL(BL108),.BLN(BLN108),.WL(WL120));
sram_cell_6t_5 inst_cell_120_109 (.BL(BL109),.BLN(BLN109),.WL(WL120));
sram_cell_6t_5 inst_cell_120_110 (.BL(BL110),.BLN(BLN110),.WL(WL120));
sram_cell_6t_5 inst_cell_120_111 (.BL(BL111),.BLN(BLN111),.WL(WL120));
sram_cell_6t_5 inst_cell_120_112 (.BL(BL112),.BLN(BLN112),.WL(WL120));
sram_cell_6t_5 inst_cell_120_113 (.BL(BL113),.BLN(BLN113),.WL(WL120));
sram_cell_6t_5 inst_cell_120_114 (.BL(BL114),.BLN(BLN114),.WL(WL120));
sram_cell_6t_5 inst_cell_120_115 (.BL(BL115),.BLN(BLN115),.WL(WL120));
sram_cell_6t_5 inst_cell_120_116 (.BL(BL116),.BLN(BLN116),.WL(WL120));
sram_cell_6t_5 inst_cell_120_117 (.BL(BL117),.BLN(BLN117),.WL(WL120));
sram_cell_6t_5 inst_cell_120_118 (.BL(BL118),.BLN(BLN118),.WL(WL120));
sram_cell_6t_5 inst_cell_120_119 (.BL(BL119),.BLN(BLN119),.WL(WL120));
sram_cell_6t_5 inst_cell_120_120 (.BL(BL120),.BLN(BLN120),.WL(WL120));
sram_cell_6t_5 inst_cell_120_121 (.BL(BL121),.BLN(BLN121),.WL(WL120));
sram_cell_6t_5 inst_cell_120_122 (.BL(BL122),.BLN(BLN122),.WL(WL120));
sram_cell_6t_5 inst_cell_120_123 (.BL(BL123),.BLN(BLN123),.WL(WL120));
sram_cell_6t_5 inst_cell_120_124 (.BL(BL124),.BLN(BLN124),.WL(WL120));
sram_cell_6t_5 inst_cell_120_125 (.BL(BL125),.BLN(BLN125),.WL(WL120));
sram_cell_6t_5 inst_cell_120_126 (.BL(BL126),.BLN(BLN126),.WL(WL120));
sram_cell_6t_5 inst_cell_120_127 (.BL(BL127),.BLN(BLN127),.WL(WL120));
sram_cell_6t_5 inst_cell_121_0 (.BL(BL0),.BLN(BLN0),.WL(WL121));
sram_cell_6t_5 inst_cell_121_1 (.BL(BL1),.BLN(BLN1),.WL(WL121));
sram_cell_6t_5 inst_cell_121_2 (.BL(BL2),.BLN(BLN2),.WL(WL121));
sram_cell_6t_5 inst_cell_121_3 (.BL(BL3),.BLN(BLN3),.WL(WL121));
sram_cell_6t_5 inst_cell_121_4 (.BL(BL4),.BLN(BLN4),.WL(WL121));
sram_cell_6t_5 inst_cell_121_5 (.BL(BL5),.BLN(BLN5),.WL(WL121));
sram_cell_6t_5 inst_cell_121_6 (.BL(BL6),.BLN(BLN6),.WL(WL121));
sram_cell_6t_5 inst_cell_121_7 (.BL(BL7),.BLN(BLN7),.WL(WL121));
sram_cell_6t_5 inst_cell_121_8 (.BL(BL8),.BLN(BLN8),.WL(WL121));
sram_cell_6t_5 inst_cell_121_9 (.BL(BL9),.BLN(BLN9),.WL(WL121));
sram_cell_6t_5 inst_cell_121_10 (.BL(BL10),.BLN(BLN10),.WL(WL121));
sram_cell_6t_5 inst_cell_121_11 (.BL(BL11),.BLN(BLN11),.WL(WL121));
sram_cell_6t_5 inst_cell_121_12 (.BL(BL12),.BLN(BLN12),.WL(WL121));
sram_cell_6t_5 inst_cell_121_13 (.BL(BL13),.BLN(BLN13),.WL(WL121));
sram_cell_6t_5 inst_cell_121_14 (.BL(BL14),.BLN(BLN14),.WL(WL121));
sram_cell_6t_5 inst_cell_121_15 (.BL(BL15),.BLN(BLN15),.WL(WL121));
sram_cell_6t_5 inst_cell_121_16 (.BL(BL16),.BLN(BLN16),.WL(WL121));
sram_cell_6t_5 inst_cell_121_17 (.BL(BL17),.BLN(BLN17),.WL(WL121));
sram_cell_6t_5 inst_cell_121_18 (.BL(BL18),.BLN(BLN18),.WL(WL121));
sram_cell_6t_5 inst_cell_121_19 (.BL(BL19),.BLN(BLN19),.WL(WL121));
sram_cell_6t_5 inst_cell_121_20 (.BL(BL20),.BLN(BLN20),.WL(WL121));
sram_cell_6t_5 inst_cell_121_21 (.BL(BL21),.BLN(BLN21),.WL(WL121));
sram_cell_6t_5 inst_cell_121_22 (.BL(BL22),.BLN(BLN22),.WL(WL121));
sram_cell_6t_5 inst_cell_121_23 (.BL(BL23),.BLN(BLN23),.WL(WL121));
sram_cell_6t_5 inst_cell_121_24 (.BL(BL24),.BLN(BLN24),.WL(WL121));
sram_cell_6t_5 inst_cell_121_25 (.BL(BL25),.BLN(BLN25),.WL(WL121));
sram_cell_6t_5 inst_cell_121_26 (.BL(BL26),.BLN(BLN26),.WL(WL121));
sram_cell_6t_5 inst_cell_121_27 (.BL(BL27),.BLN(BLN27),.WL(WL121));
sram_cell_6t_5 inst_cell_121_28 (.BL(BL28),.BLN(BLN28),.WL(WL121));
sram_cell_6t_5 inst_cell_121_29 (.BL(BL29),.BLN(BLN29),.WL(WL121));
sram_cell_6t_5 inst_cell_121_30 (.BL(BL30),.BLN(BLN30),.WL(WL121));
sram_cell_6t_5 inst_cell_121_31 (.BL(BL31),.BLN(BLN31),.WL(WL121));
sram_cell_6t_5 inst_cell_121_32 (.BL(BL32),.BLN(BLN32),.WL(WL121));
sram_cell_6t_5 inst_cell_121_33 (.BL(BL33),.BLN(BLN33),.WL(WL121));
sram_cell_6t_5 inst_cell_121_34 (.BL(BL34),.BLN(BLN34),.WL(WL121));
sram_cell_6t_5 inst_cell_121_35 (.BL(BL35),.BLN(BLN35),.WL(WL121));
sram_cell_6t_5 inst_cell_121_36 (.BL(BL36),.BLN(BLN36),.WL(WL121));
sram_cell_6t_5 inst_cell_121_37 (.BL(BL37),.BLN(BLN37),.WL(WL121));
sram_cell_6t_5 inst_cell_121_38 (.BL(BL38),.BLN(BLN38),.WL(WL121));
sram_cell_6t_5 inst_cell_121_39 (.BL(BL39),.BLN(BLN39),.WL(WL121));
sram_cell_6t_5 inst_cell_121_40 (.BL(BL40),.BLN(BLN40),.WL(WL121));
sram_cell_6t_5 inst_cell_121_41 (.BL(BL41),.BLN(BLN41),.WL(WL121));
sram_cell_6t_5 inst_cell_121_42 (.BL(BL42),.BLN(BLN42),.WL(WL121));
sram_cell_6t_5 inst_cell_121_43 (.BL(BL43),.BLN(BLN43),.WL(WL121));
sram_cell_6t_5 inst_cell_121_44 (.BL(BL44),.BLN(BLN44),.WL(WL121));
sram_cell_6t_5 inst_cell_121_45 (.BL(BL45),.BLN(BLN45),.WL(WL121));
sram_cell_6t_5 inst_cell_121_46 (.BL(BL46),.BLN(BLN46),.WL(WL121));
sram_cell_6t_5 inst_cell_121_47 (.BL(BL47),.BLN(BLN47),.WL(WL121));
sram_cell_6t_5 inst_cell_121_48 (.BL(BL48),.BLN(BLN48),.WL(WL121));
sram_cell_6t_5 inst_cell_121_49 (.BL(BL49),.BLN(BLN49),.WL(WL121));
sram_cell_6t_5 inst_cell_121_50 (.BL(BL50),.BLN(BLN50),.WL(WL121));
sram_cell_6t_5 inst_cell_121_51 (.BL(BL51),.BLN(BLN51),.WL(WL121));
sram_cell_6t_5 inst_cell_121_52 (.BL(BL52),.BLN(BLN52),.WL(WL121));
sram_cell_6t_5 inst_cell_121_53 (.BL(BL53),.BLN(BLN53),.WL(WL121));
sram_cell_6t_5 inst_cell_121_54 (.BL(BL54),.BLN(BLN54),.WL(WL121));
sram_cell_6t_5 inst_cell_121_55 (.BL(BL55),.BLN(BLN55),.WL(WL121));
sram_cell_6t_5 inst_cell_121_56 (.BL(BL56),.BLN(BLN56),.WL(WL121));
sram_cell_6t_5 inst_cell_121_57 (.BL(BL57),.BLN(BLN57),.WL(WL121));
sram_cell_6t_5 inst_cell_121_58 (.BL(BL58),.BLN(BLN58),.WL(WL121));
sram_cell_6t_5 inst_cell_121_59 (.BL(BL59),.BLN(BLN59),.WL(WL121));
sram_cell_6t_5 inst_cell_121_60 (.BL(BL60),.BLN(BLN60),.WL(WL121));
sram_cell_6t_5 inst_cell_121_61 (.BL(BL61),.BLN(BLN61),.WL(WL121));
sram_cell_6t_5 inst_cell_121_62 (.BL(BL62),.BLN(BLN62),.WL(WL121));
sram_cell_6t_5 inst_cell_121_63 (.BL(BL63),.BLN(BLN63),.WL(WL121));
sram_cell_6t_5 inst_cell_121_64 (.BL(BL64),.BLN(BLN64),.WL(WL121));
sram_cell_6t_5 inst_cell_121_65 (.BL(BL65),.BLN(BLN65),.WL(WL121));
sram_cell_6t_5 inst_cell_121_66 (.BL(BL66),.BLN(BLN66),.WL(WL121));
sram_cell_6t_5 inst_cell_121_67 (.BL(BL67),.BLN(BLN67),.WL(WL121));
sram_cell_6t_5 inst_cell_121_68 (.BL(BL68),.BLN(BLN68),.WL(WL121));
sram_cell_6t_5 inst_cell_121_69 (.BL(BL69),.BLN(BLN69),.WL(WL121));
sram_cell_6t_5 inst_cell_121_70 (.BL(BL70),.BLN(BLN70),.WL(WL121));
sram_cell_6t_5 inst_cell_121_71 (.BL(BL71),.BLN(BLN71),.WL(WL121));
sram_cell_6t_5 inst_cell_121_72 (.BL(BL72),.BLN(BLN72),.WL(WL121));
sram_cell_6t_5 inst_cell_121_73 (.BL(BL73),.BLN(BLN73),.WL(WL121));
sram_cell_6t_5 inst_cell_121_74 (.BL(BL74),.BLN(BLN74),.WL(WL121));
sram_cell_6t_5 inst_cell_121_75 (.BL(BL75),.BLN(BLN75),.WL(WL121));
sram_cell_6t_5 inst_cell_121_76 (.BL(BL76),.BLN(BLN76),.WL(WL121));
sram_cell_6t_5 inst_cell_121_77 (.BL(BL77),.BLN(BLN77),.WL(WL121));
sram_cell_6t_5 inst_cell_121_78 (.BL(BL78),.BLN(BLN78),.WL(WL121));
sram_cell_6t_5 inst_cell_121_79 (.BL(BL79),.BLN(BLN79),.WL(WL121));
sram_cell_6t_5 inst_cell_121_80 (.BL(BL80),.BLN(BLN80),.WL(WL121));
sram_cell_6t_5 inst_cell_121_81 (.BL(BL81),.BLN(BLN81),.WL(WL121));
sram_cell_6t_5 inst_cell_121_82 (.BL(BL82),.BLN(BLN82),.WL(WL121));
sram_cell_6t_5 inst_cell_121_83 (.BL(BL83),.BLN(BLN83),.WL(WL121));
sram_cell_6t_5 inst_cell_121_84 (.BL(BL84),.BLN(BLN84),.WL(WL121));
sram_cell_6t_5 inst_cell_121_85 (.BL(BL85),.BLN(BLN85),.WL(WL121));
sram_cell_6t_5 inst_cell_121_86 (.BL(BL86),.BLN(BLN86),.WL(WL121));
sram_cell_6t_5 inst_cell_121_87 (.BL(BL87),.BLN(BLN87),.WL(WL121));
sram_cell_6t_5 inst_cell_121_88 (.BL(BL88),.BLN(BLN88),.WL(WL121));
sram_cell_6t_5 inst_cell_121_89 (.BL(BL89),.BLN(BLN89),.WL(WL121));
sram_cell_6t_5 inst_cell_121_90 (.BL(BL90),.BLN(BLN90),.WL(WL121));
sram_cell_6t_5 inst_cell_121_91 (.BL(BL91),.BLN(BLN91),.WL(WL121));
sram_cell_6t_5 inst_cell_121_92 (.BL(BL92),.BLN(BLN92),.WL(WL121));
sram_cell_6t_5 inst_cell_121_93 (.BL(BL93),.BLN(BLN93),.WL(WL121));
sram_cell_6t_5 inst_cell_121_94 (.BL(BL94),.BLN(BLN94),.WL(WL121));
sram_cell_6t_5 inst_cell_121_95 (.BL(BL95),.BLN(BLN95),.WL(WL121));
sram_cell_6t_5 inst_cell_121_96 (.BL(BL96),.BLN(BLN96),.WL(WL121));
sram_cell_6t_5 inst_cell_121_97 (.BL(BL97),.BLN(BLN97),.WL(WL121));
sram_cell_6t_5 inst_cell_121_98 (.BL(BL98),.BLN(BLN98),.WL(WL121));
sram_cell_6t_5 inst_cell_121_99 (.BL(BL99),.BLN(BLN99),.WL(WL121));
sram_cell_6t_5 inst_cell_121_100 (.BL(BL100),.BLN(BLN100),.WL(WL121));
sram_cell_6t_5 inst_cell_121_101 (.BL(BL101),.BLN(BLN101),.WL(WL121));
sram_cell_6t_5 inst_cell_121_102 (.BL(BL102),.BLN(BLN102),.WL(WL121));
sram_cell_6t_5 inst_cell_121_103 (.BL(BL103),.BLN(BLN103),.WL(WL121));
sram_cell_6t_5 inst_cell_121_104 (.BL(BL104),.BLN(BLN104),.WL(WL121));
sram_cell_6t_5 inst_cell_121_105 (.BL(BL105),.BLN(BLN105),.WL(WL121));
sram_cell_6t_5 inst_cell_121_106 (.BL(BL106),.BLN(BLN106),.WL(WL121));
sram_cell_6t_5 inst_cell_121_107 (.BL(BL107),.BLN(BLN107),.WL(WL121));
sram_cell_6t_5 inst_cell_121_108 (.BL(BL108),.BLN(BLN108),.WL(WL121));
sram_cell_6t_5 inst_cell_121_109 (.BL(BL109),.BLN(BLN109),.WL(WL121));
sram_cell_6t_5 inst_cell_121_110 (.BL(BL110),.BLN(BLN110),.WL(WL121));
sram_cell_6t_5 inst_cell_121_111 (.BL(BL111),.BLN(BLN111),.WL(WL121));
sram_cell_6t_5 inst_cell_121_112 (.BL(BL112),.BLN(BLN112),.WL(WL121));
sram_cell_6t_5 inst_cell_121_113 (.BL(BL113),.BLN(BLN113),.WL(WL121));
sram_cell_6t_5 inst_cell_121_114 (.BL(BL114),.BLN(BLN114),.WL(WL121));
sram_cell_6t_5 inst_cell_121_115 (.BL(BL115),.BLN(BLN115),.WL(WL121));
sram_cell_6t_5 inst_cell_121_116 (.BL(BL116),.BLN(BLN116),.WL(WL121));
sram_cell_6t_5 inst_cell_121_117 (.BL(BL117),.BLN(BLN117),.WL(WL121));
sram_cell_6t_5 inst_cell_121_118 (.BL(BL118),.BLN(BLN118),.WL(WL121));
sram_cell_6t_5 inst_cell_121_119 (.BL(BL119),.BLN(BLN119),.WL(WL121));
sram_cell_6t_5 inst_cell_121_120 (.BL(BL120),.BLN(BLN120),.WL(WL121));
sram_cell_6t_5 inst_cell_121_121 (.BL(BL121),.BLN(BLN121),.WL(WL121));
sram_cell_6t_5 inst_cell_121_122 (.BL(BL122),.BLN(BLN122),.WL(WL121));
sram_cell_6t_5 inst_cell_121_123 (.BL(BL123),.BLN(BLN123),.WL(WL121));
sram_cell_6t_5 inst_cell_121_124 (.BL(BL124),.BLN(BLN124),.WL(WL121));
sram_cell_6t_5 inst_cell_121_125 (.BL(BL125),.BLN(BLN125),.WL(WL121));
sram_cell_6t_5 inst_cell_121_126 (.BL(BL126),.BLN(BLN126),.WL(WL121));
sram_cell_6t_5 inst_cell_121_127 (.BL(BL127),.BLN(BLN127),.WL(WL121));
sram_cell_6t_5 inst_cell_122_0 (.BL(BL0),.BLN(BLN0),.WL(WL122));
sram_cell_6t_5 inst_cell_122_1 (.BL(BL1),.BLN(BLN1),.WL(WL122));
sram_cell_6t_5 inst_cell_122_2 (.BL(BL2),.BLN(BLN2),.WL(WL122));
sram_cell_6t_5 inst_cell_122_3 (.BL(BL3),.BLN(BLN3),.WL(WL122));
sram_cell_6t_5 inst_cell_122_4 (.BL(BL4),.BLN(BLN4),.WL(WL122));
sram_cell_6t_5 inst_cell_122_5 (.BL(BL5),.BLN(BLN5),.WL(WL122));
sram_cell_6t_5 inst_cell_122_6 (.BL(BL6),.BLN(BLN6),.WL(WL122));
sram_cell_6t_5 inst_cell_122_7 (.BL(BL7),.BLN(BLN7),.WL(WL122));
sram_cell_6t_5 inst_cell_122_8 (.BL(BL8),.BLN(BLN8),.WL(WL122));
sram_cell_6t_5 inst_cell_122_9 (.BL(BL9),.BLN(BLN9),.WL(WL122));
sram_cell_6t_5 inst_cell_122_10 (.BL(BL10),.BLN(BLN10),.WL(WL122));
sram_cell_6t_5 inst_cell_122_11 (.BL(BL11),.BLN(BLN11),.WL(WL122));
sram_cell_6t_5 inst_cell_122_12 (.BL(BL12),.BLN(BLN12),.WL(WL122));
sram_cell_6t_5 inst_cell_122_13 (.BL(BL13),.BLN(BLN13),.WL(WL122));
sram_cell_6t_5 inst_cell_122_14 (.BL(BL14),.BLN(BLN14),.WL(WL122));
sram_cell_6t_5 inst_cell_122_15 (.BL(BL15),.BLN(BLN15),.WL(WL122));
sram_cell_6t_5 inst_cell_122_16 (.BL(BL16),.BLN(BLN16),.WL(WL122));
sram_cell_6t_5 inst_cell_122_17 (.BL(BL17),.BLN(BLN17),.WL(WL122));
sram_cell_6t_5 inst_cell_122_18 (.BL(BL18),.BLN(BLN18),.WL(WL122));
sram_cell_6t_5 inst_cell_122_19 (.BL(BL19),.BLN(BLN19),.WL(WL122));
sram_cell_6t_5 inst_cell_122_20 (.BL(BL20),.BLN(BLN20),.WL(WL122));
sram_cell_6t_5 inst_cell_122_21 (.BL(BL21),.BLN(BLN21),.WL(WL122));
sram_cell_6t_5 inst_cell_122_22 (.BL(BL22),.BLN(BLN22),.WL(WL122));
sram_cell_6t_5 inst_cell_122_23 (.BL(BL23),.BLN(BLN23),.WL(WL122));
sram_cell_6t_5 inst_cell_122_24 (.BL(BL24),.BLN(BLN24),.WL(WL122));
sram_cell_6t_5 inst_cell_122_25 (.BL(BL25),.BLN(BLN25),.WL(WL122));
sram_cell_6t_5 inst_cell_122_26 (.BL(BL26),.BLN(BLN26),.WL(WL122));
sram_cell_6t_5 inst_cell_122_27 (.BL(BL27),.BLN(BLN27),.WL(WL122));
sram_cell_6t_5 inst_cell_122_28 (.BL(BL28),.BLN(BLN28),.WL(WL122));
sram_cell_6t_5 inst_cell_122_29 (.BL(BL29),.BLN(BLN29),.WL(WL122));
sram_cell_6t_5 inst_cell_122_30 (.BL(BL30),.BLN(BLN30),.WL(WL122));
sram_cell_6t_5 inst_cell_122_31 (.BL(BL31),.BLN(BLN31),.WL(WL122));
sram_cell_6t_5 inst_cell_122_32 (.BL(BL32),.BLN(BLN32),.WL(WL122));
sram_cell_6t_5 inst_cell_122_33 (.BL(BL33),.BLN(BLN33),.WL(WL122));
sram_cell_6t_5 inst_cell_122_34 (.BL(BL34),.BLN(BLN34),.WL(WL122));
sram_cell_6t_5 inst_cell_122_35 (.BL(BL35),.BLN(BLN35),.WL(WL122));
sram_cell_6t_5 inst_cell_122_36 (.BL(BL36),.BLN(BLN36),.WL(WL122));
sram_cell_6t_5 inst_cell_122_37 (.BL(BL37),.BLN(BLN37),.WL(WL122));
sram_cell_6t_5 inst_cell_122_38 (.BL(BL38),.BLN(BLN38),.WL(WL122));
sram_cell_6t_5 inst_cell_122_39 (.BL(BL39),.BLN(BLN39),.WL(WL122));
sram_cell_6t_5 inst_cell_122_40 (.BL(BL40),.BLN(BLN40),.WL(WL122));
sram_cell_6t_5 inst_cell_122_41 (.BL(BL41),.BLN(BLN41),.WL(WL122));
sram_cell_6t_5 inst_cell_122_42 (.BL(BL42),.BLN(BLN42),.WL(WL122));
sram_cell_6t_5 inst_cell_122_43 (.BL(BL43),.BLN(BLN43),.WL(WL122));
sram_cell_6t_5 inst_cell_122_44 (.BL(BL44),.BLN(BLN44),.WL(WL122));
sram_cell_6t_5 inst_cell_122_45 (.BL(BL45),.BLN(BLN45),.WL(WL122));
sram_cell_6t_5 inst_cell_122_46 (.BL(BL46),.BLN(BLN46),.WL(WL122));
sram_cell_6t_5 inst_cell_122_47 (.BL(BL47),.BLN(BLN47),.WL(WL122));
sram_cell_6t_5 inst_cell_122_48 (.BL(BL48),.BLN(BLN48),.WL(WL122));
sram_cell_6t_5 inst_cell_122_49 (.BL(BL49),.BLN(BLN49),.WL(WL122));
sram_cell_6t_5 inst_cell_122_50 (.BL(BL50),.BLN(BLN50),.WL(WL122));
sram_cell_6t_5 inst_cell_122_51 (.BL(BL51),.BLN(BLN51),.WL(WL122));
sram_cell_6t_5 inst_cell_122_52 (.BL(BL52),.BLN(BLN52),.WL(WL122));
sram_cell_6t_5 inst_cell_122_53 (.BL(BL53),.BLN(BLN53),.WL(WL122));
sram_cell_6t_5 inst_cell_122_54 (.BL(BL54),.BLN(BLN54),.WL(WL122));
sram_cell_6t_5 inst_cell_122_55 (.BL(BL55),.BLN(BLN55),.WL(WL122));
sram_cell_6t_5 inst_cell_122_56 (.BL(BL56),.BLN(BLN56),.WL(WL122));
sram_cell_6t_5 inst_cell_122_57 (.BL(BL57),.BLN(BLN57),.WL(WL122));
sram_cell_6t_5 inst_cell_122_58 (.BL(BL58),.BLN(BLN58),.WL(WL122));
sram_cell_6t_5 inst_cell_122_59 (.BL(BL59),.BLN(BLN59),.WL(WL122));
sram_cell_6t_5 inst_cell_122_60 (.BL(BL60),.BLN(BLN60),.WL(WL122));
sram_cell_6t_5 inst_cell_122_61 (.BL(BL61),.BLN(BLN61),.WL(WL122));
sram_cell_6t_5 inst_cell_122_62 (.BL(BL62),.BLN(BLN62),.WL(WL122));
sram_cell_6t_5 inst_cell_122_63 (.BL(BL63),.BLN(BLN63),.WL(WL122));
sram_cell_6t_5 inst_cell_122_64 (.BL(BL64),.BLN(BLN64),.WL(WL122));
sram_cell_6t_5 inst_cell_122_65 (.BL(BL65),.BLN(BLN65),.WL(WL122));
sram_cell_6t_5 inst_cell_122_66 (.BL(BL66),.BLN(BLN66),.WL(WL122));
sram_cell_6t_5 inst_cell_122_67 (.BL(BL67),.BLN(BLN67),.WL(WL122));
sram_cell_6t_5 inst_cell_122_68 (.BL(BL68),.BLN(BLN68),.WL(WL122));
sram_cell_6t_5 inst_cell_122_69 (.BL(BL69),.BLN(BLN69),.WL(WL122));
sram_cell_6t_5 inst_cell_122_70 (.BL(BL70),.BLN(BLN70),.WL(WL122));
sram_cell_6t_5 inst_cell_122_71 (.BL(BL71),.BLN(BLN71),.WL(WL122));
sram_cell_6t_5 inst_cell_122_72 (.BL(BL72),.BLN(BLN72),.WL(WL122));
sram_cell_6t_5 inst_cell_122_73 (.BL(BL73),.BLN(BLN73),.WL(WL122));
sram_cell_6t_5 inst_cell_122_74 (.BL(BL74),.BLN(BLN74),.WL(WL122));
sram_cell_6t_5 inst_cell_122_75 (.BL(BL75),.BLN(BLN75),.WL(WL122));
sram_cell_6t_5 inst_cell_122_76 (.BL(BL76),.BLN(BLN76),.WL(WL122));
sram_cell_6t_5 inst_cell_122_77 (.BL(BL77),.BLN(BLN77),.WL(WL122));
sram_cell_6t_5 inst_cell_122_78 (.BL(BL78),.BLN(BLN78),.WL(WL122));
sram_cell_6t_5 inst_cell_122_79 (.BL(BL79),.BLN(BLN79),.WL(WL122));
sram_cell_6t_5 inst_cell_122_80 (.BL(BL80),.BLN(BLN80),.WL(WL122));
sram_cell_6t_5 inst_cell_122_81 (.BL(BL81),.BLN(BLN81),.WL(WL122));
sram_cell_6t_5 inst_cell_122_82 (.BL(BL82),.BLN(BLN82),.WL(WL122));
sram_cell_6t_5 inst_cell_122_83 (.BL(BL83),.BLN(BLN83),.WL(WL122));
sram_cell_6t_5 inst_cell_122_84 (.BL(BL84),.BLN(BLN84),.WL(WL122));
sram_cell_6t_5 inst_cell_122_85 (.BL(BL85),.BLN(BLN85),.WL(WL122));
sram_cell_6t_5 inst_cell_122_86 (.BL(BL86),.BLN(BLN86),.WL(WL122));
sram_cell_6t_5 inst_cell_122_87 (.BL(BL87),.BLN(BLN87),.WL(WL122));
sram_cell_6t_5 inst_cell_122_88 (.BL(BL88),.BLN(BLN88),.WL(WL122));
sram_cell_6t_5 inst_cell_122_89 (.BL(BL89),.BLN(BLN89),.WL(WL122));
sram_cell_6t_5 inst_cell_122_90 (.BL(BL90),.BLN(BLN90),.WL(WL122));
sram_cell_6t_5 inst_cell_122_91 (.BL(BL91),.BLN(BLN91),.WL(WL122));
sram_cell_6t_5 inst_cell_122_92 (.BL(BL92),.BLN(BLN92),.WL(WL122));
sram_cell_6t_5 inst_cell_122_93 (.BL(BL93),.BLN(BLN93),.WL(WL122));
sram_cell_6t_5 inst_cell_122_94 (.BL(BL94),.BLN(BLN94),.WL(WL122));
sram_cell_6t_5 inst_cell_122_95 (.BL(BL95),.BLN(BLN95),.WL(WL122));
sram_cell_6t_5 inst_cell_122_96 (.BL(BL96),.BLN(BLN96),.WL(WL122));
sram_cell_6t_5 inst_cell_122_97 (.BL(BL97),.BLN(BLN97),.WL(WL122));
sram_cell_6t_5 inst_cell_122_98 (.BL(BL98),.BLN(BLN98),.WL(WL122));
sram_cell_6t_5 inst_cell_122_99 (.BL(BL99),.BLN(BLN99),.WL(WL122));
sram_cell_6t_5 inst_cell_122_100 (.BL(BL100),.BLN(BLN100),.WL(WL122));
sram_cell_6t_5 inst_cell_122_101 (.BL(BL101),.BLN(BLN101),.WL(WL122));
sram_cell_6t_5 inst_cell_122_102 (.BL(BL102),.BLN(BLN102),.WL(WL122));
sram_cell_6t_5 inst_cell_122_103 (.BL(BL103),.BLN(BLN103),.WL(WL122));
sram_cell_6t_5 inst_cell_122_104 (.BL(BL104),.BLN(BLN104),.WL(WL122));
sram_cell_6t_5 inst_cell_122_105 (.BL(BL105),.BLN(BLN105),.WL(WL122));
sram_cell_6t_5 inst_cell_122_106 (.BL(BL106),.BLN(BLN106),.WL(WL122));
sram_cell_6t_5 inst_cell_122_107 (.BL(BL107),.BLN(BLN107),.WL(WL122));
sram_cell_6t_5 inst_cell_122_108 (.BL(BL108),.BLN(BLN108),.WL(WL122));
sram_cell_6t_5 inst_cell_122_109 (.BL(BL109),.BLN(BLN109),.WL(WL122));
sram_cell_6t_5 inst_cell_122_110 (.BL(BL110),.BLN(BLN110),.WL(WL122));
sram_cell_6t_5 inst_cell_122_111 (.BL(BL111),.BLN(BLN111),.WL(WL122));
sram_cell_6t_5 inst_cell_122_112 (.BL(BL112),.BLN(BLN112),.WL(WL122));
sram_cell_6t_5 inst_cell_122_113 (.BL(BL113),.BLN(BLN113),.WL(WL122));
sram_cell_6t_5 inst_cell_122_114 (.BL(BL114),.BLN(BLN114),.WL(WL122));
sram_cell_6t_5 inst_cell_122_115 (.BL(BL115),.BLN(BLN115),.WL(WL122));
sram_cell_6t_5 inst_cell_122_116 (.BL(BL116),.BLN(BLN116),.WL(WL122));
sram_cell_6t_5 inst_cell_122_117 (.BL(BL117),.BLN(BLN117),.WL(WL122));
sram_cell_6t_5 inst_cell_122_118 (.BL(BL118),.BLN(BLN118),.WL(WL122));
sram_cell_6t_5 inst_cell_122_119 (.BL(BL119),.BLN(BLN119),.WL(WL122));
sram_cell_6t_5 inst_cell_122_120 (.BL(BL120),.BLN(BLN120),.WL(WL122));
sram_cell_6t_5 inst_cell_122_121 (.BL(BL121),.BLN(BLN121),.WL(WL122));
sram_cell_6t_5 inst_cell_122_122 (.BL(BL122),.BLN(BLN122),.WL(WL122));
sram_cell_6t_5 inst_cell_122_123 (.BL(BL123),.BLN(BLN123),.WL(WL122));
sram_cell_6t_5 inst_cell_122_124 (.BL(BL124),.BLN(BLN124),.WL(WL122));
sram_cell_6t_5 inst_cell_122_125 (.BL(BL125),.BLN(BLN125),.WL(WL122));
sram_cell_6t_5 inst_cell_122_126 (.BL(BL126),.BLN(BLN126),.WL(WL122));
sram_cell_6t_5 inst_cell_122_127 (.BL(BL127),.BLN(BLN127),.WL(WL122));
sram_cell_6t_5 inst_cell_123_0 (.BL(BL0),.BLN(BLN0),.WL(WL123));
sram_cell_6t_5 inst_cell_123_1 (.BL(BL1),.BLN(BLN1),.WL(WL123));
sram_cell_6t_5 inst_cell_123_2 (.BL(BL2),.BLN(BLN2),.WL(WL123));
sram_cell_6t_5 inst_cell_123_3 (.BL(BL3),.BLN(BLN3),.WL(WL123));
sram_cell_6t_5 inst_cell_123_4 (.BL(BL4),.BLN(BLN4),.WL(WL123));
sram_cell_6t_5 inst_cell_123_5 (.BL(BL5),.BLN(BLN5),.WL(WL123));
sram_cell_6t_5 inst_cell_123_6 (.BL(BL6),.BLN(BLN6),.WL(WL123));
sram_cell_6t_5 inst_cell_123_7 (.BL(BL7),.BLN(BLN7),.WL(WL123));
sram_cell_6t_5 inst_cell_123_8 (.BL(BL8),.BLN(BLN8),.WL(WL123));
sram_cell_6t_5 inst_cell_123_9 (.BL(BL9),.BLN(BLN9),.WL(WL123));
sram_cell_6t_5 inst_cell_123_10 (.BL(BL10),.BLN(BLN10),.WL(WL123));
sram_cell_6t_5 inst_cell_123_11 (.BL(BL11),.BLN(BLN11),.WL(WL123));
sram_cell_6t_5 inst_cell_123_12 (.BL(BL12),.BLN(BLN12),.WL(WL123));
sram_cell_6t_5 inst_cell_123_13 (.BL(BL13),.BLN(BLN13),.WL(WL123));
sram_cell_6t_5 inst_cell_123_14 (.BL(BL14),.BLN(BLN14),.WL(WL123));
sram_cell_6t_5 inst_cell_123_15 (.BL(BL15),.BLN(BLN15),.WL(WL123));
sram_cell_6t_5 inst_cell_123_16 (.BL(BL16),.BLN(BLN16),.WL(WL123));
sram_cell_6t_5 inst_cell_123_17 (.BL(BL17),.BLN(BLN17),.WL(WL123));
sram_cell_6t_5 inst_cell_123_18 (.BL(BL18),.BLN(BLN18),.WL(WL123));
sram_cell_6t_5 inst_cell_123_19 (.BL(BL19),.BLN(BLN19),.WL(WL123));
sram_cell_6t_5 inst_cell_123_20 (.BL(BL20),.BLN(BLN20),.WL(WL123));
sram_cell_6t_5 inst_cell_123_21 (.BL(BL21),.BLN(BLN21),.WL(WL123));
sram_cell_6t_5 inst_cell_123_22 (.BL(BL22),.BLN(BLN22),.WL(WL123));
sram_cell_6t_5 inst_cell_123_23 (.BL(BL23),.BLN(BLN23),.WL(WL123));
sram_cell_6t_5 inst_cell_123_24 (.BL(BL24),.BLN(BLN24),.WL(WL123));
sram_cell_6t_5 inst_cell_123_25 (.BL(BL25),.BLN(BLN25),.WL(WL123));
sram_cell_6t_5 inst_cell_123_26 (.BL(BL26),.BLN(BLN26),.WL(WL123));
sram_cell_6t_5 inst_cell_123_27 (.BL(BL27),.BLN(BLN27),.WL(WL123));
sram_cell_6t_5 inst_cell_123_28 (.BL(BL28),.BLN(BLN28),.WL(WL123));
sram_cell_6t_5 inst_cell_123_29 (.BL(BL29),.BLN(BLN29),.WL(WL123));
sram_cell_6t_5 inst_cell_123_30 (.BL(BL30),.BLN(BLN30),.WL(WL123));
sram_cell_6t_5 inst_cell_123_31 (.BL(BL31),.BLN(BLN31),.WL(WL123));
sram_cell_6t_5 inst_cell_123_32 (.BL(BL32),.BLN(BLN32),.WL(WL123));
sram_cell_6t_5 inst_cell_123_33 (.BL(BL33),.BLN(BLN33),.WL(WL123));
sram_cell_6t_5 inst_cell_123_34 (.BL(BL34),.BLN(BLN34),.WL(WL123));
sram_cell_6t_5 inst_cell_123_35 (.BL(BL35),.BLN(BLN35),.WL(WL123));
sram_cell_6t_5 inst_cell_123_36 (.BL(BL36),.BLN(BLN36),.WL(WL123));
sram_cell_6t_5 inst_cell_123_37 (.BL(BL37),.BLN(BLN37),.WL(WL123));
sram_cell_6t_5 inst_cell_123_38 (.BL(BL38),.BLN(BLN38),.WL(WL123));
sram_cell_6t_5 inst_cell_123_39 (.BL(BL39),.BLN(BLN39),.WL(WL123));
sram_cell_6t_5 inst_cell_123_40 (.BL(BL40),.BLN(BLN40),.WL(WL123));
sram_cell_6t_5 inst_cell_123_41 (.BL(BL41),.BLN(BLN41),.WL(WL123));
sram_cell_6t_5 inst_cell_123_42 (.BL(BL42),.BLN(BLN42),.WL(WL123));
sram_cell_6t_5 inst_cell_123_43 (.BL(BL43),.BLN(BLN43),.WL(WL123));
sram_cell_6t_5 inst_cell_123_44 (.BL(BL44),.BLN(BLN44),.WL(WL123));
sram_cell_6t_5 inst_cell_123_45 (.BL(BL45),.BLN(BLN45),.WL(WL123));
sram_cell_6t_5 inst_cell_123_46 (.BL(BL46),.BLN(BLN46),.WL(WL123));
sram_cell_6t_5 inst_cell_123_47 (.BL(BL47),.BLN(BLN47),.WL(WL123));
sram_cell_6t_5 inst_cell_123_48 (.BL(BL48),.BLN(BLN48),.WL(WL123));
sram_cell_6t_5 inst_cell_123_49 (.BL(BL49),.BLN(BLN49),.WL(WL123));
sram_cell_6t_5 inst_cell_123_50 (.BL(BL50),.BLN(BLN50),.WL(WL123));
sram_cell_6t_5 inst_cell_123_51 (.BL(BL51),.BLN(BLN51),.WL(WL123));
sram_cell_6t_5 inst_cell_123_52 (.BL(BL52),.BLN(BLN52),.WL(WL123));
sram_cell_6t_5 inst_cell_123_53 (.BL(BL53),.BLN(BLN53),.WL(WL123));
sram_cell_6t_5 inst_cell_123_54 (.BL(BL54),.BLN(BLN54),.WL(WL123));
sram_cell_6t_5 inst_cell_123_55 (.BL(BL55),.BLN(BLN55),.WL(WL123));
sram_cell_6t_5 inst_cell_123_56 (.BL(BL56),.BLN(BLN56),.WL(WL123));
sram_cell_6t_5 inst_cell_123_57 (.BL(BL57),.BLN(BLN57),.WL(WL123));
sram_cell_6t_5 inst_cell_123_58 (.BL(BL58),.BLN(BLN58),.WL(WL123));
sram_cell_6t_5 inst_cell_123_59 (.BL(BL59),.BLN(BLN59),.WL(WL123));
sram_cell_6t_5 inst_cell_123_60 (.BL(BL60),.BLN(BLN60),.WL(WL123));
sram_cell_6t_5 inst_cell_123_61 (.BL(BL61),.BLN(BLN61),.WL(WL123));
sram_cell_6t_5 inst_cell_123_62 (.BL(BL62),.BLN(BLN62),.WL(WL123));
sram_cell_6t_5 inst_cell_123_63 (.BL(BL63),.BLN(BLN63),.WL(WL123));
sram_cell_6t_5 inst_cell_123_64 (.BL(BL64),.BLN(BLN64),.WL(WL123));
sram_cell_6t_5 inst_cell_123_65 (.BL(BL65),.BLN(BLN65),.WL(WL123));
sram_cell_6t_5 inst_cell_123_66 (.BL(BL66),.BLN(BLN66),.WL(WL123));
sram_cell_6t_5 inst_cell_123_67 (.BL(BL67),.BLN(BLN67),.WL(WL123));
sram_cell_6t_5 inst_cell_123_68 (.BL(BL68),.BLN(BLN68),.WL(WL123));
sram_cell_6t_5 inst_cell_123_69 (.BL(BL69),.BLN(BLN69),.WL(WL123));
sram_cell_6t_5 inst_cell_123_70 (.BL(BL70),.BLN(BLN70),.WL(WL123));
sram_cell_6t_5 inst_cell_123_71 (.BL(BL71),.BLN(BLN71),.WL(WL123));
sram_cell_6t_5 inst_cell_123_72 (.BL(BL72),.BLN(BLN72),.WL(WL123));
sram_cell_6t_5 inst_cell_123_73 (.BL(BL73),.BLN(BLN73),.WL(WL123));
sram_cell_6t_5 inst_cell_123_74 (.BL(BL74),.BLN(BLN74),.WL(WL123));
sram_cell_6t_5 inst_cell_123_75 (.BL(BL75),.BLN(BLN75),.WL(WL123));
sram_cell_6t_5 inst_cell_123_76 (.BL(BL76),.BLN(BLN76),.WL(WL123));
sram_cell_6t_5 inst_cell_123_77 (.BL(BL77),.BLN(BLN77),.WL(WL123));
sram_cell_6t_5 inst_cell_123_78 (.BL(BL78),.BLN(BLN78),.WL(WL123));
sram_cell_6t_5 inst_cell_123_79 (.BL(BL79),.BLN(BLN79),.WL(WL123));
sram_cell_6t_5 inst_cell_123_80 (.BL(BL80),.BLN(BLN80),.WL(WL123));
sram_cell_6t_5 inst_cell_123_81 (.BL(BL81),.BLN(BLN81),.WL(WL123));
sram_cell_6t_5 inst_cell_123_82 (.BL(BL82),.BLN(BLN82),.WL(WL123));
sram_cell_6t_5 inst_cell_123_83 (.BL(BL83),.BLN(BLN83),.WL(WL123));
sram_cell_6t_5 inst_cell_123_84 (.BL(BL84),.BLN(BLN84),.WL(WL123));
sram_cell_6t_5 inst_cell_123_85 (.BL(BL85),.BLN(BLN85),.WL(WL123));
sram_cell_6t_5 inst_cell_123_86 (.BL(BL86),.BLN(BLN86),.WL(WL123));
sram_cell_6t_5 inst_cell_123_87 (.BL(BL87),.BLN(BLN87),.WL(WL123));
sram_cell_6t_5 inst_cell_123_88 (.BL(BL88),.BLN(BLN88),.WL(WL123));
sram_cell_6t_5 inst_cell_123_89 (.BL(BL89),.BLN(BLN89),.WL(WL123));
sram_cell_6t_5 inst_cell_123_90 (.BL(BL90),.BLN(BLN90),.WL(WL123));
sram_cell_6t_5 inst_cell_123_91 (.BL(BL91),.BLN(BLN91),.WL(WL123));
sram_cell_6t_5 inst_cell_123_92 (.BL(BL92),.BLN(BLN92),.WL(WL123));
sram_cell_6t_5 inst_cell_123_93 (.BL(BL93),.BLN(BLN93),.WL(WL123));
sram_cell_6t_5 inst_cell_123_94 (.BL(BL94),.BLN(BLN94),.WL(WL123));
sram_cell_6t_5 inst_cell_123_95 (.BL(BL95),.BLN(BLN95),.WL(WL123));
sram_cell_6t_5 inst_cell_123_96 (.BL(BL96),.BLN(BLN96),.WL(WL123));
sram_cell_6t_5 inst_cell_123_97 (.BL(BL97),.BLN(BLN97),.WL(WL123));
sram_cell_6t_5 inst_cell_123_98 (.BL(BL98),.BLN(BLN98),.WL(WL123));
sram_cell_6t_5 inst_cell_123_99 (.BL(BL99),.BLN(BLN99),.WL(WL123));
sram_cell_6t_5 inst_cell_123_100 (.BL(BL100),.BLN(BLN100),.WL(WL123));
sram_cell_6t_5 inst_cell_123_101 (.BL(BL101),.BLN(BLN101),.WL(WL123));
sram_cell_6t_5 inst_cell_123_102 (.BL(BL102),.BLN(BLN102),.WL(WL123));
sram_cell_6t_5 inst_cell_123_103 (.BL(BL103),.BLN(BLN103),.WL(WL123));
sram_cell_6t_5 inst_cell_123_104 (.BL(BL104),.BLN(BLN104),.WL(WL123));
sram_cell_6t_5 inst_cell_123_105 (.BL(BL105),.BLN(BLN105),.WL(WL123));
sram_cell_6t_5 inst_cell_123_106 (.BL(BL106),.BLN(BLN106),.WL(WL123));
sram_cell_6t_5 inst_cell_123_107 (.BL(BL107),.BLN(BLN107),.WL(WL123));
sram_cell_6t_5 inst_cell_123_108 (.BL(BL108),.BLN(BLN108),.WL(WL123));
sram_cell_6t_5 inst_cell_123_109 (.BL(BL109),.BLN(BLN109),.WL(WL123));
sram_cell_6t_5 inst_cell_123_110 (.BL(BL110),.BLN(BLN110),.WL(WL123));
sram_cell_6t_5 inst_cell_123_111 (.BL(BL111),.BLN(BLN111),.WL(WL123));
sram_cell_6t_5 inst_cell_123_112 (.BL(BL112),.BLN(BLN112),.WL(WL123));
sram_cell_6t_5 inst_cell_123_113 (.BL(BL113),.BLN(BLN113),.WL(WL123));
sram_cell_6t_5 inst_cell_123_114 (.BL(BL114),.BLN(BLN114),.WL(WL123));
sram_cell_6t_5 inst_cell_123_115 (.BL(BL115),.BLN(BLN115),.WL(WL123));
sram_cell_6t_5 inst_cell_123_116 (.BL(BL116),.BLN(BLN116),.WL(WL123));
sram_cell_6t_5 inst_cell_123_117 (.BL(BL117),.BLN(BLN117),.WL(WL123));
sram_cell_6t_5 inst_cell_123_118 (.BL(BL118),.BLN(BLN118),.WL(WL123));
sram_cell_6t_5 inst_cell_123_119 (.BL(BL119),.BLN(BLN119),.WL(WL123));
sram_cell_6t_5 inst_cell_123_120 (.BL(BL120),.BLN(BLN120),.WL(WL123));
sram_cell_6t_5 inst_cell_123_121 (.BL(BL121),.BLN(BLN121),.WL(WL123));
sram_cell_6t_5 inst_cell_123_122 (.BL(BL122),.BLN(BLN122),.WL(WL123));
sram_cell_6t_5 inst_cell_123_123 (.BL(BL123),.BLN(BLN123),.WL(WL123));
sram_cell_6t_5 inst_cell_123_124 (.BL(BL124),.BLN(BLN124),.WL(WL123));
sram_cell_6t_5 inst_cell_123_125 (.BL(BL125),.BLN(BLN125),.WL(WL123));
sram_cell_6t_5 inst_cell_123_126 (.BL(BL126),.BLN(BLN126),.WL(WL123));
sram_cell_6t_5 inst_cell_123_127 (.BL(BL127),.BLN(BLN127),.WL(WL123));
sram_cell_6t_5 inst_cell_124_0 (.BL(BL0),.BLN(BLN0),.WL(WL124));
sram_cell_6t_5 inst_cell_124_1 (.BL(BL1),.BLN(BLN1),.WL(WL124));
sram_cell_6t_5 inst_cell_124_2 (.BL(BL2),.BLN(BLN2),.WL(WL124));
sram_cell_6t_5 inst_cell_124_3 (.BL(BL3),.BLN(BLN3),.WL(WL124));
sram_cell_6t_5 inst_cell_124_4 (.BL(BL4),.BLN(BLN4),.WL(WL124));
sram_cell_6t_5 inst_cell_124_5 (.BL(BL5),.BLN(BLN5),.WL(WL124));
sram_cell_6t_5 inst_cell_124_6 (.BL(BL6),.BLN(BLN6),.WL(WL124));
sram_cell_6t_5 inst_cell_124_7 (.BL(BL7),.BLN(BLN7),.WL(WL124));
sram_cell_6t_5 inst_cell_124_8 (.BL(BL8),.BLN(BLN8),.WL(WL124));
sram_cell_6t_5 inst_cell_124_9 (.BL(BL9),.BLN(BLN9),.WL(WL124));
sram_cell_6t_5 inst_cell_124_10 (.BL(BL10),.BLN(BLN10),.WL(WL124));
sram_cell_6t_5 inst_cell_124_11 (.BL(BL11),.BLN(BLN11),.WL(WL124));
sram_cell_6t_5 inst_cell_124_12 (.BL(BL12),.BLN(BLN12),.WL(WL124));
sram_cell_6t_5 inst_cell_124_13 (.BL(BL13),.BLN(BLN13),.WL(WL124));
sram_cell_6t_5 inst_cell_124_14 (.BL(BL14),.BLN(BLN14),.WL(WL124));
sram_cell_6t_5 inst_cell_124_15 (.BL(BL15),.BLN(BLN15),.WL(WL124));
sram_cell_6t_5 inst_cell_124_16 (.BL(BL16),.BLN(BLN16),.WL(WL124));
sram_cell_6t_5 inst_cell_124_17 (.BL(BL17),.BLN(BLN17),.WL(WL124));
sram_cell_6t_5 inst_cell_124_18 (.BL(BL18),.BLN(BLN18),.WL(WL124));
sram_cell_6t_5 inst_cell_124_19 (.BL(BL19),.BLN(BLN19),.WL(WL124));
sram_cell_6t_5 inst_cell_124_20 (.BL(BL20),.BLN(BLN20),.WL(WL124));
sram_cell_6t_5 inst_cell_124_21 (.BL(BL21),.BLN(BLN21),.WL(WL124));
sram_cell_6t_5 inst_cell_124_22 (.BL(BL22),.BLN(BLN22),.WL(WL124));
sram_cell_6t_5 inst_cell_124_23 (.BL(BL23),.BLN(BLN23),.WL(WL124));
sram_cell_6t_5 inst_cell_124_24 (.BL(BL24),.BLN(BLN24),.WL(WL124));
sram_cell_6t_5 inst_cell_124_25 (.BL(BL25),.BLN(BLN25),.WL(WL124));
sram_cell_6t_5 inst_cell_124_26 (.BL(BL26),.BLN(BLN26),.WL(WL124));
sram_cell_6t_5 inst_cell_124_27 (.BL(BL27),.BLN(BLN27),.WL(WL124));
sram_cell_6t_5 inst_cell_124_28 (.BL(BL28),.BLN(BLN28),.WL(WL124));
sram_cell_6t_5 inst_cell_124_29 (.BL(BL29),.BLN(BLN29),.WL(WL124));
sram_cell_6t_5 inst_cell_124_30 (.BL(BL30),.BLN(BLN30),.WL(WL124));
sram_cell_6t_5 inst_cell_124_31 (.BL(BL31),.BLN(BLN31),.WL(WL124));
sram_cell_6t_5 inst_cell_124_32 (.BL(BL32),.BLN(BLN32),.WL(WL124));
sram_cell_6t_5 inst_cell_124_33 (.BL(BL33),.BLN(BLN33),.WL(WL124));
sram_cell_6t_5 inst_cell_124_34 (.BL(BL34),.BLN(BLN34),.WL(WL124));
sram_cell_6t_5 inst_cell_124_35 (.BL(BL35),.BLN(BLN35),.WL(WL124));
sram_cell_6t_5 inst_cell_124_36 (.BL(BL36),.BLN(BLN36),.WL(WL124));
sram_cell_6t_5 inst_cell_124_37 (.BL(BL37),.BLN(BLN37),.WL(WL124));
sram_cell_6t_5 inst_cell_124_38 (.BL(BL38),.BLN(BLN38),.WL(WL124));
sram_cell_6t_5 inst_cell_124_39 (.BL(BL39),.BLN(BLN39),.WL(WL124));
sram_cell_6t_5 inst_cell_124_40 (.BL(BL40),.BLN(BLN40),.WL(WL124));
sram_cell_6t_5 inst_cell_124_41 (.BL(BL41),.BLN(BLN41),.WL(WL124));
sram_cell_6t_5 inst_cell_124_42 (.BL(BL42),.BLN(BLN42),.WL(WL124));
sram_cell_6t_5 inst_cell_124_43 (.BL(BL43),.BLN(BLN43),.WL(WL124));
sram_cell_6t_5 inst_cell_124_44 (.BL(BL44),.BLN(BLN44),.WL(WL124));
sram_cell_6t_5 inst_cell_124_45 (.BL(BL45),.BLN(BLN45),.WL(WL124));
sram_cell_6t_5 inst_cell_124_46 (.BL(BL46),.BLN(BLN46),.WL(WL124));
sram_cell_6t_5 inst_cell_124_47 (.BL(BL47),.BLN(BLN47),.WL(WL124));
sram_cell_6t_5 inst_cell_124_48 (.BL(BL48),.BLN(BLN48),.WL(WL124));
sram_cell_6t_5 inst_cell_124_49 (.BL(BL49),.BLN(BLN49),.WL(WL124));
sram_cell_6t_5 inst_cell_124_50 (.BL(BL50),.BLN(BLN50),.WL(WL124));
sram_cell_6t_5 inst_cell_124_51 (.BL(BL51),.BLN(BLN51),.WL(WL124));
sram_cell_6t_5 inst_cell_124_52 (.BL(BL52),.BLN(BLN52),.WL(WL124));
sram_cell_6t_5 inst_cell_124_53 (.BL(BL53),.BLN(BLN53),.WL(WL124));
sram_cell_6t_5 inst_cell_124_54 (.BL(BL54),.BLN(BLN54),.WL(WL124));
sram_cell_6t_5 inst_cell_124_55 (.BL(BL55),.BLN(BLN55),.WL(WL124));
sram_cell_6t_5 inst_cell_124_56 (.BL(BL56),.BLN(BLN56),.WL(WL124));
sram_cell_6t_5 inst_cell_124_57 (.BL(BL57),.BLN(BLN57),.WL(WL124));
sram_cell_6t_5 inst_cell_124_58 (.BL(BL58),.BLN(BLN58),.WL(WL124));
sram_cell_6t_5 inst_cell_124_59 (.BL(BL59),.BLN(BLN59),.WL(WL124));
sram_cell_6t_5 inst_cell_124_60 (.BL(BL60),.BLN(BLN60),.WL(WL124));
sram_cell_6t_5 inst_cell_124_61 (.BL(BL61),.BLN(BLN61),.WL(WL124));
sram_cell_6t_5 inst_cell_124_62 (.BL(BL62),.BLN(BLN62),.WL(WL124));
sram_cell_6t_5 inst_cell_124_63 (.BL(BL63),.BLN(BLN63),.WL(WL124));
sram_cell_6t_5 inst_cell_124_64 (.BL(BL64),.BLN(BLN64),.WL(WL124));
sram_cell_6t_5 inst_cell_124_65 (.BL(BL65),.BLN(BLN65),.WL(WL124));
sram_cell_6t_5 inst_cell_124_66 (.BL(BL66),.BLN(BLN66),.WL(WL124));
sram_cell_6t_5 inst_cell_124_67 (.BL(BL67),.BLN(BLN67),.WL(WL124));
sram_cell_6t_5 inst_cell_124_68 (.BL(BL68),.BLN(BLN68),.WL(WL124));
sram_cell_6t_5 inst_cell_124_69 (.BL(BL69),.BLN(BLN69),.WL(WL124));
sram_cell_6t_5 inst_cell_124_70 (.BL(BL70),.BLN(BLN70),.WL(WL124));
sram_cell_6t_5 inst_cell_124_71 (.BL(BL71),.BLN(BLN71),.WL(WL124));
sram_cell_6t_5 inst_cell_124_72 (.BL(BL72),.BLN(BLN72),.WL(WL124));
sram_cell_6t_5 inst_cell_124_73 (.BL(BL73),.BLN(BLN73),.WL(WL124));
sram_cell_6t_5 inst_cell_124_74 (.BL(BL74),.BLN(BLN74),.WL(WL124));
sram_cell_6t_5 inst_cell_124_75 (.BL(BL75),.BLN(BLN75),.WL(WL124));
sram_cell_6t_5 inst_cell_124_76 (.BL(BL76),.BLN(BLN76),.WL(WL124));
sram_cell_6t_5 inst_cell_124_77 (.BL(BL77),.BLN(BLN77),.WL(WL124));
sram_cell_6t_5 inst_cell_124_78 (.BL(BL78),.BLN(BLN78),.WL(WL124));
sram_cell_6t_5 inst_cell_124_79 (.BL(BL79),.BLN(BLN79),.WL(WL124));
sram_cell_6t_5 inst_cell_124_80 (.BL(BL80),.BLN(BLN80),.WL(WL124));
sram_cell_6t_5 inst_cell_124_81 (.BL(BL81),.BLN(BLN81),.WL(WL124));
sram_cell_6t_5 inst_cell_124_82 (.BL(BL82),.BLN(BLN82),.WL(WL124));
sram_cell_6t_5 inst_cell_124_83 (.BL(BL83),.BLN(BLN83),.WL(WL124));
sram_cell_6t_5 inst_cell_124_84 (.BL(BL84),.BLN(BLN84),.WL(WL124));
sram_cell_6t_5 inst_cell_124_85 (.BL(BL85),.BLN(BLN85),.WL(WL124));
sram_cell_6t_5 inst_cell_124_86 (.BL(BL86),.BLN(BLN86),.WL(WL124));
sram_cell_6t_5 inst_cell_124_87 (.BL(BL87),.BLN(BLN87),.WL(WL124));
sram_cell_6t_5 inst_cell_124_88 (.BL(BL88),.BLN(BLN88),.WL(WL124));
sram_cell_6t_5 inst_cell_124_89 (.BL(BL89),.BLN(BLN89),.WL(WL124));
sram_cell_6t_5 inst_cell_124_90 (.BL(BL90),.BLN(BLN90),.WL(WL124));
sram_cell_6t_5 inst_cell_124_91 (.BL(BL91),.BLN(BLN91),.WL(WL124));
sram_cell_6t_5 inst_cell_124_92 (.BL(BL92),.BLN(BLN92),.WL(WL124));
sram_cell_6t_5 inst_cell_124_93 (.BL(BL93),.BLN(BLN93),.WL(WL124));
sram_cell_6t_5 inst_cell_124_94 (.BL(BL94),.BLN(BLN94),.WL(WL124));
sram_cell_6t_5 inst_cell_124_95 (.BL(BL95),.BLN(BLN95),.WL(WL124));
sram_cell_6t_5 inst_cell_124_96 (.BL(BL96),.BLN(BLN96),.WL(WL124));
sram_cell_6t_5 inst_cell_124_97 (.BL(BL97),.BLN(BLN97),.WL(WL124));
sram_cell_6t_5 inst_cell_124_98 (.BL(BL98),.BLN(BLN98),.WL(WL124));
sram_cell_6t_5 inst_cell_124_99 (.BL(BL99),.BLN(BLN99),.WL(WL124));
sram_cell_6t_5 inst_cell_124_100 (.BL(BL100),.BLN(BLN100),.WL(WL124));
sram_cell_6t_5 inst_cell_124_101 (.BL(BL101),.BLN(BLN101),.WL(WL124));
sram_cell_6t_5 inst_cell_124_102 (.BL(BL102),.BLN(BLN102),.WL(WL124));
sram_cell_6t_5 inst_cell_124_103 (.BL(BL103),.BLN(BLN103),.WL(WL124));
sram_cell_6t_5 inst_cell_124_104 (.BL(BL104),.BLN(BLN104),.WL(WL124));
sram_cell_6t_5 inst_cell_124_105 (.BL(BL105),.BLN(BLN105),.WL(WL124));
sram_cell_6t_5 inst_cell_124_106 (.BL(BL106),.BLN(BLN106),.WL(WL124));
sram_cell_6t_5 inst_cell_124_107 (.BL(BL107),.BLN(BLN107),.WL(WL124));
sram_cell_6t_5 inst_cell_124_108 (.BL(BL108),.BLN(BLN108),.WL(WL124));
sram_cell_6t_5 inst_cell_124_109 (.BL(BL109),.BLN(BLN109),.WL(WL124));
sram_cell_6t_5 inst_cell_124_110 (.BL(BL110),.BLN(BLN110),.WL(WL124));
sram_cell_6t_5 inst_cell_124_111 (.BL(BL111),.BLN(BLN111),.WL(WL124));
sram_cell_6t_5 inst_cell_124_112 (.BL(BL112),.BLN(BLN112),.WL(WL124));
sram_cell_6t_5 inst_cell_124_113 (.BL(BL113),.BLN(BLN113),.WL(WL124));
sram_cell_6t_5 inst_cell_124_114 (.BL(BL114),.BLN(BLN114),.WL(WL124));
sram_cell_6t_5 inst_cell_124_115 (.BL(BL115),.BLN(BLN115),.WL(WL124));
sram_cell_6t_5 inst_cell_124_116 (.BL(BL116),.BLN(BLN116),.WL(WL124));
sram_cell_6t_5 inst_cell_124_117 (.BL(BL117),.BLN(BLN117),.WL(WL124));
sram_cell_6t_5 inst_cell_124_118 (.BL(BL118),.BLN(BLN118),.WL(WL124));
sram_cell_6t_5 inst_cell_124_119 (.BL(BL119),.BLN(BLN119),.WL(WL124));
sram_cell_6t_5 inst_cell_124_120 (.BL(BL120),.BLN(BLN120),.WL(WL124));
sram_cell_6t_5 inst_cell_124_121 (.BL(BL121),.BLN(BLN121),.WL(WL124));
sram_cell_6t_5 inst_cell_124_122 (.BL(BL122),.BLN(BLN122),.WL(WL124));
sram_cell_6t_5 inst_cell_124_123 (.BL(BL123),.BLN(BLN123),.WL(WL124));
sram_cell_6t_5 inst_cell_124_124 (.BL(BL124),.BLN(BLN124),.WL(WL124));
sram_cell_6t_5 inst_cell_124_125 (.BL(BL125),.BLN(BLN125),.WL(WL124));
sram_cell_6t_5 inst_cell_124_126 (.BL(BL126),.BLN(BLN126),.WL(WL124));
sram_cell_6t_5 inst_cell_124_127 (.BL(BL127),.BLN(BLN127),.WL(WL124));
sram_cell_6t_5 inst_cell_125_0 (.BL(BL0),.BLN(BLN0),.WL(WL125));
sram_cell_6t_5 inst_cell_125_1 (.BL(BL1),.BLN(BLN1),.WL(WL125));
sram_cell_6t_5 inst_cell_125_2 (.BL(BL2),.BLN(BLN2),.WL(WL125));
sram_cell_6t_5 inst_cell_125_3 (.BL(BL3),.BLN(BLN3),.WL(WL125));
sram_cell_6t_5 inst_cell_125_4 (.BL(BL4),.BLN(BLN4),.WL(WL125));
sram_cell_6t_5 inst_cell_125_5 (.BL(BL5),.BLN(BLN5),.WL(WL125));
sram_cell_6t_5 inst_cell_125_6 (.BL(BL6),.BLN(BLN6),.WL(WL125));
sram_cell_6t_5 inst_cell_125_7 (.BL(BL7),.BLN(BLN7),.WL(WL125));
sram_cell_6t_5 inst_cell_125_8 (.BL(BL8),.BLN(BLN8),.WL(WL125));
sram_cell_6t_5 inst_cell_125_9 (.BL(BL9),.BLN(BLN9),.WL(WL125));
sram_cell_6t_5 inst_cell_125_10 (.BL(BL10),.BLN(BLN10),.WL(WL125));
sram_cell_6t_5 inst_cell_125_11 (.BL(BL11),.BLN(BLN11),.WL(WL125));
sram_cell_6t_5 inst_cell_125_12 (.BL(BL12),.BLN(BLN12),.WL(WL125));
sram_cell_6t_5 inst_cell_125_13 (.BL(BL13),.BLN(BLN13),.WL(WL125));
sram_cell_6t_5 inst_cell_125_14 (.BL(BL14),.BLN(BLN14),.WL(WL125));
sram_cell_6t_5 inst_cell_125_15 (.BL(BL15),.BLN(BLN15),.WL(WL125));
sram_cell_6t_5 inst_cell_125_16 (.BL(BL16),.BLN(BLN16),.WL(WL125));
sram_cell_6t_5 inst_cell_125_17 (.BL(BL17),.BLN(BLN17),.WL(WL125));
sram_cell_6t_5 inst_cell_125_18 (.BL(BL18),.BLN(BLN18),.WL(WL125));
sram_cell_6t_5 inst_cell_125_19 (.BL(BL19),.BLN(BLN19),.WL(WL125));
sram_cell_6t_5 inst_cell_125_20 (.BL(BL20),.BLN(BLN20),.WL(WL125));
sram_cell_6t_5 inst_cell_125_21 (.BL(BL21),.BLN(BLN21),.WL(WL125));
sram_cell_6t_5 inst_cell_125_22 (.BL(BL22),.BLN(BLN22),.WL(WL125));
sram_cell_6t_5 inst_cell_125_23 (.BL(BL23),.BLN(BLN23),.WL(WL125));
sram_cell_6t_5 inst_cell_125_24 (.BL(BL24),.BLN(BLN24),.WL(WL125));
sram_cell_6t_5 inst_cell_125_25 (.BL(BL25),.BLN(BLN25),.WL(WL125));
sram_cell_6t_5 inst_cell_125_26 (.BL(BL26),.BLN(BLN26),.WL(WL125));
sram_cell_6t_5 inst_cell_125_27 (.BL(BL27),.BLN(BLN27),.WL(WL125));
sram_cell_6t_5 inst_cell_125_28 (.BL(BL28),.BLN(BLN28),.WL(WL125));
sram_cell_6t_5 inst_cell_125_29 (.BL(BL29),.BLN(BLN29),.WL(WL125));
sram_cell_6t_5 inst_cell_125_30 (.BL(BL30),.BLN(BLN30),.WL(WL125));
sram_cell_6t_5 inst_cell_125_31 (.BL(BL31),.BLN(BLN31),.WL(WL125));
sram_cell_6t_5 inst_cell_125_32 (.BL(BL32),.BLN(BLN32),.WL(WL125));
sram_cell_6t_5 inst_cell_125_33 (.BL(BL33),.BLN(BLN33),.WL(WL125));
sram_cell_6t_5 inst_cell_125_34 (.BL(BL34),.BLN(BLN34),.WL(WL125));
sram_cell_6t_5 inst_cell_125_35 (.BL(BL35),.BLN(BLN35),.WL(WL125));
sram_cell_6t_5 inst_cell_125_36 (.BL(BL36),.BLN(BLN36),.WL(WL125));
sram_cell_6t_5 inst_cell_125_37 (.BL(BL37),.BLN(BLN37),.WL(WL125));
sram_cell_6t_5 inst_cell_125_38 (.BL(BL38),.BLN(BLN38),.WL(WL125));
sram_cell_6t_5 inst_cell_125_39 (.BL(BL39),.BLN(BLN39),.WL(WL125));
sram_cell_6t_5 inst_cell_125_40 (.BL(BL40),.BLN(BLN40),.WL(WL125));
sram_cell_6t_5 inst_cell_125_41 (.BL(BL41),.BLN(BLN41),.WL(WL125));
sram_cell_6t_5 inst_cell_125_42 (.BL(BL42),.BLN(BLN42),.WL(WL125));
sram_cell_6t_5 inst_cell_125_43 (.BL(BL43),.BLN(BLN43),.WL(WL125));
sram_cell_6t_5 inst_cell_125_44 (.BL(BL44),.BLN(BLN44),.WL(WL125));
sram_cell_6t_5 inst_cell_125_45 (.BL(BL45),.BLN(BLN45),.WL(WL125));
sram_cell_6t_5 inst_cell_125_46 (.BL(BL46),.BLN(BLN46),.WL(WL125));
sram_cell_6t_5 inst_cell_125_47 (.BL(BL47),.BLN(BLN47),.WL(WL125));
sram_cell_6t_5 inst_cell_125_48 (.BL(BL48),.BLN(BLN48),.WL(WL125));
sram_cell_6t_5 inst_cell_125_49 (.BL(BL49),.BLN(BLN49),.WL(WL125));
sram_cell_6t_5 inst_cell_125_50 (.BL(BL50),.BLN(BLN50),.WL(WL125));
sram_cell_6t_5 inst_cell_125_51 (.BL(BL51),.BLN(BLN51),.WL(WL125));
sram_cell_6t_5 inst_cell_125_52 (.BL(BL52),.BLN(BLN52),.WL(WL125));
sram_cell_6t_5 inst_cell_125_53 (.BL(BL53),.BLN(BLN53),.WL(WL125));
sram_cell_6t_5 inst_cell_125_54 (.BL(BL54),.BLN(BLN54),.WL(WL125));
sram_cell_6t_5 inst_cell_125_55 (.BL(BL55),.BLN(BLN55),.WL(WL125));
sram_cell_6t_5 inst_cell_125_56 (.BL(BL56),.BLN(BLN56),.WL(WL125));
sram_cell_6t_5 inst_cell_125_57 (.BL(BL57),.BLN(BLN57),.WL(WL125));
sram_cell_6t_5 inst_cell_125_58 (.BL(BL58),.BLN(BLN58),.WL(WL125));
sram_cell_6t_5 inst_cell_125_59 (.BL(BL59),.BLN(BLN59),.WL(WL125));
sram_cell_6t_5 inst_cell_125_60 (.BL(BL60),.BLN(BLN60),.WL(WL125));
sram_cell_6t_5 inst_cell_125_61 (.BL(BL61),.BLN(BLN61),.WL(WL125));
sram_cell_6t_5 inst_cell_125_62 (.BL(BL62),.BLN(BLN62),.WL(WL125));
sram_cell_6t_5 inst_cell_125_63 (.BL(BL63),.BLN(BLN63),.WL(WL125));
sram_cell_6t_5 inst_cell_125_64 (.BL(BL64),.BLN(BLN64),.WL(WL125));
sram_cell_6t_5 inst_cell_125_65 (.BL(BL65),.BLN(BLN65),.WL(WL125));
sram_cell_6t_5 inst_cell_125_66 (.BL(BL66),.BLN(BLN66),.WL(WL125));
sram_cell_6t_5 inst_cell_125_67 (.BL(BL67),.BLN(BLN67),.WL(WL125));
sram_cell_6t_5 inst_cell_125_68 (.BL(BL68),.BLN(BLN68),.WL(WL125));
sram_cell_6t_5 inst_cell_125_69 (.BL(BL69),.BLN(BLN69),.WL(WL125));
sram_cell_6t_5 inst_cell_125_70 (.BL(BL70),.BLN(BLN70),.WL(WL125));
sram_cell_6t_5 inst_cell_125_71 (.BL(BL71),.BLN(BLN71),.WL(WL125));
sram_cell_6t_5 inst_cell_125_72 (.BL(BL72),.BLN(BLN72),.WL(WL125));
sram_cell_6t_5 inst_cell_125_73 (.BL(BL73),.BLN(BLN73),.WL(WL125));
sram_cell_6t_5 inst_cell_125_74 (.BL(BL74),.BLN(BLN74),.WL(WL125));
sram_cell_6t_5 inst_cell_125_75 (.BL(BL75),.BLN(BLN75),.WL(WL125));
sram_cell_6t_5 inst_cell_125_76 (.BL(BL76),.BLN(BLN76),.WL(WL125));
sram_cell_6t_5 inst_cell_125_77 (.BL(BL77),.BLN(BLN77),.WL(WL125));
sram_cell_6t_5 inst_cell_125_78 (.BL(BL78),.BLN(BLN78),.WL(WL125));
sram_cell_6t_5 inst_cell_125_79 (.BL(BL79),.BLN(BLN79),.WL(WL125));
sram_cell_6t_5 inst_cell_125_80 (.BL(BL80),.BLN(BLN80),.WL(WL125));
sram_cell_6t_5 inst_cell_125_81 (.BL(BL81),.BLN(BLN81),.WL(WL125));
sram_cell_6t_5 inst_cell_125_82 (.BL(BL82),.BLN(BLN82),.WL(WL125));
sram_cell_6t_5 inst_cell_125_83 (.BL(BL83),.BLN(BLN83),.WL(WL125));
sram_cell_6t_5 inst_cell_125_84 (.BL(BL84),.BLN(BLN84),.WL(WL125));
sram_cell_6t_5 inst_cell_125_85 (.BL(BL85),.BLN(BLN85),.WL(WL125));
sram_cell_6t_5 inst_cell_125_86 (.BL(BL86),.BLN(BLN86),.WL(WL125));
sram_cell_6t_5 inst_cell_125_87 (.BL(BL87),.BLN(BLN87),.WL(WL125));
sram_cell_6t_5 inst_cell_125_88 (.BL(BL88),.BLN(BLN88),.WL(WL125));
sram_cell_6t_5 inst_cell_125_89 (.BL(BL89),.BLN(BLN89),.WL(WL125));
sram_cell_6t_5 inst_cell_125_90 (.BL(BL90),.BLN(BLN90),.WL(WL125));
sram_cell_6t_5 inst_cell_125_91 (.BL(BL91),.BLN(BLN91),.WL(WL125));
sram_cell_6t_5 inst_cell_125_92 (.BL(BL92),.BLN(BLN92),.WL(WL125));
sram_cell_6t_5 inst_cell_125_93 (.BL(BL93),.BLN(BLN93),.WL(WL125));
sram_cell_6t_5 inst_cell_125_94 (.BL(BL94),.BLN(BLN94),.WL(WL125));
sram_cell_6t_5 inst_cell_125_95 (.BL(BL95),.BLN(BLN95),.WL(WL125));
sram_cell_6t_5 inst_cell_125_96 (.BL(BL96),.BLN(BLN96),.WL(WL125));
sram_cell_6t_5 inst_cell_125_97 (.BL(BL97),.BLN(BLN97),.WL(WL125));
sram_cell_6t_5 inst_cell_125_98 (.BL(BL98),.BLN(BLN98),.WL(WL125));
sram_cell_6t_5 inst_cell_125_99 (.BL(BL99),.BLN(BLN99),.WL(WL125));
sram_cell_6t_5 inst_cell_125_100 (.BL(BL100),.BLN(BLN100),.WL(WL125));
sram_cell_6t_5 inst_cell_125_101 (.BL(BL101),.BLN(BLN101),.WL(WL125));
sram_cell_6t_5 inst_cell_125_102 (.BL(BL102),.BLN(BLN102),.WL(WL125));
sram_cell_6t_5 inst_cell_125_103 (.BL(BL103),.BLN(BLN103),.WL(WL125));
sram_cell_6t_5 inst_cell_125_104 (.BL(BL104),.BLN(BLN104),.WL(WL125));
sram_cell_6t_5 inst_cell_125_105 (.BL(BL105),.BLN(BLN105),.WL(WL125));
sram_cell_6t_5 inst_cell_125_106 (.BL(BL106),.BLN(BLN106),.WL(WL125));
sram_cell_6t_5 inst_cell_125_107 (.BL(BL107),.BLN(BLN107),.WL(WL125));
sram_cell_6t_5 inst_cell_125_108 (.BL(BL108),.BLN(BLN108),.WL(WL125));
sram_cell_6t_5 inst_cell_125_109 (.BL(BL109),.BLN(BLN109),.WL(WL125));
sram_cell_6t_5 inst_cell_125_110 (.BL(BL110),.BLN(BLN110),.WL(WL125));
sram_cell_6t_5 inst_cell_125_111 (.BL(BL111),.BLN(BLN111),.WL(WL125));
sram_cell_6t_5 inst_cell_125_112 (.BL(BL112),.BLN(BLN112),.WL(WL125));
sram_cell_6t_5 inst_cell_125_113 (.BL(BL113),.BLN(BLN113),.WL(WL125));
sram_cell_6t_5 inst_cell_125_114 (.BL(BL114),.BLN(BLN114),.WL(WL125));
sram_cell_6t_5 inst_cell_125_115 (.BL(BL115),.BLN(BLN115),.WL(WL125));
sram_cell_6t_5 inst_cell_125_116 (.BL(BL116),.BLN(BLN116),.WL(WL125));
sram_cell_6t_5 inst_cell_125_117 (.BL(BL117),.BLN(BLN117),.WL(WL125));
sram_cell_6t_5 inst_cell_125_118 (.BL(BL118),.BLN(BLN118),.WL(WL125));
sram_cell_6t_5 inst_cell_125_119 (.BL(BL119),.BLN(BLN119),.WL(WL125));
sram_cell_6t_5 inst_cell_125_120 (.BL(BL120),.BLN(BLN120),.WL(WL125));
sram_cell_6t_5 inst_cell_125_121 (.BL(BL121),.BLN(BLN121),.WL(WL125));
sram_cell_6t_5 inst_cell_125_122 (.BL(BL122),.BLN(BLN122),.WL(WL125));
sram_cell_6t_5 inst_cell_125_123 (.BL(BL123),.BLN(BLN123),.WL(WL125));
sram_cell_6t_5 inst_cell_125_124 (.BL(BL124),.BLN(BLN124),.WL(WL125));
sram_cell_6t_5 inst_cell_125_125 (.BL(BL125),.BLN(BLN125),.WL(WL125));
sram_cell_6t_5 inst_cell_125_126 (.BL(BL126),.BLN(BLN126),.WL(WL125));
sram_cell_6t_5 inst_cell_125_127 (.BL(BL127),.BLN(BLN127),.WL(WL125));
sram_cell_6t_5 inst_cell_126_0 (.BL(BL0),.BLN(BLN0),.WL(WL126));
sram_cell_6t_5 inst_cell_126_1 (.BL(BL1),.BLN(BLN1),.WL(WL126));
sram_cell_6t_5 inst_cell_126_2 (.BL(BL2),.BLN(BLN2),.WL(WL126));
sram_cell_6t_5 inst_cell_126_3 (.BL(BL3),.BLN(BLN3),.WL(WL126));
sram_cell_6t_5 inst_cell_126_4 (.BL(BL4),.BLN(BLN4),.WL(WL126));
sram_cell_6t_5 inst_cell_126_5 (.BL(BL5),.BLN(BLN5),.WL(WL126));
sram_cell_6t_5 inst_cell_126_6 (.BL(BL6),.BLN(BLN6),.WL(WL126));
sram_cell_6t_5 inst_cell_126_7 (.BL(BL7),.BLN(BLN7),.WL(WL126));
sram_cell_6t_5 inst_cell_126_8 (.BL(BL8),.BLN(BLN8),.WL(WL126));
sram_cell_6t_5 inst_cell_126_9 (.BL(BL9),.BLN(BLN9),.WL(WL126));
sram_cell_6t_5 inst_cell_126_10 (.BL(BL10),.BLN(BLN10),.WL(WL126));
sram_cell_6t_5 inst_cell_126_11 (.BL(BL11),.BLN(BLN11),.WL(WL126));
sram_cell_6t_5 inst_cell_126_12 (.BL(BL12),.BLN(BLN12),.WL(WL126));
sram_cell_6t_5 inst_cell_126_13 (.BL(BL13),.BLN(BLN13),.WL(WL126));
sram_cell_6t_5 inst_cell_126_14 (.BL(BL14),.BLN(BLN14),.WL(WL126));
sram_cell_6t_5 inst_cell_126_15 (.BL(BL15),.BLN(BLN15),.WL(WL126));
sram_cell_6t_5 inst_cell_126_16 (.BL(BL16),.BLN(BLN16),.WL(WL126));
sram_cell_6t_5 inst_cell_126_17 (.BL(BL17),.BLN(BLN17),.WL(WL126));
sram_cell_6t_5 inst_cell_126_18 (.BL(BL18),.BLN(BLN18),.WL(WL126));
sram_cell_6t_5 inst_cell_126_19 (.BL(BL19),.BLN(BLN19),.WL(WL126));
sram_cell_6t_5 inst_cell_126_20 (.BL(BL20),.BLN(BLN20),.WL(WL126));
sram_cell_6t_5 inst_cell_126_21 (.BL(BL21),.BLN(BLN21),.WL(WL126));
sram_cell_6t_5 inst_cell_126_22 (.BL(BL22),.BLN(BLN22),.WL(WL126));
sram_cell_6t_5 inst_cell_126_23 (.BL(BL23),.BLN(BLN23),.WL(WL126));
sram_cell_6t_5 inst_cell_126_24 (.BL(BL24),.BLN(BLN24),.WL(WL126));
sram_cell_6t_5 inst_cell_126_25 (.BL(BL25),.BLN(BLN25),.WL(WL126));
sram_cell_6t_5 inst_cell_126_26 (.BL(BL26),.BLN(BLN26),.WL(WL126));
sram_cell_6t_5 inst_cell_126_27 (.BL(BL27),.BLN(BLN27),.WL(WL126));
sram_cell_6t_5 inst_cell_126_28 (.BL(BL28),.BLN(BLN28),.WL(WL126));
sram_cell_6t_5 inst_cell_126_29 (.BL(BL29),.BLN(BLN29),.WL(WL126));
sram_cell_6t_5 inst_cell_126_30 (.BL(BL30),.BLN(BLN30),.WL(WL126));
sram_cell_6t_5 inst_cell_126_31 (.BL(BL31),.BLN(BLN31),.WL(WL126));
sram_cell_6t_5 inst_cell_126_32 (.BL(BL32),.BLN(BLN32),.WL(WL126));
sram_cell_6t_5 inst_cell_126_33 (.BL(BL33),.BLN(BLN33),.WL(WL126));
sram_cell_6t_5 inst_cell_126_34 (.BL(BL34),.BLN(BLN34),.WL(WL126));
sram_cell_6t_5 inst_cell_126_35 (.BL(BL35),.BLN(BLN35),.WL(WL126));
sram_cell_6t_5 inst_cell_126_36 (.BL(BL36),.BLN(BLN36),.WL(WL126));
sram_cell_6t_5 inst_cell_126_37 (.BL(BL37),.BLN(BLN37),.WL(WL126));
sram_cell_6t_5 inst_cell_126_38 (.BL(BL38),.BLN(BLN38),.WL(WL126));
sram_cell_6t_5 inst_cell_126_39 (.BL(BL39),.BLN(BLN39),.WL(WL126));
sram_cell_6t_5 inst_cell_126_40 (.BL(BL40),.BLN(BLN40),.WL(WL126));
sram_cell_6t_5 inst_cell_126_41 (.BL(BL41),.BLN(BLN41),.WL(WL126));
sram_cell_6t_5 inst_cell_126_42 (.BL(BL42),.BLN(BLN42),.WL(WL126));
sram_cell_6t_5 inst_cell_126_43 (.BL(BL43),.BLN(BLN43),.WL(WL126));
sram_cell_6t_5 inst_cell_126_44 (.BL(BL44),.BLN(BLN44),.WL(WL126));
sram_cell_6t_5 inst_cell_126_45 (.BL(BL45),.BLN(BLN45),.WL(WL126));
sram_cell_6t_5 inst_cell_126_46 (.BL(BL46),.BLN(BLN46),.WL(WL126));
sram_cell_6t_5 inst_cell_126_47 (.BL(BL47),.BLN(BLN47),.WL(WL126));
sram_cell_6t_5 inst_cell_126_48 (.BL(BL48),.BLN(BLN48),.WL(WL126));
sram_cell_6t_5 inst_cell_126_49 (.BL(BL49),.BLN(BLN49),.WL(WL126));
sram_cell_6t_5 inst_cell_126_50 (.BL(BL50),.BLN(BLN50),.WL(WL126));
sram_cell_6t_5 inst_cell_126_51 (.BL(BL51),.BLN(BLN51),.WL(WL126));
sram_cell_6t_5 inst_cell_126_52 (.BL(BL52),.BLN(BLN52),.WL(WL126));
sram_cell_6t_5 inst_cell_126_53 (.BL(BL53),.BLN(BLN53),.WL(WL126));
sram_cell_6t_5 inst_cell_126_54 (.BL(BL54),.BLN(BLN54),.WL(WL126));
sram_cell_6t_5 inst_cell_126_55 (.BL(BL55),.BLN(BLN55),.WL(WL126));
sram_cell_6t_5 inst_cell_126_56 (.BL(BL56),.BLN(BLN56),.WL(WL126));
sram_cell_6t_5 inst_cell_126_57 (.BL(BL57),.BLN(BLN57),.WL(WL126));
sram_cell_6t_5 inst_cell_126_58 (.BL(BL58),.BLN(BLN58),.WL(WL126));
sram_cell_6t_5 inst_cell_126_59 (.BL(BL59),.BLN(BLN59),.WL(WL126));
sram_cell_6t_5 inst_cell_126_60 (.BL(BL60),.BLN(BLN60),.WL(WL126));
sram_cell_6t_5 inst_cell_126_61 (.BL(BL61),.BLN(BLN61),.WL(WL126));
sram_cell_6t_5 inst_cell_126_62 (.BL(BL62),.BLN(BLN62),.WL(WL126));
sram_cell_6t_5 inst_cell_126_63 (.BL(BL63),.BLN(BLN63),.WL(WL126));
sram_cell_6t_5 inst_cell_126_64 (.BL(BL64),.BLN(BLN64),.WL(WL126));
sram_cell_6t_5 inst_cell_126_65 (.BL(BL65),.BLN(BLN65),.WL(WL126));
sram_cell_6t_5 inst_cell_126_66 (.BL(BL66),.BLN(BLN66),.WL(WL126));
sram_cell_6t_5 inst_cell_126_67 (.BL(BL67),.BLN(BLN67),.WL(WL126));
sram_cell_6t_5 inst_cell_126_68 (.BL(BL68),.BLN(BLN68),.WL(WL126));
sram_cell_6t_5 inst_cell_126_69 (.BL(BL69),.BLN(BLN69),.WL(WL126));
sram_cell_6t_5 inst_cell_126_70 (.BL(BL70),.BLN(BLN70),.WL(WL126));
sram_cell_6t_5 inst_cell_126_71 (.BL(BL71),.BLN(BLN71),.WL(WL126));
sram_cell_6t_5 inst_cell_126_72 (.BL(BL72),.BLN(BLN72),.WL(WL126));
sram_cell_6t_5 inst_cell_126_73 (.BL(BL73),.BLN(BLN73),.WL(WL126));
sram_cell_6t_5 inst_cell_126_74 (.BL(BL74),.BLN(BLN74),.WL(WL126));
sram_cell_6t_5 inst_cell_126_75 (.BL(BL75),.BLN(BLN75),.WL(WL126));
sram_cell_6t_5 inst_cell_126_76 (.BL(BL76),.BLN(BLN76),.WL(WL126));
sram_cell_6t_5 inst_cell_126_77 (.BL(BL77),.BLN(BLN77),.WL(WL126));
sram_cell_6t_5 inst_cell_126_78 (.BL(BL78),.BLN(BLN78),.WL(WL126));
sram_cell_6t_5 inst_cell_126_79 (.BL(BL79),.BLN(BLN79),.WL(WL126));
sram_cell_6t_5 inst_cell_126_80 (.BL(BL80),.BLN(BLN80),.WL(WL126));
sram_cell_6t_5 inst_cell_126_81 (.BL(BL81),.BLN(BLN81),.WL(WL126));
sram_cell_6t_5 inst_cell_126_82 (.BL(BL82),.BLN(BLN82),.WL(WL126));
sram_cell_6t_5 inst_cell_126_83 (.BL(BL83),.BLN(BLN83),.WL(WL126));
sram_cell_6t_5 inst_cell_126_84 (.BL(BL84),.BLN(BLN84),.WL(WL126));
sram_cell_6t_5 inst_cell_126_85 (.BL(BL85),.BLN(BLN85),.WL(WL126));
sram_cell_6t_5 inst_cell_126_86 (.BL(BL86),.BLN(BLN86),.WL(WL126));
sram_cell_6t_5 inst_cell_126_87 (.BL(BL87),.BLN(BLN87),.WL(WL126));
sram_cell_6t_5 inst_cell_126_88 (.BL(BL88),.BLN(BLN88),.WL(WL126));
sram_cell_6t_5 inst_cell_126_89 (.BL(BL89),.BLN(BLN89),.WL(WL126));
sram_cell_6t_5 inst_cell_126_90 (.BL(BL90),.BLN(BLN90),.WL(WL126));
sram_cell_6t_5 inst_cell_126_91 (.BL(BL91),.BLN(BLN91),.WL(WL126));
sram_cell_6t_5 inst_cell_126_92 (.BL(BL92),.BLN(BLN92),.WL(WL126));
sram_cell_6t_5 inst_cell_126_93 (.BL(BL93),.BLN(BLN93),.WL(WL126));
sram_cell_6t_5 inst_cell_126_94 (.BL(BL94),.BLN(BLN94),.WL(WL126));
sram_cell_6t_5 inst_cell_126_95 (.BL(BL95),.BLN(BLN95),.WL(WL126));
sram_cell_6t_5 inst_cell_126_96 (.BL(BL96),.BLN(BLN96),.WL(WL126));
sram_cell_6t_5 inst_cell_126_97 (.BL(BL97),.BLN(BLN97),.WL(WL126));
sram_cell_6t_5 inst_cell_126_98 (.BL(BL98),.BLN(BLN98),.WL(WL126));
sram_cell_6t_5 inst_cell_126_99 (.BL(BL99),.BLN(BLN99),.WL(WL126));
sram_cell_6t_5 inst_cell_126_100 (.BL(BL100),.BLN(BLN100),.WL(WL126));
sram_cell_6t_5 inst_cell_126_101 (.BL(BL101),.BLN(BLN101),.WL(WL126));
sram_cell_6t_5 inst_cell_126_102 (.BL(BL102),.BLN(BLN102),.WL(WL126));
sram_cell_6t_5 inst_cell_126_103 (.BL(BL103),.BLN(BLN103),.WL(WL126));
sram_cell_6t_5 inst_cell_126_104 (.BL(BL104),.BLN(BLN104),.WL(WL126));
sram_cell_6t_5 inst_cell_126_105 (.BL(BL105),.BLN(BLN105),.WL(WL126));
sram_cell_6t_5 inst_cell_126_106 (.BL(BL106),.BLN(BLN106),.WL(WL126));
sram_cell_6t_5 inst_cell_126_107 (.BL(BL107),.BLN(BLN107),.WL(WL126));
sram_cell_6t_5 inst_cell_126_108 (.BL(BL108),.BLN(BLN108),.WL(WL126));
sram_cell_6t_5 inst_cell_126_109 (.BL(BL109),.BLN(BLN109),.WL(WL126));
sram_cell_6t_5 inst_cell_126_110 (.BL(BL110),.BLN(BLN110),.WL(WL126));
sram_cell_6t_5 inst_cell_126_111 (.BL(BL111),.BLN(BLN111),.WL(WL126));
sram_cell_6t_5 inst_cell_126_112 (.BL(BL112),.BLN(BLN112),.WL(WL126));
sram_cell_6t_5 inst_cell_126_113 (.BL(BL113),.BLN(BLN113),.WL(WL126));
sram_cell_6t_5 inst_cell_126_114 (.BL(BL114),.BLN(BLN114),.WL(WL126));
sram_cell_6t_5 inst_cell_126_115 (.BL(BL115),.BLN(BLN115),.WL(WL126));
sram_cell_6t_5 inst_cell_126_116 (.BL(BL116),.BLN(BLN116),.WL(WL126));
sram_cell_6t_5 inst_cell_126_117 (.BL(BL117),.BLN(BLN117),.WL(WL126));
sram_cell_6t_5 inst_cell_126_118 (.BL(BL118),.BLN(BLN118),.WL(WL126));
sram_cell_6t_5 inst_cell_126_119 (.BL(BL119),.BLN(BLN119),.WL(WL126));
sram_cell_6t_5 inst_cell_126_120 (.BL(BL120),.BLN(BLN120),.WL(WL126));
sram_cell_6t_5 inst_cell_126_121 (.BL(BL121),.BLN(BLN121),.WL(WL126));
sram_cell_6t_5 inst_cell_126_122 (.BL(BL122),.BLN(BLN122),.WL(WL126));
sram_cell_6t_5 inst_cell_126_123 (.BL(BL123),.BLN(BLN123),.WL(WL126));
sram_cell_6t_5 inst_cell_126_124 (.BL(BL124),.BLN(BLN124),.WL(WL126));
sram_cell_6t_5 inst_cell_126_125 (.BL(BL125),.BLN(BLN125),.WL(WL126));
sram_cell_6t_5 inst_cell_126_126 (.BL(BL126),.BLN(BLN126),.WL(WL126));
sram_cell_6t_5 inst_cell_126_127 (.BL(BL127),.BLN(BLN127),.WL(WL126));
sram_cell_6t_5 inst_cell_127_0 (.BL(BL0),.BLN(BLN0),.WL(WL127));
sram_cell_6t_5 inst_cell_127_1 (.BL(BL1),.BLN(BLN1),.WL(WL127));
sram_cell_6t_5 inst_cell_127_2 (.BL(BL2),.BLN(BLN2),.WL(WL127));
sram_cell_6t_5 inst_cell_127_3 (.BL(BL3),.BLN(BLN3),.WL(WL127));
sram_cell_6t_5 inst_cell_127_4 (.BL(BL4),.BLN(BLN4),.WL(WL127));
sram_cell_6t_5 inst_cell_127_5 (.BL(BL5),.BLN(BLN5),.WL(WL127));
sram_cell_6t_5 inst_cell_127_6 (.BL(BL6),.BLN(BLN6),.WL(WL127));
sram_cell_6t_5 inst_cell_127_7 (.BL(BL7),.BLN(BLN7),.WL(WL127));
sram_cell_6t_5 inst_cell_127_8 (.BL(BL8),.BLN(BLN8),.WL(WL127));
sram_cell_6t_5 inst_cell_127_9 (.BL(BL9),.BLN(BLN9),.WL(WL127));
sram_cell_6t_5 inst_cell_127_10 (.BL(BL10),.BLN(BLN10),.WL(WL127));
sram_cell_6t_5 inst_cell_127_11 (.BL(BL11),.BLN(BLN11),.WL(WL127));
sram_cell_6t_5 inst_cell_127_12 (.BL(BL12),.BLN(BLN12),.WL(WL127));
sram_cell_6t_5 inst_cell_127_13 (.BL(BL13),.BLN(BLN13),.WL(WL127));
sram_cell_6t_5 inst_cell_127_14 (.BL(BL14),.BLN(BLN14),.WL(WL127));
sram_cell_6t_5 inst_cell_127_15 (.BL(BL15),.BLN(BLN15),.WL(WL127));
sram_cell_6t_5 inst_cell_127_16 (.BL(BL16),.BLN(BLN16),.WL(WL127));
sram_cell_6t_5 inst_cell_127_17 (.BL(BL17),.BLN(BLN17),.WL(WL127));
sram_cell_6t_5 inst_cell_127_18 (.BL(BL18),.BLN(BLN18),.WL(WL127));
sram_cell_6t_5 inst_cell_127_19 (.BL(BL19),.BLN(BLN19),.WL(WL127));
sram_cell_6t_5 inst_cell_127_20 (.BL(BL20),.BLN(BLN20),.WL(WL127));
sram_cell_6t_5 inst_cell_127_21 (.BL(BL21),.BLN(BLN21),.WL(WL127));
sram_cell_6t_5 inst_cell_127_22 (.BL(BL22),.BLN(BLN22),.WL(WL127));
sram_cell_6t_5 inst_cell_127_23 (.BL(BL23),.BLN(BLN23),.WL(WL127));
sram_cell_6t_5 inst_cell_127_24 (.BL(BL24),.BLN(BLN24),.WL(WL127));
sram_cell_6t_5 inst_cell_127_25 (.BL(BL25),.BLN(BLN25),.WL(WL127));
sram_cell_6t_5 inst_cell_127_26 (.BL(BL26),.BLN(BLN26),.WL(WL127));
sram_cell_6t_5 inst_cell_127_27 (.BL(BL27),.BLN(BLN27),.WL(WL127));
sram_cell_6t_5 inst_cell_127_28 (.BL(BL28),.BLN(BLN28),.WL(WL127));
sram_cell_6t_5 inst_cell_127_29 (.BL(BL29),.BLN(BLN29),.WL(WL127));
sram_cell_6t_5 inst_cell_127_30 (.BL(BL30),.BLN(BLN30),.WL(WL127));
sram_cell_6t_5 inst_cell_127_31 (.BL(BL31),.BLN(BLN31),.WL(WL127));
sram_cell_6t_5 inst_cell_127_32 (.BL(BL32),.BLN(BLN32),.WL(WL127));
sram_cell_6t_5 inst_cell_127_33 (.BL(BL33),.BLN(BLN33),.WL(WL127));
sram_cell_6t_5 inst_cell_127_34 (.BL(BL34),.BLN(BLN34),.WL(WL127));
sram_cell_6t_5 inst_cell_127_35 (.BL(BL35),.BLN(BLN35),.WL(WL127));
sram_cell_6t_5 inst_cell_127_36 (.BL(BL36),.BLN(BLN36),.WL(WL127));
sram_cell_6t_5 inst_cell_127_37 (.BL(BL37),.BLN(BLN37),.WL(WL127));
sram_cell_6t_5 inst_cell_127_38 (.BL(BL38),.BLN(BLN38),.WL(WL127));
sram_cell_6t_5 inst_cell_127_39 (.BL(BL39),.BLN(BLN39),.WL(WL127));
sram_cell_6t_5 inst_cell_127_40 (.BL(BL40),.BLN(BLN40),.WL(WL127));
sram_cell_6t_5 inst_cell_127_41 (.BL(BL41),.BLN(BLN41),.WL(WL127));
sram_cell_6t_5 inst_cell_127_42 (.BL(BL42),.BLN(BLN42),.WL(WL127));
sram_cell_6t_5 inst_cell_127_43 (.BL(BL43),.BLN(BLN43),.WL(WL127));
sram_cell_6t_5 inst_cell_127_44 (.BL(BL44),.BLN(BLN44),.WL(WL127));
sram_cell_6t_5 inst_cell_127_45 (.BL(BL45),.BLN(BLN45),.WL(WL127));
sram_cell_6t_5 inst_cell_127_46 (.BL(BL46),.BLN(BLN46),.WL(WL127));
sram_cell_6t_5 inst_cell_127_47 (.BL(BL47),.BLN(BLN47),.WL(WL127));
sram_cell_6t_5 inst_cell_127_48 (.BL(BL48),.BLN(BLN48),.WL(WL127));
sram_cell_6t_5 inst_cell_127_49 (.BL(BL49),.BLN(BLN49),.WL(WL127));
sram_cell_6t_5 inst_cell_127_50 (.BL(BL50),.BLN(BLN50),.WL(WL127));
sram_cell_6t_5 inst_cell_127_51 (.BL(BL51),.BLN(BLN51),.WL(WL127));
sram_cell_6t_5 inst_cell_127_52 (.BL(BL52),.BLN(BLN52),.WL(WL127));
sram_cell_6t_5 inst_cell_127_53 (.BL(BL53),.BLN(BLN53),.WL(WL127));
sram_cell_6t_5 inst_cell_127_54 (.BL(BL54),.BLN(BLN54),.WL(WL127));
sram_cell_6t_5 inst_cell_127_55 (.BL(BL55),.BLN(BLN55),.WL(WL127));
sram_cell_6t_5 inst_cell_127_56 (.BL(BL56),.BLN(BLN56),.WL(WL127));
sram_cell_6t_5 inst_cell_127_57 (.BL(BL57),.BLN(BLN57),.WL(WL127));
sram_cell_6t_5 inst_cell_127_58 (.BL(BL58),.BLN(BLN58),.WL(WL127));
sram_cell_6t_5 inst_cell_127_59 (.BL(BL59),.BLN(BLN59),.WL(WL127));
sram_cell_6t_5 inst_cell_127_60 (.BL(BL60),.BLN(BLN60),.WL(WL127));
sram_cell_6t_5 inst_cell_127_61 (.BL(BL61),.BLN(BLN61),.WL(WL127));
sram_cell_6t_5 inst_cell_127_62 (.BL(BL62),.BLN(BLN62),.WL(WL127));
sram_cell_6t_5 inst_cell_127_63 (.BL(BL63),.BLN(BLN63),.WL(WL127));
sram_cell_6t_5 inst_cell_127_64 (.BL(BL64),.BLN(BLN64),.WL(WL127));
sram_cell_6t_5 inst_cell_127_65 (.BL(BL65),.BLN(BLN65),.WL(WL127));
sram_cell_6t_5 inst_cell_127_66 (.BL(BL66),.BLN(BLN66),.WL(WL127));
sram_cell_6t_5 inst_cell_127_67 (.BL(BL67),.BLN(BLN67),.WL(WL127));
sram_cell_6t_5 inst_cell_127_68 (.BL(BL68),.BLN(BLN68),.WL(WL127));
sram_cell_6t_5 inst_cell_127_69 (.BL(BL69),.BLN(BLN69),.WL(WL127));
sram_cell_6t_5 inst_cell_127_70 (.BL(BL70),.BLN(BLN70),.WL(WL127));
sram_cell_6t_5 inst_cell_127_71 (.BL(BL71),.BLN(BLN71),.WL(WL127));
sram_cell_6t_5 inst_cell_127_72 (.BL(BL72),.BLN(BLN72),.WL(WL127));
sram_cell_6t_5 inst_cell_127_73 (.BL(BL73),.BLN(BLN73),.WL(WL127));
sram_cell_6t_5 inst_cell_127_74 (.BL(BL74),.BLN(BLN74),.WL(WL127));
sram_cell_6t_5 inst_cell_127_75 (.BL(BL75),.BLN(BLN75),.WL(WL127));
sram_cell_6t_5 inst_cell_127_76 (.BL(BL76),.BLN(BLN76),.WL(WL127));
sram_cell_6t_5 inst_cell_127_77 (.BL(BL77),.BLN(BLN77),.WL(WL127));
sram_cell_6t_5 inst_cell_127_78 (.BL(BL78),.BLN(BLN78),.WL(WL127));
sram_cell_6t_5 inst_cell_127_79 (.BL(BL79),.BLN(BLN79),.WL(WL127));
sram_cell_6t_5 inst_cell_127_80 (.BL(BL80),.BLN(BLN80),.WL(WL127));
sram_cell_6t_5 inst_cell_127_81 (.BL(BL81),.BLN(BLN81),.WL(WL127));
sram_cell_6t_5 inst_cell_127_82 (.BL(BL82),.BLN(BLN82),.WL(WL127));
sram_cell_6t_5 inst_cell_127_83 (.BL(BL83),.BLN(BLN83),.WL(WL127));
sram_cell_6t_5 inst_cell_127_84 (.BL(BL84),.BLN(BLN84),.WL(WL127));
sram_cell_6t_5 inst_cell_127_85 (.BL(BL85),.BLN(BLN85),.WL(WL127));
sram_cell_6t_5 inst_cell_127_86 (.BL(BL86),.BLN(BLN86),.WL(WL127));
sram_cell_6t_5 inst_cell_127_87 (.BL(BL87),.BLN(BLN87),.WL(WL127));
sram_cell_6t_5 inst_cell_127_88 (.BL(BL88),.BLN(BLN88),.WL(WL127));
sram_cell_6t_5 inst_cell_127_89 (.BL(BL89),.BLN(BLN89),.WL(WL127));
sram_cell_6t_5 inst_cell_127_90 (.BL(BL90),.BLN(BLN90),.WL(WL127));
sram_cell_6t_5 inst_cell_127_91 (.BL(BL91),.BLN(BLN91),.WL(WL127));
sram_cell_6t_5 inst_cell_127_92 (.BL(BL92),.BLN(BLN92),.WL(WL127));
sram_cell_6t_5 inst_cell_127_93 (.BL(BL93),.BLN(BLN93),.WL(WL127));
sram_cell_6t_5 inst_cell_127_94 (.BL(BL94),.BLN(BLN94),.WL(WL127));
sram_cell_6t_5 inst_cell_127_95 (.BL(BL95),.BLN(BLN95),.WL(WL127));
sram_cell_6t_5 inst_cell_127_96 (.BL(BL96),.BLN(BLN96),.WL(WL127));
sram_cell_6t_5 inst_cell_127_97 (.BL(BL97),.BLN(BLN97),.WL(WL127));
sram_cell_6t_5 inst_cell_127_98 (.BL(BL98),.BLN(BLN98),.WL(WL127));
sram_cell_6t_5 inst_cell_127_99 (.BL(BL99),.BLN(BLN99),.WL(WL127));
sram_cell_6t_5 inst_cell_127_100 (.BL(BL100),.BLN(BLN100),.WL(WL127));
sram_cell_6t_5 inst_cell_127_101 (.BL(BL101),.BLN(BLN101),.WL(WL127));
sram_cell_6t_5 inst_cell_127_102 (.BL(BL102),.BLN(BLN102),.WL(WL127));
sram_cell_6t_5 inst_cell_127_103 (.BL(BL103),.BLN(BLN103),.WL(WL127));
sram_cell_6t_5 inst_cell_127_104 (.BL(BL104),.BLN(BLN104),.WL(WL127));
sram_cell_6t_5 inst_cell_127_105 (.BL(BL105),.BLN(BLN105),.WL(WL127));
sram_cell_6t_5 inst_cell_127_106 (.BL(BL106),.BLN(BLN106),.WL(WL127));
sram_cell_6t_5 inst_cell_127_107 (.BL(BL107),.BLN(BLN107),.WL(WL127));
sram_cell_6t_5 inst_cell_127_108 (.BL(BL108),.BLN(BLN108),.WL(WL127));
sram_cell_6t_5 inst_cell_127_109 (.BL(BL109),.BLN(BLN109),.WL(WL127));
sram_cell_6t_5 inst_cell_127_110 (.BL(BL110),.BLN(BLN110),.WL(WL127));
sram_cell_6t_5 inst_cell_127_111 (.BL(BL111),.BLN(BLN111),.WL(WL127));
sram_cell_6t_5 inst_cell_127_112 (.BL(BL112),.BLN(BLN112),.WL(WL127));
sram_cell_6t_5 inst_cell_127_113 (.BL(BL113),.BLN(BLN113),.WL(WL127));
sram_cell_6t_5 inst_cell_127_114 (.BL(BL114),.BLN(BLN114),.WL(WL127));
sram_cell_6t_5 inst_cell_127_115 (.BL(BL115),.BLN(BLN115),.WL(WL127));
sram_cell_6t_5 inst_cell_127_116 (.BL(BL116),.BLN(BLN116),.WL(WL127));
sram_cell_6t_5 inst_cell_127_117 (.BL(BL117),.BLN(BLN117),.WL(WL127));
sram_cell_6t_5 inst_cell_127_118 (.BL(BL118),.BLN(BLN118),.WL(WL127));
sram_cell_6t_5 inst_cell_127_119 (.BL(BL119),.BLN(BLN119),.WL(WL127));
sram_cell_6t_5 inst_cell_127_120 (.BL(BL120),.BLN(BLN120),.WL(WL127));
sram_cell_6t_5 inst_cell_127_121 (.BL(BL121),.BLN(BLN121),.WL(WL127));
sram_cell_6t_5 inst_cell_127_122 (.BL(BL122),.BLN(BLN122),.WL(WL127));
sram_cell_6t_5 inst_cell_127_123 (.BL(BL123),.BLN(BLN123),.WL(WL127));
sram_cell_6t_5 inst_cell_127_124 (.BL(BL124),.BLN(BLN124),.WL(WL127));
sram_cell_6t_5 inst_cell_127_125 (.BL(BL125),.BLN(BLN125),.WL(WL127));
sram_cell_6t_5 inst_cell_127_126 (.BL(BL126),.BLN(BLN126),.WL(WL127));
sram_cell_6t_5 inst_cell_127_127 (.BL(BL127),.BLN(BLN127),.WL(WL127));
sram_cell_6t_5 inst_cell_128_0 (.BL(BL0),.BLN(BLN0),.WL(WL128));
sram_cell_6t_5 inst_cell_128_1 (.BL(BL1),.BLN(BLN1),.WL(WL128));
sram_cell_6t_5 inst_cell_128_2 (.BL(BL2),.BLN(BLN2),.WL(WL128));
sram_cell_6t_5 inst_cell_128_3 (.BL(BL3),.BLN(BLN3),.WL(WL128));
sram_cell_6t_5 inst_cell_128_4 (.BL(BL4),.BLN(BLN4),.WL(WL128));
sram_cell_6t_5 inst_cell_128_5 (.BL(BL5),.BLN(BLN5),.WL(WL128));
sram_cell_6t_5 inst_cell_128_6 (.BL(BL6),.BLN(BLN6),.WL(WL128));
sram_cell_6t_5 inst_cell_128_7 (.BL(BL7),.BLN(BLN7),.WL(WL128));
sram_cell_6t_5 inst_cell_128_8 (.BL(BL8),.BLN(BLN8),.WL(WL128));
sram_cell_6t_5 inst_cell_128_9 (.BL(BL9),.BLN(BLN9),.WL(WL128));
sram_cell_6t_5 inst_cell_128_10 (.BL(BL10),.BLN(BLN10),.WL(WL128));
sram_cell_6t_5 inst_cell_128_11 (.BL(BL11),.BLN(BLN11),.WL(WL128));
sram_cell_6t_5 inst_cell_128_12 (.BL(BL12),.BLN(BLN12),.WL(WL128));
sram_cell_6t_5 inst_cell_128_13 (.BL(BL13),.BLN(BLN13),.WL(WL128));
sram_cell_6t_5 inst_cell_128_14 (.BL(BL14),.BLN(BLN14),.WL(WL128));
sram_cell_6t_5 inst_cell_128_15 (.BL(BL15),.BLN(BLN15),.WL(WL128));
sram_cell_6t_5 inst_cell_128_16 (.BL(BL16),.BLN(BLN16),.WL(WL128));
sram_cell_6t_5 inst_cell_128_17 (.BL(BL17),.BLN(BLN17),.WL(WL128));
sram_cell_6t_5 inst_cell_128_18 (.BL(BL18),.BLN(BLN18),.WL(WL128));
sram_cell_6t_5 inst_cell_128_19 (.BL(BL19),.BLN(BLN19),.WL(WL128));
sram_cell_6t_5 inst_cell_128_20 (.BL(BL20),.BLN(BLN20),.WL(WL128));
sram_cell_6t_5 inst_cell_128_21 (.BL(BL21),.BLN(BLN21),.WL(WL128));
sram_cell_6t_5 inst_cell_128_22 (.BL(BL22),.BLN(BLN22),.WL(WL128));
sram_cell_6t_5 inst_cell_128_23 (.BL(BL23),.BLN(BLN23),.WL(WL128));
sram_cell_6t_5 inst_cell_128_24 (.BL(BL24),.BLN(BLN24),.WL(WL128));
sram_cell_6t_5 inst_cell_128_25 (.BL(BL25),.BLN(BLN25),.WL(WL128));
sram_cell_6t_5 inst_cell_128_26 (.BL(BL26),.BLN(BLN26),.WL(WL128));
sram_cell_6t_5 inst_cell_128_27 (.BL(BL27),.BLN(BLN27),.WL(WL128));
sram_cell_6t_5 inst_cell_128_28 (.BL(BL28),.BLN(BLN28),.WL(WL128));
sram_cell_6t_5 inst_cell_128_29 (.BL(BL29),.BLN(BLN29),.WL(WL128));
sram_cell_6t_5 inst_cell_128_30 (.BL(BL30),.BLN(BLN30),.WL(WL128));
sram_cell_6t_5 inst_cell_128_31 (.BL(BL31),.BLN(BLN31),.WL(WL128));
sram_cell_6t_5 inst_cell_128_32 (.BL(BL32),.BLN(BLN32),.WL(WL128));
sram_cell_6t_5 inst_cell_128_33 (.BL(BL33),.BLN(BLN33),.WL(WL128));
sram_cell_6t_5 inst_cell_128_34 (.BL(BL34),.BLN(BLN34),.WL(WL128));
sram_cell_6t_5 inst_cell_128_35 (.BL(BL35),.BLN(BLN35),.WL(WL128));
sram_cell_6t_5 inst_cell_128_36 (.BL(BL36),.BLN(BLN36),.WL(WL128));
sram_cell_6t_5 inst_cell_128_37 (.BL(BL37),.BLN(BLN37),.WL(WL128));
sram_cell_6t_5 inst_cell_128_38 (.BL(BL38),.BLN(BLN38),.WL(WL128));
sram_cell_6t_5 inst_cell_128_39 (.BL(BL39),.BLN(BLN39),.WL(WL128));
sram_cell_6t_5 inst_cell_128_40 (.BL(BL40),.BLN(BLN40),.WL(WL128));
sram_cell_6t_5 inst_cell_128_41 (.BL(BL41),.BLN(BLN41),.WL(WL128));
sram_cell_6t_5 inst_cell_128_42 (.BL(BL42),.BLN(BLN42),.WL(WL128));
sram_cell_6t_5 inst_cell_128_43 (.BL(BL43),.BLN(BLN43),.WL(WL128));
sram_cell_6t_5 inst_cell_128_44 (.BL(BL44),.BLN(BLN44),.WL(WL128));
sram_cell_6t_5 inst_cell_128_45 (.BL(BL45),.BLN(BLN45),.WL(WL128));
sram_cell_6t_5 inst_cell_128_46 (.BL(BL46),.BLN(BLN46),.WL(WL128));
sram_cell_6t_5 inst_cell_128_47 (.BL(BL47),.BLN(BLN47),.WL(WL128));
sram_cell_6t_5 inst_cell_128_48 (.BL(BL48),.BLN(BLN48),.WL(WL128));
sram_cell_6t_5 inst_cell_128_49 (.BL(BL49),.BLN(BLN49),.WL(WL128));
sram_cell_6t_5 inst_cell_128_50 (.BL(BL50),.BLN(BLN50),.WL(WL128));
sram_cell_6t_5 inst_cell_128_51 (.BL(BL51),.BLN(BLN51),.WL(WL128));
sram_cell_6t_5 inst_cell_128_52 (.BL(BL52),.BLN(BLN52),.WL(WL128));
sram_cell_6t_5 inst_cell_128_53 (.BL(BL53),.BLN(BLN53),.WL(WL128));
sram_cell_6t_5 inst_cell_128_54 (.BL(BL54),.BLN(BLN54),.WL(WL128));
sram_cell_6t_5 inst_cell_128_55 (.BL(BL55),.BLN(BLN55),.WL(WL128));
sram_cell_6t_5 inst_cell_128_56 (.BL(BL56),.BLN(BLN56),.WL(WL128));
sram_cell_6t_5 inst_cell_128_57 (.BL(BL57),.BLN(BLN57),.WL(WL128));
sram_cell_6t_5 inst_cell_128_58 (.BL(BL58),.BLN(BLN58),.WL(WL128));
sram_cell_6t_5 inst_cell_128_59 (.BL(BL59),.BLN(BLN59),.WL(WL128));
sram_cell_6t_5 inst_cell_128_60 (.BL(BL60),.BLN(BLN60),.WL(WL128));
sram_cell_6t_5 inst_cell_128_61 (.BL(BL61),.BLN(BLN61),.WL(WL128));
sram_cell_6t_5 inst_cell_128_62 (.BL(BL62),.BLN(BLN62),.WL(WL128));
sram_cell_6t_5 inst_cell_128_63 (.BL(BL63),.BLN(BLN63),.WL(WL128));
sram_cell_6t_5 inst_cell_128_64 (.BL(BL64),.BLN(BLN64),.WL(WL128));
sram_cell_6t_5 inst_cell_128_65 (.BL(BL65),.BLN(BLN65),.WL(WL128));
sram_cell_6t_5 inst_cell_128_66 (.BL(BL66),.BLN(BLN66),.WL(WL128));
sram_cell_6t_5 inst_cell_128_67 (.BL(BL67),.BLN(BLN67),.WL(WL128));
sram_cell_6t_5 inst_cell_128_68 (.BL(BL68),.BLN(BLN68),.WL(WL128));
sram_cell_6t_5 inst_cell_128_69 (.BL(BL69),.BLN(BLN69),.WL(WL128));
sram_cell_6t_5 inst_cell_128_70 (.BL(BL70),.BLN(BLN70),.WL(WL128));
sram_cell_6t_5 inst_cell_128_71 (.BL(BL71),.BLN(BLN71),.WL(WL128));
sram_cell_6t_5 inst_cell_128_72 (.BL(BL72),.BLN(BLN72),.WL(WL128));
sram_cell_6t_5 inst_cell_128_73 (.BL(BL73),.BLN(BLN73),.WL(WL128));
sram_cell_6t_5 inst_cell_128_74 (.BL(BL74),.BLN(BLN74),.WL(WL128));
sram_cell_6t_5 inst_cell_128_75 (.BL(BL75),.BLN(BLN75),.WL(WL128));
sram_cell_6t_5 inst_cell_128_76 (.BL(BL76),.BLN(BLN76),.WL(WL128));
sram_cell_6t_5 inst_cell_128_77 (.BL(BL77),.BLN(BLN77),.WL(WL128));
sram_cell_6t_5 inst_cell_128_78 (.BL(BL78),.BLN(BLN78),.WL(WL128));
sram_cell_6t_5 inst_cell_128_79 (.BL(BL79),.BLN(BLN79),.WL(WL128));
sram_cell_6t_5 inst_cell_128_80 (.BL(BL80),.BLN(BLN80),.WL(WL128));
sram_cell_6t_5 inst_cell_128_81 (.BL(BL81),.BLN(BLN81),.WL(WL128));
sram_cell_6t_5 inst_cell_128_82 (.BL(BL82),.BLN(BLN82),.WL(WL128));
sram_cell_6t_5 inst_cell_128_83 (.BL(BL83),.BLN(BLN83),.WL(WL128));
sram_cell_6t_5 inst_cell_128_84 (.BL(BL84),.BLN(BLN84),.WL(WL128));
sram_cell_6t_5 inst_cell_128_85 (.BL(BL85),.BLN(BLN85),.WL(WL128));
sram_cell_6t_5 inst_cell_128_86 (.BL(BL86),.BLN(BLN86),.WL(WL128));
sram_cell_6t_5 inst_cell_128_87 (.BL(BL87),.BLN(BLN87),.WL(WL128));
sram_cell_6t_5 inst_cell_128_88 (.BL(BL88),.BLN(BLN88),.WL(WL128));
sram_cell_6t_5 inst_cell_128_89 (.BL(BL89),.BLN(BLN89),.WL(WL128));
sram_cell_6t_5 inst_cell_128_90 (.BL(BL90),.BLN(BLN90),.WL(WL128));
sram_cell_6t_5 inst_cell_128_91 (.BL(BL91),.BLN(BLN91),.WL(WL128));
sram_cell_6t_5 inst_cell_128_92 (.BL(BL92),.BLN(BLN92),.WL(WL128));
sram_cell_6t_5 inst_cell_128_93 (.BL(BL93),.BLN(BLN93),.WL(WL128));
sram_cell_6t_5 inst_cell_128_94 (.BL(BL94),.BLN(BLN94),.WL(WL128));
sram_cell_6t_5 inst_cell_128_95 (.BL(BL95),.BLN(BLN95),.WL(WL128));
sram_cell_6t_5 inst_cell_128_96 (.BL(BL96),.BLN(BLN96),.WL(WL128));
sram_cell_6t_5 inst_cell_128_97 (.BL(BL97),.BLN(BLN97),.WL(WL128));
sram_cell_6t_5 inst_cell_128_98 (.BL(BL98),.BLN(BLN98),.WL(WL128));
sram_cell_6t_5 inst_cell_128_99 (.BL(BL99),.BLN(BLN99),.WL(WL128));
sram_cell_6t_5 inst_cell_128_100 (.BL(BL100),.BLN(BLN100),.WL(WL128));
sram_cell_6t_5 inst_cell_128_101 (.BL(BL101),.BLN(BLN101),.WL(WL128));
sram_cell_6t_5 inst_cell_128_102 (.BL(BL102),.BLN(BLN102),.WL(WL128));
sram_cell_6t_5 inst_cell_128_103 (.BL(BL103),.BLN(BLN103),.WL(WL128));
sram_cell_6t_5 inst_cell_128_104 (.BL(BL104),.BLN(BLN104),.WL(WL128));
sram_cell_6t_5 inst_cell_128_105 (.BL(BL105),.BLN(BLN105),.WL(WL128));
sram_cell_6t_5 inst_cell_128_106 (.BL(BL106),.BLN(BLN106),.WL(WL128));
sram_cell_6t_5 inst_cell_128_107 (.BL(BL107),.BLN(BLN107),.WL(WL128));
sram_cell_6t_5 inst_cell_128_108 (.BL(BL108),.BLN(BLN108),.WL(WL128));
sram_cell_6t_5 inst_cell_128_109 (.BL(BL109),.BLN(BLN109),.WL(WL128));
sram_cell_6t_5 inst_cell_128_110 (.BL(BL110),.BLN(BLN110),.WL(WL128));
sram_cell_6t_5 inst_cell_128_111 (.BL(BL111),.BLN(BLN111),.WL(WL128));
sram_cell_6t_5 inst_cell_128_112 (.BL(BL112),.BLN(BLN112),.WL(WL128));
sram_cell_6t_5 inst_cell_128_113 (.BL(BL113),.BLN(BLN113),.WL(WL128));
sram_cell_6t_5 inst_cell_128_114 (.BL(BL114),.BLN(BLN114),.WL(WL128));
sram_cell_6t_5 inst_cell_128_115 (.BL(BL115),.BLN(BLN115),.WL(WL128));
sram_cell_6t_5 inst_cell_128_116 (.BL(BL116),.BLN(BLN116),.WL(WL128));
sram_cell_6t_5 inst_cell_128_117 (.BL(BL117),.BLN(BLN117),.WL(WL128));
sram_cell_6t_5 inst_cell_128_118 (.BL(BL118),.BLN(BLN118),.WL(WL128));
sram_cell_6t_5 inst_cell_128_119 (.BL(BL119),.BLN(BLN119),.WL(WL128));
sram_cell_6t_5 inst_cell_128_120 (.BL(BL120),.BLN(BLN120),.WL(WL128));
sram_cell_6t_5 inst_cell_128_121 (.BL(BL121),.BLN(BLN121),.WL(WL128));
sram_cell_6t_5 inst_cell_128_122 (.BL(BL122),.BLN(BLN122),.WL(WL128));
sram_cell_6t_5 inst_cell_128_123 (.BL(BL123),.BLN(BLN123),.WL(WL128));
sram_cell_6t_5 inst_cell_128_124 (.BL(BL124),.BLN(BLN124),.WL(WL128));
sram_cell_6t_5 inst_cell_128_125 (.BL(BL125),.BLN(BLN125),.WL(WL128));
sram_cell_6t_5 inst_cell_128_126 (.BL(BL126),.BLN(BLN126),.WL(WL128));
sram_cell_6t_5 inst_cell_128_127 (.BL(BL127),.BLN(BLN127),.WL(WL128));
sram_cell_6t_5 inst_cell_129_0 (.BL(BL0),.BLN(BLN0),.WL(WL129));
sram_cell_6t_5 inst_cell_129_1 (.BL(BL1),.BLN(BLN1),.WL(WL129));
sram_cell_6t_5 inst_cell_129_2 (.BL(BL2),.BLN(BLN2),.WL(WL129));
sram_cell_6t_5 inst_cell_129_3 (.BL(BL3),.BLN(BLN3),.WL(WL129));
sram_cell_6t_5 inst_cell_129_4 (.BL(BL4),.BLN(BLN4),.WL(WL129));
sram_cell_6t_5 inst_cell_129_5 (.BL(BL5),.BLN(BLN5),.WL(WL129));
sram_cell_6t_5 inst_cell_129_6 (.BL(BL6),.BLN(BLN6),.WL(WL129));
sram_cell_6t_5 inst_cell_129_7 (.BL(BL7),.BLN(BLN7),.WL(WL129));
sram_cell_6t_5 inst_cell_129_8 (.BL(BL8),.BLN(BLN8),.WL(WL129));
sram_cell_6t_5 inst_cell_129_9 (.BL(BL9),.BLN(BLN9),.WL(WL129));
sram_cell_6t_5 inst_cell_129_10 (.BL(BL10),.BLN(BLN10),.WL(WL129));
sram_cell_6t_5 inst_cell_129_11 (.BL(BL11),.BLN(BLN11),.WL(WL129));
sram_cell_6t_5 inst_cell_129_12 (.BL(BL12),.BLN(BLN12),.WL(WL129));
sram_cell_6t_5 inst_cell_129_13 (.BL(BL13),.BLN(BLN13),.WL(WL129));
sram_cell_6t_5 inst_cell_129_14 (.BL(BL14),.BLN(BLN14),.WL(WL129));
sram_cell_6t_5 inst_cell_129_15 (.BL(BL15),.BLN(BLN15),.WL(WL129));
sram_cell_6t_5 inst_cell_129_16 (.BL(BL16),.BLN(BLN16),.WL(WL129));
sram_cell_6t_5 inst_cell_129_17 (.BL(BL17),.BLN(BLN17),.WL(WL129));
sram_cell_6t_5 inst_cell_129_18 (.BL(BL18),.BLN(BLN18),.WL(WL129));
sram_cell_6t_5 inst_cell_129_19 (.BL(BL19),.BLN(BLN19),.WL(WL129));
sram_cell_6t_5 inst_cell_129_20 (.BL(BL20),.BLN(BLN20),.WL(WL129));
sram_cell_6t_5 inst_cell_129_21 (.BL(BL21),.BLN(BLN21),.WL(WL129));
sram_cell_6t_5 inst_cell_129_22 (.BL(BL22),.BLN(BLN22),.WL(WL129));
sram_cell_6t_5 inst_cell_129_23 (.BL(BL23),.BLN(BLN23),.WL(WL129));
sram_cell_6t_5 inst_cell_129_24 (.BL(BL24),.BLN(BLN24),.WL(WL129));
sram_cell_6t_5 inst_cell_129_25 (.BL(BL25),.BLN(BLN25),.WL(WL129));
sram_cell_6t_5 inst_cell_129_26 (.BL(BL26),.BLN(BLN26),.WL(WL129));
sram_cell_6t_5 inst_cell_129_27 (.BL(BL27),.BLN(BLN27),.WL(WL129));
sram_cell_6t_5 inst_cell_129_28 (.BL(BL28),.BLN(BLN28),.WL(WL129));
sram_cell_6t_5 inst_cell_129_29 (.BL(BL29),.BLN(BLN29),.WL(WL129));
sram_cell_6t_5 inst_cell_129_30 (.BL(BL30),.BLN(BLN30),.WL(WL129));
sram_cell_6t_5 inst_cell_129_31 (.BL(BL31),.BLN(BLN31),.WL(WL129));
sram_cell_6t_5 inst_cell_129_32 (.BL(BL32),.BLN(BLN32),.WL(WL129));
sram_cell_6t_5 inst_cell_129_33 (.BL(BL33),.BLN(BLN33),.WL(WL129));
sram_cell_6t_5 inst_cell_129_34 (.BL(BL34),.BLN(BLN34),.WL(WL129));
sram_cell_6t_5 inst_cell_129_35 (.BL(BL35),.BLN(BLN35),.WL(WL129));
sram_cell_6t_5 inst_cell_129_36 (.BL(BL36),.BLN(BLN36),.WL(WL129));
sram_cell_6t_5 inst_cell_129_37 (.BL(BL37),.BLN(BLN37),.WL(WL129));
sram_cell_6t_5 inst_cell_129_38 (.BL(BL38),.BLN(BLN38),.WL(WL129));
sram_cell_6t_5 inst_cell_129_39 (.BL(BL39),.BLN(BLN39),.WL(WL129));
sram_cell_6t_5 inst_cell_129_40 (.BL(BL40),.BLN(BLN40),.WL(WL129));
sram_cell_6t_5 inst_cell_129_41 (.BL(BL41),.BLN(BLN41),.WL(WL129));
sram_cell_6t_5 inst_cell_129_42 (.BL(BL42),.BLN(BLN42),.WL(WL129));
sram_cell_6t_5 inst_cell_129_43 (.BL(BL43),.BLN(BLN43),.WL(WL129));
sram_cell_6t_5 inst_cell_129_44 (.BL(BL44),.BLN(BLN44),.WL(WL129));
sram_cell_6t_5 inst_cell_129_45 (.BL(BL45),.BLN(BLN45),.WL(WL129));
sram_cell_6t_5 inst_cell_129_46 (.BL(BL46),.BLN(BLN46),.WL(WL129));
sram_cell_6t_5 inst_cell_129_47 (.BL(BL47),.BLN(BLN47),.WL(WL129));
sram_cell_6t_5 inst_cell_129_48 (.BL(BL48),.BLN(BLN48),.WL(WL129));
sram_cell_6t_5 inst_cell_129_49 (.BL(BL49),.BLN(BLN49),.WL(WL129));
sram_cell_6t_5 inst_cell_129_50 (.BL(BL50),.BLN(BLN50),.WL(WL129));
sram_cell_6t_5 inst_cell_129_51 (.BL(BL51),.BLN(BLN51),.WL(WL129));
sram_cell_6t_5 inst_cell_129_52 (.BL(BL52),.BLN(BLN52),.WL(WL129));
sram_cell_6t_5 inst_cell_129_53 (.BL(BL53),.BLN(BLN53),.WL(WL129));
sram_cell_6t_5 inst_cell_129_54 (.BL(BL54),.BLN(BLN54),.WL(WL129));
sram_cell_6t_5 inst_cell_129_55 (.BL(BL55),.BLN(BLN55),.WL(WL129));
sram_cell_6t_5 inst_cell_129_56 (.BL(BL56),.BLN(BLN56),.WL(WL129));
sram_cell_6t_5 inst_cell_129_57 (.BL(BL57),.BLN(BLN57),.WL(WL129));
sram_cell_6t_5 inst_cell_129_58 (.BL(BL58),.BLN(BLN58),.WL(WL129));
sram_cell_6t_5 inst_cell_129_59 (.BL(BL59),.BLN(BLN59),.WL(WL129));
sram_cell_6t_5 inst_cell_129_60 (.BL(BL60),.BLN(BLN60),.WL(WL129));
sram_cell_6t_5 inst_cell_129_61 (.BL(BL61),.BLN(BLN61),.WL(WL129));
sram_cell_6t_5 inst_cell_129_62 (.BL(BL62),.BLN(BLN62),.WL(WL129));
sram_cell_6t_5 inst_cell_129_63 (.BL(BL63),.BLN(BLN63),.WL(WL129));
sram_cell_6t_5 inst_cell_129_64 (.BL(BL64),.BLN(BLN64),.WL(WL129));
sram_cell_6t_5 inst_cell_129_65 (.BL(BL65),.BLN(BLN65),.WL(WL129));
sram_cell_6t_5 inst_cell_129_66 (.BL(BL66),.BLN(BLN66),.WL(WL129));
sram_cell_6t_5 inst_cell_129_67 (.BL(BL67),.BLN(BLN67),.WL(WL129));
sram_cell_6t_5 inst_cell_129_68 (.BL(BL68),.BLN(BLN68),.WL(WL129));
sram_cell_6t_5 inst_cell_129_69 (.BL(BL69),.BLN(BLN69),.WL(WL129));
sram_cell_6t_5 inst_cell_129_70 (.BL(BL70),.BLN(BLN70),.WL(WL129));
sram_cell_6t_5 inst_cell_129_71 (.BL(BL71),.BLN(BLN71),.WL(WL129));
sram_cell_6t_5 inst_cell_129_72 (.BL(BL72),.BLN(BLN72),.WL(WL129));
sram_cell_6t_5 inst_cell_129_73 (.BL(BL73),.BLN(BLN73),.WL(WL129));
sram_cell_6t_5 inst_cell_129_74 (.BL(BL74),.BLN(BLN74),.WL(WL129));
sram_cell_6t_5 inst_cell_129_75 (.BL(BL75),.BLN(BLN75),.WL(WL129));
sram_cell_6t_5 inst_cell_129_76 (.BL(BL76),.BLN(BLN76),.WL(WL129));
sram_cell_6t_5 inst_cell_129_77 (.BL(BL77),.BLN(BLN77),.WL(WL129));
sram_cell_6t_5 inst_cell_129_78 (.BL(BL78),.BLN(BLN78),.WL(WL129));
sram_cell_6t_5 inst_cell_129_79 (.BL(BL79),.BLN(BLN79),.WL(WL129));
sram_cell_6t_5 inst_cell_129_80 (.BL(BL80),.BLN(BLN80),.WL(WL129));
sram_cell_6t_5 inst_cell_129_81 (.BL(BL81),.BLN(BLN81),.WL(WL129));
sram_cell_6t_5 inst_cell_129_82 (.BL(BL82),.BLN(BLN82),.WL(WL129));
sram_cell_6t_5 inst_cell_129_83 (.BL(BL83),.BLN(BLN83),.WL(WL129));
sram_cell_6t_5 inst_cell_129_84 (.BL(BL84),.BLN(BLN84),.WL(WL129));
sram_cell_6t_5 inst_cell_129_85 (.BL(BL85),.BLN(BLN85),.WL(WL129));
sram_cell_6t_5 inst_cell_129_86 (.BL(BL86),.BLN(BLN86),.WL(WL129));
sram_cell_6t_5 inst_cell_129_87 (.BL(BL87),.BLN(BLN87),.WL(WL129));
sram_cell_6t_5 inst_cell_129_88 (.BL(BL88),.BLN(BLN88),.WL(WL129));
sram_cell_6t_5 inst_cell_129_89 (.BL(BL89),.BLN(BLN89),.WL(WL129));
sram_cell_6t_5 inst_cell_129_90 (.BL(BL90),.BLN(BLN90),.WL(WL129));
sram_cell_6t_5 inst_cell_129_91 (.BL(BL91),.BLN(BLN91),.WL(WL129));
sram_cell_6t_5 inst_cell_129_92 (.BL(BL92),.BLN(BLN92),.WL(WL129));
sram_cell_6t_5 inst_cell_129_93 (.BL(BL93),.BLN(BLN93),.WL(WL129));
sram_cell_6t_5 inst_cell_129_94 (.BL(BL94),.BLN(BLN94),.WL(WL129));
sram_cell_6t_5 inst_cell_129_95 (.BL(BL95),.BLN(BLN95),.WL(WL129));
sram_cell_6t_5 inst_cell_129_96 (.BL(BL96),.BLN(BLN96),.WL(WL129));
sram_cell_6t_5 inst_cell_129_97 (.BL(BL97),.BLN(BLN97),.WL(WL129));
sram_cell_6t_5 inst_cell_129_98 (.BL(BL98),.BLN(BLN98),.WL(WL129));
sram_cell_6t_5 inst_cell_129_99 (.BL(BL99),.BLN(BLN99),.WL(WL129));
sram_cell_6t_5 inst_cell_129_100 (.BL(BL100),.BLN(BLN100),.WL(WL129));
sram_cell_6t_5 inst_cell_129_101 (.BL(BL101),.BLN(BLN101),.WL(WL129));
sram_cell_6t_5 inst_cell_129_102 (.BL(BL102),.BLN(BLN102),.WL(WL129));
sram_cell_6t_5 inst_cell_129_103 (.BL(BL103),.BLN(BLN103),.WL(WL129));
sram_cell_6t_5 inst_cell_129_104 (.BL(BL104),.BLN(BLN104),.WL(WL129));
sram_cell_6t_5 inst_cell_129_105 (.BL(BL105),.BLN(BLN105),.WL(WL129));
sram_cell_6t_5 inst_cell_129_106 (.BL(BL106),.BLN(BLN106),.WL(WL129));
sram_cell_6t_5 inst_cell_129_107 (.BL(BL107),.BLN(BLN107),.WL(WL129));
sram_cell_6t_5 inst_cell_129_108 (.BL(BL108),.BLN(BLN108),.WL(WL129));
sram_cell_6t_5 inst_cell_129_109 (.BL(BL109),.BLN(BLN109),.WL(WL129));
sram_cell_6t_5 inst_cell_129_110 (.BL(BL110),.BLN(BLN110),.WL(WL129));
sram_cell_6t_5 inst_cell_129_111 (.BL(BL111),.BLN(BLN111),.WL(WL129));
sram_cell_6t_5 inst_cell_129_112 (.BL(BL112),.BLN(BLN112),.WL(WL129));
sram_cell_6t_5 inst_cell_129_113 (.BL(BL113),.BLN(BLN113),.WL(WL129));
sram_cell_6t_5 inst_cell_129_114 (.BL(BL114),.BLN(BLN114),.WL(WL129));
sram_cell_6t_5 inst_cell_129_115 (.BL(BL115),.BLN(BLN115),.WL(WL129));
sram_cell_6t_5 inst_cell_129_116 (.BL(BL116),.BLN(BLN116),.WL(WL129));
sram_cell_6t_5 inst_cell_129_117 (.BL(BL117),.BLN(BLN117),.WL(WL129));
sram_cell_6t_5 inst_cell_129_118 (.BL(BL118),.BLN(BLN118),.WL(WL129));
sram_cell_6t_5 inst_cell_129_119 (.BL(BL119),.BLN(BLN119),.WL(WL129));
sram_cell_6t_5 inst_cell_129_120 (.BL(BL120),.BLN(BLN120),.WL(WL129));
sram_cell_6t_5 inst_cell_129_121 (.BL(BL121),.BLN(BLN121),.WL(WL129));
sram_cell_6t_5 inst_cell_129_122 (.BL(BL122),.BLN(BLN122),.WL(WL129));
sram_cell_6t_5 inst_cell_129_123 (.BL(BL123),.BLN(BLN123),.WL(WL129));
sram_cell_6t_5 inst_cell_129_124 (.BL(BL124),.BLN(BLN124),.WL(WL129));
sram_cell_6t_5 inst_cell_129_125 (.BL(BL125),.BLN(BLN125),.WL(WL129));
sram_cell_6t_5 inst_cell_129_126 (.BL(BL126),.BLN(BLN126),.WL(WL129));
sram_cell_6t_5 inst_cell_129_127 (.BL(BL127),.BLN(BLN127),.WL(WL129));
sram_cell_6t_5 inst_cell_130_0 (.BL(BL0),.BLN(BLN0),.WL(WL130));
sram_cell_6t_5 inst_cell_130_1 (.BL(BL1),.BLN(BLN1),.WL(WL130));
sram_cell_6t_5 inst_cell_130_2 (.BL(BL2),.BLN(BLN2),.WL(WL130));
sram_cell_6t_5 inst_cell_130_3 (.BL(BL3),.BLN(BLN3),.WL(WL130));
sram_cell_6t_5 inst_cell_130_4 (.BL(BL4),.BLN(BLN4),.WL(WL130));
sram_cell_6t_5 inst_cell_130_5 (.BL(BL5),.BLN(BLN5),.WL(WL130));
sram_cell_6t_5 inst_cell_130_6 (.BL(BL6),.BLN(BLN6),.WL(WL130));
sram_cell_6t_5 inst_cell_130_7 (.BL(BL7),.BLN(BLN7),.WL(WL130));
sram_cell_6t_5 inst_cell_130_8 (.BL(BL8),.BLN(BLN8),.WL(WL130));
sram_cell_6t_5 inst_cell_130_9 (.BL(BL9),.BLN(BLN9),.WL(WL130));
sram_cell_6t_5 inst_cell_130_10 (.BL(BL10),.BLN(BLN10),.WL(WL130));
sram_cell_6t_5 inst_cell_130_11 (.BL(BL11),.BLN(BLN11),.WL(WL130));
sram_cell_6t_5 inst_cell_130_12 (.BL(BL12),.BLN(BLN12),.WL(WL130));
sram_cell_6t_5 inst_cell_130_13 (.BL(BL13),.BLN(BLN13),.WL(WL130));
sram_cell_6t_5 inst_cell_130_14 (.BL(BL14),.BLN(BLN14),.WL(WL130));
sram_cell_6t_5 inst_cell_130_15 (.BL(BL15),.BLN(BLN15),.WL(WL130));
sram_cell_6t_5 inst_cell_130_16 (.BL(BL16),.BLN(BLN16),.WL(WL130));
sram_cell_6t_5 inst_cell_130_17 (.BL(BL17),.BLN(BLN17),.WL(WL130));
sram_cell_6t_5 inst_cell_130_18 (.BL(BL18),.BLN(BLN18),.WL(WL130));
sram_cell_6t_5 inst_cell_130_19 (.BL(BL19),.BLN(BLN19),.WL(WL130));
sram_cell_6t_5 inst_cell_130_20 (.BL(BL20),.BLN(BLN20),.WL(WL130));
sram_cell_6t_5 inst_cell_130_21 (.BL(BL21),.BLN(BLN21),.WL(WL130));
sram_cell_6t_5 inst_cell_130_22 (.BL(BL22),.BLN(BLN22),.WL(WL130));
sram_cell_6t_5 inst_cell_130_23 (.BL(BL23),.BLN(BLN23),.WL(WL130));
sram_cell_6t_5 inst_cell_130_24 (.BL(BL24),.BLN(BLN24),.WL(WL130));
sram_cell_6t_5 inst_cell_130_25 (.BL(BL25),.BLN(BLN25),.WL(WL130));
sram_cell_6t_5 inst_cell_130_26 (.BL(BL26),.BLN(BLN26),.WL(WL130));
sram_cell_6t_5 inst_cell_130_27 (.BL(BL27),.BLN(BLN27),.WL(WL130));
sram_cell_6t_5 inst_cell_130_28 (.BL(BL28),.BLN(BLN28),.WL(WL130));
sram_cell_6t_5 inst_cell_130_29 (.BL(BL29),.BLN(BLN29),.WL(WL130));
sram_cell_6t_5 inst_cell_130_30 (.BL(BL30),.BLN(BLN30),.WL(WL130));
sram_cell_6t_5 inst_cell_130_31 (.BL(BL31),.BLN(BLN31),.WL(WL130));
sram_cell_6t_5 inst_cell_130_32 (.BL(BL32),.BLN(BLN32),.WL(WL130));
sram_cell_6t_5 inst_cell_130_33 (.BL(BL33),.BLN(BLN33),.WL(WL130));
sram_cell_6t_5 inst_cell_130_34 (.BL(BL34),.BLN(BLN34),.WL(WL130));
sram_cell_6t_5 inst_cell_130_35 (.BL(BL35),.BLN(BLN35),.WL(WL130));
sram_cell_6t_5 inst_cell_130_36 (.BL(BL36),.BLN(BLN36),.WL(WL130));
sram_cell_6t_5 inst_cell_130_37 (.BL(BL37),.BLN(BLN37),.WL(WL130));
sram_cell_6t_5 inst_cell_130_38 (.BL(BL38),.BLN(BLN38),.WL(WL130));
sram_cell_6t_5 inst_cell_130_39 (.BL(BL39),.BLN(BLN39),.WL(WL130));
sram_cell_6t_5 inst_cell_130_40 (.BL(BL40),.BLN(BLN40),.WL(WL130));
sram_cell_6t_5 inst_cell_130_41 (.BL(BL41),.BLN(BLN41),.WL(WL130));
sram_cell_6t_5 inst_cell_130_42 (.BL(BL42),.BLN(BLN42),.WL(WL130));
sram_cell_6t_5 inst_cell_130_43 (.BL(BL43),.BLN(BLN43),.WL(WL130));
sram_cell_6t_5 inst_cell_130_44 (.BL(BL44),.BLN(BLN44),.WL(WL130));
sram_cell_6t_5 inst_cell_130_45 (.BL(BL45),.BLN(BLN45),.WL(WL130));
sram_cell_6t_5 inst_cell_130_46 (.BL(BL46),.BLN(BLN46),.WL(WL130));
sram_cell_6t_5 inst_cell_130_47 (.BL(BL47),.BLN(BLN47),.WL(WL130));
sram_cell_6t_5 inst_cell_130_48 (.BL(BL48),.BLN(BLN48),.WL(WL130));
sram_cell_6t_5 inst_cell_130_49 (.BL(BL49),.BLN(BLN49),.WL(WL130));
sram_cell_6t_5 inst_cell_130_50 (.BL(BL50),.BLN(BLN50),.WL(WL130));
sram_cell_6t_5 inst_cell_130_51 (.BL(BL51),.BLN(BLN51),.WL(WL130));
sram_cell_6t_5 inst_cell_130_52 (.BL(BL52),.BLN(BLN52),.WL(WL130));
sram_cell_6t_5 inst_cell_130_53 (.BL(BL53),.BLN(BLN53),.WL(WL130));
sram_cell_6t_5 inst_cell_130_54 (.BL(BL54),.BLN(BLN54),.WL(WL130));
sram_cell_6t_5 inst_cell_130_55 (.BL(BL55),.BLN(BLN55),.WL(WL130));
sram_cell_6t_5 inst_cell_130_56 (.BL(BL56),.BLN(BLN56),.WL(WL130));
sram_cell_6t_5 inst_cell_130_57 (.BL(BL57),.BLN(BLN57),.WL(WL130));
sram_cell_6t_5 inst_cell_130_58 (.BL(BL58),.BLN(BLN58),.WL(WL130));
sram_cell_6t_5 inst_cell_130_59 (.BL(BL59),.BLN(BLN59),.WL(WL130));
sram_cell_6t_5 inst_cell_130_60 (.BL(BL60),.BLN(BLN60),.WL(WL130));
sram_cell_6t_5 inst_cell_130_61 (.BL(BL61),.BLN(BLN61),.WL(WL130));
sram_cell_6t_5 inst_cell_130_62 (.BL(BL62),.BLN(BLN62),.WL(WL130));
sram_cell_6t_5 inst_cell_130_63 (.BL(BL63),.BLN(BLN63),.WL(WL130));
sram_cell_6t_5 inst_cell_130_64 (.BL(BL64),.BLN(BLN64),.WL(WL130));
sram_cell_6t_5 inst_cell_130_65 (.BL(BL65),.BLN(BLN65),.WL(WL130));
sram_cell_6t_5 inst_cell_130_66 (.BL(BL66),.BLN(BLN66),.WL(WL130));
sram_cell_6t_5 inst_cell_130_67 (.BL(BL67),.BLN(BLN67),.WL(WL130));
sram_cell_6t_5 inst_cell_130_68 (.BL(BL68),.BLN(BLN68),.WL(WL130));
sram_cell_6t_5 inst_cell_130_69 (.BL(BL69),.BLN(BLN69),.WL(WL130));
sram_cell_6t_5 inst_cell_130_70 (.BL(BL70),.BLN(BLN70),.WL(WL130));
sram_cell_6t_5 inst_cell_130_71 (.BL(BL71),.BLN(BLN71),.WL(WL130));
sram_cell_6t_5 inst_cell_130_72 (.BL(BL72),.BLN(BLN72),.WL(WL130));
sram_cell_6t_5 inst_cell_130_73 (.BL(BL73),.BLN(BLN73),.WL(WL130));
sram_cell_6t_5 inst_cell_130_74 (.BL(BL74),.BLN(BLN74),.WL(WL130));
sram_cell_6t_5 inst_cell_130_75 (.BL(BL75),.BLN(BLN75),.WL(WL130));
sram_cell_6t_5 inst_cell_130_76 (.BL(BL76),.BLN(BLN76),.WL(WL130));
sram_cell_6t_5 inst_cell_130_77 (.BL(BL77),.BLN(BLN77),.WL(WL130));
sram_cell_6t_5 inst_cell_130_78 (.BL(BL78),.BLN(BLN78),.WL(WL130));
sram_cell_6t_5 inst_cell_130_79 (.BL(BL79),.BLN(BLN79),.WL(WL130));
sram_cell_6t_5 inst_cell_130_80 (.BL(BL80),.BLN(BLN80),.WL(WL130));
sram_cell_6t_5 inst_cell_130_81 (.BL(BL81),.BLN(BLN81),.WL(WL130));
sram_cell_6t_5 inst_cell_130_82 (.BL(BL82),.BLN(BLN82),.WL(WL130));
sram_cell_6t_5 inst_cell_130_83 (.BL(BL83),.BLN(BLN83),.WL(WL130));
sram_cell_6t_5 inst_cell_130_84 (.BL(BL84),.BLN(BLN84),.WL(WL130));
sram_cell_6t_5 inst_cell_130_85 (.BL(BL85),.BLN(BLN85),.WL(WL130));
sram_cell_6t_5 inst_cell_130_86 (.BL(BL86),.BLN(BLN86),.WL(WL130));
sram_cell_6t_5 inst_cell_130_87 (.BL(BL87),.BLN(BLN87),.WL(WL130));
sram_cell_6t_5 inst_cell_130_88 (.BL(BL88),.BLN(BLN88),.WL(WL130));
sram_cell_6t_5 inst_cell_130_89 (.BL(BL89),.BLN(BLN89),.WL(WL130));
sram_cell_6t_5 inst_cell_130_90 (.BL(BL90),.BLN(BLN90),.WL(WL130));
sram_cell_6t_5 inst_cell_130_91 (.BL(BL91),.BLN(BLN91),.WL(WL130));
sram_cell_6t_5 inst_cell_130_92 (.BL(BL92),.BLN(BLN92),.WL(WL130));
sram_cell_6t_5 inst_cell_130_93 (.BL(BL93),.BLN(BLN93),.WL(WL130));
sram_cell_6t_5 inst_cell_130_94 (.BL(BL94),.BLN(BLN94),.WL(WL130));
sram_cell_6t_5 inst_cell_130_95 (.BL(BL95),.BLN(BLN95),.WL(WL130));
sram_cell_6t_5 inst_cell_130_96 (.BL(BL96),.BLN(BLN96),.WL(WL130));
sram_cell_6t_5 inst_cell_130_97 (.BL(BL97),.BLN(BLN97),.WL(WL130));
sram_cell_6t_5 inst_cell_130_98 (.BL(BL98),.BLN(BLN98),.WL(WL130));
sram_cell_6t_5 inst_cell_130_99 (.BL(BL99),.BLN(BLN99),.WL(WL130));
sram_cell_6t_5 inst_cell_130_100 (.BL(BL100),.BLN(BLN100),.WL(WL130));
sram_cell_6t_5 inst_cell_130_101 (.BL(BL101),.BLN(BLN101),.WL(WL130));
sram_cell_6t_5 inst_cell_130_102 (.BL(BL102),.BLN(BLN102),.WL(WL130));
sram_cell_6t_5 inst_cell_130_103 (.BL(BL103),.BLN(BLN103),.WL(WL130));
sram_cell_6t_5 inst_cell_130_104 (.BL(BL104),.BLN(BLN104),.WL(WL130));
sram_cell_6t_5 inst_cell_130_105 (.BL(BL105),.BLN(BLN105),.WL(WL130));
sram_cell_6t_5 inst_cell_130_106 (.BL(BL106),.BLN(BLN106),.WL(WL130));
sram_cell_6t_5 inst_cell_130_107 (.BL(BL107),.BLN(BLN107),.WL(WL130));
sram_cell_6t_5 inst_cell_130_108 (.BL(BL108),.BLN(BLN108),.WL(WL130));
sram_cell_6t_5 inst_cell_130_109 (.BL(BL109),.BLN(BLN109),.WL(WL130));
sram_cell_6t_5 inst_cell_130_110 (.BL(BL110),.BLN(BLN110),.WL(WL130));
sram_cell_6t_5 inst_cell_130_111 (.BL(BL111),.BLN(BLN111),.WL(WL130));
sram_cell_6t_5 inst_cell_130_112 (.BL(BL112),.BLN(BLN112),.WL(WL130));
sram_cell_6t_5 inst_cell_130_113 (.BL(BL113),.BLN(BLN113),.WL(WL130));
sram_cell_6t_5 inst_cell_130_114 (.BL(BL114),.BLN(BLN114),.WL(WL130));
sram_cell_6t_5 inst_cell_130_115 (.BL(BL115),.BLN(BLN115),.WL(WL130));
sram_cell_6t_5 inst_cell_130_116 (.BL(BL116),.BLN(BLN116),.WL(WL130));
sram_cell_6t_5 inst_cell_130_117 (.BL(BL117),.BLN(BLN117),.WL(WL130));
sram_cell_6t_5 inst_cell_130_118 (.BL(BL118),.BLN(BLN118),.WL(WL130));
sram_cell_6t_5 inst_cell_130_119 (.BL(BL119),.BLN(BLN119),.WL(WL130));
sram_cell_6t_5 inst_cell_130_120 (.BL(BL120),.BLN(BLN120),.WL(WL130));
sram_cell_6t_5 inst_cell_130_121 (.BL(BL121),.BLN(BLN121),.WL(WL130));
sram_cell_6t_5 inst_cell_130_122 (.BL(BL122),.BLN(BLN122),.WL(WL130));
sram_cell_6t_5 inst_cell_130_123 (.BL(BL123),.BLN(BLN123),.WL(WL130));
sram_cell_6t_5 inst_cell_130_124 (.BL(BL124),.BLN(BLN124),.WL(WL130));
sram_cell_6t_5 inst_cell_130_125 (.BL(BL125),.BLN(BLN125),.WL(WL130));
sram_cell_6t_5 inst_cell_130_126 (.BL(BL126),.BLN(BLN126),.WL(WL130));
sram_cell_6t_5 inst_cell_130_127 (.BL(BL127),.BLN(BLN127),.WL(WL130));
sram_cell_6t_5 inst_cell_131_0 (.BL(BL0),.BLN(BLN0),.WL(WL131));
sram_cell_6t_5 inst_cell_131_1 (.BL(BL1),.BLN(BLN1),.WL(WL131));
sram_cell_6t_5 inst_cell_131_2 (.BL(BL2),.BLN(BLN2),.WL(WL131));
sram_cell_6t_5 inst_cell_131_3 (.BL(BL3),.BLN(BLN3),.WL(WL131));
sram_cell_6t_5 inst_cell_131_4 (.BL(BL4),.BLN(BLN4),.WL(WL131));
sram_cell_6t_5 inst_cell_131_5 (.BL(BL5),.BLN(BLN5),.WL(WL131));
sram_cell_6t_5 inst_cell_131_6 (.BL(BL6),.BLN(BLN6),.WL(WL131));
sram_cell_6t_5 inst_cell_131_7 (.BL(BL7),.BLN(BLN7),.WL(WL131));
sram_cell_6t_5 inst_cell_131_8 (.BL(BL8),.BLN(BLN8),.WL(WL131));
sram_cell_6t_5 inst_cell_131_9 (.BL(BL9),.BLN(BLN9),.WL(WL131));
sram_cell_6t_5 inst_cell_131_10 (.BL(BL10),.BLN(BLN10),.WL(WL131));
sram_cell_6t_5 inst_cell_131_11 (.BL(BL11),.BLN(BLN11),.WL(WL131));
sram_cell_6t_5 inst_cell_131_12 (.BL(BL12),.BLN(BLN12),.WL(WL131));
sram_cell_6t_5 inst_cell_131_13 (.BL(BL13),.BLN(BLN13),.WL(WL131));
sram_cell_6t_5 inst_cell_131_14 (.BL(BL14),.BLN(BLN14),.WL(WL131));
sram_cell_6t_5 inst_cell_131_15 (.BL(BL15),.BLN(BLN15),.WL(WL131));
sram_cell_6t_5 inst_cell_131_16 (.BL(BL16),.BLN(BLN16),.WL(WL131));
sram_cell_6t_5 inst_cell_131_17 (.BL(BL17),.BLN(BLN17),.WL(WL131));
sram_cell_6t_5 inst_cell_131_18 (.BL(BL18),.BLN(BLN18),.WL(WL131));
sram_cell_6t_5 inst_cell_131_19 (.BL(BL19),.BLN(BLN19),.WL(WL131));
sram_cell_6t_5 inst_cell_131_20 (.BL(BL20),.BLN(BLN20),.WL(WL131));
sram_cell_6t_5 inst_cell_131_21 (.BL(BL21),.BLN(BLN21),.WL(WL131));
sram_cell_6t_5 inst_cell_131_22 (.BL(BL22),.BLN(BLN22),.WL(WL131));
sram_cell_6t_5 inst_cell_131_23 (.BL(BL23),.BLN(BLN23),.WL(WL131));
sram_cell_6t_5 inst_cell_131_24 (.BL(BL24),.BLN(BLN24),.WL(WL131));
sram_cell_6t_5 inst_cell_131_25 (.BL(BL25),.BLN(BLN25),.WL(WL131));
sram_cell_6t_5 inst_cell_131_26 (.BL(BL26),.BLN(BLN26),.WL(WL131));
sram_cell_6t_5 inst_cell_131_27 (.BL(BL27),.BLN(BLN27),.WL(WL131));
sram_cell_6t_5 inst_cell_131_28 (.BL(BL28),.BLN(BLN28),.WL(WL131));
sram_cell_6t_5 inst_cell_131_29 (.BL(BL29),.BLN(BLN29),.WL(WL131));
sram_cell_6t_5 inst_cell_131_30 (.BL(BL30),.BLN(BLN30),.WL(WL131));
sram_cell_6t_5 inst_cell_131_31 (.BL(BL31),.BLN(BLN31),.WL(WL131));
sram_cell_6t_5 inst_cell_131_32 (.BL(BL32),.BLN(BLN32),.WL(WL131));
sram_cell_6t_5 inst_cell_131_33 (.BL(BL33),.BLN(BLN33),.WL(WL131));
sram_cell_6t_5 inst_cell_131_34 (.BL(BL34),.BLN(BLN34),.WL(WL131));
sram_cell_6t_5 inst_cell_131_35 (.BL(BL35),.BLN(BLN35),.WL(WL131));
sram_cell_6t_5 inst_cell_131_36 (.BL(BL36),.BLN(BLN36),.WL(WL131));
sram_cell_6t_5 inst_cell_131_37 (.BL(BL37),.BLN(BLN37),.WL(WL131));
sram_cell_6t_5 inst_cell_131_38 (.BL(BL38),.BLN(BLN38),.WL(WL131));
sram_cell_6t_5 inst_cell_131_39 (.BL(BL39),.BLN(BLN39),.WL(WL131));
sram_cell_6t_5 inst_cell_131_40 (.BL(BL40),.BLN(BLN40),.WL(WL131));
sram_cell_6t_5 inst_cell_131_41 (.BL(BL41),.BLN(BLN41),.WL(WL131));
sram_cell_6t_5 inst_cell_131_42 (.BL(BL42),.BLN(BLN42),.WL(WL131));
sram_cell_6t_5 inst_cell_131_43 (.BL(BL43),.BLN(BLN43),.WL(WL131));
sram_cell_6t_5 inst_cell_131_44 (.BL(BL44),.BLN(BLN44),.WL(WL131));
sram_cell_6t_5 inst_cell_131_45 (.BL(BL45),.BLN(BLN45),.WL(WL131));
sram_cell_6t_5 inst_cell_131_46 (.BL(BL46),.BLN(BLN46),.WL(WL131));
sram_cell_6t_5 inst_cell_131_47 (.BL(BL47),.BLN(BLN47),.WL(WL131));
sram_cell_6t_5 inst_cell_131_48 (.BL(BL48),.BLN(BLN48),.WL(WL131));
sram_cell_6t_5 inst_cell_131_49 (.BL(BL49),.BLN(BLN49),.WL(WL131));
sram_cell_6t_5 inst_cell_131_50 (.BL(BL50),.BLN(BLN50),.WL(WL131));
sram_cell_6t_5 inst_cell_131_51 (.BL(BL51),.BLN(BLN51),.WL(WL131));
sram_cell_6t_5 inst_cell_131_52 (.BL(BL52),.BLN(BLN52),.WL(WL131));
sram_cell_6t_5 inst_cell_131_53 (.BL(BL53),.BLN(BLN53),.WL(WL131));
sram_cell_6t_5 inst_cell_131_54 (.BL(BL54),.BLN(BLN54),.WL(WL131));
sram_cell_6t_5 inst_cell_131_55 (.BL(BL55),.BLN(BLN55),.WL(WL131));
sram_cell_6t_5 inst_cell_131_56 (.BL(BL56),.BLN(BLN56),.WL(WL131));
sram_cell_6t_5 inst_cell_131_57 (.BL(BL57),.BLN(BLN57),.WL(WL131));
sram_cell_6t_5 inst_cell_131_58 (.BL(BL58),.BLN(BLN58),.WL(WL131));
sram_cell_6t_5 inst_cell_131_59 (.BL(BL59),.BLN(BLN59),.WL(WL131));
sram_cell_6t_5 inst_cell_131_60 (.BL(BL60),.BLN(BLN60),.WL(WL131));
sram_cell_6t_5 inst_cell_131_61 (.BL(BL61),.BLN(BLN61),.WL(WL131));
sram_cell_6t_5 inst_cell_131_62 (.BL(BL62),.BLN(BLN62),.WL(WL131));
sram_cell_6t_5 inst_cell_131_63 (.BL(BL63),.BLN(BLN63),.WL(WL131));
sram_cell_6t_5 inst_cell_131_64 (.BL(BL64),.BLN(BLN64),.WL(WL131));
sram_cell_6t_5 inst_cell_131_65 (.BL(BL65),.BLN(BLN65),.WL(WL131));
sram_cell_6t_5 inst_cell_131_66 (.BL(BL66),.BLN(BLN66),.WL(WL131));
sram_cell_6t_5 inst_cell_131_67 (.BL(BL67),.BLN(BLN67),.WL(WL131));
sram_cell_6t_5 inst_cell_131_68 (.BL(BL68),.BLN(BLN68),.WL(WL131));
sram_cell_6t_5 inst_cell_131_69 (.BL(BL69),.BLN(BLN69),.WL(WL131));
sram_cell_6t_5 inst_cell_131_70 (.BL(BL70),.BLN(BLN70),.WL(WL131));
sram_cell_6t_5 inst_cell_131_71 (.BL(BL71),.BLN(BLN71),.WL(WL131));
sram_cell_6t_5 inst_cell_131_72 (.BL(BL72),.BLN(BLN72),.WL(WL131));
sram_cell_6t_5 inst_cell_131_73 (.BL(BL73),.BLN(BLN73),.WL(WL131));
sram_cell_6t_5 inst_cell_131_74 (.BL(BL74),.BLN(BLN74),.WL(WL131));
sram_cell_6t_5 inst_cell_131_75 (.BL(BL75),.BLN(BLN75),.WL(WL131));
sram_cell_6t_5 inst_cell_131_76 (.BL(BL76),.BLN(BLN76),.WL(WL131));
sram_cell_6t_5 inst_cell_131_77 (.BL(BL77),.BLN(BLN77),.WL(WL131));
sram_cell_6t_5 inst_cell_131_78 (.BL(BL78),.BLN(BLN78),.WL(WL131));
sram_cell_6t_5 inst_cell_131_79 (.BL(BL79),.BLN(BLN79),.WL(WL131));
sram_cell_6t_5 inst_cell_131_80 (.BL(BL80),.BLN(BLN80),.WL(WL131));
sram_cell_6t_5 inst_cell_131_81 (.BL(BL81),.BLN(BLN81),.WL(WL131));
sram_cell_6t_5 inst_cell_131_82 (.BL(BL82),.BLN(BLN82),.WL(WL131));
sram_cell_6t_5 inst_cell_131_83 (.BL(BL83),.BLN(BLN83),.WL(WL131));
sram_cell_6t_5 inst_cell_131_84 (.BL(BL84),.BLN(BLN84),.WL(WL131));
sram_cell_6t_5 inst_cell_131_85 (.BL(BL85),.BLN(BLN85),.WL(WL131));
sram_cell_6t_5 inst_cell_131_86 (.BL(BL86),.BLN(BLN86),.WL(WL131));
sram_cell_6t_5 inst_cell_131_87 (.BL(BL87),.BLN(BLN87),.WL(WL131));
sram_cell_6t_5 inst_cell_131_88 (.BL(BL88),.BLN(BLN88),.WL(WL131));
sram_cell_6t_5 inst_cell_131_89 (.BL(BL89),.BLN(BLN89),.WL(WL131));
sram_cell_6t_5 inst_cell_131_90 (.BL(BL90),.BLN(BLN90),.WL(WL131));
sram_cell_6t_5 inst_cell_131_91 (.BL(BL91),.BLN(BLN91),.WL(WL131));
sram_cell_6t_5 inst_cell_131_92 (.BL(BL92),.BLN(BLN92),.WL(WL131));
sram_cell_6t_5 inst_cell_131_93 (.BL(BL93),.BLN(BLN93),.WL(WL131));
sram_cell_6t_5 inst_cell_131_94 (.BL(BL94),.BLN(BLN94),.WL(WL131));
sram_cell_6t_5 inst_cell_131_95 (.BL(BL95),.BLN(BLN95),.WL(WL131));
sram_cell_6t_5 inst_cell_131_96 (.BL(BL96),.BLN(BLN96),.WL(WL131));
sram_cell_6t_5 inst_cell_131_97 (.BL(BL97),.BLN(BLN97),.WL(WL131));
sram_cell_6t_5 inst_cell_131_98 (.BL(BL98),.BLN(BLN98),.WL(WL131));
sram_cell_6t_5 inst_cell_131_99 (.BL(BL99),.BLN(BLN99),.WL(WL131));
sram_cell_6t_5 inst_cell_131_100 (.BL(BL100),.BLN(BLN100),.WL(WL131));
sram_cell_6t_5 inst_cell_131_101 (.BL(BL101),.BLN(BLN101),.WL(WL131));
sram_cell_6t_5 inst_cell_131_102 (.BL(BL102),.BLN(BLN102),.WL(WL131));
sram_cell_6t_5 inst_cell_131_103 (.BL(BL103),.BLN(BLN103),.WL(WL131));
sram_cell_6t_5 inst_cell_131_104 (.BL(BL104),.BLN(BLN104),.WL(WL131));
sram_cell_6t_5 inst_cell_131_105 (.BL(BL105),.BLN(BLN105),.WL(WL131));
sram_cell_6t_5 inst_cell_131_106 (.BL(BL106),.BLN(BLN106),.WL(WL131));
sram_cell_6t_5 inst_cell_131_107 (.BL(BL107),.BLN(BLN107),.WL(WL131));
sram_cell_6t_5 inst_cell_131_108 (.BL(BL108),.BLN(BLN108),.WL(WL131));
sram_cell_6t_5 inst_cell_131_109 (.BL(BL109),.BLN(BLN109),.WL(WL131));
sram_cell_6t_5 inst_cell_131_110 (.BL(BL110),.BLN(BLN110),.WL(WL131));
sram_cell_6t_5 inst_cell_131_111 (.BL(BL111),.BLN(BLN111),.WL(WL131));
sram_cell_6t_5 inst_cell_131_112 (.BL(BL112),.BLN(BLN112),.WL(WL131));
sram_cell_6t_5 inst_cell_131_113 (.BL(BL113),.BLN(BLN113),.WL(WL131));
sram_cell_6t_5 inst_cell_131_114 (.BL(BL114),.BLN(BLN114),.WL(WL131));
sram_cell_6t_5 inst_cell_131_115 (.BL(BL115),.BLN(BLN115),.WL(WL131));
sram_cell_6t_5 inst_cell_131_116 (.BL(BL116),.BLN(BLN116),.WL(WL131));
sram_cell_6t_5 inst_cell_131_117 (.BL(BL117),.BLN(BLN117),.WL(WL131));
sram_cell_6t_5 inst_cell_131_118 (.BL(BL118),.BLN(BLN118),.WL(WL131));
sram_cell_6t_5 inst_cell_131_119 (.BL(BL119),.BLN(BLN119),.WL(WL131));
sram_cell_6t_5 inst_cell_131_120 (.BL(BL120),.BLN(BLN120),.WL(WL131));
sram_cell_6t_5 inst_cell_131_121 (.BL(BL121),.BLN(BLN121),.WL(WL131));
sram_cell_6t_5 inst_cell_131_122 (.BL(BL122),.BLN(BLN122),.WL(WL131));
sram_cell_6t_5 inst_cell_131_123 (.BL(BL123),.BLN(BLN123),.WL(WL131));
sram_cell_6t_5 inst_cell_131_124 (.BL(BL124),.BLN(BLN124),.WL(WL131));
sram_cell_6t_5 inst_cell_131_125 (.BL(BL125),.BLN(BLN125),.WL(WL131));
sram_cell_6t_5 inst_cell_131_126 (.BL(BL126),.BLN(BLN126),.WL(WL131));
sram_cell_6t_5 inst_cell_131_127 (.BL(BL127),.BLN(BLN127),.WL(WL131));
sram_cell_6t_5 inst_cell_132_0 (.BL(BL0),.BLN(BLN0),.WL(WL132));
sram_cell_6t_5 inst_cell_132_1 (.BL(BL1),.BLN(BLN1),.WL(WL132));
sram_cell_6t_5 inst_cell_132_2 (.BL(BL2),.BLN(BLN2),.WL(WL132));
sram_cell_6t_5 inst_cell_132_3 (.BL(BL3),.BLN(BLN3),.WL(WL132));
sram_cell_6t_5 inst_cell_132_4 (.BL(BL4),.BLN(BLN4),.WL(WL132));
sram_cell_6t_5 inst_cell_132_5 (.BL(BL5),.BLN(BLN5),.WL(WL132));
sram_cell_6t_5 inst_cell_132_6 (.BL(BL6),.BLN(BLN6),.WL(WL132));
sram_cell_6t_5 inst_cell_132_7 (.BL(BL7),.BLN(BLN7),.WL(WL132));
sram_cell_6t_5 inst_cell_132_8 (.BL(BL8),.BLN(BLN8),.WL(WL132));
sram_cell_6t_5 inst_cell_132_9 (.BL(BL9),.BLN(BLN9),.WL(WL132));
sram_cell_6t_5 inst_cell_132_10 (.BL(BL10),.BLN(BLN10),.WL(WL132));
sram_cell_6t_5 inst_cell_132_11 (.BL(BL11),.BLN(BLN11),.WL(WL132));
sram_cell_6t_5 inst_cell_132_12 (.BL(BL12),.BLN(BLN12),.WL(WL132));
sram_cell_6t_5 inst_cell_132_13 (.BL(BL13),.BLN(BLN13),.WL(WL132));
sram_cell_6t_5 inst_cell_132_14 (.BL(BL14),.BLN(BLN14),.WL(WL132));
sram_cell_6t_5 inst_cell_132_15 (.BL(BL15),.BLN(BLN15),.WL(WL132));
sram_cell_6t_5 inst_cell_132_16 (.BL(BL16),.BLN(BLN16),.WL(WL132));
sram_cell_6t_5 inst_cell_132_17 (.BL(BL17),.BLN(BLN17),.WL(WL132));
sram_cell_6t_5 inst_cell_132_18 (.BL(BL18),.BLN(BLN18),.WL(WL132));
sram_cell_6t_5 inst_cell_132_19 (.BL(BL19),.BLN(BLN19),.WL(WL132));
sram_cell_6t_5 inst_cell_132_20 (.BL(BL20),.BLN(BLN20),.WL(WL132));
sram_cell_6t_5 inst_cell_132_21 (.BL(BL21),.BLN(BLN21),.WL(WL132));
sram_cell_6t_5 inst_cell_132_22 (.BL(BL22),.BLN(BLN22),.WL(WL132));
sram_cell_6t_5 inst_cell_132_23 (.BL(BL23),.BLN(BLN23),.WL(WL132));
sram_cell_6t_5 inst_cell_132_24 (.BL(BL24),.BLN(BLN24),.WL(WL132));
sram_cell_6t_5 inst_cell_132_25 (.BL(BL25),.BLN(BLN25),.WL(WL132));
sram_cell_6t_5 inst_cell_132_26 (.BL(BL26),.BLN(BLN26),.WL(WL132));
sram_cell_6t_5 inst_cell_132_27 (.BL(BL27),.BLN(BLN27),.WL(WL132));
sram_cell_6t_5 inst_cell_132_28 (.BL(BL28),.BLN(BLN28),.WL(WL132));
sram_cell_6t_5 inst_cell_132_29 (.BL(BL29),.BLN(BLN29),.WL(WL132));
sram_cell_6t_5 inst_cell_132_30 (.BL(BL30),.BLN(BLN30),.WL(WL132));
sram_cell_6t_5 inst_cell_132_31 (.BL(BL31),.BLN(BLN31),.WL(WL132));
sram_cell_6t_5 inst_cell_132_32 (.BL(BL32),.BLN(BLN32),.WL(WL132));
sram_cell_6t_5 inst_cell_132_33 (.BL(BL33),.BLN(BLN33),.WL(WL132));
sram_cell_6t_5 inst_cell_132_34 (.BL(BL34),.BLN(BLN34),.WL(WL132));
sram_cell_6t_5 inst_cell_132_35 (.BL(BL35),.BLN(BLN35),.WL(WL132));
sram_cell_6t_5 inst_cell_132_36 (.BL(BL36),.BLN(BLN36),.WL(WL132));
sram_cell_6t_5 inst_cell_132_37 (.BL(BL37),.BLN(BLN37),.WL(WL132));
sram_cell_6t_5 inst_cell_132_38 (.BL(BL38),.BLN(BLN38),.WL(WL132));
sram_cell_6t_5 inst_cell_132_39 (.BL(BL39),.BLN(BLN39),.WL(WL132));
sram_cell_6t_5 inst_cell_132_40 (.BL(BL40),.BLN(BLN40),.WL(WL132));
sram_cell_6t_5 inst_cell_132_41 (.BL(BL41),.BLN(BLN41),.WL(WL132));
sram_cell_6t_5 inst_cell_132_42 (.BL(BL42),.BLN(BLN42),.WL(WL132));
sram_cell_6t_5 inst_cell_132_43 (.BL(BL43),.BLN(BLN43),.WL(WL132));
sram_cell_6t_5 inst_cell_132_44 (.BL(BL44),.BLN(BLN44),.WL(WL132));
sram_cell_6t_5 inst_cell_132_45 (.BL(BL45),.BLN(BLN45),.WL(WL132));
sram_cell_6t_5 inst_cell_132_46 (.BL(BL46),.BLN(BLN46),.WL(WL132));
sram_cell_6t_5 inst_cell_132_47 (.BL(BL47),.BLN(BLN47),.WL(WL132));
sram_cell_6t_5 inst_cell_132_48 (.BL(BL48),.BLN(BLN48),.WL(WL132));
sram_cell_6t_5 inst_cell_132_49 (.BL(BL49),.BLN(BLN49),.WL(WL132));
sram_cell_6t_5 inst_cell_132_50 (.BL(BL50),.BLN(BLN50),.WL(WL132));
sram_cell_6t_5 inst_cell_132_51 (.BL(BL51),.BLN(BLN51),.WL(WL132));
sram_cell_6t_5 inst_cell_132_52 (.BL(BL52),.BLN(BLN52),.WL(WL132));
sram_cell_6t_5 inst_cell_132_53 (.BL(BL53),.BLN(BLN53),.WL(WL132));
sram_cell_6t_5 inst_cell_132_54 (.BL(BL54),.BLN(BLN54),.WL(WL132));
sram_cell_6t_5 inst_cell_132_55 (.BL(BL55),.BLN(BLN55),.WL(WL132));
sram_cell_6t_5 inst_cell_132_56 (.BL(BL56),.BLN(BLN56),.WL(WL132));
sram_cell_6t_5 inst_cell_132_57 (.BL(BL57),.BLN(BLN57),.WL(WL132));
sram_cell_6t_5 inst_cell_132_58 (.BL(BL58),.BLN(BLN58),.WL(WL132));
sram_cell_6t_5 inst_cell_132_59 (.BL(BL59),.BLN(BLN59),.WL(WL132));
sram_cell_6t_5 inst_cell_132_60 (.BL(BL60),.BLN(BLN60),.WL(WL132));
sram_cell_6t_5 inst_cell_132_61 (.BL(BL61),.BLN(BLN61),.WL(WL132));
sram_cell_6t_5 inst_cell_132_62 (.BL(BL62),.BLN(BLN62),.WL(WL132));
sram_cell_6t_5 inst_cell_132_63 (.BL(BL63),.BLN(BLN63),.WL(WL132));
sram_cell_6t_5 inst_cell_132_64 (.BL(BL64),.BLN(BLN64),.WL(WL132));
sram_cell_6t_5 inst_cell_132_65 (.BL(BL65),.BLN(BLN65),.WL(WL132));
sram_cell_6t_5 inst_cell_132_66 (.BL(BL66),.BLN(BLN66),.WL(WL132));
sram_cell_6t_5 inst_cell_132_67 (.BL(BL67),.BLN(BLN67),.WL(WL132));
sram_cell_6t_5 inst_cell_132_68 (.BL(BL68),.BLN(BLN68),.WL(WL132));
sram_cell_6t_5 inst_cell_132_69 (.BL(BL69),.BLN(BLN69),.WL(WL132));
sram_cell_6t_5 inst_cell_132_70 (.BL(BL70),.BLN(BLN70),.WL(WL132));
sram_cell_6t_5 inst_cell_132_71 (.BL(BL71),.BLN(BLN71),.WL(WL132));
sram_cell_6t_5 inst_cell_132_72 (.BL(BL72),.BLN(BLN72),.WL(WL132));
sram_cell_6t_5 inst_cell_132_73 (.BL(BL73),.BLN(BLN73),.WL(WL132));
sram_cell_6t_5 inst_cell_132_74 (.BL(BL74),.BLN(BLN74),.WL(WL132));
sram_cell_6t_5 inst_cell_132_75 (.BL(BL75),.BLN(BLN75),.WL(WL132));
sram_cell_6t_5 inst_cell_132_76 (.BL(BL76),.BLN(BLN76),.WL(WL132));
sram_cell_6t_5 inst_cell_132_77 (.BL(BL77),.BLN(BLN77),.WL(WL132));
sram_cell_6t_5 inst_cell_132_78 (.BL(BL78),.BLN(BLN78),.WL(WL132));
sram_cell_6t_5 inst_cell_132_79 (.BL(BL79),.BLN(BLN79),.WL(WL132));
sram_cell_6t_5 inst_cell_132_80 (.BL(BL80),.BLN(BLN80),.WL(WL132));
sram_cell_6t_5 inst_cell_132_81 (.BL(BL81),.BLN(BLN81),.WL(WL132));
sram_cell_6t_5 inst_cell_132_82 (.BL(BL82),.BLN(BLN82),.WL(WL132));
sram_cell_6t_5 inst_cell_132_83 (.BL(BL83),.BLN(BLN83),.WL(WL132));
sram_cell_6t_5 inst_cell_132_84 (.BL(BL84),.BLN(BLN84),.WL(WL132));
sram_cell_6t_5 inst_cell_132_85 (.BL(BL85),.BLN(BLN85),.WL(WL132));
sram_cell_6t_5 inst_cell_132_86 (.BL(BL86),.BLN(BLN86),.WL(WL132));
sram_cell_6t_5 inst_cell_132_87 (.BL(BL87),.BLN(BLN87),.WL(WL132));
sram_cell_6t_5 inst_cell_132_88 (.BL(BL88),.BLN(BLN88),.WL(WL132));
sram_cell_6t_5 inst_cell_132_89 (.BL(BL89),.BLN(BLN89),.WL(WL132));
sram_cell_6t_5 inst_cell_132_90 (.BL(BL90),.BLN(BLN90),.WL(WL132));
sram_cell_6t_5 inst_cell_132_91 (.BL(BL91),.BLN(BLN91),.WL(WL132));
sram_cell_6t_5 inst_cell_132_92 (.BL(BL92),.BLN(BLN92),.WL(WL132));
sram_cell_6t_5 inst_cell_132_93 (.BL(BL93),.BLN(BLN93),.WL(WL132));
sram_cell_6t_5 inst_cell_132_94 (.BL(BL94),.BLN(BLN94),.WL(WL132));
sram_cell_6t_5 inst_cell_132_95 (.BL(BL95),.BLN(BLN95),.WL(WL132));
sram_cell_6t_5 inst_cell_132_96 (.BL(BL96),.BLN(BLN96),.WL(WL132));
sram_cell_6t_5 inst_cell_132_97 (.BL(BL97),.BLN(BLN97),.WL(WL132));
sram_cell_6t_5 inst_cell_132_98 (.BL(BL98),.BLN(BLN98),.WL(WL132));
sram_cell_6t_5 inst_cell_132_99 (.BL(BL99),.BLN(BLN99),.WL(WL132));
sram_cell_6t_5 inst_cell_132_100 (.BL(BL100),.BLN(BLN100),.WL(WL132));
sram_cell_6t_5 inst_cell_132_101 (.BL(BL101),.BLN(BLN101),.WL(WL132));
sram_cell_6t_5 inst_cell_132_102 (.BL(BL102),.BLN(BLN102),.WL(WL132));
sram_cell_6t_5 inst_cell_132_103 (.BL(BL103),.BLN(BLN103),.WL(WL132));
sram_cell_6t_5 inst_cell_132_104 (.BL(BL104),.BLN(BLN104),.WL(WL132));
sram_cell_6t_5 inst_cell_132_105 (.BL(BL105),.BLN(BLN105),.WL(WL132));
sram_cell_6t_5 inst_cell_132_106 (.BL(BL106),.BLN(BLN106),.WL(WL132));
sram_cell_6t_5 inst_cell_132_107 (.BL(BL107),.BLN(BLN107),.WL(WL132));
sram_cell_6t_5 inst_cell_132_108 (.BL(BL108),.BLN(BLN108),.WL(WL132));
sram_cell_6t_5 inst_cell_132_109 (.BL(BL109),.BLN(BLN109),.WL(WL132));
sram_cell_6t_5 inst_cell_132_110 (.BL(BL110),.BLN(BLN110),.WL(WL132));
sram_cell_6t_5 inst_cell_132_111 (.BL(BL111),.BLN(BLN111),.WL(WL132));
sram_cell_6t_5 inst_cell_132_112 (.BL(BL112),.BLN(BLN112),.WL(WL132));
sram_cell_6t_5 inst_cell_132_113 (.BL(BL113),.BLN(BLN113),.WL(WL132));
sram_cell_6t_5 inst_cell_132_114 (.BL(BL114),.BLN(BLN114),.WL(WL132));
sram_cell_6t_5 inst_cell_132_115 (.BL(BL115),.BLN(BLN115),.WL(WL132));
sram_cell_6t_5 inst_cell_132_116 (.BL(BL116),.BLN(BLN116),.WL(WL132));
sram_cell_6t_5 inst_cell_132_117 (.BL(BL117),.BLN(BLN117),.WL(WL132));
sram_cell_6t_5 inst_cell_132_118 (.BL(BL118),.BLN(BLN118),.WL(WL132));
sram_cell_6t_5 inst_cell_132_119 (.BL(BL119),.BLN(BLN119),.WL(WL132));
sram_cell_6t_5 inst_cell_132_120 (.BL(BL120),.BLN(BLN120),.WL(WL132));
sram_cell_6t_5 inst_cell_132_121 (.BL(BL121),.BLN(BLN121),.WL(WL132));
sram_cell_6t_5 inst_cell_132_122 (.BL(BL122),.BLN(BLN122),.WL(WL132));
sram_cell_6t_5 inst_cell_132_123 (.BL(BL123),.BLN(BLN123),.WL(WL132));
sram_cell_6t_5 inst_cell_132_124 (.BL(BL124),.BLN(BLN124),.WL(WL132));
sram_cell_6t_5 inst_cell_132_125 (.BL(BL125),.BLN(BLN125),.WL(WL132));
sram_cell_6t_5 inst_cell_132_126 (.BL(BL126),.BLN(BLN126),.WL(WL132));
sram_cell_6t_5 inst_cell_132_127 (.BL(BL127),.BLN(BLN127),.WL(WL132));
sram_cell_6t_5 inst_cell_133_0 (.BL(BL0),.BLN(BLN0),.WL(WL133));
sram_cell_6t_5 inst_cell_133_1 (.BL(BL1),.BLN(BLN1),.WL(WL133));
sram_cell_6t_5 inst_cell_133_2 (.BL(BL2),.BLN(BLN2),.WL(WL133));
sram_cell_6t_5 inst_cell_133_3 (.BL(BL3),.BLN(BLN3),.WL(WL133));
sram_cell_6t_5 inst_cell_133_4 (.BL(BL4),.BLN(BLN4),.WL(WL133));
sram_cell_6t_5 inst_cell_133_5 (.BL(BL5),.BLN(BLN5),.WL(WL133));
sram_cell_6t_5 inst_cell_133_6 (.BL(BL6),.BLN(BLN6),.WL(WL133));
sram_cell_6t_5 inst_cell_133_7 (.BL(BL7),.BLN(BLN7),.WL(WL133));
sram_cell_6t_5 inst_cell_133_8 (.BL(BL8),.BLN(BLN8),.WL(WL133));
sram_cell_6t_5 inst_cell_133_9 (.BL(BL9),.BLN(BLN9),.WL(WL133));
sram_cell_6t_5 inst_cell_133_10 (.BL(BL10),.BLN(BLN10),.WL(WL133));
sram_cell_6t_5 inst_cell_133_11 (.BL(BL11),.BLN(BLN11),.WL(WL133));
sram_cell_6t_5 inst_cell_133_12 (.BL(BL12),.BLN(BLN12),.WL(WL133));
sram_cell_6t_5 inst_cell_133_13 (.BL(BL13),.BLN(BLN13),.WL(WL133));
sram_cell_6t_5 inst_cell_133_14 (.BL(BL14),.BLN(BLN14),.WL(WL133));
sram_cell_6t_5 inst_cell_133_15 (.BL(BL15),.BLN(BLN15),.WL(WL133));
sram_cell_6t_5 inst_cell_133_16 (.BL(BL16),.BLN(BLN16),.WL(WL133));
sram_cell_6t_5 inst_cell_133_17 (.BL(BL17),.BLN(BLN17),.WL(WL133));
sram_cell_6t_5 inst_cell_133_18 (.BL(BL18),.BLN(BLN18),.WL(WL133));
sram_cell_6t_5 inst_cell_133_19 (.BL(BL19),.BLN(BLN19),.WL(WL133));
sram_cell_6t_5 inst_cell_133_20 (.BL(BL20),.BLN(BLN20),.WL(WL133));
sram_cell_6t_5 inst_cell_133_21 (.BL(BL21),.BLN(BLN21),.WL(WL133));
sram_cell_6t_5 inst_cell_133_22 (.BL(BL22),.BLN(BLN22),.WL(WL133));
sram_cell_6t_5 inst_cell_133_23 (.BL(BL23),.BLN(BLN23),.WL(WL133));
sram_cell_6t_5 inst_cell_133_24 (.BL(BL24),.BLN(BLN24),.WL(WL133));
sram_cell_6t_5 inst_cell_133_25 (.BL(BL25),.BLN(BLN25),.WL(WL133));
sram_cell_6t_5 inst_cell_133_26 (.BL(BL26),.BLN(BLN26),.WL(WL133));
sram_cell_6t_5 inst_cell_133_27 (.BL(BL27),.BLN(BLN27),.WL(WL133));
sram_cell_6t_5 inst_cell_133_28 (.BL(BL28),.BLN(BLN28),.WL(WL133));
sram_cell_6t_5 inst_cell_133_29 (.BL(BL29),.BLN(BLN29),.WL(WL133));
sram_cell_6t_5 inst_cell_133_30 (.BL(BL30),.BLN(BLN30),.WL(WL133));
sram_cell_6t_5 inst_cell_133_31 (.BL(BL31),.BLN(BLN31),.WL(WL133));
sram_cell_6t_5 inst_cell_133_32 (.BL(BL32),.BLN(BLN32),.WL(WL133));
sram_cell_6t_5 inst_cell_133_33 (.BL(BL33),.BLN(BLN33),.WL(WL133));
sram_cell_6t_5 inst_cell_133_34 (.BL(BL34),.BLN(BLN34),.WL(WL133));
sram_cell_6t_5 inst_cell_133_35 (.BL(BL35),.BLN(BLN35),.WL(WL133));
sram_cell_6t_5 inst_cell_133_36 (.BL(BL36),.BLN(BLN36),.WL(WL133));
sram_cell_6t_5 inst_cell_133_37 (.BL(BL37),.BLN(BLN37),.WL(WL133));
sram_cell_6t_5 inst_cell_133_38 (.BL(BL38),.BLN(BLN38),.WL(WL133));
sram_cell_6t_5 inst_cell_133_39 (.BL(BL39),.BLN(BLN39),.WL(WL133));
sram_cell_6t_5 inst_cell_133_40 (.BL(BL40),.BLN(BLN40),.WL(WL133));
sram_cell_6t_5 inst_cell_133_41 (.BL(BL41),.BLN(BLN41),.WL(WL133));
sram_cell_6t_5 inst_cell_133_42 (.BL(BL42),.BLN(BLN42),.WL(WL133));
sram_cell_6t_5 inst_cell_133_43 (.BL(BL43),.BLN(BLN43),.WL(WL133));
sram_cell_6t_5 inst_cell_133_44 (.BL(BL44),.BLN(BLN44),.WL(WL133));
sram_cell_6t_5 inst_cell_133_45 (.BL(BL45),.BLN(BLN45),.WL(WL133));
sram_cell_6t_5 inst_cell_133_46 (.BL(BL46),.BLN(BLN46),.WL(WL133));
sram_cell_6t_5 inst_cell_133_47 (.BL(BL47),.BLN(BLN47),.WL(WL133));
sram_cell_6t_5 inst_cell_133_48 (.BL(BL48),.BLN(BLN48),.WL(WL133));
sram_cell_6t_5 inst_cell_133_49 (.BL(BL49),.BLN(BLN49),.WL(WL133));
sram_cell_6t_5 inst_cell_133_50 (.BL(BL50),.BLN(BLN50),.WL(WL133));
sram_cell_6t_5 inst_cell_133_51 (.BL(BL51),.BLN(BLN51),.WL(WL133));
sram_cell_6t_5 inst_cell_133_52 (.BL(BL52),.BLN(BLN52),.WL(WL133));
sram_cell_6t_5 inst_cell_133_53 (.BL(BL53),.BLN(BLN53),.WL(WL133));
sram_cell_6t_5 inst_cell_133_54 (.BL(BL54),.BLN(BLN54),.WL(WL133));
sram_cell_6t_5 inst_cell_133_55 (.BL(BL55),.BLN(BLN55),.WL(WL133));
sram_cell_6t_5 inst_cell_133_56 (.BL(BL56),.BLN(BLN56),.WL(WL133));
sram_cell_6t_5 inst_cell_133_57 (.BL(BL57),.BLN(BLN57),.WL(WL133));
sram_cell_6t_5 inst_cell_133_58 (.BL(BL58),.BLN(BLN58),.WL(WL133));
sram_cell_6t_5 inst_cell_133_59 (.BL(BL59),.BLN(BLN59),.WL(WL133));
sram_cell_6t_5 inst_cell_133_60 (.BL(BL60),.BLN(BLN60),.WL(WL133));
sram_cell_6t_5 inst_cell_133_61 (.BL(BL61),.BLN(BLN61),.WL(WL133));
sram_cell_6t_5 inst_cell_133_62 (.BL(BL62),.BLN(BLN62),.WL(WL133));
sram_cell_6t_5 inst_cell_133_63 (.BL(BL63),.BLN(BLN63),.WL(WL133));
sram_cell_6t_5 inst_cell_133_64 (.BL(BL64),.BLN(BLN64),.WL(WL133));
sram_cell_6t_5 inst_cell_133_65 (.BL(BL65),.BLN(BLN65),.WL(WL133));
sram_cell_6t_5 inst_cell_133_66 (.BL(BL66),.BLN(BLN66),.WL(WL133));
sram_cell_6t_5 inst_cell_133_67 (.BL(BL67),.BLN(BLN67),.WL(WL133));
sram_cell_6t_5 inst_cell_133_68 (.BL(BL68),.BLN(BLN68),.WL(WL133));
sram_cell_6t_5 inst_cell_133_69 (.BL(BL69),.BLN(BLN69),.WL(WL133));
sram_cell_6t_5 inst_cell_133_70 (.BL(BL70),.BLN(BLN70),.WL(WL133));
sram_cell_6t_5 inst_cell_133_71 (.BL(BL71),.BLN(BLN71),.WL(WL133));
sram_cell_6t_5 inst_cell_133_72 (.BL(BL72),.BLN(BLN72),.WL(WL133));
sram_cell_6t_5 inst_cell_133_73 (.BL(BL73),.BLN(BLN73),.WL(WL133));
sram_cell_6t_5 inst_cell_133_74 (.BL(BL74),.BLN(BLN74),.WL(WL133));
sram_cell_6t_5 inst_cell_133_75 (.BL(BL75),.BLN(BLN75),.WL(WL133));
sram_cell_6t_5 inst_cell_133_76 (.BL(BL76),.BLN(BLN76),.WL(WL133));
sram_cell_6t_5 inst_cell_133_77 (.BL(BL77),.BLN(BLN77),.WL(WL133));
sram_cell_6t_5 inst_cell_133_78 (.BL(BL78),.BLN(BLN78),.WL(WL133));
sram_cell_6t_5 inst_cell_133_79 (.BL(BL79),.BLN(BLN79),.WL(WL133));
sram_cell_6t_5 inst_cell_133_80 (.BL(BL80),.BLN(BLN80),.WL(WL133));
sram_cell_6t_5 inst_cell_133_81 (.BL(BL81),.BLN(BLN81),.WL(WL133));
sram_cell_6t_5 inst_cell_133_82 (.BL(BL82),.BLN(BLN82),.WL(WL133));
sram_cell_6t_5 inst_cell_133_83 (.BL(BL83),.BLN(BLN83),.WL(WL133));
sram_cell_6t_5 inst_cell_133_84 (.BL(BL84),.BLN(BLN84),.WL(WL133));
sram_cell_6t_5 inst_cell_133_85 (.BL(BL85),.BLN(BLN85),.WL(WL133));
sram_cell_6t_5 inst_cell_133_86 (.BL(BL86),.BLN(BLN86),.WL(WL133));
sram_cell_6t_5 inst_cell_133_87 (.BL(BL87),.BLN(BLN87),.WL(WL133));
sram_cell_6t_5 inst_cell_133_88 (.BL(BL88),.BLN(BLN88),.WL(WL133));
sram_cell_6t_5 inst_cell_133_89 (.BL(BL89),.BLN(BLN89),.WL(WL133));
sram_cell_6t_5 inst_cell_133_90 (.BL(BL90),.BLN(BLN90),.WL(WL133));
sram_cell_6t_5 inst_cell_133_91 (.BL(BL91),.BLN(BLN91),.WL(WL133));
sram_cell_6t_5 inst_cell_133_92 (.BL(BL92),.BLN(BLN92),.WL(WL133));
sram_cell_6t_5 inst_cell_133_93 (.BL(BL93),.BLN(BLN93),.WL(WL133));
sram_cell_6t_5 inst_cell_133_94 (.BL(BL94),.BLN(BLN94),.WL(WL133));
sram_cell_6t_5 inst_cell_133_95 (.BL(BL95),.BLN(BLN95),.WL(WL133));
sram_cell_6t_5 inst_cell_133_96 (.BL(BL96),.BLN(BLN96),.WL(WL133));
sram_cell_6t_5 inst_cell_133_97 (.BL(BL97),.BLN(BLN97),.WL(WL133));
sram_cell_6t_5 inst_cell_133_98 (.BL(BL98),.BLN(BLN98),.WL(WL133));
sram_cell_6t_5 inst_cell_133_99 (.BL(BL99),.BLN(BLN99),.WL(WL133));
sram_cell_6t_5 inst_cell_133_100 (.BL(BL100),.BLN(BLN100),.WL(WL133));
sram_cell_6t_5 inst_cell_133_101 (.BL(BL101),.BLN(BLN101),.WL(WL133));
sram_cell_6t_5 inst_cell_133_102 (.BL(BL102),.BLN(BLN102),.WL(WL133));
sram_cell_6t_5 inst_cell_133_103 (.BL(BL103),.BLN(BLN103),.WL(WL133));
sram_cell_6t_5 inst_cell_133_104 (.BL(BL104),.BLN(BLN104),.WL(WL133));
sram_cell_6t_5 inst_cell_133_105 (.BL(BL105),.BLN(BLN105),.WL(WL133));
sram_cell_6t_5 inst_cell_133_106 (.BL(BL106),.BLN(BLN106),.WL(WL133));
sram_cell_6t_5 inst_cell_133_107 (.BL(BL107),.BLN(BLN107),.WL(WL133));
sram_cell_6t_5 inst_cell_133_108 (.BL(BL108),.BLN(BLN108),.WL(WL133));
sram_cell_6t_5 inst_cell_133_109 (.BL(BL109),.BLN(BLN109),.WL(WL133));
sram_cell_6t_5 inst_cell_133_110 (.BL(BL110),.BLN(BLN110),.WL(WL133));
sram_cell_6t_5 inst_cell_133_111 (.BL(BL111),.BLN(BLN111),.WL(WL133));
sram_cell_6t_5 inst_cell_133_112 (.BL(BL112),.BLN(BLN112),.WL(WL133));
sram_cell_6t_5 inst_cell_133_113 (.BL(BL113),.BLN(BLN113),.WL(WL133));
sram_cell_6t_5 inst_cell_133_114 (.BL(BL114),.BLN(BLN114),.WL(WL133));
sram_cell_6t_5 inst_cell_133_115 (.BL(BL115),.BLN(BLN115),.WL(WL133));
sram_cell_6t_5 inst_cell_133_116 (.BL(BL116),.BLN(BLN116),.WL(WL133));
sram_cell_6t_5 inst_cell_133_117 (.BL(BL117),.BLN(BLN117),.WL(WL133));
sram_cell_6t_5 inst_cell_133_118 (.BL(BL118),.BLN(BLN118),.WL(WL133));
sram_cell_6t_5 inst_cell_133_119 (.BL(BL119),.BLN(BLN119),.WL(WL133));
sram_cell_6t_5 inst_cell_133_120 (.BL(BL120),.BLN(BLN120),.WL(WL133));
sram_cell_6t_5 inst_cell_133_121 (.BL(BL121),.BLN(BLN121),.WL(WL133));
sram_cell_6t_5 inst_cell_133_122 (.BL(BL122),.BLN(BLN122),.WL(WL133));
sram_cell_6t_5 inst_cell_133_123 (.BL(BL123),.BLN(BLN123),.WL(WL133));
sram_cell_6t_5 inst_cell_133_124 (.BL(BL124),.BLN(BLN124),.WL(WL133));
sram_cell_6t_5 inst_cell_133_125 (.BL(BL125),.BLN(BLN125),.WL(WL133));
sram_cell_6t_5 inst_cell_133_126 (.BL(BL126),.BLN(BLN126),.WL(WL133));
sram_cell_6t_5 inst_cell_133_127 (.BL(BL127),.BLN(BLN127),.WL(WL133));
sram_cell_6t_5 inst_cell_134_0 (.BL(BL0),.BLN(BLN0),.WL(WL134));
sram_cell_6t_5 inst_cell_134_1 (.BL(BL1),.BLN(BLN1),.WL(WL134));
sram_cell_6t_5 inst_cell_134_2 (.BL(BL2),.BLN(BLN2),.WL(WL134));
sram_cell_6t_5 inst_cell_134_3 (.BL(BL3),.BLN(BLN3),.WL(WL134));
sram_cell_6t_5 inst_cell_134_4 (.BL(BL4),.BLN(BLN4),.WL(WL134));
sram_cell_6t_5 inst_cell_134_5 (.BL(BL5),.BLN(BLN5),.WL(WL134));
sram_cell_6t_5 inst_cell_134_6 (.BL(BL6),.BLN(BLN6),.WL(WL134));
sram_cell_6t_5 inst_cell_134_7 (.BL(BL7),.BLN(BLN7),.WL(WL134));
sram_cell_6t_5 inst_cell_134_8 (.BL(BL8),.BLN(BLN8),.WL(WL134));
sram_cell_6t_5 inst_cell_134_9 (.BL(BL9),.BLN(BLN9),.WL(WL134));
sram_cell_6t_5 inst_cell_134_10 (.BL(BL10),.BLN(BLN10),.WL(WL134));
sram_cell_6t_5 inst_cell_134_11 (.BL(BL11),.BLN(BLN11),.WL(WL134));
sram_cell_6t_5 inst_cell_134_12 (.BL(BL12),.BLN(BLN12),.WL(WL134));
sram_cell_6t_5 inst_cell_134_13 (.BL(BL13),.BLN(BLN13),.WL(WL134));
sram_cell_6t_5 inst_cell_134_14 (.BL(BL14),.BLN(BLN14),.WL(WL134));
sram_cell_6t_5 inst_cell_134_15 (.BL(BL15),.BLN(BLN15),.WL(WL134));
sram_cell_6t_5 inst_cell_134_16 (.BL(BL16),.BLN(BLN16),.WL(WL134));
sram_cell_6t_5 inst_cell_134_17 (.BL(BL17),.BLN(BLN17),.WL(WL134));
sram_cell_6t_5 inst_cell_134_18 (.BL(BL18),.BLN(BLN18),.WL(WL134));
sram_cell_6t_5 inst_cell_134_19 (.BL(BL19),.BLN(BLN19),.WL(WL134));
sram_cell_6t_5 inst_cell_134_20 (.BL(BL20),.BLN(BLN20),.WL(WL134));
sram_cell_6t_5 inst_cell_134_21 (.BL(BL21),.BLN(BLN21),.WL(WL134));
sram_cell_6t_5 inst_cell_134_22 (.BL(BL22),.BLN(BLN22),.WL(WL134));
sram_cell_6t_5 inst_cell_134_23 (.BL(BL23),.BLN(BLN23),.WL(WL134));
sram_cell_6t_5 inst_cell_134_24 (.BL(BL24),.BLN(BLN24),.WL(WL134));
sram_cell_6t_5 inst_cell_134_25 (.BL(BL25),.BLN(BLN25),.WL(WL134));
sram_cell_6t_5 inst_cell_134_26 (.BL(BL26),.BLN(BLN26),.WL(WL134));
sram_cell_6t_5 inst_cell_134_27 (.BL(BL27),.BLN(BLN27),.WL(WL134));
sram_cell_6t_5 inst_cell_134_28 (.BL(BL28),.BLN(BLN28),.WL(WL134));
sram_cell_6t_5 inst_cell_134_29 (.BL(BL29),.BLN(BLN29),.WL(WL134));
sram_cell_6t_5 inst_cell_134_30 (.BL(BL30),.BLN(BLN30),.WL(WL134));
sram_cell_6t_5 inst_cell_134_31 (.BL(BL31),.BLN(BLN31),.WL(WL134));
sram_cell_6t_5 inst_cell_134_32 (.BL(BL32),.BLN(BLN32),.WL(WL134));
sram_cell_6t_5 inst_cell_134_33 (.BL(BL33),.BLN(BLN33),.WL(WL134));
sram_cell_6t_5 inst_cell_134_34 (.BL(BL34),.BLN(BLN34),.WL(WL134));
sram_cell_6t_5 inst_cell_134_35 (.BL(BL35),.BLN(BLN35),.WL(WL134));
sram_cell_6t_5 inst_cell_134_36 (.BL(BL36),.BLN(BLN36),.WL(WL134));
sram_cell_6t_5 inst_cell_134_37 (.BL(BL37),.BLN(BLN37),.WL(WL134));
sram_cell_6t_5 inst_cell_134_38 (.BL(BL38),.BLN(BLN38),.WL(WL134));
sram_cell_6t_5 inst_cell_134_39 (.BL(BL39),.BLN(BLN39),.WL(WL134));
sram_cell_6t_5 inst_cell_134_40 (.BL(BL40),.BLN(BLN40),.WL(WL134));
sram_cell_6t_5 inst_cell_134_41 (.BL(BL41),.BLN(BLN41),.WL(WL134));
sram_cell_6t_5 inst_cell_134_42 (.BL(BL42),.BLN(BLN42),.WL(WL134));
sram_cell_6t_5 inst_cell_134_43 (.BL(BL43),.BLN(BLN43),.WL(WL134));
sram_cell_6t_5 inst_cell_134_44 (.BL(BL44),.BLN(BLN44),.WL(WL134));
sram_cell_6t_5 inst_cell_134_45 (.BL(BL45),.BLN(BLN45),.WL(WL134));
sram_cell_6t_5 inst_cell_134_46 (.BL(BL46),.BLN(BLN46),.WL(WL134));
sram_cell_6t_5 inst_cell_134_47 (.BL(BL47),.BLN(BLN47),.WL(WL134));
sram_cell_6t_5 inst_cell_134_48 (.BL(BL48),.BLN(BLN48),.WL(WL134));
sram_cell_6t_5 inst_cell_134_49 (.BL(BL49),.BLN(BLN49),.WL(WL134));
sram_cell_6t_5 inst_cell_134_50 (.BL(BL50),.BLN(BLN50),.WL(WL134));
sram_cell_6t_5 inst_cell_134_51 (.BL(BL51),.BLN(BLN51),.WL(WL134));
sram_cell_6t_5 inst_cell_134_52 (.BL(BL52),.BLN(BLN52),.WL(WL134));
sram_cell_6t_5 inst_cell_134_53 (.BL(BL53),.BLN(BLN53),.WL(WL134));
sram_cell_6t_5 inst_cell_134_54 (.BL(BL54),.BLN(BLN54),.WL(WL134));
sram_cell_6t_5 inst_cell_134_55 (.BL(BL55),.BLN(BLN55),.WL(WL134));
sram_cell_6t_5 inst_cell_134_56 (.BL(BL56),.BLN(BLN56),.WL(WL134));
sram_cell_6t_5 inst_cell_134_57 (.BL(BL57),.BLN(BLN57),.WL(WL134));
sram_cell_6t_5 inst_cell_134_58 (.BL(BL58),.BLN(BLN58),.WL(WL134));
sram_cell_6t_5 inst_cell_134_59 (.BL(BL59),.BLN(BLN59),.WL(WL134));
sram_cell_6t_5 inst_cell_134_60 (.BL(BL60),.BLN(BLN60),.WL(WL134));
sram_cell_6t_5 inst_cell_134_61 (.BL(BL61),.BLN(BLN61),.WL(WL134));
sram_cell_6t_5 inst_cell_134_62 (.BL(BL62),.BLN(BLN62),.WL(WL134));
sram_cell_6t_5 inst_cell_134_63 (.BL(BL63),.BLN(BLN63),.WL(WL134));
sram_cell_6t_5 inst_cell_134_64 (.BL(BL64),.BLN(BLN64),.WL(WL134));
sram_cell_6t_5 inst_cell_134_65 (.BL(BL65),.BLN(BLN65),.WL(WL134));
sram_cell_6t_5 inst_cell_134_66 (.BL(BL66),.BLN(BLN66),.WL(WL134));
sram_cell_6t_5 inst_cell_134_67 (.BL(BL67),.BLN(BLN67),.WL(WL134));
sram_cell_6t_5 inst_cell_134_68 (.BL(BL68),.BLN(BLN68),.WL(WL134));
sram_cell_6t_5 inst_cell_134_69 (.BL(BL69),.BLN(BLN69),.WL(WL134));
sram_cell_6t_5 inst_cell_134_70 (.BL(BL70),.BLN(BLN70),.WL(WL134));
sram_cell_6t_5 inst_cell_134_71 (.BL(BL71),.BLN(BLN71),.WL(WL134));
sram_cell_6t_5 inst_cell_134_72 (.BL(BL72),.BLN(BLN72),.WL(WL134));
sram_cell_6t_5 inst_cell_134_73 (.BL(BL73),.BLN(BLN73),.WL(WL134));
sram_cell_6t_5 inst_cell_134_74 (.BL(BL74),.BLN(BLN74),.WL(WL134));
sram_cell_6t_5 inst_cell_134_75 (.BL(BL75),.BLN(BLN75),.WL(WL134));
sram_cell_6t_5 inst_cell_134_76 (.BL(BL76),.BLN(BLN76),.WL(WL134));
sram_cell_6t_5 inst_cell_134_77 (.BL(BL77),.BLN(BLN77),.WL(WL134));
sram_cell_6t_5 inst_cell_134_78 (.BL(BL78),.BLN(BLN78),.WL(WL134));
sram_cell_6t_5 inst_cell_134_79 (.BL(BL79),.BLN(BLN79),.WL(WL134));
sram_cell_6t_5 inst_cell_134_80 (.BL(BL80),.BLN(BLN80),.WL(WL134));
sram_cell_6t_5 inst_cell_134_81 (.BL(BL81),.BLN(BLN81),.WL(WL134));
sram_cell_6t_5 inst_cell_134_82 (.BL(BL82),.BLN(BLN82),.WL(WL134));
sram_cell_6t_5 inst_cell_134_83 (.BL(BL83),.BLN(BLN83),.WL(WL134));
sram_cell_6t_5 inst_cell_134_84 (.BL(BL84),.BLN(BLN84),.WL(WL134));
sram_cell_6t_5 inst_cell_134_85 (.BL(BL85),.BLN(BLN85),.WL(WL134));
sram_cell_6t_5 inst_cell_134_86 (.BL(BL86),.BLN(BLN86),.WL(WL134));
sram_cell_6t_5 inst_cell_134_87 (.BL(BL87),.BLN(BLN87),.WL(WL134));
sram_cell_6t_5 inst_cell_134_88 (.BL(BL88),.BLN(BLN88),.WL(WL134));
sram_cell_6t_5 inst_cell_134_89 (.BL(BL89),.BLN(BLN89),.WL(WL134));
sram_cell_6t_5 inst_cell_134_90 (.BL(BL90),.BLN(BLN90),.WL(WL134));
sram_cell_6t_5 inst_cell_134_91 (.BL(BL91),.BLN(BLN91),.WL(WL134));
sram_cell_6t_5 inst_cell_134_92 (.BL(BL92),.BLN(BLN92),.WL(WL134));
sram_cell_6t_5 inst_cell_134_93 (.BL(BL93),.BLN(BLN93),.WL(WL134));
sram_cell_6t_5 inst_cell_134_94 (.BL(BL94),.BLN(BLN94),.WL(WL134));
sram_cell_6t_5 inst_cell_134_95 (.BL(BL95),.BLN(BLN95),.WL(WL134));
sram_cell_6t_5 inst_cell_134_96 (.BL(BL96),.BLN(BLN96),.WL(WL134));
sram_cell_6t_5 inst_cell_134_97 (.BL(BL97),.BLN(BLN97),.WL(WL134));
sram_cell_6t_5 inst_cell_134_98 (.BL(BL98),.BLN(BLN98),.WL(WL134));
sram_cell_6t_5 inst_cell_134_99 (.BL(BL99),.BLN(BLN99),.WL(WL134));
sram_cell_6t_5 inst_cell_134_100 (.BL(BL100),.BLN(BLN100),.WL(WL134));
sram_cell_6t_5 inst_cell_134_101 (.BL(BL101),.BLN(BLN101),.WL(WL134));
sram_cell_6t_5 inst_cell_134_102 (.BL(BL102),.BLN(BLN102),.WL(WL134));
sram_cell_6t_5 inst_cell_134_103 (.BL(BL103),.BLN(BLN103),.WL(WL134));
sram_cell_6t_5 inst_cell_134_104 (.BL(BL104),.BLN(BLN104),.WL(WL134));
sram_cell_6t_5 inst_cell_134_105 (.BL(BL105),.BLN(BLN105),.WL(WL134));
sram_cell_6t_5 inst_cell_134_106 (.BL(BL106),.BLN(BLN106),.WL(WL134));
sram_cell_6t_5 inst_cell_134_107 (.BL(BL107),.BLN(BLN107),.WL(WL134));
sram_cell_6t_5 inst_cell_134_108 (.BL(BL108),.BLN(BLN108),.WL(WL134));
sram_cell_6t_5 inst_cell_134_109 (.BL(BL109),.BLN(BLN109),.WL(WL134));
sram_cell_6t_5 inst_cell_134_110 (.BL(BL110),.BLN(BLN110),.WL(WL134));
sram_cell_6t_5 inst_cell_134_111 (.BL(BL111),.BLN(BLN111),.WL(WL134));
sram_cell_6t_5 inst_cell_134_112 (.BL(BL112),.BLN(BLN112),.WL(WL134));
sram_cell_6t_5 inst_cell_134_113 (.BL(BL113),.BLN(BLN113),.WL(WL134));
sram_cell_6t_5 inst_cell_134_114 (.BL(BL114),.BLN(BLN114),.WL(WL134));
sram_cell_6t_5 inst_cell_134_115 (.BL(BL115),.BLN(BLN115),.WL(WL134));
sram_cell_6t_5 inst_cell_134_116 (.BL(BL116),.BLN(BLN116),.WL(WL134));
sram_cell_6t_5 inst_cell_134_117 (.BL(BL117),.BLN(BLN117),.WL(WL134));
sram_cell_6t_5 inst_cell_134_118 (.BL(BL118),.BLN(BLN118),.WL(WL134));
sram_cell_6t_5 inst_cell_134_119 (.BL(BL119),.BLN(BLN119),.WL(WL134));
sram_cell_6t_5 inst_cell_134_120 (.BL(BL120),.BLN(BLN120),.WL(WL134));
sram_cell_6t_5 inst_cell_134_121 (.BL(BL121),.BLN(BLN121),.WL(WL134));
sram_cell_6t_5 inst_cell_134_122 (.BL(BL122),.BLN(BLN122),.WL(WL134));
sram_cell_6t_5 inst_cell_134_123 (.BL(BL123),.BLN(BLN123),.WL(WL134));
sram_cell_6t_5 inst_cell_134_124 (.BL(BL124),.BLN(BLN124),.WL(WL134));
sram_cell_6t_5 inst_cell_134_125 (.BL(BL125),.BLN(BLN125),.WL(WL134));
sram_cell_6t_5 inst_cell_134_126 (.BL(BL126),.BLN(BLN126),.WL(WL134));
sram_cell_6t_5 inst_cell_134_127 (.BL(BL127),.BLN(BLN127),.WL(WL134));
sram_cell_6t_5 inst_cell_135_0 (.BL(BL0),.BLN(BLN0),.WL(WL135));
sram_cell_6t_5 inst_cell_135_1 (.BL(BL1),.BLN(BLN1),.WL(WL135));
sram_cell_6t_5 inst_cell_135_2 (.BL(BL2),.BLN(BLN2),.WL(WL135));
sram_cell_6t_5 inst_cell_135_3 (.BL(BL3),.BLN(BLN3),.WL(WL135));
sram_cell_6t_5 inst_cell_135_4 (.BL(BL4),.BLN(BLN4),.WL(WL135));
sram_cell_6t_5 inst_cell_135_5 (.BL(BL5),.BLN(BLN5),.WL(WL135));
sram_cell_6t_5 inst_cell_135_6 (.BL(BL6),.BLN(BLN6),.WL(WL135));
sram_cell_6t_5 inst_cell_135_7 (.BL(BL7),.BLN(BLN7),.WL(WL135));
sram_cell_6t_5 inst_cell_135_8 (.BL(BL8),.BLN(BLN8),.WL(WL135));
sram_cell_6t_5 inst_cell_135_9 (.BL(BL9),.BLN(BLN9),.WL(WL135));
sram_cell_6t_5 inst_cell_135_10 (.BL(BL10),.BLN(BLN10),.WL(WL135));
sram_cell_6t_5 inst_cell_135_11 (.BL(BL11),.BLN(BLN11),.WL(WL135));
sram_cell_6t_5 inst_cell_135_12 (.BL(BL12),.BLN(BLN12),.WL(WL135));
sram_cell_6t_5 inst_cell_135_13 (.BL(BL13),.BLN(BLN13),.WL(WL135));
sram_cell_6t_5 inst_cell_135_14 (.BL(BL14),.BLN(BLN14),.WL(WL135));
sram_cell_6t_5 inst_cell_135_15 (.BL(BL15),.BLN(BLN15),.WL(WL135));
sram_cell_6t_5 inst_cell_135_16 (.BL(BL16),.BLN(BLN16),.WL(WL135));
sram_cell_6t_5 inst_cell_135_17 (.BL(BL17),.BLN(BLN17),.WL(WL135));
sram_cell_6t_5 inst_cell_135_18 (.BL(BL18),.BLN(BLN18),.WL(WL135));
sram_cell_6t_5 inst_cell_135_19 (.BL(BL19),.BLN(BLN19),.WL(WL135));
sram_cell_6t_5 inst_cell_135_20 (.BL(BL20),.BLN(BLN20),.WL(WL135));
sram_cell_6t_5 inst_cell_135_21 (.BL(BL21),.BLN(BLN21),.WL(WL135));
sram_cell_6t_5 inst_cell_135_22 (.BL(BL22),.BLN(BLN22),.WL(WL135));
sram_cell_6t_5 inst_cell_135_23 (.BL(BL23),.BLN(BLN23),.WL(WL135));
sram_cell_6t_5 inst_cell_135_24 (.BL(BL24),.BLN(BLN24),.WL(WL135));
sram_cell_6t_5 inst_cell_135_25 (.BL(BL25),.BLN(BLN25),.WL(WL135));
sram_cell_6t_5 inst_cell_135_26 (.BL(BL26),.BLN(BLN26),.WL(WL135));
sram_cell_6t_5 inst_cell_135_27 (.BL(BL27),.BLN(BLN27),.WL(WL135));
sram_cell_6t_5 inst_cell_135_28 (.BL(BL28),.BLN(BLN28),.WL(WL135));
sram_cell_6t_5 inst_cell_135_29 (.BL(BL29),.BLN(BLN29),.WL(WL135));
sram_cell_6t_5 inst_cell_135_30 (.BL(BL30),.BLN(BLN30),.WL(WL135));
sram_cell_6t_5 inst_cell_135_31 (.BL(BL31),.BLN(BLN31),.WL(WL135));
sram_cell_6t_5 inst_cell_135_32 (.BL(BL32),.BLN(BLN32),.WL(WL135));
sram_cell_6t_5 inst_cell_135_33 (.BL(BL33),.BLN(BLN33),.WL(WL135));
sram_cell_6t_5 inst_cell_135_34 (.BL(BL34),.BLN(BLN34),.WL(WL135));
sram_cell_6t_5 inst_cell_135_35 (.BL(BL35),.BLN(BLN35),.WL(WL135));
sram_cell_6t_5 inst_cell_135_36 (.BL(BL36),.BLN(BLN36),.WL(WL135));
sram_cell_6t_5 inst_cell_135_37 (.BL(BL37),.BLN(BLN37),.WL(WL135));
sram_cell_6t_5 inst_cell_135_38 (.BL(BL38),.BLN(BLN38),.WL(WL135));
sram_cell_6t_5 inst_cell_135_39 (.BL(BL39),.BLN(BLN39),.WL(WL135));
sram_cell_6t_5 inst_cell_135_40 (.BL(BL40),.BLN(BLN40),.WL(WL135));
sram_cell_6t_5 inst_cell_135_41 (.BL(BL41),.BLN(BLN41),.WL(WL135));
sram_cell_6t_5 inst_cell_135_42 (.BL(BL42),.BLN(BLN42),.WL(WL135));
sram_cell_6t_5 inst_cell_135_43 (.BL(BL43),.BLN(BLN43),.WL(WL135));
sram_cell_6t_5 inst_cell_135_44 (.BL(BL44),.BLN(BLN44),.WL(WL135));
sram_cell_6t_5 inst_cell_135_45 (.BL(BL45),.BLN(BLN45),.WL(WL135));
sram_cell_6t_5 inst_cell_135_46 (.BL(BL46),.BLN(BLN46),.WL(WL135));
sram_cell_6t_5 inst_cell_135_47 (.BL(BL47),.BLN(BLN47),.WL(WL135));
sram_cell_6t_5 inst_cell_135_48 (.BL(BL48),.BLN(BLN48),.WL(WL135));
sram_cell_6t_5 inst_cell_135_49 (.BL(BL49),.BLN(BLN49),.WL(WL135));
sram_cell_6t_5 inst_cell_135_50 (.BL(BL50),.BLN(BLN50),.WL(WL135));
sram_cell_6t_5 inst_cell_135_51 (.BL(BL51),.BLN(BLN51),.WL(WL135));
sram_cell_6t_5 inst_cell_135_52 (.BL(BL52),.BLN(BLN52),.WL(WL135));
sram_cell_6t_5 inst_cell_135_53 (.BL(BL53),.BLN(BLN53),.WL(WL135));
sram_cell_6t_5 inst_cell_135_54 (.BL(BL54),.BLN(BLN54),.WL(WL135));
sram_cell_6t_5 inst_cell_135_55 (.BL(BL55),.BLN(BLN55),.WL(WL135));
sram_cell_6t_5 inst_cell_135_56 (.BL(BL56),.BLN(BLN56),.WL(WL135));
sram_cell_6t_5 inst_cell_135_57 (.BL(BL57),.BLN(BLN57),.WL(WL135));
sram_cell_6t_5 inst_cell_135_58 (.BL(BL58),.BLN(BLN58),.WL(WL135));
sram_cell_6t_5 inst_cell_135_59 (.BL(BL59),.BLN(BLN59),.WL(WL135));
sram_cell_6t_5 inst_cell_135_60 (.BL(BL60),.BLN(BLN60),.WL(WL135));
sram_cell_6t_5 inst_cell_135_61 (.BL(BL61),.BLN(BLN61),.WL(WL135));
sram_cell_6t_5 inst_cell_135_62 (.BL(BL62),.BLN(BLN62),.WL(WL135));
sram_cell_6t_5 inst_cell_135_63 (.BL(BL63),.BLN(BLN63),.WL(WL135));
sram_cell_6t_5 inst_cell_135_64 (.BL(BL64),.BLN(BLN64),.WL(WL135));
sram_cell_6t_5 inst_cell_135_65 (.BL(BL65),.BLN(BLN65),.WL(WL135));
sram_cell_6t_5 inst_cell_135_66 (.BL(BL66),.BLN(BLN66),.WL(WL135));
sram_cell_6t_5 inst_cell_135_67 (.BL(BL67),.BLN(BLN67),.WL(WL135));
sram_cell_6t_5 inst_cell_135_68 (.BL(BL68),.BLN(BLN68),.WL(WL135));
sram_cell_6t_5 inst_cell_135_69 (.BL(BL69),.BLN(BLN69),.WL(WL135));
sram_cell_6t_5 inst_cell_135_70 (.BL(BL70),.BLN(BLN70),.WL(WL135));
sram_cell_6t_5 inst_cell_135_71 (.BL(BL71),.BLN(BLN71),.WL(WL135));
sram_cell_6t_5 inst_cell_135_72 (.BL(BL72),.BLN(BLN72),.WL(WL135));
sram_cell_6t_5 inst_cell_135_73 (.BL(BL73),.BLN(BLN73),.WL(WL135));
sram_cell_6t_5 inst_cell_135_74 (.BL(BL74),.BLN(BLN74),.WL(WL135));
sram_cell_6t_5 inst_cell_135_75 (.BL(BL75),.BLN(BLN75),.WL(WL135));
sram_cell_6t_5 inst_cell_135_76 (.BL(BL76),.BLN(BLN76),.WL(WL135));
sram_cell_6t_5 inst_cell_135_77 (.BL(BL77),.BLN(BLN77),.WL(WL135));
sram_cell_6t_5 inst_cell_135_78 (.BL(BL78),.BLN(BLN78),.WL(WL135));
sram_cell_6t_5 inst_cell_135_79 (.BL(BL79),.BLN(BLN79),.WL(WL135));
sram_cell_6t_5 inst_cell_135_80 (.BL(BL80),.BLN(BLN80),.WL(WL135));
sram_cell_6t_5 inst_cell_135_81 (.BL(BL81),.BLN(BLN81),.WL(WL135));
sram_cell_6t_5 inst_cell_135_82 (.BL(BL82),.BLN(BLN82),.WL(WL135));
sram_cell_6t_5 inst_cell_135_83 (.BL(BL83),.BLN(BLN83),.WL(WL135));
sram_cell_6t_5 inst_cell_135_84 (.BL(BL84),.BLN(BLN84),.WL(WL135));
sram_cell_6t_5 inst_cell_135_85 (.BL(BL85),.BLN(BLN85),.WL(WL135));
sram_cell_6t_5 inst_cell_135_86 (.BL(BL86),.BLN(BLN86),.WL(WL135));
sram_cell_6t_5 inst_cell_135_87 (.BL(BL87),.BLN(BLN87),.WL(WL135));
sram_cell_6t_5 inst_cell_135_88 (.BL(BL88),.BLN(BLN88),.WL(WL135));
sram_cell_6t_5 inst_cell_135_89 (.BL(BL89),.BLN(BLN89),.WL(WL135));
sram_cell_6t_5 inst_cell_135_90 (.BL(BL90),.BLN(BLN90),.WL(WL135));
sram_cell_6t_5 inst_cell_135_91 (.BL(BL91),.BLN(BLN91),.WL(WL135));
sram_cell_6t_5 inst_cell_135_92 (.BL(BL92),.BLN(BLN92),.WL(WL135));
sram_cell_6t_5 inst_cell_135_93 (.BL(BL93),.BLN(BLN93),.WL(WL135));
sram_cell_6t_5 inst_cell_135_94 (.BL(BL94),.BLN(BLN94),.WL(WL135));
sram_cell_6t_5 inst_cell_135_95 (.BL(BL95),.BLN(BLN95),.WL(WL135));
sram_cell_6t_5 inst_cell_135_96 (.BL(BL96),.BLN(BLN96),.WL(WL135));
sram_cell_6t_5 inst_cell_135_97 (.BL(BL97),.BLN(BLN97),.WL(WL135));
sram_cell_6t_5 inst_cell_135_98 (.BL(BL98),.BLN(BLN98),.WL(WL135));
sram_cell_6t_5 inst_cell_135_99 (.BL(BL99),.BLN(BLN99),.WL(WL135));
sram_cell_6t_5 inst_cell_135_100 (.BL(BL100),.BLN(BLN100),.WL(WL135));
sram_cell_6t_5 inst_cell_135_101 (.BL(BL101),.BLN(BLN101),.WL(WL135));
sram_cell_6t_5 inst_cell_135_102 (.BL(BL102),.BLN(BLN102),.WL(WL135));
sram_cell_6t_5 inst_cell_135_103 (.BL(BL103),.BLN(BLN103),.WL(WL135));
sram_cell_6t_5 inst_cell_135_104 (.BL(BL104),.BLN(BLN104),.WL(WL135));
sram_cell_6t_5 inst_cell_135_105 (.BL(BL105),.BLN(BLN105),.WL(WL135));
sram_cell_6t_5 inst_cell_135_106 (.BL(BL106),.BLN(BLN106),.WL(WL135));
sram_cell_6t_5 inst_cell_135_107 (.BL(BL107),.BLN(BLN107),.WL(WL135));
sram_cell_6t_5 inst_cell_135_108 (.BL(BL108),.BLN(BLN108),.WL(WL135));
sram_cell_6t_5 inst_cell_135_109 (.BL(BL109),.BLN(BLN109),.WL(WL135));
sram_cell_6t_5 inst_cell_135_110 (.BL(BL110),.BLN(BLN110),.WL(WL135));
sram_cell_6t_5 inst_cell_135_111 (.BL(BL111),.BLN(BLN111),.WL(WL135));
sram_cell_6t_5 inst_cell_135_112 (.BL(BL112),.BLN(BLN112),.WL(WL135));
sram_cell_6t_5 inst_cell_135_113 (.BL(BL113),.BLN(BLN113),.WL(WL135));
sram_cell_6t_5 inst_cell_135_114 (.BL(BL114),.BLN(BLN114),.WL(WL135));
sram_cell_6t_5 inst_cell_135_115 (.BL(BL115),.BLN(BLN115),.WL(WL135));
sram_cell_6t_5 inst_cell_135_116 (.BL(BL116),.BLN(BLN116),.WL(WL135));
sram_cell_6t_5 inst_cell_135_117 (.BL(BL117),.BLN(BLN117),.WL(WL135));
sram_cell_6t_5 inst_cell_135_118 (.BL(BL118),.BLN(BLN118),.WL(WL135));
sram_cell_6t_5 inst_cell_135_119 (.BL(BL119),.BLN(BLN119),.WL(WL135));
sram_cell_6t_5 inst_cell_135_120 (.BL(BL120),.BLN(BLN120),.WL(WL135));
sram_cell_6t_5 inst_cell_135_121 (.BL(BL121),.BLN(BLN121),.WL(WL135));
sram_cell_6t_5 inst_cell_135_122 (.BL(BL122),.BLN(BLN122),.WL(WL135));
sram_cell_6t_5 inst_cell_135_123 (.BL(BL123),.BLN(BLN123),.WL(WL135));
sram_cell_6t_5 inst_cell_135_124 (.BL(BL124),.BLN(BLN124),.WL(WL135));
sram_cell_6t_5 inst_cell_135_125 (.BL(BL125),.BLN(BLN125),.WL(WL135));
sram_cell_6t_5 inst_cell_135_126 (.BL(BL126),.BLN(BLN126),.WL(WL135));
sram_cell_6t_5 inst_cell_135_127 (.BL(BL127),.BLN(BLN127),.WL(WL135));
sram_cell_6t_5 inst_cell_136_0 (.BL(BL0),.BLN(BLN0),.WL(WL136));
sram_cell_6t_5 inst_cell_136_1 (.BL(BL1),.BLN(BLN1),.WL(WL136));
sram_cell_6t_5 inst_cell_136_2 (.BL(BL2),.BLN(BLN2),.WL(WL136));
sram_cell_6t_5 inst_cell_136_3 (.BL(BL3),.BLN(BLN3),.WL(WL136));
sram_cell_6t_5 inst_cell_136_4 (.BL(BL4),.BLN(BLN4),.WL(WL136));
sram_cell_6t_5 inst_cell_136_5 (.BL(BL5),.BLN(BLN5),.WL(WL136));
sram_cell_6t_5 inst_cell_136_6 (.BL(BL6),.BLN(BLN6),.WL(WL136));
sram_cell_6t_5 inst_cell_136_7 (.BL(BL7),.BLN(BLN7),.WL(WL136));
sram_cell_6t_5 inst_cell_136_8 (.BL(BL8),.BLN(BLN8),.WL(WL136));
sram_cell_6t_5 inst_cell_136_9 (.BL(BL9),.BLN(BLN9),.WL(WL136));
sram_cell_6t_5 inst_cell_136_10 (.BL(BL10),.BLN(BLN10),.WL(WL136));
sram_cell_6t_5 inst_cell_136_11 (.BL(BL11),.BLN(BLN11),.WL(WL136));
sram_cell_6t_5 inst_cell_136_12 (.BL(BL12),.BLN(BLN12),.WL(WL136));
sram_cell_6t_5 inst_cell_136_13 (.BL(BL13),.BLN(BLN13),.WL(WL136));
sram_cell_6t_5 inst_cell_136_14 (.BL(BL14),.BLN(BLN14),.WL(WL136));
sram_cell_6t_5 inst_cell_136_15 (.BL(BL15),.BLN(BLN15),.WL(WL136));
sram_cell_6t_5 inst_cell_136_16 (.BL(BL16),.BLN(BLN16),.WL(WL136));
sram_cell_6t_5 inst_cell_136_17 (.BL(BL17),.BLN(BLN17),.WL(WL136));
sram_cell_6t_5 inst_cell_136_18 (.BL(BL18),.BLN(BLN18),.WL(WL136));
sram_cell_6t_5 inst_cell_136_19 (.BL(BL19),.BLN(BLN19),.WL(WL136));
sram_cell_6t_5 inst_cell_136_20 (.BL(BL20),.BLN(BLN20),.WL(WL136));
sram_cell_6t_5 inst_cell_136_21 (.BL(BL21),.BLN(BLN21),.WL(WL136));
sram_cell_6t_5 inst_cell_136_22 (.BL(BL22),.BLN(BLN22),.WL(WL136));
sram_cell_6t_5 inst_cell_136_23 (.BL(BL23),.BLN(BLN23),.WL(WL136));
sram_cell_6t_5 inst_cell_136_24 (.BL(BL24),.BLN(BLN24),.WL(WL136));
sram_cell_6t_5 inst_cell_136_25 (.BL(BL25),.BLN(BLN25),.WL(WL136));
sram_cell_6t_5 inst_cell_136_26 (.BL(BL26),.BLN(BLN26),.WL(WL136));
sram_cell_6t_5 inst_cell_136_27 (.BL(BL27),.BLN(BLN27),.WL(WL136));
sram_cell_6t_5 inst_cell_136_28 (.BL(BL28),.BLN(BLN28),.WL(WL136));
sram_cell_6t_5 inst_cell_136_29 (.BL(BL29),.BLN(BLN29),.WL(WL136));
sram_cell_6t_5 inst_cell_136_30 (.BL(BL30),.BLN(BLN30),.WL(WL136));
sram_cell_6t_5 inst_cell_136_31 (.BL(BL31),.BLN(BLN31),.WL(WL136));
sram_cell_6t_5 inst_cell_136_32 (.BL(BL32),.BLN(BLN32),.WL(WL136));
sram_cell_6t_5 inst_cell_136_33 (.BL(BL33),.BLN(BLN33),.WL(WL136));
sram_cell_6t_5 inst_cell_136_34 (.BL(BL34),.BLN(BLN34),.WL(WL136));
sram_cell_6t_5 inst_cell_136_35 (.BL(BL35),.BLN(BLN35),.WL(WL136));
sram_cell_6t_5 inst_cell_136_36 (.BL(BL36),.BLN(BLN36),.WL(WL136));
sram_cell_6t_5 inst_cell_136_37 (.BL(BL37),.BLN(BLN37),.WL(WL136));
sram_cell_6t_5 inst_cell_136_38 (.BL(BL38),.BLN(BLN38),.WL(WL136));
sram_cell_6t_5 inst_cell_136_39 (.BL(BL39),.BLN(BLN39),.WL(WL136));
sram_cell_6t_5 inst_cell_136_40 (.BL(BL40),.BLN(BLN40),.WL(WL136));
sram_cell_6t_5 inst_cell_136_41 (.BL(BL41),.BLN(BLN41),.WL(WL136));
sram_cell_6t_5 inst_cell_136_42 (.BL(BL42),.BLN(BLN42),.WL(WL136));
sram_cell_6t_5 inst_cell_136_43 (.BL(BL43),.BLN(BLN43),.WL(WL136));
sram_cell_6t_5 inst_cell_136_44 (.BL(BL44),.BLN(BLN44),.WL(WL136));
sram_cell_6t_5 inst_cell_136_45 (.BL(BL45),.BLN(BLN45),.WL(WL136));
sram_cell_6t_5 inst_cell_136_46 (.BL(BL46),.BLN(BLN46),.WL(WL136));
sram_cell_6t_5 inst_cell_136_47 (.BL(BL47),.BLN(BLN47),.WL(WL136));
sram_cell_6t_5 inst_cell_136_48 (.BL(BL48),.BLN(BLN48),.WL(WL136));
sram_cell_6t_5 inst_cell_136_49 (.BL(BL49),.BLN(BLN49),.WL(WL136));
sram_cell_6t_5 inst_cell_136_50 (.BL(BL50),.BLN(BLN50),.WL(WL136));
sram_cell_6t_5 inst_cell_136_51 (.BL(BL51),.BLN(BLN51),.WL(WL136));
sram_cell_6t_5 inst_cell_136_52 (.BL(BL52),.BLN(BLN52),.WL(WL136));
sram_cell_6t_5 inst_cell_136_53 (.BL(BL53),.BLN(BLN53),.WL(WL136));
sram_cell_6t_5 inst_cell_136_54 (.BL(BL54),.BLN(BLN54),.WL(WL136));
sram_cell_6t_5 inst_cell_136_55 (.BL(BL55),.BLN(BLN55),.WL(WL136));
sram_cell_6t_5 inst_cell_136_56 (.BL(BL56),.BLN(BLN56),.WL(WL136));
sram_cell_6t_5 inst_cell_136_57 (.BL(BL57),.BLN(BLN57),.WL(WL136));
sram_cell_6t_5 inst_cell_136_58 (.BL(BL58),.BLN(BLN58),.WL(WL136));
sram_cell_6t_5 inst_cell_136_59 (.BL(BL59),.BLN(BLN59),.WL(WL136));
sram_cell_6t_5 inst_cell_136_60 (.BL(BL60),.BLN(BLN60),.WL(WL136));
sram_cell_6t_5 inst_cell_136_61 (.BL(BL61),.BLN(BLN61),.WL(WL136));
sram_cell_6t_5 inst_cell_136_62 (.BL(BL62),.BLN(BLN62),.WL(WL136));
sram_cell_6t_5 inst_cell_136_63 (.BL(BL63),.BLN(BLN63),.WL(WL136));
sram_cell_6t_5 inst_cell_136_64 (.BL(BL64),.BLN(BLN64),.WL(WL136));
sram_cell_6t_5 inst_cell_136_65 (.BL(BL65),.BLN(BLN65),.WL(WL136));
sram_cell_6t_5 inst_cell_136_66 (.BL(BL66),.BLN(BLN66),.WL(WL136));
sram_cell_6t_5 inst_cell_136_67 (.BL(BL67),.BLN(BLN67),.WL(WL136));
sram_cell_6t_5 inst_cell_136_68 (.BL(BL68),.BLN(BLN68),.WL(WL136));
sram_cell_6t_5 inst_cell_136_69 (.BL(BL69),.BLN(BLN69),.WL(WL136));
sram_cell_6t_5 inst_cell_136_70 (.BL(BL70),.BLN(BLN70),.WL(WL136));
sram_cell_6t_5 inst_cell_136_71 (.BL(BL71),.BLN(BLN71),.WL(WL136));
sram_cell_6t_5 inst_cell_136_72 (.BL(BL72),.BLN(BLN72),.WL(WL136));
sram_cell_6t_5 inst_cell_136_73 (.BL(BL73),.BLN(BLN73),.WL(WL136));
sram_cell_6t_5 inst_cell_136_74 (.BL(BL74),.BLN(BLN74),.WL(WL136));
sram_cell_6t_5 inst_cell_136_75 (.BL(BL75),.BLN(BLN75),.WL(WL136));
sram_cell_6t_5 inst_cell_136_76 (.BL(BL76),.BLN(BLN76),.WL(WL136));
sram_cell_6t_5 inst_cell_136_77 (.BL(BL77),.BLN(BLN77),.WL(WL136));
sram_cell_6t_5 inst_cell_136_78 (.BL(BL78),.BLN(BLN78),.WL(WL136));
sram_cell_6t_5 inst_cell_136_79 (.BL(BL79),.BLN(BLN79),.WL(WL136));
sram_cell_6t_5 inst_cell_136_80 (.BL(BL80),.BLN(BLN80),.WL(WL136));
sram_cell_6t_5 inst_cell_136_81 (.BL(BL81),.BLN(BLN81),.WL(WL136));
sram_cell_6t_5 inst_cell_136_82 (.BL(BL82),.BLN(BLN82),.WL(WL136));
sram_cell_6t_5 inst_cell_136_83 (.BL(BL83),.BLN(BLN83),.WL(WL136));
sram_cell_6t_5 inst_cell_136_84 (.BL(BL84),.BLN(BLN84),.WL(WL136));
sram_cell_6t_5 inst_cell_136_85 (.BL(BL85),.BLN(BLN85),.WL(WL136));
sram_cell_6t_5 inst_cell_136_86 (.BL(BL86),.BLN(BLN86),.WL(WL136));
sram_cell_6t_5 inst_cell_136_87 (.BL(BL87),.BLN(BLN87),.WL(WL136));
sram_cell_6t_5 inst_cell_136_88 (.BL(BL88),.BLN(BLN88),.WL(WL136));
sram_cell_6t_5 inst_cell_136_89 (.BL(BL89),.BLN(BLN89),.WL(WL136));
sram_cell_6t_5 inst_cell_136_90 (.BL(BL90),.BLN(BLN90),.WL(WL136));
sram_cell_6t_5 inst_cell_136_91 (.BL(BL91),.BLN(BLN91),.WL(WL136));
sram_cell_6t_5 inst_cell_136_92 (.BL(BL92),.BLN(BLN92),.WL(WL136));
sram_cell_6t_5 inst_cell_136_93 (.BL(BL93),.BLN(BLN93),.WL(WL136));
sram_cell_6t_5 inst_cell_136_94 (.BL(BL94),.BLN(BLN94),.WL(WL136));
sram_cell_6t_5 inst_cell_136_95 (.BL(BL95),.BLN(BLN95),.WL(WL136));
sram_cell_6t_5 inst_cell_136_96 (.BL(BL96),.BLN(BLN96),.WL(WL136));
sram_cell_6t_5 inst_cell_136_97 (.BL(BL97),.BLN(BLN97),.WL(WL136));
sram_cell_6t_5 inst_cell_136_98 (.BL(BL98),.BLN(BLN98),.WL(WL136));
sram_cell_6t_5 inst_cell_136_99 (.BL(BL99),.BLN(BLN99),.WL(WL136));
sram_cell_6t_5 inst_cell_136_100 (.BL(BL100),.BLN(BLN100),.WL(WL136));
sram_cell_6t_5 inst_cell_136_101 (.BL(BL101),.BLN(BLN101),.WL(WL136));
sram_cell_6t_5 inst_cell_136_102 (.BL(BL102),.BLN(BLN102),.WL(WL136));
sram_cell_6t_5 inst_cell_136_103 (.BL(BL103),.BLN(BLN103),.WL(WL136));
sram_cell_6t_5 inst_cell_136_104 (.BL(BL104),.BLN(BLN104),.WL(WL136));
sram_cell_6t_5 inst_cell_136_105 (.BL(BL105),.BLN(BLN105),.WL(WL136));
sram_cell_6t_5 inst_cell_136_106 (.BL(BL106),.BLN(BLN106),.WL(WL136));
sram_cell_6t_5 inst_cell_136_107 (.BL(BL107),.BLN(BLN107),.WL(WL136));
sram_cell_6t_5 inst_cell_136_108 (.BL(BL108),.BLN(BLN108),.WL(WL136));
sram_cell_6t_5 inst_cell_136_109 (.BL(BL109),.BLN(BLN109),.WL(WL136));
sram_cell_6t_5 inst_cell_136_110 (.BL(BL110),.BLN(BLN110),.WL(WL136));
sram_cell_6t_5 inst_cell_136_111 (.BL(BL111),.BLN(BLN111),.WL(WL136));
sram_cell_6t_5 inst_cell_136_112 (.BL(BL112),.BLN(BLN112),.WL(WL136));
sram_cell_6t_5 inst_cell_136_113 (.BL(BL113),.BLN(BLN113),.WL(WL136));
sram_cell_6t_5 inst_cell_136_114 (.BL(BL114),.BLN(BLN114),.WL(WL136));
sram_cell_6t_5 inst_cell_136_115 (.BL(BL115),.BLN(BLN115),.WL(WL136));
sram_cell_6t_5 inst_cell_136_116 (.BL(BL116),.BLN(BLN116),.WL(WL136));
sram_cell_6t_5 inst_cell_136_117 (.BL(BL117),.BLN(BLN117),.WL(WL136));
sram_cell_6t_5 inst_cell_136_118 (.BL(BL118),.BLN(BLN118),.WL(WL136));
sram_cell_6t_5 inst_cell_136_119 (.BL(BL119),.BLN(BLN119),.WL(WL136));
sram_cell_6t_5 inst_cell_136_120 (.BL(BL120),.BLN(BLN120),.WL(WL136));
sram_cell_6t_5 inst_cell_136_121 (.BL(BL121),.BLN(BLN121),.WL(WL136));
sram_cell_6t_5 inst_cell_136_122 (.BL(BL122),.BLN(BLN122),.WL(WL136));
sram_cell_6t_5 inst_cell_136_123 (.BL(BL123),.BLN(BLN123),.WL(WL136));
sram_cell_6t_5 inst_cell_136_124 (.BL(BL124),.BLN(BLN124),.WL(WL136));
sram_cell_6t_5 inst_cell_136_125 (.BL(BL125),.BLN(BLN125),.WL(WL136));
sram_cell_6t_5 inst_cell_136_126 (.BL(BL126),.BLN(BLN126),.WL(WL136));
sram_cell_6t_5 inst_cell_136_127 (.BL(BL127),.BLN(BLN127),.WL(WL136));
sram_cell_6t_5 inst_cell_137_0 (.BL(BL0),.BLN(BLN0),.WL(WL137));
sram_cell_6t_5 inst_cell_137_1 (.BL(BL1),.BLN(BLN1),.WL(WL137));
sram_cell_6t_5 inst_cell_137_2 (.BL(BL2),.BLN(BLN2),.WL(WL137));
sram_cell_6t_5 inst_cell_137_3 (.BL(BL3),.BLN(BLN3),.WL(WL137));
sram_cell_6t_5 inst_cell_137_4 (.BL(BL4),.BLN(BLN4),.WL(WL137));
sram_cell_6t_5 inst_cell_137_5 (.BL(BL5),.BLN(BLN5),.WL(WL137));
sram_cell_6t_5 inst_cell_137_6 (.BL(BL6),.BLN(BLN6),.WL(WL137));
sram_cell_6t_5 inst_cell_137_7 (.BL(BL7),.BLN(BLN7),.WL(WL137));
sram_cell_6t_5 inst_cell_137_8 (.BL(BL8),.BLN(BLN8),.WL(WL137));
sram_cell_6t_5 inst_cell_137_9 (.BL(BL9),.BLN(BLN9),.WL(WL137));
sram_cell_6t_5 inst_cell_137_10 (.BL(BL10),.BLN(BLN10),.WL(WL137));
sram_cell_6t_5 inst_cell_137_11 (.BL(BL11),.BLN(BLN11),.WL(WL137));
sram_cell_6t_5 inst_cell_137_12 (.BL(BL12),.BLN(BLN12),.WL(WL137));
sram_cell_6t_5 inst_cell_137_13 (.BL(BL13),.BLN(BLN13),.WL(WL137));
sram_cell_6t_5 inst_cell_137_14 (.BL(BL14),.BLN(BLN14),.WL(WL137));
sram_cell_6t_5 inst_cell_137_15 (.BL(BL15),.BLN(BLN15),.WL(WL137));
sram_cell_6t_5 inst_cell_137_16 (.BL(BL16),.BLN(BLN16),.WL(WL137));
sram_cell_6t_5 inst_cell_137_17 (.BL(BL17),.BLN(BLN17),.WL(WL137));
sram_cell_6t_5 inst_cell_137_18 (.BL(BL18),.BLN(BLN18),.WL(WL137));
sram_cell_6t_5 inst_cell_137_19 (.BL(BL19),.BLN(BLN19),.WL(WL137));
sram_cell_6t_5 inst_cell_137_20 (.BL(BL20),.BLN(BLN20),.WL(WL137));
sram_cell_6t_5 inst_cell_137_21 (.BL(BL21),.BLN(BLN21),.WL(WL137));
sram_cell_6t_5 inst_cell_137_22 (.BL(BL22),.BLN(BLN22),.WL(WL137));
sram_cell_6t_5 inst_cell_137_23 (.BL(BL23),.BLN(BLN23),.WL(WL137));
sram_cell_6t_5 inst_cell_137_24 (.BL(BL24),.BLN(BLN24),.WL(WL137));
sram_cell_6t_5 inst_cell_137_25 (.BL(BL25),.BLN(BLN25),.WL(WL137));
sram_cell_6t_5 inst_cell_137_26 (.BL(BL26),.BLN(BLN26),.WL(WL137));
sram_cell_6t_5 inst_cell_137_27 (.BL(BL27),.BLN(BLN27),.WL(WL137));
sram_cell_6t_5 inst_cell_137_28 (.BL(BL28),.BLN(BLN28),.WL(WL137));
sram_cell_6t_5 inst_cell_137_29 (.BL(BL29),.BLN(BLN29),.WL(WL137));
sram_cell_6t_5 inst_cell_137_30 (.BL(BL30),.BLN(BLN30),.WL(WL137));
sram_cell_6t_5 inst_cell_137_31 (.BL(BL31),.BLN(BLN31),.WL(WL137));
sram_cell_6t_5 inst_cell_137_32 (.BL(BL32),.BLN(BLN32),.WL(WL137));
sram_cell_6t_5 inst_cell_137_33 (.BL(BL33),.BLN(BLN33),.WL(WL137));
sram_cell_6t_5 inst_cell_137_34 (.BL(BL34),.BLN(BLN34),.WL(WL137));
sram_cell_6t_5 inst_cell_137_35 (.BL(BL35),.BLN(BLN35),.WL(WL137));
sram_cell_6t_5 inst_cell_137_36 (.BL(BL36),.BLN(BLN36),.WL(WL137));
sram_cell_6t_5 inst_cell_137_37 (.BL(BL37),.BLN(BLN37),.WL(WL137));
sram_cell_6t_5 inst_cell_137_38 (.BL(BL38),.BLN(BLN38),.WL(WL137));
sram_cell_6t_5 inst_cell_137_39 (.BL(BL39),.BLN(BLN39),.WL(WL137));
sram_cell_6t_5 inst_cell_137_40 (.BL(BL40),.BLN(BLN40),.WL(WL137));
sram_cell_6t_5 inst_cell_137_41 (.BL(BL41),.BLN(BLN41),.WL(WL137));
sram_cell_6t_5 inst_cell_137_42 (.BL(BL42),.BLN(BLN42),.WL(WL137));
sram_cell_6t_5 inst_cell_137_43 (.BL(BL43),.BLN(BLN43),.WL(WL137));
sram_cell_6t_5 inst_cell_137_44 (.BL(BL44),.BLN(BLN44),.WL(WL137));
sram_cell_6t_5 inst_cell_137_45 (.BL(BL45),.BLN(BLN45),.WL(WL137));
sram_cell_6t_5 inst_cell_137_46 (.BL(BL46),.BLN(BLN46),.WL(WL137));
sram_cell_6t_5 inst_cell_137_47 (.BL(BL47),.BLN(BLN47),.WL(WL137));
sram_cell_6t_5 inst_cell_137_48 (.BL(BL48),.BLN(BLN48),.WL(WL137));
sram_cell_6t_5 inst_cell_137_49 (.BL(BL49),.BLN(BLN49),.WL(WL137));
sram_cell_6t_5 inst_cell_137_50 (.BL(BL50),.BLN(BLN50),.WL(WL137));
sram_cell_6t_5 inst_cell_137_51 (.BL(BL51),.BLN(BLN51),.WL(WL137));
sram_cell_6t_5 inst_cell_137_52 (.BL(BL52),.BLN(BLN52),.WL(WL137));
sram_cell_6t_5 inst_cell_137_53 (.BL(BL53),.BLN(BLN53),.WL(WL137));
sram_cell_6t_5 inst_cell_137_54 (.BL(BL54),.BLN(BLN54),.WL(WL137));
sram_cell_6t_5 inst_cell_137_55 (.BL(BL55),.BLN(BLN55),.WL(WL137));
sram_cell_6t_5 inst_cell_137_56 (.BL(BL56),.BLN(BLN56),.WL(WL137));
sram_cell_6t_5 inst_cell_137_57 (.BL(BL57),.BLN(BLN57),.WL(WL137));
sram_cell_6t_5 inst_cell_137_58 (.BL(BL58),.BLN(BLN58),.WL(WL137));
sram_cell_6t_5 inst_cell_137_59 (.BL(BL59),.BLN(BLN59),.WL(WL137));
sram_cell_6t_5 inst_cell_137_60 (.BL(BL60),.BLN(BLN60),.WL(WL137));
sram_cell_6t_5 inst_cell_137_61 (.BL(BL61),.BLN(BLN61),.WL(WL137));
sram_cell_6t_5 inst_cell_137_62 (.BL(BL62),.BLN(BLN62),.WL(WL137));
sram_cell_6t_5 inst_cell_137_63 (.BL(BL63),.BLN(BLN63),.WL(WL137));
sram_cell_6t_5 inst_cell_137_64 (.BL(BL64),.BLN(BLN64),.WL(WL137));
sram_cell_6t_5 inst_cell_137_65 (.BL(BL65),.BLN(BLN65),.WL(WL137));
sram_cell_6t_5 inst_cell_137_66 (.BL(BL66),.BLN(BLN66),.WL(WL137));
sram_cell_6t_5 inst_cell_137_67 (.BL(BL67),.BLN(BLN67),.WL(WL137));
sram_cell_6t_5 inst_cell_137_68 (.BL(BL68),.BLN(BLN68),.WL(WL137));
sram_cell_6t_5 inst_cell_137_69 (.BL(BL69),.BLN(BLN69),.WL(WL137));
sram_cell_6t_5 inst_cell_137_70 (.BL(BL70),.BLN(BLN70),.WL(WL137));
sram_cell_6t_5 inst_cell_137_71 (.BL(BL71),.BLN(BLN71),.WL(WL137));
sram_cell_6t_5 inst_cell_137_72 (.BL(BL72),.BLN(BLN72),.WL(WL137));
sram_cell_6t_5 inst_cell_137_73 (.BL(BL73),.BLN(BLN73),.WL(WL137));
sram_cell_6t_5 inst_cell_137_74 (.BL(BL74),.BLN(BLN74),.WL(WL137));
sram_cell_6t_5 inst_cell_137_75 (.BL(BL75),.BLN(BLN75),.WL(WL137));
sram_cell_6t_5 inst_cell_137_76 (.BL(BL76),.BLN(BLN76),.WL(WL137));
sram_cell_6t_5 inst_cell_137_77 (.BL(BL77),.BLN(BLN77),.WL(WL137));
sram_cell_6t_5 inst_cell_137_78 (.BL(BL78),.BLN(BLN78),.WL(WL137));
sram_cell_6t_5 inst_cell_137_79 (.BL(BL79),.BLN(BLN79),.WL(WL137));
sram_cell_6t_5 inst_cell_137_80 (.BL(BL80),.BLN(BLN80),.WL(WL137));
sram_cell_6t_5 inst_cell_137_81 (.BL(BL81),.BLN(BLN81),.WL(WL137));
sram_cell_6t_5 inst_cell_137_82 (.BL(BL82),.BLN(BLN82),.WL(WL137));
sram_cell_6t_5 inst_cell_137_83 (.BL(BL83),.BLN(BLN83),.WL(WL137));
sram_cell_6t_5 inst_cell_137_84 (.BL(BL84),.BLN(BLN84),.WL(WL137));
sram_cell_6t_5 inst_cell_137_85 (.BL(BL85),.BLN(BLN85),.WL(WL137));
sram_cell_6t_5 inst_cell_137_86 (.BL(BL86),.BLN(BLN86),.WL(WL137));
sram_cell_6t_5 inst_cell_137_87 (.BL(BL87),.BLN(BLN87),.WL(WL137));
sram_cell_6t_5 inst_cell_137_88 (.BL(BL88),.BLN(BLN88),.WL(WL137));
sram_cell_6t_5 inst_cell_137_89 (.BL(BL89),.BLN(BLN89),.WL(WL137));
sram_cell_6t_5 inst_cell_137_90 (.BL(BL90),.BLN(BLN90),.WL(WL137));
sram_cell_6t_5 inst_cell_137_91 (.BL(BL91),.BLN(BLN91),.WL(WL137));
sram_cell_6t_5 inst_cell_137_92 (.BL(BL92),.BLN(BLN92),.WL(WL137));
sram_cell_6t_5 inst_cell_137_93 (.BL(BL93),.BLN(BLN93),.WL(WL137));
sram_cell_6t_5 inst_cell_137_94 (.BL(BL94),.BLN(BLN94),.WL(WL137));
sram_cell_6t_5 inst_cell_137_95 (.BL(BL95),.BLN(BLN95),.WL(WL137));
sram_cell_6t_5 inst_cell_137_96 (.BL(BL96),.BLN(BLN96),.WL(WL137));
sram_cell_6t_5 inst_cell_137_97 (.BL(BL97),.BLN(BLN97),.WL(WL137));
sram_cell_6t_5 inst_cell_137_98 (.BL(BL98),.BLN(BLN98),.WL(WL137));
sram_cell_6t_5 inst_cell_137_99 (.BL(BL99),.BLN(BLN99),.WL(WL137));
sram_cell_6t_5 inst_cell_137_100 (.BL(BL100),.BLN(BLN100),.WL(WL137));
sram_cell_6t_5 inst_cell_137_101 (.BL(BL101),.BLN(BLN101),.WL(WL137));
sram_cell_6t_5 inst_cell_137_102 (.BL(BL102),.BLN(BLN102),.WL(WL137));
sram_cell_6t_5 inst_cell_137_103 (.BL(BL103),.BLN(BLN103),.WL(WL137));
sram_cell_6t_5 inst_cell_137_104 (.BL(BL104),.BLN(BLN104),.WL(WL137));
sram_cell_6t_5 inst_cell_137_105 (.BL(BL105),.BLN(BLN105),.WL(WL137));
sram_cell_6t_5 inst_cell_137_106 (.BL(BL106),.BLN(BLN106),.WL(WL137));
sram_cell_6t_5 inst_cell_137_107 (.BL(BL107),.BLN(BLN107),.WL(WL137));
sram_cell_6t_5 inst_cell_137_108 (.BL(BL108),.BLN(BLN108),.WL(WL137));
sram_cell_6t_5 inst_cell_137_109 (.BL(BL109),.BLN(BLN109),.WL(WL137));
sram_cell_6t_5 inst_cell_137_110 (.BL(BL110),.BLN(BLN110),.WL(WL137));
sram_cell_6t_5 inst_cell_137_111 (.BL(BL111),.BLN(BLN111),.WL(WL137));
sram_cell_6t_5 inst_cell_137_112 (.BL(BL112),.BLN(BLN112),.WL(WL137));
sram_cell_6t_5 inst_cell_137_113 (.BL(BL113),.BLN(BLN113),.WL(WL137));
sram_cell_6t_5 inst_cell_137_114 (.BL(BL114),.BLN(BLN114),.WL(WL137));
sram_cell_6t_5 inst_cell_137_115 (.BL(BL115),.BLN(BLN115),.WL(WL137));
sram_cell_6t_5 inst_cell_137_116 (.BL(BL116),.BLN(BLN116),.WL(WL137));
sram_cell_6t_5 inst_cell_137_117 (.BL(BL117),.BLN(BLN117),.WL(WL137));
sram_cell_6t_5 inst_cell_137_118 (.BL(BL118),.BLN(BLN118),.WL(WL137));
sram_cell_6t_5 inst_cell_137_119 (.BL(BL119),.BLN(BLN119),.WL(WL137));
sram_cell_6t_5 inst_cell_137_120 (.BL(BL120),.BLN(BLN120),.WL(WL137));
sram_cell_6t_5 inst_cell_137_121 (.BL(BL121),.BLN(BLN121),.WL(WL137));
sram_cell_6t_5 inst_cell_137_122 (.BL(BL122),.BLN(BLN122),.WL(WL137));
sram_cell_6t_5 inst_cell_137_123 (.BL(BL123),.BLN(BLN123),.WL(WL137));
sram_cell_6t_5 inst_cell_137_124 (.BL(BL124),.BLN(BLN124),.WL(WL137));
sram_cell_6t_5 inst_cell_137_125 (.BL(BL125),.BLN(BLN125),.WL(WL137));
sram_cell_6t_5 inst_cell_137_126 (.BL(BL126),.BLN(BLN126),.WL(WL137));
sram_cell_6t_5 inst_cell_137_127 (.BL(BL127),.BLN(BLN127),.WL(WL137));
sram_cell_6t_5 inst_cell_138_0 (.BL(BL0),.BLN(BLN0),.WL(WL138));
sram_cell_6t_5 inst_cell_138_1 (.BL(BL1),.BLN(BLN1),.WL(WL138));
sram_cell_6t_5 inst_cell_138_2 (.BL(BL2),.BLN(BLN2),.WL(WL138));
sram_cell_6t_5 inst_cell_138_3 (.BL(BL3),.BLN(BLN3),.WL(WL138));
sram_cell_6t_5 inst_cell_138_4 (.BL(BL4),.BLN(BLN4),.WL(WL138));
sram_cell_6t_5 inst_cell_138_5 (.BL(BL5),.BLN(BLN5),.WL(WL138));
sram_cell_6t_5 inst_cell_138_6 (.BL(BL6),.BLN(BLN6),.WL(WL138));
sram_cell_6t_5 inst_cell_138_7 (.BL(BL7),.BLN(BLN7),.WL(WL138));
sram_cell_6t_5 inst_cell_138_8 (.BL(BL8),.BLN(BLN8),.WL(WL138));
sram_cell_6t_5 inst_cell_138_9 (.BL(BL9),.BLN(BLN9),.WL(WL138));
sram_cell_6t_5 inst_cell_138_10 (.BL(BL10),.BLN(BLN10),.WL(WL138));
sram_cell_6t_5 inst_cell_138_11 (.BL(BL11),.BLN(BLN11),.WL(WL138));
sram_cell_6t_5 inst_cell_138_12 (.BL(BL12),.BLN(BLN12),.WL(WL138));
sram_cell_6t_5 inst_cell_138_13 (.BL(BL13),.BLN(BLN13),.WL(WL138));
sram_cell_6t_5 inst_cell_138_14 (.BL(BL14),.BLN(BLN14),.WL(WL138));
sram_cell_6t_5 inst_cell_138_15 (.BL(BL15),.BLN(BLN15),.WL(WL138));
sram_cell_6t_5 inst_cell_138_16 (.BL(BL16),.BLN(BLN16),.WL(WL138));
sram_cell_6t_5 inst_cell_138_17 (.BL(BL17),.BLN(BLN17),.WL(WL138));
sram_cell_6t_5 inst_cell_138_18 (.BL(BL18),.BLN(BLN18),.WL(WL138));
sram_cell_6t_5 inst_cell_138_19 (.BL(BL19),.BLN(BLN19),.WL(WL138));
sram_cell_6t_5 inst_cell_138_20 (.BL(BL20),.BLN(BLN20),.WL(WL138));
sram_cell_6t_5 inst_cell_138_21 (.BL(BL21),.BLN(BLN21),.WL(WL138));
sram_cell_6t_5 inst_cell_138_22 (.BL(BL22),.BLN(BLN22),.WL(WL138));
sram_cell_6t_5 inst_cell_138_23 (.BL(BL23),.BLN(BLN23),.WL(WL138));
sram_cell_6t_5 inst_cell_138_24 (.BL(BL24),.BLN(BLN24),.WL(WL138));
sram_cell_6t_5 inst_cell_138_25 (.BL(BL25),.BLN(BLN25),.WL(WL138));
sram_cell_6t_5 inst_cell_138_26 (.BL(BL26),.BLN(BLN26),.WL(WL138));
sram_cell_6t_5 inst_cell_138_27 (.BL(BL27),.BLN(BLN27),.WL(WL138));
sram_cell_6t_5 inst_cell_138_28 (.BL(BL28),.BLN(BLN28),.WL(WL138));
sram_cell_6t_5 inst_cell_138_29 (.BL(BL29),.BLN(BLN29),.WL(WL138));
sram_cell_6t_5 inst_cell_138_30 (.BL(BL30),.BLN(BLN30),.WL(WL138));
sram_cell_6t_5 inst_cell_138_31 (.BL(BL31),.BLN(BLN31),.WL(WL138));
sram_cell_6t_5 inst_cell_138_32 (.BL(BL32),.BLN(BLN32),.WL(WL138));
sram_cell_6t_5 inst_cell_138_33 (.BL(BL33),.BLN(BLN33),.WL(WL138));
sram_cell_6t_5 inst_cell_138_34 (.BL(BL34),.BLN(BLN34),.WL(WL138));
sram_cell_6t_5 inst_cell_138_35 (.BL(BL35),.BLN(BLN35),.WL(WL138));
sram_cell_6t_5 inst_cell_138_36 (.BL(BL36),.BLN(BLN36),.WL(WL138));
sram_cell_6t_5 inst_cell_138_37 (.BL(BL37),.BLN(BLN37),.WL(WL138));
sram_cell_6t_5 inst_cell_138_38 (.BL(BL38),.BLN(BLN38),.WL(WL138));
sram_cell_6t_5 inst_cell_138_39 (.BL(BL39),.BLN(BLN39),.WL(WL138));
sram_cell_6t_5 inst_cell_138_40 (.BL(BL40),.BLN(BLN40),.WL(WL138));
sram_cell_6t_5 inst_cell_138_41 (.BL(BL41),.BLN(BLN41),.WL(WL138));
sram_cell_6t_5 inst_cell_138_42 (.BL(BL42),.BLN(BLN42),.WL(WL138));
sram_cell_6t_5 inst_cell_138_43 (.BL(BL43),.BLN(BLN43),.WL(WL138));
sram_cell_6t_5 inst_cell_138_44 (.BL(BL44),.BLN(BLN44),.WL(WL138));
sram_cell_6t_5 inst_cell_138_45 (.BL(BL45),.BLN(BLN45),.WL(WL138));
sram_cell_6t_5 inst_cell_138_46 (.BL(BL46),.BLN(BLN46),.WL(WL138));
sram_cell_6t_5 inst_cell_138_47 (.BL(BL47),.BLN(BLN47),.WL(WL138));
sram_cell_6t_5 inst_cell_138_48 (.BL(BL48),.BLN(BLN48),.WL(WL138));
sram_cell_6t_5 inst_cell_138_49 (.BL(BL49),.BLN(BLN49),.WL(WL138));
sram_cell_6t_5 inst_cell_138_50 (.BL(BL50),.BLN(BLN50),.WL(WL138));
sram_cell_6t_5 inst_cell_138_51 (.BL(BL51),.BLN(BLN51),.WL(WL138));
sram_cell_6t_5 inst_cell_138_52 (.BL(BL52),.BLN(BLN52),.WL(WL138));
sram_cell_6t_5 inst_cell_138_53 (.BL(BL53),.BLN(BLN53),.WL(WL138));
sram_cell_6t_5 inst_cell_138_54 (.BL(BL54),.BLN(BLN54),.WL(WL138));
sram_cell_6t_5 inst_cell_138_55 (.BL(BL55),.BLN(BLN55),.WL(WL138));
sram_cell_6t_5 inst_cell_138_56 (.BL(BL56),.BLN(BLN56),.WL(WL138));
sram_cell_6t_5 inst_cell_138_57 (.BL(BL57),.BLN(BLN57),.WL(WL138));
sram_cell_6t_5 inst_cell_138_58 (.BL(BL58),.BLN(BLN58),.WL(WL138));
sram_cell_6t_5 inst_cell_138_59 (.BL(BL59),.BLN(BLN59),.WL(WL138));
sram_cell_6t_5 inst_cell_138_60 (.BL(BL60),.BLN(BLN60),.WL(WL138));
sram_cell_6t_5 inst_cell_138_61 (.BL(BL61),.BLN(BLN61),.WL(WL138));
sram_cell_6t_5 inst_cell_138_62 (.BL(BL62),.BLN(BLN62),.WL(WL138));
sram_cell_6t_5 inst_cell_138_63 (.BL(BL63),.BLN(BLN63),.WL(WL138));
sram_cell_6t_5 inst_cell_138_64 (.BL(BL64),.BLN(BLN64),.WL(WL138));
sram_cell_6t_5 inst_cell_138_65 (.BL(BL65),.BLN(BLN65),.WL(WL138));
sram_cell_6t_5 inst_cell_138_66 (.BL(BL66),.BLN(BLN66),.WL(WL138));
sram_cell_6t_5 inst_cell_138_67 (.BL(BL67),.BLN(BLN67),.WL(WL138));
sram_cell_6t_5 inst_cell_138_68 (.BL(BL68),.BLN(BLN68),.WL(WL138));
sram_cell_6t_5 inst_cell_138_69 (.BL(BL69),.BLN(BLN69),.WL(WL138));
sram_cell_6t_5 inst_cell_138_70 (.BL(BL70),.BLN(BLN70),.WL(WL138));
sram_cell_6t_5 inst_cell_138_71 (.BL(BL71),.BLN(BLN71),.WL(WL138));
sram_cell_6t_5 inst_cell_138_72 (.BL(BL72),.BLN(BLN72),.WL(WL138));
sram_cell_6t_5 inst_cell_138_73 (.BL(BL73),.BLN(BLN73),.WL(WL138));
sram_cell_6t_5 inst_cell_138_74 (.BL(BL74),.BLN(BLN74),.WL(WL138));
sram_cell_6t_5 inst_cell_138_75 (.BL(BL75),.BLN(BLN75),.WL(WL138));
sram_cell_6t_5 inst_cell_138_76 (.BL(BL76),.BLN(BLN76),.WL(WL138));
sram_cell_6t_5 inst_cell_138_77 (.BL(BL77),.BLN(BLN77),.WL(WL138));
sram_cell_6t_5 inst_cell_138_78 (.BL(BL78),.BLN(BLN78),.WL(WL138));
sram_cell_6t_5 inst_cell_138_79 (.BL(BL79),.BLN(BLN79),.WL(WL138));
sram_cell_6t_5 inst_cell_138_80 (.BL(BL80),.BLN(BLN80),.WL(WL138));
sram_cell_6t_5 inst_cell_138_81 (.BL(BL81),.BLN(BLN81),.WL(WL138));
sram_cell_6t_5 inst_cell_138_82 (.BL(BL82),.BLN(BLN82),.WL(WL138));
sram_cell_6t_5 inst_cell_138_83 (.BL(BL83),.BLN(BLN83),.WL(WL138));
sram_cell_6t_5 inst_cell_138_84 (.BL(BL84),.BLN(BLN84),.WL(WL138));
sram_cell_6t_5 inst_cell_138_85 (.BL(BL85),.BLN(BLN85),.WL(WL138));
sram_cell_6t_5 inst_cell_138_86 (.BL(BL86),.BLN(BLN86),.WL(WL138));
sram_cell_6t_5 inst_cell_138_87 (.BL(BL87),.BLN(BLN87),.WL(WL138));
sram_cell_6t_5 inst_cell_138_88 (.BL(BL88),.BLN(BLN88),.WL(WL138));
sram_cell_6t_5 inst_cell_138_89 (.BL(BL89),.BLN(BLN89),.WL(WL138));
sram_cell_6t_5 inst_cell_138_90 (.BL(BL90),.BLN(BLN90),.WL(WL138));
sram_cell_6t_5 inst_cell_138_91 (.BL(BL91),.BLN(BLN91),.WL(WL138));
sram_cell_6t_5 inst_cell_138_92 (.BL(BL92),.BLN(BLN92),.WL(WL138));
sram_cell_6t_5 inst_cell_138_93 (.BL(BL93),.BLN(BLN93),.WL(WL138));
sram_cell_6t_5 inst_cell_138_94 (.BL(BL94),.BLN(BLN94),.WL(WL138));
sram_cell_6t_5 inst_cell_138_95 (.BL(BL95),.BLN(BLN95),.WL(WL138));
sram_cell_6t_5 inst_cell_138_96 (.BL(BL96),.BLN(BLN96),.WL(WL138));
sram_cell_6t_5 inst_cell_138_97 (.BL(BL97),.BLN(BLN97),.WL(WL138));
sram_cell_6t_5 inst_cell_138_98 (.BL(BL98),.BLN(BLN98),.WL(WL138));
sram_cell_6t_5 inst_cell_138_99 (.BL(BL99),.BLN(BLN99),.WL(WL138));
sram_cell_6t_5 inst_cell_138_100 (.BL(BL100),.BLN(BLN100),.WL(WL138));
sram_cell_6t_5 inst_cell_138_101 (.BL(BL101),.BLN(BLN101),.WL(WL138));
sram_cell_6t_5 inst_cell_138_102 (.BL(BL102),.BLN(BLN102),.WL(WL138));
sram_cell_6t_5 inst_cell_138_103 (.BL(BL103),.BLN(BLN103),.WL(WL138));
sram_cell_6t_5 inst_cell_138_104 (.BL(BL104),.BLN(BLN104),.WL(WL138));
sram_cell_6t_5 inst_cell_138_105 (.BL(BL105),.BLN(BLN105),.WL(WL138));
sram_cell_6t_5 inst_cell_138_106 (.BL(BL106),.BLN(BLN106),.WL(WL138));
sram_cell_6t_5 inst_cell_138_107 (.BL(BL107),.BLN(BLN107),.WL(WL138));
sram_cell_6t_5 inst_cell_138_108 (.BL(BL108),.BLN(BLN108),.WL(WL138));
sram_cell_6t_5 inst_cell_138_109 (.BL(BL109),.BLN(BLN109),.WL(WL138));
sram_cell_6t_5 inst_cell_138_110 (.BL(BL110),.BLN(BLN110),.WL(WL138));
sram_cell_6t_5 inst_cell_138_111 (.BL(BL111),.BLN(BLN111),.WL(WL138));
sram_cell_6t_5 inst_cell_138_112 (.BL(BL112),.BLN(BLN112),.WL(WL138));
sram_cell_6t_5 inst_cell_138_113 (.BL(BL113),.BLN(BLN113),.WL(WL138));
sram_cell_6t_5 inst_cell_138_114 (.BL(BL114),.BLN(BLN114),.WL(WL138));
sram_cell_6t_5 inst_cell_138_115 (.BL(BL115),.BLN(BLN115),.WL(WL138));
sram_cell_6t_5 inst_cell_138_116 (.BL(BL116),.BLN(BLN116),.WL(WL138));
sram_cell_6t_5 inst_cell_138_117 (.BL(BL117),.BLN(BLN117),.WL(WL138));
sram_cell_6t_5 inst_cell_138_118 (.BL(BL118),.BLN(BLN118),.WL(WL138));
sram_cell_6t_5 inst_cell_138_119 (.BL(BL119),.BLN(BLN119),.WL(WL138));
sram_cell_6t_5 inst_cell_138_120 (.BL(BL120),.BLN(BLN120),.WL(WL138));
sram_cell_6t_5 inst_cell_138_121 (.BL(BL121),.BLN(BLN121),.WL(WL138));
sram_cell_6t_5 inst_cell_138_122 (.BL(BL122),.BLN(BLN122),.WL(WL138));
sram_cell_6t_5 inst_cell_138_123 (.BL(BL123),.BLN(BLN123),.WL(WL138));
sram_cell_6t_5 inst_cell_138_124 (.BL(BL124),.BLN(BLN124),.WL(WL138));
sram_cell_6t_5 inst_cell_138_125 (.BL(BL125),.BLN(BLN125),.WL(WL138));
sram_cell_6t_5 inst_cell_138_126 (.BL(BL126),.BLN(BLN126),.WL(WL138));
sram_cell_6t_5 inst_cell_138_127 (.BL(BL127),.BLN(BLN127),.WL(WL138));
sram_cell_6t_5 inst_cell_139_0 (.BL(BL0),.BLN(BLN0),.WL(WL139));
sram_cell_6t_5 inst_cell_139_1 (.BL(BL1),.BLN(BLN1),.WL(WL139));
sram_cell_6t_5 inst_cell_139_2 (.BL(BL2),.BLN(BLN2),.WL(WL139));
sram_cell_6t_5 inst_cell_139_3 (.BL(BL3),.BLN(BLN3),.WL(WL139));
sram_cell_6t_5 inst_cell_139_4 (.BL(BL4),.BLN(BLN4),.WL(WL139));
sram_cell_6t_5 inst_cell_139_5 (.BL(BL5),.BLN(BLN5),.WL(WL139));
sram_cell_6t_5 inst_cell_139_6 (.BL(BL6),.BLN(BLN6),.WL(WL139));
sram_cell_6t_5 inst_cell_139_7 (.BL(BL7),.BLN(BLN7),.WL(WL139));
sram_cell_6t_5 inst_cell_139_8 (.BL(BL8),.BLN(BLN8),.WL(WL139));
sram_cell_6t_5 inst_cell_139_9 (.BL(BL9),.BLN(BLN9),.WL(WL139));
sram_cell_6t_5 inst_cell_139_10 (.BL(BL10),.BLN(BLN10),.WL(WL139));
sram_cell_6t_5 inst_cell_139_11 (.BL(BL11),.BLN(BLN11),.WL(WL139));
sram_cell_6t_5 inst_cell_139_12 (.BL(BL12),.BLN(BLN12),.WL(WL139));
sram_cell_6t_5 inst_cell_139_13 (.BL(BL13),.BLN(BLN13),.WL(WL139));
sram_cell_6t_5 inst_cell_139_14 (.BL(BL14),.BLN(BLN14),.WL(WL139));
sram_cell_6t_5 inst_cell_139_15 (.BL(BL15),.BLN(BLN15),.WL(WL139));
sram_cell_6t_5 inst_cell_139_16 (.BL(BL16),.BLN(BLN16),.WL(WL139));
sram_cell_6t_5 inst_cell_139_17 (.BL(BL17),.BLN(BLN17),.WL(WL139));
sram_cell_6t_5 inst_cell_139_18 (.BL(BL18),.BLN(BLN18),.WL(WL139));
sram_cell_6t_5 inst_cell_139_19 (.BL(BL19),.BLN(BLN19),.WL(WL139));
sram_cell_6t_5 inst_cell_139_20 (.BL(BL20),.BLN(BLN20),.WL(WL139));
sram_cell_6t_5 inst_cell_139_21 (.BL(BL21),.BLN(BLN21),.WL(WL139));
sram_cell_6t_5 inst_cell_139_22 (.BL(BL22),.BLN(BLN22),.WL(WL139));
sram_cell_6t_5 inst_cell_139_23 (.BL(BL23),.BLN(BLN23),.WL(WL139));
sram_cell_6t_5 inst_cell_139_24 (.BL(BL24),.BLN(BLN24),.WL(WL139));
sram_cell_6t_5 inst_cell_139_25 (.BL(BL25),.BLN(BLN25),.WL(WL139));
sram_cell_6t_5 inst_cell_139_26 (.BL(BL26),.BLN(BLN26),.WL(WL139));
sram_cell_6t_5 inst_cell_139_27 (.BL(BL27),.BLN(BLN27),.WL(WL139));
sram_cell_6t_5 inst_cell_139_28 (.BL(BL28),.BLN(BLN28),.WL(WL139));
sram_cell_6t_5 inst_cell_139_29 (.BL(BL29),.BLN(BLN29),.WL(WL139));
sram_cell_6t_5 inst_cell_139_30 (.BL(BL30),.BLN(BLN30),.WL(WL139));
sram_cell_6t_5 inst_cell_139_31 (.BL(BL31),.BLN(BLN31),.WL(WL139));
sram_cell_6t_5 inst_cell_139_32 (.BL(BL32),.BLN(BLN32),.WL(WL139));
sram_cell_6t_5 inst_cell_139_33 (.BL(BL33),.BLN(BLN33),.WL(WL139));
sram_cell_6t_5 inst_cell_139_34 (.BL(BL34),.BLN(BLN34),.WL(WL139));
sram_cell_6t_5 inst_cell_139_35 (.BL(BL35),.BLN(BLN35),.WL(WL139));
sram_cell_6t_5 inst_cell_139_36 (.BL(BL36),.BLN(BLN36),.WL(WL139));
sram_cell_6t_5 inst_cell_139_37 (.BL(BL37),.BLN(BLN37),.WL(WL139));
sram_cell_6t_5 inst_cell_139_38 (.BL(BL38),.BLN(BLN38),.WL(WL139));
sram_cell_6t_5 inst_cell_139_39 (.BL(BL39),.BLN(BLN39),.WL(WL139));
sram_cell_6t_5 inst_cell_139_40 (.BL(BL40),.BLN(BLN40),.WL(WL139));
sram_cell_6t_5 inst_cell_139_41 (.BL(BL41),.BLN(BLN41),.WL(WL139));
sram_cell_6t_5 inst_cell_139_42 (.BL(BL42),.BLN(BLN42),.WL(WL139));
sram_cell_6t_5 inst_cell_139_43 (.BL(BL43),.BLN(BLN43),.WL(WL139));
sram_cell_6t_5 inst_cell_139_44 (.BL(BL44),.BLN(BLN44),.WL(WL139));
sram_cell_6t_5 inst_cell_139_45 (.BL(BL45),.BLN(BLN45),.WL(WL139));
sram_cell_6t_5 inst_cell_139_46 (.BL(BL46),.BLN(BLN46),.WL(WL139));
sram_cell_6t_5 inst_cell_139_47 (.BL(BL47),.BLN(BLN47),.WL(WL139));
sram_cell_6t_5 inst_cell_139_48 (.BL(BL48),.BLN(BLN48),.WL(WL139));
sram_cell_6t_5 inst_cell_139_49 (.BL(BL49),.BLN(BLN49),.WL(WL139));
sram_cell_6t_5 inst_cell_139_50 (.BL(BL50),.BLN(BLN50),.WL(WL139));
sram_cell_6t_5 inst_cell_139_51 (.BL(BL51),.BLN(BLN51),.WL(WL139));
sram_cell_6t_5 inst_cell_139_52 (.BL(BL52),.BLN(BLN52),.WL(WL139));
sram_cell_6t_5 inst_cell_139_53 (.BL(BL53),.BLN(BLN53),.WL(WL139));
sram_cell_6t_5 inst_cell_139_54 (.BL(BL54),.BLN(BLN54),.WL(WL139));
sram_cell_6t_5 inst_cell_139_55 (.BL(BL55),.BLN(BLN55),.WL(WL139));
sram_cell_6t_5 inst_cell_139_56 (.BL(BL56),.BLN(BLN56),.WL(WL139));
sram_cell_6t_5 inst_cell_139_57 (.BL(BL57),.BLN(BLN57),.WL(WL139));
sram_cell_6t_5 inst_cell_139_58 (.BL(BL58),.BLN(BLN58),.WL(WL139));
sram_cell_6t_5 inst_cell_139_59 (.BL(BL59),.BLN(BLN59),.WL(WL139));
sram_cell_6t_5 inst_cell_139_60 (.BL(BL60),.BLN(BLN60),.WL(WL139));
sram_cell_6t_5 inst_cell_139_61 (.BL(BL61),.BLN(BLN61),.WL(WL139));
sram_cell_6t_5 inst_cell_139_62 (.BL(BL62),.BLN(BLN62),.WL(WL139));
sram_cell_6t_5 inst_cell_139_63 (.BL(BL63),.BLN(BLN63),.WL(WL139));
sram_cell_6t_5 inst_cell_139_64 (.BL(BL64),.BLN(BLN64),.WL(WL139));
sram_cell_6t_5 inst_cell_139_65 (.BL(BL65),.BLN(BLN65),.WL(WL139));
sram_cell_6t_5 inst_cell_139_66 (.BL(BL66),.BLN(BLN66),.WL(WL139));
sram_cell_6t_5 inst_cell_139_67 (.BL(BL67),.BLN(BLN67),.WL(WL139));
sram_cell_6t_5 inst_cell_139_68 (.BL(BL68),.BLN(BLN68),.WL(WL139));
sram_cell_6t_5 inst_cell_139_69 (.BL(BL69),.BLN(BLN69),.WL(WL139));
sram_cell_6t_5 inst_cell_139_70 (.BL(BL70),.BLN(BLN70),.WL(WL139));
sram_cell_6t_5 inst_cell_139_71 (.BL(BL71),.BLN(BLN71),.WL(WL139));
sram_cell_6t_5 inst_cell_139_72 (.BL(BL72),.BLN(BLN72),.WL(WL139));
sram_cell_6t_5 inst_cell_139_73 (.BL(BL73),.BLN(BLN73),.WL(WL139));
sram_cell_6t_5 inst_cell_139_74 (.BL(BL74),.BLN(BLN74),.WL(WL139));
sram_cell_6t_5 inst_cell_139_75 (.BL(BL75),.BLN(BLN75),.WL(WL139));
sram_cell_6t_5 inst_cell_139_76 (.BL(BL76),.BLN(BLN76),.WL(WL139));
sram_cell_6t_5 inst_cell_139_77 (.BL(BL77),.BLN(BLN77),.WL(WL139));
sram_cell_6t_5 inst_cell_139_78 (.BL(BL78),.BLN(BLN78),.WL(WL139));
sram_cell_6t_5 inst_cell_139_79 (.BL(BL79),.BLN(BLN79),.WL(WL139));
sram_cell_6t_5 inst_cell_139_80 (.BL(BL80),.BLN(BLN80),.WL(WL139));
sram_cell_6t_5 inst_cell_139_81 (.BL(BL81),.BLN(BLN81),.WL(WL139));
sram_cell_6t_5 inst_cell_139_82 (.BL(BL82),.BLN(BLN82),.WL(WL139));
sram_cell_6t_5 inst_cell_139_83 (.BL(BL83),.BLN(BLN83),.WL(WL139));
sram_cell_6t_5 inst_cell_139_84 (.BL(BL84),.BLN(BLN84),.WL(WL139));
sram_cell_6t_5 inst_cell_139_85 (.BL(BL85),.BLN(BLN85),.WL(WL139));
sram_cell_6t_5 inst_cell_139_86 (.BL(BL86),.BLN(BLN86),.WL(WL139));
sram_cell_6t_5 inst_cell_139_87 (.BL(BL87),.BLN(BLN87),.WL(WL139));
sram_cell_6t_5 inst_cell_139_88 (.BL(BL88),.BLN(BLN88),.WL(WL139));
sram_cell_6t_5 inst_cell_139_89 (.BL(BL89),.BLN(BLN89),.WL(WL139));
sram_cell_6t_5 inst_cell_139_90 (.BL(BL90),.BLN(BLN90),.WL(WL139));
sram_cell_6t_5 inst_cell_139_91 (.BL(BL91),.BLN(BLN91),.WL(WL139));
sram_cell_6t_5 inst_cell_139_92 (.BL(BL92),.BLN(BLN92),.WL(WL139));
sram_cell_6t_5 inst_cell_139_93 (.BL(BL93),.BLN(BLN93),.WL(WL139));
sram_cell_6t_5 inst_cell_139_94 (.BL(BL94),.BLN(BLN94),.WL(WL139));
sram_cell_6t_5 inst_cell_139_95 (.BL(BL95),.BLN(BLN95),.WL(WL139));
sram_cell_6t_5 inst_cell_139_96 (.BL(BL96),.BLN(BLN96),.WL(WL139));
sram_cell_6t_5 inst_cell_139_97 (.BL(BL97),.BLN(BLN97),.WL(WL139));
sram_cell_6t_5 inst_cell_139_98 (.BL(BL98),.BLN(BLN98),.WL(WL139));
sram_cell_6t_5 inst_cell_139_99 (.BL(BL99),.BLN(BLN99),.WL(WL139));
sram_cell_6t_5 inst_cell_139_100 (.BL(BL100),.BLN(BLN100),.WL(WL139));
sram_cell_6t_5 inst_cell_139_101 (.BL(BL101),.BLN(BLN101),.WL(WL139));
sram_cell_6t_5 inst_cell_139_102 (.BL(BL102),.BLN(BLN102),.WL(WL139));
sram_cell_6t_5 inst_cell_139_103 (.BL(BL103),.BLN(BLN103),.WL(WL139));
sram_cell_6t_5 inst_cell_139_104 (.BL(BL104),.BLN(BLN104),.WL(WL139));
sram_cell_6t_5 inst_cell_139_105 (.BL(BL105),.BLN(BLN105),.WL(WL139));
sram_cell_6t_5 inst_cell_139_106 (.BL(BL106),.BLN(BLN106),.WL(WL139));
sram_cell_6t_5 inst_cell_139_107 (.BL(BL107),.BLN(BLN107),.WL(WL139));
sram_cell_6t_5 inst_cell_139_108 (.BL(BL108),.BLN(BLN108),.WL(WL139));
sram_cell_6t_5 inst_cell_139_109 (.BL(BL109),.BLN(BLN109),.WL(WL139));
sram_cell_6t_5 inst_cell_139_110 (.BL(BL110),.BLN(BLN110),.WL(WL139));
sram_cell_6t_5 inst_cell_139_111 (.BL(BL111),.BLN(BLN111),.WL(WL139));
sram_cell_6t_5 inst_cell_139_112 (.BL(BL112),.BLN(BLN112),.WL(WL139));
sram_cell_6t_5 inst_cell_139_113 (.BL(BL113),.BLN(BLN113),.WL(WL139));
sram_cell_6t_5 inst_cell_139_114 (.BL(BL114),.BLN(BLN114),.WL(WL139));
sram_cell_6t_5 inst_cell_139_115 (.BL(BL115),.BLN(BLN115),.WL(WL139));
sram_cell_6t_5 inst_cell_139_116 (.BL(BL116),.BLN(BLN116),.WL(WL139));
sram_cell_6t_5 inst_cell_139_117 (.BL(BL117),.BLN(BLN117),.WL(WL139));
sram_cell_6t_5 inst_cell_139_118 (.BL(BL118),.BLN(BLN118),.WL(WL139));
sram_cell_6t_5 inst_cell_139_119 (.BL(BL119),.BLN(BLN119),.WL(WL139));
sram_cell_6t_5 inst_cell_139_120 (.BL(BL120),.BLN(BLN120),.WL(WL139));
sram_cell_6t_5 inst_cell_139_121 (.BL(BL121),.BLN(BLN121),.WL(WL139));
sram_cell_6t_5 inst_cell_139_122 (.BL(BL122),.BLN(BLN122),.WL(WL139));
sram_cell_6t_5 inst_cell_139_123 (.BL(BL123),.BLN(BLN123),.WL(WL139));
sram_cell_6t_5 inst_cell_139_124 (.BL(BL124),.BLN(BLN124),.WL(WL139));
sram_cell_6t_5 inst_cell_139_125 (.BL(BL125),.BLN(BLN125),.WL(WL139));
sram_cell_6t_5 inst_cell_139_126 (.BL(BL126),.BLN(BLN126),.WL(WL139));
sram_cell_6t_5 inst_cell_139_127 (.BL(BL127),.BLN(BLN127),.WL(WL139));
sram_cell_6t_5 inst_cell_140_0 (.BL(BL0),.BLN(BLN0),.WL(WL140));
sram_cell_6t_5 inst_cell_140_1 (.BL(BL1),.BLN(BLN1),.WL(WL140));
sram_cell_6t_5 inst_cell_140_2 (.BL(BL2),.BLN(BLN2),.WL(WL140));
sram_cell_6t_5 inst_cell_140_3 (.BL(BL3),.BLN(BLN3),.WL(WL140));
sram_cell_6t_5 inst_cell_140_4 (.BL(BL4),.BLN(BLN4),.WL(WL140));
sram_cell_6t_5 inst_cell_140_5 (.BL(BL5),.BLN(BLN5),.WL(WL140));
sram_cell_6t_5 inst_cell_140_6 (.BL(BL6),.BLN(BLN6),.WL(WL140));
sram_cell_6t_5 inst_cell_140_7 (.BL(BL7),.BLN(BLN7),.WL(WL140));
sram_cell_6t_5 inst_cell_140_8 (.BL(BL8),.BLN(BLN8),.WL(WL140));
sram_cell_6t_5 inst_cell_140_9 (.BL(BL9),.BLN(BLN9),.WL(WL140));
sram_cell_6t_5 inst_cell_140_10 (.BL(BL10),.BLN(BLN10),.WL(WL140));
sram_cell_6t_5 inst_cell_140_11 (.BL(BL11),.BLN(BLN11),.WL(WL140));
sram_cell_6t_5 inst_cell_140_12 (.BL(BL12),.BLN(BLN12),.WL(WL140));
sram_cell_6t_5 inst_cell_140_13 (.BL(BL13),.BLN(BLN13),.WL(WL140));
sram_cell_6t_5 inst_cell_140_14 (.BL(BL14),.BLN(BLN14),.WL(WL140));
sram_cell_6t_5 inst_cell_140_15 (.BL(BL15),.BLN(BLN15),.WL(WL140));
sram_cell_6t_5 inst_cell_140_16 (.BL(BL16),.BLN(BLN16),.WL(WL140));
sram_cell_6t_5 inst_cell_140_17 (.BL(BL17),.BLN(BLN17),.WL(WL140));
sram_cell_6t_5 inst_cell_140_18 (.BL(BL18),.BLN(BLN18),.WL(WL140));
sram_cell_6t_5 inst_cell_140_19 (.BL(BL19),.BLN(BLN19),.WL(WL140));
sram_cell_6t_5 inst_cell_140_20 (.BL(BL20),.BLN(BLN20),.WL(WL140));
sram_cell_6t_5 inst_cell_140_21 (.BL(BL21),.BLN(BLN21),.WL(WL140));
sram_cell_6t_5 inst_cell_140_22 (.BL(BL22),.BLN(BLN22),.WL(WL140));
sram_cell_6t_5 inst_cell_140_23 (.BL(BL23),.BLN(BLN23),.WL(WL140));
sram_cell_6t_5 inst_cell_140_24 (.BL(BL24),.BLN(BLN24),.WL(WL140));
sram_cell_6t_5 inst_cell_140_25 (.BL(BL25),.BLN(BLN25),.WL(WL140));
sram_cell_6t_5 inst_cell_140_26 (.BL(BL26),.BLN(BLN26),.WL(WL140));
sram_cell_6t_5 inst_cell_140_27 (.BL(BL27),.BLN(BLN27),.WL(WL140));
sram_cell_6t_5 inst_cell_140_28 (.BL(BL28),.BLN(BLN28),.WL(WL140));
sram_cell_6t_5 inst_cell_140_29 (.BL(BL29),.BLN(BLN29),.WL(WL140));
sram_cell_6t_5 inst_cell_140_30 (.BL(BL30),.BLN(BLN30),.WL(WL140));
sram_cell_6t_5 inst_cell_140_31 (.BL(BL31),.BLN(BLN31),.WL(WL140));
sram_cell_6t_5 inst_cell_140_32 (.BL(BL32),.BLN(BLN32),.WL(WL140));
sram_cell_6t_5 inst_cell_140_33 (.BL(BL33),.BLN(BLN33),.WL(WL140));
sram_cell_6t_5 inst_cell_140_34 (.BL(BL34),.BLN(BLN34),.WL(WL140));
sram_cell_6t_5 inst_cell_140_35 (.BL(BL35),.BLN(BLN35),.WL(WL140));
sram_cell_6t_5 inst_cell_140_36 (.BL(BL36),.BLN(BLN36),.WL(WL140));
sram_cell_6t_5 inst_cell_140_37 (.BL(BL37),.BLN(BLN37),.WL(WL140));
sram_cell_6t_5 inst_cell_140_38 (.BL(BL38),.BLN(BLN38),.WL(WL140));
sram_cell_6t_5 inst_cell_140_39 (.BL(BL39),.BLN(BLN39),.WL(WL140));
sram_cell_6t_5 inst_cell_140_40 (.BL(BL40),.BLN(BLN40),.WL(WL140));
sram_cell_6t_5 inst_cell_140_41 (.BL(BL41),.BLN(BLN41),.WL(WL140));
sram_cell_6t_5 inst_cell_140_42 (.BL(BL42),.BLN(BLN42),.WL(WL140));
sram_cell_6t_5 inst_cell_140_43 (.BL(BL43),.BLN(BLN43),.WL(WL140));
sram_cell_6t_5 inst_cell_140_44 (.BL(BL44),.BLN(BLN44),.WL(WL140));
sram_cell_6t_5 inst_cell_140_45 (.BL(BL45),.BLN(BLN45),.WL(WL140));
sram_cell_6t_5 inst_cell_140_46 (.BL(BL46),.BLN(BLN46),.WL(WL140));
sram_cell_6t_5 inst_cell_140_47 (.BL(BL47),.BLN(BLN47),.WL(WL140));
sram_cell_6t_5 inst_cell_140_48 (.BL(BL48),.BLN(BLN48),.WL(WL140));
sram_cell_6t_5 inst_cell_140_49 (.BL(BL49),.BLN(BLN49),.WL(WL140));
sram_cell_6t_5 inst_cell_140_50 (.BL(BL50),.BLN(BLN50),.WL(WL140));
sram_cell_6t_5 inst_cell_140_51 (.BL(BL51),.BLN(BLN51),.WL(WL140));
sram_cell_6t_5 inst_cell_140_52 (.BL(BL52),.BLN(BLN52),.WL(WL140));
sram_cell_6t_5 inst_cell_140_53 (.BL(BL53),.BLN(BLN53),.WL(WL140));
sram_cell_6t_5 inst_cell_140_54 (.BL(BL54),.BLN(BLN54),.WL(WL140));
sram_cell_6t_5 inst_cell_140_55 (.BL(BL55),.BLN(BLN55),.WL(WL140));
sram_cell_6t_5 inst_cell_140_56 (.BL(BL56),.BLN(BLN56),.WL(WL140));
sram_cell_6t_5 inst_cell_140_57 (.BL(BL57),.BLN(BLN57),.WL(WL140));
sram_cell_6t_5 inst_cell_140_58 (.BL(BL58),.BLN(BLN58),.WL(WL140));
sram_cell_6t_5 inst_cell_140_59 (.BL(BL59),.BLN(BLN59),.WL(WL140));
sram_cell_6t_5 inst_cell_140_60 (.BL(BL60),.BLN(BLN60),.WL(WL140));
sram_cell_6t_5 inst_cell_140_61 (.BL(BL61),.BLN(BLN61),.WL(WL140));
sram_cell_6t_5 inst_cell_140_62 (.BL(BL62),.BLN(BLN62),.WL(WL140));
sram_cell_6t_5 inst_cell_140_63 (.BL(BL63),.BLN(BLN63),.WL(WL140));
sram_cell_6t_5 inst_cell_140_64 (.BL(BL64),.BLN(BLN64),.WL(WL140));
sram_cell_6t_5 inst_cell_140_65 (.BL(BL65),.BLN(BLN65),.WL(WL140));
sram_cell_6t_5 inst_cell_140_66 (.BL(BL66),.BLN(BLN66),.WL(WL140));
sram_cell_6t_5 inst_cell_140_67 (.BL(BL67),.BLN(BLN67),.WL(WL140));
sram_cell_6t_5 inst_cell_140_68 (.BL(BL68),.BLN(BLN68),.WL(WL140));
sram_cell_6t_5 inst_cell_140_69 (.BL(BL69),.BLN(BLN69),.WL(WL140));
sram_cell_6t_5 inst_cell_140_70 (.BL(BL70),.BLN(BLN70),.WL(WL140));
sram_cell_6t_5 inst_cell_140_71 (.BL(BL71),.BLN(BLN71),.WL(WL140));
sram_cell_6t_5 inst_cell_140_72 (.BL(BL72),.BLN(BLN72),.WL(WL140));
sram_cell_6t_5 inst_cell_140_73 (.BL(BL73),.BLN(BLN73),.WL(WL140));
sram_cell_6t_5 inst_cell_140_74 (.BL(BL74),.BLN(BLN74),.WL(WL140));
sram_cell_6t_5 inst_cell_140_75 (.BL(BL75),.BLN(BLN75),.WL(WL140));
sram_cell_6t_5 inst_cell_140_76 (.BL(BL76),.BLN(BLN76),.WL(WL140));
sram_cell_6t_5 inst_cell_140_77 (.BL(BL77),.BLN(BLN77),.WL(WL140));
sram_cell_6t_5 inst_cell_140_78 (.BL(BL78),.BLN(BLN78),.WL(WL140));
sram_cell_6t_5 inst_cell_140_79 (.BL(BL79),.BLN(BLN79),.WL(WL140));
sram_cell_6t_5 inst_cell_140_80 (.BL(BL80),.BLN(BLN80),.WL(WL140));
sram_cell_6t_5 inst_cell_140_81 (.BL(BL81),.BLN(BLN81),.WL(WL140));
sram_cell_6t_5 inst_cell_140_82 (.BL(BL82),.BLN(BLN82),.WL(WL140));
sram_cell_6t_5 inst_cell_140_83 (.BL(BL83),.BLN(BLN83),.WL(WL140));
sram_cell_6t_5 inst_cell_140_84 (.BL(BL84),.BLN(BLN84),.WL(WL140));
sram_cell_6t_5 inst_cell_140_85 (.BL(BL85),.BLN(BLN85),.WL(WL140));
sram_cell_6t_5 inst_cell_140_86 (.BL(BL86),.BLN(BLN86),.WL(WL140));
sram_cell_6t_5 inst_cell_140_87 (.BL(BL87),.BLN(BLN87),.WL(WL140));
sram_cell_6t_5 inst_cell_140_88 (.BL(BL88),.BLN(BLN88),.WL(WL140));
sram_cell_6t_5 inst_cell_140_89 (.BL(BL89),.BLN(BLN89),.WL(WL140));
sram_cell_6t_5 inst_cell_140_90 (.BL(BL90),.BLN(BLN90),.WL(WL140));
sram_cell_6t_5 inst_cell_140_91 (.BL(BL91),.BLN(BLN91),.WL(WL140));
sram_cell_6t_5 inst_cell_140_92 (.BL(BL92),.BLN(BLN92),.WL(WL140));
sram_cell_6t_5 inst_cell_140_93 (.BL(BL93),.BLN(BLN93),.WL(WL140));
sram_cell_6t_5 inst_cell_140_94 (.BL(BL94),.BLN(BLN94),.WL(WL140));
sram_cell_6t_5 inst_cell_140_95 (.BL(BL95),.BLN(BLN95),.WL(WL140));
sram_cell_6t_5 inst_cell_140_96 (.BL(BL96),.BLN(BLN96),.WL(WL140));
sram_cell_6t_5 inst_cell_140_97 (.BL(BL97),.BLN(BLN97),.WL(WL140));
sram_cell_6t_5 inst_cell_140_98 (.BL(BL98),.BLN(BLN98),.WL(WL140));
sram_cell_6t_5 inst_cell_140_99 (.BL(BL99),.BLN(BLN99),.WL(WL140));
sram_cell_6t_5 inst_cell_140_100 (.BL(BL100),.BLN(BLN100),.WL(WL140));
sram_cell_6t_5 inst_cell_140_101 (.BL(BL101),.BLN(BLN101),.WL(WL140));
sram_cell_6t_5 inst_cell_140_102 (.BL(BL102),.BLN(BLN102),.WL(WL140));
sram_cell_6t_5 inst_cell_140_103 (.BL(BL103),.BLN(BLN103),.WL(WL140));
sram_cell_6t_5 inst_cell_140_104 (.BL(BL104),.BLN(BLN104),.WL(WL140));
sram_cell_6t_5 inst_cell_140_105 (.BL(BL105),.BLN(BLN105),.WL(WL140));
sram_cell_6t_5 inst_cell_140_106 (.BL(BL106),.BLN(BLN106),.WL(WL140));
sram_cell_6t_5 inst_cell_140_107 (.BL(BL107),.BLN(BLN107),.WL(WL140));
sram_cell_6t_5 inst_cell_140_108 (.BL(BL108),.BLN(BLN108),.WL(WL140));
sram_cell_6t_5 inst_cell_140_109 (.BL(BL109),.BLN(BLN109),.WL(WL140));
sram_cell_6t_5 inst_cell_140_110 (.BL(BL110),.BLN(BLN110),.WL(WL140));
sram_cell_6t_5 inst_cell_140_111 (.BL(BL111),.BLN(BLN111),.WL(WL140));
sram_cell_6t_5 inst_cell_140_112 (.BL(BL112),.BLN(BLN112),.WL(WL140));
sram_cell_6t_5 inst_cell_140_113 (.BL(BL113),.BLN(BLN113),.WL(WL140));
sram_cell_6t_5 inst_cell_140_114 (.BL(BL114),.BLN(BLN114),.WL(WL140));
sram_cell_6t_5 inst_cell_140_115 (.BL(BL115),.BLN(BLN115),.WL(WL140));
sram_cell_6t_5 inst_cell_140_116 (.BL(BL116),.BLN(BLN116),.WL(WL140));
sram_cell_6t_5 inst_cell_140_117 (.BL(BL117),.BLN(BLN117),.WL(WL140));
sram_cell_6t_5 inst_cell_140_118 (.BL(BL118),.BLN(BLN118),.WL(WL140));
sram_cell_6t_5 inst_cell_140_119 (.BL(BL119),.BLN(BLN119),.WL(WL140));
sram_cell_6t_5 inst_cell_140_120 (.BL(BL120),.BLN(BLN120),.WL(WL140));
sram_cell_6t_5 inst_cell_140_121 (.BL(BL121),.BLN(BLN121),.WL(WL140));
sram_cell_6t_5 inst_cell_140_122 (.BL(BL122),.BLN(BLN122),.WL(WL140));
sram_cell_6t_5 inst_cell_140_123 (.BL(BL123),.BLN(BLN123),.WL(WL140));
sram_cell_6t_5 inst_cell_140_124 (.BL(BL124),.BLN(BLN124),.WL(WL140));
sram_cell_6t_5 inst_cell_140_125 (.BL(BL125),.BLN(BLN125),.WL(WL140));
sram_cell_6t_5 inst_cell_140_126 (.BL(BL126),.BLN(BLN126),.WL(WL140));
sram_cell_6t_5 inst_cell_140_127 (.BL(BL127),.BLN(BLN127),.WL(WL140));
sram_cell_6t_5 inst_cell_141_0 (.BL(BL0),.BLN(BLN0),.WL(WL141));
sram_cell_6t_5 inst_cell_141_1 (.BL(BL1),.BLN(BLN1),.WL(WL141));
sram_cell_6t_5 inst_cell_141_2 (.BL(BL2),.BLN(BLN2),.WL(WL141));
sram_cell_6t_5 inst_cell_141_3 (.BL(BL3),.BLN(BLN3),.WL(WL141));
sram_cell_6t_5 inst_cell_141_4 (.BL(BL4),.BLN(BLN4),.WL(WL141));
sram_cell_6t_5 inst_cell_141_5 (.BL(BL5),.BLN(BLN5),.WL(WL141));
sram_cell_6t_5 inst_cell_141_6 (.BL(BL6),.BLN(BLN6),.WL(WL141));
sram_cell_6t_5 inst_cell_141_7 (.BL(BL7),.BLN(BLN7),.WL(WL141));
sram_cell_6t_5 inst_cell_141_8 (.BL(BL8),.BLN(BLN8),.WL(WL141));
sram_cell_6t_5 inst_cell_141_9 (.BL(BL9),.BLN(BLN9),.WL(WL141));
sram_cell_6t_5 inst_cell_141_10 (.BL(BL10),.BLN(BLN10),.WL(WL141));
sram_cell_6t_5 inst_cell_141_11 (.BL(BL11),.BLN(BLN11),.WL(WL141));
sram_cell_6t_5 inst_cell_141_12 (.BL(BL12),.BLN(BLN12),.WL(WL141));
sram_cell_6t_5 inst_cell_141_13 (.BL(BL13),.BLN(BLN13),.WL(WL141));
sram_cell_6t_5 inst_cell_141_14 (.BL(BL14),.BLN(BLN14),.WL(WL141));
sram_cell_6t_5 inst_cell_141_15 (.BL(BL15),.BLN(BLN15),.WL(WL141));
sram_cell_6t_5 inst_cell_141_16 (.BL(BL16),.BLN(BLN16),.WL(WL141));
sram_cell_6t_5 inst_cell_141_17 (.BL(BL17),.BLN(BLN17),.WL(WL141));
sram_cell_6t_5 inst_cell_141_18 (.BL(BL18),.BLN(BLN18),.WL(WL141));
sram_cell_6t_5 inst_cell_141_19 (.BL(BL19),.BLN(BLN19),.WL(WL141));
sram_cell_6t_5 inst_cell_141_20 (.BL(BL20),.BLN(BLN20),.WL(WL141));
sram_cell_6t_5 inst_cell_141_21 (.BL(BL21),.BLN(BLN21),.WL(WL141));
sram_cell_6t_5 inst_cell_141_22 (.BL(BL22),.BLN(BLN22),.WL(WL141));
sram_cell_6t_5 inst_cell_141_23 (.BL(BL23),.BLN(BLN23),.WL(WL141));
sram_cell_6t_5 inst_cell_141_24 (.BL(BL24),.BLN(BLN24),.WL(WL141));
sram_cell_6t_5 inst_cell_141_25 (.BL(BL25),.BLN(BLN25),.WL(WL141));
sram_cell_6t_5 inst_cell_141_26 (.BL(BL26),.BLN(BLN26),.WL(WL141));
sram_cell_6t_5 inst_cell_141_27 (.BL(BL27),.BLN(BLN27),.WL(WL141));
sram_cell_6t_5 inst_cell_141_28 (.BL(BL28),.BLN(BLN28),.WL(WL141));
sram_cell_6t_5 inst_cell_141_29 (.BL(BL29),.BLN(BLN29),.WL(WL141));
sram_cell_6t_5 inst_cell_141_30 (.BL(BL30),.BLN(BLN30),.WL(WL141));
sram_cell_6t_5 inst_cell_141_31 (.BL(BL31),.BLN(BLN31),.WL(WL141));
sram_cell_6t_5 inst_cell_141_32 (.BL(BL32),.BLN(BLN32),.WL(WL141));
sram_cell_6t_5 inst_cell_141_33 (.BL(BL33),.BLN(BLN33),.WL(WL141));
sram_cell_6t_5 inst_cell_141_34 (.BL(BL34),.BLN(BLN34),.WL(WL141));
sram_cell_6t_5 inst_cell_141_35 (.BL(BL35),.BLN(BLN35),.WL(WL141));
sram_cell_6t_5 inst_cell_141_36 (.BL(BL36),.BLN(BLN36),.WL(WL141));
sram_cell_6t_5 inst_cell_141_37 (.BL(BL37),.BLN(BLN37),.WL(WL141));
sram_cell_6t_5 inst_cell_141_38 (.BL(BL38),.BLN(BLN38),.WL(WL141));
sram_cell_6t_5 inst_cell_141_39 (.BL(BL39),.BLN(BLN39),.WL(WL141));
sram_cell_6t_5 inst_cell_141_40 (.BL(BL40),.BLN(BLN40),.WL(WL141));
sram_cell_6t_5 inst_cell_141_41 (.BL(BL41),.BLN(BLN41),.WL(WL141));
sram_cell_6t_5 inst_cell_141_42 (.BL(BL42),.BLN(BLN42),.WL(WL141));
sram_cell_6t_5 inst_cell_141_43 (.BL(BL43),.BLN(BLN43),.WL(WL141));
sram_cell_6t_5 inst_cell_141_44 (.BL(BL44),.BLN(BLN44),.WL(WL141));
sram_cell_6t_5 inst_cell_141_45 (.BL(BL45),.BLN(BLN45),.WL(WL141));
sram_cell_6t_5 inst_cell_141_46 (.BL(BL46),.BLN(BLN46),.WL(WL141));
sram_cell_6t_5 inst_cell_141_47 (.BL(BL47),.BLN(BLN47),.WL(WL141));
sram_cell_6t_5 inst_cell_141_48 (.BL(BL48),.BLN(BLN48),.WL(WL141));
sram_cell_6t_5 inst_cell_141_49 (.BL(BL49),.BLN(BLN49),.WL(WL141));
sram_cell_6t_5 inst_cell_141_50 (.BL(BL50),.BLN(BLN50),.WL(WL141));
sram_cell_6t_5 inst_cell_141_51 (.BL(BL51),.BLN(BLN51),.WL(WL141));
sram_cell_6t_5 inst_cell_141_52 (.BL(BL52),.BLN(BLN52),.WL(WL141));
sram_cell_6t_5 inst_cell_141_53 (.BL(BL53),.BLN(BLN53),.WL(WL141));
sram_cell_6t_5 inst_cell_141_54 (.BL(BL54),.BLN(BLN54),.WL(WL141));
sram_cell_6t_5 inst_cell_141_55 (.BL(BL55),.BLN(BLN55),.WL(WL141));
sram_cell_6t_5 inst_cell_141_56 (.BL(BL56),.BLN(BLN56),.WL(WL141));
sram_cell_6t_5 inst_cell_141_57 (.BL(BL57),.BLN(BLN57),.WL(WL141));
sram_cell_6t_5 inst_cell_141_58 (.BL(BL58),.BLN(BLN58),.WL(WL141));
sram_cell_6t_5 inst_cell_141_59 (.BL(BL59),.BLN(BLN59),.WL(WL141));
sram_cell_6t_5 inst_cell_141_60 (.BL(BL60),.BLN(BLN60),.WL(WL141));
sram_cell_6t_5 inst_cell_141_61 (.BL(BL61),.BLN(BLN61),.WL(WL141));
sram_cell_6t_5 inst_cell_141_62 (.BL(BL62),.BLN(BLN62),.WL(WL141));
sram_cell_6t_5 inst_cell_141_63 (.BL(BL63),.BLN(BLN63),.WL(WL141));
sram_cell_6t_5 inst_cell_141_64 (.BL(BL64),.BLN(BLN64),.WL(WL141));
sram_cell_6t_5 inst_cell_141_65 (.BL(BL65),.BLN(BLN65),.WL(WL141));
sram_cell_6t_5 inst_cell_141_66 (.BL(BL66),.BLN(BLN66),.WL(WL141));
sram_cell_6t_5 inst_cell_141_67 (.BL(BL67),.BLN(BLN67),.WL(WL141));
sram_cell_6t_5 inst_cell_141_68 (.BL(BL68),.BLN(BLN68),.WL(WL141));
sram_cell_6t_5 inst_cell_141_69 (.BL(BL69),.BLN(BLN69),.WL(WL141));
sram_cell_6t_5 inst_cell_141_70 (.BL(BL70),.BLN(BLN70),.WL(WL141));
sram_cell_6t_5 inst_cell_141_71 (.BL(BL71),.BLN(BLN71),.WL(WL141));
sram_cell_6t_5 inst_cell_141_72 (.BL(BL72),.BLN(BLN72),.WL(WL141));
sram_cell_6t_5 inst_cell_141_73 (.BL(BL73),.BLN(BLN73),.WL(WL141));
sram_cell_6t_5 inst_cell_141_74 (.BL(BL74),.BLN(BLN74),.WL(WL141));
sram_cell_6t_5 inst_cell_141_75 (.BL(BL75),.BLN(BLN75),.WL(WL141));
sram_cell_6t_5 inst_cell_141_76 (.BL(BL76),.BLN(BLN76),.WL(WL141));
sram_cell_6t_5 inst_cell_141_77 (.BL(BL77),.BLN(BLN77),.WL(WL141));
sram_cell_6t_5 inst_cell_141_78 (.BL(BL78),.BLN(BLN78),.WL(WL141));
sram_cell_6t_5 inst_cell_141_79 (.BL(BL79),.BLN(BLN79),.WL(WL141));
sram_cell_6t_5 inst_cell_141_80 (.BL(BL80),.BLN(BLN80),.WL(WL141));
sram_cell_6t_5 inst_cell_141_81 (.BL(BL81),.BLN(BLN81),.WL(WL141));
sram_cell_6t_5 inst_cell_141_82 (.BL(BL82),.BLN(BLN82),.WL(WL141));
sram_cell_6t_5 inst_cell_141_83 (.BL(BL83),.BLN(BLN83),.WL(WL141));
sram_cell_6t_5 inst_cell_141_84 (.BL(BL84),.BLN(BLN84),.WL(WL141));
sram_cell_6t_5 inst_cell_141_85 (.BL(BL85),.BLN(BLN85),.WL(WL141));
sram_cell_6t_5 inst_cell_141_86 (.BL(BL86),.BLN(BLN86),.WL(WL141));
sram_cell_6t_5 inst_cell_141_87 (.BL(BL87),.BLN(BLN87),.WL(WL141));
sram_cell_6t_5 inst_cell_141_88 (.BL(BL88),.BLN(BLN88),.WL(WL141));
sram_cell_6t_5 inst_cell_141_89 (.BL(BL89),.BLN(BLN89),.WL(WL141));
sram_cell_6t_5 inst_cell_141_90 (.BL(BL90),.BLN(BLN90),.WL(WL141));
sram_cell_6t_5 inst_cell_141_91 (.BL(BL91),.BLN(BLN91),.WL(WL141));
sram_cell_6t_5 inst_cell_141_92 (.BL(BL92),.BLN(BLN92),.WL(WL141));
sram_cell_6t_5 inst_cell_141_93 (.BL(BL93),.BLN(BLN93),.WL(WL141));
sram_cell_6t_5 inst_cell_141_94 (.BL(BL94),.BLN(BLN94),.WL(WL141));
sram_cell_6t_5 inst_cell_141_95 (.BL(BL95),.BLN(BLN95),.WL(WL141));
sram_cell_6t_5 inst_cell_141_96 (.BL(BL96),.BLN(BLN96),.WL(WL141));
sram_cell_6t_5 inst_cell_141_97 (.BL(BL97),.BLN(BLN97),.WL(WL141));
sram_cell_6t_5 inst_cell_141_98 (.BL(BL98),.BLN(BLN98),.WL(WL141));
sram_cell_6t_5 inst_cell_141_99 (.BL(BL99),.BLN(BLN99),.WL(WL141));
sram_cell_6t_5 inst_cell_141_100 (.BL(BL100),.BLN(BLN100),.WL(WL141));
sram_cell_6t_5 inst_cell_141_101 (.BL(BL101),.BLN(BLN101),.WL(WL141));
sram_cell_6t_5 inst_cell_141_102 (.BL(BL102),.BLN(BLN102),.WL(WL141));
sram_cell_6t_5 inst_cell_141_103 (.BL(BL103),.BLN(BLN103),.WL(WL141));
sram_cell_6t_5 inst_cell_141_104 (.BL(BL104),.BLN(BLN104),.WL(WL141));
sram_cell_6t_5 inst_cell_141_105 (.BL(BL105),.BLN(BLN105),.WL(WL141));
sram_cell_6t_5 inst_cell_141_106 (.BL(BL106),.BLN(BLN106),.WL(WL141));
sram_cell_6t_5 inst_cell_141_107 (.BL(BL107),.BLN(BLN107),.WL(WL141));
sram_cell_6t_5 inst_cell_141_108 (.BL(BL108),.BLN(BLN108),.WL(WL141));
sram_cell_6t_5 inst_cell_141_109 (.BL(BL109),.BLN(BLN109),.WL(WL141));
sram_cell_6t_5 inst_cell_141_110 (.BL(BL110),.BLN(BLN110),.WL(WL141));
sram_cell_6t_5 inst_cell_141_111 (.BL(BL111),.BLN(BLN111),.WL(WL141));
sram_cell_6t_5 inst_cell_141_112 (.BL(BL112),.BLN(BLN112),.WL(WL141));
sram_cell_6t_5 inst_cell_141_113 (.BL(BL113),.BLN(BLN113),.WL(WL141));
sram_cell_6t_5 inst_cell_141_114 (.BL(BL114),.BLN(BLN114),.WL(WL141));
sram_cell_6t_5 inst_cell_141_115 (.BL(BL115),.BLN(BLN115),.WL(WL141));
sram_cell_6t_5 inst_cell_141_116 (.BL(BL116),.BLN(BLN116),.WL(WL141));
sram_cell_6t_5 inst_cell_141_117 (.BL(BL117),.BLN(BLN117),.WL(WL141));
sram_cell_6t_5 inst_cell_141_118 (.BL(BL118),.BLN(BLN118),.WL(WL141));
sram_cell_6t_5 inst_cell_141_119 (.BL(BL119),.BLN(BLN119),.WL(WL141));
sram_cell_6t_5 inst_cell_141_120 (.BL(BL120),.BLN(BLN120),.WL(WL141));
sram_cell_6t_5 inst_cell_141_121 (.BL(BL121),.BLN(BLN121),.WL(WL141));
sram_cell_6t_5 inst_cell_141_122 (.BL(BL122),.BLN(BLN122),.WL(WL141));
sram_cell_6t_5 inst_cell_141_123 (.BL(BL123),.BLN(BLN123),.WL(WL141));
sram_cell_6t_5 inst_cell_141_124 (.BL(BL124),.BLN(BLN124),.WL(WL141));
sram_cell_6t_5 inst_cell_141_125 (.BL(BL125),.BLN(BLN125),.WL(WL141));
sram_cell_6t_5 inst_cell_141_126 (.BL(BL126),.BLN(BLN126),.WL(WL141));
sram_cell_6t_5 inst_cell_141_127 (.BL(BL127),.BLN(BLN127),.WL(WL141));
sram_cell_6t_5 inst_cell_142_0 (.BL(BL0),.BLN(BLN0),.WL(WL142));
sram_cell_6t_5 inst_cell_142_1 (.BL(BL1),.BLN(BLN1),.WL(WL142));
sram_cell_6t_5 inst_cell_142_2 (.BL(BL2),.BLN(BLN2),.WL(WL142));
sram_cell_6t_5 inst_cell_142_3 (.BL(BL3),.BLN(BLN3),.WL(WL142));
sram_cell_6t_5 inst_cell_142_4 (.BL(BL4),.BLN(BLN4),.WL(WL142));
sram_cell_6t_5 inst_cell_142_5 (.BL(BL5),.BLN(BLN5),.WL(WL142));
sram_cell_6t_5 inst_cell_142_6 (.BL(BL6),.BLN(BLN6),.WL(WL142));
sram_cell_6t_5 inst_cell_142_7 (.BL(BL7),.BLN(BLN7),.WL(WL142));
sram_cell_6t_5 inst_cell_142_8 (.BL(BL8),.BLN(BLN8),.WL(WL142));
sram_cell_6t_5 inst_cell_142_9 (.BL(BL9),.BLN(BLN9),.WL(WL142));
sram_cell_6t_5 inst_cell_142_10 (.BL(BL10),.BLN(BLN10),.WL(WL142));
sram_cell_6t_5 inst_cell_142_11 (.BL(BL11),.BLN(BLN11),.WL(WL142));
sram_cell_6t_5 inst_cell_142_12 (.BL(BL12),.BLN(BLN12),.WL(WL142));
sram_cell_6t_5 inst_cell_142_13 (.BL(BL13),.BLN(BLN13),.WL(WL142));
sram_cell_6t_5 inst_cell_142_14 (.BL(BL14),.BLN(BLN14),.WL(WL142));
sram_cell_6t_5 inst_cell_142_15 (.BL(BL15),.BLN(BLN15),.WL(WL142));
sram_cell_6t_5 inst_cell_142_16 (.BL(BL16),.BLN(BLN16),.WL(WL142));
sram_cell_6t_5 inst_cell_142_17 (.BL(BL17),.BLN(BLN17),.WL(WL142));
sram_cell_6t_5 inst_cell_142_18 (.BL(BL18),.BLN(BLN18),.WL(WL142));
sram_cell_6t_5 inst_cell_142_19 (.BL(BL19),.BLN(BLN19),.WL(WL142));
sram_cell_6t_5 inst_cell_142_20 (.BL(BL20),.BLN(BLN20),.WL(WL142));
sram_cell_6t_5 inst_cell_142_21 (.BL(BL21),.BLN(BLN21),.WL(WL142));
sram_cell_6t_5 inst_cell_142_22 (.BL(BL22),.BLN(BLN22),.WL(WL142));
sram_cell_6t_5 inst_cell_142_23 (.BL(BL23),.BLN(BLN23),.WL(WL142));
sram_cell_6t_5 inst_cell_142_24 (.BL(BL24),.BLN(BLN24),.WL(WL142));
sram_cell_6t_5 inst_cell_142_25 (.BL(BL25),.BLN(BLN25),.WL(WL142));
sram_cell_6t_5 inst_cell_142_26 (.BL(BL26),.BLN(BLN26),.WL(WL142));
sram_cell_6t_5 inst_cell_142_27 (.BL(BL27),.BLN(BLN27),.WL(WL142));
sram_cell_6t_5 inst_cell_142_28 (.BL(BL28),.BLN(BLN28),.WL(WL142));
sram_cell_6t_5 inst_cell_142_29 (.BL(BL29),.BLN(BLN29),.WL(WL142));
sram_cell_6t_5 inst_cell_142_30 (.BL(BL30),.BLN(BLN30),.WL(WL142));
sram_cell_6t_5 inst_cell_142_31 (.BL(BL31),.BLN(BLN31),.WL(WL142));
sram_cell_6t_5 inst_cell_142_32 (.BL(BL32),.BLN(BLN32),.WL(WL142));
sram_cell_6t_5 inst_cell_142_33 (.BL(BL33),.BLN(BLN33),.WL(WL142));
sram_cell_6t_5 inst_cell_142_34 (.BL(BL34),.BLN(BLN34),.WL(WL142));
sram_cell_6t_5 inst_cell_142_35 (.BL(BL35),.BLN(BLN35),.WL(WL142));
sram_cell_6t_5 inst_cell_142_36 (.BL(BL36),.BLN(BLN36),.WL(WL142));
sram_cell_6t_5 inst_cell_142_37 (.BL(BL37),.BLN(BLN37),.WL(WL142));
sram_cell_6t_5 inst_cell_142_38 (.BL(BL38),.BLN(BLN38),.WL(WL142));
sram_cell_6t_5 inst_cell_142_39 (.BL(BL39),.BLN(BLN39),.WL(WL142));
sram_cell_6t_5 inst_cell_142_40 (.BL(BL40),.BLN(BLN40),.WL(WL142));
sram_cell_6t_5 inst_cell_142_41 (.BL(BL41),.BLN(BLN41),.WL(WL142));
sram_cell_6t_5 inst_cell_142_42 (.BL(BL42),.BLN(BLN42),.WL(WL142));
sram_cell_6t_5 inst_cell_142_43 (.BL(BL43),.BLN(BLN43),.WL(WL142));
sram_cell_6t_5 inst_cell_142_44 (.BL(BL44),.BLN(BLN44),.WL(WL142));
sram_cell_6t_5 inst_cell_142_45 (.BL(BL45),.BLN(BLN45),.WL(WL142));
sram_cell_6t_5 inst_cell_142_46 (.BL(BL46),.BLN(BLN46),.WL(WL142));
sram_cell_6t_5 inst_cell_142_47 (.BL(BL47),.BLN(BLN47),.WL(WL142));
sram_cell_6t_5 inst_cell_142_48 (.BL(BL48),.BLN(BLN48),.WL(WL142));
sram_cell_6t_5 inst_cell_142_49 (.BL(BL49),.BLN(BLN49),.WL(WL142));
sram_cell_6t_5 inst_cell_142_50 (.BL(BL50),.BLN(BLN50),.WL(WL142));
sram_cell_6t_5 inst_cell_142_51 (.BL(BL51),.BLN(BLN51),.WL(WL142));
sram_cell_6t_5 inst_cell_142_52 (.BL(BL52),.BLN(BLN52),.WL(WL142));
sram_cell_6t_5 inst_cell_142_53 (.BL(BL53),.BLN(BLN53),.WL(WL142));
sram_cell_6t_5 inst_cell_142_54 (.BL(BL54),.BLN(BLN54),.WL(WL142));
sram_cell_6t_5 inst_cell_142_55 (.BL(BL55),.BLN(BLN55),.WL(WL142));
sram_cell_6t_5 inst_cell_142_56 (.BL(BL56),.BLN(BLN56),.WL(WL142));
sram_cell_6t_5 inst_cell_142_57 (.BL(BL57),.BLN(BLN57),.WL(WL142));
sram_cell_6t_5 inst_cell_142_58 (.BL(BL58),.BLN(BLN58),.WL(WL142));
sram_cell_6t_5 inst_cell_142_59 (.BL(BL59),.BLN(BLN59),.WL(WL142));
sram_cell_6t_5 inst_cell_142_60 (.BL(BL60),.BLN(BLN60),.WL(WL142));
sram_cell_6t_5 inst_cell_142_61 (.BL(BL61),.BLN(BLN61),.WL(WL142));
sram_cell_6t_5 inst_cell_142_62 (.BL(BL62),.BLN(BLN62),.WL(WL142));
sram_cell_6t_5 inst_cell_142_63 (.BL(BL63),.BLN(BLN63),.WL(WL142));
sram_cell_6t_5 inst_cell_142_64 (.BL(BL64),.BLN(BLN64),.WL(WL142));
sram_cell_6t_5 inst_cell_142_65 (.BL(BL65),.BLN(BLN65),.WL(WL142));
sram_cell_6t_5 inst_cell_142_66 (.BL(BL66),.BLN(BLN66),.WL(WL142));
sram_cell_6t_5 inst_cell_142_67 (.BL(BL67),.BLN(BLN67),.WL(WL142));
sram_cell_6t_5 inst_cell_142_68 (.BL(BL68),.BLN(BLN68),.WL(WL142));
sram_cell_6t_5 inst_cell_142_69 (.BL(BL69),.BLN(BLN69),.WL(WL142));
sram_cell_6t_5 inst_cell_142_70 (.BL(BL70),.BLN(BLN70),.WL(WL142));
sram_cell_6t_5 inst_cell_142_71 (.BL(BL71),.BLN(BLN71),.WL(WL142));
sram_cell_6t_5 inst_cell_142_72 (.BL(BL72),.BLN(BLN72),.WL(WL142));
sram_cell_6t_5 inst_cell_142_73 (.BL(BL73),.BLN(BLN73),.WL(WL142));
sram_cell_6t_5 inst_cell_142_74 (.BL(BL74),.BLN(BLN74),.WL(WL142));
sram_cell_6t_5 inst_cell_142_75 (.BL(BL75),.BLN(BLN75),.WL(WL142));
sram_cell_6t_5 inst_cell_142_76 (.BL(BL76),.BLN(BLN76),.WL(WL142));
sram_cell_6t_5 inst_cell_142_77 (.BL(BL77),.BLN(BLN77),.WL(WL142));
sram_cell_6t_5 inst_cell_142_78 (.BL(BL78),.BLN(BLN78),.WL(WL142));
sram_cell_6t_5 inst_cell_142_79 (.BL(BL79),.BLN(BLN79),.WL(WL142));
sram_cell_6t_5 inst_cell_142_80 (.BL(BL80),.BLN(BLN80),.WL(WL142));
sram_cell_6t_5 inst_cell_142_81 (.BL(BL81),.BLN(BLN81),.WL(WL142));
sram_cell_6t_5 inst_cell_142_82 (.BL(BL82),.BLN(BLN82),.WL(WL142));
sram_cell_6t_5 inst_cell_142_83 (.BL(BL83),.BLN(BLN83),.WL(WL142));
sram_cell_6t_5 inst_cell_142_84 (.BL(BL84),.BLN(BLN84),.WL(WL142));
sram_cell_6t_5 inst_cell_142_85 (.BL(BL85),.BLN(BLN85),.WL(WL142));
sram_cell_6t_5 inst_cell_142_86 (.BL(BL86),.BLN(BLN86),.WL(WL142));
sram_cell_6t_5 inst_cell_142_87 (.BL(BL87),.BLN(BLN87),.WL(WL142));
sram_cell_6t_5 inst_cell_142_88 (.BL(BL88),.BLN(BLN88),.WL(WL142));
sram_cell_6t_5 inst_cell_142_89 (.BL(BL89),.BLN(BLN89),.WL(WL142));
sram_cell_6t_5 inst_cell_142_90 (.BL(BL90),.BLN(BLN90),.WL(WL142));
sram_cell_6t_5 inst_cell_142_91 (.BL(BL91),.BLN(BLN91),.WL(WL142));
sram_cell_6t_5 inst_cell_142_92 (.BL(BL92),.BLN(BLN92),.WL(WL142));
sram_cell_6t_5 inst_cell_142_93 (.BL(BL93),.BLN(BLN93),.WL(WL142));
sram_cell_6t_5 inst_cell_142_94 (.BL(BL94),.BLN(BLN94),.WL(WL142));
sram_cell_6t_5 inst_cell_142_95 (.BL(BL95),.BLN(BLN95),.WL(WL142));
sram_cell_6t_5 inst_cell_142_96 (.BL(BL96),.BLN(BLN96),.WL(WL142));
sram_cell_6t_5 inst_cell_142_97 (.BL(BL97),.BLN(BLN97),.WL(WL142));
sram_cell_6t_5 inst_cell_142_98 (.BL(BL98),.BLN(BLN98),.WL(WL142));
sram_cell_6t_5 inst_cell_142_99 (.BL(BL99),.BLN(BLN99),.WL(WL142));
sram_cell_6t_5 inst_cell_142_100 (.BL(BL100),.BLN(BLN100),.WL(WL142));
sram_cell_6t_5 inst_cell_142_101 (.BL(BL101),.BLN(BLN101),.WL(WL142));
sram_cell_6t_5 inst_cell_142_102 (.BL(BL102),.BLN(BLN102),.WL(WL142));
sram_cell_6t_5 inst_cell_142_103 (.BL(BL103),.BLN(BLN103),.WL(WL142));
sram_cell_6t_5 inst_cell_142_104 (.BL(BL104),.BLN(BLN104),.WL(WL142));
sram_cell_6t_5 inst_cell_142_105 (.BL(BL105),.BLN(BLN105),.WL(WL142));
sram_cell_6t_5 inst_cell_142_106 (.BL(BL106),.BLN(BLN106),.WL(WL142));
sram_cell_6t_5 inst_cell_142_107 (.BL(BL107),.BLN(BLN107),.WL(WL142));
sram_cell_6t_5 inst_cell_142_108 (.BL(BL108),.BLN(BLN108),.WL(WL142));
sram_cell_6t_5 inst_cell_142_109 (.BL(BL109),.BLN(BLN109),.WL(WL142));
sram_cell_6t_5 inst_cell_142_110 (.BL(BL110),.BLN(BLN110),.WL(WL142));
sram_cell_6t_5 inst_cell_142_111 (.BL(BL111),.BLN(BLN111),.WL(WL142));
sram_cell_6t_5 inst_cell_142_112 (.BL(BL112),.BLN(BLN112),.WL(WL142));
sram_cell_6t_5 inst_cell_142_113 (.BL(BL113),.BLN(BLN113),.WL(WL142));
sram_cell_6t_5 inst_cell_142_114 (.BL(BL114),.BLN(BLN114),.WL(WL142));
sram_cell_6t_5 inst_cell_142_115 (.BL(BL115),.BLN(BLN115),.WL(WL142));
sram_cell_6t_5 inst_cell_142_116 (.BL(BL116),.BLN(BLN116),.WL(WL142));
sram_cell_6t_5 inst_cell_142_117 (.BL(BL117),.BLN(BLN117),.WL(WL142));
sram_cell_6t_5 inst_cell_142_118 (.BL(BL118),.BLN(BLN118),.WL(WL142));
sram_cell_6t_5 inst_cell_142_119 (.BL(BL119),.BLN(BLN119),.WL(WL142));
sram_cell_6t_5 inst_cell_142_120 (.BL(BL120),.BLN(BLN120),.WL(WL142));
sram_cell_6t_5 inst_cell_142_121 (.BL(BL121),.BLN(BLN121),.WL(WL142));
sram_cell_6t_5 inst_cell_142_122 (.BL(BL122),.BLN(BLN122),.WL(WL142));
sram_cell_6t_5 inst_cell_142_123 (.BL(BL123),.BLN(BLN123),.WL(WL142));
sram_cell_6t_5 inst_cell_142_124 (.BL(BL124),.BLN(BLN124),.WL(WL142));
sram_cell_6t_5 inst_cell_142_125 (.BL(BL125),.BLN(BLN125),.WL(WL142));
sram_cell_6t_5 inst_cell_142_126 (.BL(BL126),.BLN(BLN126),.WL(WL142));
sram_cell_6t_5 inst_cell_142_127 (.BL(BL127),.BLN(BLN127),.WL(WL142));
sram_cell_6t_5 inst_cell_143_0 (.BL(BL0),.BLN(BLN0),.WL(WL143));
sram_cell_6t_5 inst_cell_143_1 (.BL(BL1),.BLN(BLN1),.WL(WL143));
sram_cell_6t_5 inst_cell_143_2 (.BL(BL2),.BLN(BLN2),.WL(WL143));
sram_cell_6t_5 inst_cell_143_3 (.BL(BL3),.BLN(BLN3),.WL(WL143));
sram_cell_6t_5 inst_cell_143_4 (.BL(BL4),.BLN(BLN4),.WL(WL143));
sram_cell_6t_5 inst_cell_143_5 (.BL(BL5),.BLN(BLN5),.WL(WL143));
sram_cell_6t_5 inst_cell_143_6 (.BL(BL6),.BLN(BLN6),.WL(WL143));
sram_cell_6t_5 inst_cell_143_7 (.BL(BL7),.BLN(BLN7),.WL(WL143));
sram_cell_6t_5 inst_cell_143_8 (.BL(BL8),.BLN(BLN8),.WL(WL143));
sram_cell_6t_5 inst_cell_143_9 (.BL(BL9),.BLN(BLN9),.WL(WL143));
sram_cell_6t_5 inst_cell_143_10 (.BL(BL10),.BLN(BLN10),.WL(WL143));
sram_cell_6t_5 inst_cell_143_11 (.BL(BL11),.BLN(BLN11),.WL(WL143));
sram_cell_6t_5 inst_cell_143_12 (.BL(BL12),.BLN(BLN12),.WL(WL143));
sram_cell_6t_5 inst_cell_143_13 (.BL(BL13),.BLN(BLN13),.WL(WL143));
sram_cell_6t_5 inst_cell_143_14 (.BL(BL14),.BLN(BLN14),.WL(WL143));
sram_cell_6t_5 inst_cell_143_15 (.BL(BL15),.BLN(BLN15),.WL(WL143));
sram_cell_6t_5 inst_cell_143_16 (.BL(BL16),.BLN(BLN16),.WL(WL143));
sram_cell_6t_5 inst_cell_143_17 (.BL(BL17),.BLN(BLN17),.WL(WL143));
sram_cell_6t_5 inst_cell_143_18 (.BL(BL18),.BLN(BLN18),.WL(WL143));
sram_cell_6t_5 inst_cell_143_19 (.BL(BL19),.BLN(BLN19),.WL(WL143));
sram_cell_6t_5 inst_cell_143_20 (.BL(BL20),.BLN(BLN20),.WL(WL143));
sram_cell_6t_5 inst_cell_143_21 (.BL(BL21),.BLN(BLN21),.WL(WL143));
sram_cell_6t_5 inst_cell_143_22 (.BL(BL22),.BLN(BLN22),.WL(WL143));
sram_cell_6t_5 inst_cell_143_23 (.BL(BL23),.BLN(BLN23),.WL(WL143));
sram_cell_6t_5 inst_cell_143_24 (.BL(BL24),.BLN(BLN24),.WL(WL143));
sram_cell_6t_5 inst_cell_143_25 (.BL(BL25),.BLN(BLN25),.WL(WL143));
sram_cell_6t_5 inst_cell_143_26 (.BL(BL26),.BLN(BLN26),.WL(WL143));
sram_cell_6t_5 inst_cell_143_27 (.BL(BL27),.BLN(BLN27),.WL(WL143));
sram_cell_6t_5 inst_cell_143_28 (.BL(BL28),.BLN(BLN28),.WL(WL143));
sram_cell_6t_5 inst_cell_143_29 (.BL(BL29),.BLN(BLN29),.WL(WL143));
sram_cell_6t_5 inst_cell_143_30 (.BL(BL30),.BLN(BLN30),.WL(WL143));
sram_cell_6t_5 inst_cell_143_31 (.BL(BL31),.BLN(BLN31),.WL(WL143));
sram_cell_6t_5 inst_cell_143_32 (.BL(BL32),.BLN(BLN32),.WL(WL143));
sram_cell_6t_5 inst_cell_143_33 (.BL(BL33),.BLN(BLN33),.WL(WL143));
sram_cell_6t_5 inst_cell_143_34 (.BL(BL34),.BLN(BLN34),.WL(WL143));
sram_cell_6t_5 inst_cell_143_35 (.BL(BL35),.BLN(BLN35),.WL(WL143));
sram_cell_6t_5 inst_cell_143_36 (.BL(BL36),.BLN(BLN36),.WL(WL143));
sram_cell_6t_5 inst_cell_143_37 (.BL(BL37),.BLN(BLN37),.WL(WL143));
sram_cell_6t_5 inst_cell_143_38 (.BL(BL38),.BLN(BLN38),.WL(WL143));
sram_cell_6t_5 inst_cell_143_39 (.BL(BL39),.BLN(BLN39),.WL(WL143));
sram_cell_6t_5 inst_cell_143_40 (.BL(BL40),.BLN(BLN40),.WL(WL143));
sram_cell_6t_5 inst_cell_143_41 (.BL(BL41),.BLN(BLN41),.WL(WL143));
sram_cell_6t_5 inst_cell_143_42 (.BL(BL42),.BLN(BLN42),.WL(WL143));
sram_cell_6t_5 inst_cell_143_43 (.BL(BL43),.BLN(BLN43),.WL(WL143));
sram_cell_6t_5 inst_cell_143_44 (.BL(BL44),.BLN(BLN44),.WL(WL143));
sram_cell_6t_5 inst_cell_143_45 (.BL(BL45),.BLN(BLN45),.WL(WL143));
sram_cell_6t_5 inst_cell_143_46 (.BL(BL46),.BLN(BLN46),.WL(WL143));
sram_cell_6t_5 inst_cell_143_47 (.BL(BL47),.BLN(BLN47),.WL(WL143));
sram_cell_6t_5 inst_cell_143_48 (.BL(BL48),.BLN(BLN48),.WL(WL143));
sram_cell_6t_5 inst_cell_143_49 (.BL(BL49),.BLN(BLN49),.WL(WL143));
sram_cell_6t_5 inst_cell_143_50 (.BL(BL50),.BLN(BLN50),.WL(WL143));
sram_cell_6t_5 inst_cell_143_51 (.BL(BL51),.BLN(BLN51),.WL(WL143));
sram_cell_6t_5 inst_cell_143_52 (.BL(BL52),.BLN(BLN52),.WL(WL143));
sram_cell_6t_5 inst_cell_143_53 (.BL(BL53),.BLN(BLN53),.WL(WL143));
sram_cell_6t_5 inst_cell_143_54 (.BL(BL54),.BLN(BLN54),.WL(WL143));
sram_cell_6t_5 inst_cell_143_55 (.BL(BL55),.BLN(BLN55),.WL(WL143));
sram_cell_6t_5 inst_cell_143_56 (.BL(BL56),.BLN(BLN56),.WL(WL143));
sram_cell_6t_5 inst_cell_143_57 (.BL(BL57),.BLN(BLN57),.WL(WL143));
sram_cell_6t_5 inst_cell_143_58 (.BL(BL58),.BLN(BLN58),.WL(WL143));
sram_cell_6t_5 inst_cell_143_59 (.BL(BL59),.BLN(BLN59),.WL(WL143));
sram_cell_6t_5 inst_cell_143_60 (.BL(BL60),.BLN(BLN60),.WL(WL143));
sram_cell_6t_5 inst_cell_143_61 (.BL(BL61),.BLN(BLN61),.WL(WL143));
sram_cell_6t_5 inst_cell_143_62 (.BL(BL62),.BLN(BLN62),.WL(WL143));
sram_cell_6t_5 inst_cell_143_63 (.BL(BL63),.BLN(BLN63),.WL(WL143));
sram_cell_6t_5 inst_cell_143_64 (.BL(BL64),.BLN(BLN64),.WL(WL143));
sram_cell_6t_5 inst_cell_143_65 (.BL(BL65),.BLN(BLN65),.WL(WL143));
sram_cell_6t_5 inst_cell_143_66 (.BL(BL66),.BLN(BLN66),.WL(WL143));
sram_cell_6t_5 inst_cell_143_67 (.BL(BL67),.BLN(BLN67),.WL(WL143));
sram_cell_6t_5 inst_cell_143_68 (.BL(BL68),.BLN(BLN68),.WL(WL143));
sram_cell_6t_5 inst_cell_143_69 (.BL(BL69),.BLN(BLN69),.WL(WL143));
sram_cell_6t_5 inst_cell_143_70 (.BL(BL70),.BLN(BLN70),.WL(WL143));
sram_cell_6t_5 inst_cell_143_71 (.BL(BL71),.BLN(BLN71),.WL(WL143));
sram_cell_6t_5 inst_cell_143_72 (.BL(BL72),.BLN(BLN72),.WL(WL143));
sram_cell_6t_5 inst_cell_143_73 (.BL(BL73),.BLN(BLN73),.WL(WL143));
sram_cell_6t_5 inst_cell_143_74 (.BL(BL74),.BLN(BLN74),.WL(WL143));
sram_cell_6t_5 inst_cell_143_75 (.BL(BL75),.BLN(BLN75),.WL(WL143));
sram_cell_6t_5 inst_cell_143_76 (.BL(BL76),.BLN(BLN76),.WL(WL143));
sram_cell_6t_5 inst_cell_143_77 (.BL(BL77),.BLN(BLN77),.WL(WL143));
sram_cell_6t_5 inst_cell_143_78 (.BL(BL78),.BLN(BLN78),.WL(WL143));
sram_cell_6t_5 inst_cell_143_79 (.BL(BL79),.BLN(BLN79),.WL(WL143));
sram_cell_6t_5 inst_cell_143_80 (.BL(BL80),.BLN(BLN80),.WL(WL143));
sram_cell_6t_5 inst_cell_143_81 (.BL(BL81),.BLN(BLN81),.WL(WL143));
sram_cell_6t_5 inst_cell_143_82 (.BL(BL82),.BLN(BLN82),.WL(WL143));
sram_cell_6t_5 inst_cell_143_83 (.BL(BL83),.BLN(BLN83),.WL(WL143));
sram_cell_6t_5 inst_cell_143_84 (.BL(BL84),.BLN(BLN84),.WL(WL143));
sram_cell_6t_5 inst_cell_143_85 (.BL(BL85),.BLN(BLN85),.WL(WL143));
sram_cell_6t_5 inst_cell_143_86 (.BL(BL86),.BLN(BLN86),.WL(WL143));
sram_cell_6t_5 inst_cell_143_87 (.BL(BL87),.BLN(BLN87),.WL(WL143));
sram_cell_6t_5 inst_cell_143_88 (.BL(BL88),.BLN(BLN88),.WL(WL143));
sram_cell_6t_5 inst_cell_143_89 (.BL(BL89),.BLN(BLN89),.WL(WL143));
sram_cell_6t_5 inst_cell_143_90 (.BL(BL90),.BLN(BLN90),.WL(WL143));
sram_cell_6t_5 inst_cell_143_91 (.BL(BL91),.BLN(BLN91),.WL(WL143));
sram_cell_6t_5 inst_cell_143_92 (.BL(BL92),.BLN(BLN92),.WL(WL143));
sram_cell_6t_5 inst_cell_143_93 (.BL(BL93),.BLN(BLN93),.WL(WL143));
sram_cell_6t_5 inst_cell_143_94 (.BL(BL94),.BLN(BLN94),.WL(WL143));
sram_cell_6t_5 inst_cell_143_95 (.BL(BL95),.BLN(BLN95),.WL(WL143));
sram_cell_6t_5 inst_cell_143_96 (.BL(BL96),.BLN(BLN96),.WL(WL143));
sram_cell_6t_5 inst_cell_143_97 (.BL(BL97),.BLN(BLN97),.WL(WL143));
sram_cell_6t_5 inst_cell_143_98 (.BL(BL98),.BLN(BLN98),.WL(WL143));
sram_cell_6t_5 inst_cell_143_99 (.BL(BL99),.BLN(BLN99),.WL(WL143));
sram_cell_6t_5 inst_cell_143_100 (.BL(BL100),.BLN(BLN100),.WL(WL143));
sram_cell_6t_5 inst_cell_143_101 (.BL(BL101),.BLN(BLN101),.WL(WL143));
sram_cell_6t_5 inst_cell_143_102 (.BL(BL102),.BLN(BLN102),.WL(WL143));
sram_cell_6t_5 inst_cell_143_103 (.BL(BL103),.BLN(BLN103),.WL(WL143));
sram_cell_6t_5 inst_cell_143_104 (.BL(BL104),.BLN(BLN104),.WL(WL143));
sram_cell_6t_5 inst_cell_143_105 (.BL(BL105),.BLN(BLN105),.WL(WL143));
sram_cell_6t_5 inst_cell_143_106 (.BL(BL106),.BLN(BLN106),.WL(WL143));
sram_cell_6t_5 inst_cell_143_107 (.BL(BL107),.BLN(BLN107),.WL(WL143));
sram_cell_6t_5 inst_cell_143_108 (.BL(BL108),.BLN(BLN108),.WL(WL143));
sram_cell_6t_5 inst_cell_143_109 (.BL(BL109),.BLN(BLN109),.WL(WL143));
sram_cell_6t_5 inst_cell_143_110 (.BL(BL110),.BLN(BLN110),.WL(WL143));
sram_cell_6t_5 inst_cell_143_111 (.BL(BL111),.BLN(BLN111),.WL(WL143));
sram_cell_6t_5 inst_cell_143_112 (.BL(BL112),.BLN(BLN112),.WL(WL143));
sram_cell_6t_5 inst_cell_143_113 (.BL(BL113),.BLN(BLN113),.WL(WL143));
sram_cell_6t_5 inst_cell_143_114 (.BL(BL114),.BLN(BLN114),.WL(WL143));
sram_cell_6t_5 inst_cell_143_115 (.BL(BL115),.BLN(BLN115),.WL(WL143));
sram_cell_6t_5 inst_cell_143_116 (.BL(BL116),.BLN(BLN116),.WL(WL143));
sram_cell_6t_5 inst_cell_143_117 (.BL(BL117),.BLN(BLN117),.WL(WL143));
sram_cell_6t_5 inst_cell_143_118 (.BL(BL118),.BLN(BLN118),.WL(WL143));
sram_cell_6t_5 inst_cell_143_119 (.BL(BL119),.BLN(BLN119),.WL(WL143));
sram_cell_6t_5 inst_cell_143_120 (.BL(BL120),.BLN(BLN120),.WL(WL143));
sram_cell_6t_5 inst_cell_143_121 (.BL(BL121),.BLN(BLN121),.WL(WL143));
sram_cell_6t_5 inst_cell_143_122 (.BL(BL122),.BLN(BLN122),.WL(WL143));
sram_cell_6t_5 inst_cell_143_123 (.BL(BL123),.BLN(BLN123),.WL(WL143));
sram_cell_6t_5 inst_cell_143_124 (.BL(BL124),.BLN(BLN124),.WL(WL143));
sram_cell_6t_5 inst_cell_143_125 (.BL(BL125),.BLN(BLN125),.WL(WL143));
sram_cell_6t_5 inst_cell_143_126 (.BL(BL126),.BLN(BLN126),.WL(WL143));
sram_cell_6t_5 inst_cell_143_127 (.BL(BL127),.BLN(BLN127),.WL(WL143));
sram_cell_6t_5 inst_cell_144_0 (.BL(BL0),.BLN(BLN0),.WL(WL144));
sram_cell_6t_5 inst_cell_144_1 (.BL(BL1),.BLN(BLN1),.WL(WL144));
sram_cell_6t_5 inst_cell_144_2 (.BL(BL2),.BLN(BLN2),.WL(WL144));
sram_cell_6t_5 inst_cell_144_3 (.BL(BL3),.BLN(BLN3),.WL(WL144));
sram_cell_6t_5 inst_cell_144_4 (.BL(BL4),.BLN(BLN4),.WL(WL144));
sram_cell_6t_5 inst_cell_144_5 (.BL(BL5),.BLN(BLN5),.WL(WL144));
sram_cell_6t_5 inst_cell_144_6 (.BL(BL6),.BLN(BLN6),.WL(WL144));
sram_cell_6t_5 inst_cell_144_7 (.BL(BL7),.BLN(BLN7),.WL(WL144));
sram_cell_6t_5 inst_cell_144_8 (.BL(BL8),.BLN(BLN8),.WL(WL144));
sram_cell_6t_5 inst_cell_144_9 (.BL(BL9),.BLN(BLN9),.WL(WL144));
sram_cell_6t_5 inst_cell_144_10 (.BL(BL10),.BLN(BLN10),.WL(WL144));
sram_cell_6t_5 inst_cell_144_11 (.BL(BL11),.BLN(BLN11),.WL(WL144));
sram_cell_6t_5 inst_cell_144_12 (.BL(BL12),.BLN(BLN12),.WL(WL144));
sram_cell_6t_5 inst_cell_144_13 (.BL(BL13),.BLN(BLN13),.WL(WL144));
sram_cell_6t_5 inst_cell_144_14 (.BL(BL14),.BLN(BLN14),.WL(WL144));
sram_cell_6t_5 inst_cell_144_15 (.BL(BL15),.BLN(BLN15),.WL(WL144));
sram_cell_6t_5 inst_cell_144_16 (.BL(BL16),.BLN(BLN16),.WL(WL144));
sram_cell_6t_5 inst_cell_144_17 (.BL(BL17),.BLN(BLN17),.WL(WL144));
sram_cell_6t_5 inst_cell_144_18 (.BL(BL18),.BLN(BLN18),.WL(WL144));
sram_cell_6t_5 inst_cell_144_19 (.BL(BL19),.BLN(BLN19),.WL(WL144));
sram_cell_6t_5 inst_cell_144_20 (.BL(BL20),.BLN(BLN20),.WL(WL144));
sram_cell_6t_5 inst_cell_144_21 (.BL(BL21),.BLN(BLN21),.WL(WL144));
sram_cell_6t_5 inst_cell_144_22 (.BL(BL22),.BLN(BLN22),.WL(WL144));
sram_cell_6t_5 inst_cell_144_23 (.BL(BL23),.BLN(BLN23),.WL(WL144));
sram_cell_6t_5 inst_cell_144_24 (.BL(BL24),.BLN(BLN24),.WL(WL144));
sram_cell_6t_5 inst_cell_144_25 (.BL(BL25),.BLN(BLN25),.WL(WL144));
sram_cell_6t_5 inst_cell_144_26 (.BL(BL26),.BLN(BLN26),.WL(WL144));
sram_cell_6t_5 inst_cell_144_27 (.BL(BL27),.BLN(BLN27),.WL(WL144));
sram_cell_6t_5 inst_cell_144_28 (.BL(BL28),.BLN(BLN28),.WL(WL144));
sram_cell_6t_5 inst_cell_144_29 (.BL(BL29),.BLN(BLN29),.WL(WL144));
sram_cell_6t_5 inst_cell_144_30 (.BL(BL30),.BLN(BLN30),.WL(WL144));
sram_cell_6t_5 inst_cell_144_31 (.BL(BL31),.BLN(BLN31),.WL(WL144));
sram_cell_6t_5 inst_cell_144_32 (.BL(BL32),.BLN(BLN32),.WL(WL144));
sram_cell_6t_5 inst_cell_144_33 (.BL(BL33),.BLN(BLN33),.WL(WL144));
sram_cell_6t_5 inst_cell_144_34 (.BL(BL34),.BLN(BLN34),.WL(WL144));
sram_cell_6t_5 inst_cell_144_35 (.BL(BL35),.BLN(BLN35),.WL(WL144));
sram_cell_6t_5 inst_cell_144_36 (.BL(BL36),.BLN(BLN36),.WL(WL144));
sram_cell_6t_5 inst_cell_144_37 (.BL(BL37),.BLN(BLN37),.WL(WL144));
sram_cell_6t_5 inst_cell_144_38 (.BL(BL38),.BLN(BLN38),.WL(WL144));
sram_cell_6t_5 inst_cell_144_39 (.BL(BL39),.BLN(BLN39),.WL(WL144));
sram_cell_6t_5 inst_cell_144_40 (.BL(BL40),.BLN(BLN40),.WL(WL144));
sram_cell_6t_5 inst_cell_144_41 (.BL(BL41),.BLN(BLN41),.WL(WL144));
sram_cell_6t_5 inst_cell_144_42 (.BL(BL42),.BLN(BLN42),.WL(WL144));
sram_cell_6t_5 inst_cell_144_43 (.BL(BL43),.BLN(BLN43),.WL(WL144));
sram_cell_6t_5 inst_cell_144_44 (.BL(BL44),.BLN(BLN44),.WL(WL144));
sram_cell_6t_5 inst_cell_144_45 (.BL(BL45),.BLN(BLN45),.WL(WL144));
sram_cell_6t_5 inst_cell_144_46 (.BL(BL46),.BLN(BLN46),.WL(WL144));
sram_cell_6t_5 inst_cell_144_47 (.BL(BL47),.BLN(BLN47),.WL(WL144));
sram_cell_6t_5 inst_cell_144_48 (.BL(BL48),.BLN(BLN48),.WL(WL144));
sram_cell_6t_5 inst_cell_144_49 (.BL(BL49),.BLN(BLN49),.WL(WL144));
sram_cell_6t_5 inst_cell_144_50 (.BL(BL50),.BLN(BLN50),.WL(WL144));
sram_cell_6t_5 inst_cell_144_51 (.BL(BL51),.BLN(BLN51),.WL(WL144));
sram_cell_6t_5 inst_cell_144_52 (.BL(BL52),.BLN(BLN52),.WL(WL144));
sram_cell_6t_5 inst_cell_144_53 (.BL(BL53),.BLN(BLN53),.WL(WL144));
sram_cell_6t_5 inst_cell_144_54 (.BL(BL54),.BLN(BLN54),.WL(WL144));
sram_cell_6t_5 inst_cell_144_55 (.BL(BL55),.BLN(BLN55),.WL(WL144));
sram_cell_6t_5 inst_cell_144_56 (.BL(BL56),.BLN(BLN56),.WL(WL144));
sram_cell_6t_5 inst_cell_144_57 (.BL(BL57),.BLN(BLN57),.WL(WL144));
sram_cell_6t_5 inst_cell_144_58 (.BL(BL58),.BLN(BLN58),.WL(WL144));
sram_cell_6t_5 inst_cell_144_59 (.BL(BL59),.BLN(BLN59),.WL(WL144));
sram_cell_6t_5 inst_cell_144_60 (.BL(BL60),.BLN(BLN60),.WL(WL144));
sram_cell_6t_5 inst_cell_144_61 (.BL(BL61),.BLN(BLN61),.WL(WL144));
sram_cell_6t_5 inst_cell_144_62 (.BL(BL62),.BLN(BLN62),.WL(WL144));
sram_cell_6t_5 inst_cell_144_63 (.BL(BL63),.BLN(BLN63),.WL(WL144));
sram_cell_6t_5 inst_cell_144_64 (.BL(BL64),.BLN(BLN64),.WL(WL144));
sram_cell_6t_5 inst_cell_144_65 (.BL(BL65),.BLN(BLN65),.WL(WL144));
sram_cell_6t_5 inst_cell_144_66 (.BL(BL66),.BLN(BLN66),.WL(WL144));
sram_cell_6t_5 inst_cell_144_67 (.BL(BL67),.BLN(BLN67),.WL(WL144));
sram_cell_6t_5 inst_cell_144_68 (.BL(BL68),.BLN(BLN68),.WL(WL144));
sram_cell_6t_5 inst_cell_144_69 (.BL(BL69),.BLN(BLN69),.WL(WL144));
sram_cell_6t_5 inst_cell_144_70 (.BL(BL70),.BLN(BLN70),.WL(WL144));
sram_cell_6t_5 inst_cell_144_71 (.BL(BL71),.BLN(BLN71),.WL(WL144));
sram_cell_6t_5 inst_cell_144_72 (.BL(BL72),.BLN(BLN72),.WL(WL144));
sram_cell_6t_5 inst_cell_144_73 (.BL(BL73),.BLN(BLN73),.WL(WL144));
sram_cell_6t_5 inst_cell_144_74 (.BL(BL74),.BLN(BLN74),.WL(WL144));
sram_cell_6t_5 inst_cell_144_75 (.BL(BL75),.BLN(BLN75),.WL(WL144));
sram_cell_6t_5 inst_cell_144_76 (.BL(BL76),.BLN(BLN76),.WL(WL144));
sram_cell_6t_5 inst_cell_144_77 (.BL(BL77),.BLN(BLN77),.WL(WL144));
sram_cell_6t_5 inst_cell_144_78 (.BL(BL78),.BLN(BLN78),.WL(WL144));
sram_cell_6t_5 inst_cell_144_79 (.BL(BL79),.BLN(BLN79),.WL(WL144));
sram_cell_6t_5 inst_cell_144_80 (.BL(BL80),.BLN(BLN80),.WL(WL144));
sram_cell_6t_5 inst_cell_144_81 (.BL(BL81),.BLN(BLN81),.WL(WL144));
sram_cell_6t_5 inst_cell_144_82 (.BL(BL82),.BLN(BLN82),.WL(WL144));
sram_cell_6t_5 inst_cell_144_83 (.BL(BL83),.BLN(BLN83),.WL(WL144));
sram_cell_6t_5 inst_cell_144_84 (.BL(BL84),.BLN(BLN84),.WL(WL144));
sram_cell_6t_5 inst_cell_144_85 (.BL(BL85),.BLN(BLN85),.WL(WL144));
sram_cell_6t_5 inst_cell_144_86 (.BL(BL86),.BLN(BLN86),.WL(WL144));
sram_cell_6t_5 inst_cell_144_87 (.BL(BL87),.BLN(BLN87),.WL(WL144));
sram_cell_6t_5 inst_cell_144_88 (.BL(BL88),.BLN(BLN88),.WL(WL144));
sram_cell_6t_5 inst_cell_144_89 (.BL(BL89),.BLN(BLN89),.WL(WL144));
sram_cell_6t_5 inst_cell_144_90 (.BL(BL90),.BLN(BLN90),.WL(WL144));
sram_cell_6t_5 inst_cell_144_91 (.BL(BL91),.BLN(BLN91),.WL(WL144));
sram_cell_6t_5 inst_cell_144_92 (.BL(BL92),.BLN(BLN92),.WL(WL144));
sram_cell_6t_5 inst_cell_144_93 (.BL(BL93),.BLN(BLN93),.WL(WL144));
sram_cell_6t_5 inst_cell_144_94 (.BL(BL94),.BLN(BLN94),.WL(WL144));
sram_cell_6t_5 inst_cell_144_95 (.BL(BL95),.BLN(BLN95),.WL(WL144));
sram_cell_6t_5 inst_cell_144_96 (.BL(BL96),.BLN(BLN96),.WL(WL144));
sram_cell_6t_5 inst_cell_144_97 (.BL(BL97),.BLN(BLN97),.WL(WL144));
sram_cell_6t_5 inst_cell_144_98 (.BL(BL98),.BLN(BLN98),.WL(WL144));
sram_cell_6t_5 inst_cell_144_99 (.BL(BL99),.BLN(BLN99),.WL(WL144));
sram_cell_6t_5 inst_cell_144_100 (.BL(BL100),.BLN(BLN100),.WL(WL144));
sram_cell_6t_5 inst_cell_144_101 (.BL(BL101),.BLN(BLN101),.WL(WL144));
sram_cell_6t_5 inst_cell_144_102 (.BL(BL102),.BLN(BLN102),.WL(WL144));
sram_cell_6t_5 inst_cell_144_103 (.BL(BL103),.BLN(BLN103),.WL(WL144));
sram_cell_6t_5 inst_cell_144_104 (.BL(BL104),.BLN(BLN104),.WL(WL144));
sram_cell_6t_5 inst_cell_144_105 (.BL(BL105),.BLN(BLN105),.WL(WL144));
sram_cell_6t_5 inst_cell_144_106 (.BL(BL106),.BLN(BLN106),.WL(WL144));
sram_cell_6t_5 inst_cell_144_107 (.BL(BL107),.BLN(BLN107),.WL(WL144));
sram_cell_6t_5 inst_cell_144_108 (.BL(BL108),.BLN(BLN108),.WL(WL144));
sram_cell_6t_5 inst_cell_144_109 (.BL(BL109),.BLN(BLN109),.WL(WL144));
sram_cell_6t_5 inst_cell_144_110 (.BL(BL110),.BLN(BLN110),.WL(WL144));
sram_cell_6t_5 inst_cell_144_111 (.BL(BL111),.BLN(BLN111),.WL(WL144));
sram_cell_6t_5 inst_cell_144_112 (.BL(BL112),.BLN(BLN112),.WL(WL144));
sram_cell_6t_5 inst_cell_144_113 (.BL(BL113),.BLN(BLN113),.WL(WL144));
sram_cell_6t_5 inst_cell_144_114 (.BL(BL114),.BLN(BLN114),.WL(WL144));
sram_cell_6t_5 inst_cell_144_115 (.BL(BL115),.BLN(BLN115),.WL(WL144));
sram_cell_6t_5 inst_cell_144_116 (.BL(BL116),.BLN(BLN116),.WL(WL144));
sram_cell_6t_5 inst_cell_144_117 (.BL(BL117),.BLN(BLN117),.WL(WL144));
sram_cell_6t_5 inst_cell_144_118 (.BL(BL118),.BLN(BLN118),.WL(WL144));
sram_cell_6t_5 inst_cell_144_119 (.BL(BL119),.BLN(BLN119),.WL(WL144));
sram_cell_6t_5 inst_cell_144_120 (.BL(BL120),.BLN(BLN120),.WL(WL144));
sram_cell_6t_5 inst_cell_144_121 (.BL(BL121),.BLN(BLN121),.WL(WL144));
sram_cell_6t_5 inst_cell_144_122 (.BL(BL122),.BLN(BLN122),.WL(WL144));
sram_cell_6t_5 inst_cell_144_123 (.BL(BL123),.BLN(BLN123),.WL(WL144));
sram_cell_6t_5 inst_cell_144_124 (.BL(BL124),.BLN(BLN124),.WL(WL144));
sram_cell_6t_5 inst_cell_144_125 (.BL(BL125),.BLN(BLN125),.WL(WL144));
sram_cell_6t_5 inst_cell_144_126 (.BL(BL126),.BLN(BLN126),.WL(WL144));
sram_cell_6t_5 inst_cell_144_127 (.BL(BL127),.BLN(BLN127),.WL(WL144));
sram_cell_6t_5 inst_cell_145_0 (.BL(BL0),.BLN(BLN0),.WL(WL145));
sram_cell_6t_5 inst_cell_145_1 (.BL(BL1),.BLN(BLN1),.WL(WL145));
sram_cell_6t_5 inst_cell_145_2 (.BL(BL2),.BLN(BLN2),.WL(WL145));
sram_cell_6t_5 inst_cell_145_3 (.BL(BL3),.BLN(BLN3),.WL(WL145));
sram_cell_6t_5 inst_cell_145_4 (.BL(BL4),.BLN(BLN4),.WL(WL145));
sram_cell_6t_5 inst_cell_145_5 (.BL(BL5),.BLN(BLN5),.WL(WL145));
sram_cell_6t_5 inst_cell_145_6 (.BL(BL6),.BLN(BLN6),.WL(WL145));
sram_cell_6t_5 inst_cell_145_7 (.BL(BL7),.BLN(BLN7),.WL(WL145));
sram_cell_6t_5 inst_cell_145_8 (.BL(BL8),.BLN(BLN8),.WL(WL145));
sram_cell_6t_5 inst_cell_145_9 (.BL(BL9),.BLN(BLN9),.WL(WL145));
sram_cell_6t_5 inst_cell_145_10 (.BL(BL10),.BLN(BLN10),.WL(WL145));
sram_cell_6t_5 inst_cell_145_11 (.BL(BL11),.BLN(BLN11),.WL(WL145));
sram_cell_6t_5 inst_cell_145_12 (.BL(BL12),.BLN(BLN12),.WL(WL145));
sram_cell_6t_5 inst_cell_145_13 (.BL(BL13),.BLN(BLN13),.WL(WL145));
sram_cell_6t_5 inst_cell_145_14 (.BL(BL14),.BLN(BLN14),.WL(WL145));
sram_cell_6t_5 inst_cell_145_15 (.BL(BL15),.BLN(BLN15),.WL(WL145));
sram_cell_6t_5 inst_cell_145_16 (.BL(BL16),.BLN(BLN16),.WL(WL145));
sram_cell_6t_5 inst_cell_145_17 (.BL(BL17),.BLN(BLN17),.WL(WL145));
sram_cell_6t_5 inst_cell_145_18 (.BL(BL18),.BLN(BLN18),.WL(WL145));
sram_cell_6t_5 inst_cell_145_19 (.BL(BL19),.BLN(BLN19),.WL(WL145));
sram_cell_6t_5 inst_cell_145_20 (.BL(BL20),.BLN(BLN20),.WL(WL145));
sram_cell_6t_5 inst_cell_145_21 (.BL(BL21),.BLN(BLN21),.WL(WL145));
sram_cell_6t_5 inst_cell_145_22 (.BL(BL22),.BLN(BLN22),.WL(WL145));
sram_cell_6t_5 inst_cell_145_23 (.BL(BL23),.BLN(BLN23),.WL(WL145));
sram_cell_6t_5 inst_cell_145_24 (.BL(BL24),.BLN(BLN24),.WL(WL145));
sram_cell_6t_5 inst_cell_145_25 (.BL(BL25),.BLN(BLN25),.WL(WL145));
sram_cell_6t_5 inst_cell_145_26 (.BL(BL26),.BLN(BLN26),.WL(WL145));
sram_cell_6t_5 inst_cell_145_27 (.BL(BL27),.BLN(BLN27),.WL(WL145));
sram_cell_6t_5 inst_cell_145_28 (.BL(BL28),.BLN(BLN28),.WL(WL145));
sram_cell_6t_5 inst_cell_145_29 (.BL(BL29),.BLN(BLN29),.WL(WL145));
sram_cell_6t_5 inst_cell_145_30 (.BL(BL30),.BLN(BLN30),.WL(WL145));
sram_cell_6t_5 inst_cell_145_31 (.BL(BL31),.BLN(BLN31),.WL(WL145));
sram_cell_6t_5 inst_cell_145_32 (.BL(BL32),.BLN(BLN32),.WL(WL145));
sram_cell_6t_5 inst_cell_145_33 (.BL(BL33),.BLN(BLN33),.WL(WL145));
sram_cell_6t_5 inst_cell_145_34 (.BL(BL34),.BLN(BLN34),.WL(WL145));
sram_cell_6t_5 inst_cell_145_35 (.BL(BL35),.BLN(BLN35),.WL(WL145));
sram_cell_6t_5 inst_cell_145_36 (.BL(BL36),.BLN(BLN36),.WL(WL145));
sram_cell_6t_5 inst_cell_145_37 (.BL(BL37),.BLN(BLN37),.WL(WL145));
sram_cell_6t_5 inst_cell_145_38 (.BL(BL38),.BLN(BLN38),.WL(WL145));
sram_cell_6t_5 inst_cell_145_39 (.BL(BL39),.BLN(BLN39),.WL(WL145));
sram_cell_6t_5 inst_cell_145_40 (.BL(BL40),.BLN(BLN40),.WL(WL145));
sram_cell_6t_5 inst_cell_145_41 (.BL(BL41),.BLN(BLN41),.WL(WL145));
sram_cell_6t_5 inst_cell_145_42 (.BL(BL42),.BLN(BLN42),.WL(WL145));
sram_cell_6t_5 inst_cell_145_43 (.BL(BL43),.BLN(BLN43),.WL(WL145));
sram_cell_6t_5 inst_cell_145_44 (.BL(BL44),.BLN(BLN44),.WL(WL145));
sram_cell_6t_5 inst_cell_145_45 (.BL(BL45),.BLN(BLN45),.WL(WL145));
sram_cell_6t_5 inst_cell_145_46 (.BL(BL46),.BLN(BLN46),.WL(WL145));
sram_cell_6t_5 inst_cell_145_47 (.BL(BL47),.BLN(BLN47),.WL(WL145));
sram_cell_6t_5 inst_cell_145_48 (.BL(BL48),.BLN(BLN48),.WL(WL145));
sram_cell_6t_5 inst_cell_145_49 (.BL(BL49),.BLN(BLN49),.WL(WL145));
sram_cell_6t_5 inst_cell_145_50 (.BL(BL50),.BLN(BLN50),.WL(WL145));
sram_cell_6t_5 inst_cell_145_51 (.BL(BL51),.BLN(BLN51),.WL(WL145));
sram_cell_6t_5 inst_cell_145_52 (.BL(BL52),.BLN(BLN52),.WL(WL145));
sram_cell_6t_5 inst_cell_145_53 (.BL(BL53),.BLN(BLN53),.WL(WL145));
sram_cell_6t_5 inst_cell_145_54 (.BL(BL54),.BLN(BLN54),.WL(WL145));
sram_cell_6t_5 inst_cell_145_55 (.BL(BL55),.BLN(BLN55),.WL(WL145));
sram_cell_6t_5 inst_cell_145_56 (.BL(BL56),.BLN(BLN56),.WL(WL145));
sram_cell_6t_5 inst_cell_145_57 (.BL(BL57),.BLN(BLN57),.WL(WL145));
sram_cell_6t_5 inst_cell_145_58 (.BL(BL58),.BLN(BLN58),.WL(WL145));
sram_cell_6t_5 inst_cell_145_59 (.BL(BL59),.BLN(BLN59),.WL(WL145));
sram_cell_6t_5 inst_cell_145_60 (.BL(BL60),.BLN(BLN60),.WL(WL145));
sram_cell_6t_5 inst_cell_145_61 (.BL(BL61),.BLN(BLN61),.WL(WL145));
sram_cell_6t_5 inst_cell_145_62 (.BL(BL62),.BLN(BLN62),.WL(WL145));
sram_cell_6t_5 inst_cell_145_63 (.BL(BL63),.BLN(BLN63),.WL(WL145));
sram_cell_6t_5 inst_cell_145_64 (.BL(BL64),.BLN(BLN64),.WL(WL145));
sram_cell_6t_5 inst_cell_145_65 (.BL(BL65),.BLN(BLN65),.WL(WL145));
sram_cell_6t_5 inst_cell_145_66 (.BL(BL66),.BLN(BLN66),.WL(WL145));
sram_cell_6t_5 inst_cell_145_67 (.BL(BL67),.BLN(BLN67),.WL(WL145));
sram_cell_6t_5 inst_cell_145_68 (.BL(BL68),.BLN(BLN68),.WL(WL145));
sram_cell_6t_5 inst_cell_145_69 (.BL(BL69),.BLN(BLN69),.WL(WL145));
sram_cell_6t_5 inst_cell_145_70 (.BL(BL70),.BLN(BLN70),.WL(WL145));
sram_cell_6t_5 inst_cell_145_71 (.BL(BL71),.BLN(BLN71),.WL(WL145));
sram_cell_6t_5 inst_cell_145_72 (.BL(BL72),.BLN(BLN72),.WL(WL145));
sram_cell_6t_5 inst_cell_145_73 (.BL(BL73),.BLN(BLN73),.WL(WL145));
sram_cell_6t_5 inst_cell_145_74 (.BL(BL74),.BLN(BLN74),.WL(WL145));
sram_cell_6t_5 inst_cell_145_75 (.BL(BL75),.BLN(BLN75),.WL(WL145));
sram_cell_6t_5 inst_cell_145_76 (.BL(BL76),.BLN(BLN76),.WL(WL145));
sram_cell_6t_5 inst_cell_145_77 (.BL(BL77),.BLN(BLN77),.WL(WL145));
sram_cell_6t_5 inst_cell_145_78 (.BL(BL78),.BLN(BLN78),.WL(WL145));
sram_cell_6t_5 inst_cell_145_79 (.BL(BL79),.BLN(BLN79),.WL(WL145));
sram_cell_6t_5 inst_cell_145_80 (.BL(BL80),.BLN(BLN80),.WL(WL145));
sram_cell_6t_5 inst_cell_145_81 (.BL(BL81),.BLN(BLN81),.WL(WL145));
sram_cell_6t_5 inst_cell_145_82 (.BL(BL82),.BLN(BLN82),.WL(WL145));
sram_cell_6t_5 inst_cell_145_83 (.BL(BL83),.BLN(BLN83),.WL(WL145));
sram_cell_6t_5 inst_cell_145_84 (.BL(BL84),.BLN(BLN84),.WL(WL145));
sram_cell_6t_5 inst_cell_145_85 (.BL(BL85),.BLN(BLN85),.WL(WL145));
sram_cell_6t_5 inst_cell_145_86 (.BL(BL86),.BLN(BLN86),.WL(WL145));
sram_cell_6t_5 inst_cell_145_87 (.BL(BL87),.BLN(BLN87),.WL(WL145));
sram_cell_6t_5 inst_cell_145_88 (.BL(BL88),.BLN(BLN88),.WL(WL145));
sram_cell_6t_5 inst_cell_145_89 (.BL(BL89),.BLN(BLN89),.WL(WL145));
sram_cell_6t_5 inst_cell_145_90 (.BL(BL90),.BLN(BLN90),.WL(WL145));
sram_cell_6t_5 inst_cell_145_91 (.BL(BL91),.BLN(BLN91),.WL(WL145));
sram_cell_6t_5 inst_cell_145_92 (.BL(BL92),.BLN(BLN92),.WL(WL145));
sram_cell_6t_5 inst_cell_145_93 (.BL(BL93),.BLN(BLN93),.WL(WL145));
sram_cell_6t_5 inst_cell_145_94 (.BL(BL94),.BLN(BLN94),.WL(WL145));
sram_cell_6t_5 inst_cell_145_95 (.BL(BL95),.BLN(BLN95),.WL(WL145));
sram_cell_6t_5 inst_cell_145_96 (.BL(BL96),.BLN(BLN96),.WL(WL145));
sram_cell_6t_5 inst_cell_145_97 (.BL(BL97),.BLN(BLN97),.WL(WL145));
sram_cell_6t_5 inst_cell_145_98 (.BL(BL98),.BLN(BLN98),.WL(WL145));
sram_cell_6t_5 inst_cell_145_99 (.BL(BL99),.BLN(BLN99),.WL(WL145));
sram_cell_6t_5 inst_cell_145_100 (.BL(BL100),.BLN(BLN100),.WL(WL145));
sram_cell_6t_5 inst_cell_145_101 (.BL(BL101),.BLN(BLN101),.WL(WL145));
sram_cell_6t_5 inst_cell_145_102 (.BL(BL102),.BLN(BLN102),.WL(WL145));
sram_cell_6t_5 inst_cell_145_103 (.BL(BL103),.BLN(BLN103),.WL(WL145));
sram_cell_6t_5 inst_cell_145_104 (.BL(BL104),.BLN(BLN104),.WL(WL145));
sram_cell_6t_5 inst_cell_145_105 (.BL(BL105),.BLN(BLN105),.WL(WL145));
sram_cell_6t_5 inst_cell_145_106 (.BL(BL106),.BLN(BLN106),.WL(WL145));
sram_cell_6t_5 inst_cell_145_107 (.BL(BL107),.BLN(BLN107),.WL(WL145));
sram_cell_6t_5 inst_cell_145_108 (.BL(BL108),.BLN(BLN108),.WL(WL145));
sram_cell_6t_5 inst_cell_145_109 (.BL(BL109),.BLN(BLN109),.WL(WL145));
sram_cell_6t_5 inst_cell_145_110 (.BL(BL110),.BLN(BLN110),.WL(WL145));
sram_cell_6t_5 inst_cell_145_111 (.BL(BL111),.BLN(BLN111),.WL(WL145));
sram_cell_6t_5 inst_cell_145_112 (.BL(BL112),.BLN(BLN112),.WL(WL145));
sram_cell_6t_5 inst_cell_145_113 (.BL(BL113),.BLN(BLN113),.WL(WL145));
sram_cell_6t_5 inst_cell_145_114 (.BL(BL114),.BLN(BLN114),.WL(WL145));
sram_cell_6t_5 inst_cell_145_115 (.BL(BL115),.BLN(BLN115),.WL(WL145));
sram_cell_6t_5 inst_cell_145_116 (.BL(BL116),.BLN(BLN116),.WL(WL145));
sram_cell_6t_5 inst_cell_145_117 (.BL(BL117),.BLN(BLN117),.WL(WL145));
sram_cell_6t_5 inst_cell_145_118 (.BL(BL118),.BLN(BLN118),.WL(WL145));
sram_cell_6t_5 inst_cell_145_119 (.BL(BL119),.BLN(BLN119),.WL(WL145));
sram_cell_6t_5 inst_cell_145_120 (.BL(BL120),.BLN(BLN120),.WL(WL145));
sram_cell_6t_5 inst_cell_145_121 (.BL(BL121),.BLN(BLN121),.WL(WL145));
sram_cell_6t_5 inst_cell_145_122 (.BL(BL122),.BLN(BLN122),.WL(WL145));
sram_cell_6t_5 inst_cell_145_123 (.BL(BL123),.BLN(BLN123),.WL(WL145));
sram_cell_6t_5 inst_cell_145_124 (.BL(BL124),.BLN(BLN124),.WL(WL145));
sram_cell_6t_5 inst_cell_145_125 (.BL(BL125),.BLN(BLN125),.WL(WL145));
sram_cell_6t_5 inst_cell_145_126 (.BL(BL126),.BLN(BLN126),.WL(WL145));
sram_cell_6t_5 inst_cell_145_127 (.BL(BL127),.BLN(BLN127),.WL(WL145));
sram_cell_6t_5 inst_cell_146_0 (.BL(BL0),.BLN(BLN0),.WL(WL146));
sram_cell_6t_5 inst_cell_146_1 (.BL(BL1),.BLN(BLN1),.WL(WL146));
sram_cell_6t_5 inst_cell_146_2 (.BL(BL2),.BLN(BLN2),.WL(WL146));
sram_cell_6t_5 inst_cell_146_3 (.BL(BL3),.BLN(BLN3),.WL(WL146));
sram_cell_6t_5 inst_cell_146_4 (.BL(BL4),.BLN(BLN4),.WL(WL146));
sram_cell_6t_5 inst_cell_146_5 (.BL(BL5),.BLN(BLN5),.WL(WL146));
sram_cell_6t_5 inst_cell_146_6 (.BL(BL6),.BLN(BLN6),.WL(WL146));
sram_cell_6t_5 inst_cell_146_7 (.BL(BL7),.BLN(BLN7),.WL(WL146));
sram_cell_6t_5 inst_cell_146_8 (.BL(BL8),.BLN(BLN8),.WL(WL146));
sram_cell_6t_5 inst_cell_146_9 (.BL(BL9),.BLN(BLN9),.WL(WL146));
sram_cell_6t_5 inst_cell_146_10 (.BL(BL10),.BLN(BLN10),.WL(WL146));
sram_cell_6t_5 inst_cell_146_11 (.BL(BL11),.BLN(BLN11),.WL(WL146));
sram_cell_6t_5 inst_cell_146_12 (.BL(BL12),.BLN(BLN12),.WL(WL146));
sram_cell_6t_5 inst_cell_146_13 (.BL(BL13),.BLN(BLN13),.WL(WL146));
sram_cell_6t_5 inst_cell_146_14 (.BL(BL14),.BLN(BLN14),.WL(WL146));
sram_cell_6t_5 inst_cell_146_15 (.BL(BL15),.BLN(BLN15),.WL(WL146));
sram_cell_6t_5 inst_cell_146_16 (.BL(BL16),.BLN(BLN16),.WL(WL146));
sram_cell_6t_5 inst_cell_146_17 (.BL(BL17),.BLN(BLN17),.WL(WL146));
sram_cell_6t_5 inst_cell_146_18 (.BL(BL18),.BLN(BLN18),.WL(WL146));
sram_cell_6t_5 inst_cell_146_19 (.BL(BL19),.BLN(BLN19),.WL(WL146));
sram_cell_6t_5 inst_cell_146_20 (.BL(BL20),.BLN(BLN20),.WL(WL146));
sram_cell_6t_5 inst_cell_146_21 (.BL(BL21),.BLN(BLN21),.WL(WL146));
sram_cell_6t_5 inst_cell_146_22 (.BL(BL22),.BLN(BLN22),.WL(WL146));
sram_cell_6t_5 inst_cell_146_23 (.BL(BL23),.BLN(BLN23),.WL(WL146));
sram_cell_6t_5 inst_cell_146_24 (.BL(BL24),.BLN(BLN24),.WL(WL146));
sram_cell_6t_5 inst_cell_146_25 (.BL(BL25),.BLN(BLN25),.WL(WL146));
sram_cell_6t_5 inst_cell_146_26 (.BL(BL26),.BLN(BLN26),.WL(WL146));
sram_cell_6t_5 inst_cell_146_27 (.BL(BL27),.BLN(BLN27),.WL(WL146));
sram_cell_6t_5 inst_cell_146_28 (.BL(BL28),.BLN(BLN28),.WL(WL146));
sram_cell_6t_5 inst_cell_146_29 (.BL(BL29),.BLN(BLN29),.WL(WL146));
sram_cell_6t_5 inst_cell_146_30 (.BL(BL30),.BLN(BLN30),.WL(WL146));
sram_cell_6t_5 inst_cell_146_31 (.BL(BL31),.BLN(BLN31),.WL(WL146));
sram_cell_6t_5 inst_cell_146_32 (.BL(BL32),.BLN(BLN32),.WL(WL146));
sram_cell_6t_5 inst_cell_146_33 (.BL(BL33),.BLN(BLN33),.WL(WL146));
sram_cell_6t_5 inst_cell_146_34 (.BL(BL34),.BLN(BLN34),.WL(WL146));
sram_cell_6t_5 inst_cell_146_35 (.BL(BL35),.BLN(BLN35),.WL(WL146));
sram_cell_6t_5 inst_cell_146_36 (.BL(BL36),.BLN(BLN36),.WL(WL146));
sram_cell_6t_5 inst_cell_146_37 (.BL(BL37),.BLN(BLN37),.WL(WL146));
sram_cell_6t_5 inst_cell_146_38 (.BL(BL38),.BLN(BLN38),.WL(WL146));
sram_cell_6t_5 inst_cell_146_39 (.BL(BL39),.BLN(BLN39),.WL(WL146));
sram_cell_6t_5 inst_cell_146_40 (.BL(BL40),.BLN(BLN40),.WL(WL146));
sram_cell_6t_5 inst_cell_146_41 (.BL(BL41),.BLN(BLN41),.WL(WL146));
sram_cell_6t_5 inst_cell_146_42 (.BL(BL42),.BLN(BLN42),.WL(WL146));
sram_cell_6t_5 inst_cell_146_43 (.BL(BL43),.BLN(BLN43),.WL(WL146));
sram_cell_6t_5 inst_cell_146_44 (.BL(BL44),.BLN(BLN44),.WL(WL146));
sram_cell_6t_5 inst_cell_146_45 (.BL(BL45),.BLN(BLN45),.WL(WL146));
sram_cell_6t_5 inst_cell_146_46 (.BL(BL46),.BLN(BLN46),.WL(WL146));
sram_cell_6t_5 inst_cell_146_47 (.BL(BL47),.BLN(BLN47),.WL(WL146));
sram_cell_6t_5 inst_cell_146_48 (.BL(BL48),.BLN(BLN48),.WL(WL146));
sram_cell_6t_5 inst_cell_146_49 (.BL(BL49),.BLN(BLN49),.WL(WL146));
sram_cell_6t_5 inst_cell_146_50 (.BL(BL50),.BLN(BLN50),.WL(WL146));
sram_cell_6t_5 inst_cell_146_51 (.BL(BL51),.BLN(BLN51),.WL(WL146));
sram_cell_6t_5 inst_cell_146_52 (.BL(BL52),.BLN(BLN52),.WL(WL146));
sram_cell_6t_5 inst_cell_146_53 (.BL(BL53),.BLN(BLN53),.WL(WL146));
sram_cell_6t_5 inst_cell_146_54 (.BL(BL54),.BLN(BLN54),.WL(WL146));
sram_cell_6t_5 inst_cell_146_55 (.BL(BL55),.BLN(BLN55),.WL(WL146));
sram_cell_6t_5 inst_cell_146_56 (.BL(BL56),.BLN(BLN56),.WL(WL146));
sram_cell_6t_5 inst_cell_146_57 (.BL(BL57),.BLN(BLN57),.WL(WL146));
sram_cell_6t_5 inst_cell_146_58 (.BL(BL58),.BLN(BLN58),.WL(WL146));
sram_cell_6t_5 inst_cell_146_59 (.BL(BL59),.BLN(BLN59),.WL(WL146));
sram_cell_6t_5 inst_cell_146_60 (.BL(BL60),.BLN(BLN60),.WL(WL146));
sram_cell_6t_5 inst_cell_146_61 (.BL(BL61),.BLN(BLN61),.WL(WL146));
sram_cell_6t_5 inst_cell_146_62 (.BL(BL62),.BLN(BLN62),.WL(WL146));
sram_cell_6t_5 inst_cell_146_63 (.BL(BL63),.BLN(BLN63),.WL(WL146));
sram_cell_6t_5 inst_cell_146_64 (.BL(BL64),.BLN(BLN64),.WL(WL146));
sram_cell_6t_5 inst_cell_146_65 (.BL(BL65),.BLN(BLN65),.WL(WL146));
sram_cell_6t_5 inst_cell_146_66 (.BL(BL66),.BLN(BLN66),.WL(WL146));
sram_cell_6t_5 inst_cell_146_67 (.BL(BL67),.BLN(BLN67),.WL(WL146));
sram_cell_6t_5 inst_cell_146_68 (.BL(BL68),.BLN(BLN68),.WL(WL146));
sram_cell_6t_5 inst_cell_146_69 (.BL(BL69),.BLN(BLN69),.WL(WL146));
sram_cell_6t_5 inst_cell_146_70 (.BL(BL70),.BLN(BLN70),.WL(WL146));
sram_cell_6t_5 inst_cell_146_71 (.BL(BL71),.BLN(BLN71),.WL(WL146));
sram_cell_6t_5 inst_cell_146_72 (.BL(BL72),.BLN(BLN72),.WL(WL146));
sram_cell_6t_5 inst_cell_146_73 (.BL(BL73),.BLN(BLN73),.WL(WL146));
sram_cell_6t_5 inst_cell_146_74 (.BL(BL74),.BLN(BLN74),.WL(WL146));
sram_cell_6t_5 inst_cell_146_75 (.BL(BL75),.BLN(BLN75),.WL(WL146));
sram_cell_6t_5 inst_cell_146_76 (.BL(BL76),.BLN(BLN76),.WL(WL146));
sram_cell_6t_5 inst_cell_146_77 (.BL(BL77),.BLN(BLN77),.WL(WL146));
sram_cell_6t_5 inst_cell_146_78 (.BL(BL78),.BLN(BLN78),.WL(WL146));
sram_cell_6t_5 inst_cell_146_79 (.BL(BL79),.BLN(BLN79),.WL(WL146));
sram_cell_6t_5 inst_cell_146_80 (.BL(BL80),.BLN(BLN80),.WL(WL146));
sram_cell_6t_5 inst_cell_146_81 (.BL(BL81),.BLN(BLN81),.WL(WL146));
sram_cell_6t_5 inst_cell_146_82 (.BL(BL82),.BLN(BLN82),.WL(WL146));
sram_cell_6t_5 inst_cell_146_83 (.BL(BL83),.BLN(BLN83),.WL(WL146));
sram_cell_6t_5 inst_cell_146_84 (.BL(BL84),.BLN(BLN84),.WL(WL146));
sram_cell_6t_5 inst_cell_146_85 (.BL(BL85),.BLN(BLN85),.WL(WL146));
sram_cell_6t_5 inst_cell_146_86 (.BL(BL86),.BLN(BLN86),.WL(WL146));
sram_cell_6t_5 inst_cell_146_87 (.BL(BL87),.BLN(BLN87),.WL(WL146));
sram_cell_6t_5 inst_cell_146_88 (.BL(BL88),.BLN(BLN88),.WL(WL146));
sram_cell_6t_5 inst_cell_146_89 (.BL(BL89),.BLN(BLN89),.WL(WL146));
sram_cell_6t_5 inst_cell_146_90 (.BL(BL90),.BLN(BLN90),.WL(WL146));
sram_cell_6t_5 inst_cell_146_91 (.BL(BL91),.BLN(BLN91),.WL(WL146));
sram_cell_6t_5 inst_cell_146_92 (.BL(BL92),.BLN(BLN92),.WL(WL146));
sram_cell_6t_5 inst_cell_146_93 (.BL(BL93),.BLN(BLN93),.WL(WL146));
sram_cell_6t_5 inst_cell_146_94 (.BL(BL94),.BLN(BLN94),.WL(WL146));
sram_cell_6t_5 inst_cell_146_95 (.BL(BL95),.BLN(BLN95),.WL(WL146));
sram_cell_6t_5 inst_cell_146_96 (.BL(BL96),.BLN(BLN96),.WL(WL146));
sram_cell_6t_5 inst_cell_146_97 (.BL(BL97),.BLN(BLN97),.WL(WL146));
sram_cell_6t_5 inst_cell_146_98 (.BL(BL98),.BLN(BLN98),.WL(WL146));
sram_cell_6t_5 inst_cell_146_99 (.BL(BL99),.BLN(BLN99),.WL(WL146));
sram_cell_6t_5 inst_cell_146_100 (.BL(BL100),.BLN(BLN100),.WL(WL146));
sram_cell_6t_5 inst_cell_146_101 (.BL(BL101),.BLN(BLN101),.WL(WL146));
sram_cell_6t_5 inst_cell_146_102 (.BL(BL102),.BLN(BLN102),.WL(WL146));
sram_cell_6t_5 inst_cell_146_103 (.BL(BL103),.BLN(BLN103),.WL(WL146));
sram_cell_6t_5 inst_cell_146_104 (.BL(BL104),.BLN(BLN104),.WL(WL146));
sram_cell_6t_5 inst_cell_146_105 (.BL(BL105),.BLN(BLN105),.WL(WL146));
sram_cell_6t_5 inst_cell_146_106 (.BL(BL106),.BLN(BLN106),.WL(WL146));
sram_cell_6t_5 inst_cell_146_107 (.BL(BL107),.BLN(BLN107),.WL(WL146));
sram_cell_6t_5 inst_cell_146_108 (.BL(BL108),.BLN(BLN108),.WL(WL146));
sram_cell_6t_5 inst_cell_146_109 (.BL(BL109),.BLN(BLN109),.WL(WL146));
sram_cell_6t_5 inst_cell_146_110 (.BL(BL110),.BLN(BLN110),.WL(WL146));
sram_cell_6t_5 inst_cell_146_111 (.BL(BL111),.BLN(BLN111),.WL(WL146));
sram_cell_6t_5 inst_cell_146_112 (.BL(BL112),.BLN(BLN112),.WL(WL146));
sram_cell_6t_5 inst_cell_146_113 (.BL(BL113),.BLN(BLN113),.WL(WL146));
sram_cell_6t_5 inst_cell_146_114 (.BL(BL114),.BLN(BLN114),.WL(WL146));
sram_cell_6t_5 inst_cell_146_115 (.BL(BL115),.BLN(BLN115),.WL(WL146));
sram_cell_6t_5 inst_cell_146_116 (.BL(BL116),.BLN(BLN116),.WL(WL146));
sram_cell_6t_5 inst_cell_146_117 (.BL(BL117),.BLN(BLN117),.WL(WL146));
sram_cell_6t_5 inst_cell_146_118 (.BL(BL118),.BLN(BLN118),.WL(WL146));
sram_cell_6t_5 inst_cell_146_119 (.BL(BL119),.BLN(BLN119),.WL(WL146));
sram_cell_6t_5 inst_cell_146_120 (.BL(BL120),.BLN(BLN120),.WL(WL146));
sram_cell_6t_5 inst_cell_146_121 (.BL(BL121),.BLN(BLN121),.WL(WL146));
sram_cell_6t_5 inst_cell_146_122 (.BL(BL122),.BLN(BLN122),.WL(WL146));
sram_cell_6t_5 inst_cell_146_123 (.BL(BL123),.BLN(BLN123),.WL(WL146));
sram_cell_6t_5 inst_cell_146_124 (.BL(BL124),.BLN(BLN124),.WL(WL146));
sram_cell_6t_5 inst_cell_146_125 (.BL(BL125),.BLN(BLN125),.WL(WL146));
sram_cell_6t_5 inst_cell_146_126 (.BL(BL126),.BLN(BLN126),.WL(WL146));
sram_cell_6t_5 inst_cell_146_127 (.BL(BL127),.BLN(BLN127),.WL(WL146));
sram_cell_6t_5 inst_cell_147_0 (.BL(BL0),.BLN(BLN0),.WL(WL147));
sram_cell_6t_5 inst_cell_147_1 (.BL(BL1),.BLN(BLN1),.WL(WL147));
sram_cell_6t_5 inst_cell_147_2 (.BL(BL2),.BLN(BLN2),.WL(WL147));
sram_cell_6t_5 inst_cell_147_3 (.BL(BL3),.BLN(BLN3),.WL(WL147));
sram_cell_6t_5 inst_cell_147_4 (.BL(BL4),.BLN(BLN4),.WL(WL147));
sram_cell_6t_5 inst_cell_147_5 (.BL(BL5),.BLN(BLN5),.WL(WL147));
sram_cell_6t_5 inst_cell_147_6 (.BL(BL6),.BLN(BLN6),.WL(WL147));
sram_cell_6t_5 inst_cell_147_7 (.BL(BL7),.BLN(BLN7),.WL(WL147));
sram_cell_6t_5 inst_cell_147_8 (.BL(BL8),.BLN(BLN8),.WL(WL147));
sram_cell_6t_5 inst_cell_147_9 (.BL(BL9),.BLN(BLN9),.WL(WL147));
sram_cell_6t_5 inst_cell_147_10 (.BL(BL10),.BLN(BLN10),.WL(WL147));
sram_cell_6t_5 inst_cell_147_11 (.BL(BL11),.BLN(BLN11),.WL(WL147));
sram_cell_6t_5 inst_cell_147_12 (.BL(BL12),.BLN(BLN12),.WL(WL147));
sram_cell_6t_5 inst_cell_147_13 (.BL(BL13),.BLN(BLN13),.WL(WL147));
sram_cell_6t_5 inst_cell_147_14 (.BL(BL14),.BLN(BLN14),.WL(WL147));
sram_cell_6t_5 inst_cell_147_15 (.BL(BL15),.BLN(BLN15),.WL(WL147));
sram_cell_6t_5 inst_cell_147_16 (.BL(BL16),.BLN(BLN16),.WL(WL147));
sram_cell_6t_5 inst_cell_147_17 (.BL(BL17),.BLN(BLN17),.WL(WL147));
sram_cell_6t_5 inst_cell_147_18 (.BL(BL18),.BLN(BLN18),.WL(WL147));
sram_cell_6t_5 inst_cell_147_19 (.BL(BL19),.BLN(BLN19),.WL(WL147));
sram_cell_6t_5 inst_cell_147_20 (.BL(BL20),.BLN(BLN20),.WL(WL147));
sram_cell_6t_5 inst_cell_147_21 (.BL(BL21),.BLN(BLN21),.WL(WL147));
sram_cell_6t_5 inst_cell_147_22 (.BL(BL22),.BLN(BLN22),.WL(WL147));
sram_cell_6t_5 inst_cell_147_23 (.BL(BL23),.BLN(BLN23),.WL(WL147));
sram_cell_6t_5 inst_cell_147_24 (.BL(BL24),.BLN(BLN24),.WL(WL147));
sram_cell_6t_5 inst_cell_147_25 (.BL(BL25),.BLN(BLN25),.WL(WL147));
sram_cell_6t_5 inst_cell_147_26 (.BL(BL26),.BLN(BLN26),.WL(WL147));
sram_cell_6t_5 inst_cell_147_27 (.BL(BL27),.BLN(BLN27),.WL(WL147));
sram_cell_6t_5 inst_cell_147_28 (.BL(BL28),.BLN(BLN28),.WL(WL147));
sram_cell_6t_5 inst_cell_147_29 (.BL(BL29),.BLN(BLN29),.WL(WL147));
sram_cell_6t_5 inst_cell_147_30 (.BL(BL30),.BLN(BLN30),.WL(WL147));
sram_cell_6t_5 inst_cell_147_31 (.BL(BL31),.BLN(BLN31),.WL(WL147));
sram_cell_6t_5 inst_cell_147_32 (.BL(BL32),.BLN(BLN32),.WL(WL147));
sram_cell_6t_5 inst_cell_147_33 (.BL(BL33),.BLN(BLN33),.WL(WL147));
sram_cell_6t_5 inst_cell_147_34 (.BL(BL34),.BLN(BLN34),.WL(WL147));
sram_cell_6t_5 inst_cell_147_35 (.BL(BL35),.BLN(BLN35),.WL(WL147));
sram_cell_6t_5 inst_cell_147_36 (.BL(BL36),.BLN(BLN36),.WL(WL147));
sram_cell_6t_5 inst_cell_147_37 (.BL(BL37),.BLN(BLN37),.WL(WL147));
sram_cell_6t_5 inst_cell_147_38 (.BL(BL38),.BLN(BLN38),.WL(WL147));
sram_cell_6t_5 inst_cell_147_39 (.BL(BL39),.BLN(BLN39),.WL(WL147));
sram_cell_6t_5 inst_cell_147_40 (.BL(BL40),.BLN(BLN40),.WL(WL147));
sram_cell_6t_5 inst_cell_147_41 (.BL(BL41),.BLN(BLN41),.WL(WL147));
sram_cell_6t_5 inst_cell_147_42 (.BL(BL42),.BLN(BLN42),.WL(WL147));
sram_cell_6t_5 inst_cell_147_43 (.BL(BL43),.BLN(BLN43),.WL(WL147));
sram_cell_6t_5 inst_cell_147_44 (.BL(BL44),.BLN(BLN44),.WL(WL147));
sram_cell_6t_5 inst_cell_147_45 (.BL(BL45),.BLN(BLN45),.WL(WL147));
sram_cell_6t_5 inst_cell_147_46 (.BL(BL46),.BLN(BLN46),.WL(WL147));
sram_cell_6t_5 inst_cell_147_47 (.BL(BL47),.BLN(BLN47),.WL(WL147));
sram_cell_6t_5 inst_cell_147_48 (.BL(BL48),.BLN(BLN48),.WL(WL147));
sram_cell_6t_5 inst_cell_147_49 (.BL(BL49),.BLN(BLN49),.WL(WL147));
sram_cell_6t_5 inst_cell_147_50 (.BL(BL50),.BLN(BLN50),.WL(WL147));
sram_cell_6t_5 inst_cell_147_51 (.BL(BL51),.BLN(BLN51),.WL(WL147));
sram_cell_6t_5 inst_cell_147_52 (.BL(BL52),.BLN(BLN52),.WL(WL147));
sram_cell_6t_5 inst_cell_147_53 (.BL(BL53),.BLN(BLN53),.WL(WL147));
sram_cell_6t_5 inst_cell_147_54 (.BL(BL54),.BLN(BLN54),.WL(WL147));
sram_cell_6t_5 inst_cell_147_55 (.BL(BL55),.BLN(BLN55),.WL(WL147));
sram_cell_6t_5 inst_cell_147_56 (.BL(BL56),.BLN(BLN56),.WL(WL147));
sram_cell_6t_5 inst_cell_147_57 (.BL(BL57),.BLN(BLN57),.WL(WL147));
sram_cell_6t_5 inst_cell_147_58 (.BL(BL58),.BLN(BLN58),.WL(WL147));
sram_cell_6t_5 inst_cell_147_59 (.BL(BL59),.BLN(BLN59),.WL(WL147));
sram_cell_6t_5 inst_cell_147_60 (.BL(BL60),.BLN(BLN60),.WL(WL147));
sram_cell_6t_5 inst_cell_147_61 (.BL(BL61),.BLN(BLN61),.WL(WL147));
sram_cell_6t_5 inst_cell_147_62 (.BL(BL62),.BLN(BLN62),.WL(WL147));
sram_cell_6t_5 inst_cell_147_63 (.BL(BL63),.BLN(BLN63),.WL(WL147));
sram_cell_6t_5 inst_cell_147_64 (.BL(BL64),.BLN(BLN64),.WL(WL147));
sram_cell_6t_5 inst_cell_147_65 (.BL(BL65),.BLN(BLN65),.WL(WL147));
sram_cell_6t_5 inst_cell_147_66 (.BL(BL66),.BLN(BLN66),.WL(WL147));
sram_cell_6t_5 inst_cell_147_67 (.BL(BL67),.BLN(BLN67),.WL(WL147));
sram_cell_6t_5 inst_cell_147_68 (.BL(BL68),.BLN(BLN68),.WL(WL147));
sram_cell_6t_5 inst_cell_147_69 (.BL(BL69),.BLN(BLN69),.WL(WL147));
sram_cell_6t_5 inst_cell_147_70 (.BL(BL70),.BLN(BLN70),.WL(WL147));
sram_cell_6t_5 inst_cell_147_71 (.BL(BL71),.BLN(BLN71),.WL(WL147));
sram_cell_6t_5 inst_cell_147_72 (.BL(BL72),.BLN(BLN72),.WL(WL147));
sram_cell_6t_5 inst_cell_147_73 (.BL(BL73),.BLN(BLN73),.WL(WL147));
sram_cell_6t_5 inst_cell_147_74 (.BL(BL74),.BLN(BLN74),.WL(WL147));
sram_cell_6t_5 inst_cell_147_75 (.BL(BL75),.BLN(BLN75),.WL(WL147));
sram_cell_6t_5 inst_cell_147_76 (.BL(BL76),.BLN(BLN76),.WL(WL147));
sram_cell_6t_5 inst_cell_147_77 (.BL(BL77),.BLN(BLN77),.WL(WL147));
sram_cell_6t_5 inst_cell_147_78 (.BL(BL78),.BLN(BLN78),.WL(WL147));
sram_cell_6t_5 inst_cell_147_79 (.BL(BL79),.BLN(BLN79),.WL(WL147));
sram_cell_6t_5 inst_cell_147_80 (.BL(BL80),.BLN(BLN80),.WL(WL147));
sram_cell_6t_5 inst_cell_147_81 (.BL(BL81),.BLN(BLN81),.WL(WL147));
sram_cell_6t_5 inst_cell_147_82 (.BL(BL82),.BLN(BLN82),.WL(WL147));
sram_cell_6t_5 inst_cell_147_83 (.BL(BL83),.BLN(BLN83),.WL(WL147));
sram_cell_6t_5 inst_cell_147_84 (.BL(BL84),.BLN(BLN84),.WL(WL147));
sram_cell_6t_5 inst_cell_147_85 (.BL(BL85),.BLN(BLN85),.WL(WL147));
sram_cell_6t_5 inst_cell_147_86 (.BL(BL86),.BLN(BLN86),.WL(WL147));
sram_cell_6t_5 inst_cell_147_87 (.BL(BL87),.BLN(BLN87),.WL(WL147));
sram_cell_6t_5 inst_cell_147_88 (.BL(BL88),.BLN(BLN88),.WL(WL147));
sram_cell_6t_5 inst_cell_147_89 (.BL(BL89),.BLN(BLN89),.WL(WL147));
sram_cell_6t_5 inst_cell_147_90 (.BL(BL90),.BLN(BLN90),.WL(WL147));
sram_cell_6t_5 inst_cell_147_91 (.BL(BL91),.BLN(BLN91),.WL(WL147));
sram_cell_6t_5 inst_cell_147_92 (.BL(BL92),.BLN(BLN92),.WL(WL147));
sram_cell_6t_5 inst_cell_147_93 (.BL(BL93),.BLN(BLN93),.WL(WL147));
sram_cell_6t_5 inst_cell_147_94 (.BL(BL94),.BLN(BLN94),.WL(WL147));
sram_cell_6t_5 inst_cell_147_95 (.BL(BL95),.BLN(BLN95),.WL(WL147));
sram_cell_6t_5 inst_cell_147_96 (.BL(BL96),.BLN(BLN96),.WL(WL147));
sram_cell_6t_5 inst_cell_147_97 (.BL(BL97),.BLN(BLN97),.WL(WL147));
sram_cell_6t_5 inst_cell_147_98 (.BL(BL98),.BLN(BLN98),.WL(WL147));
sram_cell_6t_5 inst_cell_147_99 (.BL(BL99),.BLN(BLN99),.WL(WL147));
sram_cell_6t_5 inst_cell_147_100 (.BL(BL100),.BLN(BLN100),.WL(WL147));
sram_cell_6t_5 inst_cell_147_101 (.BL(BL101),.BLN(BLN101),.WL(WL147));
sram_cell_6t_5 inst_cell_147_102 (.BL(BL102),.BLN(BLN102),.WL(WL147));
sram_cell_6t_5 inst_cell_147_103 (.BL(BL103),.BLN(BLN103),.WL(WL147));
sram_cell_6t_5 inst_cell_147_104 (.BL(BL104),.BLN(BLN104),.WL(WL147));
sram_cell_6t_5 inst_cell_147_105 (.BL(BL105),.BLN(BLN105),.WL(WL147));
sram_cell_6t_5 inst_cell_147_106 (.BL(BL106),.BLN(BLN106),.WL(WL147));
sram_cell_6t_5 inst_cell_147_107 (.BL(BL107),.BLN(BLN107),.WL(WL147));
sram_cell_6t_5 inst_cell_147_108 (.BL(BL108),.BLN(BLN108),.WL(WL147));
sram_cell_6t_5 inst_cell_147_109 (.BL(BL109),.BLN(BLN109),.WL(WL147));
sram_cell_6t_5 inst_cell_147_110 (.BL(BL110),.BLN(BLN110),.WL(WL147));
sram_cell_6t_5 inst_cell_147_111 (.BL(BL111),.BLN(BLN111),.WL(WL147));
sram_cell_6t_5 inst_cell_147_112 (.BL(BL112),.BLN(BLN112),.WL(WL147));
sram_cell_6t_5 inst_cell_147_113 (.BL(BL113),.BLN(BLN113),.WL(WL147));
sram_cell_6t_5 inst_cell_147_114 (.BL(BL114),.BLN(BLN114),.WL(WL147));
sram_cell_6t_5 inst_cell_147_115 (.BL(BL115),.BLN(BLN115),.WL(WL147));
sram_cell_6t_5 inst_cell_147_116 (.BL(BL116),.BLN(BLN116),.WL(WL147));
sram_cell_6t_5 inst_cell_147_117 (.BL(BL117),.BLN(BLN117),.WL(WL147));
sram_cell_6t_5 inst_cell_147_118 (.BL(BL118),.BLN(BLN118),.WL(WL147));
sram_cell_6t_5 inst_cell_147_119 (.BL(BL119),.BLN(BLN119),.WL(WL147));
sram_cell_6t_5 inst_cell_147_120 (.BL(BL120),.BLN(BLN120),.WL(WL147));
sram_cell_6t_5 inst_cell_147_121 (.BL(BL121),.BLN(BLN121),.WL(WL147));
sram_cell_6t_5 inst_cell_147_122 (.BL(BL122),.BLN(BLN122),.WL(WL147));
sram_cell_6t_5 inst_cell_147_123 (.BL(BL123),.BLN(BLN123),.WL(WL147));
sram_cell_6t_5 inst_cell_147_124 (.BL(BL124),.BLN(BLN124),.WL(WL147));
sram_cell_6t_5 inst_cell_147_125 (.BL(BL125),.BLN(BLN125),.WL(WL147));
sram_cell_6t_5 inst_cell_147_126 (.BL(BL126),.BLN(BLN126),.WL(WL147));
sram_cell_6t_5 inst_cell_147_127 (.BL(BL127),.BLN(BLN127),.WL(WL147));
sram_cell_6t_5 inst_cell_148_0 (.BL(BL0),.BLN(BLN0),.WL(WL148));
sram_cell_6t_5 inst_cell_148_1 (.BL(BL1),.BLN(BLN1),.WL(WL148));
sram_cell_6t_5 inst_cell_148_2 (.BL(BL2),.BLN(BLN2),.WL(WL148));
sram_cell_6t_5 inst_cell_148_3 (.BL(BL3),.BLN(BLN3),.WL(WL148));
sram_cell_6t_5 inst_cell_148_4 (.BL(BL4),.BLN(BLN4),.WL(WL148));
sram_cell_6t_5 inst_cell_148_5 (.BL(BL5),.BLN(BLN5),.WL(WL148));
sram_cell_6t_5 inst_cell_148_6 (.BL(BL6),.BLN(BLN6),.WL(WL148));
sram_cell_6t_5 inst_cell_148_7 (.BL(BL7),.BLN(BLN7),.WL(WL148));
sram_cell_6t_5 inst_cell_148_8 (.BL(BL8),.BLN(BLN8),.WL(WL148));
sram_cell_6t_5 inst_cell_148_9 (.BL(BL9),.BLN(BLN9),.WL(WL148));
sram_cell_6t_5 inst_cell_148_10 (.BL(BL10),.BLN(BLN10),.WL(WL148));
sram_cell_6t_5 inst_cell_148_11 (.BL(BL11),.BLN(BLN11),.WL(WL148));
sram_cell_6t_5 inst_cell_148_12 (.BL(BL12),.BLN(BLN12),.WL(WL148));
sram_cell_6t_5 inst_cell_148_13 (.BL(BL13),.BLN(BLN13),.WL(WL148));
sram_cell_6t_5 inst_cell_148_14 (.BL(BL14),.BLN(BLN14),.WL(WL148));
sram_cell_6t_5 inst_cell_148_15 (.BL(BL15),.BLN(BLN15),.WL(WL148));
sram_cell_6t_5 inst_cell_148_16 (.BL(BL16),.BLN(BLN16),.WL(WL148));
sram_cell_6t_5 inst_cell_148_17 (.BL(BL17),.BLN(BLN17),.WL(WL148));
sram_cell_6t_5 inst_cell_148_18 (.BL(BL18),.BLN(BLN18),.WL(WL148));
sram_cell_6t_5 inst_cell_148_19 (.BL(BL19),.BLN(BLN19),.WL(WL148));
sram_cell_6t_5 inst_cell_148_20 (.BL(BL20),.BLN(BLN20),.WL(WL148));
sram_cell_6t_5 inst_cell_148_21 (.BL(BL21),.BLN(BLN21),.WL(WL148));
sram_cell_6t_5 inst_cell_148_22 (.BL(BL22),.BLN(BLN22),.WL(WL148));
sram_cell_6t_5 inst_cell_148_23 (.BL(BL23),.BLN(BLN23),.WL(WL148));
sram_cell_6t_5 inst_cell_148_24 (.BL(BL24),.BLN(BLN24),.WL(WL148));
sram_cell_6t_5 inst_cell_148_25 (.BL(BL25),.BLN(BLN25),.WL(WL148));
sram_cell_6t_5 inst_cell_148_26 (.BL(BL26),.BLN(BLN26),.WL(WL148));
sram_cell_6t_5 inst_cell_148_27 (.BL(BL27),.BLN(BLN27),.WL(WL148));
sram_cell_6t_5 inst_cell_148_28 (.BL(BL28),.BLN(BLN28),.WL(WL148));
sram_cell_6t_5 inst_cell_148_29 (.BL(BL29),.BLN(BLN29),.WL(WL148));
sram_cell_6t_5 inst_cell_148_30 (.BL(BL30),.BLN(BLN30),.WL(WL148));
sram_cell_6t_5 inst_cell_148_31 (.BL(BL31),.BLN(BLN31),.WL(WL148));
sram_cell_6t_5 inst_cell_148_32 (.BL(BL32),.BLN(BLN32),.WL(WL148));
sram_cell_6t_5 inst_cell_148_33 (.BL(BL33),.BLN(BLN33),.WL(WL148));
sram_cell_6t_5 inst_cell_148_34 (.BL(BL34),.BLN(BLN34),.WL(WL148));
sram_cell_6t_5 inst_cell_148_35 (.BL(BL35),.BLN(BLN35),.WL(WL148));
sram_cell_6t_5 inst_cell_148_36 (.BL(BL36),.BLN(BLN36),.WL(WL148));
sram_cell_6t_5 inst_cell_148_37 (.BL(BL37),.BLN(BLN37),.WL(WL148));
sram_cell_6t_5 inst_cell_148_38 (.BL(BL38),.BLN(BLN38),.WL(WL148));
sram_cell_6t_5 inst_cell_148_39 (.BL(BL39),.BLN(BLN39),.WL(WL148));
sram_cell_6t_5 inst_cell_148_40 (.BL(BL40),.BLN(BLN40),.WL(WL148));
sram_cell_6t_5 inst_cell_148_41 (.BL(BL41),.BLN(BLN41),.WL(WL148));
sram_cell_6t_5 inst_cell_148_42 (.BL(BL42),.BLN(BLN42),.WL(WL148));
sram_cell_6t_5 inst_cell_148_43 (.BL(BL43),.BLN(BLN43),.WL(WL148));
sram_cell_6t_5 inst_cell_148_44 (.BL(BL44),.BLN(BLN44),.WL(WL148));
sram_cell_6t_5 inst_cell_148_45 (.BL(BL45),.BLN(BLN45),.WL(WL148));
sram_cell_6t_5 inst_cell_148_46 (.BL(BL46),.BLN(BLN46),.WL(WL148));
sram_cell_6t_5 inst_cell_148_47 (.BL(BL47),.BLN(BLN47),.WL(WL148));
sram_cell_6t_5 inst_cell_148_48 (.BL(BL48),.BLN(BLN48),.WL(WL148));
sram_cell_6t_5 inst_cell_148_49 (.BL(BL49),.BLN(BLN49),.WL(WL148));
sram_cell_6t_5 inst_cell_148_50 (.BL(BL50),.BLN(BLN50),.WL(WL148));
sram_cell_6t_5 inst_cell_148_51 (.BL(BL51),.BLN(BLN51),.WL(WL148));
sram_cell_6t_5 inst_cell_148_52 (.BL(BL52),.BLN(BLN52),.WL(WL148));
sram_cell_6t_5 inst_cell_148_53 (.BL(BL53),.BLN(BLN53),.WL(WL148));
sram_cell_6t_5 inst_cell_148_54 (.BL(BL54),.BLN(BLN54),.WL(WL148));
sram_cell_6t_5 inst_cell_148_55 (.BL(BL55),.BLN(BLN55),.WL(WL148));
sram_cell_6t_5 inst_cell_148_56 (.BL(BL56),.BLN(BLN56),.WL(WL148));
sram_cell_6t_5 inst_cell_148_57 (.BL(BL57),.BLN(BLN57),.WL(WL148));
sram_cell_6t_5 inst_cell_148_58 (.BL(BL58),.BLN(BLN58),.WL(WL148));
sram_cell_6t_5 inst_cell_148_59 (.BL(BL59),.BLN(BLN59),.WL(WL148));
sram_cell_6t_5 inst_cell_148_60 (.BL(BL60),.BLN(BLN60),.WL(WL148));
sram_cell_6t_5 inst_cell_148_61 (.BL(BL61),.BLN(BLN61),.WL(WL148));
sram_cell_6t_5 inst_cell_148_62 (.BL(BL62),.BLN(BLN62),.WL(WL148));
sram_cell_6t_5 inst_cell_148_63 (.BL(BL63),.BLN(BLN63),.WL(WL148));
sram_cell_6t_5 inst_cell_148_64 (.BL(BL64),.BLN(BLN64),.WL(WL148));
sram_cell_6t_5 inst_cell_148_65 (.BL(BL65),.BLN(BLN65),.WL(WL148));
sram_cell_6t_5 inst_cell_148_66 (.BL(BL66),.BLN(BLN66),.WL(WL148));
sram_cell_6t_5 inst_cell_148_67 (.BL(BL67),.BLN(BLN67),.WL(WL148));
sram_cell_6t_5 inst_cell_148_68 (.BL(BL68),.BLN(BLN68),.WL(WL148));
sram_cell_6t_5 inst_cell_148_69 (.BL(BL69),.BLN(BLN69),.WL(WL148));
sram_cell_6t_5 inst_cell_148_70 (.BL(BL70),.BLN(BLN70),.WL(WL148));
sram_cell_6t_5 inst_cell_148_71 (.BL(BL71),.BLN(BLN71),.WL(WL148));
sram_cell_6t_5 inst_cell_148_72 (.BL(BL72),.BLN(BLN72),.WL(WL148));
sram_cell_6t_5 inst_cell_148_73 (.BL(BL73),.BLN(BLN73),.WL(WL148));
sram_cell_6t_5 inst_cell_148_74 (.BL(BL74),.BLN(BLN74),.WL(WL148));
sram_cell_6t_5 inst_cell_148_75 (.BL(BL75),.BLN(BLN75),.WL(WL148));
sram_cell_6t_5 inst_cell_148_76 (.BL(BL76),.BLN(BLN76),.WL(WL148));
sram_cell_6t_5 inst_cell_148_77 (.BL(BL77),.BLN(BLN77),.WL(WL148));
sram_cell_6t_5 inst_cell_148_78 (.BL(BL78),.BLN(BLN78),.WL(WL148));
sram_cell_6t_5 inst_cell_148_79 (.BL(BL79),.BLN(BLN79),.WL(WL148));
sram_cell_6t_5 inst_cell_148_80 (.BL(BL80),.BLN(BLN80),.WL(WL148));
sram_cell_6t_5 inst_cell_148_81 (.BL(BL81),.BLN(BLN81),.WL(WL148));
sram_cell_6t_5 inst_cell_148_82 (.BL(BL82),.BLN(BLN82),.WL(WL148));
sram_cell_6t_5 inst_cell_148_83 (.BL(BL83),.BLN(BLN83),.WL(WL148));
sram_cell_6t_5 inst_cell_148_84 (.BL(BL84),.BLN(BLN84),.WL(WL148));
sram_cell_6t_5 inst_cell_148_85 (.BL(BL85),.BLN(BLN85),.WL(WL148));
sram_cell_6t_5 inst_cell_148_86 (.BL(BL86),.BLN(BLN86),.WL(WL148));
sram_cell_6t_5 inst_cell_148_87 (.BL(BL87),.BLN(BLN87),.WL(WL148));
sram_cell_6t_5 inst_cell_148_88 (.BL(BL88),.BLN(BLN88),.WL(WL148));
sram_cell_6t_5 inst_cell_148_89 (.BL(BL89),.BLN(BLN89),.WL(WL148));
sram_cell_6t_5 inst_cell_148_90 (.BL(BL90),.BLN(BLN90),.WL(WL148));
sram_cell_6t_5 inst_cell_148_91 (.BL(BL91),.BLN(BLN91),.WL(WL148));
sram_cell_6t_5 inst_cell_148_92 (.BL(BL92),.BLN(BLN92),.WL(WL148));
sram_cell_6t_5 inst_cell_148_93 (.BL(BL93),.BLN(BLN93),.WL(WL148));
sram_cell_6t_5 inst_cell_148_94 (.BL(BL94),.BLN(BLN94),.WL(WL148));
sram_cell_6t_5 inst_cell_148_95 (.BL(BL95),.BLN(BLN95),.WL(WL148));
sram_cell_6t_5 inst_cell_148_96 (.BL(BL96),.BLN(BLN96),.WL(WL148));
sram_cell_6t_5 inst_cell_148_97 (.BL(BL97),.BLN(BLN97),.WL(WL148));
sram_cell_6t_5 inst_cell_148_98 (.BL(BL98),.BLN(BLN98),.WL(WL148));
sram_cell_6t_5 inst_cell_148_99 (.BL(BL99),.BLN(BLN99),.WL(WL148));
sram_cell_6t_5 inst_cell_148_100 (.BL(BL100),.BLN(BLN100),.WL(WL148));
sram_cell_6t_5 inst_cell_148_101 (.BL(BL101),.BLN(BLN101),.WL(WL148));
sram_cell_6t_5 inst_cell_148_102 (.BL(BL102),.BLN(BLN102),.WL(WL148));
sram_cell_6t_5 inst_cell_148_103 (.BL(BL103),.BLN(BLN103),.WL(WL148));
sram_cell_6t_5 inst_cell_148_104 (.BL(BL104),.BLN(BLN104),.WL(WL148));
sram_cell_6t_5 inst_cell_148_105 (.BL(BL105),.BLN(BLN105),.WL(WL148));
sram_cell_6t_5 inst_cell_148_106 (.BL(BL106),.BLN(BLN106),.WL(WL148));
sram_cell_6t_5 inst_cell_148_107 (.BL(BL107),.BLN(BLN107),.WL(WL148));
sram_cell_6t_5 inst_cell_148_108 (.BL(BL108),.BLN(BLN108),.WL(WL148));
sram_cell_6t_5 inst_cell_148_109 (.BL(BL109),.BLN(BLN109),.WL(WL148));
sram_cell_6t_5 inst_cell_148_110 (.BL(BL110),.BLN(BLN110),.WL(WL148));
sram_cell_6t_5 inst_cell_148_111 (.BL(BL111),.BLN(BLN111),.WL(WL148));
sram_cell_6t_5 inst_cell_148_112 (.BL(BL112),.BLN(BLN112),.WL(WL148));
sram_cell_6t_5 inst_cell_148_113 (.BL(BL113),.BLN(BLN113),.WL(WL148));
sram_cell_6t_5 inst_cell_148_114 (.BL(BL114),.BLN(BLN114),.WL(WL148));
sram_cell_6t_5 inst_cell_148_115 (.BL(BL115),.BLN(BLN115),.WL(WL148));
sram_cell_6t_5 inst_cell_148_116 (.BL(BL116),.BLN(BLN116),.WL(WL148));
sram_cell_6t_5 inst_cell_148_117 (.BL(BL117),.BLN(BLN117),.WL(WL148));
sram_cell_6t_5 inst_cell_148_118 (.BL(BL118),.BLN(BLN118),.WL(WL148));
sram_cell_6t_5 inst_cell_148_119 (.BL(BL119),.BLN(BLN119),.WL(WL148));
sram_cell_6t_5 inst_cell_148_120 (.BL(BL120),.BLN(BLN120),.WL(WL148));
sram_cell_6t_5 inst_cell_148_121 (.BL(BL121),.BLN(BLN121),.WL(WL148));
sram_cell_6t_5 inst_cell_148_122 (.BL(BL122),.BLN(BLN122),.WL(WL148));
sram_cell_6t_5 inst_cell_148_123 (.BL(BL123),.BLN(BLN123),.WL(WL148));
sram_cell_6t_5 inst_cell_148_124 (.BL(BL124),.BLN(BLN124),.WL(WL148));
sram_cell_6t_5 inst_cell_148_125 (.BL(BL125),.BLN(BLN125),.WL(WL148));
sram_cell_6t_5 inst_cell_148_126 (.BL(BL126),.BLN(BLN126),.WL(WL148));
sram_cell_6t_5 inst_cell_148_127 (.BL(BL127),.BLN(BLN127),.WL(WL148));
sram_cell_6t_5 inst_cell_149_0 (.BL(BL0),.BLN(BLN0),.WL(WL149));
sram_cell_6t_5 inst_cell_149_1 (.BL(BL1),.BLN(BLN1),.WL(WL149));
sram_cell_6t_5 inst_cell_149_2 (.BL(BL2),.BLN(BLN2),.WL(WL149));
sram_cell_6t_5 inst_cell_149_3 (.BL(BL3),.BLN(BLN3),.WL(WL149));
sram_cell_6t_5 inst_cell_149_4 (.BL(BL4),.BLN(BLN4),.WL(WL149));
sram_cell_6t_5 inst_cell_149_5 (.BL(BL5),.BLN(BLN5),.WL(WL149));
sram_cell_6t_5 inst_cell_149_6 (.BL(BL6),.BLN(BLN6),.WL(WL149));
sram_cell_6t_5 inst_cell_149_7 (.BL(BL7),.BLN(BLN7),.WL(WL149));
sram_cell_6t_5 inst_cell_149_8 (.BL(BL8),.BLN(BLN8),.WL(WL149));
sram_cell_6t_5 inst_cell_149_9 (.BL(BL9),.BLN(BLN9),.WL(WL149));
sram_cell_6t_5 inst_cell_149_10 (.BL(BL10),.BLN(BLN10),.WL(WL149));
sram_cell_6t_5 inst_cell_149_11 (.BL(BL11),.BLN(BLN11),.WL(WL149));
sram_cell_6t_5 inst_cell_149_12 (.BL(BL12),.BLN(BLN12),.WL(WL149));
sram_cell_6t_5 inst_cell_149_13 (.BL(BL13),.BLN(BLN13),.WL(WL149));
sram_cell_6t_5 inst_cell_149_14 (.BL(BL14),.BLN(BLN14),.WL(WL149));
sram_cell_6t_5 inst_cell_149_15 (.BL(BL15),.BLN(BLN15),.WL(WL149));
sram_cell_6t_5 inst_cell_149_16 (.BL(BL16),.BLN(BLN16),.WL(WL149));
sram_cell_6t_5 inst_cell_149_17 (.BL(BL17),.BLN(BLN17),.WL(WL149));
sram_cell_6t_5 inst_cell_149_18 (.BL(BL18),.BLN(BLN18),.WL(WL149));
sram_cell_6t_5 inst_cell_149_19 (.BL(BL19),.BLN(BLN19),.WL(WL149));
sram_cell_6t_5 inst_cell_149_20 (.BL(BL20),.BLN(BLN20),.WL(WL149));
sram_cell_6t_5 inst_cell_149_21 (.BL(BL21),.BLN(BLN21),.WL(WL149));
sram_cell_6t_5 inst_cell_149_22 (.BL(BL22),.BLN(BLN22),.WL(WL149));
sram_cell_6t_5 inst_cell_149_23 (.BL(BL23),.BLN(BLN23),.WL(WL149));
sram_cell_6t_5 inst_cell_149_24 (.BL(BL24),.BLN(BLN24),.WL(WL149));
sram_cell_6t_5 inst_cell_149_25 (.BL(BL25),.BLN(BLN25),.WL(WL149));
sram_cell_6t_5 inst_cell_149_26 (.BL(BL26),.BLN(BLN26),.WL(WL149));
sram_cell_6t_5 inst_cell_149_27 (.BL(BL27),.BLN(BLN27),.WL(WL149));
sram_cell_6t_5 inst_cell_149_28 (.BL(BL28),.BLN(BLN28),.WL(WL149));
sram_cell_6t_5 inst_cell_149_29 (.BL(BL29),.BLN(BLN29),.WL(WL149));
sram_cell_6t_5 inst_cell_149_30 (.BL(BL30),.BLN(BLN30),.WL(WL149));
sram_cell_6t_5 inst_cell_149_31 (.BL(BL31),.BLN(BLN31),.WL(WL149));
sram_cell_6t_5 inst_cell_149_32 (.BL(BL32),.BLN(BLN32),.WL(WL149));
sram_cell_6t_5 inst_cell_149_33 (.BL(BL33),.BLN(BLN33),.WL(WL149));
sram_cell_6t_5 inst_cell_149_34 (.BL(BL34),.BLN(BLN34),.WL(WL149));
sram_cell_6t_5 inst_cell_149_35 (.BL(BL35),.BLN(BLN35),.WL(WL149));
sram_cell_6t_5 inst_cell_149_36 (.BL(BL36),.BLN(BLN36),.WL(WL149));
sram_cell_6t_5 inst_cell_149_37 (.BL(BL37),.BLN(BLN37),.WL(WL149));
sram_cell_6t_5 inst_cell_149_38 (.BL(BL38),.BLN(BLN38),.WL(WL149));
sram_cell_6t_5 inst_cell_149_39 (.BL(BL39),.BLN(BLN39),.WL(WL149));
sram_cell_6t_5 inst_cell_149_40 (.BL(BL40),.BLN(BLN40),.WL(WL149));
sram_cell_6t_5 inst_cell_149_41 (.BL(BL41),.BLN(BLN41),.WL(WL149));
sram_cell_6t_5 inst_cell_149_42 (.BL(BL42),.BLN(BLN42),.WL(WL149));
sram_cell_6t_5 inst_cell_149_43 (.BL(BL43),.BLN(BLN43),.WL(WL149));
sram_cell_6t_5 inst_cell_149_44 (.BL(BL44),.BLN(BLN44),.WL(WL149));
sram_cell_6t_5 inst_cell_149_45 (.BL(BL45),.BLN(BLN45),.WL(WL149));
sram_cell_6t_5 inst_cell_149_46 (.BL(BL46),.BLN(BLN46),.WL(WL149));
sram_cell_6t_5 inst_cell_149_47 (.BL(BL47),.BLN(BLN47),.WL(WL149));
sram_cell_6t_5 inst_cell_149_48 (.BL(BL48),.BLN(BLN48),.WL(WL149));
sram_cell_6t_5 inst_cell_149_49 (.BL(BL49),.BLN(BLN49),.WL(WL149));
sram_cell_6t_5 inst_cell_149_50 (.BL(BL50),.BLN(BLN50),.WL(WL149));
sram_cell_6t_5 inst_cell_149_51 (.BL(BL51),.BLN(BLN51),.WL(WL149));
sram_cell_6t_5 inst_cell_149_52 (.BL(BL52),.BLN(BLN52),.WL(WL149));
sram_cell_6t_5 inst_cell_149_53 (.BL(BL53),.BLN(BLN53),.WL(WL149));
sram_cell_6t_5 inst_cell_149_54 (.BL(BL54),.BLN(BLN54),.WL(WL149));
sram_cell_6t_5 inst_cell_149_55 (.BL(BL55),.BLN(BLN55),.WL(WL149));
sram_cell_6t_5 inst_cell_149_56 (.BL(BL56),.BLN(BLN56),.WL(WL149));
sram_cell_6t_5 inst_cell_149_57 (.BL(BL57),.BLN(BLN57),.WL(WL149));
sram_cell_6t_5 inst_cell_149_58 (.BL(BL58),.BLN(BLN58),.WL(WL149));
sram_cell_6t_5 inst_cell_149_59 (.BL(BL59),.BLN(BLN59),.WL(WL149));
sram_cell_6t_5 inst_cell_149_60 (.BL(BL60),.BLN(BLN60),.WL(WL149));
sram_cell_6t_5 inst_cell_149_61 (.BL(BL61),.BLN(BLN61),.WL(WL149));
sram_cell_6t_5 inst_cell_149_62 (.BL(BL62),.BLN(BLN62),.WL(WL149));
sram_cell_6t_5 inst_cell_149_63 (.BL(BL63),.BLN(BLN63),.WL(WL149));
sram_cell_6t_5 inst_cell_149_64 (.BL(BL64),.BLN(BLN64),.WL(WL149));
sram_cell_6t_5 inst_cell_149_65 (.BL(BL65),.BLN(BLN65),.WL(WL149));
sram_cell_6t_5 inst_cell_149_66 (.BL(BL66),.BLN(BLN66),.WL(WL149));
sram_cell_6t_5 inst_cell_149_67 (.BL(BL67),.BLN(BLN67),.WL(WL149));
sram_cell_6t_5 inst_cell_149_68 (.BL(BL68),.BLN(BLN68),.WL(WL149));
sram_cell_6t_5 inst_cell_149_69 (.BL(BL69),.BLN(BLN69),.WL(WL149));
sram_cell_6t_5 inst_cell_149_70 (.BL(BL70),.BLN(BLN70),.WL(WL149));
sram_cell_6t_5 inst_cell_149_71 (.BL(BL71),.BLN(BLN71),.WL(WL149));
sram_cell_6t_5 inst_cell_149_72 (.BL(BL72),.BLN(BLN72),.WL(WL149));
sram_cell_6t_5 inst_cell_149_73 (.BL(BL73),.BLN(BLN73),.WL(WL149));
sram_cell_6t_5 inst_cell_149_74 (.BL(BL74),.BLN(BLN74),.WL(WL149));
sram_cell_6t_5 inst_cell_149_75 (.BL(BL75),.BLN(BLN75),.WL(WL149));
sram_cell_6t_5 inst_cell_149_76 (.BL(BL76),.BLN(BLN76),.WL(WL149));
sram_cell_6t_5 inst_cell_149_77 (.BL(BL77),.BLN(BLN77),.WL(WL149));
sram_cell_6t_5 inst_cell_149_78 (.BL(BL78),.BLN(BLN78),.WL(WL149));
sram_cell_6t_5 inst_cell_149_79 (.BL(BL79),.BLN(BLN79),.WL(WL149));
sram_cell_6t_5 inst_cell_149_80 (.BL(BL80),.BLN(BLN80),.WL(WL149));
sram_cell_6t_5 inst_cell_149_81 (.BL(BL81),.BLN(BLN81),.WL(WL149));
sram_cell_6t_5 inst_cell_149_82 (.BL(BL82),.BLN(BLN82),.WL(WL149));
sram_cell_6t_5 inst_cell_149_83 (.BL(BL83),.BLN(BLN83),.WL(WL149));
sram_cell_6t_5 inst_cell_149_84 (.BL(BL84),.BLN(BLN84),.WL(WL149));
sram_cell_6t_5 inst_cell_149_85 (.BL(BL85),.BLN(BLN85),.WL(WL149));
sram_cell_6t_5 inst_cell_149_86 (.BL(BL86),.BLN(BLN86),.WL(WL149));
sram_cell_6t_5 inst_cell_149_87 (.BL(BL87),.BLN(BLN87),.WL(WL149));
sram_cell_6t_5 inst_cell_149_88 (.BL(BL88),.BLN(BLN88),.WL(WL149));
sram_cell_6t_5 inst_cell_149_89 (.BL(BL89),.BLN(BLN89),.WL(WL149));
sram_cell_6t_5 inst_cell_149_90 (.BL(BL90),.BLN(BLN90),.WL(WL149));
sram_cell_6t_5 inst_cell_149_91 (.BL(BL91),.BLN(BLN91),.WL(WL149));
sram_cell_6t_5 inst_cell_149_92 (.BL(BL92),.BLN(BLN92),.WL(WL149));
sram_cell_6t_5 inst_cell_149_93 (.BL(BL93),.BLN(BLN93),.WL(WL149));
sram_cell_6t_5 inst_cell_149_94 (.BL(BL94),.BLN(BLN94),.WL(WL149));
sram_cell_6t_5 inst_cell_149_95 (.BL(BL95),.BLN(BLN95),.WL(WL149));
sram_cell_6t_5 inst_cell_149_96 (.BL(BL96),.BLN(BLN96),.WL(WL149));
sram_cell_6t_5 inst_cell_149_97 (.BL(BL97),.BLN(BLN97),.WL(WL149));
sram_cell_6t_5 inst_cell_149_98 (.BL(BL98),.BLN(BLN98),.WL(WL149));
sram_cell_6t_5 inst_cell_149_99 (.BL(BL99),.BLN(BLN99),.WL(WL149));
sram_cell_6t_5 inst_cell_149_100 (.BL(BL100),.BLN(BLN100),.WL(WL149));
sram_cell_6t_5 inst_cell_149_101 (.BL(BL101),.BLN(BLN101),.WL(WL149));
sram_cell_6t_5 inst_cell_149_102 (.BL(BL102),.BLN(BLN102),.WL(WL149));
sram_cell_6t_5 inst_cell_149_103 (.BL(BL103),.BLN(BLN103),.WL(WL149));
sram_cell_6t_5 inst_cell_149_104 (.BL(BL104),.BLN(BLN104),.WL(WL149));
sram_cell_6t_5 inst_cell_149_105 (.BL(BL105),.BLN(BLN105),.WL(WL149));
sram_cell_6t_5 inst_cell_149_106 (.BL(BL106),.BLN(BLN106),.WL(WL149));
sram_cell_6t_5 inst_cell_149_107 (.BL(BL107),.BLN(BLN107),.WL(WL149));
sram_cell_6t_5 inst_cell_149_108 (.BL(BL108),.BLN(BLN108),.WL(WL149));
sram_cell_6t_5 inst_cell_149_109 (.BL(BL109),.BLN(BLN109),.WL(WL149));
sram_cell_6t_5 inst_cell_149_110 (.BL(BL110),.BLN(BLN110),.WL(WL149));
sram_cell_6t_5 inst_cell_149_111 (.BL(BL111),.BLN(BLN111),.WL(WL149));
sram_cell_6t_5 inst_cell_149_112 (.BL(BL112),.BLN(BLN112),.WL(WL149));
sram_cell_6t_5 inst_cell_149_113 (.BL(BL113),.BLN(BLN113),.WL(WL149));
sram_cell_6t_5 inst_cell_149_114 (.BL(BL114),.BLN(BLN114),.WL(WL149));
sram_cell_6t_5 inst_cell_149_115 (.BL(BL115),.BLN(BLN115),.WL(WL149));
sram_cell_6t_5 inst_cell_149_116 (.BL(BL116),.BLN(BLN116),.WL(WL149));
sram_cell_6t_5 inst_cell_149_117 (.BL(BL117),.BLN(BLN117),.WL(WL149));
sram_cell_6t_5 inst_cell_149_118 (.BL(BL118),.BLN(BLN118),.WL(WL149));
sram_cell_6t_5 inst_cell_149_119 (.BL(BL119),.BLN(BLN119),.WL(WL149));
sram_cell_6t_5 inst_cell_149_120 (.BL(BL120),.BLN(BLN120),.WL(WL149));
sram_cell_6t_5 inst_cell_149_121 (.BL(BL121),.BLN(BLN121),.WL(WL149));
sram_cell_6t_5 inst_cell_149_122 (.BL(BL122),.BLN(BLN122),.WL(WL149));
sram_cell_6t_5 inst_cell_149_123 (.BL(BL123),.BLN(BLN123),.WL(WL149));
sram_cell_6t_5 inst_cell_149_124 (.BL(BL124),.BLN(BLN124),.WL(WL149));
sram_cell_6t_5 inst_cell_149_125 (.BL(BL125),.BLN(BLN125),.WL(WL149));
sram_cell_6t_5 inst_cell_149_126 (.BL(BL126),.BLN(BLN126),.WL(WL149));
sram_cell_6t_5 inst_cell_149_127 (.BL(BL127),.BLN(BLN127),.WL(WL149));
sram_cell_6t_5 inst_cell_150_0 (.BL(BL0),.BLN(BLN0),.WL(WL150));
sram_cell_6t_5 inst_cell_150_1 (.BL(BL1),.BLN(BLN1),.WL(WL150));
sram_cell_6t_5 inst_cell_150_2 (.BL(BL2),.BLN(BLN2),.WL(WL150));
sram_cell_6t_5 inst_cell_150_3 (.BL(BL3),.BLN(BLN3),.WL(WL150));
sram_cell_6t_5 inst_cell_150_4 (.BL(BL4),.BLN(BLN4),.WL(WL150));
sram_cell_6t_5 inst_cell_150_5 (.BL(BL5),.BLN(BLN5),.WL(WL150));
sram_cell_6t_5 inst_cell_150_6 (.BL(BL6),.BLN(BLN6),.WL(WL150));
sram_cell_6t_5 inst_cell_150_7 (.BL(BL7),.BLN(BLN7),.WL(WL150));
sram_cell_6t_5 inst_cell_150_8 (.BL(BL8),.BLN(BLN8),.WL(WL150));
sram_cell_6t_5 inst_cell_150_9 (.BL(BL9),.BLN(BLN9),.WL(WL150));
sram_cell_6t_5 inst_cell_150_10 (.BL(BL10),.BLN(BLN10),.WL(WL150));
sram_cell_6t_5 inst_cell_150_11 (.BL(BL11),.BLN(BLN11),.WL(WL150));
sram_cell_6t_5 inst_cell_150_12 (.BL(BL12),.BLN(BLN12),.WL(WL150));
sram_cell_6t_5 inst_cell_150_13 (.BL(BL13),.BLN(BLN13),.WL(WL150));
sram_cell_6t_5 inst_cell_150_14 (.BL(BL14),.BLN(BLN14),.WL(WL150));
sram_cell_6t_5 inst_cell_150_15 (.BL(BL15),.BLN(BLN15),.WL(WL150));
sram_cell_6t_5 inst_cell_150_16 (.BL(BL16),.BLN(BLN16),.WL(WL150));
sram_cell_6t_5 inst_cell_150_17 (.BL(BL17),.BLN(BLN17),.WL(WL150));
sram_cell_6t_5 inst_cell_150_18 (.BL(BL18),.BLN(BLN18),.WL(WL150));
sram_cell_6t_5 inst_cell_150_19 (.BL(BL19),.BLN(BLN19),.WL(WL150));
sram_cell_6t_5 inst_cell_150_20 (.BL(BL20),.BLN(BLN20),.WL(WL150));
sram_cell_6t_5 inst_cell_150_21 (.BL(BL21),.BLN(BLN21),.WL(WL150));
sram_cell_6t_5 inst_cell_150_22 (.BL(BL22),.BLN(BLN22),.WL(WL150));
sram_cell_6t_5 inst_cell_150_23 (.BL(BL23),.BLN(BLN23),.WL(WL150));
sram_cell_6t_5 inst_cell_150_24 (.BL(BL24),.BLN(BLN24),.WL(WL150));
sram_cell_6t_5 inst_cell_150_25 (.BL(BL25),.BLN(BLN25),.WL(WL150));
sram_cell_6t_5 inst_cell_150_26 (.BL(BL26),.BLN(BLN26),.WL(WL150));
sram_cell_6t_5 inst_cell_150_27 (.BL(BL27),.BLN(BLN27),.WL(WL150));
sram_cell_6t_5 inst_cell_150_28 (.BL(BL28),.BLN(BLN28),.WL(WL150));
sram_cell_6t_5 inst_cell_150_29 (.BL(BL29),.BLN(BLN29),.WL(WL150));
sram_cell_6t_5 inst_cell_150_30 (.BL(BL30),.BLN(BLN30),.WL(WL150));
sram_cell_6t_5 inst_cell_150_31 (.BL(BL31),.BLN(BLN31),.WL(WL150));
sram_cell_6t_5 inst_cell_150_32 (.BL(BL32),.BLN(BLN32),.WL(WL150));
sram_cell_6t_5 inst_cell_150_33 (.BL(BL33),.BLN(BLN33),.WL(WL150));
sram_cell_6t_5 inst_cell_150_34 (.BL(BL34),.BLN(BLN34),.WL(WL150));
sram_cell_6t_5 inst_cell_150_35 (.BL(BL35),.BLN(BLN35),.WL(WL150));
sram_cell_6t_5 inst_cell_150_36 (.BL(BL36),.BLN(BLN36),.WL(WL150));
sram_cell_6t_5 inst_cell_150_37 (.BL(BL37),.BLN(BLN37),.WL(WL150));
sram_cell_6t_5 inst_cell_150_38 (.BL(BL38),.BLN(BLN38),.WL(WL150));
sram_cell_6t_5 inst_cell_150_39 (.BL(BL39),.BLN(BLN39),.WL(WL150));
sram_cell_6t_5 inst_cell_150_40 (.BL(BL40),.BLN(BLN40),.WL(WL150));
sram_cell_6t_5 inst_cell_150_41 (.BL(BL41),.BLN(BLN41),.WL(WL150));
sram_cell_6t_5 inst_cell_150_42 (.BL(BL42),.BLN(BLN42),.WL(WL150));
sram_cell_6t_5 inst_cell_150_43 (.BL(BL43),.BLN(BLN43),.WL(WL150));
sram_cell_6t_5 inst_cell_150_44 (.BL(BL44),.BLN(BLN44),.WL(WL150));
sram_cell_6t_5 inst_cell_150_45 (.BL(BL45),.BLN(BLN45),.WL(WL150));
sram_cell_6t_5 inst_cell_150_46 (.BL(BL46),.BLN(BLN46),.WL(WL150));
sram_cell_6t_5 inst_cell_150_47 (.BL(BL47),.BLN(BLN47),.WL(WL150));
sram_cell_6t_5 inst_cell_150_48 (.BL(BL48),.BLN(BLN48),.WL(WL150));
sram_cell_6t_5 inst_cell_150_49 (.BL(BL49),.BLN(BLN49),.WL(WL150));
sram_cell_6t_5 inst_cell_150_50 (.BL(BL50),.BLN(BLN50),.WL(WL150));
sram_cell_6t_5 inst_cell_150_51 (.BL(BL51),.BLN(BLN51),.WL(WL150));
sram_cell_6t_5 inst_cell_150_52 (.BL(BL52),.BLN(BLN52),.WL(WL150));
sram_cell_6t_5 inst_cell_150_53 (.BL(BL53),.BLN(BLN53),.WL(WL150));
sram_cell_6t_5 inst_cell_150_54 (.BL(BL54),.BLN(BLN54),.WL(WL150));
sram_cell_6t_5 inst_cell_150_55 (.BL(BL55),.BLN(BLN55),.WL(WL150));
sram_cell_6t_5 inst_cell_150_56 (.BL(BL56),.BLN(BLN56),.WL(WL150));
sram_cell_6t_5 inst_cell_150_57 (.BL(BL57),.BLN(BLN57),.WL(WL150));
sram_cell_6t_5 inst_cell_150_58 (.BL(BL58),.BLN(BLN58),.WL(WL150));
sram_cell_6t_5 inst_cell_150_59 (.BL(BL59),.BLN(BLN59),.WL(WL150));
sram_cell_6t_5 inst_cell_150_60 (.BL(BL60),.BLN(BLN60),.WL(WL150));
sram_cell_6t_5 inst_cell_150_61 (.BL(BL61),.BLN(BLN61),.WL(WL150));
sram_cell_6t_5 inst_cell_150_62 (.BL(BL62),.BLN(BLN62),.WL(WL150));
sram_cell_6t_5 inst_cell_150_63 (.BL(BL63),.BLN(BLN63),.WL(WL150));
sram_cell_6t_5 inst_cell_150_64 (.BL(BL64),.BLN(BLN64),.WL(WL150));
sram_cell_6t_5 inst_cell_150_65 (.BL(BL65),.BLN(BLN65),.WL(WL150));
sram_cell_6t_5 inst_cell_150_66 (.BL(BL66),.BLN(BLN66),.WL(WL150));
sram_cell_6t_5 inst_cell_150_67 (.BL(BL67),.BLN(BLN67),.WL(WL150));
sram_cell_6t_5 inst_cell_150_68 (.BL(BL68),.BLN(BLN68),.WL(WL150));
sram_cell_6t_5 inst_cell_150_69 (.BL(BL69),.BLN(BLN69),.WL(WL150));
sram_cell_6t_5 inst_cell_150_70 (.BL(BL70),.BLN(BLN70),.WL(WL150));
sram_cell_6t_5 inst_cell_150_71 (.BL(BL71),.BLN(BLN71),.WL(WL150));
sram_cell_6t_5 inst_cell_150_72 (.BL(BL72),.BLN(BLN72),.WL(WL150));
sram_cell_6t_5 inst_cell_150_73 (.BL(BL73),.BLN(BLN73),.WL(WL150));
sram_cell_6t_5 inst_cell_150_74 (.BL(BL74),.BLN(BLN74),.WL(WL150));
sram_cell_6t_5 inst_cell_150_75 (.BL(BL75),.BLN(BLN75),.WL(WL150));
sram_cell_6t_5 inst_cell_150_76 (.BL(BL76),.BLN(BLN76),.WL(WL150));
sram_cell_6t_5 inst_cell_150_77 (.BL(BL77),.BLN(BLN77),.WL(WL150));
sram_cell_6t_5 inst_cell_150_78 (.BL(BL78),.BLN(BLN78),.WL(WL150));
sram_cell_6t_5 inst_cell_150_79 (.BL(BL79),.BLN(BLN79),.WL(WL150));
sram_cell_6t_5 inst_cell_150_80 (.BL(BL80),.BLN(BLN80),.WL(WL150));
sram_cell_6t_5 inst_cell_150_81 (.BL(BL81),.BLN(BLN81),.WL(WL150));
sram_cell_6t_5 inst_cell_150_82 (.BL(BL82),.BLN(BLN82),.WL(WL150));
sram_cell_6t_5 inst_cell_150_83 (.BL(BL83),.BLN(BLN83),.WL(WL150));
sram_cell_6t_5 inst_cell_150_84 (.BL(BL84),.BLN(BLN84),.WL(WL150));
sram_cell_6t_5 inst_cell_150_85 (.BL(BL85),.BLN(BLN85),.WL(WL150));
sram_cell_6t_5 inst_cell_150_86 (.BL(BL86),.BLN(BLN86),.WL(WL150));
sram_cell_6t_5 inst_cell_150_87 (.BL(BL87),.BLN(BLN87),.WL(WL150));
sram_cell_6t_5 inst_cell_150_88 (.BL(BL88),.BLN(BLN88),.WL(WL150));
sram_cell_6t_5 inst_cell_150_89 (.BL(BL89),.BLN(BLN89),.WL(WL150));
sram_cell_6t_5 inst_cell_150_90 (.BL(BL90),.BLN(BLN90),.WL(WL150));
sram_cell_6t_5 inst_cell_150_91 (.BL(BL91),.BLN(BLN91),.WL(WL150));
sram_cell_6t_5 inst_cell_150_92 (.BL(BL92),.BLN(BLN92),.WL(WL150));
sram_cell_6t_5 inst_cell_150_93 (.BL(BL93),.BLN(BLN93),.WL(WL150));
sram_cell_6t_5 inst_cell_150_94 (.BL(BL94),.BLN(BLN94),.WL(WL150));
sram_cell_6t_5 inst_cell_150_95 (.BL(BL95),.BLN(BLN95),.WL(WL150));
sram_cell_6t_5 inst_cell_150_96 (.BL(BL96),.BLN(BLN96),.WL(WL150));
sram_cell_6t_5 inst_cell_150_97 (.BL(BL97),.BLN(BLN97),.WL(WL150));
sram_cell_6t_5 inst_cell_150_98 (.BL(BL98),.BLN(BLN98),.WL(WL150));
sram_cell_6t_5 inst_cell_150_99 (.BL(BL99),.BLN(BLN99),.WL(WL150));
sram_cell_6t_5 inst_cell_150_100 (.BL(BL100),.BLN(BLN100),.WL(WL150));
sram_cell_6t_5 inst_cell_150_101 (.BL(BL101),.BLN(BLN101),.WL(WL150));
sram_cell_6t_5 inst_cell_150_102 (.BL(BL102),.BLN(BLN102),.WL(WL150));
sram_cell_6t_5 inst_cell_150_103 (.BL(BL103),.BLN(BLN103),.WL(WL150));
sram_cell_6t_5 inst_cell_150_104 (.BL(BL104),.BLN(BLN104),.WL(WL150));
sram_cell_6t_5 inst_cell_150_105 (.BL(BL105),.BLN(BLN105),.WL(WL150));
sram_cell_6t_5 inst_cell_150_106 (.BL(BL106),.BLN(BLN106),.WL(WL150));
sram_cell_6t_5 inst_cell_150_107 (.BL(BL107),.BLN(BLN107),.WL(WL150));
sram_cell_6t_5 inst_cell_150_108 (.BL(BL108),.BLN(BLN108),.WL(WL150));
sram_cell_6t_5 inst_cell_150_109 (.BL(BL109),.BLN(BLN109),.WL(WL150));
sram_cell_6t_5 inst_cell_150_110 (.BL(BL110),.BLN(BLN110),.WL(WL150));
sram_cell_6t_5 inst_cell_150_111 (.BL(BL111),.BLN(BLN111),.WL(WL150));
sram_cell_6t_5 inst_cell_150_112 (.BL(BL112),.BLN(BLN112),.WL(WL150));
sram_cell_6t_5 inst_cell_150_113 (.BL(BL113),.BLN(BLN113),.WL(WL150));
sram_cell_6t_5 inst_cell_150_114 (.BL(BL114),.BLN(BLN114),.WL(WL150));
sram_cell_6t_5 inst_cell_150_115 (.BL(BL115),.BLN(BLN115),.WL(WL150));
sram_cell_6t_5 inst_cell_150_116 (.BL(BL116),.BLN(BLN116),.WL(WL150));
sram_cell_6t_5 inst_cell_150_117 (.BL(BL117),.BLN(BLN117),.WL(WL150));
sram_cell_6t_5 inst_cell_150_118 (.BL(BL118),.BLN(BLN118),.WL(WL150));
sram_cell_6t_5 inst_cell_150_119 (.BL(BL119),.BLN(BLN119),.WL(WL150));
sram_cell_6t_5 inst_cell_150_120 (.BL(BL120),.BLN(BLN120),.WL(WL150));
sram_cell_6t_5 inst_cell_150_121 (.BL(BL121),.BLN(BLN121),.WL(WL150));
sram_cell_6t_5 inst_cell_150_122 (.BL(BL122),.BLN(BLN122),.WL(WL150));
sram_cell_6t_5 inst_cell_150_123 (.BL(BL123),.BLN(BLN123),.WL(WL150));
sram_cell_6t_5 inst_cell_150_124 (.BL(BL124),.BLN(BLN124),.WL(WL150));
sram_cell_6t_5 inst_cell_150_125 (.BL(BL125),.BLN(BLN125),.WL(WL150));
sram_cell_6t_5 inst_cell_150_126 (.BL(BL126),.BLN(BLN126),.WL(WL150));
sram_cell_6t_5 inst_cell_150_127 (.BL(BL127),.BLN(BLN127),.WL(WL150));
sram_cell_6t_5 inst_cell_151_0 (.BL(BL0),.BLN(BLN0),.WL(WL151));
sram_cell_6t_5 inst_cell_151_1 (.BL(BL1),.BLN(BLN1),.WL(WL151));
sram_cell_6t_5 inst_cell_151_2 (.BL(BL2),.BLN(BLN2),.WL(WL151));
sram_cell_6t_5 inst_cell_151_3 (.BL(BL3),.BLN(BLN3),.WL(WL151));
sram_cell_6t_5 inst_cell_151_4 (.BL(BL4),.BLN(BLN4),.WL(WL151));
sram_cell_6t_5 inst_cell_151_5 (.BL(BL5),.BLN(BLN5),.WL(WL151));
sram_cell_6t_5 inst_cell_151_6 (.BL(BL6),.BLN(BLN6),.WL(WL151));
sram_cell_6t_5 inst_cell_151_7 (.BL(BL7),.BLN(BLN7),.WL(WL151));
sram_cell_6t_5 inst_cell_151_8 (.BL(BL8),.BLN(BLN8),.WL(WL151));
sram_cell_6t_5 inst_cell_151_9 (.BL(BL9),.BLN(BLN9),.WL(WL151));
sram_cell_6t_5 inst_cell_151_10 (.BL(BL10),.BLN(BLN10),.WL(WL151));
sram_cell_6t_5 inst_cell_151_11 (.BL(BL11),.BLN(BLN11),.WL(WL151));
sram_cell_6t_5 inst_cell_151_12 (.BL(BL12),.BLN(BLN12),.WL(WL151));
sram_cell_6t_5 inst_cell_151_13 (.BL(BL13),.BLN(BLN13),.WL(WL151));
sram_cell_6t_5 inst_cell_151_14 (.BL(BL14),.BLN(BLN14),.WL(WL151));
sram_cell_6t_5 inst_cell_151_15 (.BL(BL15),.BLN(BLN15),.WL(WL151));
sram_cell_6t_5 inst_cell_151_16 (.BL(BL16),.BLN(BLN16),.WL(WL151));
sram_cell_6t_5 inst_cell_151_17 (.BL(BL17),.BLN(BLN17),.WL(WL151));
sram_cell_6t_5 inst_cell_151_18 (.BL(BL18),.BLN(BLN18),.WL(WL151));
sram_cell_6t_5 inst_cell_151_19 (.BL(BL19),.BLN(BLN19),.WL(WL151));
sram_cell_6t_5 inst_cell_151_20 (.BL(BL20),.BLN(BLN20),.WL(WL151));
sram_cell_6t_5 inst_cell_151_21 (.BL(BL21),.BLN(BLN21),.WL(WL151));
sram_cell_6t_5 inst_cell_151_22 (.BL(BL22),.BLN(BLN22),.WL(WL151));
sram_cell_6t_5 inst_cell_151_23 (.BL(BL23),.BLN(BLN23),.WL(WL151));
sram_cell_6t_5 inst_cell_151_24 (.BL(BL24),.BLN(BLN24),.WL(WL151));
sram_cell_6t_5 inst_cell_151_25 (.BL(BL25),.BLN(BLN25),.WL(WL151));
sram_cell_6t_5 inst_cell_151_26 (.BL(BL26),.BLN(BLN26),.WL(WL151));
sram_cell_6t_5 inst_cell_151_27 (.BL(BL27),.BLN(BLN27),.WL(WL151));
sram_cell_6t_5 inst_cell_151_28 (.BL(BL28),.BLN(BLN28),.WL(WL151));
sram_cell_6t_5 inst_cell_151_29 (.BL(BL29),.BLN(BLN29),.WL(WL151));
sram_cell_6t_5 inst_cell_151_30 (.BL(BL30),.BLN(BLN30),.WL(WL151));
sram_cell_6t_5 inst_cell_151_31 (.BL(BL31),.BLN(BLN31),.WL(WL151));
sram_cell_6t_5 inst_cell_151_32 (.BL(BL32),.BLN(BLN32),.WL(WL151));
sram_cell_6t_5 inst_cell_151_33 (.BL(BL33),.BLN(BLN33),.WL(WL151));
sram_cell_6t_5 inst_cell_151_34 (.BL(BL34),.BLN(BLN34),.WL(WL151));
sram_cell_6t_5 inst_cell_151_35 (.BL(BL35),.BLN(BLN35),.WL(WL151));
sram_cell_6t_5 inst_cell_151_36 (.BL(BL36),.BLN(BLN36),.WL(WL151));
sram_cell_6t_5 inst_cell_151_37 (.BL(BL37),.BLN(BLN37),.WL(WL151));
sram_cell_6t_5 inst_cell_151_38 (.BL(BL38),.BLN(BLN38),.WL(WL151));
sram_cell_6t_5 inst_cell_151_39 (.BL(BL39),.BLN(BLN39),.WL(WL151));
sram_cell_6t_5 inst_cell_151_40 (.BL(BL40),.BLN(BLN40),.WL(WL151));
sram_cell_6t_5 inst_cell_151_41 (.BL(BL41),.BLN(BLN41),.WL(WL151));
sram_cell_6t_5 inst_cell_151_42 (.BL(BL42),.BLN(BLN42),.WL(WL151));
sram_cell_6t_5 inst_cell_151_43 (.BL(BL43),.BLN(BLN43),.WL(WL151));
sram_cell_6t_5 inst_cell_151_44 (.BL(BL44),.BLN(BLN44),.WL(WL151));
sram_cell_6t_5 inst_cell_151_45 (.BL(BL45),.BLN(BLN45),.WL(WL151));
sram_cell_6t_5 inst_cell_151_46 (.BL(BL46),.BLN(BLN46),.WL(WL151));
sram_cell_6t_5 inst_cell_151_47 (.BL(BL47),.BLN(BLN47),.WL(WL151));
sram_cell_6t_5 inst_cell_151_48 (.BL(BL48),.BLN(BLN48),.WL(WL151));
sram_cell_6t_5 inst_cell_151_49 (.BL(BL49),.BLN(BLN49),.WL(WL151));
sram_cell_6t_5 inst_cell_151_50 (.BL(BL50),.BLN(BLN50),.WL(WL151));
sram_cell_6t_5 inst_cell_151_51 (.BL(BL51),.BLN(BLN51),.WL(WL151));
sram_cell_6t_5 inst_cell_151_52 (.BL(BL52),.BLN(BLN52),.WL(WL151));
sram_cell_6t_5 inst_cell_151_53 (.BL(BL53),.BLN(BLN53),.WL(WL151));
sram_cell_6t_5 inst_cell_151_54 (.BL(BL54),.BLN(BLN54),.WL(WL151));
sram_cell_6t_5 inst_cell_151_55 (.BL(BL55),.BLN(BLN55),.WL(WL151));
sram_cell_6t_5 inst_cell_151_56 (.BL(BL56),.BLN(BLN56),.WL(WL151));
sram_cell_6t_5 inst_cell_151_57 (.BL(BL57),.BLN(BLN57),.WL(WL151));
sram_cell_6t_5 inst_cell_151_58 (.BL(BL58),.BLN(BLN58),.WL(WL151));
sram_cell_6t_5 inst_cell_151_59 (.BL(BL59),.BLN(BLN59),.WL(WL151));
sram_cell_6t_5 inst_cell_151_60 (.BL(BL60),.BLN(BLN60),.WL(WL151));
sram_cell_6t_5 inst_cell_151_61 (.BL(BL61),.BLN(BLN61),.WL(WL151));
sram_cell_6t_5 inst_cell_151_62 (.BL(BL62),.BLN(BLN62),.WL(WL151));
sram_cell_6t_5 inst_cell_151_63 (.BL(BL63),.BLN(BLN63),.WL(WL151));
sram_cell_6t_5 inst_cell_151_64 (.BL(BL64),.BLN(BLN64),.WL(WL151));
sram_cell_6t_5 inst_cell_151_65 (.BL(BL65),.BLN(BLN65),.WL(WL151));
sram_cell_6t_5 inst_cell_151_66 (.BL(BL66),.BLN(BLN66),.WL(WL151));
sram_cell_6t_5 inst_cell_151_67 (.BL(BL67),.BLN(BLN67),.WL(WL151));
sram_cell_6t_5 inst_cell_151_68 (.BL(BL68),.BLN(BLN68),.WL(WL151));
sram_cell_6t_5 inst_cell_151_69 (.BL(BL69),.BLN(BLN69),.WL(WL151));
sram_cell_6t_5 inst_cell_151_70 (.BL(BL70),.BLN(BLN70),.WL(WL151));
sram_cell_6t_5 inst_cell_151_71 (.BL(BL71),.BLN(BLN71),.WL(WL151));
sram_cell_6t_5 inst_cell_151_72 (.BL(BL72),.BLN(BLN72),.WL(WL151));
sram_cell_6t_5 inst_cell_151_73 (.BL(BL73),.BLN(BLN73),.WL(WL151));
sram_cell_6t_5 inst_cell_151_74 (.BL(BL74),.BLN(BLN74),.WL(WL151));
sram_cell_6t_5 inst_cell_151_75 (.BL(BL75),.BLN(BLN75),.WL(WL151));
sram_cell_6t_5 inst_cell_151_76 (.BL(BL76),.BLN(BLN76),.WL(WL151));
sram_cell_6t_5 inst_cell_151_77 (.BL(BL77),.BLN(BLN77),.WL(WL151));
sram_cell_6t_5 inst_cell_151_78 (.BL(BL78),.BLN(BLN78),.WL(WL151));
sram_cell_6t_5 inst_cell_151_79 (.BL(BL79),.BLN(BLN79),.WL(WL151));
sram_cell_6t_5 inst_cell_151_80 (.BL(BL80),.BLN(BLN80),.WL(WL151));
sram_cell_6t_5 inst_cell_151_81 (.BL(BL81),.BLN(BLN81),.WL(WL151));
sram_cell_6t_5 inst_cell_151_82 (.BL(BL82),.BLN(BLN82),.WL(WL151));
sram_cell_6t_5 inst_cell_151_83 (.BL(BL83),.BLN(BLN83),.WL(WL151));
sram_cell_6t_5 inst_cell_151_84 (.BL(BL84),.BLN(BLN84),.WL(WL151));
sram_cell_6t_5 inst_cell_151_85 (.BL(BL85),.BLN(BLN85),.WL(WL151));
sram_cell_6t_5 inst_cell_151_86 (.BL(BL86),.BLN(BLN86),.WL(WL151));
sram_cell_6t_5 inst_cell_151_87 (.BL(BL87),.BLN(BLN87),.WL(WL151));
sram_cell_6t_5 inst_cell_151_88 (.BL(BL88),.BLN(BLN88),.WL(WL151));
sram_cell_6t_5 inst_cell_151_89 (.BL(BL89),.BLN(BLN89),.WL(WL151));
sram_cell_6t_5 inst_cell_151_90 (.BL(BL90),.BLN(BLN90),.WL(WL151));
sram_cell_6t_5 inst_cell_151_91 (.BL(BL91),.BLN(BLN91),.WL(WL151));
sram_cell_6t_5 inst_cell_151_92 (.BL(BL92),.BLN(BLN92),.WL(WL151));
sram_cell_6t_5 inst_cell_151_93 (.BL(BL93),.BLN(BLN93),.WL(WL151));
sram_cell_6t_5 inst_cell_151_94 (.BL(BL94),.BLN(BLN94),.WL(WL151));
sram_cell_6t_5 inst_cell_151_95 (.BL(BL95),.BLN(BLN95),.WL(WL151));
sram_cell_6t_5 inst_cell_151_96 (.BL(BL96),.BLN(BLN96),.WL(WL151));
sram_cell_6t_5 inst_cell_151_97 (.BL(BL97),.BLN(BLN97),.WL(WL151));
sram_cell_6t_5 inst_cell_151_98 (.BL(BL98),.BLN(BLN98),.WL(WL151));
sram_cell_6t_5 inst_cell_151_99 (.BL(BL99),.BLN(BLN99),.WL(WL151));
sram_cell_6t_5 inst_cell_151_100 (.BL(BL100),.BLN(BLN100),.WL(WL151));
sram_cell_6t_5 inst_cell_151_101 (.BL(BL101),.BLN(BLN101),.WL(WL151));
sram_cell_6t_5 inst_cell_151_102 (.BL(BL102),.BLN(BLN102),.WL(WL151));
sram_cell_6t_5 inst_cell_151_103 (.BL(BL103),.BLN(BLN103),.WL(WL151));
sram_cell_6t_5 inst_cell_151_104 (.BL(BL104),.BLN(BLN104),.WL(WL151));
sram_cell_6t_5 inst_cell_151_105 (.BL(BL105),.BLN(BLN105),.WL(WL151));
sram_cell_6t_5 inst_cell_151_106 (.BL(BL106),.BLN(BLN106),.WL(WL151));
sram_cell_6t_5 inst_cell_151_107 (.BL(BL107),.BLN(BLN107),.WL(WL151));
sram_cell_6t_5 inst_cell_151_108 (.BL(BL108),.BLN(BLN108),.WL(WL151));
sram_cell_6t_5 inst_cell_151_109 (.BL(BL109),.BLN(BLN109),.WL(WL151));
sram_cell_6t_5 inst_cell_151_110 (.BL(BL110),.BLN(BLN110),.WL(WL151));
sram_cell_6t_5 inst_cell_151_111 (.BL(BL111),.BLN(BLN111),.WL(WL151));
sram_cell_6t_5 inst_cell_151_112 (.BL(BL112),.BLN(BLN112),.WL(WL151));
sram_cell_6t_5 inst_cell_151_113 (.BL(BL113),.BLN(BLN113),.WL(WL151));
sram_cell_6t_5 inst_cell_151_114 (.BL(BL114),.BLN(BLN114),.WL(WL151));
sram_cell_6t_5 inst_cell_151_115 (.BL(BL115),.BLN(BLN115),.WL(WL151));
sram_cell_6t_5 inst_cell_151_116 (.BL(BL116),.BLN(BLN116),.WL(WL151));
sram_cell_6t_5 inst_cell_151_117 (.BL(BL117),.BLN(BLN117),.WL(WL151));
sram_cell_6t_5 inst_cell_151_118 (.BL(BL118),.BLN(BLN118),.WL(WL151));
sram_cell_6t_5 inst_cell_151_119 (.BL(BL119),.BLN(BLN119),.WL(WL151));
sram_cell_6t_5 inst_cell_151_120 (.BL(BL120),.BLN(BLN120),.WL(WL151));
sram_cell_6t_5 inst_cell_151_121 (.BL(BL121),.BLN(BLN121),.WL(WL151));
sram_cell_6t_5 inst_cell_151_122 (.BL(BL122),.BLN(BLN122),.WL(WL151));
sram_cell_6t_5 inst_cell_151_123 (.BL(BL123),.BLN(BLN123),.WL(WL151));
sram_cell_6t_5 inst_cell_151_124 (.BL(BL124),.BLN(BLN124),.WL(WL151));
sram_cell_6t_5 inst_cell_151_125 (.BL(BL125),.BLN(BLN125),.WL(WL151));
sram_cell_6t_5 inst_cell_151_126 (.BL(BL126),.BLN(BLN126),.WL(WL151));
sram_cell_6t_5 inst_cell_151_127 (.BL(BL127),.BLN(BLN127),.WL(WL151));
sram_cell_6t_5 inst_cell_152_0 (.BL(BL0),.BLN(BLN0),.WL(WL152));
sram_cell_6t_5 inst_cell_152_1 (.BL(BL1),.BLN(BLN1),.WL(WL152));
sram_cell_6t_5 inst_cell_152_2 (.BL(BL2),.BLN(BLN2),.WL(WL152));
sram_cell_6t_5 inst_cell_152_3 (.BL(BL3),.BLN(BLN3),.WL(WL152));
sram_cell_6t_5 inst_cell_152_4 (.BL(BL4),.BLN(BLN4),.WL(WL152));
sram_cell_6t_5 inst_cell_152_5 (.BL(BL5),.BLN(BLN5),.WL(WL152));
sram_cell_6t_5 inst_cell_152_6 (.BL(BL6),.BLN(BLN6),.WL(WL152));
sram_cell_6t_5 inst_cell_152_7 (.BL(BL7),.BLN(BLN7),.WL(WL152));
sram_cell_6t_5 inst_cell_152_8 (.BL(BL8),.BLN(BLN8),.WL(WL152));
sram_cell_6t_5 inst_cell_152_9 (.BL(BL9),.BLN(BLN9),.WL(WL152));
sram_cell_6t_5 inst_cell_152_10 (.BL(BL10),.BLN(BLN10),.WL(WL152));
sram_cell_6t_5 inst_cell_152_11 (.BL(BL11),.BLN(BLN11),.WL(WL152));
sram_cell_6t_5 inst_cell_152_12 (.BL(BL12),.BLN(BLN12),.WL(WL152));
sram_cell_6t_5 inst_cell_152_13 (.BL(BL13),.BLN(BLN13),.WL(WL152));
sram_cell_6t_5 inst_cell_152_14 (.BL(BL14),.BLN(BLN14),.WL(WL152));
sram_cell_6t_5 inst_cell_152_15 (.BL(BL15),.BLN(BLN15),.WL(WL152));
sram_cell_6t_5 inst_cell_152_16 (.BL(BL16),.BLN(BLN16),.WL(WL152));
sram_cell_6t_5 inst_cell_152_17 (.BL(BL17),.BLN(BLN17),.WL(WL152));
sram_cell_6t_5 inst_cell_152_18 (.BL(BL18),.BLN(BLN18),.WL(WL152));
sram_cell_6t_5 inst_cell_152_19 (.BL(BL19),.BLN(BLN19),.WL(WL152));
sram_cell_6t_5 inst_cell_152_20 (.BL(BL20),.BLN(BLN20),.WL(WL152));
sram_cell_6t_5 inst_cell_152_21 (.BL(BL21),.BLN(BLN21),.WL(WL152));
sram_cell_6t_5 inst_cell_152_22 (.BL(BL22),.BLN(BLN22),.WL(WL152));
sram_cell_6t_5 inst_cell_152_23 (.BL(BL23),.BLN(BLN23),.WL(WL152));
sram_cell_6t_5 inst_cell_152_24 (.BL(BL24),.BLN(BLN24),.WL(WL152));
sram_cell_6t_5 inst_cell_152_25 (.BL(BL25),.BLN(BLN25),.WL(WL152));
sram_cell_6t_5 inst_cell_152_26 (.BL(BL26),.BLN(BLN26),.WL(WL152));
sram_cell_6t_5 inst_cell_152_27 (.BL(BL27),.BLN(BLN27),.WL(WL152));
sram_cell_6t_5 inst_cell_152_28 (.BL(BL28),.BLN(BLN28),.WL(WL152));
sram_cell_6t_5 inst_cell_152_29 (.BL(BL29),.BLN(BLN29),.WL(WL152));
sram_cell_6t_5 inst_cell_152_30 (.BL(BL30),.BLN(BLN30),.WL(WL152));
sram_cell_6t_5 inst_cell_152_31 (.BL(BL31),.BLN(BLN31),.WL(WL152));
sram_cell_6t_5 inst_cell_152_32 (.BL(BL32),.BLN(BLN32),.WL(WL152));
sram_cell_6t_5 inst_cell_152_33 (.BL(BL33),.BLN(BLN33),.WL(WL152));
sram_cell_6t_5 inst_cell_152_34 (.BL(BL34),.BLN(BLN34),.WL(WL152));
sram_cell_6t_5 inst_cell_152_35 (.BL(BL35),.BLN(BLN35),.WL(WL152));
sram_cell_6t_5 inst_cell_152_36 (.BL(BL36),.BLN(BLN36),.WL(WL152));
sram_cell_6t_5 inst_cell_152_37 (.BL(BL37),.BLN(BLN37),.WL(WL152));
sram_cell_6t_5 inst_cell_152_38 (.BL(BL38),.BLN(BLN38),.WL(WL152));
sram_cell_6t_5 inst_cell_152_39 (.BL(BL39),.BLN(BLN39),.WL(WL152));
sram_cell_6t_5 inst_cell_152_40 (.BL(BL40),.BLN(BLN40),.WL(WL152));
sram_cell_6t_5 inst_cell_152_41 (.BL(BL41),.BLN(BLN41),.WL(WL152));
sram_cell_6t_5 inst_cell_152_42 (.BL(BL42),.BLN(BLN42),.WL(WL152));
sram_cell_6t_5 inst_cell_152_43 (.BL(BL43),.BLN(BLN43),.WL(WL152));
sram_cell_6t_5 inst_cell_152_44 (.BL(BL44),.BLN(BLN44),.WL(WL152));
sram_cell_6t_5 inst_cell_152_45 (.BL(BL45),.BLN(BLN45),.WL(WL152));
sram_cell_6t_5 inst_cell_152_46 (.BL(BL46),.BLN(BLN46),.WL(WL152));
sram_cell_6t_5 inst_cell_152_47 (.BL(BL47),.BLN(BLN47),.WL(WL152));
sram_cell_6t_5 inst_cell_152_48 (.BL(BL48),.BLN(BLN48),.WL(WL152));
sram_cell_6t_5 inst_cell_152_49 (.BL(BL49),.BLN(BLN49),.WL(WL152));
sram_cell_6t_5 inst_cell_152_50 (.BL(BL50),.BLN(BLN50),.WL(WL152));
sram_cell_6t_5 inst_cell_152_51 (.BL(BL51),.BLN(BLN51),.WL(WL152));
sram_cell_6t_5 inst_cell_152_52 (.BL(BL52),.BLN(BLN52),.WL(WL152));
sram_cell_6t_5 inst_cell_152_53 (.BL(BL53),.BLN(BLN53),.WL(WL152));
sram_cell_6t_5 inst_cell_152_54 (.BL(BL54),.BLN(BLN54),.WL(WL152));
sram_cell_6t_5 inst_cell_152_55 (.BL(BL55),.BLN(BLN55),.WL(WL152));
sram_cell_6t_5 inst_cell_152_56 (.BL(BL56),.BLN(BLN56),.WL(WL152));
sram_cell_6t_5 inst_cell_152_57 (.BL(BL57),.BLN(BLN57),.WL(WL152));
sram_cell_6t_5 inst_cell_152_58 (.BL(BL58),.BLN(BLN58),.WL(WL152));
sram_cell_6t_5 inst_cell_152_59 (.BL(BL59),.BLN(BLN59),.WL(WL152));
sram_cell_6t_5 inst_cell_152_60 (.BL(BL60),.BLN(BLN60),.WL(WL152));
sram_cell_6t_5 inst_cell_152_61 (.BL(BL61),.BLN(BLN61),.WL(WL152));
sram_cell_6t_5 inst_cell_152_62 (.BL(BL62),.BLN(BLN62),.WL(WL152));
sram_cell_6t_5 inst_cell_152_63 (.BL(BL63),.BLN(BLN63),.WL(WL152));
sram_cell_6t_5 inst_cell_152_64 (.BL(BL64),.BLN(BLN64),.WL(WL152));
sram_cell_6t_5 inst_cell_152_65 (.BL(BL65),.BLN(BLN65),.WL(WL152));
sram_cell_6t_5 inst_cell_152_66 (.BL(BL66),.BLN(BLN66),.WL(WL152));
sram_cell_6t_5 inst_cell_152_67 (.BL(BL67),.BLN(BLN67),.WL(WL152));
sram_cell_6t_5 inst_cell_152_68 (.BL(BL68),.BLN(BLN68),.WL(WL152));
sram_cell_6t_5 inst_cell_152_69 (.BL(BL69),.BLN(BLN69),.WL(WL152));
sram_cell_6t_5 inst_cell_152_70 (.BL(BL70),.BLN(BLN70),.WL(WL152));
sram_cell_6t_5 inst_cell_152_71 (.BL(BL71),.BLN(BLN71),.WL(WL152));
sram_cell_6t_5 inst_cell_152_72 (.BL(BL72),.BLN(BLN72),.WL(WL152));
sram_cell_6t_5 inst_cell_152_73 (.BL(BL73),.BLN(BLN73),.WL(WL152));
sram_cell_6t_5 inst_cell_152_74 (.BL(BL74),.BLN(BLN74),.WL(WL152));
sram_cell_6t_5 inst_cell_152_75 (.BL(BL75),.BLN(BLN75),.WL(WL152));
sram_cell_6t_5 inst_cell_152_76 (.BL(BL76),.BLN(BLN76),.WL(WL152));
sram_cell_6t_5 inst_cell_152_77 (.BL(BL77),.BLN(BLN77),.WL(WL152));
sram_cell_6t_5 inst_cell_152_78 (.BL(BL78),.BLN(BLN78),.WL(WL152));
sram_cell_6t_5 inst_cell_152_79 (.BL(BL79),.BLN(BLN79),.WL(WL152));
sram_cell_6t_5 inst_cell_152_80 (.BL(BL80),.BLN(BLN80),.WL(WL152));
sram_cell_6t_5 inst_cell_152_81 (.BL(BL81),.BLN(BLN81),.WL(WL152));
sram_cell_6t_5 inst_cell_152_82 (.BL(BL82),.BLN(BLN82),.WL(WL152));
sram_cell_6t_5 inst_cell_152_83 (.BL(BL83),.BLN(BLN83),.WL(WL152));
sram_cell_6t_5 inst_cell_152_84 (.BL(BL84),.BLN(BLN84),.WL(WL152));
sram_cell_6t_5 inst_cell_152_85 (.BL(BL85),.BLN(BLN85),.WL(WL152));
sram_cell_6t_5 inst_cell_152_86 (.BL(BL86),.BLN(BLN86),.WL(WL152));
sram_cell_6t_5 inst_cell_152_87 (.BL(BL87),.BLN(BLN87),.WL(WL152));
sram_cell_6t_5 inst_cell_152_88 (.BL(BL88),.BLN(BLN88),.WL(WL152));
sram_cell_6t_5 inst_cell_152_89 (.BL(BL89),.BLN(BLN89),.WL(WL152));
sram_cell_6t_5 inst_cell_152_90 (.BL(BL90),.BLN(BLN90),.WL(WL152));
sram_cell_6t_5 inst_cell_152_91 (.BL(BL91),.BLN(BLN91),.WL(WL152));
sram_cell_6t_5 inst_cell_152_92 (.BL(BL92),.BLN(BLN92),.WL(WL152));
sram_cell_6t_5 inst_cell_152_93 (.BL(BL93),.BLN(BLN93),.WL(WL152));
sram_cell_6t_5 inst_cell_152_94 (.BL(BL94),.BLN(BLN94),.WL(WL152));
sram_cell_6t_5 inst_cell_152_95 (.BL(BL95),.BLN(BLN95),.WL(WL152));
sram_cell_6t_5 inst_cell_152_96 (.BL(BL96),.BLN(BLN96),.WL(WL152));
sram_cell_6t_5 inst_cell_152_97 (.BL(BL97),.BLN(BLN97),.WL(WL152));
sram_cell_6t_5 inst_cell_152_98 (.BL(BL98),.BLN(BLN98),.WL(WL152));
sram_cell_6t_5 inst_cell_152_99 (.BL(BL99),.BLN(BLN99),.WL(WL152));
sram_cell_6t_5 inst_cell_152_100 (.BL(BL100),.BLN(BLN100),.WL(WL152));
sram_cell_6t_5 inst_cell_152_101 (.BL(BL101),.BLN(BLN101),.WL(WL152));
sram_cell_6t_5 inst_cell_152_102 (.BL(BL102),.BLN(BLN102),.WL(WL152));
sram_cell_6t_5 inst_cell_152_103 (.BL(BL103),.BLN(BLN103),.WL(WL152));
sram_cell_6t_5 inst_cell_152_104 (.BL(BL104),.BLN(BLN104),.WL(WL152));
sram_cell_6t_5 inst_cell_152_105 (.BL(BL105),.BLN(BLN105),.WL(WL152));
sram_cell_6t_5 inst_cell_152_106 (.BL(BL106),.BLN(BLN106),.WL(WL152));
sram_cell_6t_5 inst_cell_152_107 (.BL(BL107),.BLN(BLN107),.WL(WL152));
sram_cell_6t_5 inst_cell_152_108 (.BL(BL108),.BLN(BLN108),.WL(WL152));
sram_cell_6t_5 inst_cell_152_109 (.BL(BL109),.BLN(BLN109),.WL(WL152));
sram_cell_6t_5 inst_cell_152_110 (.BL(BL110),.BLN(BLN110),.WL(WL152));
sram_cell_6t_5 inst_cell_152_111 (.BL(BL111),.BLN(BLN111),.WL(WL152));
sram_cell_6t_5 inst_cell_152_112 (.BL(BL112),.BLN(BLN112),.WL(WL152));
sram_cell_6t_5 inst_cell_152_113 (.BL(BL113),.BLN(BLN113),.WL(WL152));
sram_cell_6t_5 inst_cell_152_114 (.BL(BL114),.BLN(BLN114),.WL(WL152));
sram_cell_6t_5 inst_cell_152_115 (.BL(BL115),.BLN(BLN115),.WL(WL152));
sram_cell_6t_5 inst_cell_152_116 (.BL(BL116),.BLN(BLN116),.WL(WL152));
sram_cell_6t_5 inst_cell_152_117 (.BL(BL117),.BLN(BLN117),.WL(WL152));
sram_cell_6t_5 inst_cell_152_118 (.BL(BL118),.BLN(BLN118),.WL(WL152));
sram_cell_6t_5 inst_cell_152_119 (.BL(BL119),.BLN(BLN119),.WL(WL152));
sram_cell_6t_5 inst_cell_152_120 (.BL(BL120),.BLN(BLN120),.WL(WL152));
sram_cell_6t_5 inst_cell_152_121 (.BL(BL121),.BLN(BLN121),.WL(WL152));
sram_cell_6t_5 inst_cell_152_122 (.BL(BL122),.BLN(BLN122),.WL(WL152));
sram_cell_6t_5 inst_cell_152_123 (.BL(BL123),.BLN(BLN123),.WL(WL152));
sram_cell_6t_5 inst_cell_152_124 (.BL(BL124),.BLN(BLN124),.WL(WL152));
sram_cell_6t_5 inst_cell_152_125 (.BL(BL125),.BLN(BLN125),.WL(WL152));
sram_cell_6t_5 inst_cell_152_126 (.BL(BL126),.BLN(BLN126),.WL(WL152));
sram_cell_6t_5 inst_cell_152_127 (.BL(BL127),.BLN(BLN127),.WL(WL152));
sram_cell_6t_5 inst_cell_153_0 (.BL(BL0),.BLN(BLN0),.WL(WL153));
sram_cell_6t_5 inst_cell_153_1 (.BL(BL1),.BLN(BLN1),.WL(WL153));
sram_cell_6t_5 inst_cell_153_2 (.BL(BL2),.BLN(BLN2),.WL(WL153));
sram_cell_6t_5 inst_cell_153_3 (.BL(BL3),.BLN(BLN3),.WL(WL153));
sram_cell_6t_5 inst_cell_153_4 (.BL(BL4),.BLN(BLN4),.WL(WL153));
sram_cell_6t_5 inst_cell_153_5 (.BL(BL5),.BLN(BLN5),.WL(WL153));
sram_cell_6t_5 inst_cell_153_6 (.BL(BL6),.BLN(BLN6),.WL(WL153));
sram_cell_6t_5 inst_cell_153_7 (.BL(BL7),.BLN(BLN7),.WL(WL153));
sram_cell_6t_5 inst_cell_153_8 (.BL(BL8),.BLN(BLN8),.WL(WL153));
sram_cell_6t_5 inst_cell_153_9 (.BL(BL9),.BLN(BLN9),.WL(WL153));
sram_cell_6t_5 inst_cell_153_10 (.BL(BL10),.BLN(BLN10),.WL(WL153));
sram_cell_6t_5 inst_cell_153_11 (.BL(BL11),.BLN(BLN11),.WL(WL153));
sram_cell_6t_5 inst_cell_153_12 (.BL(BL12),.BLN(BLN12),.WL(WL153));
sram_cell_6t_5 inst_cell_153_13 (.BL(BL13),.BLN(BLN13),.WL(WL153));
sram_cell_6t_5 inst_cell_153_14 (.BL(BL14),.BLN(BLN14),.WL(WL153));
sram_cell_6t_5 inst_cell_153_15 (.BL(BL15),.BLN(BLN15),.WL(WL153));
sram_cell_6t_5 inst_cell_153_16 (.BL(BL16),.BLN(BLN16),.WL(WL153));
sram_cell_6t_5 inst_cell_153_17 (.BL(BL17),.BLN(BLN17),.WL(WL153));
sram_cell_6t_5 inst_cell_153_18 (.BL(BL18),.BLN(BLN18),.WL(WL153));
sram_cell_6t_5 inst_cell_153_19 (.BL(BL19),.BLN(BLN19),.WL(WL153));
sram_cell_6t_5 inst_cell_153_20 (.BL(BL20),.BLN(BLN20),.WL(WL153));
sram_cell_6t_5 inst_cell_153_21 (.BL(BL21),.BLN(BLN21),.WL(WL153));
sram_cell_6t_5 inst_cell_153_22 (.BL(BL22),.BLN(BLN22),.WL(WL153));
sram_cell_6t_5 inst_cell_153_23 (.BL(BL23),.BLN(BLN23),.WL(WL153));
sram_cell_6t_5 inst_cell_153_24 (.BL(BL24),.BLN(BLN24),.WL(WL153));
sram_cell_6t_5 inst_cell_153_25 (.BL(BL25),.BLN(BLN25),.WL(WL153));
sram_cell_6t_5 inst_cell_153_26 (.BL(BL26),.BLN(BLN26),.WL(WL153));
sram_cell_6t_5 inst_cell_153_27 (.BL(BL27),.BLN(BLN27),.WL(WL153));
sram_cell_6t_5 inst_cell_153_28 (.BL(BL28),.BLN(BLN28),.WL(WL153));
sram_cell_6t_5 inst_cell_153_29 (.BL(BL29),.BLN(BLN29),.WL(WL153));
sram_cell_6t_5 inst_cell_153_30 (.BL(BL30),.BLN(BLN30),.WL(WL153));
sram_cell_6t_5 inst_cell_153_31 (.BL(BL31),.BLN(BLN31),.WL(WL153));
sram_cell_6t_5 inst_cell_153_32 (.BL(BL32),.BLN(BLN32),.WL(WL153));
sram_cell_6t_5 inst_cell_153_33 (.BL(BL33),.BLN(BLN33),.WL(WL153));
sram_cell_6t_5 inst_cell_153_34 (.BL(BL34),.BLN(BLN34),.WL(WL153));
sram_cell_6t_5 inst_cell_153_35 (.BL(BL35),.BLN(BLN35),.WL(WL153));
sram_cell_6t_5 inst_cell_153_36 (.BL(BL36),.BLN(BLN36),.WL(WL153));
sram_cell_6t_5 inst_cell_153_37 (.BL(BL37),.BLN(BLN37),.WL(WL153));
sram_cell_6t_5 inst_cell_153_38 (.BL(BL38),.BLN(BLN38),.WL(WL153));
sram_cell_6t_5 inst_cell_153_39 (.BL(BL39),.BLN(BLN39),.WL(WL153));
sram_cell_6t_5 inst_cell_153_40 (.BL(BL40),.BLN(BLN40),.WL(WL153));
sram_cell_6t_5 inst_cell_153_41 (.BL(BL41),.BLN(BLN41),.WL(WL153));
sram_cell_6t_5 inst_cell_153_42 (.BL(BL42),.BLN(BLN42),.WL(WL153));
sram_cell_6t_5 inst_cell_153_43 (.BL(BL43),.BLN(BLN43),.WL(WL153));
sram_cell_6t_5 inst_cell_153_44 (.BL(BL44),.BLN(BLN44),.WL(WL153));
sram_cell_6t_5 inst_cell_153_45 (.BL(BL45),.BLN(BLN45),.WL(WL153));
sram_cell_6t_5 inst_cell_153_46 (.BL(BL46),.BLN(BLN46),.WL(WL153));
sram_cell_6t_5 inst_cell_153_47 (.BL(BL47),.BLN(BLN47),.WL(WL153));
sram_cell_6t_5 inst_cell_153_48 (.BL(BL48),.BLN(BLN48),.WL(WL153));
sram_cell_6t_5 inst_cell_153_49 (.BL(BL49),.BLN(BLN49),.WL(WL153));
sram_cell_6t_5 inst_cell_153_50 (.BL(BL50),.BLN(BLN50),.WL(WL153));
sram_cell_6t_5 inst_cell_153_51 (.BL(BL51),.BLN(BLN51),.WL(WL153));
sram_cell_6t_5 inst_cell_153_52 (.BL(BL52),.BLN(BLN52),.WL(WL153));
sram_cell_6t_5 inst_cell_153_53 (.BL(BL53),.BLN(BLN53),.WL(WL153));
sram_cell_6t_5 inst_cell_153_54 (.BL(BL54),.BLN(BLN54),.WL(WL153));
sram_cell_6t_5 inst_cell_153_55 (.BL(BL55),.BLN(BLN55),.WL(WL153));
sram_cell_6t_5 inst_cell_153_56 (.BL(BL56),.BLN(BLN56),.WL(WL153));
sram_cell_6t_5 inst_cell_153_57 (.BL(BL57),.BLN(BLN57),.WL(WL153));
sram_cell_6t_5 inst_cell_153_58 (.BL(BL58),.BLN(BLN58),.WL(WL153));
sram_cell_6t_5 inst_cell_153_59 (.BL(BL59),.BLN(BLN59),.WL(WL153));
sram_cell_6t_5 inst_cell_153_60 (.BL(BL60),.BLN(BLN60),.WL(WL153));
sram_cell_6t_5 inst_cell_153_61 (.BL(BL61),.BLN(BLN61),.WL(WL153));
sram_cell_6t_5 inst_cell_153_62 (.BL(BL62),.BLN(BLN62),.WL(WL153));
sram_cell_6t_5 inst_cell_153_63 (.BL(BL63),.BLN(BLN63),.WL(WL153));
sram_cell_6t_5 inst_cell_153_64 (.BL(BL64),.BLN(BLN64),.WL(WL153));
sram_cell_6t_5 inst_cell_153_65 (.BL(BL65),.BLN(BLN65),.WL(WL153));
sram_cell_6t_5 inst_cell_153_66 (.BL(BL66),.BLN(BLN66),.WL(WL153));
sram_cell_6t_5 inst_cell_153_67 (.BL(BL67),.BLN(BLN67),.WL(WL153));
sram_cell_6t_5 inst_cell_153_68 (.BL(BL68),.BLN(BLN68),.WL(WL153));
sram_cell_6t_5 inst_cell_153_69 (.BL(BL69),.BLN(BLN69),.WL(WL153));
sram_cell_6t_5 inst_cell_153_70 (.BL(BL70),.BLN(BLN70),.WL(WL153));
sram_cell_6t_5 inst_cell_153_71 (.BL(BL71),.BLN(BLN71),.WL(WL153));
sram_cell_6t_5 inst_cell_153_72 (.BL(BL72),.BLN(BLN72),.WL(WL153));
sram_cell_6t_5 inst_cell_153_73 (.BL(BL73),.BLN(BLN73),.WL(WL153));
sram_cell_6t_5 inst_cell_153_74 (.BL(BL74),.BLN(BLN74),.WL(WL153));
sram_cell_6t_5 inst_cell_153_75 (.BL(BL75),.BLN(BLN75),.WL(WL153));
sram_cell_6t_5 inst_cell_153_76 (.BL(BL76),.BLN(BLN76),.WL(WL153));
sram_cell_6t_5 inst_cell_153_77 (.BL(BL77),.BLN(BLN77),.WL(WL153));
sram_cell_6t_5 inst_cell_153_78 (.BL(BL78),.BLN(BLN78),.WL(WL153));
sram_cell_6t_5 inst_cell_153_79 (.BL(BL79),.BLN(BLN79),.WL(WL153));
sram_cell_6t_5 inst_cell_153_80 (.BL(BL80),.BLN(BLN80),.WL(WL153));
sram_cell_6t_5 inst_cell_153_81 (.BL(BL81),.BLN(BLN81),.WL(WL153));
sram_cell_6t_5 inst_cell_153_82 (.BL(BL82),.BLN(BLN82),.WL(WL153));
sram_cell_6t_5 inst_cell_153_83 (.BL(BL83),.BLN(BLN83),.WL(WL153));
sram_cell_6t_5 inst_cell_153_84 (.BL(BL84),.BLN(BLN84),.WL(WL153));
sram_cell_6t_5 inst_cell_153_85 (.BL(BL85),.BLN(BLN85),.WL(WL153));
sram_cell_6t_5 inst_cell_153_86 (.BL(BL86),.BLN(BLN86),.WL(WL153));
sram_cell_6t_5 inst_cell_153_87 (.BL(BL87),.BLN(BLN87),.WL(WL153));
sram_cell_6t_5 inst_cell_153_88 (.BL(BL88),.BLN(BLN88),.WL(WL153));
sram_cell_6t_5 inst_cell_153_89 (.BL(BL89),.BLN(BLN89),.WL(WL153));
sram_cell_6t_5 inst_cell_153_90 (.BL(BL90),.BLN(BLN90),.WL(WL153));
sram_cell_6t_5 inst_cell_153_91 (.BL(BL91),.BLN(BLN91),.WL(WL153));
sram_cell_6t_5 inst_cell_153_92 (.BL(BL92),.BLN(BLN92),.WL(WL153));
sram_cell_6t_5 inst_cell_153_93 (.BL(BL93),.BLN(BLN93),.WL(WL153));
sram_cell_6t_5 inst_cell_153_94 (.BL(BL94),.BLN(BLN94),.WL(WL153));
sram_cell_6t_5 inst_cell_153_95 (.BL(BL95),.BLN(BLN95),.WL(WL153));
sram_cell_6t_5 inst_cell_153_96 (.BL(BL96),.BLN(BLN96),.WL(WL153));
sram_cell_6t_5 inst_cell_153_97 (.BL(BL97),.BLN(BLN97),.WL(WL153));
sram_cell_6t_5 inst_cell_153_98 (.BL(BL98),.BLN(BLN98),.WL(WL153));
sram_cell_6t_5 inst_cell_153_99 (.BL(BL99),.BLN(BLN99),.WL(WL153));
sram_cell_6t_5 inst_cell_153_100 (.BL(BL100),.BLN(BLN100),.WL(WL153));
sram_cell_6t_5 inst_cell_153_101 (.BL(BL101),.BLN(BLN101),.WL(WL153));
sram_cell_6t_5 inst_cell_153_102 (.BL(BL102),.BLN(BLN102),.WL(WL153));
sram_cell_6t_5 inst_cell_153_103 (.BL(BL103),.BLN(BLN103),.WL(WL153));
sram_cell_6t_5 inst_cell_153_104 (.BL(BL104),.BLN(BLN104),.WL(WL153));
sram_cell_6t_5 inst_cell_153_105 (.BL(BL105),.BLN(BLN105),.WL(WL153));
sram_cell_6t_5 inst_cell_153_106 (.BL(BL106),.BLN(BLN106),.WL(WL153));
sram_cell_6t_5 inst_cell_153_107 (.BL(BL107),.BLN(BLN107),.WL(WL153));
sram_cell_6t_5 inst_cell_153_108 (.BL(BL108),.BLN(BLN108),.WL(WL153));
sram_cell_6t_5 inst_cell_153_109 (.BL(BL109),.BLN(BLN109),.WL(WL153));
sram_cell_6t_5 inst_cell_153_110 (.BL(BL110),.BLN(BLN110),.WL(WL153));
sram_cell_6t_5 inst_cell_153_111 (.BL(BL111),.BLN(BLN111),.WL(WL153));
sram_cell_6t_5 inst_cell_153_112 (.BL(BL112),.BLN(BLN112),.WL(WL153));
sram_cell_6t_5 inst_cell_153_113 (.BL(BL113),.BLN(BLN113),.WL(WL153));
sram_cell_6t_5 inst_cell_153_114 (.BL(BL114),.BLN(BLN114),.WL(WL153));
sram_cell_6t_5 inst_cell_153_115 (.BL(BL115),.BLN(BLN115),.WL(WL153));
sram_cell_6t_5 inst_cell_153_116 (.BL(BL116),.BLN(BLN116),.WL(WL153));
sram_cell_6t_5 inst_cell_153_117 (.BL(BL117),.BLN(BLN117),.WL(WL153));
sram_cell_6t_5 inst_cell_153_118 (.BL(BL118),.BLN(BLN118),.WL(WL153));
sram_cell_6t_5 inst_cell_153_119 (.BL(BL119),.BLN(BLN119),.WL(WL153));
sram_cell_6t_5 inst_cell_153_120 (.BL(BL120),.BLN(BLN120),.WL(WL153));
sram_cell_6t_5 inst_cell_153_121 (.BL(BL121),.BLN(BLN121),.WL(WL153));
sram_cell_6t_5 inst_cell_153_122 (.BL(BL122),.BLN(BLN122),.WL(WL153));
sram_cell_6t_5 inst_cell_153_123 (.BL(BL123),.BLN(BLN123),.WL(WL153));
sram_cell_6t_5 inst_cell_153_124 (.BL(BL124),.BLN(BLN124),.WL(WL153));
sram_cell_6t_5 inst_cell_153_125 (.BL(BL125),.BLN(BLN125),.WL(WL153));
sram_cell_6t_5 inst_cell_153_126 (.BL(BL126),.BLN(BLN126),.WL(WL153));
sram_cell_6t_5 inst_cell_153_127 (.BL(BL127),.BLN(BLN127),.WL(WL153));
sram_cell_6t_5 inst_cell_154_0 (.BL(BL0),.BLN(BLN0),.WL(WL154));
sram_cell_6t_5 inst_cell_154_1 (.BL(BL1),.BLN(BLN1),.WL(WL154));
sram_cell_6t_5 inst_cell_154_2 (.BL(BL2),.BLN(BLN2),.WL(WL154));
sram_cell_6t_5 inst_cell_154_3 (.BL(BL3),.BLN(BLN3),.WL(WL154));
sram_cell_6t_5 inst_cell_154_4 (.BL(BL4),.BLN(BLN4),.WL(WL154));
sram_cell_6t_5 inst_cell_154_5 (.BL(BL5),.BLN(BLN5),.WL(WL154));
sram_cell_6t_5 inst_cell_154_6 (.BL(BL6),.BLN(BLN6),.WL(WL154));
sram_cell_6t_5 inst_cell_154_7 (.BL(BL7),.BLN(BLN7),.WL(WL154));
sram_cell_6t_5 inst_cell_154_8 (.BL(BL8),.BLN(BLN8),.WL(WL154));
sram_cell_6t_5 inst_cell_154_9 (.BL(BL9),.BLN(BLN9),.WL(WL154));
sram_cell_6t_5 inst_cell_154_10 (.BL(BL10),.BLN(BLN10),.WL(WL154));
sram_cell_6t_5 inst_cell_154_11 (.BL(BL11),.BLN(BLN11),.WL(WL154));
sram_cell_6t_5 inst_cell_154_12 (.BL(BL12),.BLN(BLN12),.WL(WL154));
sram_cell_6t_5 inst_cell_154_13 (.BL(BL13),.BLN(BLN13),.WL(WL154));
sram_cell_6t_5 inst_cell_154_14 (.BL(BL14),.BLN(BLN14),.WL(WL154));
sram_cell_6t_5 inst_cell_154_15 (.BL(BL15),.BLN(BLN15),.WL(WL154));
sram_cell_6t_5 inst_cell_154_16 (.BL(BL16),.BLN(BLN16),.WL(WL154));
sram_cell_6t_5 inst_cell_154_17 (.BL(BL17),.BLN(BLN17),.WL(WL154));
sram_cell_6t_5 inst_cell_154_18 (.BL(BL18),.BLN(BLN18),.WL(WL154));
sram_cell_6t_5 inst_cell_154_19 (.BL(BL19),.BLN(BLN19),.WL(WL154));
sram_cell_6t_5 inst_cell_154_20 (.BL(BL20),.BLN(BLN20),.WL(WL154));
sram_cell_6t_5 inst_cell_154_21 (.BL(BL21),.BLN(BLN21),.WL(WL154));
sram_cell_6t_5 inst_cell_154_22 (.BL(BL22),.BLN(BLN22),.WL(WL154));
sram_cell_6t_5 inst_cell_154_23 (.BL(BL23),.BLN(BLN23),.WL(WL154));
sram_cell_6t_5 inst_cell_154_24 (.BL(BL24),.BLN(BLN24),.WL(WL154));
sram_cell_6t_5 inst_cell_154_25 (.BL(BL25),.BLN(BLN25),.WL(WL154));
sram_cell_6t_5 inst_cell_154_26 (.BL(BL26),.BLN(BLN26),.WL(WL154));
sram_cell_6t_5 inst_cell_154_27 (.BL(BL27),.BLN(BLN27),.WL(WL154));
sram_cell_6t_5 inst_cell_154_28 (.BL(BL28),.BLN(BLN28),.WL(WL154));
sram_cell_6t_5 inst_cell_154_29 (.BL(BL29),.BLN(BLN29),.WL(WL154));
sram_cell_6t_5 inst_cell_154_30 (.BL(BL30),.BLN(BLN30),.WL(WL154));
sram_cell_6t_5 inst_cell_154_31 (.BL(BL31),.BLN(BLN31),.WL(WL154));
sram_cell_6t_5 inst_cell_154_32 (.BL(BL32),.BLN(BLN32),.WL(WL154));
sram_cell_6t_5 inst_cell_154_33 (.BL(BL33),.BLN(BLN33),.WL(WL154));
sram_cell_6t_5 inst_cell_154_34 (.BL(BL34),.BLN(BLN34),.WL(WL154));
sram_cell_6t_5 inst_cell_154_35 (.BL(BL35),.BLN(BLN35),.WL(WL154));
sram_cell_6t_5 inst_cell_154_36 (.BL(BL36),.BLN(BLN36),.WL(WL154));
sram_cell_6t_5 inst_cell_154_37 (.BL(BL37),.BLN(BLN37),.WL(WL154));
sram_cell_6t_5 inst_cell_154_38 (.BL(BL38),.BLN(BLN38),.WL(WL154));
sram_cell_6t_5 inst_cell_154_39 (.BL(BL39),.BLN(BLN39),.WL(WL154));
sram_cell_6t_5 inst_cell_154_40 (.BL(BL40),.BLN(BLN40),.WL(WL154));
sram_cell_6t_5 inst_cell_154_41 (.BL(BL41),.BLN(BLN41),.WL(WL154));
sram_cell_6t_5 inst_cell_154_42 (.BL(BL42),.BLN(BLN42),.WL(WL154));
sram_cell_6t_5 inst_cell_154_43 (.BL(BL43),.BLN(BLN43),.WL(WL154));
sram_cell_6t_5 inst_cell_154_44 (.BL(BL44),.BLN(BLN44),.WL(WL154));
sram_cell_6t_5 inst_cell_154_45 (.BL(BL45),.BLN(BLN45),.WL(WL154));
sram_cell_6t_5 inst_cell_154_46 (.BL(BL46),.BLN(BLN46),.WL(WL154));
sram_cell_6t_5 inst_cell_154_47 (.BL(BL47),.BLN(BLN47),.WL(WL154));
sram_cell_6t_5 inst_cell_154_48 (.BL(BL48),.BLN(BLN48),.WL(WL154));
sram_cell_6t_5 inst_cell_154_49 (.BL(BL49),.BLN(BLN49),.WL(WL154));
sram_cell_6t_5 inst_cell_154_50 (.BL(BL50),.BLN(BLN50),.WL(WL154));
sram_cell_6t_5 inst_cell_154_51 (.BL(BL51),.BLN(BLN51),.WL(WL154));
sram_cell_6t_5 inst_cell_154_52 (.BL(BL52),.BLN(BLN52),.WL(WL154));
sram_cell_6t_5 inst_cell_154_53 (.BL(BL53),.BLN(BLN53),.WL(WL154));
sram_cell_6t_5 inst_cell_154_54 (.BL(BL54),.BLN(BLN54),.WL(WL154));
sram_cell_6t_5 inst_cell_154_55 (.BL(BL55),.BLN(BLN55),.WL(WL154));
sram_cell_6t_5 inst_cell_154_56 (.BL(BL56),.BLN(BLN56),.WL(WL154));
sram_cell_6t_5 inst_cell_154_57 (.BL(BL57),.BLN(BLN57),.WL(WL154));
sram_cell_6t_5 inst_cell_154_58 (.BL(BL58),.BLN(BLN58),.WL(WL154));
sram_cell_6t_5 inst_cell_154_59 (.BL(BL59),.BLN(BLN59),.WL(WL154));
sram_cell_6t_5 inst_cell_154_60 (.BL(BL60),.BLN(BLN60),.WL(WL154));
sram_cell_6t_5 inst_cell_154_61 (.BL(BL61),.BLN(BLN61),.WL(WL154));
sram_cell_6t_5 inst_cell_154_62 (.BL(BL62),.BLN(BLN62),.WL(WL154));
sram_cell_6t_5 inst_cell_154_63 (.BL(BL63),.BLN(BLN63),.WL(WL154));
sram_cell_6t_5 inst_cell_154_64 (.BL(BL64),.BLN(BLN64),.WL(WL154));
sram_cell_6t_5 inst_cell_154_65 (.BL(BL65),.BLN(BLN65),.WL(WL154));
sram_cell_6t_5 inst_cell_154_66 (.BL(BL66),.BLN(BLN66),.WL(WL154));
sram_cell_6t_5 inst_cell_154_67 (.BL(BL67),.BLN(BLN67),.WL(WL154));
sram_cell_6t_5 inst_cell_154_68 (.BL(BL68),.BLN(BLN68),.WL(WL154));
sram_cell_6t_5 inst_cell_154_69 (.BL(BL69),.BLN(BLN69),.WL(WL154));
sram_cell_6t_5 inst_cell_154_70 (.BL(BL70),.BLN(BLN70),.WL(WL154));
sram_cell_6t_5 inst_cell_154_71 (.BL(BL71),.BLN(BLN71),.WL(WL154));
sram_cell_6t_5 inst_cell_154_72 (.BL(BL72),.BLN(BLN72),.WL(WL154));
sram_cell_6t_5 inst_cell_154_73 (.BL(BL73),.BLN(BLN73),.WL(WL154));
sram_cell_6t_5 inst_cell_154_74 (.BL(BL74),.BLN(BLN74),.WL(WL154));
sram_cell_6t_5 inst_cell_154_75 (.BL(BL75),.BLN(BLN75),.WL(WL154));
sram_cell_6t_5 inst_cell_154_76 (.BL(BL76),.BLN(BLN76),.WL(WL154));
sram_cell_6t_5 inst_cell_154_77 (.BL(BL77),.BLN(BLN77),.WL(WL154));
sram_cell_6t_5 inst_cell_154_78 (.BL(BL78),.BLN(BLN78),.WL(WL154));
sram_cell_6t_5 inst_cell_154_79 (.BL(BL79),.BLN(BLN79),.WL(WL154));
sram_cell_6t_5 inst_cell_154_80 (.BL(BL80),.BLN(BLN80),.WL(WL154));
sram_cell_6t_5 inst_cell_154_81 (.BL(BL81),.BLN(BLN81),.WL(WL154));
sram_cell_6t_5 inst_cell_154_82 (.BL(BL82),.BLN(BLN82),.WL(WL154));
sram_cell_6t_5 inst_cell_154_83 (.BL(BL83),.BLN(BLN83),.WL(WL154));
sram_cell_6t_5 inst_cell_154_84 (.BL(BL84),.BLN(BLN84),.WL(WL154));
sram_cell_6t_5 inst_cell_154_85 (.BL(BL85),.BLN(BLN85),.WL(WL154));
sram_cell_6t_5 inst_cell_154_86 (.BL(BL86),.BLN(BLN86),.WL(WL154));
sram_cell_6t_5 inst_cell_154_87 (.BL(BL87),.BLN(BLN87),.WL(WL154));
sram_cell_6t_5 inst_cell_154_88 (.BL(BL88),.BLN(BLN88),.WL(WL154));
sram_cell_6t_5 inst_cell_154_89 (.BL(BL89),.BLN(BLN89),.WL(WL154));
sram_cell_6t_5 inst_cell_154_90 (.BL(BL90),.BLN(BLN90),.WL(WL154));
sram_cell_6t_5 inst_cell_154_91 (.BL(BL91),.BLN(BLN91),.WL(WL154));
sram_cell_6t_5 inst_cell_154_92 (.BL(BL92),.BLN(BLN92),.WL(WL154));
sram_cell_6t_5 inst_cell_154_93 (.BL(BL93),.BLN(BLN93),.WL(WL154));
sram_cell_6t_5 inst_cell_154_94 (.BL(BL94),.BLN(BLN94),.WL(WL154));
sram_cell_6t_5 inst_cell_154_95 (.BL(BL95),.BLN(BLN95),.WL(WL154));
sram_cell_6t_5 inst_cell_154_96 (.BL(BL96),.BLN(BLN96),.WL(WL154));
sram_cell_6t_5 inst_cell_154_97 (.BL(BL97),.BLN(BLN97),.WL(WL154));
sram_cell_6t_5 inst_cell_154_98 (.BL(BL98),.BLN(BLN98),.WL(WL154));
sram_cell_6t_5 inst_cell_154_99 (.BL(BL99),.BLN(BLN99),.WL(WL154));
sram_cell_6t_5 inst_cell_154_100 (.BL(BL100),.BLN(BLN100),.WL(WL154));
sram_cell_6t_5 inst_cell_154_101 (.BL(BL101),.BLN(BLN101),.WL(WL154));
sram_cell_6t_5 inst_cell_154_102 (.BL(BL102),.BLN(BLN102),.WL(WL154));
sram_cell_6t_5 inst_cell_154_103 (.BL(BL103),.BLN(BLN103),.WL(WL154));
sram_cell_6t_5 inst_cell_154_104 (.BL(BL104),.BLN(BLN104),.WL(WL154));
sram_cell_6t_5 inst_cell_154_105 (.BL(BL105),.BLN(BLN105),.WL(WL154));
sram_cell_6t_5 inst_cell_154_106 (.BL(BL106),.BLN(BLN106),.WL(WL154));
sram_cell_6t_5 inst_cell_154_107 (.BL(BL107),.BLN(BLN107),.WL(WL154));
sram_cell_6t_5 inst_cell_154_108 (.BL(BL108),.BLN(BLN108),.WL(WL154));
sram_cell_6t_5 inst_cell_154_109 (.BL(BL109),.BLN(BLN109),.WL(WL154));
sram_cell_6t_5 inst_cell_154_110 (.BL(BL110),.BLN(BLN110),.WL(WL154));
sram_cell_6t_5 inst_cell_154_111 (.BL(BL111),.BLN(BLN111),.WL(WL154));
sram_cell_6t_5 inst_cell_154_112 (.BL(BL112),.BLN(BLN112),.WL(WL154));
sram_cell_6t_5 inst_cell_154_113 (.BL(BL113),.BLN(BLN113),.WL(WL154));
sram_cell_6t_5 inst_cell_154_114 (.BL(BL114),.BLN(BLN114),.WL(WL154));
sram_cell_6t_5 inst_cell_154_115 (.BL(BL115),.BLN(BLN115),.WL(WL154));
sram_cell_6t_5 inst_cell_154_116 (.BL(BL116),.BLN(BLN116),.WL(WL154));
sram_cell_6t_5 inst_cell_154_117 (.BL(BL117),.BLN(BLN117),.WL(WL154));
sram_cell_6t_5 inst_cell_154_118 (.BL(BL118),.BLN(BLN118),.WL(WL154));
sram_cell_6t_5 inst_cell_154_119 (.BL(BL119),.BLN(BLN119),.WL(WL154));
sram_cell_6t_5 inst_cell_154_120 (.BL(BL120),.BLN(BLN120),.WL(WL154));
sram_cell_6t_5 inst_cell_154_121 (.BL(BL121),.BLN(BLN121),.WL(WL154));
sram_cell_6t_5 inst_cell_154_122 (.BL(BL122),.BLN(BLN122),.WL(WL154));
sram_cell_6t_5 inst_cell_154_123 (.BL(BL123),.BLN(BLN123),.WL(WL154));
sram_cell_6t_5 inst_cell_154_124 (.BL(BL124),.BLN(BLN124),.WL(WL154));
sram_cell_6t_5 inst_cell_154_125 (.BL(BL125),.BLN(BLN125),.WL(WL154));
sram_cell_6t_5 inst_cell_154_126 (.BL(BL126),.BLN(BLN126),.WL(WL154));
sram_cell_6t_5 inst_cell_154_127 (.BL(BL127),.BLN(BLN127),.WL(WL154));
sram_cell_6t_5 inst_cell_155_0 (.BL(BL0),.BLN(BLN0),.WL(WL155));
sram_cell_6t_5 inst_cell_155_1 (.BL(BL1),.BLN(BLN1),.WL(WL155));
sram_cell_6t_5 inst_cell_155_2 (.BL(BL2),.BLN(BLN2),.WL(WL155));
sram_cell_6t_5 inst_cell_155_3 (.BL(BL3),.BLN(BLN3),.WL(WL155));
sram_cell_6t_5 inst_cell_155_4 (.BL(BL4),.BLN(BLN4),.WL(WL155));
sram_cell_6t_5 inst_cell_155_5 (.BL(BL5),.BLN(BLN5),.WL(WL155));
sram_cell_6t_5 inst_cell_155_6 (.BL(BL6),.BLN(BLN6),.WL(WL155));
sram_cell_6t_5 inst_cell_155_7 (.BL(BL7),.BLN(BLN7),.WL(WL155));
sram_cell_6t_5 inst_cell_155_8 (.BL(BL8),.BLN(BLN8),.WL(WL155));
sram_cell_6t_5 inst_cell_155_9 (.BL(BL9),.BLN(BLN9),.WL(WL155));
sram_cell_6t_5 inst_cell_155_10 (.BL(BL10),.BLN(BLN10),.WL(WL155));
sram_cell_6t_5 inst_cell_155_11 (.BL(BL11),.BLN(BLN11),.WL(WL155));
sram_cell_6t_5 inst_cell_155_12 (.BL(BL12),.BLN(BLN12),.WL(WL155));
sram_cell_6t_5 inst_cell_155_13 (.BL(BL13),.BLN(BLN13),.WL(WL155));
sram_cell_6t_5 inst_cell_155_14 (.BL(BL14),.BLN(BLN14),.WL(WL155));
sram_cell_6t_5 inst_cell_155_15 (.BL(BL15),.BLN(BLN15),.WL(WL155));
sram_cell_6t_5 inst_cell_155_16 (.BL(BL16),.BLN(BLN16),.WL(WL155));
sram_cell_6t_5 inst_cell_155_17 (.BL(BL17),.BLN(BLN17),.WL(WL155));
sram_cell_6t_5 inst_cell_155_18 (.BL(BL18),.BLN(BLN18),.WL(WL155));
sram_cell_6t_5 inst_cell_155_19 (.BL(BL19),.BLN(BLN19),.WL(WL155));
sram_cell_6t_5 inst_cell_155_20 (.BL(BL20),.BLN(BLN20),.WL(WL155));
sram_cell_6t_5 inst_cell_155_21 (.BL(BL21),.BLN(BLN21),.WL(WL155));
sram_cell_6t_5 inst_cell_155_22 (.BL(BL22),.BLN(BLN22),.WL(WL155));
sram_cell_6t_5 inst_cell_155_23 (.BL(BL23),.BLN(BLN23),.WL(WL155));
sram_cell_6t_5 inst_cell_155_24 (.BL(BL24),.BLN(BLN24),.WL(WL155));
sram_cell_6t_5 inst_cell_155_25 (.BL(BL25),.BLN(BLN25),.WL(WL155));
sram_cell_6t_5 inst_cell_155_26 (.BL(BL26),.BLN(BLN26),.WL(WL155));
sram_cell_6t_5 inst_cell_155_27 (.BL(BL27),.BLN(BLN27),.WL(WL155));
sram_cell_6t_5 inst_cell_155_28 (.BL(BL28),.BLN(BLN28),.WL(WL155));
sram_cell_6t_5 inst_cell_155_29 (.BL(BL29),.BLN(BLN29),.WL(WL155));
sram_cell_6t_5 inst_cell_155_30 (.BL(BL30),.BLN(BLN30),.WL(WL155));
sram_cell_6t_5 inst_cell_155_31 (.BL(BL31),.BLN(BLN31),.WL(WL155));
sram_cell_6t_5 inst_cell_155_32 (.BL(BL32),.BLN(BLN32),.WL(WL155));
sram_cell_6t_5 inst_cell_155_33 (.BL(BL33),.BLN(BLN33),.WL(WL155));
sram_cell_6t_5 inst_cell_155_34 (.BL(BL34),.BLN(BLN34),.WL(WL155));
sram_cell_6t_5 inst_cell_155_35 (.BL(BL35),.BLN(BLN35),.WL(WL155));
sram_cell_6t_5 inst_cell_155_36 (.BL(BL36),.BLN(BLN36),.WL(WL155));
sram_cell_6t_5 inst_cell_155_37 (.BL(BL37),.BLN(BLN37),.WL(WL155));
sram_cell_6t_5 inst_cell_155_38 (.BL(BL38),.BLN(BLN38),.WL(WL155));
sram_cell_6t_5 inst_cell_155_39 (.BL(BL39),.BLN(BLN39),.WL(WL155));
sram_cell_6t_5 inst_cell_155_40 (.BL(BL40),.BLN(BLN40),.WL(WL155));
sram_cell_6t_5 inst_cell_155_41 (.BL(BL41),.BLN(BLN41),.WL(WL155));
sram_cell_6t_5 inst_cell_155_42 (.BL(BL42),.BLN(BLN42),.WL(WL155));
sram_cell_6t_5 inst_cell_155_43 (.BL(BL43),.BLN(BLN43),.WL(WL155));
sram_cell_6t_5 inst_cell_155_44 (.BL(BL44),.BLN(BLN44),.WL(WL155));
sram_cell_6t_5 inst_cell_155_45 (.BL(BL45),.BLN(BLN45),.WL(WL155));
sram_cell_6t_5 inst_cell_155_46 (.BL(BL46),.BLN(BLN46),.WL(WL155));
sram_cell_6t_5 inst_cell_155_47 (.BL(BL47),.BLN(BLN47),.WL(WL155));
sram_cell_6t_5 inst_cell_155_48 (.BL(BL48),.BLN(BLN48),.WL(WL155));
sram_cell_6t_5 inst_cell_155_49 (.BL(BL49),.BLN(BLN49),.WL(WL155));
sram_cell_6t_5 inst_cell_155_50 (.BL(BL50),.BLN(BLN50),.WL(WL155));
sram_cell_6t_5 inst_cell_155_51 (.BL(BL51),.BLN(BLN51),.WL(WL155));
sram_cell_6t_5 inst_cell_155_52 (.BL(BL52),.BLN(BLN52),.WL(WL155));
sram_cell_6t_5 inst_cell_155_53 (.BL(BL53),.BLN(BLN53),.WL(WL155));
sram_cell_6t_5 inst_cell_155_54 (.BL(BL54),.BLN(BLN54),.WL(WL155));
sram_cell_6t_5 inst_cell_155_55 (.BL(BL55),.BLN(BLN55),.WL(WL155));
sram_cell_6t_5 inst_cell_155_56 (.BL(BL56),.BLN(BLN56),.WL(WL155));
sram_cell_6t_5 inst_cell_155_57 (.BL(BL57),.BLN(BLN57),.WL(WL155));
sram_cell_6t_5 inst_cell_155_58 (.BL(BL58),.BLN(BLN58),.WL(WL155));
sram_cell_6t_5 inst_cell_155_59 (.BL(BL59),.BLN(BLN59),.WL(WL155));
sram_cell_6t_5 inst_cell_155_60 (.BL(BL60),.BLN(BLN60),.WL(WL155));
sram_cell_6t_5 inst_cell_155_61 (.BL(BL61),.BLN(BLN61),.WL(WL155));
sram_cell_6t_5 inst_cell_155_62 (.BL(BL62),.BLN(BLN62),.WL(WL155));
sram_cell_6t_5 inst_cell_155_63 (.BL(BL63),.BLN(BLN63),.WL(WL155));
sram_cell_6t_5 inst_cell_155_64 (.BL(BL64),.BLN(BLN64),.WL(WL155));
sram_cell_6t_5 inst_cell_155_65 (.BL(BL65),.BLN(BLN65),.WL(WL155));
sram_cell_6t_5 inst_cell_155_66 (.BL(BL66),.BLN(BLN66),.WL(WL155));
sram_cell_6t_5 inst_cell_155_67 (.BL(BL67),.BLN(BLN67),.WL(WL155));
sram_cell_6t_5 inst_cell_155_68 (.BL(BL68),.BLN(BLN68),.WL(WL155));
sram_cell_6t_5 inst_cell_155_69 (.BL(BL69),.BLN(BLN69),.WL(WL155));
sram_cell_6t_5 inst_cell_155_70 (.BL(BL70),.BLN(BLN70),.WL(WL155));
sram_cell_6t_5 inst_cell_155_71 (.BL(BL71),.BLN(BLN71),.WL(WL155));
sram_cell_6t_5 inst_cell_155_72 (.BL(BL72),.BLN(BLN72),.WL(WL155));
sram_cell_6t_5 inst_cell_155_73 (.BL(BL73),.BLN(BLN73),.WL(WL155));
sram_cell_6t_5 inst_cell_155_74 (.BL(BL74),.BLN(BLN74),.WL(WL155));
sram_cell_6t_5 inst_cell_155_75 (.BL(BL75),.BLN(BLN75),.WL(WL155));
sram_cell_6t_5 inst_cell_155_76 (.BL(BL76),.BLN(BLN76),.WL(WL155));
sram_cell_6t_5 inst_cell_155_77 (.BL(BL77),.BLN(BLN77),.WL(WL155));
sram_cell_6t_5 inst_cell_155_78 (.BL(BL78),.BLN(BLN78),.WL(WL155));
sram_cell_6t_5 inst_cell_155_79 (.BL(BL79),.BLN(BLN79),.WL(WL155));
sram_cell_6t_5 inst_cell_155_80 (.BL(BL80),.BLN(BLN80),.WL(WL155));
sram_cell_6t_5 inst_cell_155_81 (.BL(BL81),.BLN(BLN81),.WL(WL155));
sram_cell_6t_5 inst_cell_155_82 (.BL(BL82),.BLN(BLN82),.WL(WL155));
sram_cell_6t_5 inst_cell_155_83 (.BL(BL83),.BLN(BLN83),.WL(WL155));
sram_cell_6t_5 inst_cell_155_84 (.BL(BL84),.BLN(BLN84),.WL(WL155));
sram_cell_6t_5 inst_cell_155_85 (.BL(BL85),.BLN(BLN85),.WL(WL155));
sram_cell_6t_5 inst_cell_155_86 (.BL(BL86),.BLN(BLN86),.WL(WL155));
sram_cell_6t_5 inst_cell_155_87 (.BL(BL87),.BLN(BLN87),.WL(WL155));
sram_cell_6t_5 inst_cell_155_88 (.BL(BL88),.BLN(BLN88),.WL(WL155));
sram_cell_6t_5 inst_cell_155_89 (.BL(BL89),.BLN(BLN89),.WL(WL155));
sram_cell_6t_5 inst_cell_155_90 (.BL(BL90),.BLN(BLN90),.WL(WL155));
sram_cell_6t_5 inst_cell_155_91 (.BL(BL91),.BLN(BLN91),.WL(WL155));
sram_cell_6t_5 inst_cell_155_92 (.BL(BL92),.BLN(BLN92),.WL(WL155));
sram_cell_6t_5 inst_cell_155_93 (.BL(BL93),.BLN(BLN93),.WL(WL155));
sram_cell_6t_5 inst_cell_155_94 (.BL(BL94),.BLN(BLN94),.WL(WL155));
sram_cell_6t_5 inst_cell_155_95 (.BL(BL95),.BLN(BLN95),.WL(WL155));
sram_cell_6t_5 inst_cell_155_96 (.BL(BL96),.BLN(BLN96),.WL(WL155));
sram_cell_6t_5 inst_cell_155_97 (.BL(BL97),.BLN(BLN97),.WL(WL155));
sram_cell_6t_5 inst_cell_155_98 (.BL(BL98),.BLN(BLN98),.WL(WL155));
sram_cell_6t_5 inst_cell_155_99 (.BL(BL99),.BLN(BLN99),.WL(WL155));
sram_cell_6t_5 inst_cell_155_100 (.BL(BL100),.BLN(BLN100),.WL(WL155));
sram_cell_6t_5 inst_cell_155_101 (.BL(BL101),.BLN(BLN101),.WL(WL155));
sram_cell_6t_5 inst_cell_155_102 (.BL(BL102),.BLN(BLN102),.WL(WL155));
sram_cell_6t_5 inst_cell_155_103 (.BL(BL103),.BLN(BLN103),.WL(WL155));
sram_cell_6t_5 inst_cell_155_104 (.BL(BL104),.BLN(BLN104),.WL(WL155));
sram_cell_6t_5 inst_cell_155_105 (.BL(BL105),.BLN(BLN105),.WL(WL155));
sram_cell_6t_5 inst_cell_155_106 (.BL(BL106),.BLN(BLN106),.WL(WL155));
sram_cell_6t_5 inst_cell_155_107 (.BL(BL107),.BLN(BLN107),.WL(WL155));
sram_cell_6t_5 inst_cell_155_108 (.BL(BL108),.BLN(BLN108),.WL(WL155));
sram_cell_6t_5 inst_cell_155_109 (.BL(BL109),.BLN(BLN109),.WL(WL155));
sram_cell_6t_5 inst_cell_155_110 (.BL(BL110),.BLN(BLN110),.WL(WL155));
sram_cell_6t_5 inst_cell_155_111 (.BL(BL111),.BLN(BLN111),.WL(WL155));
sram_cell_6t_5 inst_cell_155_112 (.BL(BL112),.BLN(BLN112),.WL(WL155));
sram_cell_6t_5 inst_cell_155_113 (.BL(BL113),.BLN(BLN113),.WL(WL155));
sram_cell_6t_5 inst_cell_155_114 (.BL(BL114),.BLN(BLN114),.WL(WL155));
sram_cell_6t_5 inst_cell_155_115 (.BL(BL115),.BLN(BLN115),.WL(WL155));
sram_cell_6t_5 inst_cell_155_116 (.BL(BL116),.BLN(BLN116),.WL(WL155));
sram_cell_6t_5 inst_cell_155_117 (.BL(BL117),.BLN(BLN117),.WL(WL155));
sram_cell_6t_5 inst_cell_155_118 (.BL(BL118),.BLN(BLN118),.WL(WL155));
sram_cell_6t_5 inst_cell_155_119 (.BL(BL119),.BLN(BLN119),.WL(WL155));
sram_cell_6t_5 inst_cell_155_120 (.BL(BL120),.BLN(BLN120),.WL(WL155));
sram_cell_6t_5 inst_cell_155_121 (.BL(BL121),.BLN(BLN121),.WL(WL155));
sram_cell_6t_5 inst_cell_155_122 (.BL(BL122),.BLN(BLN122),.WL(WL155));
sram_cell_6t_5 inst_cell_155_123 (.BL(BL123),.BLN(BLN123),.WL(WL155));
sram_cell_6t_5 inst_cell_155_124 (.BL(BL124),.BLN(BLN124),.WL(WL155));
sram_cell_6t_5 inst_cell_155_125 (.BL(BL125),.BLN(BLN125),.WL(WL155));
sram_cell_6t_5 inst_cell_155_126 (.BL(BL126),.BLN(BLN126),.WL(WL155));
sram_cell_6t_5 inst_cell_155_127 (.BL(BL127),.BLN(BLN127),.WL(WL155));
sram_cell_6t_5 inst_cell_156_0 (.BL(BL0),.BLN(BLN0),.WL(WL156));
sram_cell_6t_5 inst_cell_156_1 (.BL(BL1),.BLN(BLN1),.WL(WL156));
sram_cell_6t_5 inst_cell_156_2 (.BL(BL2),.BLN(BLN2),.WL(WL156));
sram_cell_6t_5 inst_cell_156_3 (.BL(BL3),.BLN(BLN3),.WL(WL156));
sram_cell_6t_5 inst_cell_156_4 (.BL(BL4),.BLN(BLN4),.WL(WL156));
sram_cell_6t_5 inst_cell_156_5 (.BL(BL5),.BLN(BLN5),.WL(WL156));
sram_cell_6t_5 inst_cell_156_6 (.BL(BL6),.BLN(BLN6),.WL(WL156));
sram_cell_6t_5 inst_cell_156_7 (.BL(BL7),.BLN(BLN7),.WL(WL156));
sram_cell_6t_5 inst_cell_156_8 (.BL(BL8),.BLN(BLN8),.WL(WL156));
sram_cell_6t_5 inst_cell_156_9 (.BL(BL9),.BLN(BLN9),.WL(WL156));
sram_cell_6t_5 inst_cell_156_10 (.BL(BL10),.BLN(BLN10),.WL(WL156));
sram_cell_6t_5 inst_cell_156_11 (.BL(BL11),.BLN(BLN11),.WL(WL156));
sram_cell_6t_5 inst_cell_156_12 (.BL(BL12),.BLN(BLN12),.WL(WL156));
sram_cell_6t_5 inst_cell_156_13 (.BL(BL13),.BLN(BLN13),.WL(WL156));
sram_cell_6t_5 inst_cell_156_14 (.BL(BL14),.BLN(BLN14),.WL(WL156));
sram_cell_6t_5 inst_cell_156_15 (.BL(BL15),.BLN(BLN15),.WL(WL156));
sram_cell_6t_5 inst_cell_156_16 (.BL(BL16),.BLN(BLN16),.WL(WL156));
sram_cell_6t_5 inst_cell_156_17 (.BL(BL17),.BLN(BLN17),.WL(WL156));
sram_cell_6t_5 inst_cell_156_18 (.BL(BL18),.BLN(BLN18),.WL(WL156));
sram_cell_6t_5 inst_cell_156_19 (.BL(BL19),.BLN(BLN19),.WL(WL156));
sram_cell_6t_5 inst_cell_156_20 (.BL(BL20),.BLN(BLN20),.WL(WL156));
sram_cell_6t_5 inst_cell_156_21 (.BL(BL21),.BLN(BLN21),.WL(WL156));
sram_cell_6t_5 inst_cell_156_22 (.BL(BL22),.BLN(BLN22),.WL(WL156));
sram_cell_6t_5 inst_cell_156_23 (.BL(BL23),.BLN(BLN23),.WL(WL156));
sram_cell_6t_5 inst_cell_156_24 (.BL(BL24),.BLN(BLN24),.WL(WL156));
sram_cell_6t_5 inst_cell_156_25 (.BL(BL25),.BLN(BLN25),.WL(WL156));
sram_cell_6t_5 inst_cell_156_26 (.BL(BL26),.BLN(BLN26),.WL(WL156));
sram_cell_6t_5 inst_cell_156_27 (.BL(BL27),.BLN(BLN27),.WL(WL156));
sram_cell_6t_5 inst_cell_156_28 (.BL(BL28),.BLN(BLN28),.WL(WL156));
sram_cell_6t_5 inst_cell_156_29 (.BL(BL29),.BLN(BLN29),.WL(WL156));
sram_cell_6t_5 inst_cell_156_30 (.BL(BL30),.BLN(BLN30),.WL(WL156));
sram_cell_6t_5 inst_cell_156_31 (.BL(BL31),.BLN(BLN31),.WL(WL156));
sram_cell_6t_5 inst_cell_156_32 (.BL(BL32),.BLN(BLN32),.WL(WL156));
sram_cell_6t_5 inst_cell_156_33 (.BL(BL33),.BLN(BLN33),.WL(WL156));
sram_cell_6t_5 inst_cell_156_34 (.BL(BL34),.BLN(BLN34),.WL(WL156));
sram_cell_6t_5 inst_cell_156_35 (.BL(BL35),.BLN(BLN35),.WL(WL156));
sram_cell_6t_5 inst_cell_156_36 (.BL(BL36),.BLN(BLN36),.WL(WL156));
sram_cell_6t_5 inst_cell_156_37 (.BL(BL37),.BLN(BLN37),.WL(WL156));
sram_cell_6t_5 inst_cell_156_38 (.BL(BL38),.BLN(BLN38),.WL(WL156));
sram_cell_6t_5 inst_cell_156_39 (.BL(BL39),.BLN(BLN39),.WL(WL156));
sram_cell_6t_5 inst_cell_156_40 (.BL(BL40),.BLN(BLN40),.WL(WL156));
sram_cell_6t_5 inst_cell_156_41 (.BL(BL41),.BLN(BLN41),.WL(WL156));
sram_cell_6t_5 inst_cell_156_42 (.BL(BL42),.BLN(BLN42),.WL(WL156));
sram_cell_6t_5 inst_cell_156_43 (.BL(BL43),.BLN(BLN43),.WL(WL156));
sram_cell_6t_5 inst_cell_156_44 (.BL(BL44),.BLN(BLN44),.WL(WL156));
sram_cell_6t_5 inst_cell_156_45 (.BL(BL45),.BLN(BLN45),.WL(WL156));
sram_cell_6t_5 inst_cell_156_46 (.BL(BL46),.BLN(BLN46),.WL(WL156));
sram_cell_6t_5 inst_cell_156_47 (.BL(BL47),.BLN(BLN47),.WL(WL156));
sram_cell_6t_5 inst_cell_156_48 (.BL(BL48),.BLN(BLN48),.WL(WL156));
sram_cell_6t_5 inst_cell_156_49 (.BL(BL49),.BLN(BLN49),.WL(WL156));
sram_cell_6t_5 inst_cell_156_50 (.BL(BL50),.BLN(BLN50),.WL(WL156));
sram_cell_6t_5 inst_cell_156_51 (.BL(BL51),.BLN(BLN51),.WL(WL156));
sram_cell_6t_5 inst_cell_156_52 (.BL(BL52),.BLN(BLN52),.WL(WL156));
sram_cell_6t_5 inst_cell_156_53 (.BL(BL53),.BLN(BLN53),.WL(WL156));
sram_cell_6t_5 inst_cell_156_54 (.BL(BL54),.BLN(BLN54),.WL(WL156));
sram_cell_6t_5 inst_cell_156_55 (.BL(BL55),.BLN(BLN55),.WL(WL156));
sram_cell_6t_5 inst_cell_156_56 (.BL(BL56),.BLN(BLN56),.WL(WL156));
sram_cell_6t_5 inst_cell_156_57 (.BL(BL57),.BLN(BLN57),.WL(WL156));
sram_cell_6t_5 inst_cell_156_58 (.BL(BL58),.BLN(BLN58),.WL(WL156));
sram_cell_6t_5 inst_cell_156_59 (.BL(BL59),.BLN(BLN59),.WL(WL156));
sram_cell_6t_5 inst_cell_156_60 (.BL(BL60),.BLN(BLN60),.WL(WL156));
sram_cell_6t_5 inst_cell_156_61 (.BL(BL61),.BLN(BLN61),.WL(WL156));
sram_cell_6t_5 inst_cell_156_62 (.BL(BL62),.BLN(BLN62),.WL(WL156));
sram_cell_6t_5 inst_cell_156_63 (.BL(BL63),.BLN(BLN63),.WL(WL156));
sram_cell_6t_5 inst_cell_156_64 (.BL(BL64),.BLN(BLN64),.WL(WL156));
sram_cell_6t_5 inst_cell_156_65 (.BL(BL65),.BLN(BLN65),.WL(WL156));
sram_cell_6t_5 inst_cell_156_66 (.BL(BL66),.BLN(BLN66),.WL(WL156));
sram_cell_6t_5 inst_cell_156_67 (.BL(BL67),.BLN(BLN67),.WL(WL156));
sram_cell_6t_5 inst_cell_156_68 (.BL(BL68),.BLN(BLN68),.WL(WL156));
sram_cell_6t_5 inst_cell_156_69 (.BL(BL69),.BLN(BLN69),.WL(WL156));
sram_cell_6t_5 inst_cell_156_70 (.BL(BL70),.BLN(BLN70),.WL(WL156));
sram_cell_6t_5 inst_cell_156_71 (.BL(BL71),.BLN(BLN71),.WL(WL156));
sram_cell_6t_5 inst_cell_156_72 (.BL(BL72),.BLN(BLN72),.WL(WL156));
sram_cell_6t_5 inst_cell_156_73 (.BL(BL73),.BLN(BLN73),.WL(WL156));
sram_cell_6t_5 inst_cell_156_74 (.BL(BL74),.BLN(BLN74),.WL(WL156));
sram_cell_6t_5 inst_cell_156_75 (.BL(BL75),.BLN(BLN75),.WL(WL156));
sram_cell_6t_5 inst_cell_156_76 (.BL(BL76),.BLN(BLN76),.WL(WL156));
sram_cell_6t_5 inst_cell_156_77 (.BL(BL77),.BLN(BLN77),.WL(WL156));
sram_cell_6t_5 inst_cell_156_78 (.BL(BL78),.BLN(BLN78),.WL(WL156));
sram_cell_6t_5 inst_cell_156_79 (.BL(BL79),.BLN(BLN79),.WL(WL156));
sram_cell_6t_5 inst_cell_156_80 (.BL(BL80),.BLN(BLN80),.WL(WL156));
sram_cell_6t_5 inst_cell_156_81 (.BL(BL81),.BLN(BLN81),.WL(WL156));
sram_cell_6t_5 inst_cell_156_82 (.BL(BL82),.BLN(BLN82),.WL(WL156));
sram_cell_6t_5 inst_cell_156_83 (.BL(BL83),.BLN(BLN83),.WL(WL156));
sram_cell_6t_5 inst_cell_156_84 (.BL(BL84),.BLN(BLN84),.WL(WL156));
sram_cell_6t_5 inst_cell_156_85 (.BL(BL85),.BLN(BLN85),.WL(WL156));
sram_cell_6t_5 inst_cell_156_86 (.BL(BL86),.BLN(BLN86),.WL(WL156));
sram_cell_6t_5 inst_cell_156_87 (.BL(BL87),.BLN(BLN87),.WL(WL156));
sram_cell_6t_5 inst_cell_156_88 (.BL(BL88),.BLN(BLN88),.WL(WL156));
sram_cell_6t_5 inst_cell_156_89 (.BL(BL89),.BLN(BLN89),.WL(WL156));
sram_cell_6t_5 inst_cell_156_90 (.BL(BL90),.BLN(BLN90),.WL(WL156));
sram_cell_6t_5 inst_cell_156_91 (.BL(BL91),.BLN(BLN91),.WL(WL156));
sram_cell_6t_5 inst_cell_156_92 (.BL(BL92),.BLN(BLN92),.WL(WL156));
sram_cell_6t_5 inst_cell_156_93 (.BL(BL93),.BLN(BLN93),.WL(WL156));
sram_cell_6t_5 inst_cell_156_94 (.BL(BL94),.BLN(BLN94),.WL(WL156));
sram_cell_6t_5 inst_cell_156_95 (.BL(BL95),.BLN(BLN95),.WL(WL156));
sram_cell_6t_5 inst_cell_156_96 (.BL(BL96),.BLN(BLN96),.WL(WL156));
sram_cell_6t_5 inst_cell_156_97 (.BL(BL97),.BLN(BLN97),.WL(WL156));
sram_cell_6t_5 inst_cell_156_98 (.BL(BL98),.BLN(BLN98),.WL(WL156));
sram_cell_6t_5 inst_cell_156_99 (.BL(BL99),.BLN(BLN99),.WL(WL156));
sram_cell_6t_5 inst_cell_156_100 (.BL(BL100),.BLN(BLN100),.WL(WL156));
sram_cell_6t_5 inst_cell_156_101 (.BL(BL101),.BLN(BLN101),.WL(WL156));
sram_cell_6t_5 inst_cell_156_102 (.BL(BL102),.BLN(BLN102),.WL(WL156));
sram_cell_6t_5 inst_cell_156_103 (.BL(BL103),.BLN(BLN103),.WL(WL156));
sram_cell_6t_5 inst_cell_156_104 (.BL(BL104),.BLN(BLN104),.WL(WL156));
sram_cell_6t_5 inst_cell_156_105 (.BL(BL105),.BLN(BLN105),.WL(WL156));
sram_cell_6t_5 inst_cell_156_106 (.BL(BL106),.BLN(BLN106),.WL(WL156));
sram_cell_6t_5 inst_cell_156_107 (.BL(BL107),.BLN(BLN107),.WL(WL156));
sram_cell_6t_5 inst_cell_156_108 (.BL(BL108),.BLN(BLN108),.WL(WL156));
sram_cell_6t_5 inst_cell_156_109 (.BL(BL109),.BLN(BLN109),.WL(WL156));
sram_cell_6t_5 inst_cell_156_110 (.BL(BL110),.BLN(BLN110),.WL(WL156));
sram_cell_6t_5 inst_cell_156_111 (.BL(BL111),.BLN(BLN111),.WL(WL156));
sram_cell_6t_5 inst_cell_156_112 (.BL(BL112),.BLN(BLN112),.WL(WL156));
sram_cell_6t_5 inst_cell_156_113 (.BL(BL113),.BLN(BLN113),.WL(WL156));
sram_cell_6t_5 inst_cell_156_114 (.BL(BL114),.BLN(BLN114),.WL(WL156));
sram_cell_6t_5 inst_cell_156_115 (.BL(BL115),.BLN(BLN115),.WL(WL156));
sram_cell_6t_5 inst_cell_156_116 (.BL(BL116),.BLN(BLN116),.WL(WL156));
sram_cell_6t_5 inst_cell_156_117 (.BL(BL117),.BLN(BLN117),.WL(WL156));
sram_cell_6t_5 inst_cell_156_118 (.BL(BL118),.BLN(BLN118),.WL(WL156));
sram_cell_6t_5 inst_cell_156_119 (.BL(BL119),.BLN(BLN119),.WL(WL156));
sram_cell_6t_5 inst_cell_156_120 (.BL(BL120),.BLN(BLN120),.WL(WL156));
sram_cell_6t_5 inst_cell_156_121 (.BL(BL121),.BLN(BLN121),.WL(WL156));
sram_cell_6t_5 inst_cell_156_122 (.BL(BL122),.BLN(BLN122),.WL(WL156));
sram_cell_6t_5 inst_cell_156_123 (.BL(BL123),.BLN(BLN123),.WL(WL156));
sram_cell_6t_5 inst_cell_156_124 (.BL(BL124),.BLN(BLN124),.WL(WL156));
sram_cell_6t_5 inst_cell_156_125 (.BL(BL125),.BLN(BLN125),.WL(WL156));
sram_cell_6t_5 inst_cell_156_126 (.BL(BL126),.BLN(BLN126),.WL(WL156));
sram_cell_6t_5 inst_cell_156_127 (.BL(BL127),.BLN(BLN127),.WL(WL156));
sram_cell_6t_5 inst_cell_157_0 (.BL(BL0),.BLN(BLN0),.WL(WL157));
sram_cell_6t_5 inst_cell_157_1 (.BL(BL1),.BLN(BLN1),.WL(WL157));
sram_cell_6t_5 inst_cell_157_2 (.BL(BL2),.BLN(BLN2),.WL(WL157));
sram_cell_6t_5 inst_cell_157_3 (.BL(BL3),.BLN(BLN3),.WL(WL157));
sram_cell_6t_5 inst_cell_157_4 (.BL(BL4),.BLN(BLN4),.WL(WL157));
sram_cell_6t_5 inst_cell_157_5 (.BL(BL5),.BLN(BLN5),.WL(WL157));
sram_cell_6t_5 inst_cell_157_6 (.BL(BL6),.BLN(BLN6),.WL(WL157));
sram_cell_6t_5 inst_cell_157_7 (.BL(BL7),.BLN(BLN7),.WL(WL157));
sram_cell_6t_5 inst_cell_157_8 (.BL(BL8),.BLN(BLN8),.WL(WL157));
sram_cell_6t_5 inst_cell_157_9 (.BL(BL9),.BLN(BLN9),.WL(WL157));
sram_cell_6t_5 inst_cell_157_10 (.BL(BL10),.BLN(BLN10),.WL(WL157));
sram_cell_6t_5 inst_cell_157_11 (.BL(BL11),.BLN(BLN11),.WL(WL157));
sram_cell_6t_5 inst_cell_157_12 (.BL(BL12),.BLN(BLN12),.WL(WL157));
sram_cell_6t_5 inst_cell_157_13 (.BL(BL13),.BLN(BLN13),.WL(WL157));
sram_cell_6t_5 inst_cell_157_14 (.BL(BL14),.BLN(BLN14),.WL(WL157));
sram_cell_6t_5 inst_cell_157_15 (.BL(BL15),.BLN(BLN15),.WL(WL157));
sram_cell_6t_5 inst_cell_157_16 (.BL(BL16),.BLN(BLN16),.WL(WL157));
sram_cell_6t_5 inst_cell_157_17 (.BL(BL17),.BLN(BLN17),.WL(WL157));
sram_cell_6t_5 inst_cell_157_18 (.BL(BL18),.BLN(BLN18),.WL(WL157));
sram_cell_6t_5 inst_cell_157_19 (.BL(BL19),.BLN(BLN19),.WL(WL157));
sram_cell_6t_5 inst_cell_157_20 (.BL(BL20),.BLN(BLN20),.WL(WL157));
sram_cell_6t_5 inst_cell_157_21 (.BL(BL21),.BLN(BLN21),.WL(WL157));
sram_cell_6t_5 inst_cell_157_22 (.BL(BL22),.BLN(BLN22),.WL(WL157));
sram_cell_6t_5 inst_cell_157_23 (.BL(BL23),.BLN(BLN23),.WL(WL157));
sram_cell_6t_5 inst_cell_157_24 (.BL(BL24),.BLN(BLN24),.WL(WL157));
sram_cell_6t_5 inst_cell_157_25 (.BL(BL25),.BLN(BLN25),.WL(WL157));
sram_cell_6t_5 inst_cell_157_26 (.BL(BL26),.BLN(BLN26),.WL(WL157));
sram_cell_6t_5 inst_cell_157_27 (.BL(BL27),.BLN(BLN27),.WL(WL157));
sram_cell_6t_5 inst_cell_157_28 (.BL(BL28),.BLN(BLN28),.WL(WL157));
sram_cell_6t_5 inst_cell_157_29 (.BL(BL29),.BLN(BLN29),.WL(WL157));
sram_cell_6t_5 inst_cell_157_30 (.BL(BL30),.BLN(BLN30),.WL(WL157));
sram_cell_6t_5 inst_cell_157_31 (.BL(BL31),.BLN(BLN31),.WL(WL157));
sram_cell_6t_5 inst_cell_157_32 (.BL(BL32),.BLN(BLN32),.WL(WL157));
sram_cell_6t_5 inst_cell_157_33 (.BL(BL33),.BLN(BLN33),.WL(WL157));
sram_cell_6t_5 inst_cell_157_34 (.BL(BL34),.BLN(BLN34),.WL(WL157));
sram_cell_6t_5 inst_cell_157_35 (.BL(BL35),.BLN(BLN35),.WL(WL157));
sram_cell_6t_5 inst_cell_157_36 (.BL(BL36),.BLN(BLN36),.WL(WL157));
sram_cell_6t_5 inst_cell_157_37 (.BL(BL37),.BLN(BLN37),.WL(WL157));
sram_cell_6t_5 inst_cell_157_38 (.BL(BL38),.BLN(BLN38),.WL(WL157));
sram_cell_6t_5 inst_cell_157_39 (.BL(BL39),.BLN(BLN39),.WL(WL157));
sram_cell_6t_5 inst_cell_157_40 (.BL(BL40),.BLN(BLN40),.WL(WL157));
sram_cell_6t_5 inst_cell_157_41 (.BL(BL41),.BLN(BLN41),.WL(WL157));
sram_cell_6t_5 inst_cell_157_42 (.BL(BL42),.BLN(BLN42),.WL(WL157));
sram_cell_6t_5 inst_cell_157_43 (.BL(BL43),.BLN(BLN43),.WL(WL157));
sram_cell_6t_5 inst_cell_157_44 (.BL(BL44),.BLN(BLN44),.WL(WL157));
sram_cell_6t_5 inst_cell_157_45 (.BL(BL45),.BLN(BLN45),.WL(WL157));
sram_cell_6t_5 inst_cell_157_46 (.BL(BL46),.BLN(BLN46),.WL(WL157));
sram_cell_6t_5 inst_cell_157_47 (.BL(BL47),.BLN(BLN47),.WL(WL157));
sram_cell_6t_5 inst_cell_157_48 (.BL(BL48),.BLN(BLN48),.WL(WL157));
sram_cell_6t_5 inst_cell_157_49 (.BL(BL49),.BLN(BLN49),.WL(WL157));
sram_cell_6t_5 inst_cell_157_50 (.BL(BL50),.BLN(BLN50),.WL(WL157));
sram_cell_6t_5 inst_cell_157_51 (.BL(BL51),.BLN(BLN51),.WL(WL157));
sram_cell_6t_5 inst_cell_157_52 (.BL(BL52),.BLN(BLN52),.WL(WL157));
sram_cell_6t_5 inst_cell_157_53 (.BL(BL53),.BLN(BLN53),.WL(WL157));
sram_cell_6t_5 inst_cell_157_54 (.BL(BL54),.BLN(BLN54),.WL(WL157));
sram_cell_6t_5 inst_cell_157_55 (.BL(BL55),.BLN(BLN55),.WL(WL157));
sram_cell_6t_5 inst_cell_157_56 (.BL(BL56),.BLN(BLN56),.WL(WL157));
sram_cell_6t_5 inst_cell_157_57 (.BL(BL57),.BLN(BLN57),.WL(WL157));
sram_cell_6t_5 inst_cell_157_58 (.BL(BL58),.BLN(BLN58),.WL(WL157));
sram_cell_6t_5 inst_cell_157_59 (.BL(BL59),.BLN(BLN59),.WL(WL157));
sram_cell_6t_5 inst_cell_157_60 (.BL(BL60),.BLN(BLN60),.WL(WL157));
sram_cell_6t_5 inst_cell_157_61 (.BL(BL61),.BLN(BLN61),.WL(WL157));
sram_cell_6t_5 inst_cell_157_62 (.BL(BL62),.BLN(BLN62),.WL(WL157));
sram_cell_6t_5 inst_cell_157_63 (.BL(BL63),.BLN(BLN63),.WL(WL157));
sram_cell_6t_5 inst_cell_157_64 (.BL(BL64),.BLN(BLN64),.WL(WL157));
sram_cell_6t_5 inst_cell_157_65 (.BL(BL65),.BLN(BLN65),.WL(WL157));
sram_cell_6t_5 inst_cell_157_66 (.BL(BL66),.BLN(BLN66),.WL(WL157));
sram_cell_6t_5 inst_cell_157_67 (.BL(BL67),.BLN(BLN67),.WL(WL157));
sram_cell_6t_5 inst_cell_157_68 (.BL(BL68),.BLN(BLN68),.WL(WL157));
sram_cell_6t_5 inst_cell_157_69 (.BL(BL69),.BLN(BLN69),.WL(WL157));
sram_cell_6t_5 inst_cell_157_70 (.BL(BL70),.BLN(BLN70),.WL(WL157));
sram_cell_6t_5 inst_cell_157_71 (.BL(BL71),.BLN(BLN71),.WL(WL157));
sram_cell_6t_5 inst_cell_157_72 (.BL(BL72),.BLN(BLN72),.WL(WL157));
sram_cell_6t_5 inst_cell_157_73 (.BL(BL73),.BLN(BLN73),.WL(WL157));
sram_cell_6t_5 inst_cell_157_74 (.BL(BL74),.BLN(BLN74),.WL(WL157));
sram_cell_6t_5 inst_cell_157_75 (.BL(BL75),.BLN(BLN75),.WL(WL157));
sram_cell_6t_5 inst_cell_157_76 (.BL(BL76),.BLN(BLN76),.WL(WL157));
sram_cell_6t_5 inst_cell_157_77 (.BL(BL77),.BLN(BLN77),.WL(WL157));
sram_cell_6t_5 inst_cell_157_78 (.BL(BL78),.BLN(BLN78),.WL(WL157));
sram_cell_6t_5 inst_cell_157_79 (.BL(BL79),.BLN(BLN79),.WL(WL157));
sram_cell_6t_5 inst_cell_157_80 (.BL(BL80),.BLN(BLN80),.WL(WL157));
sram_cell_6t_5 inst_cell_157_81 (.BL(BL81),.BLN(BLN81),.WL(WL157));
sram_cell_6t_5 inst_cell_157_82 (.BL(BL82),.BLN(BLN82),.WL(WL157));
sram_cell_6t_5 inst_cell_157_83 (.BL(BL83),.BLN(BLN83),.WL(WL157));
sram_cell_6t_5 inst_cell_157_84 (.BL(BL84),.BLN(BLN84),.WL(WL157));
sram_cell_6t_5 inst_cell_157_85 (.BL(BL85),.BLN(BLN85),.WL(WL157));
sram_cell_6t_5 inst_cell_157_86 (.BL(BL86),.BLN(BLN86),.WL(WL157));
sram_cell_6t_5 inst_cell_157_87 (.BL(BL87),.BLN(BLN87),.WL(WL157));
sram_cell_6t_5 inst_cell_157_88 (.BL(BL88),.BLN(BLN88),.WL(WL157));
sram_cell_6t_5 inst_cell_157_89 (.BL(BL89),.BLN(BLN89),.WL(WL157));
sram_cell_6t_5 inst_cell_157_90 (.BL(BL90),.BLN(BLN90),.WL(WL157));
sram_cell_6t_5 inst_cell_157_91 (.BL(BL91),.BLN(BLN91),.WL(WL157));
sram_cell_6t_5 inst_cell_157_92 (.BL(BL92),.BLN(BLN92),.WL(WL157));
sram_cell_6t_5 inst_cell_157_93 (.BL(BL93),.BLN(BLN93),.WL(WL157));
sram_cell_6t_5 inst_cell_157_94 (.BL(BL94),.BLN(BLN94),.WL(WL157));
sram_cell_6t_5 inst_cell_157_95 (.BL(BL95),.BLN(BLN95),.WL(WL157));
sram_cell_6t_5 inst_cell_157_96 (.BL(BL96),.BLN(BLN96),.WL(WL157));
sram_cell_6t_5 inst_cell_157_97 (.BL(BL97),.BLN(BLN97),.WL(WL157));
sram_cell_6t_5 inst_cell_157_98 (.BL(BL98),.BLN(BLN98),.WL(WL157));
sram_cell_6t_5 inst_cell_157_99 (.BL(BL99),.BLN(BLN99),.WL(WL157));
sram_cell_6t_5 inst_cell_157_100 (.BL(BL100),.BLN(BLN100),.WL(WL157));
sram_cell_6t_5 inst_cell_157_101 (.BL(BL101),.BLN(BLN101),.WL(WL157));
sram_cell_6t_5 inst_cell_157_102 (.BL(BL102),.BLN(BLN102),.WL(WL157));
sram_cell_6t_5 inst_cell_157_103 (.BL(BL103),.BLN(BLN103),.WL(WL157));
sram_cell_6t_5 inst_cell_157_104 (.BL(BL104),.BLN(BLN104),.WL(WL157));
sram_cell_6t_5 inst_cell_157_105 (.BL(BL105),.BLN(BLN105),.WL(WL157));
sram_cell_6t_5 inst_cell_157_106 (.BL(BL106),.BLN(BLN106),.WL(WL157));
sram_cell_6t_5 inst_cell_157_107 (.BL(BL107),.BLN(BLN107),.WL(WL157));
sram_cell_6t_5 inst_cell_157_108 (.BL(BL108),.BLN(BLN108),.WL(WL157));
sram_cell_6t_5 inst_cell_157_109 (.BL(BL109),.BLN(BLN109),.WL(WL157));
sram_cell_6t_5 inst_cell_157_110 (.BL(BL110),.BLN(BLN110),.WL(WL157));
sram_cell_6t_5 inst_cell_157_111 (.BL(BL111),.BLN(BLN111),.WL(WL157));
sram_cell_6t_5 inst_cell_157_112 (.BL(BL112),.BLN(BLN112),.WL(WL157));
sram_cell_6t_5 inst_cell_157_113 (.BL(BL113),.BLN(BLN113),.WL(WL157));
sram_cell_6t_5 inst_cell_157_114 (.BL(BL114),.BLN(BLN114),.WL(WL157));
sram_cell_6t_5 inst_cell_157_115 (.BL(BL115),.BLN(BLN115),.WL(WL157));
sram_cell_6t_5 inst_cell_157_116 (.BL(BL116),.BLN(BLN116),.WL(WL157));
sram_cell_6t_5 inst_cell_157_117 (.BL(BL117),.BLN(BLN117),.WL(WL157));
sram_cell_6t_5 inst_cell_157_118 (.BL(BL118),.BLN(BLN118),.WL(WL157));
sram_cell_6t_5 inst_cell_157_119 (.BL(BL119),.BLN(BLN119),.WL(WL157));
sram_cell_6t_5 inst_cell_157_120 (.BL(BL120),.BLN(BLN120),.WL(WL157));
sram_cell_6t_5 inst_cell_157_121 (.BL(BL121),.BLN(BLN121),.WL(WL157));
sram_cell_6t_5 inst_cell_157_122 (.BL(BL122),.BLN(BLN122),.WL(WL157));
sram_cell_6t_5 inst_cell_157_123 (.BL(BL123),.BLN(BLN123),.WL(WL157));
sram_cell_6t_5 inst_cell_157_124 (.BL(BL124),.BLN(BLN124),.WL(WL157));
sram_cell_6t_5 inst_cell_157_125 (.BL(BL125),.BLN(BLN125),.WL(WL157));
sram_cell_6t_5 inst_cell_157_126 (.BL(BL126),.BLN(BLN126),.WL(WL157));
sram_cell_6t_5 inst_cell_157_127 (.BL(BL127),.BLN(BLN127),.WL(WL157));
sram_cell_6t_5 inst_cell_158_0 (.BL(BL0),.BLN(BLN0),.WL(WL158));
sram_cell_6t_5 inst_cell_158_1 (.BL(BL1),.BLN(BLN1),.WL(WL158));
sram_cell_6t_5 inst_cell_158_2 (.BL(BL2),.BLN(BLN2),.WL(WL158));
sram_cell_6t_5 inst_cell_158_3 (.BL(BL3),.BLN(BLN3),.WL(WL158));
sram_cell_6t_5 inst_cell_158_4 (.BL(BL4),.BLN(BLN4),.WL(WL158));
sram_cell_6t_5 inst_cell_158_5 (.BL(BL5),.BLN(BLN5),.WL(WL158));
sram_cell_6t_5 inst_cell_158_6 (.BL(BL6),.BLN(BLN6),.WL(WL158));
sram_cell_6t_5 inst_cell_158_7 (.BL(BL7),.BLN(BLN7),.WL(WL158));
sram_cell_6t_5 inst_cell_158_8 (.BL(BL8),.BLN(BLN8),.WL(WL158));
sram_cell_6t_5 inst_cell_158_9 (.BL(BL9),.BLN(BLN9),.WL(WL158));
sram_cell_6t_5 inst_cell_158_10 (.BL(BL10),.BLN(BLN10),.WL(WL158));
sram_cell_6t_5 inst_cell_158_11 (.BL(BL11),.BLN(BLN11),.WL(WL158));
sram_cell_6t_5 inst_cell_158_12 (.BL(BL12),.BLN(BLN12),.WL(WL158));
sram_cell_6t_5 inst_cell_158_13 (.BL(BL13),.BLN(BLN13),.WL(WL158));
sram_cell_6t_5 inst_cell_158_14 (.BL(BL14),.BLN(BLN14),.WL(WL158));
sram_cell_6t_5 inst_cell_158_15 (.BL(BL15),.BLN(BLN15),.WL(WL158));
sram_cell_6t_5 inst_cell_158_16 (.BL(BL16),.BLN(BLN16),.WL(WL158));
sram_cell_6t_5 inst_cell_158_17 (.BL(BL17),.BLN(BLN17),.WL(WL158));
sram_cell_6t_5 inst_cell_158_18 (.BL(BL18),.BLN(BLN18),.WL(WL158));
sram_cell_6t_5 inst_cell_158_19 (.BL(BL19),.BLN(BLN19),.WL(WL158));
sram_cell_6t_5 inst_cell_158_20 (.BL(BL20),.BLN(BLN20),.WL(WL158));
sram_cell_6t_5 inst_cell_158_21 (.BL(BL21),.BLN(BLN21),.WL(WL158));
sram_cell_6t_5 inst_cell_158_22 (.BL(BL22),.BLN(BLN22),.WL(WL158));
sram_cell_6t_5 inst_cell_158_23 (.BL(BL23),.BLN(BLN23),.WL(WL158));
sram_cell_6t_5 inst_cell_158_24 (.BL(BL24),.BLN(BLN24),.WL(WL158));
sram_cell_6t_5 inst_cell_158_25 (.BL(BL25),.BLN(BLN25),.WL(WL158));
sram_cell_6t_5 inst_cell_158_26 (.BL(BL26),.BLN(BLN26),.WL(WL158));
sram_cell_6t_5 inst_cell_158_27 (.BL(BL27),.BLN(BLN27),.WL(WL158));
sram_cell_6t_5 inst_cell_158_28 (.BL(BL28),.BLN(BLN28),.WL(WL158));
sram_cell_6t_5 inst_cell_158_29 (.BL(BL29),.BLN(BLN29),.WL(WL158));
sram_cell_6t_5 inst_cell_158_30 (.BL(BL30),.BLN(BLN30),.WL(WL158));
sram_cell_6t_5 inst_cell_158_31 (.BL(BL31),.BLN(BLN31),.WL(WL158));
sram_cell_6t_5 inst_cell_158_32 (.BL(BL32),.BLN(BLN32),.WL(WL158));
sram_cell_6t_5 inst_cell_158_33 (.BL(BL33),.BLN(BLN33),.WL(WL158));
sram_cell_6t_5 inst_cell_158_34 (.BL(BL34),.BLN(BLN34),.WL(WL158));
sram_cell_6t_5 inst_cell_158_35 (.BL(BL35),.BLN(BLN35),.WL(WL158));
sram_cell_6t_5 inst_cell_158_36 (.BL(BL36),.BLN(BLN36),.WL(WL158));
sram_cell_6t_5 inst_cell_158_37 (.BL(BL37),.BLN(BLN37),.WL(WL158));
sram_cell_6t_5 inst_cell_158_38 (.BL(BL38),.BLN(BLN38),.WL(WL158));
sram_cell_6t_5 inst_cell_158_39 (.BL(BL39),.BLN(BLN39),.WL(WL158));
sram_cell_6t_5 inst_cell_158_40 (.BL(BL40),.BLN(BLN40),.WL(WL158));
sram_cell_6t_5 inst_cell_158_41 (.BL(BL41),.BLN(BLN41),.WL(WL158));
sram_cell_6t_5 inst_cell_158_42 (.BL(BL42),.BLN(BLN42),.WL(WL158));
sram_cell_6t_5 inst_cell_158_43 (.BL(BL43),.BLN(BLN43),.WL(WL158));
sram_cell_6t_5 inst_cell_158_44 (.BL(BL44),.BLN(BLN44),.WL(WL158));
sram_cell_6t_5 inst_cell_158_45 (.BL(BL45),.BLN(BLN45),.WL(WL158));
sram_cell_6t_5 inst_cell_158_46 (.BL(BL46),.BLN(BLN46),.WL(WL158));
sram_cell_6t_5 inst_cell_158_47 (.BL(BL47),.BLN(BLN47),.WL(WL158));
sram_cell_6t_5 inst_cell_158_48 (.BL(BL48),.BLN(BLN48),.WL(WL158));
sram_cell_6t_5 inst_cell_158_49 (.BL(BL49),.BLN(BLN49),.WL(WL158));
sram_cell_6t_5 inst_cell_158_50 (.BL(BL50),.BLN(BLN50),.WL(WL158));
sram_cell_6t_5 inst_cell_158_51 (.BL(BL51),.BLN(BLN51),.WL(WL158));
sram_cell_6t_5 inst_cell_158_52 (.BL(BL52),.BLN(BLN52),.WL(WL158));
sram_cell_6t_5 inst_cell_158_53 (.BL(BL53),.BLN(BLN53),.WL(WL158));
sram_cell_6t_5 inst_cell_158_54 (.BL(BL54),.BLN(BLN54),.WL(WL158));
sram_cell_6t_5 inst_cell_158_55 (.BL(BL55),.BLN(BLN55),.WL(WL158));
sram_cell_6t_5 inst_cell_158_56 (.BL(BL56),.BLN(BLN56),.WL(WL158));
sram_cell_6t_5 inst_cell_158_57 (.BL(BL57),.BLN(BLN57),.WL(WL158));
sram_cell_6t_5 inst_cell_158_58 (.BL(BL58),.BLN(BLN58),.WL(WL158));
sram_cell_6t_5 inst_cell_158_59 (.BL(BL59),.BLN(BLN59),.WL(WL158));
sram_cell_6t_5 inst_cell_158_60 (.BL(BL60),.BLN(BLN60),.WL(WL158));
sram_cell_6t_5 inst_cell_158_61 (.BL(BL61),.BLN(BLN61),.WL(WL158));
sram_cell_6t_5 inst_cell_158_62 (.BL(BL62),.BLN(BLN62),.WL(WL158));
sram_cell_6t_5 inst_cell_158_63 (.BL(BL63),.BLN(BLN63),.WL(WL158));
sram_cell_6t_5 inst_cell_158_64 (.BL(BL64),.BLN(BLN64),.WL(WL158));
sram_cell_6t_5 inst_cell_158_65 (.BL(BL65),.BLN(BLN65),.WL(WL158));
sram_cell_6t_5 inst_cell_158_66 (.BL(BL66),.BLN(BLN66),.WL(WL158));
sram_cell_6t_5 inst_cell_158_67 (.BL(BL67),.BLN(BLN67),.WL(WL158));
sram_cell_6t_5 inst_cell_158_68 (.BL(BL68),.BLN(BLN68),.WL(WL158));
sram_cell_6t_5 inst_cell_158_69 (.BL(BL69),.BLN(BLN69),.WL(WL158));
sram_cell_6t_5 inst_cell_158_70 (.BL(BL70),.BLN(BLN70),.WL(WL158));
sram_cell_6t_5 inst_cell_158_71 (.BL(BL71),.BLN(BLN71),.WL(WL158));
sram_cell_6t_5 inst_cell_158_72 (.BL(BL72),.BLN(BLN72),.WL(WL158));
sram_cell_6t_5 inst_cell_158_73 (.BL(BL73),.BLN(BLN73),.WL(WL158));
sram_cell_6t_5 inst_cell_158_74 (.BL(BL74),.BLN(BLN74),.WL(WL158));
sram_cell_6t_5 inst_cell_158_75 (.BL(BL75),.BLN(BLN75),.WL(WL158));
sram_cell_6t_5 inst_cell_158_76 (.BL(BL76),.BLN(BLN76),.WL(WL158));
sram_cell_6t_5 inst_cell_158_77 (.BL(BL77),.BLN(BLN77),.WL(WL158));
sram_cell_6t_5 inst_cell_158_78 (.BL(BL78),.BLN(BLN78),.WL(WL158));
sram_cell_6t_5 inst_cell_158_79 (.BL(BL79),.BLN(BLN79),.WL(WL158));
sram_cell_6t_5 inst_cell_158_80 (.BL(BL80),.BLN(BLN80),.WL(WL158));
sram_cell_6t_5 inst_cell_158_81 (.BL(BL81),.BLN(BLN81),.WL(WL158));
sram_cell_6t_5 inst_cell_158_82 (.BL(BL82),.BLN(BLN82),.WL(WL158));
sram_cell_6t_5 inst_cell_158_83 (.BL(BL83),.BLN(BLN83),.WL(WL158));
sram_cell_6t_5 inst_cell_158_84 (.BL(BL84),.BLN(BLN84),.WL(WL158));
sram_cell_6t_5 inst_cell_158_85 (.BL(BL85),.BLN(BLN85),.WL(WL158));
sram_cell_6t_5 inst_cell_158_86 (.BL(BL86),.BLN(BLN86),.WL(WL158));
sram_cell_6t_5 inst_cell_158_87 (.BL(BL87),.BLN(BLN87),.WL(WL158));
sram_cell_6t_5 inst_cell_158_88 (.BL(BL88),.BLN(BLN88),.WL(WL158));
sram_cell_6t_5 inst_cell_158_89 (.BL(BL89),.BLN(BLN89),.WL(WL158));
sram_cell_6t_5 inst_cell_158_90 (.BL(BL90),.BLN(BLN90),.WL(WL158));
sram_cell_6t_5 inst_cell_158_91 (.BL(BL91),.BLN(BLN91),.WL(WL158));
sram_cell_6t_5 inst_cell_158_92 (.BL(BL92),.BLN(BLN92),.WL(WL158));
sram_cell_6t_5 inst_cell_158_93 (.BL(BL93),.BLN(BLN93),.WL(WL158));
sram_cell_6t_5 inst_cell_158_94 (.BL(BL94),.BLN(BLN94),.WL(WL158));
sram_cell_6t_5 inst_cell_158_95 (.BL(BL95),.BLN(BLN95),.WL(WL158));
sram_cell_6t_5 inst_cell_158_96 (.BL(BL96),.BLN(BLN96),.WL(WL158));
sram_cell_6t_5 inst_cell_158_97 (.BL(BL97),.BLN(BLN97),.WL(WL158));
sram_cell_6t_5 inst_cell_158_98 (.BL(BL98),.BLN(BLN98),.WL(WL158));
sram_cell_6t_5 inst_cell_158_99 (.BL(BL99),.BLN(BLN99),.WL(WL158));
sram_cell_6t_5 inst_cell_158_100 (.BL(BL100),.BLN(BLN100),.WL(WL158));
sram_cell_6t_5 inst_cell_158_101 (.BL(BL101),.BLN(BLN101),.WL(WL158));
sram_cell_6t_5 inst_cell_158_102 (.BL(BL102),.BLN(BLN102),.WL(WL158));
sram_cell_6t_5 inst_cell_158_103 (.BL(BL103),.BLN(BLN103),.WL(WL158));
sram_cell_6t_5 inst_cell_158_104 (.BL(BL104),.BLN(BLN104),.WL(WL158));
sram_cell_6t_5 inst_cell_158_105 (.BL(BL105),.BLN(BLN105),.WL(WL158));
sram_cell_6t_5 inst_cell_158_106 (.BL(BL106),.BLN(BLN106),.WL(WL158));
sram_cell_6t_5 inst_cell_158_107 (.BL(BL107),.BLN(BLN107),.WL(WL158));
sram_cell_6t_5 inst_cell_158_108 (.BL(BL108),.BLN(BLN108),.WL(WL158));
sram_cell_6t_5 inst_cell_158_109 (.BL(BL109),.BLN(BLN109),.WL(WL158));
sram_cell_6t_5 inst_cell_158_110 (.BL(BL110),.BLN(BLN110),.WL(WL158));
sram_cell_6t_5 inst_cell_158_111 (.BL(BL111),.BLN(BLN111),.WL(WL158));
sram_cell_6t_5 inst_cell_158_112 (.BL(BL112),.BLN(BLN112),.WL(WL158));
sram_cell_6t_5 inst_cell_158_113 (.BL(BL113),.BLN(BLN113),.WL(WL158));
sram_cell_6t_5 inst_cell_158_114 (.BL(BL114),.BLN(BLN114),.WL(WL158));
sram_cell_6t_5 inst_cell_158_115 (.BL(BL115),.BLN(BLN115),.WL(WL158));
sram_cell_6t_5 inst_cell_158_116 (.BL(BL116),.BLN(BLN116),.WL(WL158));
sram_cell_6t_5 inst_cell_158_117 (.BL(BL117),.BLN(BLN117),.WL(WL158));
sram_cell_6t_5 inst_cell_158_118 (.BL(BL118),.BLN(BLN118),.WL(WL158));
sram_cell_6t_5 inst_cell_158_119 (.BL(BL119),.BLN(BLN119),.WL(WL158));
sram_cell_6t_5 inst_cell_158_120 (.BL(BL120),.BLN(BLN120),.WL(WL158));
sram_cell_6t_5 inst_cell_158_121 (.BL(BL121),.BLN(BLN121),.WL(WL158));
sram_cell_6t_5 inst_cell_158_122 (.BL(BL122),.BLN(BLN122),.WL(WL158));
sram_cell_6t_5 inst_cell_158_123 (.BL(BL123),.BLN(BLN123),.WL(WL158));
sram_cell_6t_5 inst_cell_158_124 (.BL(BL124),.BLN(BLN124),.WL(WL158));
sram_cell_6t_5 inst_cell_158_125 (.BL(BL125),.BLN(BLN125),.WL(WL158));
sram_cell_6t_5 inst_cell_158_126 (.BL(BL126),.BLN(BLN126),.WL(WL158));
sram_cell_6t_5 inst_cell_158_127 (.BL(BL127),.BLN(BLN127),.WL(WL158));
sram_cell_6t_5 inst_cell_159_0 (.BL(BL0),.BLN(BLN0),.WL(WL159));
sram_cell_6t_5 inst_cell_159_1 (.BL(BL1),.BLN(BLN1),.WL(WL159));
sram_cell_6t_5 inst_cell_159_2 (.BL(BL2),.BLN(BLN2),.WL(WL159));
sram_cell_6t_5 inst_cell_159_3 (.BL(BL3),.BLN(BLN3),.WL(WL159));
sram_cell_6t_5 inst_cell_159_4 (.BL(BL4),.BLN(BLN4),.WL(WL159));
sram_cell_6t_5 inst_cell_159_5 (.BL(BL5),.BLN(BLN5),.WL(WL159));
sram_cell_6t_5 inst_cell_159_6 (.BL(BL6),.BLN(BLN6),.WL(WL159));
sram_cell_6t_5 inst_cell_159_7 (.BL(BL7),.BLN(BLN7),.WL(WL159));
sram_cell_6t_5 inst_cell_159_8 (.BL(BL8),.BLN(BLN8),.WL(WL159));
sram_cell_6t_5 inst_cell_159_9 (.BL(BL9),.BLN(BLN9),.WL(WL159));
sram_cell_6t_5 inst_cell_159_10 (.BL(BL10),.BLN(BLN10),.WL(WL159));
sram_cell_6t_5 inst_cell_159_11 (.BL(BL11),.BLN(BLN11),.WL(WL159));
sram_cell_6t_5 inst_cell_159_12 (.BL(BL12),.BLN(BLN12),.WL(WL159));
sram_cell_6t_5 inst_cell_159_13 (.BL(BL13),.BLN(BLN13),.WL(WL159));
sram_cell_6t_5 inst_cell_159_14 (.BL(BL14),.BLN(BLN14),.WL(WL159));
sram_cell_6t_5 inst_cell_159_15 (.BL(BL15),.BLN(BLN15),.WL(WL159));
sram_cell_6t_5 inst_cell_159_16 (.BL(BL16),.BLN(BLN16),.WL(WL159));
sram_cell_6t_5 inst_cell_159_17 (.BL(BL17),.BLN(BLN17),.WL(WL159));
sram_cell_6t_5 inst_cell_159_18 (.BL(BL18),.BLN(BLN18),.WL(WL159));
sram_cell_6t_5 inst_cell_159_19 (.BL(BL19),.BLN(BLN19),.WL(WL159));
sram_cell_6t_5 inst_cell_159_20 (.BL(BL20),.BLN(BLN20),.WL(WL159));
sram_cell_6t_5 inst_cell_159_21 (.BL(BL21),.BLN(BLN21),.WL(WL159));
sram_cell_6t_5 inst_cell_159_22 (.BL(BL22),.BLN(BLN22),.WL(WL159));
sram_cell_6t_5 inst_cell_159_23 (.BL(BL23),.BLN(BLN23),.WL(WL159));
sram_cell_6t_5 inst_cell_159_24 (.BL(BL24),.BLN(BLN24),.WL(WL159));
sram_cell_6t_5 inst_cell_159_25 (.BL(BL25),.BLN(BLN25),.WL(WL159));
sram_cell_6t_5 inst_cell_159_26 (.BL(BL26),.BLN(BLN26),.WL(WL159));
sram_cell_6t_5 inst_cell_159_27 (.BL(BL27),.BLN(BLN27),.WL(WL159));
sram_cell_6t_5 inst_cell_159_28 (.BL(BL28),.BLN(BLN28),.WL(WL159));
sram_cell_6t_5 inst_cell_159_29 (.BL(BL29),.BLN(BLN29),.WL(WL159));
sram_cell_6t_5 inst_cell_159_30 (.BL(BL30),.BLN(BLN30),.WL(WL159));
sram_cell_6t_5 inst_cell_159_31 (.BL(BL31),.BLN(BLN31),.WL(WL159));
sram_cell_6t_5 inst_cell_159_32 (.BL(BL32),.BLN(BLN32),.WL(WL159));
sram_cell_6t_5 inst_cell_159_33 (.BL(BL33),.BLN(BLN33),.WL(WL159));
sram_cell_6t_5 inst_cell_159_34 (.BL(BL34),.BLN(BLN34),.WL(WL159));
sram_cell_6t_5 inst_cell_159_35 (.BL(BL35),.BLN(BLN35),.WL(WL159));
sram_cell_6t_5 inst_cell_159_36 (.BL(BL36),.BLN(BLN36),.WL(WL159));
sram_cell_6t_5 inst_cell_159_37 (.BL(BL37),.BLN(BLN37),.WL(WL159));
sram_cell_6t_5 inst_cell_159_38 (.BL(BL38),.BLN(BLN38),.WL(WL159));
sram_cell_6t_5 inst_cell_159_39 (.BL(BL39),.BLN(BLN39),.WL(WL159));
sram_cell_6t_5 inst_cell_159_40 (.BL(BL40),.BLN(BLN40),.WL(WL159));
sram_cell_6t_5 inst_cell_159_41 (.BL(BL41),.BLN(BLN41),.WL(WL159));
sram_cell_6t_5 inst_cell_159_42 (.BL(BL42),.BLN(BLN42),.WL(WL159));
sram_cell_6t_5 inst_cell_159_43 (.BL(BL43),.BLN(BLN43),.WL(WL159));
sram_cell_6t_5 inst_cell_159_44 (.BL(BL44),.BLN(BLN44),.WL(WL159));
sram_cell_6t_5 inst_cell_159_45 (.BL(BL45),.BLN(BLN45),.WL(WL159));
sram_cell_6t_5 inst_cell_159_46 (.BL(BL46),.BLN(BLN46),.WL(WL159));
sram_cell_6t_5 inst_cell_159_47 (.BL(BL47),.BLN(BLN47),.WL(WL159));
sram_cell_6t_5 inst_cell_159_48 (.BL(BL48),.BLN(BLN48),.WL(WL159));
sram_cell_6t_5 inst_cell_159_49 (.BL(BL49),.BLN(BLN49),.WL(WL159));
sram_cell_6t_5 inst_cell_159_50 (.BL(BL50),.BLN(BLN50),.WL(WL159));
sram_cell_6t_5 inst_cell_159_51 (.BL(BL51),.BLN(BLN51),.WL(WL159));
sram_cell_6t_5 inst_cell_159_52 (.BL(BL52),.BLN(BLN52),.WL(WL159));
sram_cell_6t_5 inst_cell_159_53 (.BL(BL53),.BLN(BLN53),.WL(WL159));
sram_cell_6t_5 inst_cell_159_54 (.BL(BL54),.BLN(BLN54),.WL(WL159));
sram_cell_6t_5 inst_cell_159_55 (.BL(BL55),.BLN(BLN55),.WL(WL159));
sram_cell_6t_5 inst_cell_159_56 (.BL(BL56),.BLN(BLN56),.WL(WL159));
sram_cell_6t_5 inst_cell_159_57 (.BL(BL57),.BLN(BLN57),.WL(WL159));
sram_cell_6t_5 inst_cell_159_58 (.BL(BL58),.BLN(BLN58),.WL(WL159));
sram_cell_6t_5 inst_cell_159_59 (.BL(BL59),.BLN(BLN59),.WL(WL159));
sram_cell_6t_5 inst_cell_159_60 (.BL(BL60),.BLN(BLN60),.WL(WL159));
sram_cell_6t_5 inst_cell_159_61 (.BL(BL61),.BLN(BLN61),.WL(WL159));
sram_cell_6t_5 inst_cell_159_62 (.BL(BL62),.BLN(BLN62),.WL(WL159));
sram_cell_6t_5 inst_cell_159_63 (.BL(BL63),.BLN(BLN63),.WL(WL159));
sram_cell_6t_5 inst_cell_159_64 (.BL(BL64),.BLN(BLN64),.WL(WL159));
sram_cell_6t_5 inst_cell_159_65 (.BL(BL65),.BLN(BLN65),.WL(WL159));
sram_cell_6t_5 inst_cell_159_66 (.BL(BL66),.BLN(BLN66),.WL(WL159));
sram_cell_6t_5 inst_cell_159_67 (.BL(BL67),.BLN(BLN67),.WL(WL159));
sram_cell_6t_5 inst_cell_159_68 (.BL(BL68),.BLN(BLN68),.WL(WL159));
sram_cell_6t_5 inst_cell_159_69 (.BL(BL69),.BLN(BLN69),.WL(WL159));
sram_cell_6t_5 inst_cell_159_70 (.BL(BL70),.BLN(BLN70),.WL(WL159));
sram_cell_6t_5 inst_cell_159_71 (.BL(BL71),.BLN(BLN71),.WL(WL159));
sram_cell_6t_5 inst_cell_159_72 (.BL(BL72),.BLN(BLN72),.WL(WL159));
sram_cell_6t_5 inst_cell_159_73 (.BL(BL73),.BLN(BLN73),.WL(WL159));
sram_cell_6t_5 inst_cell_159_74 (.BL(BL74),.BLN(BLN74),.WL(WL159));
sram_cell_6t_5 inst_cell_159_75 (.BL(BL75),.BLN(BLN75),.WL(WL159));
sram_cell_6t_5 inst_cell_159_76 (.BL(BL76),.BLN(BLN76),.WL(WL159));
sram_cell_6t_5 inst_cell_159_77 (.BL(BL77),.BLN(BLN77),.WL(WL159));
sram_cell_6t_5 inst_cell_159_78 (.BL(BL78),.BLN(BLN78),.WL(WL159));
sram_cell_6t_5 inst_cell_159_79 (.BL(BL79),.BLN(BLN79),.WL(WL159));
sram_cell_6t_5 inst_cell_159_80 (.BL(BL80),.BLN(BLN80),.WL(WL159));
sram_cell_6t_5 inst_cell_159_81 (.BL(BL81),.BLN(BLN81),.WL(WL159));
sram_cell_6t_5 inst_cell_159_82 (.BL(BL82),.BLN(BLN82),.WL(WL159));
sram_cell_6t_5 inst_cell_159_83 (.BL(BL83),.BLN(BLN83),.WL(WL159));
sram_cell_6t_5 inst_cell_159_84 (.BL(BL84),.BLN(BLN84),.WL(WL159));
sram_cell_6t_5 inst_cell_159_85 (.BL(BL85),.BLN(BLN85),.WL(WL159));
sram_cell_6t_5 inst_cell_159_86 (.BL(BL86),.BLN(BLN86),.WL(WL159));
sram_cell_6t_5 inst_cell_159_87 (.BL(BL87),.BLN(BLN87),.WL(WL159));
sram_cell_6t_5 inst_cell_159_88 (.BL(BL88),.BLN(BLN88),.WL(WL159));
sram_cell_6t_5 inst_cell_159_89 (.BL(BL89),.BLN(BLN89),.WL(WL159));
sram_cell_6t_5 inst_cell_159_90 (.BL(BL90),.BLN(BLN90),.WL(WL159));
sram_cell_6t_5 inst_cell_159_91 (.BL(BL91),.BLN(BLN91),.WL(WL159));
sram_cell_6t_5 inst_cell_159_92 (.BL(BL92),.BLN(BLN92),.WL(WL159));
sram_cell_6t_5 inst_cell_159_93 (.BL(BL93),.BLN(BLN93),.WL(WL159));
sram_cell_6t_5 inst_cell_159_94 (.BL(BL94),.BLN(BLN94),.WL(WL159));
sram_cell_6t_5 inst_cell_159_95 (.BL(BL95),.BLN(BLN95),.WL(WL159));
sram_cell_6t_5 inst_cell_159_96 (.BL(BL96),.BLN(BLN96),.WL(WL159));
sram_cell_6t_5 inst_cell_159_97 (.BL(BL97),.BLN(BLN97),.WL(WL159));
sram_cell_6t_5 inst_cell_159_98 (.BL(BL98),.BLN(BLN98),.WL(WL159));
sram_cell_6t_5 inst_cell_159_99 (.BL(BL99),.BLN(BLN99),.WL(WL159));
sram_cell_6t_5 inst_cell_159_100 (.BL(BL100),.BLN(BLN100),.WL(WL159));
sram_cell_6t_5 inst_cell_159_101 (.BL(BL101),.BLN(BLN101),.WL(WL159));
sram_cell_6t_5 inst_cell_159_102 (.BL(BL102),.BLN(BLN102),.WL(WL159));
sram_cell_6t_5 inst_cell_159_103 (.BL(BL103),.BLN(BLN103),.WL(WL159));
sram_cell_6t_5 inst_cell_159_104 (.BL(BL104),.BLN(BLN104),.WL(WL159));
sram_cell_6t_5 inst_cell_159_105 (.BL(BL105),.BLN(BLN105),.WL(WL159));
sram_cell_6t_5 inst_cell_159_106 (.BL(BL106),.BLN(BLN106),.WL(WL159));
sram_cell_6t_5 inst_cell_159_107 (.BL(BL107),.BLN(BLN107),.WL(WL159));
sram_cell_6t_5 inst_cell_159_108 (.BL(BL108),.BLN(BLN108),.WL(WL159));
sram_cell_6t_5 inst_cell_159_109 (.BL(BL109),.BLN(BLN109),.WL(WL159));
sram_cell_6t_5 inst_cell_159_110 (.BL(BL110),.BLN(BLN110),.WL(WL159));
sram_cell_6t_5 inst_cell_159_111 (.BL(BL111),.BLN(BLN111),.WL(WL159));
sram_cell_6t_5 inst_cell_159_112 (.BL(BL112),.BLN(BLN112),.WL(WL159));
sram_cell_6t_5 inst_cell_159_113 (.BL(BL113),.BLN(BLN113),.WL(WL159));
sram_cell_6t_5 inst_cell_159_114 (.BL(BL114),.BLN(BLN114),.WL(WL159));
sram_cell_6t_5 inst_cell_159_115 (.BL(BL115),.BLN(BLN115),.WL(WL159));
sram_cell_6t_5 inst_cell_159_116 (.BL(BL116),.BLN(BLN116),.WL(WL159));
sram_cell_6t_5 inst_cell_159_117 (.BL(BL117),.BLN(BLN117),.WL(WL159));
sram_cell_6t_5 inst_cell_159_118 (.BL(BL118),.BLN(BLN118),.WL(WL159));
sram_cell_6t_5 inst_cell_159_119 (.BL(BL119),.BLN(BLN119),.WL(WL159));
sram_cell_6t_5 inst_cell_159_120 (.BL(BL120),.BLN(BLN120),.WL(WL159));
sram_cell_6t_5 inst_cell_159_121 (.BL(BL121),.BLN(BLN121),.WL(WL159));
sram_cell_6t_5 inst_cell_159_122 (.BL(BL122),.BLN(BLN122),.WL(WL159));
sram_cell_6t_5 inst_cell_159_123 (.BL(BL123),.BLN(BLN123),.WL(WL159));
sram_cell_6t_5 inst_cell_159_124 (.BL(BL124),.BLN(BLN124),.WL(WL159));
sram_cell_6t_5 inst_cell_159_125 (.BL(BL125),.BLN(BLN125),.WL(WL159));
sram_cell_6t_5 inst_cell_159_126 (.BL(BL126),.BLN(BLN126),.WL(WL159));
sram_cell_6t_5 inst_cell_159_127 (.BL(BL127),.BLN(BLN127),.WL(WL159));
sram_cell_6t_5 inst_cell_160_0 (.BL(BL0),.BLN(BLN0),.WL(WL160));
sram_cell_6t_5 inst_cell_160_1 (.BL(BL1),.BLN(BLN1),.WL(WL160));
sram_cell_6t_5 inst_cell_160_2 (.BL(BL2),.BLN(BLN2),.WL(WL160));
sram_cell_6t_5 inst_cell_160_3 (.BL(BL3),.BLN(BLN3),.WL(WL160));
sram_cell_6t_5 inst_cell_160_4 (.BL(BL4),.BLN(BLN4),.WL(WL160));
sram_cell_6t_5 inst_cell_160_5 (.BL(BL5),.BLN(BLN5),.WL(WL160));
sram_cell_6t_5 inst_cell_160_6 (.BL(BL6),.BLN(BLN6),.WL(WL160));
sram_cell_6t_5 inst_cell_160_7 (.BL(BL7),.BLN(BLN7),.WL(WL160));
sram_cell_6t_5 inst_cell_160_8 (.BL(BL8),.BLN(BLN8),.WL(WL160));
sram_cell_6t_5 inst_cell_160_9 (.BL(BL9),.BLN(BLN9),.WL(WL160));
sram_cell_6t_5 inst_cell_160_10 (.BL(BL10),.BLN(BLN10),.WL(WL160));
sram_cell_6t_5 inst_cell_160_11 (.BL(BL11),.BLN(BLN11),.WL(WL160));
sram_cell_6t_5 inst_cell_160_12 (.BL(BL12),.BLN(BLN12),.WL(WL160));
sram_cell_6t_5 inst_cell_160_13 (.BL(BL13),.BLN(BLN13),.WL(WL160));
sram_cell_6t_5 inst_cell_160_14 (.BL(BL14),.BLN(BLN14),.WL(WL160));
sram_cell_6t_5 inst_cell_160_15 (.BL(BL15),.BLN(BLN15),.WL(WL160));
sram_cell_6t_5 inst_cell_160_16 (.BL(BL16),.BLN(BLN16),.WL(WL160));
sram_cell_6t_5 inst_cell_160_17 (.BL(BL17),.BLN(BLN17),.WL(WL160));
sram_cell_6t_5 inst_cell_160_18 (.BL(BL18),.BLN(BLN18),.WL(WL160));
sram_cell_6t_5 inst_cell_160_19 (.BL(BL19),.BLN(BLN19),.WL(WL160));
sram_cell_6t_5 inst_cell_160_20 (.BL(BL20),.BLN(BLN20),.WL(WL160));
sram_cell_6t_5 inst_cell_160_21 (.BL(BL21),.BLN(BLN21),.WL(WL160));
sram_cell_6t_5 inst_cell_160_22 (.BL(BL22),.BLN(BLN22),.WL(WL160));
sram_cell_6t_5 inst_cell_160_23 (.BL(BL23),.BLN(BLN23),.WL(WL160));
sram_cell_6t_5 inst_cell_160_24 (.BL(BL24),.BLN(BLN24),.WL(WL160));
sram_cell_6t_5 inst_cell_160_25 (.BL(BL25),.BLN(BLN25),.WL(WL160));
sram_cell_6t_5 inst_cell_160_26 (.BL(BL26),.BLN(BLN26),.WL(WL160));
sram_cell_6t_5 inst_cell_160_27 (.BL(BL27),.BLN(BLN27),.WL(WL160));
sram_cell_6t_5 inst_cell_160_28 (.BL(BL28),.BLN(BLN28),.WL(WL160));
sram_cell_6t_5 inst_cell_160_29 (.BL(BL29),.BLN(BLN29),.WL(WL160));
sram_cell_6t_5 inst_cell_160_30 (.BL(BL30),.BLN(BLN30),.WL(WL160));
sram_cell_6t_5 inst_cell_160_31 (.BL(BL31),.BLN(BLN31),.WL(WL160));
sram_cell_6t_5 inst_cell_160_32 (.BL(BL32),.BLN(BLN32),.WL(WL160));
sram_cell_6t_5 inst_cell_160_33 (.BL(BL33),.BLN(BLN33),.WL(WL160));
sram_cell_6t_5 inst_cell_160_34 (.BL(BL34),.BLN(BLN34),.WL(WL160));
sram_cell_6t_5 inst_cell_160_35 (.BL(BL35),.BLN(BLN35),.WL(WL160));
sram_cell_6t_5 inst_cell_160_36 (.BL(BL36),.BLN(BLN36),.WL(WL160));
sram_cell_6t_5 inst_cell_160_37 (.BL(BL37),.BLN(BLN37),.WL(WL160));
sram_cell_6t_5 inst_cell_160_38 (.BL(BL38),.BLN(BLN38),.WL(WL160));
sram_cell_6t_5 inst_cell_160_39 (.BL(BL39),.BLN(BLN39),.WL(WL160));
sram_cell_6t_5 inst_cell_160_40 (.BL(BL40),.BLN(BLN40),.WL(WL160));
sram_cell_6t_5 inst_cell_160_41 (.BL(BL41),.BLN(BLN41),.WL(WL160));
sram_cell_6t_5 inst_cell_160_42 (.BL(BL42),.BLN(BLN42),.WL(WL160));
sram_cell_6t_5 inst_cell_160_43 (.BL(BL43),.BLN(BLN43),.WL(WL160));
sram_cell_6t_5 inst_cell_160_44 (.BL(BL44),.BLN(BLN44),.WL(WL160));
sram_cell_6t_5 inst_cell_160_45 (.BL(BL45),.BLN(BLN45),.WL(WL160));
sram_cell_6t_5 inst_cell_160_46 (.BL(BL46),.BLN(BLN46),.WL(WL160));
sram_cell_6t_5 inst_cell_160_47 (.BL(BL47),.BLN(BLN47),.WL(WL160));
sram_cell_6t_5 inst_cell_160_48 (.BL(BL48),.BLN(BLN48),.WL(WL160));
sram_cell_6t_5 inst_cell_160_49 (.BL(BL49),.BLN(BLN49),.WL(WL160));
sram_cell_6t_5 inst_cell_160_50 (.BL(BL50),.BLN(BLN50),.WL(WL160));
sram_cell_6t_5 inst_cell_160_51 (.BL(BL51),.BLN(BLN51),.WL(WL160));
sram_cell_6t_5 inst_cell_160_52 (.BL(BL52),.BLN(BLN52),.WL(WL160));
sram_cell_6t_5 inst_cell_160_53 (.BL(BL53),.BLN(BLN53),.WL(WL160));
sram_cell_6t_5 inst_cell_160_54 (.BL(BL54),.BLN(BLN54),.WL(WL160));
sram_cell_6t_5 inst_cell_160_55 (.BL(BL55),.BLN(BLN55),.WL(WL160));
sram_cell_6t_5 inst_cell_160_56 (.BL(BL56),.BLN(BLN56),.WL(WL160));
sram_cell_6t_5 inst_cell_160_57 (.BL(BL57),.BLN(BLN57),.WL(WL160));
sram_cell_6t_5 inst_cell_160_58 (.BL(BL58),.BLN(BLN58),.WL(WL160));
sram_cell_6t_5 inst_cell_160_59 (.BL(BL59),.BLN(BLN59),.WL(WL160));
sram_cell_6t_5 inst_cell_160_60 (.BL(BL60),.BLN(BLN60),.WL(WL160));
sram_cell_6t_5 inst_cell_160_61 (.BL(BL61),.BLN(BLN61),.WL(WL160));
sram_cell_6t_5 inst_cell_160_62 (.BL(BL62),.BLN(BLN62),.WL(WL160));
sram_cell_6t_5 inst_cell_160_63 (.BL(BL63),.BLN(BLN63),.WL(WL160));
sram_cell_6t_5 inst_cell_160_64 (.BL(BL64),.BLN(BLN64),.WL(WL160));
sram_cell_6t_5 inst_cell_160_65 (.BL(BL65),.BLN(BLN65),.WL(WL160));
sram_cell_6t_5 inst_cell_160_66 (.BL(BL66),.BLN(BLN66),.WL(WL160));
sram_cell_6t_5 inst_cell_160_67 (.BL(BL67),.BLN(BLN67),.WL(WL160));
sram_cell_6t_5 inst_cell_160_68 (.BL(BL68),.BLN(BLN68),.WL(WL160));
sram_cell_6t_5 inst_cell_160_69 (.BL(BL69),.BLN(BLN69),.WL(WL160));
sram_cell_6t_5 inst_cell_160_70 (.BL(BL70),.BLN(BLN70),.WL(WL160));
sram_cell_6t_5 inst_cell_160_71 (.BL(BL71),.BLN(BLN71),.WL(WL160));
sram_cell_6t_5 inst_cell_160_72 (.BL(BL72),.BLN(BLN72),.WL(WL160));
sram_cell_6t_5 inst_cell_160_73 (.BL(BL73),.BLN(BLN73),.WL(WL160));
sram_cell_6t_5 inst_cell_160_74 (.BL(BL74),.BLN(BLN74),.WL(WL160));
sram_cell_6t_5 inst_cell_160_75 (.BL(BL75),.BLN(BLN75),.WL(WL160));
sram_cell_6t_5 inst_cell_160_76 (.BL(BL76),.BLN(BLN76),.WL(WL160));
sram_cell_6t_5 inst_cell_160_77 (.BL(BL77),.BLN(BLN77),.WL(WL160));
sram_cell_6t_5 inst_cell_160_78 (.BL(BL78),.BLN(BLN78),.WL(WL160));
sram_cell_6t_5 inst_cell_160_79 (.BL(BL79),.BLN(BLN79),.WL(WL160));
sram_cell_6t_5 inst_cell_160_80 (.BL(BL80),.BLN(BLN80),.WL(WL160));
sram_cell_6t_5 inst_cell_160_81 (.BL(BL81),.BLN(BLN81),.WL(WL160));
sram_cell_6t_5 inst_cell_160_82 (.BL(BL82),.BLN(BLN82),.WL(WL160));
sram_cell_6t_5 inst_cell_160_83 (.BL(BL83),.BLN(BLN83),.WL(WL160));
sram_cell_6t_5 inst_cell_160_84 (.BL(BL84),.BLN(BLN84),.WL(WL160));
sram_cell_6t_5 inst_cell_160_85 (.BL(BL85),.BLN(BLN85),.WL(WL160));
sram_cell_6t_5 inst_cell_160_86 (.BL(BL86),.BLN(BLN86),.WL(WL160));
sram_cell_6t_5 inst_cell_160_87 (.BL(BL87),.BLN(BLN87),.WL(WL160));
sram_cell_6t_5 inst_cell_160_88 (.BL(BL88),.BLN(BLN88),.WL(WL160));
sram_cell_6t_5 inst_cell_160_89 (.BL(BL89),.BLN(BLN89),.WL(WL160));
sram_cell_6t_5 inst_cell_160_90 (.BL(BL90),.BLN(BLN90),.WL(WL160));
sram_cell_6t_5 inst_cell_160_91 (.BL(BL91),.BLN(BLN91),.WL(WL160));
sram_cell_6t_5 inst_cell_160_92 (.BL(BL92),.BLN(BLN92),.WL(WL160));
sram_cell_6t_5 inst_cell_160_93 (.BL(BL93),.BLN(BLN93),.WL(WL160));
sram_cell_6t_5 inst_cell_160_94 (.BL(BL94),.BLN(BLN94),.WL(WL160));
sram_cell_6t_5 inst_cell_160_95 (.BL(BL95),.BLN(BLN95),.WL(WL160));
sram_cell_6t_5 inst_cell_160_96 (.BL(BL96),.BLN(BLN96),.WL(WL160));
sram_cell_6t_5 inst_cell_160_97 (.BL(BL97),.BLN(BLN97),.WL(WL160));
sram_cell_6t_5 inst_cell_160_98 (.BL(BL98),.BLN(BLN98),.WL(WL160));
sram_cell_6t_5 inst_cell_160_99 (.BL(BL99),.BLN(BLN99),.WL(WL160));
sram_cell_6t_5 inst_cell_160_100 (.BL(BL100),.BLN(BLN100),.WL(WL160));
sram_cell_6t_5 inst_cell_160_101 (.BL(BL101),.BLN(BLN101),.WL(WL160));
sram_cell_6t_5 inst_cell_160_102 (.BL(BL102),.BLN(BLN102),.WL(WL160));
sram_cell_6t_5 inst_cell_160_103 (.BL(BL103),.BLN(BLN103),.WL(WL160));
sram_cell_6t_5 inst_cell_160_104 (.BL(BL104),.BLN(BLN104),.WL(WL160));
sram_cell_6t_5 inst_cell_160_105 (.BL(BL105),.BLN(BLN105),.WL(WL160));
sram_cell_6t_5 inst_cell_160_106 (.BL(BL106),.BLN(BLN106),.WL(WL160));
sram_cell_6t_5 inst_cell_160_107 (.BL(BL107),.BLN(BLN107),.WL(WL160));
sram_cell_6t_5 inst_cell_160_108 (.BL(BL108),.BLN(BLN108),.WL(WL160));
sram_cell_6t_5 inst_cell_160_109 (.BL(BL109),.BLN(BLN109),.WL(WL160));
sram_cell_6t_5 inst_cell_160_110 (.BL(BL110),.BLN(BLN110),.WL(WL160));
sram_cell_6t_5 inst_cell_160_111 (.BL(BL111),.BLN(BLN111),.WL(WL160));
sram_cell_6t_5 inst_cell_160_112 (.BL(BL112),.BLN(BLN112),.WL(WL160));
sram_cell_6t_5 inst_cell_160_113 (.BL(BL113),.BLN(BLN113),.WL(WL160));
sram_cell_6t_5 inst_cell_160_114 (.BL(BL114),.BLN(BLN114),.WL(WL160));
sram_cell_6t_5 inst_cell_160_115 (.BL(BL115),.BLN(BLN115),.WL(WL160));
sram_cell_6t_5 inst_cell_160_116 (.BL(BL116),.BLN(BLN116),.WL(WL160));
sram_cell_6t_5 inst_cell_160_117 (.BL(BL117),.BLN(BLN117),.WL(WL160));
sram_cell_6t_5 inst_cell_160_118 (.BL(BL118),.BLN(BLN118),.WL(WL160));
sram_cell_6t_5 inst_cell_160_119 (.BL(BL119),.BLN(BLN119),.WL(WL160));
sram_cell_6t_5 inst_cell_160_120 (.BL(BL120),.BLN(BLN120),.WL(WL160));
sram_cell_6t_5 inst_cell_160_121 (.BL(BL121),.BLN(BLN121),.WL(WL160));
sram_cell_6t_5 inst_cell_160_122 (.BL(BL122),.BLN(BLN122),.WL(WL160));
sram_cell_6t_5 inst_cell_160_123 (.BL(BL123),.BLN(BLN123),.WL(WL160));
sram_cell_6t_5 inst_cell_160_124 (.BL(BL124),.BLN(BLN124),.WL(WL160));
sram_cell_6t_5 inst_cell_160_125 (.BL(BL125),.BLN(BLN125),.WL(WL160));
sram_cell_6t_5 inst_cell_160_126 (.BL(BL126),.BLN(BLN126),.WL(WL160));
sram_cell_6t_5 inst_cell_160_127 (.BL(BL127),.BLN(BLN127),.WL(WL160));
sram_cell_6t_5 inst_cell_161_0 (.BL(BL0),.BLN(BLN0),.WL(WL161));
sram_cell_6t_5 inst_cell_161_1 (.BL(BL1),.BLN(BLN1),.WL(WL161));
sram_cell_6t_5 inst_cell_161_2 (.BL(BL2),.BLN(BLN2),.WL(WL161));
sram_cell_6t_5 inst_cell_161_3 (.BL(BL3),.BLN(BLN3),.WL(WL161));
sram_cell_6t_5 inst_cell_161_4 (.BL(BL4),.BLN(BLN4),.WL(WL161));
sram_cell_6t_5 inst_cell_161_5 (.BL(BL5),.BLN(BLN5),.WL(WL161));
sram_cell_6t_5 inst_cell_161_6 (.BL(BL6),.BLN(BLN6),.WL(WL161));
sram_cell_6t_5 inst_cell_161_7 (.BL(BL7),.BLN(BLN7),.WL(WL161));
sram_cell_6t_5 inst_cell_161_8 (.BL(BL8),.BLN(BLN8),.WL(WL161));
sram_cell_6t_5 inst_cell_161_9 (.BL(BL9),.BLN(BLN9),.WL(WL161));
sram_cell_6t_5 inst_cell_161_10 (.BL(BL10),.BLN(BLN10),.WL(WL161));
sram_cell_6t_5 inst_cell_161_11 (.BL(BL11),.BLN(BLN11),.WL(WL161));
sram_cell_6t_5 inst_cell_161_12 (.BL(BL12),.BLN(BLN12),.WL(WL161));
sram_cell_6t_5 inst_cell_161_13 (.BL(BL13),.BLN(BLN13),.WL(WL161));
sram_cell_6t_5 inst_cell_161_14 (.BL(BL14),.BLN(BLN14),.WL(WL161));
sram_cell_6t_5 inst_cell_161_15 (.BL(BL15),.BLN(BLN15),.WL(WL161));
sram_cell_6t_5 inst_cell_161_16 (.BL(BL16),.BLN(BLN16),.WL(WL161));
sram_cell_6t_5 inst_cell_161_17 (.BL(BL17),.BLN(BLN17),.WL(WL161));
sram_cell_6t_5 inst_cell_161_18 (.BL(BL18),.BLN(BLN18),.WL(WL161));
sram_cell_6t_5 inst_cell_161_19 (.BL(BL19),.BLN(BLN19),.WL(WL161));
sram_cell_6t_5 inst_cell_161_20 (.BL(BL20),.BLN(BLN20),.WL(WL161));
sram_cell_6t_5 inst_cell_161_21 (.BL(BL21),.BLN(BLN21),.WL(WL161));
sram_cell_6t_5 inst_cell_161_22 (.BL(BL22),.BLN(BLN22),.WL(WL161));
sram_cell_6t_5 inst_cell_161_23 (.BL(BL23),.BLN(BLN23),.WL(WL161));
sram_cell_6t_5 inst_cell_161_24 (.BL(BL24),.BLN(BLN24),.WL(WL161));
sram_cell_6t_5 inst_cell_161_25 (.BL(BL25),.BLN(BLN25),.WL(WL161));
sram_cell_6t_5 inst_cell_161_26 (.BL(BL26),.BLN(BLN26),.WL(WL161));
sram_cell_6t_5 inst_cell_161_27 (.BL(BL27),.BLN(BLN27),.WL(WL161));
sram_cell_6t_5 inst_cell_161_28 (.BL(BL28),.BLN(BLN28),.WL(WL161));
sram_cell_6t_5 inst_cell_161_29 (.BL(BL29),.BLN(BLN29),.WL(WL161));
sram_cell_6t_5 inst_cell_161_30 (.BL(BL30),.BLN(BLN30),.WL(WL161));
sram_cell_6t_5 inst_cell_161_31 (.BL(BL31),.BLN(BLN31),.WL(WL161));
sram_cell_6t_5 inst_cell_161_32 (.BL(BL32),.BLN(BLN32),.WL(WL161));
sram_cell_6t_5 inst_cell_161_33 (.BL(BL33),.BLN(BLN33),.WL(WL161));
sram_cell_6t_5 inst_cell_161_34 (.BL(BL34),.BLN(BLN34),.WL(WL161));
sram_cell_6t_5 inst_cell_161_35 (.BL(BL35),.BLN(BLN35),.WL(WL161));
sram_cell_6t_5 inst_cell_161_36 (.BL(BL36),.BLN(BLN36),.WL(WL161));
sram_cell_6t_5 inst_cell_161_37 (.BL(BL37),.BLN(BLN37),.WL(WL161));
sram_cell_6t_5 inst_cell_161_38 (.BL(BL38),.BLN(BLN38),.WL(WL161));
sram_cell_6t_5 inst_cell_161_39 (.BL(BL39),.BLN(BLN39),.WL(WL161));
sram_cell_6t_5 inst_cell_161_40 (.BL(BL40),.BLN(BLN40),.WL(WL161));
sram_cell_6t_5 inst_cell_161_41 (.BL(BL41),.BLN(BLN41),.WL(WL161));
sram_cell_6t_5 inst_cell_161_42 (.BL(BL42),.BLN(BLN42),.WL(WL161));
sram_cell_6t_5 inst_cell_161_43 (.BL(BL43),.BLN(BLN43),.WL(WL161));
sram_cell_6t_5 inst_cell_161_44 (.BL(BL44),.BLN(BLN44),.WL(WL161));
sram_cell_6t_5 inst_cell_161_45 (.BL(BL45),.BLN(BLN45),.WL(WL161));
sram_cell_6t_5 inst_cell_161_46 (.BL(BL46),.BLN(BLN46),.WL(WL161));
sram_cell_6t_5 inst_cell_161_47 (.BL(BL47),.BLN(BLN47),.WL(WL161));
sram_cell_6t_5 inst_cell_161_48 (.BL(BL48),.BLN(BLN48),.WL(WL161));
sram_cell_6t_5 inst_cell_161_49 (.BL(BL49),.BLN(BLN49),.WL(WL161));
sram_cell_6t_5 inst_cell_161_50 (.BL(BL50),.BLN(BLN50),.WL(WL161));
sram_cell_6t_5 inst_cell_161_51 (.BL(BL51),.BLN(BLN51),.WL(WL161));
sram_cell_6t_5 inst_cell_161_52 (.BL(BL52),.BLN(BLN52),.WL(WL161));
sram_cell_6t_5 inst_cell_161_53 (.BL(BL53),.BLN(BLN53),.WL(WL161));
sram_cell_6t_5 inst_cell_161_54 (.BL(BL54),.BLN(BLN54),.WL(WL161));
sram_cell_6t_5 inst_cell_161_55 (.BL(BL55),.BLN(BLN55),.WL(WL161));
sram_cell_6t_5 inst_cell_161_56 (.BL(BL56),.BLN(BLN56),.WL(WL161));
sram_cell_6t_5 inst_cell_161_57 (.BL(BL57),.BLN(BLN57),.WL(WL161));
sram_cell_6t_5 inst_cell_161_58 (.BL(BL58),.BLN(BLN58),.WL(WL161));
sram_cell_6t_5 inst_cell_161_59 (.BL(BL59),.BLN(BLN59),.WL(WL161));
sram_cell_6t_5 inst_cell_161_60 (.BL(BL60),.BLN(BLN60),.WL(WL161));
sram_cell_6t_5 inst_cell_161_61 (.BL(BL61),.BLN(BLN61),.WL(WL161));
sram_cell_6t_5 inst_cell_161_62 (.BL(BL62),.BLN(BLN62),.WL(WL161));
sram_cell_6t_5 inst_cell_161_63 (.BL(BL63),.BLN(BLN63),.WL(WL161));
sram_cell_6t_5 inst_cell_161_64 (.BL(BL64),.BLN(BLN64),.WL(WL161));
sram_cell_6t_5 inst_cell_161_65 (.BL(BL65),.BLN(BLN65),.WL(WL161));
sram_cell_6t_5 inst_cell_161_66 (.BL(BL66),.BLN(BLN66),.WL(WL161));
sram_cell_6t_5 inst_cell_161_67 (.BL(BL67),.BLN(BLN67),.WL(WL161));
sram_cell_6t_5 inst_cell_161_68 (.BL(BL68),.BLN(BLN68),.WL(WL161));
sram_cell_6t_5 inst_cell_161_69 (.BL(BL69),.BLN(BLN69),.WL(WL161));
sram_cell_6t_5 inst_cell_161_70 (.BL(BL70),.BLN(BLN70),.WL(WL161));
sram_cell_6t_5 inst_cell_161_71 (.BL(BL71),.BLN(BLN71),.WL(WL161));
sram_cell_6t_5 inst_cell_161_72 (.BL(BL72),.BLN(BLN72),.WL(WL161));
sram_cell_6t_5 inst_cell_161_73 (.BL(BL73),.BLN(BLN73),.WL(WL161));
sram_cell_6t_5 inst_cell_161_74 (.BL(BL74),.BLN(BLN74),.WL(WL161));
sram_cell_6t_5 inst_cell_161_75 (.BL(BL75),.BLN(BLN75),.WL(WL161));
sram_cell_6t_5 inst_cell_161_76 (.BL(BL76),.BLN(BLN76),.WL(WL161));
sram_cell_6t_5 inst_cell_161_77 (.BL(BL77),.BLN(BLN77),.WL(WL161));
sram_cell_6t_5 inst_cell_161_78 (.BL(BL78),.BLN(BLN78),.WL(WL161));
sram_cell_6t_5 inst_cell_161_79 (.BL(BL79),.BLN(BLN79),.WL(WL161));
sram_cell_6t_5 inst_cell_161_80 (.BL(BL80),.BLN(BLN80),.WL(WL161));
sram_cell_6t_5 inst_cell_161_81 (.BL(BL81),.BLN(BLN81),.WL(WL161));
sram_cell_6t_5 inst_cell_161_82 (.BL(BL82),.BLN(BLN82),.WL(WL161));
sram_cell_6t_5 inst_cell_161_83 (.BL(BL83),.BLN(BLN83),.WL(WL161));
sram_cell_6t_5 inst_cell_161_84 (.BL(BL84),.BLN(BLN84),.WL(WL161));
sram_cell_6t_5 inst_cell_161_85 (.BL(BL85),.BLN(BLN85),.WL(WL161));
sram_cell_6t_5 inst_cell_161_86 (.BL(BL86),.BLN(BLN86),.WL(WL161));
sram_cell_6t_5 inst_cell_161_87 (.BL(BL87),.BLN(BLN87),.WL(WL161));
sram_cell_6t_5 inst_cell_161_88 (.BL(BL88),.BLN(BLN88),.WL(WL161));
sram_cell_6t_5 inst_cell_161_89 (.BL(BL89),.BLN(BLN89),.WL(WL161));
sram_cell_6t_5 inst_cell_161_90 (.BL(BL90),.BLN(BLN90),.WL(WL161));
sram_cell_6t_5 inst_cell_161_91 (.BL(BL91),.BLN(BLN91),.WL(WL161));
sram_cell_6t_5 inst_cell_161_92 (.BL(BL92),.BLN(BLN92),.WL(WL161));
sram_cell_6t_5 inst_cell_161_93 (.BL(BL93),.BLN(BLN93),.WL(WL161));
sram_cell_6t_5 inst_cell_161_94 (.BL(BL94),.BLN(BLN94),.WL(WL161));
sram_cell_6t_5 inst_cell_161_95 (.BL(BL95),.BLN(BLN95),.WL(WL161));
sram_cell_6t_5 inst_cell_161_96 (.BL(BL96),.BLN(BLN96),.WL(WL161));
sram_cell_6t_5 inst_cell_161_97 (.BL(BL97),.BLN(BLN97),.WL(WL161));
sram_cell_6t_5 inst_cell_161_98 (.BL(BL98),.BLN(BLN98),.WL(WL161));
sram_cell_6t_5 inst_cell_161_99 (.BL(BL99),.BLN(BLN99),.WL(WL161));
sram_cell_6t_5 inst_cell_161_100 (.BL(BL100),.BLN(BLN100),.WL(WL161));
sram_cell_6t_5 inst_cell_161_101 (.BL(BL101),.BLN(BLN101),.WL(WL161));
sram_cell_6t_5 inst_cell_161_102 (.BL(BL102),.BLN(BLN102),.WL(WL161));
sram_cell_6t_5 inst_cell_161_103 (.BL(BL103),.BLN(BLN103),.WL(WL161));
sram_cell_6t_5 inst_cell_161_104 (.BL(BL104),.BLN(BLN104),.WL(WL161));
sram_cell_6t_5 inst_cell_161_105 (.BL(BL105),.BLN(BLN105),.WL(WL161));
sram_cell_6t_5 inst_cell_161_106 (.BL(BL106),.BLN(BLN106),.WL(WL161));
sram_cell_6t_5 inst_cell_161_107 (.BL(BL107),.BLN(BLN107),.WL(WL161));
sram_cell_6t_5 inst_cell_161_108 (.BL(BL108),.BLN(BLN108),.WL(WL161));
sram_cell_6t_5 inst_cell_161_109 (.BL(BL109),.BLN(BLN109),.WL(WL161));
sram_cell_6t_5 inst_cell_161_110 (.BL(BL110),.BLN(BLN110),.WL(WL161));
sram_cell_6t_5 inst_cell_161_111 (.BL(BL111),.BLN(BLN111),.WL(WL161));
sram_cell_6t_5 inst_cell_161_112 (.BL(BL112),.BLN(BLN112),.WL(WL161));
sram_cell_6t_5 inst_cell_161_113 (.BL(BL113),.BLN(BLN113),.WL(WL161));
sram_cell_6t_5 inst_cell_161_114 (.BL(BL114),.BLN(BLN114),.WL(WL161));
sram_cell_6t_5 inst_cell_161_115 (.BL(BL115),.BLN(BLN115),.WL(WL161));
sram_cell_6t_5 inst_cell_161_116 (.BL(BL116),.BLN(BLN116),.WL(WL161));
sram_cell_6t_5 inst_cell_161_117 (.BL(BL117),.BLN(BLN117),.WL(WL161));
sram_cell_6t_5 inst_cell_161_118 (.BL(BL118),.BLN(BLN118),.WL(WL161));
sram_cell_6t_5 inst_cell_161_119 (.BL(BL119),.BLN(BLN119),.WL(WL161));
sram_cell_6t_5 inst_cell_161_120 (.BL(BL120),.BLN(BLN120),.WL(WL161));
sram_cell_6t_5 inst_cell_161_121 (.BL(BL121),.BLN(BLN121),.WL(WL161));
sram_cell_6t_5 inst_cell_161_122 (.BL(BL122),.BLN(BLN122),.WL(WL161));
sram_cell_6t_5 inst_cell_161_123 (.BL(BL123),.BLN(BLN123),.WL(WL161));
sram_cell_6t_5 inst_cell_161_124 (.BL(BL124),.BLN(BLN124),.WL(WL161));
sram_cell_6t_5 inst_cell_161_125 (.BL(BL125),.BLN(BLN125),.WL(WL161));
sram_cell_6t_5 inst_cell_161_126 (.BL(BL126),.BLN(BLN126),.WL(WL161));
sram_cell_6t_5 inst_cell_161_127 (.BL(BL127),.BLN(BLN127),.WL(WL161));
sram_cell_6t_5 inst_cell_162_0 (.BL(BL0),.BLN(BLN0),.WL(WL162));
sram_cell_6t_5 inst_cell_162_1 (.BL(BL1),.BLN(BLN1),.WL(WL162));
sram_cell_6t_5 inst_cell_162_2 (.BL(BL2),.BLN(BLN2),.WL(WL162));
sram_cell_6t_5 inst_cell_162_3 (.BL(BL3),.BLN(BLN3),.WL(WL162));
sram_cell_6t_5 inst_cell_162_4 (.BL(BL4),.BLN(BLN4),.WL(WL162));
sram_cell_6t_5 inst_cell_162_5 (.BL(BL5),.BLN(BLN5),.WL(WL162));
sram_cell_6t_5 inst_cell_162_6 (.BL(BL6),.BLN(BLN6),.WL(WL162));
sram_cell_6t_5 inst_cell_162_7 (.BL(BL7),.BLN(BLN7),.WL(WL162));
sram_cell_6t_5 inst_cell_162_8 (.BL(BL8),.BLN(BLN8),.WL(WL162));
sram_cell_6t_5 inst_cell_162_9 (.BL(BL9),.BLN(BLN9),.WL(WL162));
sram_cell_6t_5 inst_cell_162_10 (.BL(BL10),.BLN(BLN10),.WL(WL162));
sram_cell_6t_5 inst_cell_162_11 (.BL(BL11),.BLN(BLN11),.WL(WL162));
sram_cell_6t_5 inst_cell_162_12 (.BL(BL12),.BLN(BLN12),.WL(WL162));
sram_cell_6t_5 inst_cell_162_13 (.BL(BL13),.BLN(BLN13),.WL(WL162));
sram_cell_6t_5 inst_cell_162_14 (.BL(BL14),.BLN(BLN14),.WL(WL162));
sram_cell_6t_5 inst_cell_162_15 (.BL(BL15),.BLN(BLN15),.WL(WL162));
sram_cell_6t_5 inst_cell_162_16 (.BL(BL16),.BLN(BLN16),.WL(WL162));
sram_cell_6t_5 inst_cell_162_17 (.BL(BL17),.BLN(BLN17),.WL(WL162));
sram_cell_6t_5 inst_cell_162_18 (.BL(BL18),.BLN(BLN18),.WL(WL162));
sram_cell_6t_5 inst_cell_162_19 (.BL(BL19),.BLN(BLN19),.WL(WL162));
sram_cell_6t_5 inst_cell_162_20 (.BL(BL20),.BLN(BLN20),.WL(WL162));
sram_cell_6t_5 inst_cell_162_21 (.BL(BL21),.BLN(BLN21),.WL(WL162));
sram_cell_6t_5 inst_cell_162_22 (.BL(BL22),.BLN(BLN22),.WL(WL162));
sram_cell_6t_5 inst_cell_162_23 (.BL(BL23),.BLN(BLN23),.WL(WL162));
sram_cell_6t_5 inst_cell_162_24 (.BL(BL24),.BLN(BLN24),.WL(WL162));
sram_cell_6t_5 inst_cell_162_25 (.BL(BL25),.BLN(BLN25),.WL(WL162));
sram_cell_6t_5 inst_cell_162_26 (.BL(BL26),.BLN(BLN26),.WL(WL162));
sram_cell_6t_5 inst_cell_162_27 (.BL(BL27),.BLN(BLN27),.WL(WL162));
sram_cell_6t_5 inst_cell_162_28 (.BL(BL28),.BLN(BLN28),.WL(WL162));
sram_cell_6t_5 inst_cell_162_29 (.BL(BL29),.BLN(BLN29),.WL(WL162));
sram_cell_6t_5 inst_cell_162_30 (.BL(BL30),.BLN(BLN30),.WL(WL162));
sram_cell_6t_5 inst_cell_162_31 (.BL(BL31),.BLN(BLN31),.WL(WL162));
sram_cell_6t_5 inst_cell_162_32 (.BL(BL32),.BLN(BLN32),.WL(WL162));
sram_cell_6t_5 inst_cell_162_33 (.BL(BL33),.BLN(BLN33),.WL(WL162));
sram_cell_6t_5 inst_cell_162_34 (.BL(BL34),.BLN(BLN34),.WL(WL162));
sram_cell_6t_5 inst_cell_162_35 (.BL(BL35),.BLN(BLN35),.WL(WL162));
sram_cell_6t_5 inst_cell_162_36 (.BL(BL36),.BLN(BLN36),.WL(WL162));
sram_cell_6t_5 inst_cell_162_37 (.BL(BL37),.BLN(BLN37),.WL(WL162));
sram_cell_6t_5 inst_cell_162_38 (.BL(BL38),.BLN(BLN38),.WL(WL162));
sram_cell_6t_5 inst_cell_162_39 (.BL(BL39),.BLN(BLN39),.WL(WL162));
sram_cell_6t_5 inst_cell_162_40 (.BL(BL40),.BLN(BLN40),.WL(WL162));
sram_cell_6t_5 inst_cell_162_41 (.BL(BL41),.BLN(BLN41),.WL(WL162));
sram_cell_6t_5 inst_cell_162_42 (.BL(BL42),.BLN(BLN42),.WL(WL162));
sram_cell_6t_5 inst_cell_162_43 (.BL(BL43),.BLN(BLN43),.WL(WL162));
sram_cell_6t_5 inst_cell_162_44 (.BL(BL44),.BLN(BLN44),.WL(WL162));
sram_cell_6t_5 inst_cell_162_45 (.BL(BL45),.BLN(BLN45),.WL(WL162));
sram_cell_6t_5 inst_cell_162_46 (.BL(BL46),.BLN(BLN46),.WL(WL162));
sram_cell_6t_5 inst_cell_162_47 (.BL(BL47),.BLN(BLN47),.WL(WL162));
sram_cell_6t_5 inst_cell_162_48 (.BL(BL48),.BLN(BLN48),.WL(WL162));
sram_cell_6t_5 inst_cell_162_49 (.BL(BL49),.BLN(BLN49),.WL(WL162));
sram_cell_6t_5 inst_cell_162_50 (.BL(BL50),.BLN(BLN50),.WL(WL162));
sram_cell_6t_5 inst_cell_162_51 (.BL(BL51),.BLN(BLN51),.WL(WL162));
sram_cell_6t_5 inst_cell_162_52 (.BL(BL52),.BLN(BLN52),.WL(WL162));
sram_cell_6t_5 inst_cell_162_53 (.BL(BL53),.BLN(BLN53),.WL(WL162));
sram_cell_6t_5 inst_cell_162_54 (.BL(BL54),.BLN(BLN54),.WL(WL162));
sram_cell_6t_5 inst_cell_162_55 (.BL(BL55),.BLN(BLN55),.WL(WL162));
sram_cell_6t_5 inst_cell_162_56 (.BL(BL56),.BLN(BLN56),.WL(WL162));
sram_cell_6t_5 inst_cell_162_57 (.BL(BL57),.BLN(BLN57),.WL(WL162));
sram_cell_6t_5 inst_cell_162_58 (.BL(BL58),.BLN(BLN58),.WL(WL162));
sram_cell_6t_5 inst_cell_162_59 (.BL(BL59),.BLN(BLN59),.WL(WL162));
sram_cell_6t_5 inst_cell_162_60 (.BL(BL60),.BLN(BLN60),.WL(WL162));
sram_cell_6t_5 inst_cell_162_61 (.BL(BL61),.BLN(BLN61),.WL(WL162));
sram_cell_6t_5 inst_cell_162_62 (.BL(BL62),.BLN(BLN62),.WL(WL162));
sram_cell_6t_5 inst_cell_162_63 (.BL(BL63),.BLN(BLN63),.WL(WL162));
sram_cell_6t_5 inst_cell_162_64 (.BL(BL64),.BLN(BLN64),.WL(WL162));
sram_cell_6t_5 inst_cell_162_65 (.BL(BL65),.BLN(BLN65),.WL(WL162));
sram_cell_6t_5 inst_cell_162_66 (.BL(BL66),.BLN(BLN66),.WL(WL162));
sram_cell_6t_5 inst_cell_162_67 (.BL(BL67),.BLN(BLN67),.WL(WL162));
sram_cell_6t_5 inst_cell_162_68 (.BL(BL68),.BLN(BLN68),.WL(WL162));
sram_cell_6t_5 inst_cell_162_69 (.BL(BL69),.BLN(BLN69),.WL(WL162));
sram_cell_6t_5 inst_cell_162_70 (.BL(BL70),.BLN(BLN70),.WL(WL162));
sram_cell_6t_5 inst_cell_162_71 (.BL(BL71),.BLN(BLN71),.WL(WL162));
sram_cell_6t_5 inst_cell_162_72 (.BL(BL72),.BLN(BLN72),.WL(WL162));
sram_cell_6t_5 inst_cell_162_73 (.BL(BL73),.BLN(BLN73),.WL(WL162));
sram_cell_6t_5 inst_cell_162_74 (.BL(BL74),.BLN(BLN74),.WL(WL162));
sram_cell_6t_5 inst_cell_162_75 (.BL(BL75),.BLN(BLN75),.WL(WL162));
sram_cell_6t_5 inst_cell_162_76 (.BL(BL76),.BLN(BLN76),.WL(WL162));
sram_cell_6t_5 inst_cell_162_77 (.BL(BL77),.BLN(BLN77),.WL(WL162));
sram_cell_6t_5 inst_cell_162_78 (.BL(BL78),.BLN(BLN78),.WL(WL162));
sram_cell_6t_5 inst_cell_162_79 (.BL(BL79),.BLN(BLN79),.WL(WL162));
sram_cell_6t_5 inst_cell_162_80 (.BL(BL80),.BLN(BLN80),.WL(WL162));
sram_cell_6t_5 inst_cell_162_81 (.BL(BL81),.BLN(BLN81),.WL(WL162));
sram_cell_6t_5 inst_cell_162_82 (.BL(BL82),.BLN(BLN82),.WL(WL162));
sram_cell_6t_5 inst_cell_162_83 (.BL(BL83),.BLN(BLN83),.WL(WL162));
sram_cell_6t_5 inst_cell_162_84 (.BL(BL84),.BLN(BLN84),.WL(WL162));
sram_cell_6t_5 inst_cell_162_85 (.BL(BL85),.BLN(BLN85),.WL(WL162));
sram_cell_6t_5 inst_cell_162_86 (.BL(BL86),.BLN(BLN86),.WL(WL162));
sram_cell_6t_5 inst_cell_162_87 (.BL(BL87),.BLN(BLN87),.WL(WL162));
sram_cell_6t_5 inst_cell_162_88 (.BL(BL88),.BLN(BLN88),.WL(WL162));
sram_cell_6t_5 inst_cell_162_89 (.BL(BL89),.BLN(BLN89),.WL(WL162));
sram_cell_6t_5 inst_cell_162_90 (.BL(BL90),.BLN(BLN90),.WL(WL162));
sram_cell_6t_5 inst_cell_162_91 (.BL(BL91),.BLN(BLN91),.WL(WL162));
sram_cell_6t_5 inst_cell_162_92 (.BL(BL92),.BLN(BLN92),.WL(WL162));
sram_cell_6t_5 inst_cell_162_93 (.BL(BL93),.BLN(BLN93),.WL(WL162));
sram_cell_6t_5 inst_cell_162_94 (.BL(BL94),.BLN(BLN94),.WL(WL162));
sram_cell_6t_5 inst_cell_162_95 (.BL(BL95),.BLN(BLN95),.WL(WL162));
sram_cell_6t_5 inst_cell_162_96 (.BL(BL96),.BLN(BLN96),.WL(WL162));
sram_cell_6t_5 inst_cell_162_97 (.BL(BL97),.BLN(BLN97),.WL(WL162));
sram_cell_6t_5 inst_cell_162_98 (.BL(BL98),.BLN(BLN98),.WL(WL162));
sram_cell_6t_5 inst_cell_162_99 (.BL(BL99),.BLN(BLN99),.WL(WL162));
sram_cell_6t_5 inst_cell_162_100 (.BL(BL100),.BLN(BLN100),.WL(WL162));
sram_cell_6t_5 inst_cell_162_101 (.BL(BL101),.BLN(BLN101),.WL(WL162));
sram_cell_6t_5 inst_cell_162_102 (.BL(BL102),.BLN(BLN102),.WL(WL162));
sram_cell_6t_5 inst_cell_162_103 (.BL(BL103),.BLN(BLN103),.WL(WL162));
sram_cell_6t_5 inst_cell_162_104 (.BL(BL104),.BLN(BLN104),.WL(WL162));
sram_cell_6t_5 inst_cell_162_105 (.BL(BL105),.BLN(BLN105),.WL(WL162));
sram_cell_6t_5 inst_cell_162_106 (.BL(BL106),.BLN(BLN106),.WL(WL162));
sram_cell_6t_5 inst_cell_162_107 (.BL(BL107),.BLN(BLN107),.WL(WL162));
sram_cell_6t_5 inst_cell_162_108 (.BL(BL108),.BLN(BLN108),.WL(WL162));
sram_cell_6t_5 inst_cell_162_109 (.BL(BL109),.BLN(BLN109),.WL(WL162));
sram_cell_6t_5 inst_cell_162_110 (.BL(BL110),.BLN(BLN110),.WL(WL162));
sram_cell_6t_5 inst_cell_162_111 (.BL(BL111),.BLN(BLN111),.WL(WL162));
sram_cell_6t_5 inst_cell_162_112 (.BL(BL112),.BLN(BLN112),.WL(WL162));
sram_cell_6t_5 inst_cell_162_113 (.BL(BL113),.BLN(BLN113),.WL(WL162));
sram_cell_6t_5 inst_cell_162_114 (.BL(BL114),.BLN(BLN114),.WL(WL162));
sram_cell_6t_5 inst_cell_162_115 (.BL(BL115),.BLN(BLN115),.WL(WL162));
sram_cell_6t_5 inst_cell_162_116 (.BL(BL116),.BLN(BLN116),.WL(WL162));
sram_cell_6t_5 inst_cell_162_117 (.BL(BL117),.BLN(BLN117),.WL(WL162));
sram_cell_6t_5 inst_cell_162_118 (.BL(BL118),.BLN(BLN118),.WL(WL162));
sram_cell_6t_5 inst_cell_162_119 (.BL(BL119),.BLN(BLN119),.WL(WL162));
sram_cell_6t_5 inst_cell_162_120 (.BL(BL120),.BLN(BLN120),.WL(WL162));
sram_cell_6t_5 inst_cell_162_121 (.BL(BL121),.BLN(BLN121),.WL(WL162));
sram_cell_6t_5 inst_cell_162_122 (.BL(BL122),.BLN(BLN122),.WL(WL162));
sram_cell_6t_5 inst_cell_162_123 (.BL(BL123),.BLN(BLN123),.WL(WL162));
sram_cell_6t_5 inst_cell_162_124 (.BL(BL124),.BLN(BLN124),.WL(WL162));
sram_cell_6t_5 inst_cell_162_125 (.BL(BL125),.BLN(BLN125),.WL(WL162));
sram_cell_6t_5 inst_cell_162_126 (.BL(BL126),.BLN(BLN126),.WL(WL162));
sram_cell_6t_5 inst_cell_162_127 (.BL(BL127),.BLN(BLN127),.WL(WL162));
sram_cell_6t_5 inst_cell_163_0 (.BL(BL0),.BLN(BLN0),.WL(WL163));
sram_cell_6t_5 inst_cell_163_1 (.BL(BL1),.BLN(BLN1),.WL(WL163));
sram_cell_6t_5 inst_cell_163_2 (.BL(BL2),.BLN(BLN2),.WL(WL163));
sram_cell_6t_5 inst_cell_163_3 (.BL(BL3),.BLN(BLN3),.WL(WL163));
sram_cell_6t_5 inst_cell_163_4 (.BL(BL4),.BLN(BLN4),.WL(WL163));
sram_cell_6t_5 inst_cell_163_5 (.BL(BL5),.BLN(BLN5),.WL(WL163));
sram_cell_6t_5 inst_cell_163_6 (.BL(BL6),.BLN(BLN6),.WL(WL163));
sram_cell_6t_5 inst_cell_163_7 (.BL(BL7),.BLN(BLN7),.WL(WL163));
sram_cell_6t_5 inst_cell_163_8 (.BL(BL8),.BLN(BLN8),.WL(WL163));
sram_cell_6t_5 inst_cell_163_9 (.BL(BL9),.BLN(BLN9),.WL(WL163));
sram_cell_6t_5 inst_cell_163_10 (.BL(BL10),.BLN(BLN10),.WL(WL163));
sram_cell_6t_5 inst_cell_163_11 (.BL(BL11),.BLN(BLN11),.WL(WL163));
sram_cell_6t_5 inst_cell_163_12 (.BL(BL12),.BLN(BLN12),.WL(WL163));
sram_cell_6t_5 inst_cell_163_13 (.BL(BL13),.BLN(BLN13),.WL(WL163));
sram_cell_6t_5 inst_cell_163_14 (.BL(BL14),.BLN(BLN14),.WL(WL163));
sram_cell_6t_5 inst_cell_163_15 (.BL(BL15),.BLN(BLN15),.WL(WL163));
sram_cell_6t_5 inst_cell_163_16 (.BL(BL16),.BLN(BLN16),.WL(WL163));
sram_cell_6t_5 inst_cell_163_17 (.BL(BL17),.BLN(BLN17),.WL(WL163));
sram_cell_6t_5 inst_cell_163_18 (.BL(BL18),.BLN(BLN18),.WL(WL163));
sram_cell_6t_5 inst_cell_163_19 (.BL(BL19),.BLN(BLN19),.WL(WL163));
sram_cell_6t_5 inst_cell_163_20 (.BL(BL20),.BLN(BLN20),.WL(WL163));
sram_cell_6t_5 inst_cell_163_21 (.BL(BL21),.BLN(BLN21),.WL(WL163));
sram_cell_6t_5 inst_cell_163_22 (.BL(BL22),.BLN(BLN22),.WL(WL163));
sram_cell_6t_5 inst_cell_163_23 (.BL(BL23),.BLN(BLN23),.WL(WL163));
sram_cell_6t_5 inst_cell_163_24 (.BL(BL24),.BLN(BLN24),.WL(WL163));
sram_cell_6t_5 inst_cell_163_25 (.BL(BL25),.BLN(BLN25),.WL(WL163));
sram_cell_6t_5 inst_cell_163_26 (.BL(BL26),.BLN(BLN26),.WL(WL163));
sram_cell_6t_5 inst_cell_163_27 (.BL(BL27),.BLN(BLN27),.WL(WL163));
sram_cell_6t_5 inst_cell_163_28 (.BL(BL28),.BLN(BLN28),.WL(WL163));
sram_cell_6t_5 inst_cell_163_29 (.BL(BL29),.BLN(BLN29),.WL(WL163));
sram_cell_6t_5 inst_cell_163_30 (.BL(BL30),.BLN(BLN30),.WL(WL163));
sram_cell_6t_5 inst_cell_163_31 (.BL(BL31),.BLN(BLN31),.WL(WL163));
sram_cell_6t_5 inst_cell_163_32 (.BL(BL32),.BLN(BLN32),.WL(WL163));
sram_cell_6t_5 inst_cell_163_33 (.BL(BL33),.BLN(BLN33),.WL(WL163));
sram_cell_6t_5 inst_cell_163_34 (.BL(BL34),.BLN(BLN34),.WL(WL163));
sram_cell_6t_5 inst_cell_163_35 (.BL(BL35),.BLN(BLN35),.WL(WL163));
sram_cell_6t_5 inst_cell_163_36 (.BL(BL36),.BLN(BLN36),.WL(WL163));
sram_cell_6t_5 inst_cell_163_37 (.BL(BL37),.BLN(BLN37),.WL(WL163));
sram_cell_6t_5 inst_cell_163_38 (.BL(BL38),.BLN(BLN38),.WL(WL163));
sram_cell_6t_5 inst_cell_163_39 (.BL(BL39),.BLN(BLN39),.WL(WL163));
sram_cell_6t_5 inst_cell_163_40 (.BL(BL40),.BLN(BLN40),.WL(WL163));
sram_cell_6t_5 inst_cell_163_41 (.BL(BL41),.BLN(BLN41),.WL(WL163));
sram_cell_6t_5 inst_cell_163_42 (.BL(BL42),.BLN(BLN42),.WL(WL163));
sram_cell_6t_5 inst_cell_163_43 (.BL(BL43),.BLN(BLN43),.WL(WL163));
sram_cell_6t_5 inst_cell_163_44 (.BL(BL44),.BLN(BLN44),.WL(WL163));
sram_cell_6t_5 inst_cell_163_45 (.BL(BL45),.BLN(BLN45),.WL(WL163));
sram_cell_6t_5 inst_cell_163_46 (.BL(BL46),.BLN(BLN46),.WL(WL163));
sram_cell_6t_5 inst_cell_163_47 (.BL(BL47),.BLN(BLN47),.WL(WL163));
sram_cell_6t_5 inst_cell_163_48 (.BL(BL48),.BLN(BLN48),.WL(WL163));
sram_cell_6t_5 inst_cell_163_49 (.BL(BL49),.BLN(BLN49),.WL(WL163));
sram_cell_6t_5 inst_cell_163_50 (.BL(BL50),.BLN(BLN50),.WL(WL163));
sram_cell_6t_5 inst_cell_163_51 (.BL(BL51),.BLN(BLN51),.WL(WL163));
sram_cell_6t_5 inst_cell_163_52 (.BL(BL52),.BLN(BLN52),.WL(WL163));
sram_cell_6t_5 inst_cell_163_53 (.BL(BL53),.BLN(BLN53),.WL(WL163));
sram_cell_6t_5 inst_cell_163_54 (.BL(BL54),.BLN(BLN54),.WL(WL163));
sram_cell_6t_5 inst_cell_163_55 (.BL(BL55),.BLN(BLN55),.WL(WL163));
sram_cell_6t_5 inst_cell_163_56 (.BL(BL56),.BLN(BLN56),.WL(WL163));
sram_cell_6t_5 inst_cell_163_57 (.BL(BL57),.BLN(BLN57),.WL(WL163));
sram_cell_6t_5 inst_cell_163_58 (.BL(BL58),.BLN(BLN58),.WL(WL163));
sram_cell_6t_5 inst_cell_163_59 (.BL(BL59),.BLN(BLN59),.WL(WL163));
sram_cell_6t_5 inst_cell_163_60 (.BL(BL60),.BLN(BLN60),.WL(WL163));
sram_cell_6t_5 inst_cell_163_61 (.BL(BL61),.BLN(BLN61),.WL(WL163));
sram_cell_6t_5 inst_cell_163_62 (.BL(BL62),.BLN(BLN62),.WL(WL163));
sram_cell_6t_5 inst_cell_163_63 (.BL(BL63),.BLN(BLN63),.WL(WL163));
sram_cell_6t_5 inst_cell_163_64 (.BL(BL64),.BLN(BLN64),.WL(WL163));
sram_cell_6t_5 inst_cell_163_65 (.BL(BL65),.BLN(BLN65),.WL(WL163));
sram_cell_6t_5 inst_cell_163_66 (.BL(BL66),.BLN(BLN66),.WL(WL163));
sram_cell_6t_5 inst_cell_163_67 (.BL(BL67),.BLN(BLN67),.WL(WL163));
sram_cell_6t_5 inst_cell_163_68 (.BL(BL68),.BLN(BLN68),.WL(WL163));
sram_cell_6t_5 inst_cell_163_69 (.BL(BL69),.BLN(BLN69),.WL(WL163));
sram_cell_6t_5 inst_cell_163_70 (.BL(BL70),.BLN(BLN70),.WL(WL163));
sram_cell_6t_5 inst_cell_163_71 (.BL(BL71),.BLN(BLN71),.WL(WL163));
sram_cell_6t_5 inst_cell_163_72 (.BL(BL72),.BLN(BLN72),.WL(WL163));
sram_cell_6t_5 inst_cell_163_73 (.BL(BL73),.BLN(BLN73),.WL(WL163));
sram_cell_6t_5 inst_cell_163_74 (.BL(BL74),.BLN(BLN74),.WL(WL163));
sram_cell_6t_5 inst_cell_163_75 (.BL(BL75),.BLN(BLN75),.WL(WL163));
sram_cell_6t_5 inst_cell_163_76 (.BL(BL76),.BLN(BLN76),.WL(WL163));
sram_cell_6t_5 inst_cell_163_77 (.BL(BL77),.BLN(BLN77),.WL(WL163));
sram_cell_6t_5 inst_cell_163_78 (.BL(BL78),.BLN(BLN78),.WL(WL163));
sram_cell_6t_5 inst_cell_163_79 (.BL(BL79),.BLN(BLN79),.WL(WL163));
sram_cell_6t_5 inst_cell_163_80 (.BL(BL80),.BLN(BLN80),.WL(WL163));
sram_cell_6t_5 inst_cell_163_81 (.BL(BL81),.BLN(BLN81),.WL(WL163));
sram_cell_6t_5 inst_cell_163_82 (.BL(BL82),.BLN(BLN82),.WL(WL163));
sram_cell_6t_5 inst_cell_163_83 (.BL(BL83),.BLN(BLN83),.WL(WL163));
sram_cell_6t_5 inst_cell_163_84 (.BL(BL84),.BLN(BLN84),.WL(WL163));
sram_cell_6t_5 inst_cell_163_85 (.BL(BL85),.BLN(BLN85),.WL(WL163));
sram_cell_6t_5 inst_cell_163_86 (.BL(BL86),.BLN(BLN86),.WL(WL163));
sram_cell_6t_5 inst_cell_163_87 (.BL(BL87),.BLN(BLN87),.WL(WL163));
sram_cell_6t_5 inst_cell_163_88 (.BL(BL88),.BLN(BLN88),.WL(WL163));
sram_cell_6t_5 inst_cell_163_89 (.BL(BL89),.BLN(BLN89),.WL(WL163));
sram_cell_6t_5 inst_cell_163_90 (.BL(BL90),.BLN(BLN90),.WL(WL163));
sram_cell_6t_5 inst_cell_163_91 (.BL(BL91),.BLN(BLN91),.WL(WL163));
sram_cell_6t_5 inst_cell_163_92 (.BL(BL92),.BLN(BLN92),.WL(WL163));
sram_cell_6t_5 inst_cell_163_93 (.BL(BL93),.BLN(BLN93),.WL(WL163));
sram_cell_6t_5 inst_cell_163_94 (.BL(BL94),.BLN(BLN94),.WL(WL163));
sram_cell_6t_5 inst_cell_163_95 (.BL(BL95),.BLN(BLN95),.WL(WL163));
sram_cell_6t_5 inst_cell_163_96 (.BL(BL96),.BLN(BLN96),.WL(WL163));
sram_cell_6t_5 inst_cell_163_97 (.BL(BL97),.BLN(BLN97),.WL(WL163));
sram_cell_6t_5 inst_cell_163_98 (.BL(BL98),.BLN(BLN98),.WL(WL163));
sram_cell_6t_5 inst_cell_163_99 (.BL(BL99),.BLN(BLN99),.WL(WL163));
sram_cell_6t_5 inst_cell_163_100 (.BL(BL100),.BLN(BLN100),.WL(WL163));
sram_cell_6t_5 inst_cell_163_101 (.BL(BL101),.BLN(BLN101),.WL(WL163));
sram_cell_6t_5 inst_cell_163_102 (.BL(BL102),.BLN(BLN102),.WL(WL163));
sram_cell_6t_5 inst_cell_163_103 (.BL(BL103),.BLN(BLN103),.WL(WL163));
sram_cell_6t_5 inst_cell_163_104 (.BL(BL104),.BLN(BLN104),.WL(WL163));
sram_cell_6t_5 inst_cell_163_105 (.BL(BL105),.BLN(BLN105),.WL(WL163));
sram_cell_6t_5 inst_cell_163_106 (.BL(BL106),.BLN(BLN106),.WL(WL163));
sram_cell_6t_5 inst_cell_163_107 (.BL(BL107),.BLN(BLN107),.WL(WL163));
sram_cell_6t_5 inst_cell_163_108 (.BL(BL108),.BLN(BLN108),.WL(WL163));
sram_cell_6t_5 inst_cell_163_109 (.BL(BL109),.BLN(BLN109),.WL(WL163));
sram_cell_6t_5 inst_cell_163_110 (.BL(BL110),.BLN(BLN110),.WL(WL163));
sram_cell_6t_5 inst_cell_163_111 (.BL(BL111),.BLN(BLN111),.WL(WL163));
sram_cell_6t_5 inst_cell_163_112 (.BL(BL112),.BLN(BLN112),.WL(WL163));
sram_cell_6t_5 inst_cell_163_113 (.BL(BL113),.BLN(BLN113),.WL(WL163));
sram_cell_6t_5 inst_cell_163_114 (.BL(BL114),.BLN(BLN114),.WL(WL163));
sram_cell_6t_5 inst_cell_163_115 (.BL(BL115),.BLN(BLN115),.WL(WL163));
sram_cell_6t_5 inst_cell_163_116 (.BL(BL116),.BLN(BLN116),.WL(WL163));
sram_cell_6t_5 inst_cell_163_117 (.BL(BL117),.BLN(BLN117),.WL(WL163));
sram_cell_6t_5 inst_cell_163_118 (.BL(BL118),.BLN(BLN118),.WL(WL163));
sram_cell_6t_5 inst_cell_163_119 (.BL(BL119),.BLN(BLN119),.WL(WL163));
sram_cell_6t_5 inst_cell_163_120 (.BL(BL120),.BLN(BLN120),.WL(WL163));
sram_cell_6t_5 inst_cell_163_121 (.BL(BL121),.BLN(BLN121),.WL(WL163));
sram_cell_6t_5 inst_cell_163_122 (.BL(BL122),.BLN(BLN122),.WL(WL163));
sram_cell_6t_5 inst_cell_163_123 (.BL(BL123),.BLN(BLN123),.WL(WL163));
sram_cell_6t_5 inst_cell_163_124 (.BL(BL124),.BLN(BLN124),.WL(WL163));
sram_cell_6t_5 inst_cell_163_125 (.BL(BL125),.BLN(BLN125),.WL(WL163));
sram_cell_6t_5 inst_cell_163_126 (.BL(BL126),.BLN(BLN126),.WL(WL163));
sram_cell_6t_5 inst_cell_163_127 (.BL(BL127),.BLN(BLN127),.WL(WL163));
sram_cell_6t_5 inst_cell_164_0 (.BL(BL0),.BLN(BLN0),.WL(WL164));
sram_cell_6t_5 inst_cell_164_1 (.BL(BL1),.BLN(BLN1),.WL(WL164));
sram_cell_6t_5 inst_cell_164_2 (.BL(BL2),.BLN(BLN2),.WL(WL164));
sram_cell_6t_5 inst_cell_164_3 (.BL(BL3),.BLN(BLN3),.WL(WL164));
sram_cell_6t_5 inst_cell_164_4 (.BL(BL4),.BLN(BLN4),.WL(WL164));
sram_cell_6t_5 inst_cell_164_5 (.BL(BL5),.BLN(BLN5),.WL(WL164));
sram_cell_6t_5 inst_cell_164_6 (.BL(BL6),.BLN(BLN6),.WL(WL164));
sram_cell_6t_5 inst_cell_164_7 (.BL(BL7),.BLN(BLN7),.WL(WL164));
sram_cell_6t_5 inst_cell_164_8 (.BL(BL8),.BLN(BLN8),.WL(WL164));
sram_cell_6t_5 inst_cell_164_9 (.BL(BL9),.BLN(BLN9),.WL(WL164));
sram_cell_6t_5 inst_cell_164_10 (.BL(BL10),.BLN(BLN10),.WL(WL164));
sram_cell_6t_5 inst_cell_164_11 (.BL(BL11),.BLN(BLN11),.WL(WL164));
sram_cell_6t_5 inst_cell_164_12 (.BL(BL12),.BLN(BLN12),.WL(WL164));
sram_cell_6t_5 inst_cell_164_13 (.BL(BL13),.BLN(BLN13),.WL(WL164));
sram_cell_6t_5 inst_cell_164_14 (.BL(BL14),.BLN(BLN14),.WL(WL164));
sram_cell_6t_5 inst_cell_164_15 (.BL(BL15),.BLN(BLN15),.WL(WL164));
sram_cell_6t_5 inst_cell_164_16 (.BL(BL16),.BLN(BLN16),.WL(WL164));
sram_cell_6t_5 inst_cell_164_17 (.BL(BL17),.BLN(BLN17),.WL(WL164));
sram_cell_6t_5 inst_cell_164_18 (.BL(BL18),.BLN(BLN18),.WL(WL164));
sram_cell_6t_5 inst_cell_164_19 (.BL(BL19),.BLN(BLN19),.WL(WL164));
sram_cell_6t_5 inst_cell_164_20 (.BL(BL20),.BLN(BLN20),.WL(WL164));
sram_cell_6t_5 inst_cell_164_21 (.BL(BL21),.BLN(BLN21),.WL(WL164));
sram_cell_6t_5 inst_cell_164_22 (.BL(BL22),.BLN(BLN22),.WL(WL164));
sram_cell_6t_5 inst_cell_164_23 (.BL(BL23),.BLN(BLN23),.WL(WL164));
sram_cell_6t_5 inst_cell_164_24 (.BL(BL24),.BLN(BLN24),.WL(WL164));
sram_cell_6t_5 inst_cell_164_25 (.BL(BL25),.BLN(BLN25),.WL(WL164));
sram_cell_6t_5 inst_cell_164_26 (.BL(BL26),.BLN(BLN26),.WL(WL164));
sram_cell_6t_5 inst_cell_164_27 (.BL(BL27),.BLN(BLN27),.WL(WL164));
sram_cell_6t_5 inst_cell_164_28 (.BL(BL28),.BLN(BLN28),.WL(WL164));
sram_cell_6t_5 inst_cell_164_29 (.BL(BL29),.BLN(BLN29),.WL(WL164));
sram_cell_6t_5 inst_cell_164_30 (.BL(BL30),.BLN(BLN30),.WL(WL164));
sram_cell_6t_5 inst_cell_164_31 (.BL(BL31),.BLN(BLN31),.WL(WL164));
sram_cell_6t_5 inst_cell_164_32 (.BL(BL32),.BLN(BLN32),.WL(WL164));
sram_cell_6t_5 inst_cell_164_33 (.BL(BL33),.BLN(BLN33),.WL(WL164));
sram_cell_6t_5 inst_cell_164_34 (.BL(BL34),.BLN(BLN34),.WL(WL164));
sram_cell_6t_5 inst_cell_164_35 (.BL(BL35),.BLN(BLN35),.WL(WL164));
sram_cell_6t_5 inst_cell_164_36 (.BL(BL36),.BLN(BLN36),.WL(WL164));
sram_cell_6t_5 inst_cell_164_37 (.BL(BL37),.BLN(BLN37),.WL(WL164));
sram_cell_6t_5 inst_cell_164_38 (.BL(BL38),.BLN(BLN38),.WL(WL164));
sram_cell_6t_5 inst_cell_164_39 (.BL(BL39),.BLN(BLN39),.WL(WL164));
sram_cell_6t_5 inst_cell_164_40 (.BL(BL40),.BLN(BLN40),.WL(WL164));
sram_cell_6t_5 inst_cell_164_41 (.BL(BL41),.BLN(BLN41),.WL(WL164));
sram_cell_6t_5 inst_cell_164_42 (.BL(BL42),.BLN(BLN42),.WL(WL164));
sram_cell_6t_5 inst_cell_164_43 (.BL(BL43),.BLN(BLN43),.WL(WL164));
sram_cell_6t_5 inst_cell_164_44 (.BL(BL44),.BLN(BLN44),.WL(WL164));
sram_cell_6t_5 inst_cell_164_45 (.BL(BL45),.BLN(BLN45),.WL(WL164));
sram_cell_6t_5 inst_cell_164_46 (.BL(BL46),.BLN(BLN46),.WL(WL164));
sram_cell_6t_5 inst_cell_164_47 (.BL(BL47),.BLN(BLN47),.WL(WL164));
sram_cell_6t_5 inst_cell_164_48 (.BL(BL48),.BLN(BLN48),.WL(WL164));
sram_cell_6t_5 inst_cell_164_49 (.BL(BL49),.BLN(BLN49),.WL(WL164));
sram_cell_6t_5 inst_cell_164_50 (.BL(BL50),.BLN(BLN50),.WL(WL164));
sram_cell_6t_5 inst_cell_164_51 (.BL(BL51),.BLN(BLN51),.WL(WL164));
sram_cell_6t_5 inst_cell_164_52 (.BL(BL52),.BLN(BLN52),.WL(WL164));
sram_cell_6t_5 inst_cell_164_53 (.BL(BL53),.BLN(BLN53),.WL(WL164));
sram_cell_6t_5 inst_cell_164_54 (.BL(BL54),.BLN(BLN54),.WL(WL164));
sram_cell_6t_5 inst_cell_164_55 (.BL(BL55),.BLN(BLN55),.WL(WL164));
sram_cell_6t_5 inst_cell_164_56 (.BL(BL56),.BLN(BLN56),.WL(WL164));
sram_cell_6t_5 inst_cell_164_57 (.BL(BL57),.BLN(BLN57),.WL(WL164));
sram_cell_6t_5 inst_cell_164_58 (.BL(BL58),.BLN(BLN58),.WL(WL164));
sram_cell_6t_5 inst_cell_164_59 (.BL(BL59),.BLN(BLN59),.WL(WL164));
sram_cell_6t_5 inst_cell_164_60 (.BL(BL60),.BLN(BLN60),.WL(WL164));
sram_cell_6t_5 inst_cell_164_61 (.BL(BL61),.BLN(BLN61),.WL(WL164));
sram_cell_6t_5 inst_cell_164_62 (.BL(BL62),.BLN(BLN62),.WL(WL164));
sram_cell_6t_5 inst_cell_164_63 (.BL(BL63),.BLN(BLN63),.WL(WL164));
sram_cell_6t_5 inst_cell_164_64 (.BL(BL64),.BLN(BLN64),.WL(WL164));
sram_cell_6t_5 inst_cell_164_65 (.BL(BL65),.BLN(BLN65),.WL(WL164));
sram_cell_6t_5 inst_cell_164_66 (.BL(BL66),.BLN(BLN66),.WL(WL164));
sram_cell_6t_5 inst_cell_164_67 (.BL(BL67),.BLN(BLN67),.WL(WL164));
sram_cell_6t_5 inst_cell_164_68 (.BL(BL68),.BLN(BLN68),.WL(WL164));
sram_cell_6t_5 inst_cell_164_69 (.BL(BL69),.BLN(BLN69),.WL(WL164));
sram_cell_6t_5 inst_cell_164_70 (.BL(BL70),.BLN(BLN70),.WL(WL164));
sram_cell_6t_5 inst_cell_164_71 (.BL(BL71),.BLN(BLN71),.WL(WL164));
sram_cell_6t_5 inst_cell_164_72 (.BL(BL72),.BLN(BLN72),.WL(WL164));
sram_cell_6t_5 inst_cell_164_73 (.BL(BL73),.BLN(BLN73),.WL(WL164));
sram_cell_6t_5 inst_cell_164_74 (.BL(BL74),.BLN(BLN74),.WL(WL164));
sram_cell_6t_5 inst_cell_164_75 (.BL(BL75),.BLN(BLN75),.WL(WL164));
sram_cell_6t_5 inst_cell_164_76 (.BL(BL76),.BLN(BLN76),.WL(WL164));
sram_cell_6t_5 inst_cell_164_77 (.BL(BL77),.BLN(BLN77),.WL(WL164));
sram_cell_6t_5 inst_cell_164_78 (.BL(BL78),.BLN(BLN78),.WL(WL164));
sram_cell_6t_5 inst_cell_164_79 (.BL(BL79),.BLN(BLN79),.WL(WL164));
sram_cell_6t_5 inst_cell_164_80 (.BL(BL80),.BLN(BLN80),.WL(WL164));
sram_cell_6t_5 inst_cell_164_81 (.BL(BL81),.BLN(BLN81),.WL(WL164));
sram_cell_6t_5 inst_cell_164_82 (.BL(BL82),.BLN(BLN82),.WL(WL164));
sram_cell_6t_5 inst_cell_164_83 (.BL(BL83),.BLN(BLN83),.WL(WL164));
sram_cell_6t_5 inst_cell_164_84 (.BL(BL84),.BLN(BLN84),.WL(WL164));
sram_cell_6t_5 inst_cell_164_85 (.BL(BL85),.BLN(BLN85),.WL(WL164));
sram_cell_6t_5 inst_cell_164_86 (.BL(BL86),.BLN(BLN86),.WL(WL164));
sram_cell_6t_5 inst_cell_164_87 (.BL(BL87),.BLN(BLN87),.WL(WL164));
sram_cell_6t_5 inst_cell_164_88 (.BL(BL88),.BLN(BLN88),.WL(WL164));
sram_cell_6t_5 inst_cell_164_89 (.BL(BL89),.BLN(BLN89),.WL(WL164));
sram_cell_6t_5 inst_cell_164_90 (.BL(BL90),.BLN(BLN90),.WL(WL164));
sram_cell_6t_5 inst_cell_164_91 (.BL(BL91),.BLN(BLN91),.WL(WL164));
sram_cell_6t_5 inst_cell_164_92 (.BL(BL92),.BLN(BLN92),.WL(WL164));
sram_cell_6t_5 inst_cell_164_93 (.BL(BL93),.BLN(BLN93),.WL(WL164));
sram_cell_6t_5 inst_cell_164_94 (.BL(BL94),.BLN(BLN94),.WL(WL164));
sram_cell_6t_5 inst_cell_164_95 (.BL(BL95),.BLN(BLN95),.WL(WL164));
sram_cell_6t_5 inst_cell_164_96 (.BL(BL96),.BLN(BLN96),.WL(WL164));
sram_cell_6t_5 inst_cell_164_97 (.BL(BL97),.BLN(BLN97),.WL(WL164));
sram_cell_6t_5 inst_cell_164_98 (.BL(BL98),.BLN(BLN98),.WL(WL164));
sram_cell_6t_5 inst_cell_164_99 (.BL(BL99),.BLN(BLN99),.WL(WL164));
sram_cell_6t_5 inst_cell_164_100 (.BL(BL100),.BLN(BLN100),.WL(WL164));
sram_cell_6t_5 inst_cell_164_101 (.BL(BL101),.BLN(BLN101),.WL(WL164));
sram_cell_6t_5 inst_cell_164_102 (.BL(BL102),.BLN(BLN102),.WL(WL164));
sram_cell_6t_5 inst_cell_164_103 (.BL(BL103),.BLN(BLN103),.WL(WL164));
sram_cell_6t_5 inst_cell_164_104 (.BL(BL104),.BLN(BLN104),.WL(WL164));
sram_cell_6t_5 inst_cell_164_105 (.BL(BL105),.BLN(BLN105),.WL(WL164));
sram_cell_6t_5 inst_cell_164_106 (.BL(BL106),.BLN(BLN106),.WL(WL164));
sram_cell_6t_5 inst_cell_164_107 (.BL(BL107),.BLN(BLN107),.WL(WL164));
sram_cell_6t_5 inst_cell_164_108 (.BL(BL108),.BLN(BLN108),.WL(WL164));
sram_cell_6t_5 inst_cell_164_109 (.BL(BL109),.BLN(BLN109),.WL(WL164));
sram_cell_6t_5 inst_cell_164_110 (.BL(BL110),.BLN(BLN110),.WL(WL164));
sram_cell_6t_5 inst_cell_164_111 (.BL(BL111),.BLN(BLN111),.WL(WL164));
sram_cell_6t_5 inst_cell_164_112 (.BL(BL112),.BLN(BLN112),.WL(WL164));
sram_cell_6t_5 inst_cell_164_113 (.BL(BL113),.BLN(BLN113),.WL(WL164));
sram_cell_6t_5 inst_cell_164_114 (.BL(BL114),.BLN(BLN114),.WL(WL164));
sram_cell_6t_5 inst_cell_164_115 (.BL(BL115),.BLN(BLN115),.WL(WL164));
sram_cell_6t_5 inst_cell_164_116 (.BL(BL116),.BLN(BLN116),.WL(WL164));
sram_cell_6t_5 inst_cell_164_117 (.BL(BL117),.BLN(BLN117),.WL(WL164));
sram_cell_6t_5 inst_cell_164_118 (.BL(BL118),.BLN(BLN118),.WL(WL164));
sram_cell_6t_5 inst_cell_164_119 (.BL(BL119),.BLN(BLN119),.WL(WL164));
sram_cell_6t_5 inst_cell_164_120 (.BL(BL120),.BLN(BLN120),.WL(WL164));
sram_cell_6t_5 inst_cell_164_121 (.BL(BL121),.BLN(BLN121),.WL(WL164));
sram_cell_6t_5 inst_cell_164_122 (.BL(BL122),.BLN(BLN122),.WL(WL164));
sram_cell_6t_5 inst_cell_164_123 (.BL(BL123),.BLN(BLN123),.WL(WL164));
sram_cell_6t_5 inst_cell_164_124 (.BL(BL124),.BLN(BLN124),.WL(WL164));
sram_cell_6t_5 inst_cell_164_125 (.BL(BL125),.BLN(BLN125),.WL(WL164));
sram_cell_6t_5 inst_cell_164_126 (.BL(BL126),.BLN(BLN126),.WL(WL164));
sram_cell_6t_5 inst_cell_164_127 (.BL(BL127),.BLN(BLN127),.WL(WL164));
sram_cell_6t_5 inst_cell_165_0 (.BL(BL0),.BLN(BLN0),.WL(WL165));
sram_cell_6t_5 inst_cell_165_1 (.BL(BL1),.BLN(BLN1),.WL(WL165));
sram_cell_6t_5 inst_cell_165_2 (.BL(BL2),.BLN(BLN2),.WL(WL165));
sram_cell_6t_5 inst_cell_165_3 (.BL(BL3),.BLN(BLN3),.WL(WL165));
sram_cell_6t_5 inst_cell_165_4 (.BL(BL4),.BLN(BLN4),.WL(WL165));
sram_cell_6t_5 inst_cell_165_5 (.BL(BL5),.BLN(BLN5),.WL(WL165));
sram_cell_6t_5 inst_cell_165_6 (.BL(BL6),.BLN(BLN6),.WL(WL165));
sram_cell_6t_5 inst_cell_165_7 (.BL(BL7),.BLN(BLN7),.WL(WL165));
sram_cell_6t_5 inst_cell_165_8 (.BL(BL8),.BLN(BLN8),.WL(WL165));
sram_cell_6t_5 inst_cell_165_9 (.BL(BL9),.BLN(BLN9),.WL(WL165));
sram_cell_6t_5 inst_cell_165_10 (.BL(BL10),.BLN(BLN10),.WL(WL165));
sram_cell_6t_5 inst_cell_165_11 (.BL(BL11),.BLN(BLN11),.WL(WL165));
sram_cell_6t_5 inst_cell_165_12 (.BL(BL12),.BLN(BLN12),.WL(WL165));
sram_cell_6t_5 inst_cell_165_13 (.BL(BL13),.BLN(BLN13),.WL(WL165));
sram_cell_6t_5 inst_cell_165_14 (.BL(BL14),.BLN(BLN14),.WL(WL165));
sram_cell_6t_5 inst_cell_165_15 (.BL(BL15),.BLN(BLN15),.WL(WL165));
sram_cell_6t_5 inst_cell_165_16 (.BL(BL16),.BLN(BLN16),.WL(WL165));
sram_cell_6t_5 inst_cell_165_17 (.BL(BL17),.BLN(BLN17),.WL(WL165));
sram_cell_6t_5 inst_cell_165_18 (.BL(BL18),.BLN(BLN18),.WL(WL165));
sram_cell_6t_5 inst_cell_165_19 (.BL(BL19),.BLN(BLN19),.WL(WL165));
sram_cell_6t_5 inst_cell_165_20 (.BL(BL20),.BLN(BLN20),.WL(WL165));
sram_cell_6t_5 inst_cell_165_21 (.BL(BL21),.BLN(BLN21),.WL(WL165));
sram_cell_6t_5 inst_cell_165_22 (.BL(BL22),.BLN(BLN22),.WL(WL165));
sram_cell_6t_5 inst_cell_165_23 (.BL(BL23),.BLN(BLN23),.WL(WL165));
sram_cell_6t_5 inst_cell_165_24 (.BL(BL24),.BLN(BLN24),.WL(WL165));
sram_cell_6t_5 inst_cell_165_25 (.BL(BL25),.BLN(BLN25),.WL(WL165));
sram_cell_6t_5 inst_cell_165_26 (.BL(BL26),.BLN(BLN26),.WL(WL165));
sram_cell_6t_5 inst_cell_165_27 (.BL(BL27),.BLN(BLN27),.WL(WL165));
sram_cell_6t_5 inst_cell_165_28 (.BL(BL28),.BLN(BLN28),.WL(WL165));
sram_cell_6t_5 inst_cell_165_29 (.BL(BL29),.BLN(BLN29),.WL(WL165));
sram_cell_6t_5 inst_cell_165_30 (.BL(BL30),.BLN(BLN30),.WL(WL165));
sram_cell_6t_5 inst_cell_165_31 (.BL(BL31),.BLN(BLN31),.WL(WL165));
sram_cell_6t_5 inst_cell_165_32 (.BL(BL32),.BLN(BLN32),.WL(WL165));
sram_cell_6t_5 inst_cell_165_33 (.BL(BL33),.BLN(BLN33),.WL(WL165));
sram_cell_6t_5 inst_cell_165_34 (.BL(BL34),.BLN(BLN34),.WL(WL165));
sram_cell_6t_5 inst_cell_165_35 (.BL(BL35),.BLN(BLN35),.WL(WL165));
sram_cell_6t_5 inst_cell_165_36 (.BL(BL36),.BLN(BLN36),.WL(WL165));
sram_cell_6t_5 inst_cell_165_37 (.BL(BL37),.BLN(BLN37),.WL(WL165));
sram_cell_6t_5 inst_cell_165_38 (.BL(BL38),.BLN(BLN38),.WL(WL165));
sram_cell_6t_5 inst_cell_165_39 (.BL(BL39),.BLN(BLN39),.WL(WL165));
sram_cell_6t_5 inst_cell_165_40 (.BL(BL40),.BLN(BLN40),.WL(WL165));
sram_cell_6t_5 inst_cell_165_41 (.BL(BL41),.BLN(BLN41),.WL(WL165));
sram_cell_6t_5 inst_cell_165_42 (.BL(BL42),.BLN(BLN42),.WL(WL165));
sram_cell_6t_5 inst_cell_165_43 (.BL(BL43),.BLN(BLN43),.WL(WL165));
sram_cell_6t_5 inst_cell_165_44 (.BL(BL44),.BLN(BLN44),.WL(WL165));
sram_cell_6t_5 inst_cell_165_45 (.BL(BL45),.BLN(BLN45),.WL(WL165));
sram_cell_6t_5 inst_cell_165_46 (.BL(BL46),.BLN(BLN46),.WL(WL165));
sram_cell_6t_5 inst_cell_165_47 (.BL(BL47),.BLN(BLN47),.WL(WL165));
sram_cell_6t_5 inst_cell_165_48 (.BL(BL48),.BLN(BLN48),.WL(WL165));
sram_cell_6t_5 inst_cell_165_49 (.BL(BL49),.BLN(BLN49),.WL(WL165));
sram_cell_6t_5 inst_cell_165_50 (.BL(BL50),.BLN(BLN50),.WL(WL165));
sram_cell_6t_5 inst_cell_165_51 (.BL(BL51),.BLN(BLN51),.WL(WL165));
sram_cell_6t_5 inst_cell_165_52 (.BL(BL52),.BLN(BLN52),.WL(WL165));
sram_cell_6t_5 inst_cell_165_53 (.BL(BL53),.BLN(BLN53),.WL(WL165));
sram_cell_6t_5 inst_cell_165_54 (.BL(BL54),.BLN(BLN54),.WL(WL165));
sram_cell_6t_5 inst_cell_165_55 (.BL(BL55),.BLN(BLN55),.WL(WL165));
sram_cell_6t_5 inst_cell_165_56 (.BL(BL56),.BLN(BLN56),.WL(WL165));
sram_cell_6t_5 inst_cell_165_57 (.BL(BL57),.BLN(BLN57),.WL(WL165));
sram_cell_6t_5 inst_cell_165_58 (.BL(BL58),.BLN(BLN58),.WL(WL165));
sram_cell_6t_5 inst_cell_165_59 (.BL(BL59),.BLN(BLN59),.WL(WL165));
sram_cell_6t_5 inst_cell_165_60 (.BL(BL60),.BLN(BLN60),.WL(WL165));
sram_cell_6t_5 inst_cell_165_61 (.BL(BL61),.BLN(BLN61),.WL(WL165));
sram_cell_6t_5 inst_cell_165_62 (.BL(BL62),.BLN(BLN62),.WL(WL165));
sram_cell_6t_5 inst_cell_165_63 (.BL(BL63),.BLN(BLN63),.WL(WL165));
sram_cell_6t_5 inst_cell_165_64 (.BL(BL64),.BLN(BLN64),.WL(WL165));
sram_cell_6t_5 inst_cell_165_65 (.BL(BL65),.BLN(BLN65),.WL(WL165));
sram_cell_6t_5 inst_cell_165_66 (.BL(BL66),.BLN(BLN66),.WL(WL165));
sram_cell_6t_5 inst_cell_165_67 (.BL(BL67),.BLN(BLN67),.WL(WL165));
sram_cell_6t_5 inst_cell_165_68 (.BL(BL68),.BLN(BLN68),.WL(WL165));
sram_cell_6t_5 inst_cell_165_69 (.BL(BL69),.BLN(BLN69),.WL(WL165));
sram_cell_6t_5 inst_cell_165_70 (.BL(BL70),.BLN(BLN70),.WL(WL165));
sram_cell_6t_5 inst_cell_165_71 (.BL(BL71),.BLN(BLN71),.WL(WL165));
sram_cell_6t_5 inst_cell_165_72 (.BL(BL72),.BLN(BLN72),.WL(WL165));
sram_cell_6t_5 inst_cell_165_73 (.BL(BL73),.BLN(BLN73),.WL(WL165));
sram_cell_6t_5 inst_cell_165_74 (.BL(BL74),.BLN(BLN74),.WL(WL165));
sram_cell_6t_5 inst_cell_165_75 (.BL(BL75),.BLN(BLN75),.WL(WL165));
sram_cell_6t_5 inst_cell_165_76 (.BL(BL76),.BLN(BLN76),.WL(WL165));
sram_cell_6t_5 inst_cell_165_77 (.BL(BL77),.BLN(BLN77),.WL(WL165));
sram_cell_6t_5 inst_cell_165_78 (.BL(BL78),.BLN(BLN78),.WL(WL165));
sram_cell_6t_5 inst_cell_165_79 (.BL(BL79),.BLN(BLN79),.WL(WL165));
sram_cell_6t_5 inst_cell_165_80 (.BL(BL80),.BLN(BLN80),.WL(WL165));
sram_cell_6t_5 inst_cell_165_81 (.BL(BL81),.BLN(BLN81),.WL(WL165));
sram_cell_6t_5 inst_cell_165_82 (.BL(BL82),.BLN(BLN82),.WL(WL165));
sram_cell_6t_5 inst_cell_165_83 (.BL(BL83),.BLN(BLN83),.WL(WL165));
sram_cell_6t_5 inst_cell_165_84 (.BL(BL84),.BLN(BLN84),.WL(WL165));
sram_cell_6t_5 inst_cell_165_85 (.BL(BL85),.BLN(BLN85),.WL(WL165));
sram_cell_6t_5 inst_cell_165_86 (.BL(BL86),.BLN(BLN86),.WL(WL165));
sram_cell_6t_5 inst_cell_165_87 (.BL(BL87),.BLN(BLN87),.WL(WL165));
sram_cell_6t_5 inst_cell_165_88 (.BL(BL88),.BLN(BLN88),.WL(WL165));
sram_cell_6t_5 inst_cell_165_89 (.BL(BL89),.BLN(BLN89),.WL(WL165));
sram_cell_6t_5 inst_cell_165_90 (.BL(BL90),.BLN(BLN90),.WL(WL165));
sram_cell_6t_5 inst_cell_165_91 (.BL(BL91),.BLN(BLN91),.WL(WL165));
sram_cell_6t_5 inst_cell_165_92 (.BL(BL92),.BLN(BLN92),.WL(WL165));
sram_cell_6t_5 inst_cell_165_93 (.BL(BL93),.BLN(BLN93),.WL(WL165));
sram_cell_6t_5 inst_cell_165_94 (.BL(BL94),.BLN(BLN94),.WL(WL165));
sram_cell_6t_5 inst_cell_165_95 (.BL(BL95),.BLN(BLN95),.WL(WL165));
sram_cell_6t_5 inst_cell_165_96 (.BL(BL96),.BLN(BLN96),.WL(WL165));
sram_cell_6t_5 inst_cell_165_97 (.BL(BL97),.BLN(BLN97),.WL(WL165));
sram_cell_6t_5 inst_cell_165_98 (.BL(BL98),.BLN(BLN98),.WL(WL165));
sram_cell_6t_5 inst_cell_165_99 (.BL(BL99),.BLN(BLN99),.WL(WL165));
sram_cell_6t_5 inst_cell_165_100 (.BL(BL100),.BLN(BLN100),.WL(WL165));
sram_cell_6t_5 inst_cell_165_101 (.BL(BL101),.BLN(BLN101),.WL(WL165));
sram_cell_6t_5 inst_cell_165_102 (.BL(BL102),.BLN(BLN102),.WL(WL165));
sram_cell_6t_5 inst_cell_165_103 (.BL(BL103),.BLN(BLN103),.WL(WL165));
sram_cell_6t_5 inst_cell_165_104 (.BL(BL104),.BLN(BLN104),.WL(WL165));
sram_cell_6t_5 inst_cell_165_105 (.BL(BL105),.BLN(BLN105),.WL(WL165));
sram_cell_6t_5 inst_cell_165_106 (.BL(BL106),.BLN(BLN106),.WL(WL165));
sram_cell_6t_5 inst_cell_165_107 (.BL(BL107),.BLN(BLN107),.WL(WL165));
sram_cell_6t_5 inst_cell_165_108 (.BL(BL108),.BLN(BLN108),.WL(WL165));
sram_cell_6t_5 inst_cell_165_109 (.BL(BL109),.BLN(BLN109),.WL(WL165));
sram_cell_6t_5 inst_cell_165_110 (.BL(BL110),.BLN(BLN110),.WL(WL165));
sram_cell_6t_5 inst_cell_165_111 (.BL(BL111),.BLN(BLN111),.WL(WL165));
sram_cell_6t_5 inst_cell_165_112 (.BL(BL112),.BLN(BLN112),.WL(WL165));
sram_cell_6t_5 inst_cell_165_113 (.BL(BL113),.BLN(BLN113),.WL(WL165));
sram_cell_6t_5 inst_cell_165_114 (.BL(BL114),.BLN(BLN114),.WL(WL165));
sram_cell_6t_5 inst_cell_165_115 (.BL(BL115),.BLN(BLN115),.WL(WL165));
sram_cell_6t_5 inst_cell_165_116 (.BL(BL116),.BLN(BLN116),.WL(WL165));
sram_cell_6t_5 inst_cell_165_117 (.BL(BL117),.BLN(BLN117),.WL(WL165));
sram_cell_6t_5 inst_cell_165_118 (.BL(BL118),.BLN(BLN118),.WL(WL165));
sram_cell_6t_5 inst_cell_165_119 (.BL(BL119),.BLN(BLN119),.WL(WL165));
sram_cell_6t_5 inst_cell_165_120 (.BL(BL120),.BLN(BLN120),.WL(WL165));
sram_cell_6t_5 inst_cell_165_121 (.BL(BL121),.BLN(BLN121),.WL(WL165));
sram_cell_6t_5 inst_cell_165_122 (.BL(BL122),.BLN(BLN122),.WL(WL165));
sram_cell_6t_5 inst_cell_165_123 (.BL(BL123),.BLN(BLN123),.WL(WL165));
sram_cell_6t_5 inst_cell_165_124 (.BL(BL124),.BLN(BLN124),.WL(WL165));
sram_cell_6t_5 inst_cell_165_125 (.BL(BL125),.BLN(BLN125),.WL(WL165));
sram_cell_6t_5 inst_cell_165_126 (.BL(BL126),.BLN(BLN126),.WL(WL165));
sram_cell_6t_5 inst_cell_165_127 (.BL(BL127),.BLN(BLN127),.WL(WL165));
sram_cell_6t_5 inst_cell_166_0 (.BL(BL0),.BLN(BLN0),.WL(WL166));
sram_cell_6t_5 inst_cell_166_1 (.BL(BL1),.BLN(BLN1),.WL(WL166));
sram_cell_6t_5 inst_cell_166_2 (.BL(BL2),.BLN(BLN2),.WL(WL166));
sram_cell_6t_5 inst_cell_166_3 (.BL(BL3),.BLN(BLN3),.WL(WL166));
sram_cell_6t_5 inst_cell_166_4 (.BL(BL4),.BLN(BLN4),.WL(WL166));
sram_cell_6t_5 inst_cell_166_5 (.BL(BL5),.BLN(BLN5),.WL(WL166));
sram_cell_6t_5 inst_cell_166_6 (.BL(BL6),.BLN(BLN6),.WL(WL166));
sram_cell_6t_5 inst_cell_166_7 (.BL(BL7),.BLN(BLN7),.WL(WL166));
sram_cell_6t_5 inst_cell_166_8 (.BL(BL8),.BLN(BLN8),.WL(WL166));
sram_cell_6t_5 inst_cell_166_9 (.BL(BL9),.BLN(BLN9),.WL(WL166));
sram_cell_6t_5 inst_cell_166_10 (.BL(BL10),.BLN(BLN10),.WL(WL166));
sram_cell_6t_5 inst_cell_166_11 (.BL(BL11),.BLN(BLN11),.WL(WL166));
sram_cell_6t_5 inst_cell_166_12 (.BL(BL12),.BLN(BLN12),.WL(WL166));
sram_cell_6t_5 inst_cell_166_13 (.BL(BL13),.BLN(BLN13),.WL(WL166));
sram_cell_6t_5 inst_cell_166_14 (.BL(BL14),.BLN(BLN14),.WL(WL166));
sram_cell_6t_5 inst_cell_166_15 (.BL(BL15),.BLN(BLN15),.WL(WL166));
sram_cell_6t_5 inst_cell_166_16 (.BL(BL16),.BLN(BLN16),.WL(WL166));
sram_cell_6t_5 inst_cell_166_17 (.BL(BL17),.BLN(BLN17),.WL(WL166));
sram_cell_6t_5 inst_cell_166_18 (.BL(BL18),.BLN(BLN18),.WL(WL166));
sram_cell_6t_5 inst_cell_166_19 (.BL(BL19),.BLN(BLN19),.WL(WL166));
sram_cell_6t_5 inst_cell_166_20 (.BL(BL20),.BLN(BLN20),.WL(WL166));
sram_cell_6t_5 inst_cell_166_21 (.BL(BL21),.BLN(BLN21),.WL(WL166));
sram_cell_6t_5 inst_cell_166_22 (.BL(BL22),.BLN(BLN22),.WL(WL166));
sram_cell_6t_5 inst_cell_166_23 (.BL(BL23),.BLN(BLN23),.WL(WL166));
sram_cell_6t_5 inst_cell_166_24 (.BL(BL24),.BLN(BLN24),.WL(WL166));
sram_cell_6t_5 inst_cell_166_25 (.BL(BL25),.BLN(BLN25),.WL(WL166));
sram_cell_6t_5 inst_cell_166_26 (.BL(BL26),.BLN(BLN26),.WL(WL166));
sram_cell_6t_5 inst_cell_166_27 (.BL(BL27),.BLN(BLN27),.WL(WL166));
sram_cell_6t_5 inst_cell_166_28 (.BL(BL28),.BLN(BLN28),.WL(WL166));
sram_cell_6t_5 inst_cell_166_29 (.BL(BL29),.BLN(BLN29),.WL(WL166));
sram_cell_6t_5 inst_cell_166_30 (.BL(BL30),.BLN(BLN30),.WL(WL166));
sram_cell_6t_5 inst_cell_166_31 (.BL(BL31),.BLN(BLN31),.WL(WL166));
sram_cell_6t_5 inst_cell_166_32 (.BL(BL32),.BLN(BLN32),.WL(WL166));
sram_cell_6t_5 inst_cell_166_33 (.BL(BL33),.BLN(BLN33),.WL(WL166));
sram_cell_6t_5 inst_cell_166_34 (.BL(BL34),.BLN(BLN34),.WL(WL166));
sram_cell_6t_5 inst_cell_166_35 (.BL(BL35),.BLN(BLN35),.WL(WL166));
sram_cell_6t_5 inst_cell_166_36 (.BL(BL36),.BLN(BLN36),.WL(WL166));
sram_cell_6t_5 inst_cell_166_37 (.BL(BL37),.BLN(BLN37),.WL(WL166));
sram_cell_6t_5 inst_cell_166_38 (.BL(BL38),.BLN(BLN38),.WL(WL166));
sram_cell_6t_5 inst_cell_166_39 (.BL(BL39),.BLN(BLN39),.WL(WL166));
sram_cell_6t_5 inst_cell_166_40 (.BL(BL40),.BLN(BLN40),.WL(WL166));
sram_cell_6t_5 inst_cell_166_41 (.BL(BL41),.BLN(BLN41),.WL(WL166));
sram_cell_6t_5 inst_cell_166_42 (.BL(BL42),.BLN(BLN42),.WL(WL166));
sram_cell_6t_5 inst_cell_166_43 (.BL(BL43),.BLN(BLN43),.WL(WL166));
sram_cell_6t_5 inst_cell_166_44 (.BL(BL44),.BLN(BLN44),.WL(WL166));
sram_cell_6t_5 inst_cell_166_45 (.BL(BL45),.BLN(BLN45),.WL(WL166));
sram_cell_6t_5 inst_cell_166_46 (.BL(BL46),.BLN(BLN46),.WL(WL166));
sram_cell_6t_5 inst_cell_166_47 (.BL(BL47),.BLN(BLN47),.WL(WL166));
sram_cell_6t_5 inst_cell_166_48 (.BL(BL48),.BLN(BLN48),.WL(WL166));
sram_cell_6t_5 inst_cell_166_49 (.BL(BL49),.BLN(BLN49),.WL(WL166));
sram_cell_6t_5 inst_cell_166_50 (.BL(BL50),.BLN(BLN50),.WL(WL166));
sram_cell_6t_5 inst_cell_166_51 (.BL(BL51),.BLN(BLN51),.WL(WL166));
sram_cell_6t_5 inst_cell_166_52 (.BL(BL52),.BLN(BLN52),.WL(WL166));
sram_cell_6t_5 inst_cell_166_53 (.BL(BL53),.BLN(BLN53),.WL(WL166));
sram_cell_6t_5 inst_cell_166_54 (.BL(BL54),.BLN(BLN54),.WL(WL166));
sram_cell_6t_5 inst_cell_166_55 (.BL(BL55),.BLN(BLN55),.WL(WL166));
sram_cell_6t_5 inst_cell_166_56 (.BL(BL56),.BLN(BLN56),.WL(WL166));
sram_cell_6t_5 inst_cell_166_57 (.BL(BL57),.BLN(BLN57),.WL(WL166));
sram_cell_6t_5 inst_cell_166_58 (.BL(BL58),.BLN(BLN58),.WL(WL166));
sram_cell_6t_5 inst_cell_166_59 (.BL(BL59),.BLN(BLN59),.WL(WL166));
sram_cell_6t_5 inst_cell_166_60 (.BL(BL60),.BLN(BLN60),.WL(WL166));
sram_cell_6t_5 inst_cell_166_61 (.BL(BL61),.BLN(BLN61),.WL(WL166));
sram_cell_6t_5 inst_cell_166_62 (.BL(BL62),.BLN(BLN62),.WL(WL166));
sram_cell_6t_5 inst_cell_166_63 (.BL(BL63),.BLN(BLN63),.WL(WL166));
sram_cell_6t_5 inst_cell_166_64 (.BL(BL64),.BLN(BLN64),.WL(WL166));
sram_cell_6t_5 inst_cell_166_65 (.BL(BL65),.BLN(BLN65),.WL(WL166));
sram_cell_6t_5 inst_cell_166_66 (.BL(BL66),.BLN(BLN66),.WL(WL166));
sram_cell_6t_5 inst_cell_166_67 (.BL(BL67),.BLN(BLN67),.WL(WL166));
sram_cell_6t_5 inst_cell_166_68 (.BL(BL68),.BLN(BLN68),.WL(WL166));
sram_cell_6t_5 inst_cell_166_69 (.BL(BL69),.BLN(BLN69),.WL(WL166));
sram_cell_6t_5 inst_cell_166_70 (.BL(BL70),.BLN(BLN70),.WL(WL166));
sram_cell_6t_5 inst_cell_166_71 (.BL(BL71),.BLN(BLN71),.WL(WL166));
sram_cell_6t_5 inst_cell_166_72 (.BL(BL72),.BLN(BLN72),.WL(WL166));
sram_cell_6t_5 inst_cell_166_73 (.BL(BL73),.BLN(BLN73),.WL(WL166));
sram_cell_6t_5 inst_cell_166_74 (.BL(BL74),.BLN(BLN74),.WL(WL166));
sram_cell_6t_5 inst_cell_166_75 (.BL(BL75),.BLN(BLN75),.WL(WL166));
sram_cell_6t_5 inst_cell_166_76 (.BL(BL76),.BLN(BLN76),.WL(WL166));
sram_cell_6t_5 inst_cell_166_77 (.BL(BL77),.BLN(BLN77),.WL(WL166));
sram_cell_6t_5 inst_cell_166_78 (.BL(BL78),.BLN(BLN78),.WL(WL166));
sram_cell_6t_5 inst_cell_166_79 (.BL(BL79),.BLN(BLN79),.WL(WL166));
sram_cell_6t_5 inst_cell_166_80 (.BL(BL80),.BLN(BLN80),.WL(WL166));
sram_cell_6t_5 inst_cell_166_81 (.BL(BL81),.BLN(BLN81),.WL(WL166));
sram_cell_6t_5 inst_cell_166_82 (.BL(BL82),.BLN(BLN82),.WL(WL166));
sram_cell_6t_5 inst_cell_166_83 (.BL(BL83),.BLN(BLN83),.WL(WL166));
sram_cell_6t_5 inst_cell_166_84 (.BL(BL84),.BLN(BLN84),.WL(WL166));
sram_cell_6t_5 inst_cell_166_85 (.BL(BL85),.BLN(BLN85),.WL(WL166));
sram_cell_6t_5 inst_cell_166_86 (.BL(BL86),.BLN(BLN86),.WL(WL166));
sram_cell_6t_5 inst_cell_166_87 (.BL(BL87),.BLN(BLN87),.WL(WL166));
sram_cell_6t_5 inst_cell_166_88 (.BL(BL88),.BLN(BLN88),.WL(WL166));
sram_cell_6t_5 inst_cell_166_89 (.BL(BL89),.BLN(BLN89),.WL(WL166));
sram_cell_6t_5 inst_cell_166_90 (.BL(BL90),.BLN(BLN90),.WL(WL166));
sram_cell_6t_5 inst_cell_166_91 (.BL(BL91),.BLN(BLN91),.WL(WL166));
sram_cell_6t_5 inst_cell_166_92 (.BL(BL92),.BLN(BLN92),.WL(WL166));
sram_cell_6t_5 inst_cell_166_93 (.BL(BL93),.BLN(BLN93),.WL(WL166));
sram_cell_6t_5 inst_cell_166_94 (.BL(BL94),.BLN(BLN94),.WL(WL166));
sram_cell_6t_5 inst_cell_166_95 (.BL(BL95),.BLN(BLN95),.WL(WL166));
sram_cell_6t_5 inst_cell_166_96 (.BL(BL96),.BLN(BLN96),.WL(WL166));
sram_cell_6t_5 inst_cell_166_97 (.BL(BL97),.BLN(BLN97),.WL(WL166));
sram_cell_6t_5 inst_cell_166_98 (.BL(BL98),.BLN(BLN98),.WL(WL166));
sram_cell_6t_5 inst_cell_166_99 (.BL(BL99),.BLN(BLN99),.WL(WL166));
sram_cell_6t_5 inst_cell_166_100 (.BL(BL100),.BLN(BLN100),.WL(WL166));
sram_cell_6t_5 inst_cell_166_101 (.BL(BL101),.BLN(BLN101),.WL(WL166));
sram_cell_6t_5 inst_cell_166_102 (.BL(BL102),.BLN(BLN102),.WL(WL166));
sram_cell_6t_5 inst_cell_166_103 (.BL(BL103),.BLN(BLN103),.WL(WL166));
sram_cell_6t_5 inst_cell_166_104 (.BL(BL104),.BLN(BLN104),.WL(WL166));
sram_cell_6t_5 inst_cell_166_105 (.BL(BL105),.BLN(BLN105),.WL(WL166));
sram_cell_6t_5 inst_cell_166_106 (.BL(BL106),.BLN(BLN106),.WL(WL166));
sram_cell_6t_5 inst_cell_166_107 (.BL(BL107),.BLN(BLN107),.WL(WL166));
sram_cell_6t_5 inst_cell_166_108 (.BL(BL108),.BLN(BLN108),.WL(WL166));
sram_cell_6t_5 inst_cell_166_109 (.BL(BL109),.BLN(BLN109),.WL(WL166));
sram_cell_6t_5 inst_cell_166_110 (.BL(BL110),.BLN(BLN110),.WL(WL166));
sram_cell_6t_5 inst_cell_166_111 (.BL(BL111),.BLN(BLN111),.WL(WL166));
sram_cell_6t_5 inst_cell_166_112 (.BL(BL112),.BLN(BLN112),.WL(WL166));
sram_cell_6t_5 inst_cell_166_113 (.BL(BL113),.BLN(BLN113),.WL(WL166));
sram_cell_6t_5 inst_cell_166_114 (.BL(BL114),.BLN(BLN114),.WL(WL166));
sram_cell_6t_5 inst_cell_166_115 (.BL(BL115),.BLN(BLN115),.WL(WL166));
sram_cell_6t_5 inst_cell_166_116 (.BL(BL116),.BLN(BLN116),.WL(WL166));
sram_cell_6t_5 inst_cell_166_117 (.BL(BL117),.BLN(BLN117),.WL(WL166));
sram_cell_6t_5 inst_cell_166_118 (.BL(BL118),.BLN(BLN118),.WL(WL166));
sram_cell_6t_5 inst_cell_166_119 (.BL(BL119),.BLN(BLN119),.WL(WL166));
sram_cell_6t_5 inst_cell_166_120 (.BL(BL120),.BLN(BLN120),.WL(WL166));
sram_cell_6t_5 inst_cell_166_121 (.BL(BL121),.BLN(BLN121),.WL(WL166));
sram_cell_6t_5 inst_cell_166_122 (.BL(BL122),.BLN(BLN122),.WL(WL166));
sram_cell_6t_5 inst_cell_166_123 (.BL(BL123),.BLN(BLN123),.WL(WL166));
sram_cell_6t_5 inst_cell_166_124 (.BL(BL124),.BLN(BLN124),.WL(WL166));
sram_cell_6t_5 inst_cell_166_125 (.BL(BL125),.BLN(BLN125),.WL(WL166));
sram_cell_6t_5 inst_cell_166_126 (.BL(BL126),.BLN(BLN126),.WL(WL166));
sram_cell_6t_5 inst_cell_166_127 (.BL(BL127),.BLN(BLN127),.WL(WL166));
sram_cell_6t_5 inst_cell_167_0 (.BL(BL0),.BLN(BLN0),.WL(WL167));
sram_cell_6t_5 inst_cell_167_1 (.BL(BL1),.BLN(BLN1),.WL(WL167));
sram_cell_6t_5 inst_cell_167_2 (.BL(BL2),.BLN(BLN2),.WL(WL167));
sram_cell_6t_5 inst_cell_167_3 (.BL(BL3),.BLN(BLN3),.WL(WL167));
sram_cell_6t_5 inst_cell_167_4 (.BL(BL4),.BLN(BLN4),.WL(WL167));
sram_cell_6t_5 inst_cell_167_5 (.BL(BL5),.BLN(BLN5),.WL(WL167));
sram_cell_6t_5 inst_cell_167_6 (.BL(BL6),.BLN(BLN6),.WL(WL167));
sram_cell_6t_5 inst_cell_167_7 (.BL(BL7),.BLN(BLN7),.WL(WL167));
sram_cell_6t_5 inst_cell_167_8 (.BL(BL8),.BLN(BLN8),.WL(WL167));
sram_cell_6t_5 inst_cell_167_9 (.BL(BL9),.BLN(BLN9),.WL(WL167));
sram_cell_6t_5 inst_cell_167_10 (.BL(BL10),.BLN(BLN10),.WL(WL167));
sram_cell_6t_5 inst_cell_167_11 (.BL(BL11),.BLN(BLN11),.WL(WL167));
sram_cell_6t_5 inst_cell_167_12 (.BL(BL12),.BLN(BLN12),.WL(WL167));
sram_cell_6t_5 inst_cell_167_13 (.BL(BL13),.BLN(BLN13),.WL(WL167));
sram_cell_6t_5 inst_cell_167_14 (.BL(BL14),.BLN(BLN14),.WL(WL167));
sram_cell_6t_5 inst_cell_167_15 (.BL(BL15),.BLN(BLN15),.WL(WL167));
sram_cell_6t_5 inst_cell_167_16 (.BL(BL16),.BLN(BLN16),.WL(WL167));
sram_cell_6t_5 inst_cell_167_17 (.BL(BL17),.BLN(BLN17),.WL(WL167));
sram_cell_6t_5 inst_cell_167_18 (.BL(BL18),.BLN(BLN18),.WL(WL167));
sram_cell_6t_5 inst_cell_167_19 (.BL(BL19),.BLN(BLN19),.WL(WL167));
sram_cell_6t_5 inst_cell_167_20 (.BL(BL20),.BLN(BLN20),.WL(WL167));
sram_cell_6t_5 inst_cell_167_21 (.BL(BL21),.BLN(BLN21),.WL(WL167));
sram_cell_6t_5 inst_cell_167_22 (.BL(BL22),.BLN(BLN22),.WL(WL167));
sram_cell_6t_5 inst_cell_167_23 (.BL(BL23),.BLN(BLN23),.WL(WL167));
sram_cell_6t_5 inst_cell_167_24 (.BL(BL24),.BLN(BLN24),.WL(WL167));
sram_cell_6t_5 inst_cell_167_25 (.BL(BL25),.BLN(BLN25),.WL(WL167));
sram_cell_6t_5 inst_cell_167_26 (.BL(BL26),.BLN(BLN26),.WL(WL167));
sram_cell_6t_5 inst_cell_167_27 (.BL(BL27),.BLN(BLN27),.WL(WL167));
sram_cell_6t_5 inst_cell_167_28 (.BL(BL28),.BLN(BLN28),.WL(WL167));
sram_cell_6t_5 inst_cell_167_29 (.BL(BL29),.BLN(BLN29),.WL(WL167));
sram_cell_6t_5 inst_cell_167_30 (.BL(BL30),.BLN(BLN30),.WL(WL167));
sram_cell_6t_5 inst_cell_167_31 (.BL(BL31),.BLN(BLN31),.WL(WL167));
sram_cell_6t_5 inst_cell_167_32 (.BL(BL32),.BLN(BLN32),.WL(WL167));
sram_cell_6t_5 inst_cell_167_33 (.BL(BL33),.BLN(BLN33),.WL(WL167));
sram_cell_6t_5 inst_cell_167_34 (.BL(BL34),.BLN(BLN34),.WL(WL167));
sram_cell_6t_5 inst_cell_167_35 (.BL(BL35),.BLN(BLN35),.WL(WL167));
sram_cell_6t_5 inst_cell_167_36 (.BL(BL36),.BLN(BLN36),.WL(WL167));
sram_cell_6t_5 inst_cell_167_37 (.BL(BL37),.BLN(BLN37),.WL(WL167));
sram_cell_6t_5 inst_cell_167_38 (.BL(BL38),.BLN(BLN38),.WL(WL167));
sram_cell_6t_5 inst_cell_167_39 (.BL(BL39),.BLN(BLN39),.WL(WL167));
sram_cell_6t_5 inst_cell_167_40 (.BL(BL40),.BLN(BLN40),.WL(WL167));
sram_cell_6t_5 inst_cell_167_41 (.BL(BL41),.BLN(BLN41),.WL(WL167));
sram_cell_6t_5 inst_cell_167_42 (.BL(BL42),.BLN(BLN42),.WL(WL167));
sram_cell_6t_5 inst_cell_167_43 (.BL(BL43),.BLN(BLN43),.WL(WL167));
sram_cell_6t_5 inst_cell_167_44 (.BL(BL44),.BLN(BLN44),.WL(WL167));
sram_cell_6t_5 inst_cell_167_45 (.BL(BL45),.BLN(BLN45),.WL(WL167));
sram_cell_6t_5 inst_cell_167_46 (.BL(BL46),.BLN(BLN46),.WL(WL167));
sram_cell_6t_5 inst_cell_167_47 (.BL(BL47),.BLN(BLN47),.WL(WL167));
sram_cell_6t_5 inst_cell_167_48 (.BL(BL48),.BLN(BLN48),.WL(WL167));
sram_cell_6t_5 inst_cell_167_49 (.BL(BL49),.BLN(BLN49),.WL(WL167));
sram_cell_6t_5 inst_cell_167_50 (.BL(BL50),.BLN(BLN50),.WL(WL167));
sram_cell_6t_5 inst_cell_167_51 (.BL(BL51),.BLN(BLN51),.WL(WL167));
sram_cell_6t_5 inst_cell_167_52 (.BL(BL52),.BLN(BLN52),.WL(WL167));
sram_cell_6t_5 inst_cell_167_53 (.BL(BL53),.BLN(BLN53),.WL(WL167));
sram_cell_6t_5 inst_cell_167_54 (.BL(BL54),.BLN(BLN54),.WL(WL167));
sram_cell_6t_5 inst_cell_167_55 (.BL(BL55),.BLN(BLN55),.WL(WL167));
sram_cell_6t_5 inst_cell_167_56 (.BL(BL56),.BLN(BLN56),.WL(WL167));
sram_cell_6t_5 inst_cell_167_57 (.BL(BL57),.BLN(BLN57),.WL(WL167));
sram_cell_6t_5 inst_cell_167_58 (.BL(BL58),.BLN(BLN58),.WL(WL167));
sram_cell_6t_5 inst_cell_167_59 (.BL(BL59),.BLN(BLN59),.WL(WL167));
sram_cell_6t_5 inst_cell_167_60 (.BL(BL60),.BLN(BLN60),.WL(WL167));
sram_cell_6t_5 inst_cell_167_61 (.BL(BL61),.BLN(BLN61),.WL(WL167));
sram_cell_6t_5 inst_cell_167_62 (.BL(BL62),.BLN(BLN62),.WL(WL167));
sram_cell_6t_5 inst_cell_167_63 (.BL(BL63),.BLN(BLN63),.WL(WL167));
sram_cell_6t_5 inst_cell_167_64 (.BL(BL64),.BLN(BLN64),.WL(WL167));
sram_cell_6t_5 inst_cell_167_65 (.BL(BL65),.BLN(BLN65),.WL(WL167));
sram_cell_6t_5 inst_cell_167_66 (.BL(BL66),.BLN(BLN66),.WL(WL167));
sram_cell_6t_5 inst_cell_167_67 (.BL(BL67),.BLN(BLN67),.WL(WL167));
sram_cell_6t_5 inst_cell_167_68 (.BL(BL68),.BLN(BLN68),.WL(WL167));
sram_cell_6t_5 inst_cell_167_69 (.BL(BL69),.BLN(BLN69),.WL(WL167));
sram_cell_6t_5 inst_cell_167_70 (.BL(BL70),.BLN(BLN70),.WL(WL167));
sram_cell_6t_5 inst_cell_167_71 (.BL(BL71),.BLN(BLN71),.WL(WL167));
sram_cell_6t_5 inst_cell_167_72 (.BL(BL72),.BLN(BLN72),.WL(WL167));
sram_cell_6t_5 inst_cell_167_73 (.BL(BL73),.BLN(BLN73),.WL(WL167));
sram_cell_6t_5 inst_cell_167_74 (.BL(BL74),.BLN(BLN74),.WL(WL167));
sram_cell_6t_5 inst_cell_167_75 (.BL(BL75),.BLN(BLN75),.WL(WL167));
sram_cell_6t_5 inst_cell_167_76 (.BL(BL76),.BLN(BLN76),.WL(WL167));
sram_cell_6t_5 inst_cell_167_77 (.BL(BL77),.BLN(BLN77),.WL(WL167));
sram_cell_6t_5 inst_cell_167_78 (.BL(BL78),.BLN(BLN78),.WL(WL167));
sram_cell_6t_5 inst_cell_167_79 (.BL(BL79),.BLN(BLN79),.WL(WL167));
sram_cell_6t_5 inst_cell_167_80 (.BL(BL80),.BLN(BLN80),.WL(WL167));
sram_cell_6t_5 inst_cell_167_81 (.BL(BL81),.BLN(BLN81),.WL(WL167));
sram_cell_6t_5 inst_cell_167_82 (.BL(BL82),.BLN(BLN82),.WL(WL167));
sram_cell_6t_5 inst_cell_167_83 (.BL(BL83),.BLN(BLN83),.WL(WL167));
sram_cell_6t_5 inst_cell_167_84 (.BL(BL84),.BLN(BLN84),.WL(WL167));
sram_cell_6t_5 inst_cell_167_85 (.BL(BL85),.BLN(BLN85),.WL(WL167));
sram_cell_6t_5 inst_cell_167_86 (.BL(BL86),.BLN(BLN86),.WL(WL167));
sram_cell_6t_5 inst_cell_167_87 (.BL(BL87),.BLN(BLN87),.WL(WL167));
sram_cell_6t_5 inst_cell_167_88 (.BL(BL88),.BLN(BLN88),.WL(WL167));
sram_cell_6t_5 inst_cell_167_89 (.BL(BL89),.BLN(BLN89),.WL(WL167));
sram_cell_6t_5 inst_cell_167_90 (.BL(BL90),.BLN(BLN90),.WL(WL167));
sram_cell_6t_5 inst_cell_167_91 (.BL(BL91),.BLN(BLN91),.WL(WL167));
sram_cell_6t_5 inst_cell_167_92 (.BL(BL92),.BLN(BLN92),.WL(WL167));
sram_cell_6t_5 inst_cell_167_93 (.BL(BL93),.BLN(BLN93),.WL(WL167));
sram_cell_6t_5 inst_cell_167_94 (.BL(BL94),.BLN(BLN94),.WL(WL167));
sram_cell_6t_5 inst_cell_167_95 (.BL(BL95),.BLN(BLN95),.WL(WL167));
sram_cell_6t_5 inst_cell_167_96 (.BL(BL96),.BLN(BLN96),.WL(WL167));
sram_cell_6t_5 inst_cell_167_97 (.BL(BL97),.BLN(BLN97),.WL(WL167));
sram_cell_6t_5 inst_cell_167_98 (.BL(BL98),.BLN(BLN98),.WL(WL167));
sram_cell_6t_5 inst_cell_167_99 (.BL(BL99),.BLN(BLN99),.WL(WL167));
sram_cell_6t_5 inst_cell_167_100 (.BL(BL100),.BLN(BLN100),.WL(WL167));
sram_cell_6t_5 inst_cell_167_101 (.BL(BL101),.BLN(BLN101),.WL(WL167));
sram_cell_6t_5 inst_cell_167_102 (.BL(BL102),.BLN(BLN102),.WL(WL167));
sram_cell_6t_5 inst_cell_167_103 (.BL(BL103),.BLN(BLN103),.WL(WL167));
sram_cell_6t_5 inst_cell_167_104 (.BL(BL104),.BLN(BLN104),.WL(WL167));
sram_cell_6t_5 inst_cell_167_105 (.BL(BL105),.BLN(BLN105),.WL(WL167));
sram_cell_6t_5 inst_cell_167_106 (.BL(BL106),.BLN(BLN106),.WL(WL167));
sram_cell_6t_5 inst_cell_167_107 (.BL(BL107),.BLN(BLN107),.WL(WL167));
sram_cell_6t_5 inst_cell_167_108 (.BL(BL108),.BLN(BLN108),.WL(WL167));
sram_cell_6t_5 inst_cell_167_109 (.BL(BL109),.BLN(BLN109),.WL(WL167));
sram_cell_6t_5 inst_cell_167_110 (.BL(BL110),.BLN(BLN110),.WL(WL167));
sram_cell_6t_5 inst_cell_167_111 (.BL(BL111),.BLN(BLN111),.WL(WL167));
sram_cell_6t_5 inst_cell_167_112 (.BL(BL112),.BLN(BLN112),.WL(WL167));
sram_cell_6t_5 inst_cell_167_113 (.BL(BL113),.BLN(BLN113),.WL(WL167));
sram_cell_6t_5 inst_cell_167_114 (.BL(BL114),.BLN(BLN114),.WL(WL167));
sram_cell_6t_5 inst_cell_167_115 (.BL(BL115),.BLN(BLN115),.WL(WL167));
sram_cell_6t_5 inst_cell_167_116 (.BL(BL116),.BLN(BLN116),.WL(WL167));
sram_cell_6t_5 inst_cell_167_117 (.BL(BL117),.BLN(BLN117),.WL(WL167));
sram_cell_6t_5 inst_cell_167_118 (.BL(BL118),.BLN(BLN118),.WL(WL167));
sram_cell_6t_5 inst_cell_167_119 (.BL(BL119),.BLN(BLN119),.WL(WL167));
sram_cell_6t_5 inst_cell_167_120 (.BL(BL120),.BLN(BLN120),.WL(WL167));
sram_cell_6t_5 inst_cell_167_121 (.BL(BL121),.BLN(BLN121),.WL(WL167));
sram_cell_6t_5 inst_cell_167_122 (.BL(BL122),.BLN(BLN122),.WL(WL167));
sram_cell_6t_5 inst_cell_167_123 (.BL(BL123),.BLN(BLN123),.WL(WL167));
sram_cell_6t_5 inst_cell_167_124 (.BL(BL124),.BLN(BLN124),.WL(WL167));
sram_cell_6t_5 inst_cell_167_125 (.BL(BL125),.BLN(BLN125),.WL(WL167));
sram_cell_6t_5 inst_cell_167_126 (.BL(BL126),.BLN(BLN126),.WL(WL167));
sram_cell_6t_5 inst_cell_167_127 (.BL(BL127),.BLN(BLN127),.WL(WL167));
sram_cell_6t_5 inst_cell_168_0 (.BL(BL0),.BLN(BLN0),.WL(WL168));
sram_cell_6t_5 inst_cell_168_1 (.BL(BL1),.BLN(BLN1),.WL(WL168));
sram_cell_6t_5 inst_cell_168_2 (.BL(BL2),.BLN(BLN2),.WL(WL168));
sram_cell_6t_5 inst_cell_168_3 (.BL(BL3),.BLN(BLN3),.WL(WL168));
sram_cell_6t_5 inst_cell_168_4 (.BL(BL4),.BLN(BLN4),.WL(WL168));
sram_cell_6t_5 inst_cell_168_5 (.BL(BL5),.BLN(BLN5),.WL(WL168));
sram_cell_6t_5 inst_cell_168_6 (.BL(BL6),.BLN(BLN6),.WL(WL168));
sram_cell_6t_5 inst_cell_168_7 (.BL(BL7),.BLN(BLN7),.WL(WL168));
sram_cell_6t_5 inst_cell_168_8 (.BL(BL8),.BLN(BLN8),.WL(WL168));
sram_cell_6t_5 inst_cell_168_9 (.BL(BL9),.BLN(BLN9),.WL(WL168));
sram_cell_6t_5 inst_cell_168_10 (.BL(BL10),.BLN(BLN10),.WL(WL168));
sram_cell_6t_5 inst_cell_168_11 (.BL(BL11),.BLN(BLN11),.WL(WL168));
sram_cell_6t_5 inst_cell_168_12 (.BL(BL12),.BLN(BLN12),.WL(WL168));
sram_cell_6t_5 inst_cell_168_13 (.BL(BL13),.BLN(BLN13),.WL(WL168));
sram_cell_6t_5 inst_cell_168_14 (.BL(BL14),.BLN(BLN14),.WL(WL168));
sram_cell_6t_5 inst_cell_168_15 (.BL(BL15),.BLN(BLN15),.WL(WL168));
sram_cell_6t_5 inst_cell_168_16 (.BL(BL16),.BLN(BLN16),.WL(WL168));
sram_cell_6t_5 inst_cell_168_17 (.BL(BL17),.BLN(BLN17),.WL(WL168));
sram_cell_6t_5 inst_cell_168_18 (.BL(BL18),.BLN(BLN18),.WL(WL168));
sram_cell_6t_5 inst_cell_168_19 (.BL(BL19),.BLN(BLN19),.WL(WL168));
sram_cell_6t_5 inst_cell_168_20 (.BL(BL20),.BLN(BLN20),.WL(WL168));
sram_cell_6t_5 inst_cell_168_21 (.BL(BL21),.BLN(BLN21),.WL(WL168));
sram_cell_6t_5 inst_cell_168_22 (.BL(BL22),.BLN(BLN22),.WL(WL168));
sram_cell_6t_5 inst_cell_168_23 (.BL(BL23),.BLN(BLN23),.WL(WL168));
sram_cell_6t_5 inst_cell_168_24 (.BL(BL24),.BLN(BLN24),.WL(WL168));
sram_cell_6t_5 inst_cell_168_25 (.BL(BL25),.BLN(BLN25),.WL(WL168));
sram_cell_6t_5 inst_cell_168_26 (.BL(BL26),.BLN(BLN26),.WL(WL168));
sram_cell_6t_5 inst_cell_168_27 (.BL(BL27),.BLN(BLN27),.WL(WL168));
sram_cell_6t_5 inst_cell_168_28 (.BL(BL28),.BLN(BLN28),.WL(WL168));
sram_cell_6t_5 inst_cell_168_29 (.BL(BL29),.BLN(BLN29),.WL(WL168));
sram_cell_6t_5 inst_cell_168_30 (.BL(BL30),.BLN(BLN30),.WL(WL168));
sram_cell_6t_5 inst_cell_168_31 (.BL(BL31),.BLN(BLN31),.WL(WL168));
sram_cell_6t_5 inst_cell_168_32 (.BL(BL32),.BLN(BLN32),.WL(WL168));
sram_cell_6t_5 inst_cell_168_33 (.BL(BL33),.BLN(BLN33),.WL(WL168));
sram_cell_6t_5 inst_cell_168_34 (.BL(BL34),.BLN(BLN34),.WL(WL168));
sram_cell_6t_5 inst_cell_168_35 (.BL(BL35),.BLN(BLN35),.WL(WL168));
sram_cell_6t_5 inst_cell_168_36 (.BL(BL36),.BLN(BLN36),.WL(WL168));
sram_cell_6t_5 inst_cell_168_37 (.BL(BL37),.BLN(BLN37),.WL(WL168));
sram_cell_6t_5 inst_cell_168_38 (.BL(BL38),.BLN(BLN38),.WL(WL168));
sram_cell_6t_5 inst_cell_168_39 (.BL(BL39),.BLN(BLN39),.WL(WL168));
sram_cell_6t_5 inst_cell_168_40 (.BL(BL40),.BLN(BLN40),.WL(WL168));
sram_cell_6t_5 inst_cell_168_41 (.BL(BL41),.BLN(BLN41),.WL(WL168));
sram_cell_6t_5 inst_cell_168_42 (.BL(BL42),.BLN(BLN42),.WL(WL168));
sram_cell_6t_5 inst_cell_168_43 (.BL(BL43),.BLN(BLN43),.WL(WL168));
sram_cell_6t_5 inst_cell_168_44 (.BL(BL44),.BLN(BLN44),.WL(WL168));
sram_cell_6t_5 inst_cell_168_45 (.BL(BL45),.BLN(BLN45),.WL(WL168));
sram_cell_6t_5 inst_cell_168_46 (.BL(BL46),.BLN(BLN46),.WL(WL168));
sram_cell_6t_5 inst_cell_168_47 (.BL(BL47),.BLN(BLN47),.WL(WL168));
sram_cell_6t_5 inst_cell_168_48 (.BL(BL48),.BLN(BLN48),.WL(WL168));
sram_cell_6t_5 inst_cell_168_49 (.BL(BL49),.BLN(BLN49),.WL(WL168));
sram_cell_6t_5 inst_cell_168_50 (.BL(BL50),.BLN(BLN50),.WL(WL168));
sram_cell_6t_5 inst_cell_168_51 (.BL(BL51),.BLN(BLN51),.WL(WL168));
sram_cell_6t_5 inst_cell_168_52 (.BL(BL52),.BLN(BLN52),.WL(WL168));
sram_cell_6t_5 inst_cell_168_53 (.BL(BL53),.BLN(BLN53),.WL(WL168));
sram_cell_6t_5 inst_cell_168_54 (.BL(BL54),.BLN(BLN54),.WL(WL168));
sram_cell_6t_5 inst_cell_168_55 (.BL(BL55),.BLN(BLN55),.WL(WL168));
sram_cell_6t_5 inst_cell_168_56 (.BL(BL56),.BLN(BLN56),.WL(WL168));
sram_cell_6t_5 inst_cell_168_57 (.BL(BL57),.BLN(BLN57),.WL(WL168));
sram_cell_6t_5 inst_cell_168_58 (.BL(BL58),.BLN(BLN58),.WL(WL168));
sram_cell_6t_5 inst_cell_168_59 (.BL(BL59),.BLN(BLN59),.WL(WL168));
sram_cell_6t_5 inst_cell_168_60 (.BL(BL60),.BLN(BLN60),.WL(WL168));
sram_cell_6t_5 inst_cell_168_61 (.BL(BL61),.BLN(BLN61),.WL(WL168));
sram_cell_6t_5 inst_cell_168_62 (.BL(BL62),.BLN(BLN62),.WL(WL168));
sram_cell_6t_5 inst_cell_168_63 (.BL(BL63),.BLN(BLN63),.WL(WL168));
sram_cell_6t_5 inst_cell_168_64 (.BL(BL64),.BLN(BLN64),.WL(WL168));
sram_cell_6t_5 inst_cell_168_65 (.BL(BL65),.BLN(BLN65),.WL(WL168));
sram_cell_6t_5 inst_cell_168_66 (.BL(BL66),.BLN(BLN66),.WL(WL168));
sram_cell_6t_5 inst_cell_168_67 (.BL(BL67),.BLN(BLN67),.WL(WL168));
sram_cell_6t_5 inst_cell_168_68 (.BL(BL68),.BLN(BLN68),.WL(WL168));
sram_cell_6t_5 inst_cell_168_69 (.BL(BL69),.BLN(BLN69),.WL(WL168));
sram_cell_6t_5 inst_cell_168_70 (.BL(BL70),.BLN(BLN70),.WL(WL168));
sram_cell_6t_5 inst_cell_168_71 (.BL(BL71),.BLN(BLN71),.WL(WL168));
sram_cell_6t_5 inst_cell_168_72 (.BL(BL72),.BLN(BLN72),.WL(WL168));
sram_cell_6t_5 inst_cell_168_73 (.BL(BL73),.BLN(BLN73),.WL(WL168));
sram_cell_6t_5 inst_cell_168_74 (.BL(BL74),.BLN(BLN74),.WL(WL168));
sram_cell_6t_5 inst_cell_168_75 (.BL(BL75),.BLN(BLN75),.WL(WL168));
sram_cell_6t_5 inst_cell_168_76 (.BL(BL76),.BLN(BLN76),.WL(WL168));
sram_cell_6t_5 inst_cell_168_77 (.BL(BL77),.BLN(BLN77),.WL(WL168));
sram_cell_6t_5 inst_cell_168_78 (.BL(BL78),.BLN(BLN78),.WL(WL168));
sram_cell_6t_5 inst_cell_168_79 (.BL(BL79),.BLN(BLN79),.WL(WL168));
sram_cell_6t_5 inst_cell_168_80 (.BL(BL80),.BLN(BLN80),.WL(WL168));
sram_cell_6t_5 inst_cell_168_81 (.BL(BL81),.BLN(BLN81),.WL(WL168));
sram_cell_6t_5 inst_cell_168_82 (.BL(BL82),.BLN(BLN82),.WL(WL168));
sram_cell_6t_5 inst_cell_168_83 (.BL(BL83),.BLN(BLN83),.WL(WL168));
sram_cell_6t_5 inst_cell_168_84 (.BL(BL84),.BLN(BLN84),.WL(WL168));
sram_cell_6t_5 inst_cell_168_85 (.BL(BL85),.BLN(BLN85),.WL(WL168));
sram_cell_6t_5 inst_cell_168_86 (.BL(BL86),.BLN(BLN86),.WL(WL168));
sram_cell_6t_5 inst_cell_168_87 (.BL(BL87),.BLN(BLN87),.WL(WL168));
sram_cell_6t_5 inst_cell_168_88 (.BL(BL88),.BLN(BLN88),.WL(WL168));
sram_cell_6t_5 inst_cell_168_89 (.BL(BL89),.BLN(BLN89),.WL(WL168));
sram_cell_6t_5 inst_cell_168_90 (.BL(BL90),.BLN(BLN90),.WL(WL168));
sram_cell_6t_5 inst_cell_168_91 (.BL(BL91),.BLN(BLN91),.WL(WL168));
sram_cell_6t_5 inst_cell_168_92 (.BL(BL92),.BLN(BLN92),.WL(WL168));
sram_cell_6t_5 inst_cell_168_93 (.BL(BL93),.BLN(BLN93),.WL(WL168));
sram_cell_6t_5 inst_cell_168_94 (.BL(BL94),.BLN(BLN94),.WL(WL168));
sram_cell_6t_5 inst_cell_168_95 (.BL(BL95),.BLN(BLN95),.WL(WL168));
sram_cell_6t_5 inst_cell_168_96 (.BL(BL96),.BLN(BLN96),.WL(WL168));
sram_cell_6t_5 inst_cell_168_97 (.BL(BL97),.BLN(BLN97),.WL(WL168));
sram_cell_6t_5 inst_cell_168_98 (.BL(BL98),.BLN(BLN98),.WL(WL168));
sram_cell_6t_5 inst_cell_168_99 (.BL(BL99),.BLN(BLN99),.WL(WL168));
sram_cell_6t_5 inst_cell_168_100 (.BL(BL100),.BLN(BLN100),.WL(WL168));
sram_cell_6t_5 inst_cell_168_101 (.BL(BL101),.BLN(BLN101),.WL(WL168));
sram_cell_6t_5 inst_cell_168_102 (.BL(BL102),.BLN(BLN102),.WL(WL168));
sram_cell_6t_5 inst_cell_168_103 (.BL(BL103),.BLN(BLN103),.WL(WL168));
sram_cell_6t_5 inst_cell_168_104 (.BL(BL104),.BLN(BLN104),.WL(WL168));
sram_cell_6t_5 inst_cell_168_105 (.BL(BL105),.BLN(BLN105),.WL(WL168));
sram_cell_6t_5 inst_cell_168_106 (.BL(BL106),.BLN(BLN106),.WL(WL168));
sram_cell_6t_5 inst_cell_168_107 (.BL(BL107),.BLN(BLN107),.WL(WL168));
sram_cell_6t_5 inst_cell_168_108 (.BL(BL108),.BLN(BLN108),.WL(WL168));
sram_cell_6t_5 inst_cell_168_109 (.BL(BL109),.BLN(BLN109),.WL(WL168));
sram_cell_6t_5 inst_cell_168_110 (.BL(BL110),.BLN(BLN110),.WL(WL168));
sram_cell_6t_5 inst_cell_168_111 (.BL(BL111),.BLN(BLN111),.WL(WL168));
sram_cell_6t_5 inst_cell_168_112 (.BL(BL112),.BLN(BLN112),.WL(WL168));
sram_cell_6t_5 inst_cell_168_113 (.BL(BL113),.BLN(BLN113),.WL(WL168));
sram_cell_6t_5 inst_cell_168_114 (.BL(BL114),.BLN(BLN114),.WL(WL168));
sram_cell_6t_5 inst_cell_168_115 (.BL(BL115),.BLN(BLN115),.WL(WL168));
sram_cell_6t_5 inst_cell_168_116 (.BL(BL116),.BLN(BLN116),.WL(WL168));
sram_cell_6t_5 inst_cell_168_117 (.BL(BL117),.BLN(BLN117),.WL(WL168));
sram_cell_6t_5 inst_cell_168_118 (.BL(BL118),.BLN(BLN118),.WL(WL168));
sram_cell_6t_5 inst_cell_168_119 (.BL(BL119),.BLN(BLN119),.WL(WL168));
sram_cell_6t_5 inst_cell_168_120 (.BL(BL120),.BLN(BLN120),.WL(WL168));
sram_cell_6t_5 inst_cell_168_121 (.BL(BL121),.BLN(BLN121),.WL(WL168));
sram_cell_6t_5 inst_cell_168_122 (.BL(BL122),.BLN(BLN122),.WL(WL168));
sram_cell_6t_5 inst_cell_168_123 (.BL(BL123),.BLN(BLN123),.WL(WL168));
sram_cell_6t_5 inst_cell_168_124 (.BL(BL124),.BLN(BLN124),.WL(WL168));
sram_cell_6t_5 inst_cell_168_125 (.BL(BL125),.BLN(BLN125),.WL(WL168));
sram_cell_6t_5 inst_cell_168_126 (.BL(BL126),.BLN(BLN126),.WL(WL168));
sram_cell_6t_5 inst_cell_168_127 (.BL(BL127),.BLN(BLN127),.WL(WL168));
sram_cell_6t_5 inst_cell_169_0 (.BL(BL0),.BLN(BLN0),.WL(WL169));
sram_cell_6t_5 inst_cell_169_1 (.BL(BL1),.BLN(BLN1),.WL(WL169));
sram_cell_6t_5 inst_cell_169_2 (.BL(BL2),.BLN(BLN2),.WL(WL169));
sram_cell_6t_5 inst_cell_169_3 (.BL(BL3),.BLN(BLN3),.WL(WL169));
sram_cell_6t_5 inst_cell_169_4 (.BL(BL4),.BLN(BLN4),.WL(WL169));
sram_cell_6t_5 inst_cell_169_5 (.BL(BL5),.BLN(BLN5),.WL(WL169));
sram_cell_6t_5 inst_cell_169_6 (.BL(BL6),.BLN(BLN6),.WL(WL169));
sram_cell_6t_5 inst_cell_169_7 (.BL(BL7),.BLN(BLN7),.WL(WL169));
sram_cell_6t_5 inst_cell_169_8 (.BL(BL8),.BLN(BLN8),.WL(WL169));
sram_cell_6t_5 inst_cell_169_9 (.BL(BL9),.BLN(BLN9),.WL(WL169));
sram_cell_6t_5 inst_cell_169_10 (.BL(BL10),.BLN(BLN10),.WL(WL169));
sram_cell_6t_5 inst_cell_169_11 (.BL(BL11),.BLN(BLN11),.WL(WL169));
sram_cell_6t_5 inst_cell_169_12 (.BL(BL12),.BLN(BLN12),.WL(WL169));
sram_cell_6t_5 inst_cell_169_13 (.BL(BL13),.BLN(BLN13),.WL(WL169));
sram_cell_6t_5 inst_cell_169_14 (.BL(BL14),.BLN(BLN14),.WL(WL169));
sram_cell_6t_5 inst_cell_169_15 (.BL(BL15),.BLN(BLN15),.WL(WL169));
sram_cell_6t_5 inst_cell_169_16 (.BL(BL16),.BLN(BLN16),.WL(WL169));
sram_cell_6t_5 inst_cell_169_17 (.BL(BL17),.BLN(BLN17),.WL(WL169));
sram_cell_6t_5 inst_cell_169_18 (.BL(BL18),.BLN(BLN18),.WL(WL169));
sram_cell_6t_5 inst_cell_169_19 (.BL(BL19),.BLN(BLN19),.WL(WL169));
sram_cell_6t_5 inst_cell_169_20 (.BL(BL20),.BLN(BLN20),.WL(WL169));
sram_cell_6t_5 inst_cell_169_21 (.BL(BL21),.BLN(BLN21),.WL(WL169));
sram_cell_6t_5 inst_cell_169_22 (.BL(BL22),.BLN(BLN22),.WL(WL169));
sram_cell_6t_5 inst_cell_169_23 (.BL(BL23),.BLN(BLN23),.WL(WL169));
sram_cell_6t_5 inst_cell_169_24 (.BL(BL24),.BLN(BLN24),.WL(WL169));
sram_cell_6t_5 inst_cell_169_25 (.BL(BL25),.BLN(BLN25),.WL(WL169));
sram_cell_6t_5 inst_cell_169_26 (.BL(BL26),.BLN(BLN26),.WL(WL169));
sram_cell_6t_5 inst_cell_169_27 (.BL(BL27),.BLN(BLN27),.WL(WL169));
sram_cell_6t_5 inst_cell_169_28 (.BL(BL28),.BLN(BLN28),.WL(WL169));
sram_cell_6t_5 inst_cell_169_29 (.BL(BL29),.BLN(BLN29),.WL(WL169));
sram_cell_6t_5 inst_cell_169_30 (.BL(BL30),.BLN(BLN30),.WL(WL169));
sram_cell_6t_5 inst_cell_169_31 (.BL(BL31),.BLN(BLN31),.WL(WL169));
sram_cell_6t_5 inst_cell_169_32 (.BL(BL32),.BLN(BLN32),.WL(WL169));
sram_cell_6t_5 inst_cell_169_33 (.BL(BL33),.BLN(BLN33),.WL(WL169));
sram_cell_6t_5 inst_cell_169_34 (.BL(BL34),.BLN(BLN34),.WL(WL169));
sram_cell_6t_5 inst_cell_169_35 (.BL(BL35),.BLN(BLN35),.WL(WL169));
sram_cell_6t_5 inst_cell_169_36 (.BL(BL36),.BLN(BLN36),.WL(WL169));
sram_cell_6t_5 inst_cell_169_37 (.BL(BL37),.BLN(BLN37),.WL(WL169));
sram_cell_6t_5 inst_cell_169_38 (.BL(BL38),.BLN(BLN38),.WL(WL169));
sram_cell_6t_5 inst_cell_169_39 (.BL(BL39),.BLN(BLN39),.WL(WL169));
sram_cell_6t_5 inst_cell_169_40 (.BL(BL40),.BLN(BLN40),.WL(WL169));
sram_cell_6t_5 inst_cell_169_41 (.BL(BL41),.BLN(BLN41),.WL(WL169));
sram_cell_6t_5 inst_cell_169_42 (.BL(BL42),.BLN(BLN42),.WL(WL169));
sram_cell_6t_5 inst_cell_169_43 (.BL(BL43),.BLN(BLN43),.WL(WL169));
sram_cell_6t_5 inst_cell_169_44 (.BL(BL44),.BLN(BLN44),.WL(WL169));
sram_cell_6t_5 inst_cell_169_45 (.BL(BL45),.BLN(BLN45),.WL(WL169));
sram_cell_6t_5 inst_cell_169_46 (.BL(BL46),.BLN(BLN46),.WL(WL169));
sram_cell_6t_5 inst_cell_169_47 (.BL(BL47),.BLN(BLN47),.WL(WL169));
sram_cell_6t_5 inst_cell_169_48 (.BL(BL48),.BLN(BLN48),.WL(WL169));
sram_cell_6t_5 inst_cell_169_49 (.BL(BL49),.BLN(BLN49),.WL(WL169));
sram_cell_6t_5 inst_cell_169_50 (.BL(BL50),.BLN(BLN50),.WL(WL169));
sram_cell_6t_5 inst_cell_169_51 (.BL(BL51),.BLN(BLN51),.WL(WL169));
sram_cell_6t_5 inst_cell_169_52 (.BL(BL52),.BLN(BLN52),.WL(WL169));
sram_cell_6t_5 inst_cell_169_53 (.BL(BL53),.BLN(BLN53),.WL(WL169));
sram_cell_6t_5 inst_cell_169_54 (.BL(BL54),.BLN(BLN54),.WL(WL169));
sram_cell_6t_5 inst_cell_169_55 (.BL(BL55),.BLN(BLN55),.WL(WL169));
sram_cell_6t_5 inst_cell_169_56 (.BL(BL56),.BLN(BLN56),.WL(WL169));
sram_cell_6t_5 inst_cell_169_57 (.BL(BL57),.BLN(BLN57),.WL(WL169));
sram_cell_6t_5 inst_cell_169_58 (.BL(BL58),.BLN(BLN58),.WL(WL169));
sram_cell_6t_5 inst_cell_169_59 (.BL(BL59),.BLN(BLN59),.WL(WL169));
sram_cell_6t_5 inst_cell_169_60 (.BL(BL60),.BLN(BLN60),.WL(WL169));
sram_cell_6t_5 inst_cell_169_61 (.BL(BL61),.BLN(BLN61),.WL(WL169));
sram_cell_6t_5 inst_cell_169_62 (.BL(BL62),.BLN(BLN62),.WL(WL169));
sram_cell_6t_5 inst_cell_169_63 (.BL(BL63),.BLN(BLN63),.WL(WL169));
sram_cell_6t_5 inst_cell_169_64 (.BL(BL64),.BLN(BLN64),.WL(WL169));
sram_cell_6t_5 inst_cell_169_65 (.BL(BL65),.BLN(BLN65),.WL(WL169));
sram_cell_6t_5 inst_cell_169_66 (.BL(BL66),.BLN(BLN66),.WL(WL169));
sram_cell_6t_5 inst_cell_169_67 (.BL(BL67),.BLN(BLN67),.WL(WL169));
sram_cell_6t_5 inst_cell_169_68 (.BL(BL68),.BLN(BLN68),.WL(WL169));
sram_cell_6t_5 inst_cell_169_69 (.BL(BL69),.BLN(BLN69),.WL(WL169));
sram_cell_6t_5 inst_cell_169_70 (.BL(BL70),.BLN(BLN70),.WL(WL169));
sram_cell_6t_5 inst_cell_169_71 (.BL(BL71),.BLN(BLN71),.WL(WL169));
sram_cell_6t_5 inst_cell_169_72 (.BL(BL72),.BLN(BLN72),.WL(WL169));
sram_cell_6t_5 inst_cell_169_73 (.BL(BL73),.BLN(BLN73),.WL(WL169));
sram_cell_6t_5 inst_cell_169_74 (.BL(BL74),.BLN(BLN74),.WL(WL169));
sram_cell_6t_5 inst_cell_169_75 (.BL(BL75),.BLN(BLN75),.WL(WL169));
sram_cell_6t_5 inst_cell_169_76 (.BL(BL76),.BLN(BLN76),.WL(WL169));
sram_cell_6t_5 inst_cell_169_77 (.BL(BL77),.BLN(BLN77),.WL(WL169));
sram_cell_6t_5 inst_cell_169_78 (.BL(BL78),.BLN(BLN78),.WL(WL169));
sram_cell_6t_5 inst_cell_169_79 (.BL(BL79),.BLN(BLN79),.WL(WL169));
sram_cell_6t_5 inst_cell_169_80 (.BL(BL80),.BLN(BLN80),.WL(WL169));
sram_cell_6t_5 inst_cell_169_81 (.BL(BL81),.BLN(BLN81),.WL(WL169));
sram_cell_6t_5 inst_cell_169_82 (.BL(BL82),.BLN(BLN82),.WL(WL169));
sram_cell_6t_5 inst_cell_169_83 (.BL(BL83),.BLN(BLN83),.WL(WL169));
sram_cell_6t_5 inst_cell_169_84 (.BL(BL84),.BLN(BLN84),.WL(WL169));
sram_cell_6t_5 inst_cell_169_85 (.BL(BL85),.BLN(BLN85),.WL(WL169));
sram_cell_6t_5 inst_cell_169_86 (.BL(BL86),.BLN(BLN86),.WL(WL169));
sram_cell_6t_5 inst_cell_169_87 (.BL(BL87),.BLN(BLN87),.WL(WL169));
sram_cell_6t_5 inst_cell_169_88 (.BL(BL88),.BLN(BLN88),.WL(WL169));
sram_cell_6t_5 inst_cell_169_89 (.BL(BL89),.BLN(BLN89),.WL(WL169));
sram_cell_6t_5 inst_cell_169_90 (.BL(BL90),.BLN(BLN90),.WL(WL169));
sram_cell_6t_5 inst_cell_169_91 (.BL(BL91),.BLN(BLN91),.WL(WL169));
sram_cell_6t_5 inst_cell_169_92 (.BL(BL92),.BLN(BLN92),.WL(WL169));
sram_cell_6t_5 inst_cell_169_93 (.BL(BL93),.BLN(BLN93),.WL(WL169));
sram_cell_6t_5 inst_cell_169_94 (.BL(BL94),.BLN(BLN94),.WL(WL169));
sram_cell_6t_5 inst_cell_169_95 (.BL(BL95),.BLN(BLN95),.WL(WL169));
sram_cell_6t_5 inst_cell_169_96 (.BL(BL96),.BLN(BLN96),.WL(WL169));
sram_cell_6t_5 inst_cell_169_97 (.BL(BL97),.BLN(BLN97),.WL(WL169));
sram_cell_6t_5 inst_cell_169_98 (.BL(BL98),.BLN(BLN98),.WL(WL169));
sram_cell_6t_5 inst_cell_169_99 (.BL(BL99),.BLN(BLN99),.WL(WL169));
sram_cell_6t_5 inst_cell_169_100 (.BL(BL100),.BLN(BLN100),.WL(WL169));
sram_cell_6t_5 inst_cell_169_101 (.BL(BL101),.BLN(BLN101),.WL(WL169));
sram_cell_6t_5 inst_cell_169_102 (.BL(BL102),.BLN(BLN102),.WL(WL169));
sram_cell_6t_5 inst_cell_169_103 (.BL(BL103),.BLN(BLN103),.WL(WL169));
sram_cell_6t_5 inst_cell_169_104 (.BL(BL104),.BLN(BLN104),.WL(WL169));
sram_cell_6t_5 inst_cell_169_105 (.BL(BL105),.BLN(BLN105),.WL(WL169));
sram_cell_6t_5 inst_cell_169_106 (.BL(BL106),.BLN(BLN106),.WL(WL169));
sram_cell_6t_5 inst_cell_169_107 (.BL(BL107),.BLN(BLN107),.WL(WL169));
sram_cell_6t_5 inst_cell_169_108 (.BL(BL108),.BLN(BLN108),.WL(WL169));
sram_cell_6t_5 inst_cell_169_109 (.BL(BL109),.BLN(BLN109),.WL(WL169));
sram_cell_6t_5 inst_cell_169_110 (.BL(BL110),.BLN(BLN110),.WL(WL169));
sram_cell_6t_5 inst_cell_169_111 (.BL(BL111),.BLN(BLN111),.WL(WL169));
sram_cell_6t_5 inst_cell_169_112 (.BL(BL112),.BLN(BLN112),.WL(WL169));
sram_cell_6t_5 inst_cell_169_113 (.BL(BL113),.BLN(BLN113),.WL(WL169));
sram_cell_6t_5 inst_cell_169_114 (.BL(BL114),.BLN(BLN114),.WL(WL169));
sram_cell_6t_5 inst_cell_169_115 (.BL(BL115),.BLN(BLN115),.WL(WL169));
sram_cell_6t_5 inst_cell_169_116 (.BL(BL116),.BLN(BLN116),.WL(WL169));
sram_cell_6t_5 inst_cell_169_117 (.BL(BL117),.BLN(BLN117),.WL(WL169));
sram_cell_6t_5 inst_cell_169_118 (.BL(BL118),.BLN(BLN118),.WL(WL169));
sram_cell_6t_5 inst_cell_169_119 (.BL(BL119),.BLN(BLN119),.WL(WL169));
sram_cell_6t_5 inst_cell_169_120 (.BL(BL120),.BLN(BLN120),.WL(WL169));
sram_cell_6t_5 inst_cell_169_121 (.BL(BL121),.BLN(BLN121),.WL(WL169));
sram_cell_6t_5 inst_cell_169_122 (.BL(BL122),.BLN(BLN122),.WL(WL169));
sram_cell_6t_5 inst_cell_169_123 (.BL(BL123),.BLN(BLN123),.WL(WL169));
sram_cell_6t_5 inst_cell_169_124 (.BL(BL124),.BLN(BLN124),.WL(WL169));
sram_cell_6t_5 inst_cell_169_125 (.BL(BL125),.BLN(BLN125),.WL(WL169));
sram_cell_6t_5 inst_cell_169_126 (.BL(BL126),.BLN(BLN126),.WL(WL169));
sram_cell_6t_5 inst_cell_169_127 (.BL(BL127),.BLN(BLN127),.WL(WL169));
sram_cell_6t_5 inst_cell_170_0 (.BL(BL0),.BLN(BLN0),.WL(WL170));
sram_cell_6t_5 inst_cell_170_1 (.BL(BL1),.BLN(BLN1),.WL(WL170));
sram_cell_6t_5 inst_cell_170_2 (.BL(BL2),.BLN(BLN2),.WL(WL170));
sram_cell_6t_5 inst_cell_170_3 (.BL(BL3),.BLN(BLN3),.WL(WL170));
sram_cell_6t_5 inst_cell_170_4 (.BL(BL4),.BLN(BLN4),.WL(WL170));
sram_cell_6t_5 inst_cell_170_5 (.BL(BL5),.BLN(BLN5),.WL(WL170));
sram_cell_6t_5 inst_cell_170_6 (.BL(BL6),.BLN(BLN6),.WL(WL170));
sram_cell_6t_5 inst_cell_170_7 (.BL(BL7),.BLN(BLN7),.WL(WL170));
sram_cell_6t_5 inst_cell_170_8 (.BL(BL8),.BLN(BLN8),.WL(WL170));
sram_cell_6t_5 inst_cell_170_9 (.BL(BL9),.BLN(BLN9),.WL(WL170));
sram_cell_6t_5 inst_cell_170_10 (.BL(BL10),.BLN(BLN10),.WL(WL170));
sram_cell_6t_5 inst_cell_170_11 (.BL(BL11),.BLN(BLN11),.WL(WL170));
sram_cell_6t_5 inst_cell_170_12 (.BL(BL12),.BLN(BLN12),.WL(WL170));
sram_cell_6t_5 inst_cell_170_13 (.BL(BL13),.BLN(BLN13),.WL(WL170));
sram_cell_6t_5 inst_cell_170_14 (.BL(BL14),.BLN(BLN14),.WL(WL170));
sram_cell_6t_5 inst_cell_170_15 (.BL(BL15),.BLN(BLN15),.WL(WL170));
sram_cell_6t_5 inst_cell_170_16 (.BL(BL16),.BLN(BLN16),.WL(WL170));
sram_cell_6t_5 inst_cell_170_17 (.BL(BL17),.BLN(BLN17),.WL(WL170));
sram_cell_6t_5 inst_cell_170_18 (.BL(BL18),.BLN(BLN18),.WL(WL170));
sram_cell_6t_5 inst_cell_170_19 (.BL(BL19),.BLN(BLN19),.WL(WL170));
sram_cell_6t_5 inst_cell_170_20 (.BL(BL20),.BLN(BLN20),.WL(WL170));
sram_cell_6t_5 inst_cell_170_21 (.BL(BL21),.BLN(BLN21),.WL(WL170));
sram_cell_6t_5 inst_cell_170_22 (.BL(BL22),.BLN(BLN22),.WL(WL170));
sram_cell_6t_5 inst_cell_170_23 (.BL(BL23),.BLN(BLN23),.WL(WL170));
sram_cell_6t_5 inst_cell_170_24 (.BL(BL24),.BLN(BLN24),.WL(WL170));
sram_cell_6t_5 inst_cell_170_25 (.BL(BL25),.BLN(BLN25),.WL(WL170));
sram_cell_6t_5 inst_cell_170_26 (.BL(BL26),.BLN(BLN26),.WL(WL170));
sram_cell_6t_5 inst_cell_170_27 (.BL(BL27),.BLN(BLN27),.WL(WL170));
sram_cell_6t_5 inst_cell_170_28 (.BL(BL28),.BLN(BLN28),.WL(WL170));
sram_cell_6t_5 inst_cell_170_29 (.BL(BL29),.BLN(BLN29),.WL(WL170));
sram_cell_6t_5 inst_cell_170_30 (.BL(BL30),.BLN(BLN30),.WL(WL170));
sram_cell_6t_5 inst_cell_170_31 (.BL(BL31),.BLN(BLN31),.WL(WL170));
sram_cell_6t_5 inst_cell_170_32 (.BL(BL32),.BLN(BLN32),.WL(WL170));
sram_cell_6t_5 inst_cell_170_33 (.BL(BL33),.BLN(BLN33),.WL(WL170));
sram_cell_6t_5 inst_cell_170_34 (.BL(BL34),.BLN(BLN34),.WL(WL170));
sram_cell_6t_5 inst_cell_170_35 (.BL(BL35),.BLN(BLN35),.WL(WL170));
sram_cell_6t_5 inst_cell_170_36 (.BL(BL36),.BLN(BLN36),.WL(WL170));
sram_cell_6t_5 inst_cell_170_37 (.BL(BL37),.BLN(BLN37),.WL(WL170));
sram_cell_6t_5 inst_cell_170_38 (.BL(BL38),.BLN(BLN38),.WL(WL170));
sram_cell_6t_5 inst_cell_170_39 (.BL(BL39),.BLN(BLN39),.WL(WL170));
sram_cell_6t_5 inst_cell_170_40 (.BL(BL40),.BLN(BLN40),.WL(WL170));
sram_cell_6t_5 inst_cell_170_41 (.BL(BL41),.BLN(BLN41),.WL(WL170));
sram_cell_6t_5 inst_cell_170_42 (.BL(BL42),.BLN(BLN42),.WL(WL170));
sram_cell_6t_5 inst_cell_170_43 (.BL(BL43),.BLN(BLN43),.WL(WL170));
sram_cell_6t_5 inst_cell_170_44 (.BL(BL44),.BLN(BLN44),.WL(WL170));
sram_cell_6t_5 inst_cell_170_45 (.BL(BL45),.BLN(BLN45),.WL(WL170));
sram_cell_6t_5 inst_cell_170_46 (.BL(BL46),.BLN(BLN46),.WL(WL170));
sram_cell_6t_5 inst_cell_170_47 (.BL(BL47),.BLN(BLN47),.WL(WL170));
sram_cell_6t_5 inst_cell_170_48 (.BL(BL48),.BLN(BLN48),.WL(WL170));
sram_cell_6t_5 inst_cell_170_49 (.BL(BL49),.BLN(BLN49),.WL(WL170));
sram_cell_6t_5 inst_cell_170_50 (.BL(BL50),.BLN(BLN50),.WL(WL170));
sram_cell_6t_5 inst_cell_170_51 (.BL(BL51),.BLN(BLN51),.WL(WL170));
sram_cell_6t_5 inst_cell_170_52 (.BL(BL52),.BLN(BLN52),.WL(WL170));
sram_cell_6t_5 inst_cell_170_53 (.BL(BL53),.BLN(BLN53),.WL(WL170));
sram_cell_6t_5 inst_cell_170_54 (.BL(BL54),.BLN(BLN54),.WL(WL170));
sram_cell_6t_5 inst_cell_170_55 (.BL(BL55),.BLN(BLN55),.WL(WL170));
sram_cell_6t_5 inst_cell_170_56 (.BL(BL56),.BLN(BLN56),.WL(WL170));
sram_cell_6t_5 inst_cell_170_57 (.BL(BL57),.BLN(BLN57),.WL(WL170));
sram_cell_6t_5 inst_cell_170_58 (.BL(BL58),.BLN(BLN58),.WL(WL170));
sram_cell_6t_5 inst_cell_170_59 (.BL(BL59),.BLN(BLN59),.WL(WL170));
sram_cell_6t_5 inst_cell_170_60 (.BL(BL60),.BLN(BLN60),.WL(WL170));
sram_cell_6t_5 inst_cell_170_61 (.BL(BL61),.BLN(BLN61),.WL(WL170));
sram_cell_6t_5 inst_cell_170_62 (.BL(BL62),.BLN(BLN62),.WL(WL170));
sram_cell_6t_5 inst_cell_170_63 (.BL(BL63),.BLN(BLN63),.WL(WL170));
sram_cell_6t_5 inst_cell_170_64 (.BL(BL64),.BLN(BLN64),.WL(WL170));
sram_cell_6t_5 inst_cell_170_65 (.BL(BL65),.BLN(BLN65),.WL(WL170));
sram_cell_6t_5 inst_cell_170_66 (.BL(BL66),.BLN(BLN66),.WL(WL170));
sram_cell_6t_5 inst_cell_170_67 (.BL(BL67),.BLN(BLN67),.WL(WL170));
sram_cell_6t_5 inst_cell_170_68 (.BL(BL68),.BLN(BLN68),.WL(WL170));
sram_cell_6t_5 inst_cell_170_69 (.BL(BL69),.BLN(BLN69),.WL(WL170));
sram_cell_6t_5 inst_cell_170_70 (.BL(BL70),.BLN(BLN70),.WL(WL170));
sram_cell_6t_5 inst_cell_170_71 (.BL(BL71),.BLN(BLN71),.WL(WL170));
sram_cell_6t_5 inst_cell_170_72 (.BL(BL72),.BLN(BLN72),.WL(WL170));
sram_cell_6t_5 inst_cell_170_73 (.BL(BL73),.BLN(BLN73),.WL(WL170));
sram_cell_6t_5 inst_cell_170_74 (.BL(BL74),.BLN(BLN74),.WL(WL170));
sram_cell_6t_5 inst_cell_170_75 (.BL(BL75),.BLN(BLN75),.WL(WL170));
sram_cell_6t_5 inst_cell_170_76 (.BL(BL76),.BLN(BLN76),.WL(WL170));
sram_cell_6t_5 inst_cell_170_77 (.BL(BL77),.BLN(BLN77),.WL(WL170));
sram_cell_6t_5 inst_cell_170_78 (.BL(BL78),.BLN(BLN78),.WL(WL170));
sram_cell_6t_5 inst_cell_170_79 (.BL(BL79),.BLN(BLN79),.WL(WL170));
sram_cell_6t_5 inst_cell_170_80 (.BL(BL80),.BLN(BLN80),.WL(WL170));
sram_cell_6t_5 inst_cell_170_81 (.BL(BL81),.BLN(BLN81),.WL(WL170));
sram_cell_6t_5 inst_cell_170_82 (.BL(BL82),.BLN(BLN82),.WL(WL170));
sram_cell_6t_5 inst_cell_170_83 (.BL(BL83),.BLN(BLN83),.WL(WL170));
sram_cell_6t_5 inst_cell_170_84 (.BL(BL84),.BLN(BLN84),.WL(WL170));
sram_cell_6t_5 inst_cell_170_85 (.BL(BL85),.BLN(BLN85),.WL(WL170));
sram_cell_6t_5 inst_cell_170_86 (.BL(BL86),.BLN(BLN86),.WL(WL170));
sram_cell_6t_5 inst_cell_170_87 (.BL(BL87),.BLN(BLN87),.WL(WL170));
sram_cell_6t_5 inst_cell_170_88 (.BL(BL88),.BLN(BLN88),.WL(WL170));
sram_cell_6t_5 inst_cell_170_89 (.BL(BL89),.BLN(BLN89),.WL(WL170));
sram_cell_6t_5 inst_cell_170_90 (.BL(BL90),.BLN(BLN90),.WL(WL170));
sram_cell_6t_5 inst_cell_170_91 (.BL(BL91),.BLN(BLN91),.WL(WL170));
sram_cell_6t_5 inst_cell_170_92 (.BL(BL92),.BLN(BLN92),.WL(WL170));
sram_cell_6t_5 inst_cell_170_93 (.BL(BL93),.BLN(BLN93),.WL(WL170));
sram_cell_6t_5 inst_cell_170_94 (.BL(BL94),.BLN(BLN94),.WL(WL170));
sram_cell_6t_5 inst_cell_170_95 (.BL(BL95),.BLN(BLN95),.WL(WL170));
sram_cell_6t_5 inst_cell_170_96 (.BL(BL96),.BLN(BLN96),.WL(WL170));
sram_cell_6t_5 inst_cell_170_97 (.BL(BL97),.BLN(BLN97),.WL(WL170));
sram_cell_6t_5 inst_cell_170_98 (.BL(BL98),.BLN(BLN98),.WL(WL170));
sram_cell_6t_5 inst_cell_170_99 (.BL(BL99),.BLN(BLN99),.WL(WL170));
sram_cell_6t_5 inst_cell_170_100 (.BL(BL100),.BLN(BLN100),.WL(WL170));
sram_cell_6t_5 inst_cell_170_101 (.BL(BL101),.BLN(BLN101),.WL(WL170));
sram_cell_6t_5 inst_cell_170_102 (.BL(BL102),.BLN(BLN102),.WL(WL170));
sram_cell_6t_5 inst_cell_170_103 (.BL(BL103),.BLN(BLN103),.WL(WL170));
sram_cell_6t_5 inst_cell_170_104 (.BL(BL104),.BLN(BLN104),.WL(WL170));
sram_cell_6t_5 inst_cell_170_105 (.BL(BL105),.BLN(BLN105),.WL(WL170));
sram_cell_6t_5 inst_cell_170_106 (.BL(BL106),.BLN(BLN106),.WL(WL170));
sram_cell_6t_5 inst_cell_170_107 (.BL(BL107),.BLN(BLN107),.WL(WL170));
sram_cell_6t_5 inst_cell_170_108 (.BL(BL108),.BLN(BLN108),.WL(WL170));
sram_cell_6t_5 inst_cell_170_109 (.BL(BL109),.BLN(BLN109),.WL(WL170));
sram_cell_6t_5 inst_cell_170_110 (.BL(BL110),.BLN(BLN110),.WL(WL170));
sram_cell_6t_5 inst_cell_170_111 (.BL(BL111),.BLN(BLN111),.WL(WL170));
sram_cell_6t_5 inst_cell_170_112 (.BL(BL112),.BLN(BLN112),.WL(WL170));
sram_cell_6t_5 inst_cell_170_113 (.BL(BL113),.BLN(BLN113),.WL(WL170));
sram_cell_6t_5 inst_cell_170_114 (.BL(BL114),.BLN(BLN114),.WL(WL170));
sram_cell_6t_5 inst_cell_170_115 (.BL(BL115),.BLN(BLN115),.WL(WL170));
sram_cell_6t_5 inst_cell_170_116 (.BL(BL116),.BLN(BLN116),.WL(WL170));
sram_cell_6t_5 inst_cell_170_117 (.BL(BL117),.BLN(BLN117),.WL(WL170));
sram_cell_6t_5 inst_cell_170_118 (.BL(BL118),.BLN(BLN118),.WL(WL170));
sram_cell_6t_5 inst_cell_170_119 (.BL(BL119),.BLN(BLN119),.WL(WL170));
sram_cell_6t_5 inst_cell_170_120 (.BL(BL120),.BLN(BLN120),.WL(WL170));
sram_cell_6t_5 inst_cell_170_121 (.BL(BL121),.BLN(BLN121),.WL(WL170));
sram_cell_6t_5 inst_cell_170_122 (.BL(BL122),.BLN(BLN122),.WL(WL170));
sram_cell_6t_5 inst_cell_170_123 (.BL(BL123),.BLN(BLN123),.WL(WL170));
sram_cell_6t_5 inst_cell_170_124 (.BL(BL124),.BLN(BLN124),.WL(WL170));
sram_cell_6t_5 inst_cell_170_125 (.BL(BL125),.BLN(BLN125),.WL(WL170));
sram_cell_6t_5 inst_cell_170_126 (.BL(BL126),.BLN(BLN126),.WL(WL170));
sram_cell_6t_5 inst_cell_170_127 (.BL(BL127),.BLN(BLN127),.WL(WL170));
sram_cell_6t_5 inst_cell_171_0 (.BL(BL0),.BLN(BLN0),.WL(WL171));
sram_cell_6t_5 inst_cell_171_1 (.BL(BL1),.BLN(BLN1),.WL(WL171));
sram_cell_6t_5 inst_cell_171_2 (.BL(BL2),.BLN(BLN2),.WL(WL171));
sram_cell_6t_5 inst_cell_171_3 (.BL(BL3),.BLN(BLN3),.WL(WL171));
sram_cell_6t_5 inst_cell_171_4 (.BL(BL4),.BLN(BLN4),.WL(WL171));
sram_cell_6t_5 inst_cell_171_5 (.BL(BL5),.BLN(BLN5),.WL(WL171));
sram_cell_6t_5 inst_cell_171_6 (.BL(BL6),.BLN(BLN6),.WL(WL171));
sram_cell_6t_5 inst_cell_171_7 (.BL(BL7),.BLN(BLN7),.WL(WL171));
sram_cell_6t_5 inst_cell_171_8 (.BL(BL8),.BLN(BLN8),.WL(WL171));
sram_cell_6t_5 inst_cell_171_9 (.BL(BL9),.BLN(BLN9),.WL(WL171));
sram_cell_6t_5 inst_cell_171_10 (.BL(BL10),.BLN(BLN10),.WL(WL171));
sram_cell_6t_5 inst_cell_171_11 (.BL(BL11),.BLN(BLN11),.WL(WL171));
sram_cell_6t_5 inst_cell_171_12 (.BL(BL12),.BLN(BLN12),.WL(WL171));
sram_cell_6t_5 inst_cell_171_13 (.BL(BL13),.BLN(BLN13),.WL(WL171));
sram_cell_6t_5 inst_cell_171_14 (.BL(BL14),.BLN(BLN14),.WL(WL171));
sram_cell_6t_5 inst_cell_171_15 (.BL(BL15),.BLN(BLN15),.WL(WL171));
sram_cell_6t_5 inst_cell_171_16 (.BL(BL16),.BLN(BLN16),.WL(WL171));
sram_cell_6t_5 inst_cell_171_17 (.BL(BL17),.BLN(BLN17),.WL(WL171));
sram_cell_6t_5 inst_cell_171_18 (.BL(BL18),.BLN(BLN18),.WL(WL171));
sram_cell_6t_5 inst_cell_171_19 (.BL(BL19),.BLN(BLN19),.WL(WL171));
sram_cell_6t_5 inst_cell_171_20 (.BL(BL20),.BLN(BLN20),.WL(WL171));
sram_cell_6t_5 inst_cell_171_21 (.BL(BL21),.BLN(BLN21),.WL(WL171));
sram_cell_6t_5 inst_cell_171_22 (.BL(BL22),.BLN(BLN22),.WL(WL171));
sram_cell_6t_5 inst_cell_171_23 (.BL(BL23),.BLN(BLN23),.WL(WL171));
sram_cell_6t_5 inst_cell_171_24 (.BL(BL24),.BLN(BLN24),.WL(WL171));
sram_cell_6t_5 inst_cell_171_25 (.BL(BL25),.BLN(BLN25),.WL(WL171));
sram_cell_6t_5 inst_cell_171_26 (.BL(BL26),.BLN(BLN26),.WL(WL171));
sram_cell_6t_5 inst_cell_171_27 (.BL(BL27),.BLN(BLN27),.WL(WL171));
sram_cell_6t_5 inst_cell_171_28 (.BL(BL28),.BLN(BLN28),.WL(WL171));
sram_cell_6t_5 inst_cell_171_29 (.BL(BL29),.BLN(BLN29),.WL(WL171));
sram_cell_6t_5 inst_cell_171_30 (.BL(BL30),.BLN(BLN30),.WL(WL171));
sram_cell_6t_5 inst_cell_171_31 (.BL(BL31),.BLN(BLN31),.WL(WL171));
sram_cell_6t_5 inst_cell_171_32 (.BL(BL32),.BLN(BLN32),.WL(WL171));
sram_cell_6t_5 inst_cell_171_33 (.BL(BL33),.BLN(BLN33),.WL(WL171));
sram_cell_6t_5 inst_cell_171_34 (.BL(BL34),.BLN(BLN34),.WL(WL171));
sram_cell_6t_5 inst_cell_171_35 (.BL(BL35),.BLN(BLN35),.WL(WL171));
sram_cell_6t_5 inst_cell_171_36 (.BL(BL36),.BLN(BLN36),.WL(WL171));
sram_cell_6t_5 inst_cell_171_37 (.BL(BL37),.BLN(BLN37),.WL(WL171));
sram_cell_6t_5 inst_cell_171_38 (.BL(BL38),.BLN(BLN38),.WL(WL171));
sram_cell_6t_5 inst_cell_171_39 (.BL(BL39),.BLN(BLN39),.WL(WL171));
sram_cell_6t_5 inst_cell_171_40 (.BL(BL40),.BLN(BLN40),.WL(WL171));
sram_cell_6t_5 inst_cell_171_41 (.BL(BL41),.BLN(BLN41),.WL(WL171));
sram_cell_6t_5 inst_cell_171_42 (.BL(BL42),.BLN(BLN42),.WL(WL171));
sram_cell_6t_5 inst_cell_171_43 (.BL(BL43),.BLN(BLN43),.WL(WL171));
sram_cell_6t_5 inst_cell_171_44 (.BL(BL44),.BLN(BLN44),.WL(WL171));
sram_cell_6t_5 inst_cell_171_45 (.BL(BL45),.BLN(BLN45),.WL(WL171));
sram_cell_6t_5 inst_cell_171_46 (.BL(BL46),.BLN(BLN46),.WL(WL171));
sram_cell_6t_5 inst_cell_171_47 (.BL(BL47),.BLN(BLN47),.WL(WL171));
sram_cell_6t_5 inst_cell_171_48 (.BL(BL48),.BLN(BLN48),.WL(WL171));
sram_cell_6t_5 inst_cell_171_49 (.BL(BL49),.BLN(BLN49),.WL(WL171));
sram_cell_6t_5 inst_cell_171_50 (.BL(BL50),.BLN(BLN50),.WL(WL171));
sram_cell_6t_5 inst_cell_171_51 (.BL(BL51),.BLN(BLN51),.WL(WL171));
sram_cell_6t_5 inst_cell_171_52 (.BL(BL52),.BLN(BLN52),.WL(WL171));
sram_cell_6t_5 inst_cell_171_53 (.BL(BL53),.BLN(BLN53),.WL(WL171));
sram_cell_6t_5 inst_cell_171_54 (.BL(BL54),.BLN(BLN54),.WL(WL171));
sram_cell_6t_5 inst_cell_171_55 (.BL(BL55),.BLN(BLN55),.WL(WL171));
sram_cell_6t_5 inst_cell_171_56 (.BL(BL56),.BLN(BLN56),.WL(WL171));
sram_cell_6t_5 inst_cell_171_57 (.BL(BL57),.BLN(BLN57),.WL(WL171));
sram_cell_6t_5 inst_cell_171_58 (.BL(BL58),.BLN(BLN58),.WL(WL171));
sram_cell_6t_5 inst_cell_171_59 (.BL(BL59),.BLN(BLN59),.WL(WL171));
sram_cell_6t_5 inst_cell_171_60 (.BL(BL60),.BLN(BLN60),.WL(WL171));
sram_cell_6t_5 inst_cell_171_61 (.BL(BL61),.BLN(BLN61),.WL(WL171));
sram_cell_6t_5 inst_cell_171_62 (.BL(BL62),.BLN(BLN62),.WL(WL171));
sram_cell_6t_5 inst_cell_171_63 (.BL(BL63),.BLN(BLN63),.WL(WL171));
sram_cell_6t_5 inst_cell_171_64 (.BL(BL64),.BLN(BLN64),.WL(WL171));
sram_cell_6t_5 inst_cell_171_65 (.BL(BL65),.BLN(BLN65),.WL(WL171));
sram_cell_6t_5 inst_cell_171_66 (.BL(BL66),.BLN(BLN66),.WL(WL171));
sram_cell_6t_5 inst_cell_171_67 (.BL(BL67),.BLN(BLN67),.WL(WL171));
sram_cell_6t_5 inst_cell_171_68 (.BL(BL68),.BLN(BLN68),.WL(WL171));
sram_cell_6t_5 inst_cell_171_69 (.BL(BL69),.BLN(BLN69),.WL(WL171));
sram_cell_6t_5 inst_cell_171_70 (.BL(BL70),.BLN(BLN70),.WL(WL171));
sram_cell_6t_5 inst_cell_171_71 (.BL(BL71),.BLN(BLN71),.WL(WL171));
sram_cell_6t_5 inst_cell_171_72 (.BL(BL72),.BLN(BLN72),.WL(WL171));
sram_cell_6t_5 inst_cell_171_73 (.BL(BL73),.BLN(BLN73),.WL(WL171));
sram_cell_6t_5 inst_cell_171_74 (.BL(BL74),.BLN(BLN74),.WL(WL171));
sram_cell_6t_5 inst_cell_171_75 (.BL(BL75),.BLN(BLN75),.WL(WL171));
sram_cell_6t_5 inst_cell_171_76 (.BL(BL76),.BLN(BLN76),.WL(WL171));
sram_cell_6t_5 inst_cell_171_77 (.BL(BL77),.BLN(BLN77),.WL(WL171));
sram_cell_6t_5 inst_cell_171_78 (.BL(BL78),.BLN(BLN78),.WL(WL171));
sram_cell_6t_5 inst_cell_171_79 (.BL(BL79),.BLN(BLN79),.WL(WL171));
sram_cell_6t_5 inst_cell_171_80 (.BL(BL80),.BLN(BLN80),.WL(WL171));
sram_cell_6t_5 inst_cell_171_81 (.BL(BL81),.BLN(BLN81),.WL(WL171));
sram_cell_6t_5 inst_cell_171_82 (.BL(BL82),.BLN(BLN82),.WL(WL171));
sram_cell_6t_5 inst_cell_171_83 (.BL(BL83),.BLN(BLN83),.WL(WL171));
sram_cell_6t_5 inst_cell_171_84 (.BL(BL84),.BLN(BLN84),.WL(WL171));
sram_cell_6t_5 inst_cell_171_85 (.BL(BL85),.BLN(BLN85),.WL(WL171));
sram_cell_6t_5 inst_cell_171_86 (.BL(BL86),.BLN(BLN86),.WL(WL171));
sram_cell_6t_5 inst_cell_171_87 (.BL(BL87),.BLN(BLN87),.WL(WL171));
sram_cell_6t_5 inst_cell_171_88 (.BL(BL88),.BLN(BLN88),.WL(WL171));
sram_cell_6t_5 inst_cell_171_89 (.BL(BL89),.BLN(BLN89),.WL(WL171));
sram_cell_6t_5 inst_cell_171_90 (.BL(BL90),.BLN(BLN90),.WL(WL171));
sram_cell_6t_5 inst_cell_171_91 (.BL(BL91),.BLN(BLN91),.WL(WL171));
sram_cell_6t_5 inst_cell_171_92 (.BL(BL92),.BLN(BLN92),.WL(WL171));
sram_cell_6t_5 inst_cell_171_93 (.BL(BL93),.BLN(BLN93),.WL(WL171));
sram_cell_6t_5 inst_cell_171_94 (.BL(BL94),.BLN(BLN94),.WL(WL171));
sram_cell_6t_5 inst_cell_171_95 (.BL(BL95),.BLN(BLN95),.WL(WL171));
sram_cell_6t_5 inst_cell_171_96 (.BL(BL96),.BLN(BLN96),.WL(WL171));
sram_cell_6t_5 inst_cell_171_97 (.BL(BL97),.BLN(BLN97),.WL(WL171));
sram_cell_6t_5 inst_cell_171_98 (.BL(BL98),.BLN(BLN98),.WL(WL171));
sram_cell_6t_5 inst_cell_171_99 (.BL(BL99),.BLN(BLN99),.WL(WL171));
sram_cell_6t_5 inst_cell_171_100 (.BL(BL100),.BLN(BLN100),.WL(WL171));
sram_cell_6t_5 inst_cell_171_101 (.BL(BL101),.BLN(BLN101),.WL(WL171));
sram_cell_6t_5 inst_cell_171_102 (.BL(BL102),.BLN(BLN102),.WL(WL171));
sram_cell_6t_5 inst_cell_171_103 (.BL(BL103),.BLN(BLN103),.WL(WL171));
sram_cell_6t_5 inst_cell_171_104 (.BL(BL104),.BLN(BLN104),.WL(WL171));
sram_cell_6t_5 inst_cell_171_105 (.BL(BL105),.BLN(BLN105),.WL(WL171));
sram_cell_6t_5 inst_cell_171_106 (.BL(BL106),.BLN(BLN106),.WL(WL171));
sram_cell_6t_5 inst_cell_171_107 (.BL(BL107),.BLN(BLN107),.WL(WL171));
sram_cell_6t_5 inst_cell_171_108 (.BL(BL108),.BLN(BLN108),.WL(WL171));
sram_cell_6t_5 inst_cell_171_109 (.BL(BL109),.BLN(BLN109),.WL(WL171));
sram_cell_6t_5 inst_cell_171_110 (.BL(BL110),.BLN(BLN110),.WL(WL171));
sram_cell_6t_5 inst_cell_171_111 (.BL(BL111),.BLN(BLN111),.WL(WL171));
sram_cell_6t_5 inst_cell_171_112 (.BL(BL112),.BLN(BLN112),.WL(WL171));
sram_cell_6t_5 inst_cell_171_113 (.BL(BL113),.BLN(BLN113),.WL(WL171));
sram_cell_6t_5 inst_cell_171_114 (.BL(BL114),.BLN(BLN114),.WL(WL171));
sram_cell_6t_5 inst_cell_171_115 (.BL(BL115),.BLN(BLN115),.WL(WL171));
sram_cell_6t_5 inst_cell_171_116 (.BL(BL116),.BLN(BLN116),.WL(WL171));
sram_cell_6t_5 inst_cell_171_117 (.BL(BL117),.BLN(BLN117),.WL(WL171));
sram_cell_6t_5 inst_cell_171_118 (.BL(BL118),.BLN(BLN118),.WL(WL171));
sram_cell_6t_5 inst_cell_171_119 (.BL(BL119),.BLN(BLN119),.WL(WL171));
sram_cell_6t_5 inst_cell_171_120 (.BL(BL120),.BLN(BLN120),.WL(WL171));
sram_cell_6t_5 inst_cell_171_121 (.BL(BL121),.BLN(BLN121),.WL(WL171));
sram_cell_6t_5 inst_cell_171_122 (.BL(BL122),.BLN(BLN122),.WL(WL171));
sram_cell_6t_5 inst_cell_171_123 (.BL(BL123),.BLN(BLN123),.WL(WL171));
sram_cell_6t_5 inst_cell_171_124 (.BL(BL124),.BLN(BLN124),.WL(WL171));
sram_cell_6t_5 inst_cell_171_125 (.BL(BL125),.BLN(BLN125),.WL(WL171));
sram_cell_6t_5 inst_cell_171_126 (.BL(BL126),.BLN(BLN126),.WL(WL171));
sram_cell_6t_5 inst_cell_171_127 (.BL(BL127),.BLN(BLN127),.WL(WL171));
sram_cell_6t_5 inst_cell_172_0 (.BL(BL0),.BLN(BLN0),.WL(WL172));
sram_cell_6t_5 inst_cell_172_1 (.BL(BL1),.BLN(BLN1),.WL(WL172));
sram_cell_6t_5 inst_cell_172_2 (.BL(BL2),.BLN(BLN2),.WL(WL172));
sram_cell_6t_5 inst_cell_172_3 (.BL(BL3),.BLN(BLN3),.WL(WL172));
sram_cell_6t_5 inst_cell_172_4 (.BL(BL4),.BLN(BLN4),.WL(WL172));
sram_cell_6t_5 inst_cell_172_5 (.BL(BL5),.BLN(BLN5),.WL(WL172));
sram_cell_6t_5 inst_cell_172_6 (.BL(BL6),.BLN(BLN6),.WL(WL172));
sram_cell_6t_5 inst_cell_172_7 (.BL(BL7),.BLN(BLN7),.WL(WL172));
sram_cell_6t_5 inst_cell_172_8 (.BL(BL8),.BLN(BLN8),.WL(WL172));
sram_cell_6t_5 inst_cell_172_9 (.BL(BL9),.BLN(BLN9),.WL(WL172));
sram_cell_6t_5 inst_cell_172_10 (.BL(BL10),.BLN(BLN10),.WL(WL172));
sram_cell_6t_5 inst_cell_172_11 (.BL(BL11),.BLN(BLN11),.WL(WL172));
sram_cell_6t_5 inst_cell_172_12 (.BL(BL12),.BLN(BLN12),.WL(WL172));
sram_cell_6t_5 inst_cell_172_13 (.BL(BL13),.BLN(BLN13),.WL(WL172));
sram_cell_6t_5 inst_cell_172_14 (.BL(BL14),.BLN(BLN14),.WL(WL172));
sram_cell_6t_5 inst_cell_172_15 (.BL(BL15),.BLN(BLN15),.WL(WL172));
sram_cell_6t_5 inst_cell_172_16 (.BL(BL16),.BLN(BLN16),.WL(WL172));
sram_cell_6t_5 inst_cell_172_17 (.BL(BL17),.BLN(BLN17),.WL(WL172));
sram_cell_6t_5 inst_cell_172_18 (.BL(BL18),.BLN(BLN18),.WL(WL172));
sram_cell_6t_5 inst_cell_172_19 (.BL(BL19),.BLN(BLN19),.WL(WL172));
sram_cell_6t_5 inst_cell_172_20 (.BL(BL20),.BLN(BLN20),.WL(WL172));
sram_cell_6t_5 inst_cell_172_21 (.BL(BL21),.BLN(BLN21),.WL(WL172));
sram_cell_6t_5 inst_cell_172_22 (.BL(BL22),.BLN(BLN22),.WL(WL172));
sram_cell_6t_5 inst_cell_172_23 (.BL(BL23),.BLN(BLN23),.WL(WL172));
sram_cell_6t_5 inst_cell_172_24 (.BL(BL24),.BLN(BLN24),.WL(WL172));
sram_cell_6t_5 inst_cell_172_25 (.BL(BL25),.BLN(BLN25),.WL(WL172));
sram_cell_6t_5 inst_cell_172_26 (.BL(BL26),.BLN(BLN26),.WL(WL172));
sram_cell_6t_5 inst_cell_172_27 (.BL(BL27),.BLN(BLN27),.WL(WL172));
sram_cell_6t_5 inst_cell_172_28 (.BL(BL28),.BLN(BLN28),.WL(WL172));
sram_cell_6t_5 inst_cell_172_29 (.BL(BL29),.BLN(BLN29),.WL(WL172));
sram_cell_6t_5 inst_cell_172_30 (.BL(BL30),.BLN(BLN30),.WL(WL172));
sram_cell_6t_5 inst_cell_172_31 (.BL(BL31),.BLN(BLN31),.WL(WL172));
sram_cell_6t_5 inst_cell_172_32 (.BL(BL32),.BLN(BLN32),.WL(WL172));
sram_cell_6t_5 inst_cell_172_33 (.BL(BL33),.BLN(BLN33),.WL(WL172));
sram_cell_6t_5 inst_cell_172_34 (.BL(BL34),.BLN(BLN34),.WL(WL172));
sram_cell_6t_5 inst_cell_172_35 (.BL(BL35),.BLN(BLN35),.WL(WL172));
sram_cell_6t_5 inst_cell_172_36 (.BL(BL36),.BLN(BLN36),.WL(WL172));
sram_cell_6t_5 inst_cell_172_37 (.BL(BL37),.BLN(BLN37),.WL(WL172));
sram_cell_6t_5 inst_cell_172_38 (.BL(BL38),.BLN(BLN38),.WL(WL172));
sram_cell_6t_5 inst_cell_172_39 (.BL(BL39),.BLN(BLN39),.WL(WL172));
sram_cell_6t_5 inst_cell_172_40 (.BL(BL40),.BLN(BLN40),.WL(WL172));
sram_cell_6t_5 inst_cell_172_41 (.BL(BL41),.BLN(BLN41),.WL(WL172));
sram_cell_6t_5 inst_cell_172_42 (.BL(BL42),.BLN(BLN42),.WL(WL172));
sram_cell_6t_5 inst_cell_172_43 (.BL(BL43),.BLN(BLN43),.WL(WL172));
sram_cell_6t_5 inst_cell_172_44 (.BL(BL44),.BLN(BLN44),.WL(WL172));
sram_cell_6t_5 inst_cell_172_45 (.BL(BL45),.BLN(BLN45),.WL(WL172));
sram_cell_6t_5 inst_cell_172_46 (.BL(BL46),.BLN(BLN46),.WL(WL172));
sram_cell_6t_5 inst_cell_172_47 (.BL(BL47),.BLN(BLN47),.WL(WL172));
sram_cell_6t_5 inst_cell_172_48 (.BL(BL48),.BLN(BLN48),.WL(WL172));
sram_cell_6t_5 inst_cell_172_49 (.BL(BL49),.BLN(BLN49),.WL(WL172));
sram_cell_6t_5 inst_cell_172_50 (.BL(BL50),.BLN(BLN50),.WL(WL172));
sram_cell_6t_5 inst_cell_172_51 (.BL(BL51),.BLN(BLN51),.WL(WL172));
sram_cell_6t_5 inst_cell_172_52 (.BL(BL52),.BLN(BLN52),.WL(WL172));
sram_cell_6t_5 inst_cell_172_53 (.BL(BL53),.BLN(BLN53),.WL(WL172));
sram_cell_6t_5 inst_cell_172_54 (.BL(BL54),.BLN(BLN54),.WL(WL172));
sram_cell_6t_5 inst_cell_172_55 (.BL(BL55),.BLN(BLN55),.WL(WL172));
sram_cell_6t_5 inst_cell_172_56 (.BL(BL56),.BLN(BLN56),.WL(WL172));
sram_cell_6t_5 inst_cell_172_57 (.BL(BL57),.BLN(BLN57),.WL(WL172));
sram_cell_6t_5 inst_cell_172_58 (.BL(BL58),.BLN(BLN58),.WL(WL172));
sram_cell_6t_5 inst_cell_172_59 (.BL(BL59),.BLN(BLN59),.WL(WL172));
sram_cell_6t_5 inst_cell_172_60 (.BL(BL60),.BLN(BLN60),.WL(WL172));
sram_cell_6t_5 inst_cell_172_61 (.BL(BL61),.BLN(BLN61),.WL(WL172));
sram_cell_6t_5 inst_cell_172_62 (.BL(BL62),.BLN(BLN62),.WL(WL172));
sram_cell_6t_5 inst_cell_172_63 (.BL(BL63),.BLN(BLN63),.WL(WL172));
sram_cell_6t_5 inst_cell_172_64 (.BL(BL64),.BLN(BLN64),.WL(WL172));
sram_cell_6t_5 inst_cell_172_65 (.BL(BL65),.BLN(BLN65),.WL(WL172));
sram_cell_6t_5 inst_cell_172_66 (.BL(BL66),.BLN(BLN66),.WL(WL172));
sram_cell_6t_5 inst_cell_172_67 (.BL(BL67),.BLN(BLN67),.WL(WL172));
sram_cell_6t_5 inst_cell_172_68 (.BL(BL68),.BLN(BLN68),.WL(WL172));
sram_cell_6t_5 inst_cell_172_69 (.BL(BL69),.BLN(BLN69),.WL(WL172));
sram_cell_6t_5 inst_cell_172_70 (.BL(BL70),.BLN(BLN70),.WL(WL172));
sram_cell_6t_5 inst_cell_172_71 (.BL(BL71),.BLN(BLN71),.WL(WL172));
sram_cell_6t_5 inst_cell_172_72 (.BL(BL72),.BLN(BLN72),.WL(WL172));
sram_cell_6t_5 inst_cell_172_73 (.BL(BL73),.BLN(BLN73),.WL(WL172));
sram_cell_6t_5 inst_cell_172_74 (.BL(BL74),.BLN(BLN74),.WL(WL172));
sram_cell_6t_5 inst_cell_172_75 (.BL(BL75),.BLN(BLN75),.WL(WL172));
sram_cell_6t_5 inst_cell_172_76 (.BL(BL76),.BLN(BLN76),.WL(WL172));
sram_cell_6t_5 inst_cell_172_77 (.BL(BL77),.BLN(BLN77),.WL(WL172));
sram_cell_6t_5 inst_cell_172_78 (.BL(BL78),.BLN(BLN78),.WL(WL172));
sram_cell_6t_5 inst_cell_172_79 (.BL(BL79),.BLN(BLN79),.WL(WL172));
sram_cell_6t_5 inst_cell_172_80 (.BL(BL80),.BLN(BLN80),.WL(WL172));
sram_cell_6t_5 inst_cell_172_81 (.BL(BL81),.BLN(BLN81),.WL(WL172));
sram_cell_6t_5 inst_cell_172_82 (.BL(BL82),.BLN(BLN82),.WL(WL172));
sram_cell_6t_5 inst_cell_172_83 (.BL(BL83),.BLN(BLN83),.WL(WL172));
sram_cell_6t_5 inst_cell_172_84 (.BL(BL84),.BLN(BLN84),.WL(WL172));
sram_cell_6t_5 inst_cell_172_85 (.BL(BL85),.BLN(BLN85),.WL(WL172));
sram_cell_6t_5 inst_cell_172_86 (.BL(BL86),.BLN(BLN86),.WL(WL172));
sram_cell_6t_5 inst_cell_172_87 (.BL(BL87),.BLN(BLN87),.WL(WL172));
sram_cell_6t_5 inst_cell_172_88 (.BL(BL88),.BLN(BLN88),.WL(WL172));
sram_cell_6t_5 inst_cell_172_89 (.BL(BL89),.BLN(BLN89),.WL(WL172));
sram_cell_6t_5 inst_cell_172_90 (.BL(BL90),.BLN(BLN90),.WL(WL172));
sram_cell_6t_5 inst_cell_172_91 (.BL(BL91),.BLN(BLN91),.WL(WL172));
sram_cell_6t_5 inst_cell_172_92 (.BL(BL92),.BLN(BLN92),.WL(WL172));
sram_cell_6t_5 inst_cell_172_93 (.BL(BL93),.BLN(BLN93),.WL(WL172));
sram_cell_6t_5 inst_cell_172_94 (.BL(BL94),.BLN(BLN94),.WL(WL172));
sram_cell_6t_5 inst_cell_172_95 (.BL(BL95),.BLN(BLN95),.WL(WL172));
sram_cell_6t_5 inst_cell_172_96 (.BL(BL96),.BLN(BLN96),.WL(WL172));
sram_cell_6t_5 inst_cell_172_97 (.BL(BL97),.BLN(BLN97),.WL(WL172));
sram_cell_6t_5 inst_cell_172_98 (.BL(BL98),.BLN(BLN98),.WL(WL172));
sram_cell_6t_5 inst_cell_172_99 (.BL(BL99),.BLN(BLN99),.WL(WL172));
sram_cell_6t_5 inst_cell_172_100 (.BL(BL100),.BLN(BLN100),.WL(WL172));
sram_cell_6t_5 inst_cell_172_101 (.BL(BL101),.BLN(BLN101),.WL(WL172));
sram_cell_6t_5 inst_cell_172_102 (.BL(BL102),.BLN(BLN102),.WL(WL172));
sram_cell_6t_5 inst_cell_172_103 (.BL(BL103),.BLN(BLN103),.WL(WL172));
sram_cell_6t_5 inst_cell_172_104 (.BL(BL104),.BLN(BLN104),.WL(WL172));
sram_cell_6t_5 inst_cell_172_105 (.BL(BL105),.BLN(BLN105),.WL(WL172));
sram_cell_6t_5 inst_cell_172_106 (.BL(BL106),.BLN(BLN106),.WL(WL172));
sram_cell_6t_5 inst_cell_172_107 (.BL(BL107),.BLN(BLN107),.WL(WL172));
sram_cell_6t_5 inst_cell_172_108 (.BL(BL108),.BLN(BLN108),.WL(WL172));
sram_cell_6t_5 inst_cell_172_109 (.BL(BL109),.BLN(BLN109),.WL(WL172));
sram_cell_6t_5 inst_cell_172_110 (.BL(BL110),.BLN(BLN110),.WL(WL172));
sram_cell_6t_5 inst_cell_172_111 (.BL(BL111),.BLN(BLN111),.WL(WL172));
sram_cell_6t_5 inst_cell_172_112 (.BL(BL112),.BLN(BLN112),.WL(WL172));
sram_cell_6t_5 inst_cell_172_113 (.BL(BL113),.BLN(BLN113),.WL(WL172));
sram_cell_6t_5 inst_cell_172_114 (.BL(BL114),.BLN(BLN114),.WL(WL172));
sram_cell_6t_5 inst_cell_172_115 (.BL(BL115),.BLN(BLN115),.WL(WL172));
sram_cell_6t_5 inst_cell_172_116 (.BL(BL116),.BLN(BLN116),.WL(WL172));
sram_cell_6t_5 inst_cell_172_117 (.BL(BL117),.BLN(BLN117),.WL(WL172));
sram_cell_6t_5 inst_cell_172_118 (.BL(BL118),.BLN(BLN118),.WL(WL172));
sram_cell_6t_5 inst_cell_172_119 (.BL(BL119),.BLN(BLN119),.WL(WL172));
sram_cell_6t_5 inst_cell_172_120 (.BL(BL120),.BLN(BLN120),.WL(WL172));
sram_cell_6t_5 inst_cell_172_121 (.BL(BL121),.BLN(BLN121),.WL(WL172));
sram_cell_6t_5 inst_cell_172_122 (.BL(BL122),.BLN(BLN122),.WL(WL172));
sram_cell_6t_5 inst_cell_172_123 (.BL(BL123),.BLN(BLN123),.WL(WL172));
sram_cell_6t_5 inst_cell_172_124 (.BL(BL124),.BLN(BLN124),.WL(WL172));
sram_cell_6t_5 inst_cell_172_125 (.BL(BL125),.BLN(BLN125),.WL(WL172));
sram_cell_6t_5 inst_cell_172_126 (.BL(BL126),.BLN(BLN126),.WL(WL172));
sram_cell_6t_5 inst_cell_172_127 (.BL(BL127),.BLN(BLN127),.WL(WL172));
sram_cell_6t_5 inst_cell_173_0 (.BL(BL0),.BLN(BLN0),.WL(WL173));
sram_cell_6t_5 inst_cell_173_1 (.BL(BL1),.BLN(BLN1),.WL(WL173));
sram_cell_6t_5 inst_cell_173_2 (.BL(BL2),.BLN(BLN2),.WL(WL173));
sram_cell_6t_5 inst_cell_173_3 (.BL(BL3),.BLN(BLN3),.WL(WL173));
sram_cell_6t_5 inst_cell_173_4 (.BL(BL4),.BLN(BLN4),.WL(WL173));
sram_cell_6t_5 inst_cell_173_5 (.BL(BL5),.BLN(BLN5),.WL(WL173));
sram_cell_6t_5 inst_cell_173_6 (.BL(BL6),.BLN(BLN6),.WL(WL173));
sram_cell_6t_5 inst_cell_173_7 (.BL(BL7),.BLN(BLN7),.WL(WL173));
sram_cell_6t_5 inst_cell_173_8 (.BL(BL8),.BLN(BLN8),.WL(WL173));
sram_cell_6t_5 inst_cell_173_9 (.BL(BL9),.BLN(BLN9),.WL(WL173));
sram_cell_6t_5 inst_cell_173_10 (.BL(BL10),.BLN(BLN10),.WL(WL173));
sram_cell_6t_5 inst_cell_173_11 (.BL(BL11),.BLN(BLN11),.WL(WL173));
sram_cell_6t_5 inst_cell_173_12 (.BL(BL12),.BLN(BLN12),.WL(WL173));
sram_cell_6t_5 inst_cell_173_13 (.BL(BL13),.BLN(BLN13),.WL(WL173));
sram_cell_6t_5 inst_cell_173_14 (.BL(BL14),.BLN(BLN14),.WL(WL173));
sram_cell_6t_5 inst_cell_173_15 (.BL(BL15),.BLN(BLN15),.WL(WL173));
sram_cell_6t_5 inst_cell_173_16 (.BL(BL16),.BLN(BLN16),.WL(WL173));
sram_cell_6t_5 inst_cell_173_17 (.BL(BL17),.BLN(BLN17),.WL(WL173));
sram_cell_6t_5 inst_cell_173_18 (.BL(BL18),.BLN(BLN18),.WL(WL173));
sram_cell_6t_5 inst_cell_173_19 (.BL(BL19),.BLN(BLN19),.WL(WL173));
sram_cell_6t_5 inst_cell_173_20 (.BL(BL20),.BLN(BLN20),.WL(WL173));
sram_cell_6t_5 inst_cell_173_21 (.BL(BL21),.BLN(BLN21),.WL(WL173));
sram_cell_6t_5 inst_cell_173_22 (.BL(BL22),.BLN(BLN22),.WL(WL173));
sram_cell_6t_5 inst_cell_173_23 (.BL(BL23),.BLN(BLN23),.WL(WL173));
sram_cell_6t_5 inst_cell_173_24 (.BL(BL24),.BLN(BLN24),.WL(WL173));
sram_cell_6t_5 inst_cell_173_25 (.BL(BL25),.BLN(BLN25),.WL(WL173));
sram_cell_6t_5 inst_cell_173_26 (.BL(BL26),.BLN(BLN26),.WL(WL173));
sram_cell_6t_5 inst_cell_173_27 (.BL(BL27),.BLN(BLN27),.WL(WL173));
sram_cell_6t_5 inst_cell_173_28 (.BL(BL28),.BLN(BLN28),.WL(WL173));
sram_cell_6t_5 inst_cell_173_29 (.BL(BL29),.BLN(BLN29),.WL(WL173));
sram_cell_6t_5 inst_cell_173_30 (.BL(BL30),.BLN(BLN30),.WL(WL173));
sram_cell_6t_5 inst_cell_173_31 (.BL(BL31),.BLN(BLN31),.WL(WL173));
sram_cell_6t_5 inst_cell_173_32 (.BL(BL32),.BLN(BLN32),.WL(WL173));
sram_cell_6t_5 inst_cell_173_33 (.BL(BL33),.BLN(BLN33),.WL(WL173));
sram_cell_6t_5 inst_cell_173_34 (.BL(BL34),.BLN(BLN34),.WL(WL173));
sram_cell_6t_5 inst_cell_173_35 (.BL(BL35),.BLN(BLN35),.WL(WL173));
sram_cell_6t_5 inst_cell_173_36 (.BL(BL36),.BLN(BLN36),.WL(WL173));
sram_cell_6t_5 inst_cell_173_37 (.BL(BL37),.BLN(BLN37),.WL(WL173));
sram_cell_6t_5 inst_cell_173_38 (.BL(BL38),.BLN(BLN38),.WL(WL173));
sram_cell_6t_5 inst_cell_173_39 (.BL(BL39),.BLN(BLN39),.WL(WL173));
sram_cell_6t_5 inst_cell_173_40 (.BL(BL40),.BLN(BLN40),.WL(WL173));
sram_cell_6t_5 inst_cell_173_41 (.BL(BL41),.BLN(BLN41),.WL(WL173));
sram_cell_6t_5 inst_cell_173_42 (.BL(BL42),.BLN(BLN42),.WL(WL173));
sram_cell_6t_5 inst_cell_173_43 (.BL(BL43),.BLN(BLN43),.WL(WL173));
sram_cell_6t_5 inst_cell_173_44 (.BL(BL44),.BLN(BLN44),.WL(WL173));
sram_cell_6t_5 inst_cell_173_45 (.BL(BL45),.BLN(BLN45),.WL(WL173));
sram_cell_6t_5 inst_cell_173_46 (.BL(BL46),.BLN(BLN46),.WL(WL173));
sram_cell_6t_5 inst_cell_173_47 (.BL(BL47),.BLN(BLN47),.WL(WL173));
sram_cell_6t_5 inst_cell_173_48 (.BL(BL48),.BLN(BLN48),.WL(WL173));
sram_cell_6t_5 inst_cell_173_49 (.BL(BL49),.BLN(BLN49),.WL(WL173));
sram_cell_6t_5 inst_cell_173_50 (.BL(BL50),.BLN(BLN50),.WL(WL173));
sram_cell_6t_5 inst_cell_173_51 (.BL(BL51),.BLN(BLN51),.WL(WL173));
sram_cell_6t_5 inst_cell_173_52 (.BL(BL52),.BLN(BLN52),.WL(WL173));
sram_cell_6t_5 inst_cell_173_53 (.BL(BL53),.BLN(BLN53),.WL(WL173));
sram_cell_6t_5 inst_cell_173_54 (.BL(BL54),.BLN(BLN54),.WL(WL173));
sram_cell_6t_5 inst_cell_173_55 (.BL(BL55),.BLN(BLN55),.WL(WL173));
sram_cell_6t_5 inst_cell_173_56 (.BL(BL56),.BLN(BLN56),.WL(WL173));
sram_cell_6t_5 inst_cell_173_57 (.BL(BL57),.BLN(BLN57),.WL(WL173));
sram_cell_6t_5 inst_cell_173_58 (.BL(BL58),.BLN(BLN58),.WL(WL173));
sram_cell_6t_5 inst_cell_173_59 (.BL(BL59),.BLN(BLN59),.WL(WL173));
sram_cell_6t_5 inst_cell_173_60 (.BL(BL60),.BLN(BLN60),.WL(WL173));
sram_cell_6t_5 inst_cell_173_61 (.BL(BL61),.BLN(BLN61),.WL(WL173));
sram_cell_6t_5 inst_cell_173_62 (.BL(BL62),.BLN(BLN62),.WL(WL173));
sram_cell_6t_5 inst_cell_173_63 (.BL(BL63),.BLN(BLN63),.WL(WL173));
sram_cell_6t_5 inst_cell_173_64 (.BL(BL64),.BLN(BLN64),.WL(WL173));
sram_cell_6t_5 inst_cell_173_65 (.BL(BL65),.BLN(BLN65),.WL(WL173));
sram_cell_6t_5 inst_cell_173_66 (.BL(BL66),.BLN(BLN66),.WL(WL173));
sram_cell_6t_5 inst_cell_173_67 (.BL(BL67),.BLN(BLN67),.WL(WL173));
sram_cell_6t_5 inst_cell_173_68 (.BL(BL68),.BLN(BLN68),.WL(WL173));
sram_cell_6t_5 inst_cell_173_69 (.BL(BL69),.BLN(BLN69),.WL(WL173));
sram_cell_6t_5 inst_cell_173_70 (.BL(BL70),.BLN(BLN70),.WL(WL173));
sram_cell_6t_5 inst_cell_173_71 (.BL(BL71),.BLN(BLN71),.WL(WL173));
sram_cell_6t_5 inst_cell_173_72 (.BL(BL72),.BLN(BLN72),.WL(WL173));
sram_cell_6t_5 inst_cell_173_73 (.BL(BL73),.BLN(BLN73),.WL(WL173));
sram_cell_6t_5 inst_cell_173_74 (.BL(BL74),.BLN(BLN74),.WL(WL173));
sram_cell_6t_5 inst_cell_173_75 (.BL(BL75),.BLN(BLN75),.WL(WL173));
sram_cell_6t_5 inst_cell_173_76 (.BL(BL76),.BLN(BLN76),.WL(WL173));
sram_cell_6t_5 inst_cell_173_77 (.BL(BL77),.BLN(BLN77),.WL(WL173));
sram_cell_6t_5 inst_cell_173_78 (.BL(BL78),.BLN(BLN78),.WL(WL173));
sram_cell_6t_5 inst_cell_173_79 (.BL(BL79),.BLN(BLN79),.WL(WL173));
sram_cell_6t_5 inst_cell_173_80 (.BL(BL80),.BLN(BLN80),.WL(WL173));
sram_cell_6t_5 inst_cell_173_81 (.BL(BL81),.BLN(BLN81),.WL(WL173));
sram_cell_6t_5 inst_cell_173_82 (.BL(BL82),.BLN(BLN82),.WL(WL173));
sram_cell_6t_5 inst_cell_173_83 (.BL(BL83),.BLN(BLN83),.WL(WL173));
sram_cell_6t_5 inst_cell_173_84 (.BL(BL84),.BLN(BLN84),.WL(WL173));
sram_cell_6t_5 inst_cell_173_85 (.BL(BL85),.BLN(BLN85),.WL(WL173));
sram_cell_6t_5 inst_cell_173_86 (.BL(BL86),.BLN(BLN86),.WL(WL173));
sram_cell_6t_5 inst_cell_173_87 (.BL(BL87),.BLN(BLN87),.WL(WL173));
sram_cell_6t_5 inst_cell_173_88 (.BL(BL88),.BLN(BLN88),.WL(WL173));
sram_cell_6t_5 inst_cell_173_89 (.BL(BL89),.BLN(BLN89),.WL(WL173));
sram_cell_6t_5 inst_cell_173_90 (.BL(BL90),.BLN(BLN90),.WL(WL173));
sram_cell_6t_5 inst_cell_173_91 (.BL(BL91),.BLN(BLN91),.WL(WL173));
sram_cell_6t_5 inst_cell_173_92 (.BL(BL92),.BLN(BLN92),.WL(WL173));
sram_cell_6t_5 inst_cell_173_93 (.BL(BL93),.BLN(BLN93),.WL(WL173));
sram_cell_6t_5 inst_cell_173_94 (.BL(BL94),.BLN(BLN94),.WL(WL173));
sram_cell_6t_5 inst_cell_173_95 (.BL(BL95),.BLN(BLN95),.WL(WL173));
sram_cell_6t_5 inst_cell_173_96 (.BL(BL96),.BLN(BLN96),.WL(WL173));
sram_cell_6t_5 inst_cell_173_97 (.BL(BL97),.BLN(BLN97),.WL(WL173));
sram_cell_6t_5 inst_cell_173_98 (.BL(BL98),.BLN(BLN98),.WL(WL173));
sram_cell_6t_5 inst_cell_173_99 (.BL(BL99),.BLN(BLN99),.WL(WL173));
sram_cell_6t_5 inst_cell_173_100 (.BL(BL100),.BLN(BLN100),.WL(WL173));
sram_cell_6t_5 inst_cell_173_101 (.BL(BL101),.BLN(BLN101),.WL(WL173));
sram_cell_6t_5 inst_cell_173_102 (.BL(BL102),.BLN(BLN102),.WL(WL173));
sram_cell_6t_5 inst_cell_173_103 (.BL(BL103),.BLN(BLN103),.WL(WL173));
sram_cell_6t_5 inst_cell_173_104 (.BL(BL104),.BLN(BLN104),.WL(WL173));
sram_cell_6t_5 inst_cell_173_105 (.BL(BL105),.BLN(BLN105),.WL(WL173));
sram_cell_6t_5 inst_cell_173_106 (.BL(BL106),.BLN(BLN106),.WL(WL173));
sram_cell_6t_5 inst_cell_173_107 (.BL(BL107),.BLN(BLN107),.WL(WL173));
sram_cell_6t_5 inst_cell_173_108 (.BL(BL108),.BLN(BLN108),.WL(WL173));
sram_cell_6t_5 inst_cell_173_109 (.BL(BL109),.BLN(BLN109),.WL(WL173));
sram_cell_6t_5 inst_cell_173_110 (.BL(BL110),.BLN(BLN110),.WL(WL173));
sram_cell_6t_5 inst_cell_173_111 (.BL(BL111),.BLN(BLN111),.WL(WL173));
sram_cell_6t_5 inst_cell_173_112 (.BL(BL112),.BLN(BLN112),.WL(WL173));
sram_cell_6t_5 inst_cell_173_113 (.BL(BL113),.BLN(BLN113),.WL(WL173));
sram_cell_6t_5 inst_cell_173_114 (.BL(BL114),.BLN(BLN114),.WL(WL173));
sram_cell_6t_5 inst_cell_173_115 (.BL(BL115),.BLN(BLN115),.WL(WL173));
sram_cell_6t_5 inst_cell_173_116 (.BL(BL116),.BLN(BLN116),.WL(WL173));
sram_cell_6t_5 inst_cell_173_117 (.BL(BL117),.BLN(BLN117),.WL(WL173));
sram_cell_6t_5 inst_cell_173_118 (.BL(BL118),.BLN(BLN118),.WL(WL173));
sram_cell_6t_5 inst_cell_173_119 (.BL(BL119),.BLN(BLN119),.WL(WL173));
sram_cell_6t_5 inst_cell_173_120 (.BL(BL120),.BLN(BLN120),.WL(WL173));
sram_cell_6t_5 inst_cell_173_121 (.BL(BL121),.BLN(BLN121),.WL(WL173));
sram_cell_6t_5 inst_cell_173_122 (.BL(BL122),.BLN(BLN122),.WL(WL173));
sram_cell_6t_5 inst_cell_173_123 (.BL(BL123),.BLN(BLN123),.WL(WL173));
sram_cell_6t_5 inst_cell_173_124 (.BL(BL124),.BLN(BLN124),.WL(WL173));
sram_cell_6t_5 inst_cell_173_125 (.BL(BL125),.BLN(BLN125),.WL(WL173));
sram_cell_6t_5 inst_cell_173_126 (.BL(BL126),.BLN(BLN126),.WL(WL173));
sram_cell_6t_5 inst_cell_173_127 (.BL(BL127),.BLN(BLN127),.WL(WL173));
sram_cell_6t_5 inst_cell_174_0 (.BL(BL0),.BLN(BLN0),.WL(WL174));
sram_cell_6t_5 inst_cell_174_1 (.BL(BL1),.BLN(BLN1),.WL(WL174));
sram_cell_6t_5 inst_cell_174_2 (.BL(BL2),.BLN(BLN2),.WL(WL174));
sram_cell_6t_5 inst_cell_174_3 (.BL(BL3),.BLN(BLN3),.WL(WL174));
sram_cell_6t_5 inst_cell_174_4 (.BL(BL4),.BLN(BLN4),.WL(WL174));
sram_cell_6t_5 inst_cell_174_5 (.BL(BL5),.BLN(BLN5),.WL(WL174));
sram_cell_6t_5 inst_cell_174_6 (.BL(BL6),.BLN(BLN6),.WL(WL174));
sram_cell_6t_5 inst_cell_174_7 (.BL(BL7),.BLN(BLN7),.WL(WL174));
sram_cell_6t_5 inst_cell_174_8 (.BL(BL8),.BLN(BLN8),.WL(WL174));
sram_cell_6t_5 inst_cell_174_9 (.BL(BL9),.BLN(BLN9),.WL(WL174));
sram_cell_6t_5 inst_cell_174_10 (.BL(BL10),.BLN(BLN10),.WL(WL174));
sram_cell_6t_5 inst_cell_174_11 (.BL(BL11),.BLN(BLN11),.WL(WL174));
sram_cell_6t_5 inst_cell_174_12 (.BL(BL12),.BLN(BLN12),.WL(WL174));
sram_cell_6t_5 inst_cell_174_13 (.BL(BL13),.BLN(BLN13),.WL(WL174));
sram_cell_6t_5 inst_cell_174_14 (.BL(BL14),.BLN(BLN14),.WL(WL174));
sram_cell_6t_5 inst_cell_174_15 (.BL(BL15),.BLN(BLN15),.WL(WL174));
sram_cell_6t_5 inst_cell_174_16 (.BL(BL16),.BLN(BLN16),.WL(WL174));
sram_cell_6t_5 inst_cell_174_17 (.BL(BL17),.BLN(BLN17),.WL(WL174));
sram_cell_6t_5 inst_cell_174_18 (.BL(BL18),.BLN(BLN18),.WL(WL174));
sram_cell_6t_5 inst_cell_174_19 (.BL(BL19),.BLN(BLN19),.WL(WL174));
sram_cell_6t_5 inst_cell_174_20 (.BL(BL20),.BLN(BLN20),.WL(WL174));
sram_cell_6t_5 inst_cell_174_21 (.BL(BL21),.BLN(BLN21),.WL(WL174));
sram_cell_6t_5 inst_cell_174_22 (.BL(BL22),.BLN(BLN22),.WL(WL174));
sram_cell_6t_5 inst_cell_174_23 (.BL(BL23),.BLN(BLN23),.WL(WL174));
sram_cell_6t_5 inst_cell_174_24 (.BL(BL24),.BLN(BLN24),.WL(WL174));
sram_cell_6t_5 inst_cell_174_25 (.BL(BL25),.BLN(BLN25),.WL(WL174));
sram_cell_6t_5 inst_cell_174_26 (.BL(BL26),.BLN(BLN26),.WL(WL174));
sram_cell_6t_5 inst_cell_174_27 (.BL(BL27),.BLN(BLN27),.WL(WL174));
sram_cell_6t_5 inst_cell_174_28 (.BL(BL28),.BLN(BLN28),.WL(WL174));
sram_cell_6t_5 inst_cell_174_29 (.BL(BL29),.BLN(BLN29),.WL(WL174));
sram_cell_6t_5 inst_cell_174_30 (.BL(BL30),.BLN(BLN30),.WL(WL174));
sram_cell_6t_5 inst_cell_174_31 (.BL(BL31),.BLN(BLN31),.WL(WL174));
sram_cell_6t_5 inst_cell_174_32 (.BL(BL32),.BLN(BLN32),.WL(WL174));
sram_cell_6t_5 inst_cell_174_33 (.BL(BL33),.BLN(BLN33),.WL(WL174));
sram_cell_6t_5 inst_cell_174_34 (.BL(BL34),.BLN(BLN34),.WL(WL174));
sram_cell_6t_5 inst_cell_174_35 (.BL(BL35),.BLN(BLN35),.WL(WL174));
sram_cell_6t_5 inst_cell_174_36 (.BL(BL36),.BLN(BLN36),.WL(WL174));
sram_cell_6t_5 inst_cell_174_37 (.BL(BL37),.BLN(BLN37),.WL(WL174));
sram_cell_6t_5 inst_cell_174_38 (.BL(BL38),.BLN(BLN38),.WL(WL174));
sram_cell_6t_5 inst_cell_174_39 (.BL(BL39),.BLN(BLN39),.WL(WL174));
sram_cell_6t_5 inst_cell_174_40 (.BL(BL40),.BLN(BLN40),.WL(WL174));
sram_cell_6t_5 inst_cell_174_41 (.BL(BL41),.BLN(BLN41),.WL(WL174));
sram_cell_6t_5 inst_cell_174_42 (.BL(BL42),.BLN(BLN42),.WL(WL174));
sram_cell_6t_5 inst_cell_174_43 (.BL(BL43),.BLN(BLN43),.WL(WL174));
sram_cell_6t_5 inst_cell_174_44 (.BL(BL44),.BLN(BLN44),.WL(WL174));
sram_cell_6t_5 inst_cell_174_45 (.BL(BL45),.BLN(BLN45),.WL(WL174));
sram_cell_6t_5 inst_cell_174_46 (.BL(BL46),.BLN(BLN46),.WL(WL174));
sram_cell_6t_5 inst_cell_174_47 (.BL(BL47),.BLN(BLN47),.WL(WL174));
sram_cell_6t_5 inst_cell_174_48 (.BL(BL48),.BLN(BLN48),.WL(WL174));
sram_cell_6t_5 inst_cell_174_49 (.BL(BL49),.BLN(BLN49),.WL(WL174));
sram_cell_6t_5 inst_cell_174_50 (.BL(BL50),.BLN(BLN50),.WL(WL174));
sram_cell_6t_5 inst_cell_174_51 (.BL(BL51),.BLN(BLN51),.WL(WL174));
sram_cell_6t_5 inst_cell_174_52 (.BL(BL52),.BLN(BLN52),.WL(WL174));
sram_cell_6t_5 inst_cell_174_53 (.BL(BL53),.BLN(BLN53),.WL(WL174));
sram_cell_6t_5 inst_cell_174_54 (.BL(BL54),.BLN(BLN54),.WL(WL174));
sram_cell_6t_5 inst_cell_174_55 (.BL(BL55),.BLN(BLN55),.WL(WL174));
sram_cell_6t_5 inst_cell_174_56 (.BL(BL56),.BLN(BLN56),.WL(WL174));
sram_cell_6t_5 inst_cell_174_57 (.BL(BL57),.BLN(BLN57),.WL(WL174));
sram_cell_6t_5 inst_cell_174_58 (.BL(BL58),.BLN(BLN58),.WL(WL174));
sram_cell_6t_5 inst_cell_174_59 (.BL(BL59),.BLN(BLN59),.WL(WL174));
sram_cell_6t_5 inst_cell_174_60 (.BL(BL60),.BLN(BLN60),.WL(WL174));
sram_cell_6t_5 inst_cell_174_61 (.BL(BL61),.BLN(BLN61),.WL(WL174));
sram_cell_6t_5 inst_cell_174_62 (.BL(BL62),.BLN(BLN62),.WL(WL174));
sram_cell_6t_5 inst_cell_174_63 (.BL(BL63),.BLN(BLN63),.WL(WL174));
sram_cell_6t_5 inst_cell_174_64 (.BL(BL64),.BLN(BLN64),.WL(WL174));
sram_cell_6t_5 inst_cell_174_65 (.BL(BL65),.BLN(BLN65),.WL(WL174));
sram_cell_6t_5 inst_cell_174_66 (.BL(BL66),.BLN(BLN66),.WL(WL174));
sram_cell_6t_5 inst_cell_174_67 (.BL(BL67),.BLN(BLN67),.WL(WL174));
sram_cell_6t_5 inst_cell_174_68 (.BL(BL68),.BLN(BLN68),.WL(WL174));
sram_cell_6t_5 inst_cell_174_69 (.BL(BL69),.BLN(BLN69),.WL(WL174));
sram_cell_6t_5 inst_cell_174_70 (.BL(BL70),.BLN(BLN70),.WL(WL174));
sram_cell_6t_5 inst_cell_174_71 (.BL(BL71),.BLN(BLN71),.WL(WL174));
sram_cell_6t_5 inst_cell_174_72 (.BL(BL72),.BLN(BLN72),.WL(WL174));
sram_cell_6t_5 inst_cell_174_73 (.BL(BL73),.BLN(BLN73),.WL(WL174));
sram_cell_6t_5 inst_cell_174_74 (.BL(BL74),.BLN(BLN74),.WL(WL174));
sram_cell_6t_5 inst_cell_174_75 (.BL(BL75),.BLN(BLN75),.WL(WL174));
sram_cell_6t_5 inst_cell_174_76 (.BL(BL76),.BLN(BLN76),.WL(WL174));
sram_cell_6t_5 inst_cell_174_77 (.BL(BL77),.BLN(BLN77),.WL(WL174));
sram_cell_6t_5 inst_cell_174_78 (.BL(BL78),.BLN(BLN78),.WL(WL174));
sram_cell_6t_5 inst_cell_174_79 (.BL(BL79),.BLN(BLN79),.WL(WL174));
sram_cell_6t_5 inst_cell_174_80 (.BL(BL80),.BLN(BLN80),.WL(WL174));
sram_cell_6t_5 inst_cell_174_81 (.BL(BL81),.BLN(BLN81),.WL(WL174));
sram_cell_6t_5 inst_cell_174_82 (.BL(BL82),.BLN(BLN82),.WL(WL174));
sram_cell_6t_5 inst_cell_174_83 (.BL(BL83),.BLN(BLN83),.WL(WL174));
sram_cell_6t_5 inst_cell_174_84 (.BL(BL84),.BLN(BLN84),.WL(WL174));
sram_cell_6t_5 inst_cell_174_85 (.BL(BL85),.BLN(BLN85),.WL(WL174));
sram_cell_6t_5 inst_cell_174_86 (.BL(BL86),.BLN(BLN86),.WL(WL174));
sram_cell_6t_5 inst_cell_174_87 (.BL(BL87),.BLN(BLN87),.WL(WL174));
sram_cell_6t_5 inst_cell_174_88 (.BL(BL88),.BLN(BLN88),.WL(WL174));
sram_cell_6t_5 inst_cell_174_89 (.BL(BL89),.BLN(BLN89),.WL(WL174));
sram_cell_6t_5 inst_cell_174_90 (.BL(BL90),.BLN(BLN90),.WL(WL174));
sram_cell_6t_5 inst_cell_174_91 (.BL(BL91),.BLN(BLN91),.WL(WL174));
sram_cell_6t_5 inst_cell_174_92 (.BL(BL92),.BLN(BLN92),.WL(WL174));
sram_cell_6t_5 inst_cell_174_93 (.BL(BL93),.BLN(BLN93),.WL(WL174));
sram_cell_6t_5 inst_cell_174_94 (.BL(BL94),.BLN(BLN94),.WL(WL174));
sram_cell_6t_5 inst_cell_174_95 (.BL(BL95),.BLN(BLN95),.WL(WL174));
sram_cell_6t_5 inst_cell_174_96 (.BL(BL96),.BLN(BLN96),.WL(WL174));
sram_cell_6t_5 inst_cell_174_97 (.BL(BL97),.BLN(BLN97),.WL(WL174));
sram_cell_6t_5 inst_cell_174_98 (.BL(BL98),.BLN(BLN98),.WL(WL174));
sram_cell_6t_5 inst_cell_174_99 (.BL(BL99),.BLN(BLN99),.WL(WL174));
sram_cell_6t_5 inst_cell_174_100 (.BL(BL100),.BLN(BLN100),.WL(WL174));
sram_cell_6t_5 inst_cell_174_101 (.BL(BL101),.BLN(BLN101),.WL(WL174));
sram_cell_6t_5 inst_cell_174_102 (.BL(BL102),.BLN(BLN102),.WL(WL174));
sram_cell_6t_5 inst_cell_174_103 (.BL(BL103),.BLN(BLN103),.WL(WL174));
sram_cell_6t_5 inst_cell_174_104 (.BL(BL104),.BLN(BLN104),.WL(WL174));
sram_cell_6t_5 inst_cell_174_105 (.BL(BL105),.BLN(BLN105),.WL(WL174));
sram_cell_6t_5 inst_cell_174_106 (.BL(BL106),.BLN(BLN106),.WL(WL174));
sram_cell_6t_5 inst_cell_174_107 (.BL(BL107),.BLN(BLN107),.WL(WL174));
sram_cell_6t_5 inst_cell_174_108 (.BL(BL108),.BLN(BLN108),.WL(WL174));
sram_cell_6t_5 inst_cell_174_109 (.BL(BL109),.BLN(BLN109),.WL(WL174));
sram_cell_6t_5 inst_cell_174_110 (.BL(BL110),.BLN(BLN110),.WL(WL174));
sram_cell_6t_5 inst_cell_174_111 (.BL(BL111),.BLN(BLN111),.WL(WL174));
sram_cell_6t_5 inst_cell_174_112 (.BL(BL112),.BLN(BLN112),.WL(WL174));
sram_cell_6t_5 inst_cell_174_113 (.BL(BL113),.BLN(BLN113),.WL(WL174));
sram_cell_6t_5 inst_cell_174_114 (.BL(BL114),.BLN(BLN114),.WL(WL174));
sram_cell_6t_5 inst_cell_174_115 (.BL(BL115),.BLN(BLN115),.WL(WL174));
sram_cell_6t_5 inst_cell_174_116 (.BL(BL116),.BLN(BLN116),.WL(WL174));
sram_cell_6t_5 inst_cell_174_117 (.BL(BL117),.BLN(BLN117),.WL(WL174));
sram_cell_6t_5 inst_cell_174_118 (.BL(BL118),.BLN(BLN118),.WL(WL174));
sram_cell_6t_5 inst_cell_174_119 (.BL(BL119),.BLN(BLN119),.WL(WL174));
sram_cell_6t_5 inst_cell_174_120 (.BL(BL120),.BLN(BLN120),.WL(WL174));
sram_cell_6t_5 inst_cell_174_121 (.BL(BL121),.BLN(BLN121),.WL(WL174));
sram_cell_6t_5 inst_cell_174_122 (.BL(BL122),.BLN(BLN122),.WL(WL174));
sram_cell_6t_5 inst_cell_174_123 (.BL(BL123),.BLN(BLN123),.WL(WL174));
sram_cell_6t_5 inst_cell_174_124 (.BL(BL124),.BLN(BLN124),.WL(WL174));
sram_cell_6t_5 inst_cell_174_125 (.BL(BL125),.BLN(BLN125),.WL(WL174));
sram_cell_6t_5 inst_cell_174_126 (.BL(BL126),.BLN(BLN126),.WL(WL174));
sram_cell_6t_5 inst_cell_174_127 (.BL(BL127),.BLN(BLN127),.WL(WL174));
sram_cell_6t_5 inst_cell_175_0 (.BL(BL0),.BLN(BLN0),.WL(WL175));
sram_cell_6t_5 inst_cell_175_1 (.BL(BL1),.BLN(BLN1),.WL(WL175));
sram_cell_6t_5 inst_cell_175_2 (.BL(BL2),.BLN(BLN2),.WL(WL175));
sram_cell_6t_5 inst_cell_175_3 (.BL(BL3),.BLN(BLN3),.WL(WL175));
sram_cell_6t_5 inst_cell_175_4 (.BL(BL4),.BLN(BLN4),.WL(WL175));
sram_cell_6t_5 inst_cell_175_5 (.BL(BL5),.BLN(BLN5),.WL(WL175));
sram_cell_6t_5 inst_cell_175_6 (.BL(BL6),.BLN(BLN6),.WL(WL175));
sram_cell_6t_5 inst_cell_175_7 (.BL(BL7),.BLN(BLN7),.WL(WL175));
sram_cell_6t_5 inst_cell_175_8 (.BL(BL8),.BLN(BLN8),.WL(WL175));
sram_cell_6t_5 inst_cell_175_9 (.BL(BL9),.BLN(BLN9),.WL(WL175));
sram_cell_6t_5 inst_cell_175_10 (.BL(BL10),.BLN(BLN10),.WL(WL175));
sram_cell_6t_5 inst_cell_175_11 (.BL(BL11),.BLN(BLN11),.WL(WL175));
sram_cell_6t_5 inst_cell_175_12 (.BL(BL12),.BLN(BLN12),.WL(WL175));
sram_cell_6t_5 inst_cell_175_13 (.BL(BL13),.BLN(BLN13),.WL(WL175));
sram_cell_6t_5 inst_cell_175_14 (.BL(BL14),.BLN(BLN14),.WL(WL175));
sram_cell_6t_5 inst_cell_175_15 (.BL(BL15),.BLN(BLN15),.WL(WL175));
sram_cell_6t_5 inst_cell_175_16 (.BL(BL16),.BLN(BLN16),.WL(WL175));
sram_cell_6t_5 inst_cell_175_17 (.BL(BL17),.BLN(BLN17),.WL(WL175));
sram_cell_6t_5 inst_cell_175_18 (.BL(BL18),.BLN(BLN18),.WL(WL175));
sram_cell_6t_5 inst_cell_175_19 (.BL(BL19),.BLN(BLN19),.WL(WL175));
sram_cell_6t_5 inst_cell_175_20 (.BL(BL20),.BLN(BLN20),.WL(WL175));
sram_cell_6t_5 inst_cell_175_21 (.BL(BL21),.BLN(BLN21),.WL(WL175));
sram_cell_6t_5 inst_cell_175_22 (.BL(BL22),.BLN(BLN22),.WL(WL175));
sram_cell_6t_5 inst_cell_175_23 (.BL(BL23),.BLN(BLN23),.WL(WL175));
sram_cell_6t_5 inst_cell_175_24 (.BL(BL24),.BLN(BLN24),.WL(WL175));
sram_cell_6t_5 inst_cell_175_25 (.BL(BL25),.BLN(BLN25),.WL(WL175));
sram_cell_6t_5 inst_cell_175_26 (.BL(BL26),.BLN(BLN26),.WL(WL175));
sram_cell_6t_5 inst_cell_175_27 (.BL(BL27),.BLN(BLN27),.WL(WL175));
sram_cell_6t_5 inst_cell_175_28 (.BL(BL28),.BLN(BLN28),.WL(WL175));
sram_cell_6t_5 inst_cell_175_29 (.BL(BL29),.BLN(BLN29),.WL(WL175));
sram_cell_6t_5 inst_cell_175_30 (.BL(BL30),.BLN(BLN30),.WL(WL175));
sram_cell_6t_5 inst_cell_175_31 (.BL(BL31),.BLN(BLN31),.WL(WL175));
sram_cell_6t_5 inst_cell_175_32 (.BL(BL32),.BLN(BLN32),.WL(WL175));
sram_cell_6t_5 inst_cell_175_33 (.BL(BL33),.BLN(BLN33),.WL(WL175));
sram_cell_6t_5 inst_cell_175_34 (.BL(BL34),.BLN(BLN34),.WL(WL175));
sram_cell_6t_5 inst_cell_175_35 (.BL(BL35),.BLN(BLN35),.WL(WL175));
sram_cell_6t_5 inst_cell_175_36 (.BL(BL36),.BLN(BLN36),.WL(WL175));
sram_cell_6t_5 inst_cell_175_37 (.BL(BL37),.BLN(BLN37),.WL(WL175));
sram_cell_6t_5 inst_cell_175_38 (.BL(BL38),.BLN(BLN38),.WL(WL175));
sram_cell_6t_5 inst_cell_175_39 (.BL(BL39),.BLN(BLN39),.WL(WL175));
sram_cell_6t_5 inst_cell_175_40 (.BL(BL40),.BLN(BLN40),.WL(WL175));
sram_cell_6t_5 inst_cell_175_41 (.BL(BL41),.BLN(BLN41),.WL(WL175));
sram_cell_6t_5 inst_cell_175_42 (.BL(BL42),.BLN(BLN42),.WL(WL175));
sram_cell_6t_5 inst_cell_175_43 (.BL(BL43),.BLN(BLN43),.WL(WL175));
sram_cell_6t_5 inst_cell_175_44 (.BL(BL44),.BLN(BLN44),.WL(WL175));
sram_cell_6t_5 inst_cell_175_45 (.BL(BL45),.BLN(BLN45),.WL(WL175));
sram_cell_6t_5 inst_cell_175_46 (.BL(BL46),.BLN(BLN46),.WL(WL175));
sram_cell_6t_5 inst_cell_175_47 (.BL(BL47),.BLN(BLN47),.WL(WL175));
sram_cell_6t_5 inst_cell_175_48 (.BL(BL48),.BLN(BLN48),.WL(WL175));
sram_cell_6t_5 inst_cell_175_49 (.BL(BL49),.BLN(BLN49),.WL(WL175));
sram_cell_6t_5 inst_cell_175_50 (.BL(BL50),.BLN(BLN50),.WL(WL175));
sram_cell_6t_5 inst_cell_175_51 (.BL(BL51),.BLN(BLN51),.WL(WL175));
sram_cell_6t_5 inst_cell_175_52 (.BL(BL52),.BLN(BLN52),.WL(WL175));
sram_cell_6t_5 inst_cell_175_53 (.BL(BL53),.BLN(BLN53),.WL(WL175));
sram_cell_6t_5 inst_cell_175_54 (.BL(BL54),.BLN(BLN54),.WL(WL175));
sram_cell_6t_5 inst_cell_175_55 (.BL(BL55),.BLN(BLN55),.WL(WL175));
sram_cell_6t_5 inst_cell_175_56 (.BL(BL56),.BLN(BLN56),.WL(WL175));
sram_cell_6t_5 inst_cell_175_57 (.BL(BL57),.BLN(BLN57),.WL(WL175));
sram_cell_6t_5 inst_cell_175_58 (.BL(BL58),.BLN(BLN58),.WL(WL175));
sram_cell_6t_5 inst_cell_175_59 (.BL(BL59),.BLN(BLN59),.WL(WL175));
sram_cell_6t_5 inst_cell_175_60 (.BL(BL60),.BLN(BLN60),.WL(WL175));
sram_cell_6t_5 inst_cell_175_61 (.BL(BL61),.BLN(BLN61),.WL(WL175));
sram_cell_6t_5 inst_cell_175_62 (.BL(BL62),.BLN(BLN62),.WL(WL175));
sram_cell_6t_5 inst_cell_175_63 (.BL(BL63),.BLN(BLN63),.WL(WL175));
sram_cell_6t_5 inst_cell_175_64 (.BL(BL64),.BLN(BLN64),.WL(WL175));
sram_cell_6t_5 inst_cell_175_65 (.BL(BL65),.BLN(BLN65),.WL(WL175));
sram_cell_6t_5 inst_cell_175_66 (.BL(BL66),.BLN(BLN66),.WL(WL175));
sram_cell_6t_5 inst_cell_175_67 (.BL(BL67),.BLN(BLN67),.WL(WL175));
sram_cell_6t_5 inst_cell_175_68 (.BL(BL68),.BLN(BLN68),.WL(WL175));
sram_cell_6t_5 inst_cell_175_69 (.BL(BL69),.BLN(BLN69),.WL(WL175));
sram_cell_6t_5 inst_cell_175_70 (.BL(BL70),.BLN(BLN70),.WL(WL175));
sram_cell_6t_5 inst_cell_175_71 (.BL(BL71),.BLN(BLN71),.WL(WL175));
sram_cell_6t_5 inst_cell_175_72 (.BL(BL72),.BLN(BLN72),.WL(WL175));
sram_cell_6t_5 inst_cell_175_73 (.BL(BL73),.BLN(BLN73),.WL(WL175));
sram_cell_6t_5 inst_cell_175_74 (.BL(BL74),.BLN(BLN74),.WL(WL175));
sram_cell_6t_5 inst_cell_175_75 (.BL(BL75),.BLN(BLN75),.WL(WL175));
sram_cell_6t_5 inst_cell_175_76 (.BL(BL76),.BLN(BLN76),.WL(WL175));
sram_cell_6t_5 inst_cell_175_77 (.BL(BL77),.BLN(BLN77),.WL(WL175));
sram_cell_6t_5 inst_cell_175_78 (.BL(BL78),.BLN(BLN78),.WL(WL175));
sram_cell_6t_5 inst_cell_175_79 (.BL(BL79),.BLN(BLN79),.WL(WL175));
sram_cell_6t_5 inst_cell_175_80 (.BL(BL80),.BLN(BLN80),.WL(WL175));
sram_cell_6t_5 inst_cell_175_81 (.BL(BL81),.BLN(BLN81),.WL(WL175));
sram_cell_6t_5 inst_cell_175_82 (.BL(BL82),.BLN(BLN82),.WL(WL175));
sram_cell_6t_5 inst_cell_175_83 (.BL(BL83),.BLN(BLN83),.WL(WL175));
sram_cell_6t_5 inst_cell_175_84 (.BL(BL84),.BLN(BLN84),.WL(WL175));
sram_cell_6t_5 inst_cell_175_85 (.BL(BL85),.BLN(BLN85),.WL(WL175));
sram_cell_6t_5 inst_cell_175_86 (.BL(BL86),.BLN(BLN86),.WL(WL175));
sram_cell_6t_5 inst_cell_175_87 (.BL(BL87),.BLN(BLN87),.WL(WL175));
sram_cell_6t_5 inst_cell_175_88 (.BL(BL88),.BLN(BLN88),.WL(WL175));
sram_cell_6t_5 inst_cell_175_89 (.BL(BL89),.BLN(BLN89),.WL(WL175));
sram_cell_6t_5 inst_cell_175_90 (.BL(BL90),.BLN(BLN90),.WL(WL175));
sram_cell_6t_5 inst_cell_175_91 (.BL(BL91),.BLN(BLN91),.WL(WL175));
sram_cell_6t_5 inst_cell_175_92 (.BL(BL92),.BLN(BLN92),.WL(WL175));
sram_cell_6t_5 inst_cell_175_93 (.BL(BL93),.BLN(BLN93),.WL(WL175));
sram_cell_6t_5 inst_cell_175_94 (.BL(BL94),.BLN(BLN94),.WL(WL175));
sram_cell_6t_5 inst_cell_175_95 (.BL(BL95),.BLN(BLN95),.WL(WL175));
sram_cell_6t_5 inst_cell_175_96 (.BL(BL96),.BLN(BLN96),.WL(WL175));
sram_cell_6t_5 inst_cell_175_97 (.BL(BL97),.BLN(BLN97),.WL(WL175));
sram_cell_6t_5 inst_cell_175_98 (.BL(BL98),.BLN(BLN98),.WL(WL175));
sram_cell_6t_5 inst_cell_175_99 (.BL(BL99),.BLN(BLN99),.WL(WL175));
sram_cell_6t_5 inst_cell_175_100 (.BL(BL100),.BLN(BLN100),.WL(WL175));
sram_cell_6t_5 inst_cell_175_101 (.BL(BL101),.BLN(BLN101),.WL(WL175));
sram_cell_6t_5 inst_cell_175_102 (.BL(BL102),.BLN(BLN102),.WL(WL175));
sram_cell_6t_5 inst_cell_175_103 (.BL(BL103),.BLN(BLN103),.WL(WL175));
sram_cell_6t_5 inst_cell_175_104 (.BL(BL104),.BLN(BLN104),.WL(WL175));
sram_cell_6t_5 inst_cell_175_105 (.BL(BL105),.BLN(BLN105),.WL(WL175));
sram_cell_6t_5 inst_cell_175_106 (.BL(BL106),.BLN(BLN106),.WL(WL175));
sram_cell_6t_5 inst_cell_175_107 (.BL(BL107),.BLN(BLN107),.WL(WL175));
sram_cell_6t_5 inst_cell_175_108 (.BL(BL108),.BLN(BLN108),.WL(WL175));
sram_cell_6t_5 inst_cell_175_109 (.BL(BL109),.BLN(BLN109),.WL(WL175));
sram_cell_6t_5 inst_cell_175_110 (.BL(BL110),.BLN(BLN110),.WL(WL175));
sram_cell_6t_5 inst_cell_175_111 (.BL(BL111),.BLN(BLN111),.WL(WL175));
sram_cell_6t_5 inst_cell_175_112 (.BL(BL112),.BLN(BLN112),.WL(WL175));
sram_cell_6t_5 inst_cell_175_113 (.BL(BL113),.BLN(BLN113),.WL(WL175));
sram_cell_6t_5 inst_cell_175_114 (.BL(BL114),.BLN(BLN114),.WL(WL175));
sram_cell_6t_5 inst_cell_175_115 (.BL(BL115),.BLN(BLN115),.WL(WL175));
sram_cell_6t_5 inst_cell_175_116 (.BL(BL116),.BLN(BLN116),.WL(WL175));
sram_cell_6t_5 inst_cell_175_117 (.BL(BL117),.BLN(BLN117),.WL(WL175));
sram_cell_6t_5 inst_cell_175_118 (.BL(BL118),.BLN(BLN118),.WL(WL175));
sram_cell_6t_5 inst_cell_175_119 (.BL(BL119),.BLN(BLN119),.WL(WL175));
sram_cell_6t_5 inst_cell_175_120 (.BL(BL120),.BLN(BLN120),.WL(WL175));
sram_cell_6t_5 inst_cell_175_121 (.BL(BL121),.BLN(BLN121),.WL(WL175));
sram_cell_6t_5 inst_cell_175_122 (.BL(BL122),.BLN(BLN122),.WL(WL175));
sram_cell_6t_5 inst_cell_175_123 (.BL(BL123),.BLN(BLN123),.WL(WL175));
sram_cell_6t_5 inst_cell_175_124 (.BL(BL124),.BLN(BLN124),.WL(WL175));
sram_cell_6t_5 inst_cell_175_125 (.BL(BL125),.BLN(BLN125),.WL(WL175));
sram_cell_6t_5 inst_cell_175_126 (.BL(BL126),.BLN(BLN126),.WL(WL175));
sram_cell_6t_5 inst_cell_175_127 (.BL(BL127),.BLN(BLN127),.WL(WL175));
sram_cell_6t_5 inst_cell_176_0 (.BL(BL0),.BLN(BLN0),.WL(WL176));
sram_cell_6t_5 inst_cell_176_1 (.BL(BL1),.BLN(BLN1),.WL(WL176));
sram_cell_6t_5 inst_cell_176_2 (.BL(BL2),.BLN(BLN2),.WL(WL176));
sram_cell_6t_5 inst_cell_176_3 (.BL(BL3),.BLN(BLN3),.WL(WL176));
sram_cell_6t_5 inst_cell_176_4 (.BL(BL4),.BLN(BLN4),.WL(WL176));
sram_cell_6t_5 inst_cell_176_5 (.BL(BL5),.BLN(BLN5),.WL(WL176));
sram_cell_6t_5 inst_cell_176_6 (.BL(BL6),.BLN(BLN6),.WL(WL176));
sram_cell_6t_5 inst_cell_176_7 (.BL(BL7),.BLN(BLN7),.WL(WL176));
sram_cell_6t_5 inst_cell_176_8 (.BL(BL8),.BLN(BLN8),.WL(WL176));
sram_cell_6t_5 inst_cell_176_9 (.BL(BL9),.BLN(BLN9),.WL(WL176));
sram_cell_6t_5 inst_cell_176_10 (.BL(BL10),.BLN(BLN10),.WL(WL176));
sram_cell_6t_5 inst_cell_176_11 (.BL(BL11),.BLN(BLN11),.WL(WL176));
sram_cell_6t_5 inst_cell_176_12 (.BL(BL12),.BLN(BLN12),.WL(WL176));
sram_cell_6t_5 inst_cell_176_13 (.BL(BL13),.BLN(BLN13),.WL(WL176));
sram_cell_6t_5 inst_cell_176_14 (.BL(BL14),.BLN(BLN14),.WL(WL176));
sram_cell_6t_5 inst_cell_176_15 (.BL(BL15),.BLN(BLN15),.WL(WL176));
sram_cell_6t_5 inst_cell_176_16 (.BL(BL16),.BLN(BLN16),.WL(WL176));
sram_cell_6t_5 inst_cell_176_17 (.BL(BL17),.BLN(BLN17),.WL(WL176));
sram_cell_6t_5 inst_cell_176_18 (.BL(BL18),.BLN(BLN18),.WL(WL176));
sram_cell_6t_5 inst_cell_176_19 (.BL(BL19),.BLN(BLN19),.WL(WL176));
sram_cell_6t_5 inst_cell_176_20 (.BL(BL20),.BLN(BLN20),.WL(WL176));
sram_cell_6t_5 inst_cell_176_21 (.BL(BL21),.BLN(BLN21),.WL(WL176));
sram_cell_6t_5 inst_cell_176_22 (.BL(BL22),.BLN(BLN22),.WL(WL176));
sram_cell_6t_5 inst_cell_176_23 (.BL(BL23),.BLN(BLN23),.WL(WL176));
sram_cell_6t_5 inst_cell_176_24 (.BL(BL24),.BLN(BLN24),.WL(WL176));
sram_cell_6t_5 inst_cell_176_25 (.BL(BL25),.BLN(BLN25),.WL(WL176));
sram_cell_6t_5 inst_cell_176_26 (.BL(BL26),.BLN(BLN26),.WL(WL176));
sram_cell_6t_5 inst_cell_176_27 (.BL(BL27),.BLN(BLN27),.WL(WL176));
sram_cell_6t_5 inst_cell_176_28 (.BL(BL28),.BLN(BLN28),.WL(WL176));
sram_cell_6t_5 inst_cell_176_29 (.BL(BL29),.BLN(BLN29),.WL(WL176));
sram_cell_6t_5 inst_cell_176_30 (.BL(BL30),.BLN(BLN30),.WL(WL176));
sram_cell_6t_5 inst_cell_176_31 (.BL(BL31),.BLN(BLN31),.WL(WL176));
sram_cell_6t_5 inst_cell_176_32 (.BL(BL32),.BLN(BLN32),.WL(WL176));
sram_cell_6t_5 inst_cell_176_33 (.BL(BL33),.BLN(BLN33),.WL(WL176));
sram_cell_6t_5 inst_cell_176_34 (.BL(BL34),.BLN(BLN34),.WL(WL176));
sram_cell_6t_5 inst_cell_176_35 (.BL(BL35),.BLN(BLN35),.WL(WL176));
sram_cell_6t_5 inst_cell_176_36 (.BL(BL36),.BLN(BLN36),.WL(WL176));
sram_cell_6t_5 inst_cell_176_37 (.BL(BL37),.BLN(BLN37),.WL(WL176));
sram_cell_6t_5 inst_cell_176_38 (.BL(BL38),.BLN(BLN38),.WL(WL176));
sram_cell_6t_5 inst_cell_176_39 (.BL(BL39),.BLN(BLN39),.WL(WL176));
sram_cell_6t_5 inst_cell_176_40 (.BL(BL40),.BLN(BLN40),.WL(WL176));
sram_cell_6t_5 inst_cell_176_41 (.BL(BL41),.BLN(BLN41),.WL(WL176));
sram_cell_6t_5 inst_cell_176_42 (.BL(BL42),.BLN(BLN42),.WL(WL176));
sram_cell_6t_5 inst_cell_176_43 (.BL(BL43),.BLN(BLN43),.WL(WL176));
sram_cell_6t_5 inst_cell_176_44 (.BL(BL44),.BLN(BLN44),.WL(WL176));
sram_cell_6t_5 inst_cell_176_45 (.BL(BL45),.BLN(BLN45),.WL(WL176));
sram_cell_6t_5 inst_cell_176_46 (.BL(BL46),.BLN(BLN46),.WL(WL176));
sram_cell_6t_5 inst_cell_176_47 (.BL(BL47),.BLN(BLN47),.WL(WL176));
sram_cell_6t_5 inst_cell_176_48 (.BL(BL48),.BLN(BLN48),.WL(WL176));
sram_cell_6t_5 inst_cell_176_49 (.BL(BL49),.BLN(BLN49),.WL(WL176));
sram_cell_6t_5 inst_cell_176_50 (.BL(BL50),.BLN(BLN50),.WL(WL176));
sram_cell_6t_5 inst_cell_176_51 (.BL(BL51),.BLN(BLN51),.WL(WL176));
sram_cell_6t_5 inst_cell_176_52 (.BL(BL52),.BLN(BLN52),.WL(WL176));
sram_cell_6t_5 inst_cell_176_53 (.BL(BL53),.BLN(BLN53),.WL(WL176));
sram_cell_6t_5 inst_cell_176_54 (.BL(BL54),.BLN(BLN54),.WL(WL176));
sram_cell_6t_5 inst_cell_176_55 (.BL(BL55),.BLN(BLN55),.WL(WL176));
sram_cell_6t_5 inst_cell_176_56 (.BL(BL56),.BLN(BLN56),.WL(WL176));
sram_cell_6t_5 inst_cell_176_57 (.BL(BL57),.BLN(BLN57),.WL(WL176));
sram_cell_6t_5 inst_cell_176_58 (.BL(BL58),.BLN(BLN58),.WL(WL176));
sram_cell_6t_5 inst_cell_176_59 (.BL(BL59),.BLN(BLN59),.WL(WL176));
sram_cell_6t_5 inst_cell_176_60 (.BL(BL60),.BLN(BLN60),.WL(WL176));
sram_cell_6t_5 inst_cell_176_61 (.BL(BL61),.BLN(BLN61),.WL(WL176));
sram_cell_6t_5 inst_cell_176_62 (.BL(BL62),.BLN(BLN62),.WL(WL176));
sram_cell_6t_5 inst_cell_176_63 (.BL(BL63),.BLN(BLN63),.WL(WL176));
sram_cell_6t_5 inst_cell_176_64 (.BL(BL64),.BLN(BLN64),.WL(WL176));
sram_cell_6t_5 inst_cell_176_65 (.BL(BL65),.BLN(BLN65),.WL(WL176));
sram_cell_6t_5 inst_cell_176_66 (.BL(BL66),.BLN(BLN66),.WL(WL176));
sram_cell_6t_5 inst_cell_176_67 (.BL(BL67),.BLN(BLN67),.WL(WL176));
sram_cell_6t_5 inst_cell_176_68 (.BL(BL68),.BLN(BLN68),.WL(WL176));
sram_cell_6t_5 inst_cell_176_69 (.BL(BL69),.BLN(BLN69),.WL(WL176));
sram_cell_6t_5 inst_cell_176_70 (.BL(BL70),.BLN(BLN70),.WL(WL176));
sram_cell_6t_5 inst_cell_176_71 (.BL(BL71),.BLN(BLN71),.WL(WL176));
sram_cell_6t_5 inst_cell_176_72 (.BL(BL72),.BLN(BLN72),.WL(WL176));
sram_cell_6t_5 inst_cell_176_73 (.BL(BL73),.BLN(BLN73),.WL(WL176));
sram_cell_6t_5 inst_cell_176_74 (.BL(BL74),.BLN(BLN74),.WL(WL176));
sram_cell_6t_5 inst_cell_176_75 (.BL(BL75),.BLN(BLN75),.WL(WL176));
sram_cell_6t_5 inst_cell_176_76 (.BL(BL76),.BLN(BLN76),.WL(WL176));
sram_cell_6t_5 inst_cell_176_77 (.BL(BL77),.BLN(BLN77),.WL(WL176));
sram_cell_6t_5 inst_cell_176_78 (.BL(BL78),.BLN(BLN78),.WL(WL176));
sram_cell_6t_5 inst_cell_176_79 (.BL(BL79),.BLN(BLN79),.WL(WL176));
sram_cell_6t_5 inst_cell_176_80 (.BL(BL80),.BLN(BLN80),.WL(WL176));
sram_cell_6t_5 inst_cell_176_81 (.BL(BL81),.BLN(BLN81),.WL(WL176));
sram_cell_6t_5 inst_cell_176_82 (.BL(BL82),.BLN(BLN82),.WL(WL176));
sram_cell_6t_5 inst_cell_176_83 (.BL(BL83),.BLN(BLN83),.WL(WL176));
sram_cell_6t_5 inst_cell_176_84 (.BL(BL84),.BLN(BLN84),.WL(WL176));
sram_cell_6t_5 inst_cell_176_85 (.BL(BL85),.BLN(BLN85),.WL(WL176));
sram_cell_6t_5 inst_cell_176_86 (.BL(BL86),.BLN(BLN86),.WL(WL176));
sram_cell_6t_5 inst_cell_176_87 (.BL(BL87),.BLN(BLN87),.WL(WL176));
sram_cell_6t_5 inst_cell_176_88 (.BL(BL88),.BLN(BLN88),.WL(WL176));
sram_cell_6t_5 inst_cell_176_89 (.BL(BL89),.BLN(BLN89),.WL(WL176));
sram_cell_6t_5 inst_cell_176_90 (.BL(BL90),.BLN(BLN90),.WL(WL176));
sram_cell_6t_5 inst_cell_176_91 (.BL(BL91),.BLN(BLN91),.WL(WL176));
sram_cell_6t_5 inst_cell_176_92 (.BL(BL92),.BLN(BLN92),.WL(WL176));
sram_cell_6t_5 inst_cell_176_93 (.BL(BL93),.BLN(BLN93),.WL(WL176));
sram_cell_6t_5 inst_cell_176_94 (.BL(BL94),.BLN(BLN94),.WL(WL176));
sram_cell_6t_5 inst_cell_176_95 (.BL(BL95),.BLN(BLN95),.WL(WL176));
sram_cell_6t_5 inst_cell_176_96 (.BL(BL96),.BLN(BLN96),.WL(WL176));
sram_cell_6t_5 inst_cell_176_97 (.BL(BL97),.BLN(BLN97),.WL(WL176));
sram_cell_6t_5 inst_cell_176_98 (.BL(BL98),.BLN(BLN98),.WL(WL176));
sram_cell_6t_5 inst_cell_176_99 (.BL(BL99),.BLN(BLN99),.WL(WL176));
sram_cell_6t_5 inst_cell_176_100 (.BL(BL100),.BLN(BLN100),.WL(WL176));
sram_cell_6t_5 inst_cell_176_101 (.BL(BL101),.BLN(BLN101),.WL(WL176));
sram_cell_6t_5 inst_cell_176_102 (.BL(BL102),.BLN(BLN102),.WL(WL176));
sram_cell_6t_5 inst_cell_176_103 (.BL(BL103),.BLN(BLN103),.WL(WL176));
sram_cell_6t_5 inst_cell_176_104 (.BL(BL104),.BLN(BLN104),.WL(WL176));
sram_cell_6t_5 inst_cell_176_105 (.BL(BL105),.BLN(BLN105),.WL(WL176));
sram_cell_6t_5 inst_cell_176_106 (.BL(BL106),.BLN(BLN106),.WL(WL176));
sram_cell_6t_5 inst_cell_176_107 (.BL(BL107),.BLN(BLN107),.WL(WL176));
sram_cell_6t_5 inst_cell_176_108 (.BL(BL108),.BLN(BLN108),.WL(WL176));
sram_cell_6t_5 inst_cell_176_109 (.BL(BL109),.BLN(BLN109),.WL(WL176));
sram_cell_6t_5 inst_cell_176_110 (.BL(BL110),.BLN(BLN110),.WL(WL176));
sram_cell_6t_5 inst_cell_176_111 (.BL(BL111),.BLN(BLN111),.WL(WL176));
sram_cell_6t_5 inst_cell_176_112 (.BL(BL112),.BLN(BLN112),.WL(WL176));
sram_cell_6t_5 inst_cell_176_113 (.BL(BL113),.BLN(BLN113),.WL(WL176));
sram_cell_6t_5 inst_cell_176_114 (.BL(BL114),.BLN(BLN114),.WL(WL176));
sram_cell_6t_5 inst_cell_176_115 (.BL(BL115),.BLN(BLN115),.WL(WL176));
sram_cell_6t_5 inst_cell_176_116 (.BL(BL116),.BLN(BLN116),.WL(WL176));
sram_cell_6t_5 inst_cell_176_117 (.BL(BL117),.BLN(BLN117),.WL(WL176));
sram_cell_6t_5 inst_cell_176_118 (.BL(BL118),.BLN(BLN118),.WL(WL176));
sram_cell_6t_5 inst_cell_176_119 (.BL(BL119),.BLN(BLN119),.WL(WL176));
sram_cell_6t_5 inst_cell_176_120 (.BL(BL120),.BLN(BLN120),.WL(WL176));
sram_cell_6t_5 inst_cell_176_121 (.BL(BL121),.BLN(BLN121),.WL(WL176));
sram_cell_6t_5 inst_cell_176_122 (.BL(BL122),.BLN(BLN122),.WL(WL176));
sram_cell_6t_5 inst_cell_176_123 (.BL(BL123),.BLN(BLN123),.WL(WL176));
sram_cell_6t_5 inst_cell_176_124 (.BL(BL124),.BLN(BLN124),.WL(WL176));
sram_cell_6t_5 inst_cell_176_125 (.BL(BL125),.BLN(BLN125),.WL(WL176));
sram_cell_6t_5 inst_cell_176_126 (.BL(BL126),.BLN(BLN126),.WL(WL176));
sram_cell_6t_5 inst_cell_176_127 (.BL(BL127),.BLN(BLN127),.WL(WL176));
sram_cell_6t_5 inst_cell_177_0 (.BL(BL0),.BLN(BLN0),.WL(WL177));
sram_cell_6t_5 inst_cell_177_1 (.BL(BL1),.BLN(BLN1),.WL(WL177));
sram_cell_6t_5 inst_cell_177_2 (.BL(BL2),.BLN(BLN2),.WL(WL177));
sram_cell_6t_5 inst_cell_177_3 (.BL(BL3),.BLN(BLN3),.WL(WL177));
sram_cell_6t_5 inst_cell_177_4 (.BL(BL4),.BLN(BLN4),.WL(WL177));
sram_cell_6t_5 inst_cell_177_5 (.BL(BL5),.BLN(BLN5),.WL(WL177));
sram_cell_6t_5 inst_cell_177_6 (.BL(BL6),.BLN(BLN6),.WL(WL177));
sram_cell_6t_5 inst_cell_177_7 (.BL(BL7),.BLN(BLN7),.WL(WL177));
sram_cell_6t_5 inst_cell_177_8 (.BL(BL8),.BLN(BLN8),.WL(WL177));
sram_cell_6t_5 inst_cell_177_9 (.BL(BL9),.BLN(BLN9),.WL(WL177));
sram_cell_6t_5 inst_cell_177_10 (.BL(BL10),.BLN(BLN10),.WL(WL177));
sram_cell_6t_5 inst_cell_177_11 (.BL(BL11),.BLN(BLN11),.WL(WL177));
sram_cell_6t_5 inst_cell_177_12 (.BL(BL12),.BLN(BLN12),.WL(WL177));
sram_cell_6t_5 inst_cell_177_13 (.BL(BL13),.BLN(BLN13),.WL(WL177));
sram_cell_6t_5 inst_cell_177_14 (.BL(BL14),.BLN(BLN14),.WL(WL177));
sram_cell_6t_5 inst_cell_177_15 (.BL(BL15),.BLN(BLN15),.WL(WL177));
sram_cell_6t_5 inst_cell_177_16 (.BL(BL16),.BLN(BLN16),.WL(WL177));
sram_cell_6t_5 inst_cell_177_17 (.BL(BL17),.BLN(BLN17),.WL(WL177));
sram_cell_6t_5 inst_cell_177_18 (.BL(BL18),.BLN(BLN18),.WL(WL177));
sram_cell_6t_5 inst_cell_177_19 (.BL(BL19),.BLN(BLN19),.WL(WL177));
sram_cell_6t_5 inst_cell_177_20 (.BL(BL20),.BLN(BLN20),.WL(WL177));
sram_cell_6t_5 inst_cell_177_21 (.BL(BL21),.BLN(BLN21),.WL(WL177));
sram_cell_6t_5 inst_cell_177_22 (.BL(BL22),.BLN(BLN22),.WL(WL177));
sram_cell_6t_5 inst_cell_177_23 (.BL(BL23),.BLN(BLN23),.WL(WL177));
sram_cell_6t_5 inst_cell_177_24 (.BL(BL24),.BLN(BLN24),.WL(WL177));
sram_cell_6t_5 inst_cell_177_25 (.BL(BL25),.BLN(BLN25),.WL(WL177));
sram_cell_6t_5 inst_cell_177_26 (.BL(BL26),.BLN(BLN26),.WL(WL177));
sram_cell_6t_5 inst_cell_177_27 (.BL(BL27),.BLN(BLN27),.WL(WL177));
sram_cell_6t_5 inst_cell_177_28 (.BL(BL28),.BLN(BLN28),.WL(WL177));
sram_cell_6t_5 inst_cell_177_29 (.BL(BL29),.BLN(BLN29),.WL(WL177));
sram_cell_6t_5 inst_cell_177_30 (.BL(BL30),.BLN(BLN30),.WL(WL177));
sram_cell_6t_5 inst_cell_177_31 (.BL(BL31),.BLN(BLN31),.WL(WL177));
sram_cell_6t_5 inst_cell_177_32 (.BL(BL32),.BLN(BLN32),.WL(WL177));
sram_cell_6t_5 inst_cell_177_33 (.BL(BL33),.BLN(BLN33),.WL(WL177));
sram_cell_6t_5 inst_cell_177_34 (.BL(BL34),.BLN(BLN34),.WL(WL177));
sram_cell_6t_5 inst_cell_177_35 (.BL(BL35),.BLN(BLN35),.WL(WL177));
sram_cell_6t_5 inst_cell_177_36 (.BL(BL36),.BLN(BLN36),.WL(WL177));
sram_cell_6t_5 inst_cell_177_37 (.BL(BL37),.BLN(BLN37),.WL(WL177));
sram_cell_6t_5 inst_cell_177_38 (.BL(BL38),.BLN(BLN38),.WL(WL177));
sram_cell_6t_5 inst_cell_177_39 (.BL(BL39),.BLN(BLN39),.WL(WL177));
sram_cell_6t_5 inst_cell_177_40 (.BL(BL40),.BLN(BLN40),.WL(WL177));
sram_cell_6t_5 inst_cell_177_41 (.BL(BL41),.BLN(BLN41),.WL(WL177));
sram_cell_6t_5 inst_cell_177_42 (.BL(BL42),.BLN(BLN42),.WL(WL177));
sram_cell_6t_5 inst_cell_177_43 (.BL(BL43),.BLN(BLN43),.WL(WL177));
sram_cell_6t_5 inst_cell_177_44 (.BL(BL44),.BLN(BLN44),.WL(WL177));
sram_cell_6t_5 inst_cell_177_45 (.BL(BL45),.BLN(BLN45),.WL(WL177));
sram_cell_6t_5 inst_cell_177_46 (.BL(BL46),.BLN(BLN46),.WL(WL177));
sram_cell_6t_5 inst_cell_177_47 (.BL(BL47),.BLN(BLN47),.WL(WL177));
sram_cell_6t_5 inst_cell_177_48 (.BL(BL48),.BLN(BLN48),.WL(WL177));
sram_cell_6t_5 inst_cell_177_49 (.BL(BL49),.BLN(BLN49),.WL(WL177));
sram_cell_6t_5 inst_cell_177_50 (.BL(BL50),.BLN(BLN50),.WL(WL177));
sram_cell_6t_5 inst_cell_177_51 (.BL(BL51),.BLN(BLN51),.WL(WL177));
sram_cell_6t_5 inst_cell_177_52 (.BL(BL52),.BLN(BLN52),.WL(WL177));
sram_cell_6t_5 inst_cell_177_53 (.BL(BL53),.BLN(BLN53),.WL(WL177));
sram_cell_6t_5 inst_cell_177_54 (.BL(BL54),.BLN(BLN54),.WL(WL177));
sram_cell_6t_5 inst_cell_177_55 (.BL(BL55),.BLN(BLN55),.WL(WL177));
sram_cell_6t_5 inst_cell_177_56 (.BL(BL56),.BLN(BLN56),.WL(WL177));
sram_cell_6t_5 inst_cell_177_57 (.BL(BL57),.BLN(BLN57),.WL(WL177));
sram_cell_6t_5 inst_cell_177_58 (.BL(BL58),.BLN(BLN58),.WL(WL177));
sram_cell_6t_5 inst_cell_177_59 (.BL(BL59),.BLN(BLN59),.WL(WL177));
sram_cell_6t_5 inst_cell_177_60 (.BL(BL60),.BLN(BLN60),.WL(WL177));
sram_cell_6t_5 inst_cell_177_61 (.BL(BL61),.BLN(BLN61),.WL(WL177));
sram_cell_6t_5 inst_cell_177_62 (.BL(BL62),.BLN(BLN62),.WL(WL177));
sram_cell_6t_5 inst_cell_177_63 (.BL(BL63),.BLN(BLN63),.WL(WL177));
sram_cell_6t_5 inst_cell_177_64 (.BL(BL64),.BLN(BLN64),.WL(WL177));
sram_cell_6t_5 inst_cell_177_65 (.BL(BL65),.BLN(BLN65),.WL(WL177));
sram_cell_6t_5 inst_cell_177_66 (.BL(BL66),.BLN(BLN66),.WL(WL177));
sram_cell_6t_5 inst_cell_177_67 (.BL(BL67),.BLN(BLN67),.WL(WL177));
sram_cell_6t_5 inst_cell_177_68 (.BL(BL68),.BLN(BLN68),.WL(WL177));
sram_cell_6t_5 inst_cell_177_69 (.BL(BL69),.BLN(BLN69),.WL(WL177));
sram_cell_6t_5 inst_cell_177_70 (.BL(BL70),.BLN(BLN70),.WL(WL177));
sram_cell_6t_5 inst_cell_177_71 (.BL(BL71),.BLN(BLN71),.WL(WL177));
sram_cell_6t_5 inst_cell_177_72 (.BL(BL72),.BLN(BLN72),.WL(WL177));
sram_cell_6t_5 inst_cell_177_73 (.BL(BL73),.BLN(BLN73),.WL(WL177));
sram_cell_6t_5 inst_cell_177_74 (.BL(BL74),.BLN(BLN74),.WL(WL177));
sram_cell_6t_5 inst_cell_177_75 (.BL(BL75),.BLN(BLN75),.WL(WL177));
sram_cell_6t_5 inst_cell_177_76 (.BL(BL76),.BLN(BLN76),.WL(WL177));
sram_cell_6t_5 inst_cell_177_77 (.BL(BL77),.BLN(BLN77),.WL(WL177));
sram_cell_6t_5 inst_cell_177_78 (.BL(BL78),.BLN(BLN78),.WL(WL177));
sram_cell_6t_5 inst_cell_177_79 (.BL(BL79),.BLN(BLN79),.WL(WL177));
sram_cell_6t_5 inst_cell_177_80 (.BL(BL80),.BLN(BLN80),.WL(WL177));
sram_cell_6t_5 inst_cell_177_81 (.BL(BL81),.BLN(BLN81),.WL(WL177));
sram_cell_6t_5 inst_cell_177_82 (.BL(BL82),.BLN(BLN82),.WL(WL177));
sram_cell_6t_5 inst_cell_177_83 (.BL(BL83),.BLN(BLN83),.WL(WL177));
sram_cell_6t_5 inst_cell_177_84 (.BL(BL84),.BLN(BLN84),.WL(WL177));
sram_cell_6t_5 inst_cell_177_85 (.BL(BL85),.BLN(BLN85),.WL(WL177));
sram_cell_6t_5 inst_cell_177_86 (.BL(BL86),.BLN(BLN86),.WL(WL177));
sram_cell_6t_5 inst_cell_177_87 (.BL(BL87),.BLN(BLN87),.WL(WL177));
sram_cell_6t_5 inst_cell_177_88 (.BL(BL88),.BLN(BLN88),.WL(WL177));
sram_cell_6t_5 inst_cell_177_89 (.BL(BL89),.BLN(BLN89),.WL(WL177));
sram_cell_6t_5 inst_cell_177_90 (.BL(BL90),.BLN(BLN90),.WL(WL177));
sram_cell_6t_5 inst_cell_177_91 (.BL(BL91),.BLN(BLN91),.WL(WL177));
sram_cell_6t_5 inst_cell_177_92 (.BL(BL92),.BLN(BLN92),.WL(WL177));
sram_cell_6t_5 inst_cell_177_93 (.BL(BL93),.BLN(BLN93),.WL(WL177));
sram_cell_6t_5 inst_cell_177_94 (.BL(BL94),.BLN(BLN94),.WL(WL177));
sram_cell_6t_5 inst_cell_177_95 (.BL(BL95),.BLN(BLN95),.WL(WL177));
sram_cell_6t_5 inst_cell_177_96 (.BL(BL96),.BLN(BLN96),.WL(WL177));
sram_cell_6t_5 inst_cell_177_97 (.BL(BL97),.BLN(BLN97),.WL(WL177));
sram_cell_6t_5 inst_cell_177_98 (.BL(BL98),.BLN(BLN98),.WL(WL177));
sram_cell_6t_5 inst_cell_177_99 (.BL(BL99),.BLN(BLN99),.WL(WL177));
sram_cell_6t_5 inst_cell_177_100 (.BL(BL100),.BLN(BLN100),.WL(WL177));
sram_cell_6t_5 inst_cell_177_101 (.BL(BL101),.BLN(BLN101),.WL(WL177));
sram_cell_6t_5 inst_cell_177_102 (.BL(BL102),.BLN(BLN102),.WL(WL177));
sram_cell_6t_5 inst_cell_177_103 (.BL(BL103),.BLN(BLN103),.WL(WL177));
sram_cell_6t_5 inst_cell_177_104 (.BL(BL104),.BLN(BLN104),.WL(WL177));
sram_cell_6t_5 inst_cell_177_105 (.BL(BL105),.BLN(BLN105),.WL(WL177));
sram_cell_6t_5 inst_cell_177_106 (.BL(BL106),.BLN(BLN106),.WL(WL177));
sram_cell_6t_5 inst_cell_177_107 (.BL(BL107),.BLN(BLN107),.WL(WL177));
sram_cell_6t_5 inst_cell_177_108 (.BL(BL108),.BLN(BLN108),.WL(WL177));
sram_cell_6t_5 inst_cell_177_109 (.BL(BL109),.BLN(BLN109),.WL(WL177));
sram_cell_6t_5 inst_cell_177_110 (.BL(BL110),.BLN(BLN110),.WL(WL177));
sram_cell_6t_5 inst_cell_177_111 (.BL(BL111),.BLN(BLN111),.WL(WL177));
sram_cell_6t_5 inst_cell_177_112 (.BL(BL112),.BLN(BLN112),.WL(WL177));
sram_cell_6t_5 inst_cell_177_113 (.BL(BL113),.BLN(BLN113),.WL(WL177));
sram_cell_6t_5 inst_cell_177_114 (.BL(BL114),.BLN(BLN114),.WL(WL177));
sram_cell_6t_5 inst_cell_177_115 (.BL(BL115),.BLN(BLN115),.WL(WL177));
sram_cell_6t_5 inst_cell_177_116 (.BL(BL116),.BLN(BLN116),.WL(WL177));
sram_cell_6t_5 inst_cell_177_117 (.BL(BL117),.BLN(BLN117),.WL(WL177));
sram_cell_6t_5 inst_cell_177_118 (.BL(BL118),.BLN(BLN118),.WL(WL177));
sram_cell_6t_5 inst_cell_177_119 (.BL(BL119),.BLN(BLN119),.WL(WL177));
sram_cell_6t_5 inst_cell_177_120 (.BL(BL120),.BLN(BLN120),.WL(WL177));
sram_cell_6t_5 inst_cell_177_121 (.BL(BL121),.BLN(BLN121),.WL(WL177));
sram_cell_6t_5 inst_cell_177_122 (.BL(BL122),.BLN(BLN122),.WL(WL177));
sram_cell_6t_5 inst_cell_177_123 (.BL(BL123),.BLN(BLN123),.WL(WL177));
sram_cell_6t_5 inst_cell_177_124 (.BL(BL124),.BLN(BLN124),.WL(WL177));
sram_cell_6t_5 inst_cell_177_125 (.BL(BL125),.BLN(BLN125),.WL(WL177));
sram_cell_6t_5 inst_cell_177_126 (.BL(BL126),.BLN(BLN126),.WL(WL177));
sram_cell_6t_5 inst_cell_177_127 (.BL(BL127),.BLN(BLN127),.WL(WL177));
sram_cell_6t_5 inst_cell_178_0 (.BL(BL0),.BLN(BLN0),.WL(WL178));
sram_cell_6t_5 inst_cell_178_1 (.BL(BL1),.BLN(BLN1),.WL(WL178));
sram_cell_6t_5 inst_cell_178_2 (.BL(BL2),.BLN(BLN2),.WL(WL178));
sram_cell_6t_5 inst_cell_178_3 (.BL(BL3),.BLN(BLN3),.WL(WL178));
sram_cell_6t_5 inst_cell_178_4 (.BL(BL4),.BLN(BLN4),.WL(WL178));
sram_cell_6t_5 inst_cell_178_5 (.BL(BL5),.BLN(BLN5),.WL(WL178));
sram_cell_6t_5 inst_cell_178_6 (.BL(BL6),.BLN(BLN6),.WL(WL178));
sram_cell_6t_5 inst_cell_178_7 (.BL(BL7),.BLN(BLN7),.WL(WL178));
sram_cell_6t_5 inst_cell_178_8 (.BL(BL8),.BLN(BLN8),.WL(WL178));
sram_cell_6t_5 inst_cell_178_9 (.BL(BL9),.BLN(BLN9),.WL(WL178));
sram_cell_6t_5 inst_cell_178_10 (.BL(BL10),.BLN(BLN10),.WL(WL178));
sram_cell_6t_5 inst_cell_178_11 (.BL(BL11),.BLN(BLN11),.WL(WL178));
sram_cell_6t_5 inst_cell_178_12 (.BL(BL12),.BLN(BLN12),.WL(WL178));
sram_cell_6t_5 inst_cell_178_13 (.BL(BL13),.BLN(BLN13),.WL(WL178));
sram_cell_6t_5 inst_cell_178_14 (.BL(BL14),.BLN(BLN14),.WL(WL178));
sram_cell_6t_5 inst_cell_178_15 (.BL(BL15),.BLN(BLN15),.WL(WL178));
sram_cell_6t_5 inst_cell_178_16 (.BL(BL16),.BLN(BLN16),.WL(WL178));
sram_cell_6t_5 inst_cell_178_17 (.BL(BL17),.BLN(BLN17),.WL(WL178));
sram_cell_6t_5 inst_cell_178_18 (.BL(BL18),.BLN(BLN18),.WL(WL178));
sram_cell_6t_5 inst_cell_178_19 (.BL(BL19),.BLN(BLN19),.WL(WL178));
sram_cell_6t_5 inst_cell_178_20 (.BL(BL20),.BLN(BLN20),.WL(WL178));
sram_cell_6t_5 inst_cell_178_21 (.BL(BL21),.BLN(BLN21),.WL(WL178));
sram_cell_6t_5 inst_cell_178_22 (.BL(BL22),.BLN(BLN22),.WL(WL178));
sram_cell_6t_5 inst_cell_178_23 (.BL(BL23),.BLN(BLN23),.WL(WL178));
sram_cell_6t_5 inst_cell_178_24 (.BL(BL24),.BLN(BLN24),.WL(WL178));
sram_cell_6t_5 inst_cell_178_25 (.BL(BL25),.BLN(BLN25),.WL(WL178));
sram_cell_6t_5 inst_cell_178_26 (.BL(BL26),.BLN(BLN26),.WL(WL178));
sram_cell_6t_5 inst_cell_178_27 (.BL(BL27),.BLN(BLN27),.WL(WL178));
sram_cell_6t_5 inst_cell_178_28 (.BL(BL28),.BLN(BLN28),.WL(WL178));
sram_cell_6t_5 inst_cell_178_29 (.BL(BL29),.BLN(BLN29),.WL(WL178));
sram_cell_6t_5 inst_cell_178_30 (.BL(BL30),.BLN(BLN30),.WL(WL178));
sram_cell_6t_5 inst_cell_178_31 (.BL(BL31),.BLN(BLN31),.WL(WL178));
sram_cell_6t_5 inst_cell_178_32 (.BL(BL32),.BLN(BLN32),.WL(WL178));
sram_cell_6t_5 inst_cell_178_33 (.BL(BL33),.BLN(BLN33),.WL(WL178));
sram_cell_6t_5 inst_cell_178_34 (.BL(BL34),.BLN(BLN34),.WL(WL178));
sram_cell_6t_5 inst_cell_178_35 (.BL(BL35),.BLN(BLN35),.WL(WL178));
sram_cell_6t_5 inst_cell_178_36 (.BL(BL36),.BLN(BLN36),.WL(WL178));
sram_cell_6t_5 inst_cell_178_37 (.BL(BL37),.BLN(BLN37),.WL(WL178));
sram_cell_6t_5 inst_cell_178_38 (.BL(BL38),.BLN(BLN38),.WL(WL178));
sram_cell_6t_5 inst_cell_178_39 (.BL(BL39),.BLN(BLN39),.WL(WL178));
sram_cell_6t_5 inst_cell_178_40 (.BL(BL40),.BLN(BLN40),.WL(WL178));
sram_cell_6t_5 inst_cell_178_41 (.BL(BL41),.BLN(BLN41),.WL(WL178));
sram_cell_6t_5 inst_cell_178_42 (.BL(BL42),.BLN(BLN42),.WL(WL178));
sram_cell_6t_5 inst_cell_178_43 (.BL(BL43),.BLN(BLN43),.WL(WL178));
sram_cell_6t_5 inst_cell_178_44 (.BL(BL44),.BLN(BLN44),.WL(WL178));
sram_cell_6t_5 inst_cell_178_45 (.BL(BL45),.BLN(BLN45),.WL(WL178));
sram_cell_6t_5 inst_cell_178_46 (.BL(BL46),.BLN(BLN46),.WL(WL178));
sram_cell_6t_5 inst_cell_178_47 (.BL(BL47),.BLN(BLN47),.WL(WL178));
sram_cell_6t_5 inst_cell_178_48 (.BL(BL48),.BLN(BLN48),.WL(WL178));
sram_cell_6t_5 inst_cell_178_49 (.BL(BL49),.BLN(BLN49),.WL(WL178));
sram_cell_6t_5 inst_cell_178_50 (.BL(BL50),.BLN(BLN50),.WL(WL178));
sram_cell_6t_5 inst_cell_178_51 (.BL(BL51),.BLN(BLN51),.WL(WL178));
sram_cell_6t_5 inst_cell_178_52 (.BL(BL52),.BLN(BLN52),.WL(WL178));
sram_cell_6t_5 inst_cell_178_53 (.BL(BL53),.BLN(BLN53),.WL(WL178));
sram_cell_6t_5 inst_cell_178_54 (.BL(BL54),.BLN(BLN54),.WL(WL178));
sram_cell_6t_5 inst_cell_178_55 (.BL(BL55),.BLN(BLN55),.WL(WL178));
sram_cell_6t_5 inst_cell_178_56 (.BL(BL56),.BLN(BLN56),.WL(WL178));
sram_cell_6t_5 inst_cell_178_57 (.BL(BL57),.BLN(BLN57),.WL(WL178));
sram_cell_6t_5 inst_cell_178_58 (.BL(BL58),.BLN(BLN58),.WL(WL178));
sram_cell_6t_5 inst_cell_178_59 (.BL(BL59),.BLN(BLN59),.WL(WL178));
sram_cell_6t_5 inst_cell_178_60 (.BL(BL60),.BLN(BLN60),.WL(WL178));
sram_cell_6t_5 inst_cell_178_61 (.BL(BL61),.BLN(BLN61),.WL(WL178));
sram_cell_6t_5 inst_cell_178_62 (.BL(BL62),.BLN(BLN62),.WL(WL178));
sram_cell_6t_5 inst_cell_178_63 (.BL(BL63),.BLN(BLN63),.WL(WL178));
sram_cell_6t_5 inst_cell_178_64 (.BL(BL64),.BLN(BLN64),.WL(WL178));
sram_cell_6t_5 inst_cell_178_65 (.BL(BL65),.BLN(BLN65),.WL(WL178));
sram_cell_6t_5 inst_cell_178_66 (.BL(BL66),.BLN(BLN66),.WL(WL178));
sram_cell_6t_5 inst_cell_178_67 (.BL(BL67),.BLN(BLN67),.WL(WL178));
sram_cell_6t_5 inst_cell_178_68 (.BL(BL68),.BLN(BLN68),.WL(WL178));
sram_cell_6t_5 inst_cell_178_69 (.BL(BL69),.BLN(BLN69),.WL(WL178));
sram_cell_6t_5 inst_cell_178_70 (.BL(BL70),.BLN(BLN70),.WL(WL178));
sram_cell_6t_5 inst_cell_178_71 (.BL(BL71),.BLN(BLN71),.WL(WL178));
sram_cell_6t_5 inst_cell_178_72 (.BL(BL72),.BLN(BLN72),.WL(WL178));
sram_cell_6t_5 inst_cell_178_73 (.BL(BL73),.BLN(BLN73),.WL(WL178));
sram_cell_6t_5 inst_cell_178_74 (.BL(BL74),.BLN(BLN74),.WL(WL178));
sram_cell_6t_5 inst_cell_178_75 (.BL(BL75),.BLN(BLN75),.WL(WL178));
sram_cell_6t_5 inst_cell_178_76 (.BL(BL76),.BLN(BLN76),.WL(WL178));
sram_cell_6t_5 inst_cell_178_77 (.BL(BL77),.BLN(BLN77),.WL(WL178));
sram_cell_6t_5 inst_cell_178_78 (.BL(BL78),.BLN(BLN78),.WL(WL178));
sram_cell_6t_5 inst_cell_178_79 (.BL(BL79),.BLN(BLN79),.WL(WL178));
sram_cell_6t_5 inst_cell_178_80 (.BL(BL80),.BLN(BLN80),.WL(WL178));
sram_cell_6t_5 inst_cell_178_81 (.BL(BL81),.BLN(BLN81),.WL(WL178));
sram_cell_6t_5 inst_cell_178_82 (.BL(BL82),.BLN(BLN82),.WL(WL178));
sram_cell_6t_5 inst_cell_178_83 (.BL(BL83),.BLN(BLN83),.WL(WL178));
sram_cell_6t_5 inst_cell_178_84 (.BL(BL84),.BLN(BLN84),.WL(WL178));
sram_cell_6t_5 inst_cell_178_85 (.BL(BL85),.BLN(BLN85),.WL(WL178));
sram_cell_6t_5 inst_cell_178_86 (.BL(BL86),.BLN(BLN86),.WL(WL178));
sram_cell_6t_5 inst_cell_178_87 (.BL(BL87),.BLN(BLN87),.WL(WL178));
sram_cell_6t_5 inst_cell_178_88 (.BL(BL88),.BLN(BLN88),.WL(WL178));
sram_cell_6t_5 inst_cell_178_89 (.BL(BL89),.BLN(BLN89),.WL(WL178));
sram_cell_6t_5 inst_cell_178_90 (.BL(BL90),.BLN(BLN90),.WL(WL178));
sram_cell_6t_5 inst_cell_178_91 (.BL(BL91),.BLN(BLN91),.WL(WL178));
sram_cell_6t_5 inst_cell_178_92 (.BL(BL92),.BLN(BLN92),.WL(WL178));
sram_cell_6t_5 inst_cell_178_93 (.BL(BL93),.BLN(BLN93),.WL(WL178));
sram_cell_6t_5 inst_cell_178_94 (.BL(BL94),.BLN(BLN94),.WL(WL178));
sram_cell_6t_5 inst_cell_178_95 (.BL(BL95),.BLN(BLN95),.WL(WL178));
sram_cell_6t_5 inst_cell_178_96 (.BL(BL96),.BLN(BLN96),.WL(WL178));
sram_cell_6t_5 inst_cell_178_97 (.BL(BL97),.BLN(BLN97),.WL(WL178));
sram_cell_6t_5 inst_cell_178_98 (.BL(BL98),.BLN(BLN98),.WL(WL178));
sram_cell_6t_5 inst_cell_178_99 (.BL(BL99),.BLN(BLN99),.WL(WL178));
sram_cell_6t_5 inst_cell_178_100 (.BL(BL100),.BLN(BLN100),.WL(WL178));
sram_cell_6t_5 inst_cell_178_101 (.BL(BL101),.BLN(BLN101),.WL(WL178));
sram_cell_6t_5 inst_cell_178_102 (.BL(BL102),.BLN(BLN102),.WL(WL178));
sram_cell_6t_5 inst_cell_178_103 (.BL(BL103),.BLN(BLN103),.WL(WL178));
sram_cell_6t_5 inst_cell_178_104 (.BL(BL104),.BLN(BLN104),.WL(WL178));
sram_cell_6t_5 inst_cell_178_105 (.BL(BL105),.BLN(BLN105),.WL(WL178));
sram_cell_6t_5 inst_cell_178_106 (.BL(BL106),.BLN(BLN106),.WL(WL178));
sram_cell_6t_5 inst_cell_178_107 (.BL(BL107),.BLN(BLN107),.WL(WL178));
sram_cell_6t_5 inst_cell_178_108 (.BL(BL108),.BLN(BLN108),.WL(WL178));
sram_cell_6t_5 inst_cell_178_109 (.BL(BL109),.BLN(BLN109),.WL(WL178));
sram_cell_6t_5 inst_cell_178_110 (.BL(BL110),.BLN(BLN110),.WL(WL178));
sram_cell_6t_5 inst_cell_178_111 (.BL(BL111),.BLN(BLN111),.WL(WL178));
sram_cell_6t_5 inst_cell_178_112 (.BL(BL112),.BLN(BLN112),.WL(WL178));
sram_cell_6t_5 inst_cell_178_113 (.BL(BL113),.BLN(BLN113),.WL(WL178));
sram_cell_6t_5 inst_cell_178_114 (.BL(BL114),.BLN(BLN114),.WL(WL178));
sram_cell_6t_5 inst_cell_178_115 (.BL(BL115),.BLN(BLN115),.WL(WL178));
sram_cell_6t_5 inst_cell_178_116 (.BL(BL116),.BLN(BLN116),.WL(WL178));
sram_cell_6t_5 inst_cell_178_117 (.BL(BL117),.BLN(BLN117),.WL(WL178));
sram_cell_6t_5 inst_cell_178_118 (.BL(BL118),.BLN(BLN118),.WL(WL178));
sram_cell_6t_5 inst_cell_178_119 (.BL(BL119),.BLN(BLN119),.WL(WL178));
sram_cell_6t_5 inst_cell_178_120 (.BL(BL120),.BLN(BLN120),.WL(WL178));
sram_cell_6t_5 inst_cell_178_121 (.BL(BL121),.BLN(BLN121),.WL(WL178));
sram_cell_6t_5 inst_cell_178_122 (.BL(BL122),.BLN(BLN122),.WL(WL178));
sram_cell_6t_5 inst_cell_178_123 (.BL(BL123),.BLN(BLN123),.WL(WL178));
sram_cell_6t_5 inst_cell_178_124 (.BL(BL124),.BLN(BLN124),.WL(WL178));
sram_cell_6t_5 inst_cell_178_125 (.BL(BL125),.BLN(BLN125),.WL(WL178));
sram_cell_6t_5 inst_cell_178_126 (.BL(BL126),.BLN(BLN126),.WL(WL178));
sram_cell_6t_5 inst_cell_178_127 (.BL(BL127),.BLN(BLN127),.WL(WL178));
sram_cell_6t_5 inst_cell_179_0 (.BL(BL0),.BLN(BLN0),.WL(WL179));
sram_cell_6t_5 inst_cell_179_1 (.BL(BL1),.BLN(BLN1),.WL(WL179));
sram_cell_6t_5 inst_cell_179_2 (.BL(BL2),.BLN(BLN2),.WL(WL179));
sram_cell_6t_5 inst_cell_179_3 (.BL(BL3),.BLN(BLN3),.WL(WL179));
sram_cell_6t_5 inst_cell_179_4 (.BL(BL4),.BLN(BLN4),.WL(WL179));
sram_cell_6t_5 inst_cell_179_5 (.BL(BL5),.BLN(BLN5),.WL(WL179));
sram_cell_6t_5 inst_cell_179_6 (.BL(BL6),.BLN(BLN6),.WL(WL179));
sram_cell_6t_5 inst_cell_179_7 (.BL(BL7),.BLN(BLN7),.WL(WL179));
sram_cell_6t_5 inst_cell_179_8 (.BL(BL8),.BLN(BLN8),.WL(WL179));
sram_cell_6t_5 inst_cell_179_9 (.BL(BL9),.BLN(BLN9),.WL(WL179));
sram_cell_6t_5 inst_cell_179_10 (.BL(BL10),.BLN(BLN10),.WL(WL179));
sram_cell_6t_5 inst_cell_179_11 (.BL(BL11),.BLN(BLN11),.WL(WL179));
sram_cell_6t_5 inst_cell_179_12 (.BL(BL12),.BLN(BLN12),.WL(WL179));
sram_cell_6t_5 inst_cell_179_13 (.BL(BL13),.BLN(BLN13),.WL(WL179));
sram_cell_6t_5 inst_cell_179_14 (.BL(BL14),.BLN(BLN14),.WL(WL179));
sram_cell_6t_5 inst_cell_179_15 (.BL(BL15),.BLN(BLN15),.WL(WL179));
sram_cell_6t_5 inst_cell_179_16 (.BL(BL16),.BLN(BLN16),.WL(WL179));
sram_cell_6t_5 inst_cell_179_17 (.BL(BL17),.BLN(BLN17),.WL(WL179));
sram_cell_6t_5 inst_cell_179_18 (.BL(BL18),.BLN(BLN18),.WL(WL179));
sram_cell_6t_5 inst_cell_179_19 (.BL(BL19),.BLN(BLN19),.WL(WL179));
sram_cell_6t_5 inst_cell_179_20 (.BL(BL20),.BLN(BLN20),.WL(WL179));
sram_cell_6t_5 inst_cell_179_21 (.BL(BL21),.BLN(BLN21),.WL(WL179));
sram_cell_6t_5 inst_cell_179_22 (.BL(BL22),.BLN(BLN22),.WL(WL179));
sram_cell_6t_5 inst_cell_179_23 (.BL(BL23),.BLN(BLN23),.WL(WL179));
sram_cell_6t_5 inst_cell_179_24 (.BL(BL24),.BLN(BLN24),.WL(WL179));
sram_cell_6t_5 inst_cell_179_25 (.BL(BL25),.BLN(BLN25),.WL(WL179));
sram_cell_6t_5 inst_cell_179_26 (.BL(BL26),.BLN(BLN26),.WL(WL179));
sram_cell_6t_5 inst_cell_179_27 (.BL(BL27),.BLN(BLN27),.WL(WL179));
sram_cell_6t_5 inst_cell_179_28 (.BL(BL28),.BLN(BLN28),.WL(WL179));
sram_cell_6t_5 inst_cell_179_29 (.BL(BL29),.BLN(BLN29),.WL(WL179));
sram_cell_6t_5 inst_cell_179_30 (.BL(BL30),.BLN(BLN30),.WL(WL179));
sram_cell_6t_5 inst_cell_179_31 (.BL(BL31),.BLN(BLN31),.WL(WL179));
sram_cell_6t_5 inst_cell_179_32 (.BL(BL32),.BLN(BLN32),.WL(WL179));
sram_cell_6t_5 inst_cell_179_33 (.BL(BL33),.BLN(BLN33),.WL(WL179));
sram_cell_6t_5 inst_cell_179_34 (.BL(BL34),.BLN(BLN34),.WL(WL179));
sram_cell_6t_5 inst_cell_179_35 (.BL(BL35),.BLN(BLN35),.WL(WL179));
sram_cell_6t_5 inst_cell_179_36 (.BL(BL36),.BLN(BLN36),.WL(WL179));
sram_cell_6t_5 inst_cell_179_37 (.BL(BL37),.BLN(BLN37),.WL(WL179));
sram_cell_6t_5 inst_cell_179_38 (.BL(BL38),.BLN(BLN38),.WL(WL179));
sram_cell_6t_5 inst_cell_179_39 (.BL(BL39),.BLN(BLN39),.WL(WL179));
sram_cell_6t_5 inst_cell_179_40 (.BL(BL40),.BLN(BLN40),.WL(WL179));
sram_cell_6t_5 inst_cell_179_41 (.BL(BL41),.BLN(BLN41),.WL(WL179));
sram_cell_6t_5 inst_cell_179_42 (.BL(BL42),.BLN(BLN42),.WL(WL179));
sram_cell_6t_5 inst_cell_179_43 (.BL(BL43),.BLN(BLN43),.WL(WL179));
sram_cell_6t_5 inst_cell_179_44 (.BL(BL44),.BLN(BLN44),.WL(WL179));
sram_cell_6t_5 inst_cell_179_45 (.BL(BL45),.BLN(BLN45),.WL(WL179));
sram_cell_6t_5 inst_cell_179_46 (.BL(BL46),.BLN(BLN46),.WL(WL179));
sram_cell_6t_5 inst_cell_179_47 (.BL(BL47),.BLN(BLN47),.WL(WL179));
sram_cell_6t_5 inst_cell_179_48 (.BL(BL48),.BLN(BLN48),.WL(WL179));
sram_cell_6t_5 inst_cell_179_49 (.BL(BL49),.BLN(BLN49),.WL(WL179));
sram_cell_6t_5 inst_cell_179_50 (.BL(BL50),.BLN(BLN50),.WL(WL179));
sram_cell_6t_5 inst_cell_179_51 (.BL(BL51),.BLN(BLN51),.WL(WL179));
sram_cell_6t_5 inst_cell_179_52 (.BL(BL52),.BLN(BLN52),.WL(WL179));
sram_cell_6t_5 inst_cell_179_53 (.BL(BL53),.BLN(BLN53),.WL(WL179));
sram_cell_6t_5 inst_cell_179_54 (.BL(BL54),.BLN(BLN54),.WL(WL179));
sram_cell_6t_5 inst_cell_179_55 (.BL(BL55),.BLN(BLN55),.WL(WL179));
sram_cell_6t_5 inst_cell_179_56 (.BL(BL56),.BLN(BLN56),.WL(WL179));
sram_cell_6t_5 inst_cell_179_57 (.BL(BL57),.BLN(BLN57),.WL(WL179));
sram_cell_6t_5 inst_cell_179_58 (.BL(BL58),.BLN(BLN58),.WL(WL179));
sram_cell_6t_5 inst_cell_179_59 (.BL(BL59),.BLN(BLN59),.WL(WL179));
sram_cell_6t_5 inst_cell_179_60 (.BL(BL60),.BLN(BLN60),.WL(WL179));
sram_cell_6t_5 inst_cell_179_61 (.BL(BL61),.BLN(BLN61),.WL(WL179));
sram_cell_6t_5 inst_cell_179_62 (.BL(BL62),.BLN(BLN62),.WL(WL179));
sram_cell_6t_5 inst_cell_179_63 (.BL(BL63),.BLN(BLN63),.WL(WL179));
sram_cell_6t_5 inst_cell_179_64 (.BL(BL64),.BLN(BLN64),.WL(WL179));
sram_cell_6t_5 inst_cell_179_65 (.BL(BL65),.BLN(BLN65),.WL(WL179));
sram_cell_6t_5 inst_cell_179_66 (.BL(BL66),.BLN(BLN66),.WL(WL179));
sram_cell_6t_5 inst_cell_179_67 (.BL(BL67),.BLN(BLN67),.WL(WL179));
sram_cell_6t_5 inst_cell_179_68 (.BL(BL68),.BLN(BLN68),.WL(WL179));
sram_cell_6t_5 inst_cell_179_69 (.BL(BL69),.BLN(BLN69),.WL(WL179));
sram_cell_6t_5 inst_cell_179_70 (.BL(BL70),.BLN(BLN70),.WL(WL179));
sram_cell_6t_5 inst_cell_179_71 (.BL(BL71),.BLN(BLN71),.WL(WL179));
sram_cell_6t_5 inst_cell_179_72 (.BL(BL72),.BLN(BLN72),.WL(WL179));
sram_cell_6t_5 inst_cell_179_73 (.BL(BL73),.BLN(BLN73),.WL(WL179));
sram_cell_6t_5 inst_cell_179_74 (.BL(BL74),.BLN(BLN74),.WL(WL179));
sram_cell_6t_5 inst_cell_179_75 (.BL(BL75),.BLN(BLN75),.WL(WL179));
sram_cell_6t_5 inst_cell_179_76 (.BL(BL76),.BLN(BLN76),.WL(WL179));
sram_cell_6t_5 inst_cell_179_77 (.BL(BL77),.BLN(BLN77),.WL(WL179));
sram_cell_6t_5 inst_cell_179_78 (.BL(BL78),.BLN(BLN78),.WL(WL179));
sram_cell_6t_5 inst_cell_179_79 (.BL(BL79),.BLN(BLN79),.WL(WL179));
sram_cell_6t_5 inst_cell_179_80 (.BL(BL80),.BLN(BLN80),.WL(WL179));
sram_cell_6t_5 inst_cell_179_81 (.BL(BL81),.BLN(BLN81),.WL(WL179));
sram_cell_6t_5 inst_cell_179_82 (.BL(BL82),.BLN(BLN82),.WL(WL179));
sram_cell_6t_5 inst_cell_179_83 (.BL(BL83),.BLN(BLN83),.WL(WL179));
sram_cell_6t_5 inst_cell_179_84 (.BL(BL84),.BLN(BLN84),.WL(WL179));
sram_cell_6t_5 inst_cell_179_85 (.BL(BL85),.BLN(BLN85),.WL(WL179));
sram_cell_6t_5 inst_cell_179_86 (.BL(BL86),.BLN(BLN86),.WL(WL179));
sram_cell_6t_5 inst_cell_179_87 (.BL(BL87),.BLN(BLN87),.WL(WL179));
sram_cell_6t_5 inst_cell_179_88 (.BL(BL88),.BLN(BLN88),.WL(WL179));
sram_cell_6t_5 inst_cell_179_89 (.BL(BL89),.BLN(BLN89),.WL(WL179));
sram_cell_6t_5 inst_cell_179_90 (.BL(BL90),.BLN(BLN90),.WL(WL179));
sram_cell_6t_5 inst_cell_179_91 (.BL(BL91),.BLN(BLN91),.WL(WL179));
sram_cell_6t_5 inst_cell_179_92 (.BL(BL92),.BLN(BLN92),.WL(WL179));
sram_cell_6t_5 inst_cell_179_93 (.BL(BL93),.BLN(BLN93),.WL(WL179));
sram_cell_6t_5 inst_cell_179_94 (.BL(BL94),.BLN(BLN94),.WL(WL179));
sram_cell_6t_5 inst_cell_179_95 (.BL(BL95),.BLN(BLN95),.WL(WL179));
sram_cell_6t_5 inst_cell_179_96 (.BL(BL96),.BLN(BLN96),.WL(WL179));
sram_cell_6t_5 inst_cell_179_97 (.BL(BL97),.BLN(BLN97),.WL(WL179));
sram_cell_6t_5 inst_cell_179_98 (.BL(BL98),.BLN(BLN98),.WL(WL179));
sram_cell_6t_5 inst_cell_179_99 (.BL(BL99),.BLN(BLN99),.WL(WL179));
sram_cell_6t_5 inst_cell_179_100 (.BL(BL100),.BLN(BLN100),.WL(WL179));
sram_cell_6t_5 inst_cell_179_101 (.BL(BL101),.BLN(BLN101),.WL(WL179));
sram_cell_6t_5 inst_cell_179_102 (.BL(BL102),.BLN(BLN102),.WL(WL179));
sram_cell_6t_5 inst_cell_179_103 (.BL(BL103),.BLN(BLN103),.WL(WL179));
sram_cell_6t_5 inst_cell_179_104 (.BL(BL104),.BLN(BLN104),.WL(WL179));
sram_cell_6t_5 inst_cell_179_105 (.BL(BL105),.BLN(BLN105),.WL(WL179));
sram_cell_6t_5 inst_cell_179_106 (.BL(BL106),.BLN(BLN106),.WL(WL179));
sram_cell_6t_5 inst_cell_179_107 (.BL(BL107),.BLN(BLN107),.WL(WL179));
sram_cell_6t_5 inst_cell_179_108 (.BL(BL108),.BLN(BLN108),.WL(WL179));
sram_cell_6t_5 inst_cell_179_109 (.BL(BL109),.BLN(BLN109),.WL(WL179));
sram_cell_6t_5 inst_cell_179_110 (.BL(BL110),.BLN(BLN110),.WL(WL179));
sram_cell_6t_5 inst_cell_179_111 (.BL(BL111),.BLN(BLN111),.WL(WL179));
sram_cell_6t_5 inst_cell_179_112 (.BL(BL112),.BLN(BLN112),.WL(WL179));
sram_cell_6t_5 inst_cell_179_113 (.BL(BL113),.BLN(BLN113),.WL(WL179));
sram_cell_6t_5 inst_cell_179_114 (.BL(BL114),.BLN(BLN114),.WL(WL179));
sram_cell_6t_5 inst_cell_179_115 (.BL(BL115),.BLN(BLN115),.WL(WL179));
sram_cell_6t_5 inst_cell_179_116 (.BL(BL116),.BLN(BLN116),.WL(WL179));
sram_cell_6t_5 inst_cell_179_117 (.BL(BL117),.BLN(BLN117),.WL(WL179));
sram_cell_6t_5 inst_cell_179_118 (.BL(BL118),.BLN(BLN118),.WL(WL179));
sram_cell_6t_5 inst_cell_179_119 (.BL(BL119),.BLN(BLN119),.WL(WL179));
sram_cell_6t_5 inst_cell_179_120 (.BL(BL120),.BLN(BLN120),.WL(WL179));
sram_cell_6t_5 inst_cell_179_121 (.BL(BL121),.BLN(BLN121),.WL(WL179));
sram_cell_6t_5 inst_cell_179_122 (.BL(BL122),.BLN(BLN122),.WL(WL179));
sram_cell_6t_5 inst_cell_179_123 (.BL(BL123),.BLN(BLN123),.WL(WL179));
sram_cell_6t_5 inst_cell_179_124 (.BL(BL124),.BLN(BLN124),.WL(WL179));
sram_cell_6t_5 inst_cell_179_125 (.BL(BL125),.BLN(BLN125),.WL(WL179));
sram_cell_6t_5 inst_cell_179_126 (.BL(BL126),.BLN(BLN126),.WL(WL179));
sram_cell_6t_5 inst_cell_179_127 (.BL(BL127),.BLN(BLN127),.WL(WL179));
sram_cell_6t_5 inst_cell_180_0 (.BL(BL0),.BLN(BLN0),.WL(WL180));
sram_cell_6t_5 inst_cell_180_1 (.BL(BL1),.BLN(BLN1),.WL(WL180));
sram_cell_6t_5 inst_cell_180_2 (.BL(BL2),.BLN(BLN2),.WL(WL180));
sram_cell_6t_5 inst_cell_180_3 (.BL(BL3),.BLN(BLN3),.WL(WL180));
sram_cell_6t_5 inst_cell_180_4 (.BL(BL4),.BLN(BLN4),.WL(WL180));
sram_cell_6t_5 inst_cell_180_5 (.BL(BL5),.BLN(BLN5),.WL(WL180));
sram_cell_6t_5 inst_cell_180_6 (.BL(BL6),.BLN(BLN6),.WL(WL180));
sram_cell_6t_5 inst_cell_180_7 (.BL(BL7),.BLN(BLN7),.WL(WL180));
sram_cell_6t_5 inst_cell_180_8 (.BL(BL8),.BLN(BLN8),.WL(WL180));
sram_cell_6t_5 inst_cell_180_9 (.BL(BL9),.BLN(BLN9),.WL(WL180));
sram_cell_6t_5 inst_cell_180_10 (.BL(BL10),.BLN(BLN10),.WL(WL180));
sram_cell_6t_5 inst_cell_180_11 (.BL(BL11),.BLN(BLN11),.WL(WL180));
sram_cell_6t_5 inst_cell_180_12 (.BL(BL12),.BLN(BLN12),.WL(WL180));
sram_cell_6t_5 inst_cell_180_13 (.BL(BL13),.BLN(BLN13),.WL(WL180));
sram_cell_6t_5 inst_cell_180_14 (.BL(BL14),.BLN(BLN14),.WL(WL180));
sram_cell_6t_5 inst_cell_180_15 (.BL(BL15),.BLN(BLN15),.WL(WL180));
sram_cell_6t_5 inst_cell_180_16 (.BL(BL16),.BLN(BLN16),.WL(WL180));
sram_cell_6t_5 inst_cell_180_17 (.BL(BL17),.BLN(BLN17),.WL(WL180));
sram_cell_6t_5 inst_cell_180_18 (.BL(BL18),.BLN(BLN18),.WL(WL180));
sram_cell_6t_5 inst_cell_180_19 (.BL(BL19),.BLN(BLN19),.WL(WL180));
sram_cell_6t_5 inst_cell_180_20 (.BL(BL20),.BLN(BLN20),.WL(WL180));
sram_cell_6t_5 inst_cell_180_21 (.BL(BL21),.BLN(BLN21),.WL(WL180));
sram_cell_6t_5 inst_cell_180_22 (.BL(BL22),.BLN(BLN22),.WL(WL180));
sram_cell_6t_5 inst_cell_180_23 (.BL(BL23),.BLN(BLN23),.WL(WL180));
sram_cell_6t_5 inst_cell_180_24 (.BL(BL24),.BLN(BLN24),.WL(WL180));
sram_cell_6t_5 inst_cell_180_25 (.BL(BL25),.BLN(BLN25),.WL(WL180));
sram_cell_6t_5 inst_cell_180_26 (.BL(BL26),.BLN(BLN26),.WL(WL180));
sram_cell_6t_5 inst_cell_180_27 (.BL(BL27),.BLN(BLN27),.WL(WL180));
sram_cell_6t_5 inst_cell_180_28 (.BL(BL28),.BLN(BLN28),.WL(WL180));
sram_cell_6t_5 inst_cell_180_29 (.BL(BL29),.BLN(BLN29),.WL(WL180));
sram_cell_6t_5 inst_cell_180_30 (.BL(BL30),.BLN(BLN30),.WL(WL180));
sram_cell_6t_5 inst_cell_180_31 (.BL(BL31),.BLN(BLN31),.WL(WL180));
sram_cell_6t_5 inst_cell_180_32 (.BL(BL32),.BLN(BLN32),.WL(WL180));
sram_cell_6t_5 inst_cell_180_33 (.BL(BL33),.BLN(BLN33),.WL(WL180));
sram_cell_6t_5 inst_cell_180_34 (.BL(BL34),.BLN(BLN34),.WL(WL180));
sram_cell_6t_5 inst_cell_180_35 (.BL(BL35),.BLN(BLN35),.WL(WL180));
sram_cell_6t_5 inst_cell_180_36 (.BL(BL36),.BLN(BLN36),.WL(WL180));
sram_cell_6t_5 inst_cell_180_37 (.BL(BL37),.BLN(BLN37),.WL(WL180));
sram_cell_6t_5 inst_cell_180_38 (.BL(BL38),.BLN(BLN38),.WL(WL180));
sram_cell_6t_5 inst_cell_180_39 (.BL(BL39),.BLN(BLN39),.WL(WL180));
sram_cell_6t_5 inst_cell_180_40 (.BL(BL40),.BLN(BLN40),.WL(WL180));
sram_cell_6t_5 inst_cell_180_41 (.BL(BL41),.BLN(BLN41),.WL(WL180));
sram_cell_6t_5 inst_cell_180_42 (.BL(BL42),.BLN(BLN42),.WL(WL180));
sram_cell_6t_5 inst_cell_180_43 (.BL(BL43),.BLN(BLN43),.WL(WL180));
sram_cell_6t_5 inst_cell_180_44 (.BL(BL44),.BLN(BLN44),.WL(WL180));
sram_cell_6t_5 inst_cell_180_45 (.BL(BL45),.BLN(BLN45),.WL(WL180));
sram_cell_6t_5 inst_cell_180_46 (.BL(BL46),.BLN(BLN46),.WL(WL180));
sram_cell_6t_5 inst_cell_180_47 (.BL(BL47),.BLN(BLN47),.WL(WL180));
sram_cell_6t_5 inst_cell_180_48 (.BL(BL48),.BLN(BLN48),.WL(WL180));
sram_cell_6t_5 inst_cell_180_49 (.BL(BL49),.BLN(BLN49),.WL(WL180));
sram_cell_6t_5 inst_cell_180_50 (.BL(BL50),.BLN(BLN50),.WL(WL180));
sram_cell_6t_5 inst_cell_180_51 (.BL(BL51),.BLN(BLN51),.WL(WL180));
sram_cell_6t_5 inst_cell_180_52 (.BL(BL52),.BLN(BLN52),.WL(WL180));
sram_cell_6t_5 inst_cell_180_53 (.BL(BL53),.BLN(BLN53),.WL(WL180));
sram_cell_6t_5 inst_cell_180_54 (.BL(BL54),.BLN(BLN54),.WL(WL180));
sram_cell_6t_5 inst_cell_180_55 (.BL(BL55),.BLN(BLN55),.WL(WL180));
sram_cell_6t_5 inst_cell_180_56 (.BL(BL56),.BLN(BLN56),.WL(WL180));
sram_cell_6t_5 inst_cell_180_57 (.BL(BL57),.BLN(BLN57),.WL(WL180));
sram_cell_6t_5 inst_cell_180_58 (.BL(BL58),.BLN(BLN58),.WL(WL180));
sram_cell_6t_5 inst_cell_180_59 (.BL(BL59),.BLN(BLN59),.WL(WL180));
sram_cell_6t_5 inst_cell_180_60 (.BL(BL60),.BLN(BLN60),.WL(WL180));
sram_cell_6t_5 inst_cell_180_61 (.BL(BL61),.BLN(BLN61),.WL(WL180));
sram_cell_6t_5 inst_cell_180_62 (.BL(BL62),.BLN(BLN62),.WL(WL180));
sram_cell_6t_5 inst_cell_180_63 (.BL(BL63),.BLN(BLN63),.WL(WL180));
sram_cell_6t_5 inst_cell_180_64 (.BL(BL64),.BLN(BLN64),.WL(WL180));
sram_cell_6t_5 inst_cell_180_65 (.BL(BL65),.BLN(BLN65),.WL(WL180));
sram_cell_6t_5 inst_cell_180_66 (.BL(BL66),.BLN(BLN66),.WL(WL180));
sram_cell_6t_5 inst_cell_180_67 (.BL(BL67),.BLN(BLN67),.WL(WL180));
sram_cell_6t_5 inst_cell_180_68 (.BL(BL68),.BLN(BLN68),.WL(WL180));
sram_cell_6t_5 inst_cell_180_69 (.BL(BL69),.BLN(BLN69),.WL(WL180));
sram_cell_6t_5 inst_cell_180_70 (.BL(BL70),.BLN(BLN70),.WL(WL180));
sram_cell_6t_5 inst_cell_180_71 (.BL(BL71),.BLN(BLN71),.WL(WL180));
sram_cell_6t_5 inst_cell_180_72 (.BL(BL72),.BLN(BLN72),.WL(WL180));
sram_cell_6t_5 inst_cell_180_73 (.BL(BL73),.BLN(BLN73),.WL(WL180));
sram_cell_6t_5 inst_cell_180_74 (.BL(BL74),.BLN(BLN74),.WL(WL180));
sram_cell_6t_5 inst_cell_180_75 (.BL(BL75),.BLN(BLN75),.WL(WL180));
sram_cell_6t_5 inst_cell_180_76 (.BL(BL76),.BLN(BLN76),.WL(WL180));
sram_cell_6t_5 inst_cell_180_77 (.BL(BL77),.BLN(BLN77),.WL(WL180));
sram_cell_6t_5 inst_cell_180_78 (.BL(BL78),.BLN(BLN78),.WL(WL180));
sram_cell_6t_5 inst_cell_180_79 (.BL(BL79),.BLN(BLN79),.WL(WL180));
sram_cell_6t_5 inst_cell_180_80 (.BL(BL80),.BLN(BLN80),.WL(WL180));
sram_cell_6t_5 inst_cell_180_81 (.BL(BL81),.BLN(BLN81),.WL(WL180));
sram_cell_6t_5 inst_cell_180_82 (.BL(BL82),.BLN(BLN82),.WL(WL180));
sram_cell_6t_5 inst_cell_180_83 (.BL(BL83),.BLN(BLN83),.WL(WL180));
sram_cell_6t_5 inst_cell_180_84 (.BL(BL84),.BLN(BLN84),.WL(WL180));
sram_cell_6t_5 inst_cell_180_85 (.BL(BL85),.BLN(BLN85),.WL(WL180));
sram_cell_6t_5 inst_cell_180_86 (.BL(BL86),.BLN(BLN86),.WL(WL180));
sram_cell_6t_5 inst_cell_180_87 (.BL(BL87),.BLN(BLN87),.WL(WL180));
sram_cell_6t_5 inst_cell_180_88 (.BL(BL88),.BLN(BLN88),.WL(WL180));
sram_cell_6t_5 inst_cell_180_89 (.BL(BL89),.BLN(BLN89),.WL(WL180));
sram_cell_6t_5 inst_cell_180_90 (.BL(BL90),.BLN(BLN90),.WL(WL180));
sram_cell_6t_5 inst_cell_180_91 (.BL(BL91),.BLN(BLN91),.WL(WL180));
sram_cell_6t_5 inst_cell_180_92 (.BL(BL92),.BLN(BLN92),.WL(WL180));
sram_cell_6t_5 inst_cell_180_93 (.BL(BL93),.BLN(BLN93),.WL(WL180));
sram_cell_6t_5 inst_cell_180_94 (.BL(BL94),.BLN(BLN94),.WL(WL180));
sram_cell_6t_5 inst_cell_180_95 (.BL(BL95),.BLN(BLN95),.WL(WL180));
sram_cell_6t_5 inst_cell_180_96 (.BL(BL96),.BLN(BLN96),.WL(WL180));
sram_cell_6t_5 inst_cell_180_97 (.BL(BL97),.BLN(BLN97),.WL(WL180));
sram_cell_6t_5 inst_cell_180_98 (.BL(BL98),.BLN(BLN98),.WL(WL180));
sram_cell_6t_5 inst_cell_180_99 (.BL(BL99),.BLN(BLN99),.WL(WL180));
sram_cell_6t_5 inst_cell_180_100 (.BL(BL100),.BLN(BLN100),.WL(WL180));
sram_cell_6t_5 inst_cell_180_101 (.BL(BL101),.BLN(BLN101),.WL(WL180));
sram_cell_6t_5 inst_cell_180_102 (.BL(BL102),.BLN(BLN102),.WL(WL180));
sram_cell_6t_5 inst_cell_180_103 (.BL(BL103),.BLN(BLN103),.WL(WL180));
sram_cell_6t_5 inst_cell_180_104 (.BL(BL104),.BLN(BLN104),.WL(WL180));
sram_cell_6t_5 inst_cell_180_105 (.BL(BL105),.BLN(BLN105),.WL(WL180));
sram_cell_6t_5 inst_cell_180_106 (.BL(BL106),.BLN(BLN106),.WL(WL180));
sram_cell_6t_5 inst_cell_180_107 (.BL(BL107),.BLN(BLN107),.WL(WL180));
sram_cell_6t_5 inst_cell_180_108 (.BL(BL108),.BLN(BLN108),.WL(WL180));
sram_cell_6t_5 inst_cell_180_109 (.BL(BL109),.BLN(BLN109),.WL(WL180));
sram_cell_6t_5 inst_cell_180_110 (.BL(BL110),.BLN(BLN110),.WL(WL180));
sram_cell_6t_5 inst_cell_180_111 (.BL(BL111),.BLN(BLN111),.WL(WL180));
sram_cell_6t_5 inst_cell_180_112 (.BL(BL112),.BLN(BLN112),.WL(WL180));
sram_cell_6t_5 inst_cell_180_113 (.BL(BL113),.BLN(BLN113),.WL(WL180));
sram_cell_6t_5 inst_cell_180_114 (.BL(BL114),.BLN(BLN114),.WL(WL180));
sram_cell_6t_5 inst_cell_180_115 (.BL(BL115),.BLN(BLN115),.WL(WL180));
sram_cell_6t_5 inst_cell_180_116 (.BL(BL116),.BLN(BLN116),.WL(WL180));
sram_cell_6t_5 inst_cell_180_117 (.BL(BL117),.BLN(BLN117),.WL(WL180));
sram_cell_6t_5 inst_cell_180_118 (.BL(BL118),.BLN(BLN118),.WL(WL180));
sram_cell_6t_5 inst_cell_180_119 (.BL(BL119),.BLN(BLN119),.WL(WL180));
sram_cell_6t_5 inst_cell_180_120 (.BL(BL120),.BLN(BLN120),.WL(WL180));
sram_cell_6t_5 inst_cell_180_121 (.BL(BL121),.BLN(BLN121),.WL(WL180));
sram_cell_6t_5 inst_cell_180_122 (.BL(BL122),.BLN(BLN122),.WL(WL180));
sram_cell_6t_5 inst_cell_180_123 (.BL(BL123),.BLN(BLN123),.WL(WL180));
sram_cell_6t_5 inst_cell_180_124 (.BL(BL124),.BLN(BLN124),.WL(WL180));
sram_cell_6t_5 inst_cell_180_125 (.BL(BL125),.BLN(BLN125),.WL(WL180));
sram_cell_6t_5 inst_cell_180_126 (.BL(BL126),.BLN(BLN126),.WL(WL180));
sram_cell_6t_5 inst_cell_180_127 (.BL(BL127),.BLN(BLN127),.WL(WL180));
sram_cell_6t_5 inst_cell_181_0 (.BL(BL0),.BLN(BLN0),.WL(WL181));
sram_cell_6t_5 inst_cell_181_1 (.BL(BL1),.BLN(BLN1),.WL(WL181));
sram_cell_6t_5 inst_cell_181_2 (.BL(BL2),.BLN(BLN2),.WL(WL181));
sram_cell_6t_5 inst_cell_181_3 (.BL(BL3),.BLN(BLN3),.WL(WL181));
sram_cell_6t_5 inst_cell_181_4 (.BL(BL4),.BLN(BLN4),.WL(WL181));
sram_cell_6t_5 inst_cell_181_5 (.BL(BL5),.BLN(BLN5),.WL(WL181));
sram_cell_6t_5 inst_cell_181_6 (.BL(BL6),.BLN(BLN6),.WL(WL181));
sram_cell_6t_5 inst_cell_181_7 (.BL(BL7),.BLN(BLN7),.WL(WL181));
sram_cell_6t_5 inst_cell_181_8 (.BL(BL8),.BLN(BLN8),.WL(WL181));
sram_cell_6t_5 inst_cell_181_9 (.BL(BL9),.BLN(BLN9),.WL(WL181));
sram_cell_6t_5 inst_cell_181_10 (.BL(BL10),.BLN(BLN10),.WL(WL181));
sram_cell_6t_5 inst_cell_181_11 (.BL(BL11),.BLN(BLN11),.WL(WL181));
sram_cell_6t_5 inst_cell_181_12 (.BL(BL12),.BLN(BLN12),.WL(WL181));
sram_cell_6t_5 inst_cell_181_13 (.BL(BL13),.BLN(BLN13),.WL(WL181));
sram_cell_6t_5 inst_cell_181_14 (.BL(BL14),.BLN(BLN14),.WL(WL181));
sram_cell_6t_5 inst_cell_181_15 (.BL(BL15),.BLN(BLN15),.WL(WL181));
sram_cell_6t_5 inst_cell_181_16 (.BL(BL16),.BLN(BLN16),.WL(WL181));
sram_cell_6t_5 inst_cell_181_17 (.BL(BL17),.BLN(BLN17),.WL(WL181));
sram_cell_6t_5 inst_cell_181_18 (.BL(BL18),.BLN(BLN18),.WL(WL181));
sram_cell_6t_5 inst_cell_181_19 (.BL(BL19),.BLN(BLN19),.WL(WL181));
sram_cell_6t_5 inst_cell_181_20 (.BL(BL20),.BLN(BLN20),.WL(WL181));
sram_cell_6t_5 inst_cell_181_21 (.BL(BL21),.BLN(BLN21),.WL(WL181));
sram_cell_6t_5 inst_cell_181_22 (.BL(BL22),.BLN(BLN22),.WL(WL181));
sram_cell_6t_5 inst_cell_181_23 (.BL(BL23),.BLN(BLN23),.WL(WL181));
sram_cell_6t_5 inst_cell_181_24 (.BL(BL24),.BLN(BLN24),.WL(WL181));
sram_cell_6t_5 inst_cell_181_25 (.BL(BL25),.BLN(BLN25),.WL(WL181));
sram_cell_6t_5 inst_cell_181_26 (.BL(BL26),.BLN(BLN26),.WL(WL181));
sram_cell_6t_5 inst_cell_181_27 (.BL(BL27),.BLN(BLN27),.WL(WL181));
sram_cell_6t_5 inst_cell_181_28 (.BL(BL28),.BLN(BLN28),.WL(WL181));
sram_cell_6t_5 inst_cell_181_29 (.BL(BL29),.BLN(BLN29),.WL(WL181));
sram_cell_6t_5 inst_cell_181_30 (.BL(BL30),.BLN(BLN30),.WL(WL181));
sram_cell_6t_5 inst_cell_181_31 (.BL(BL31),.BLN(BLN31),.WL(WL181));
sram_cell_6t_5 inst_cell_181_32 (.BL(BL32),.BLN(BLN32),.WL(WL181));
sram_cell_6t_5 inst_cell_181_33 (.BL(BL33),.BLN(BLN33),.WL(WL181));
sram_cell_6t_5 inst_cell_181_34 (.BL(BL34),.BLN(BLN34),.WL(WL181));
sram_cell_6t_5 inst_cell_181_35 (.BL(BL35),.BLN(BLN35),.WL(WL181));
sram_cell_6t_5 inst_cell_181_36 (.BL(BL36),.BLN(BLN36),.WL(WL181));
sram_cell_6t_5 inst_cell_181_37 (.BL(BL37),.BLN(BLN37),.WL(WL181));
sram_cell_6t_5 inst_cell_181_38 (.BL(BL38),.BLN(BLN38),.WL(WL181));
sram_cell_6t_5 inst_cell_181_39 (.BL(BL39),.BLN(BLN39),.WL(WL181));
sram_cell_6t_5 inst_cell_181_40 (.BL(BL40),.BLN(BLN40),.WL(WL181));
sram_cell_6t_5 inst_cell_181_41 (.BL(BL41),.BLN(BLN41),.WL(WL181));
sram_cell_6t_5 inst_cell_181_42 (.BL(BL42),.BLN(BLN42),.WL(WL181));
sram_cell_6t_5 inst_cell_181_43 (.BL(BL43),.BLN(BLN43),.WL(WL181));
sram_cell_6t_5 inst_cell_181_44 (.BL(BL44),.BLN(BLN44),.WL(WL181));
sram_cell_6t_5 inst_cell_181_45 (.BL(BL45),.BLN(BLN45),.WL(WL181));
sram_cell_6t_5 inst_cell_181_46 (.BL(BL46),.BLN(BLN46),.WL(WL181));
sram_cell_6t_5 inst_cell_181_47 (.BL(BL47),.BLN(BLN47),.WL(WL181));
sram_cell_6t_5 inst_cell_181_48 (.BL(BL48),.BLN(BLN48),.WL(WL181));
sram_cell_6t_5 inst_cell_181_49 (.BL(BL49),.BLN(BLN49),.WL(WL181));
sram_cell_6t_5 inst_cell_181_50 (.BL(BL50),.BLN(BLN50),.WL(WL181));
sram_cell_6t_5 inst_cell_181_51 (.BL(BL51),.BLN(BLN51),.WL(WL181));
sram_cell_6t_5 inst_cell_181_52 (.BL(BL52),.BLN(BLN52),.WL(WL181));
sram_cell_6t_5 inst_cell_181_53 (.BL(BL53),.BLN(BLN53),.WL(WL181));
sram_cell_6t_5 inst_cell_181_54 (.BL(BL54),.BLN(BLN54),.WL(WL181));
sram_cell_6t_5 inst_cell_181_55 (.BL(BL55),.BLN(BLN55),.WL(WL181));
sram_cell_6t_5 inst_cell_181_56 (.BL(BL56),.BLN(BLN56),.WL(WL181));
sram_cell_6t_5 inst_cell_181_57 (.BL(BL57),.BLN(BLN57),.WL(WL181));
sram_cell_6t_5 inst_cell_181_58 (.BL(BL58),.BLN(BLN58),.WL(WL181));
sram_cell_6t_5 inst_cell_181_59 (.BL(BL59),.BLN(BLN59),.WL(WL181));
sram_cell_6t_5 inst_cell_181_60 (.BL(BL60),.BLN(BLN60),.WL(WL181));
sram_cell_6t_5 inst_cell_181_61 (.BL(BL61),.BLN(BLN61),.WL(WL181));
sram_cell_6t_5 inst_cell_181_62 (.BL(BL62),.BLN(BLN62),.WL(WL181));
sram_cell_6t_5 inst_cell_181_63 (.BL(BL63),.BLN(BLN63),.WL(WL181));
sram_cell_6t_5 inst_cell_181_64 (.BL(BL64),.BLN(BLN64),.WL(WL181));
sram_cell_6t_5 inst_cell_181_65 (.BL(BL65),.BLN(BLN65),.WL(WL181));
sram_cell_6t_5 inst_cell_181_66 (.BL(BL66),.BLN(BLN66),.WL(WL181));
sram_cell_6t_5 inst_cell_181_67 (.BL(BL67),.BLN(BLN67),.WL(WL181));
sram_cell_6t_5 inst_cell_181_68 (.BL(BL68),.BLN(BLN68),.WL(WL181));
sram_cell_6t_5 inst_cell_181_69 (.BL(BL69),.BLN(BLN69),.WL(WL181));
sram_cell_6t_5 inst_cell_181_70 (.BL(BL70),.BLN(BLN70),.WL(WL181));
sram_cell_6t_5 inst_cell_181_71 (.BL(BL71),.BLN(BLN71),.WL(WL181));
sram_cell_6t_5 inst_cell_181_72 (.BL(BL72),.BLN(BLN72),.WL(WL181));
sram_cell_6t_5 inst_cell_181_73 (.BL(BL73),.BLN(BLN73),.WL(WL181));
sram_cell_6t_5 inst_cell_181_74 (.BL(BL74),.BLN(BLN74),.WL(WL181));
sram_cell_6t_5 inst_cell_181_75 (.BL(BL75),.BLN(BLN75),.WL(WL181));
sram_cell_6t_5 inst_cell_181_76 (.BL(BL76),.BLN(BLN76),.WL(WL181));
sram_cell_6t_5 inst_cell_181_77 (.BL(BL77),.BLN(BLN77),.WL(WL181));
sram_cell_6t_5 inst_cell_181_78 (.BL(BL78),.BLN(BLN78),.WL(WL181));
sram_cell_6t_5 inst_cell_181_79 (.BL(BL79),.BLN(BLN79),.WL(WL181));
sram_cell_6t_5 inst_cell_181_80 (.BL(BL80),.BLN(BLN80),.WL(WL181));
sram_cell_6t_5 inst_cell_181_81 (.BL(BL81),.BLN(BLN81),.WL(WL181));
sram_cell_6t_5 inst_cell_181_82 (.BL(BL82),.BLN(BLN82),.WL(WL181));
sram_cell_6t_5 inst_cell_181_83 (.BL(BL83),.BLN(BLN83),.WL(WL181));
sram_cell_6t_5 inst_cell_181_84 (.BL(BL84),.BLN(BLN84),.WL(WL181));
sram_cell_6t_5 inst_cell_181_85 (.BL(BL85),.BLN(BLN85),.WL(WL181));
sram_cell_6t_5 inst_cell_181_86 (.BL(BL86),.BLN(BLN86),.WL(WL181));
sram_cell_6t_5 inst_cell_181_87 (.BL(BL87),.BLN(BLN87),.WL(WL181));
sram_cell_6t_5 inst_cell_181_88 (.BL(BL88),.BLN(BLN88),.WL(WL181));
sram_cell_6t_5 inst_cell_181_89 (.BL(BL89),.BLN(BLN89),.WL(WL181));
sram_cell_6t_5 inst_cell_181_90 (.BL(BL90),.BLN(BLN90),.WL(WL181));
sram_cell_6t_5 inst_cell_181_91 (.BL(BL91),.BLN(BLN91),.WL(WL181));
sram_cell_6t_5 inst_cell_181_92 (.BL(BL92),.BLN(BLN92),.WL(WL181));
sram_cell_6t_5 inst_cell_181_93 (.BL(BL93),.BLN(BLN93),.WL(WL181));
sram_cell_6t_5 inst_cell_181_94 (.BL(BL94),.BLN(BLN94),.WL(WL181));
sram_cell_6t_5 inst_cell_181_95 (.BL(BL95),.BLN(BLN95),.WL(WL181));
sram_cell_6t_5 inst_cell_181_96 (.BL(BL96),.BLN(BLN96),.WL(WL181));
sram_cell_6t_5 inst_cell_181_97 (.BL(BL97),.BLN(BLN97),.WL(WL181));
sram_cell_6t_5 inst_cell_181_98 (.BL(BL98),.BLN(BLN98),.WL(WL181));
sram_cell_6t_5 inst_cell_181_99 (.BL(BL99),.BLN(BLN99),.WL(WL181));
sram_cell_6t_5 inst_cell_181_100 (.BL(BL100),.BLN(BLN100),.WL(WL181));
sram_cell_6t_5 inst_cell_181_101 (.BL(BL101),.BLN(BLN101),.WL(WL181));
sram_cell_6t_5 inst_cell_181_102 (.BL(BL102),.BLN(BLN102),.WL(WL181));
sram_cell_6t_5 inst_cell_181_103 (.BL(BL103),.BLN(BLN103),.WL(WL181));
sram_cell_6t_5 inst_cell_181_104 (.BL(BL104),.BLN(BLN104),.WL(WL181));
sram_cell_6t_5 inst_cell_181_105 (.BL(BL105),.BLN(BLN105),.WL(WL181));
sram_cell_6t_5 inst_cell_181_106 (.BL(BL106),.BLN(BLN106),.WL(WL181));
sram_cell_6t_5 inst_cell_181_107 (.BL(BL107),.BLN(BLN107),.WL(WL181));
sram_cell_6t_5 inst_cell_181_108 (.BL(BL108),.BLN(BLN108),.WL(WL181));
sram_cell_6t_5 inst_cell_181_109 (.BL(BL109),.BLN(BLN109),.WL(WL181));
sram_cell_6t_5 inst_cell_181_110 (.BL(BL110),.BLN(BLN110),.WL(WL181));
sram_cell_6t_5 inst_cell_181_111 (.BL(BL111),.BLN(BLN111),.WL(WL181));
sram_cell_6t_5 inst_cell_181_112 (.BL(BL112),.BLN(BLN112),.WL(WL181));
sram_cell_6t_5 inst_cell_181_113 (.BL(BL113),.BLN(BLN113),.WL(WL181));
sram_cell_6t_5 inst_cell_181_114 (.BL(BL114),.BLN(BLN114),.WL(WL181));
sram_cell_6t_5 inst_cell_181_115 (.BL(BL115),.BLN(BLN115),.WL(WL181));
sram_cell_6t_5 inst_cell_181_116 (.BL(BL116),.BLN(BLN116),.WL(WL181));
sram_cell_6t_5 inst_cell_181_117 (.BL(BL117),.BLN(BLN117),.WL(WL181));
sram_cell_6t_5 inst_cell_181_118 (.BL(BL118),.BLN(BLN118),.WL(WL181));
sram_cell_6t_5 inst_cell_181_119 (.BL(BL119),.BLN(BLN119),.WL(WL181));
sram_cell_6t_5 inst_cell_181_120 (.BL(BL120),.BLN(BLN120),.WL(WL181));
sram_cell_6t_5 inst_cell_181_121 (.BL(BL121),.BLN(BLN121),.WL(WL181));
sram_cell_6t_5 inst_cell_181_122 (.BL(BL122),.BLN(BLN122),.WL(WL181));
sram_cell_6t_5 inst_cell_181_123 (.BL(BL123),.BLN(BLN123),.WL(WL181));
sram_cell_6t_5 inst_cell_181_124 (.BL(BL124),.BLN(BLN124),.WL(WL181));
sram_cell_6t_5 inst_cell_181_125 (.BL(BL125),.BLN(BLN125),.WL(WL181));
sram_cell_6t_5 inst_cell_181_126 (.BL(BL126),.BLN(BLN126),.WL(WL181));
sram_cell_6t_5 inst_cell_181_127 (.BL(BL127),.BLN(BLN127),.WL(WL181));
sram_cell_6t_5 inst_cell_182_0 (.BL(BL0),.BLN(BLN0),.WL(WL182));
sram_cell_6t_5 inst_cell_182_1 (.BL(BL1),.BLN(BLN1),.WL(WL182));
sram_cell_6t_5 inst_cell_182_2 (.BL(BL2),.BLN(BLN2),.WL(WL182));
sram_cell_6t_5 inst_cell_182_3 (.BL(BL3),.BLN(BLN3),.WL(WL182));
sram_cell_6t_5 inst_cell_182_4 (.BL(BL4),.BLN(BLN4),.WL(WL182));
sram_cell_6t_5 inst_cell_182_5 (.BL(BL5),.BLN(BLN5),.WL(WL182));
sram_cell_6t_5 inst_cell_182_6 (.BL(BL6),.BLN(BLN6),.WL(WL182));
sram_cell_6t_5 inst_cell_182_7 (.BL(BL7),.BLN(BLN7),.WL(WL182));
sram_cell_6t_5 inst_cell_182_8 (.BL(BL8),.BLN(BLN8),.WL(WL182));
sram_cell_6t_5 inst_cell_182_9 (.BL(BL9),.BLN(BLN9),.WL(WL182));
sram_cell_6t_5 inst_cell_182_10 (.BL(BL10),.BLN(BLN10),.WL(WL182));
sram_cell_6t_5 inst_cell_182_11 (.BL(BL11),.BLN(BLN11),.WL(WL182));
sram_cell_6t_5 inst_cell_182_12 (.BL(BL12),.BLN(BLN12),.WL(WL182));
sram_cell_6t_5 inst_cell_182_13 (.BL(BL13),.BLN(BLN13),.WL(WL182));
sram_cell_6t_5 inst_cell_182_14 (.BL(BL14),.BLN(BLN14),.WL(WL182));
sram_cell_6t_5 inst_cell_182_15 (.BL(BL15),.BLN(BLN15),.WL(WL182));
sram_cell_6t_5 inst_cell_182_16 (.BL(BL16),.BLN(BLN16),.WL(WL182));
sram_cell_6t_5 inst_cell_182_17 (.BL(BL17),.BLN(BLN17),.WL(WL182));
sram_cell_6t_5 inst_cell_182_18 (.BL(BL18),.BLN(BLN18),.WL(WL182));
sram_cell_6t_5 inst_cell_182_19 (.BL(BL19),.BLN(BLN19),.WL(WL182));
sram_cell_6t_5 inst_cell_182_20 (.BL(BL20),.BLN(BLN20),.WL(WL182));
sram_cell_6t_5 inst_cell_182_21 (.BL(BL21),.BLN(BLN21),.WL(WL182));
sram_cell_6t_5 inst_cell_182_22 (.BL(BL22),.BLN(BLN22),.WL(WL182));
sram_cell_6t_5 inst_cell_182_23 (.BL(BL23),.BLN(BLN23),.WL(WL182));
sram_cell_6t_5 inst_cell_182_24 (.BL(BL24),.BLN(BLN24),.WL(WL182));
sram_cell_6t_5 inst_cell_182_25 (.BL(BL25),.BLN(BLN25),.WL(WL182));
sram_cell_6t_5 inst_cell_182_26 (.BL(BL26),.BLN(BLN26),.WL(WL182));
sram_cell_6t_5 inst_cell_182_27 (.BL(BL27),.BLN(BLN27),.WL(WL182));
sram_cell_6t_5 inst_cell_182_28 (.BL(BL28),.BLN(BLN28),.WL(WL182));
sram_cell_6t_5 inst_cell_182_29 (.BL(BL29),.BLN(BLN29),.WL(WL182));
sram_cell_6t_5 inst_cell_182_30 (.BL(BL30),.BLN(BLN30),.WL(WL182));
sram_cell_6t_5 inst_cell_182_31 (.BL(BL31),.BLN(BLN31),.WL(WL182));
sram_cell_6t_5 inst_cell_182_32 (.BL(BL32),.BLN(BLN32),.WL(WL182));
sram_cell_6t_5 inst_cell_182_33 (.BL(BL33),.BLN(BLN33),.WL(WL182));
sram_cell_6t_5 inst_cell_182_34 (.BL(BL34),.BLN(BLN34),.WL(WL182));
sram_cell_6t_5 inst_cell_182_35 (.BL(BL35),.BLN(BLN35),.WL(WL182));
sram_cell_6t_5 inst_cell_182_36 (.BL(BL36),.BLN(BLN36),.WL(WL182));
sram_cell_6t_5 inst_cell_182_37 (.BL(BL37),.BLN(BLN37),.WL(WL182));
sram_cell_6t_5 inst_cell_182_38 (.BL(BL38),.BLN(BLN38),.WL(WL182));
sram_cell_6t_5 inst_cell_182_39 (.BL(BL39),.BLN(BLN39),.WL(WL182));
sram_cell_6t_5 inst_cell_182_40 (.BL(BL40),.BLN(BLN40),.WL(WL182));
sram_cell_6t_5 inst_cell_182_41 (.BL(BL41),.BLN(BLN41),.WL(WL182));
sram_cell_6t_5 inst_cell_182_42 (.BL(BL42),.BLN(BLN42),.WL(WL182));
sram_cell_6t_5 inst_cell_182_43 (.BL(BL43),.BLN(BLN43),.WL(WL182));
sram_cell_6t_5 inst_cell_182_44 (.BL(BL44),.BLN(BLN44),.WL(WL182));
sram_cell_6t_5 inst_cell_182_45 (.BL(BL45),.BLN(BLN45),.WL(WL182));
sram_cell_6t_5 inst_cell_182_46 (.BL(BL46),.BLN(BLN46),.WL(WL182));
sram_cell_6t_5 inst_cell_182_47 (.BL(BL47),.BLN(BLN47),.WL(WL182));
sram_cell_6t_5 inst_cell_182_48 (.BL(BL48),.BLN(BLN48),.WL(WL182));
sram_cell_6t_5 inst_cell_182_49 (.BL(BL49),.BLN(BLN49),.WL(WL182));
sram_cell_6t_5 inst_cell_182_50 (.BL(BL50),.BLN(BLN50),.WL(WL182));
sram_cell_6t_5 inst_cell_182_51 (.BL(BL51),.BLN(BLN51),.WL(WL182));
sram_cell_6t_5 inst_cell_182_52 (.BL(BL52),.BLN(BLN52),.WL(WL182));
sram_cell_6t_5 inst_cell_182_53 (.BL(BL53),.BLN(BLN53),.WL(WL182));
sram_cell_6t_5 inst_cell_182_54 (.BL(BL54),.BLN(BLN54),.WL(WL182));
sram_cell_6t_5 inst_cell_182_55 (.BL(BL55),.BLN(BLN55),.WL(WL182));
sram_cell_6t_5 inst_cell_182_56 (.BL(BL56),.BLN(BLN56),.WL(WL182));
sram_cell_6t_5 inst_cell_182_57 (.BL(BL57),.BLN(BLN57),.WL(WL182));
sram_cell_6t_5 inst_cell_182_58 (.BL(BL58),.BLN(BLN58),.WL(WL182));
sram_cell_6t_5 inst_cell_182_59 (.BL(BL59),.BLN(BLN59),.WL(WL182));
sram_cell_6t_5 inst_cell_182_60 (.BL(BL60),.BLN(BLN60),.WL(WL182));
sram_cell_6t_5 inst_cell_182_61 (.BL(BL61),.BLN(BLN61),.WL(WL182));
sram_cell_6t_5 inst_cell_182_62 (.BL(BL62),.BLN(BLN62),.WL(WL182));
sram_cell_6t_5 inst_cell_182_63 (.BL(BL63),.BLN(BLN63),.WL(WL182));
sram_cell_6t_5 inst_cell_182_64 (.BL(BL64),.BLN(BLN64),.WL(WL182));
sram_cell_6t_5 inst_cell_182_65 (.BL(BL65),.BLN(BLN65),.WL(WL182));
sram_cell_6t_5 inst_cell_182_66 (.BL(BL66),.BLN(BLN66),.WL(WL182));
sram_cell_6t_5 inst_cell_182_67 (.BL(BL67),.BLN(BLN67),.WL(WL182));
sram_cell_6t_5 inst_cell_182_68 (.BL(BL68),.BLN(BLN68),.WL(WL182));
sram_cell_6t_5 inst_cell_182_69 (.BL(BL69),.BLN(BLN69),.WL(WL182));
sram_cell_6t_5 inst_cell_182_70 (.BL(BL70),.BLN(BLN70),.WL(WL182));
sram_cell_6t_5 inst_cell_182_71 (.BL(BL71),.BLN(BLN71),.WL(WL182));
sram_cell_6t_5 inst_cell_182_72 (.BL(BL72),.BLN(BLN72),.WL(WL182));
sram_cell_6t_5 inst_cell_182_73 (.BL(BL73),.BLN(BLN73),.WL(WL182));
sram_cell_6t_5 inst_cell_182_74 (.BL(BL74),.BLN(BLN74),.WL(WL182));
sram_cell_6t_5 inst_cell_182_75 (.BL(BL75),.BLN(BLN75),.WL(WL182));
sram_cell_6t_5 inst_cell_182_76 (.BL(BL76),.BLN(BLN76),.WL(WL182));
sram_cell_6t_5 inst_cell_182_77 (.BL(BL77),.BLN(BLN77),.WL(WL182));
sram_cell_6t_5 inst_cell_182_78 (.BL(BL78),.BLN(BLN78),.WL(WL182));
sram_cell_6t_5 inst_cell_182_79 (.BL(BL79),.BLN(BLN79),.WL(WL182));
sram_cell_6t_5 inst_cell_182_80 (.BL(BL80),.BLN(BLN80),.WL(WL182));
sram_cell_6t_5 inst_cell_182_81 (.BL(BL81),.BLN(BLN81),.WL(WL182));
sram_cell_6t_5 inst_cell_182_82 (.BL(BL82),.BLN(BLN82),.WL(WL182));
sram_cell_6t_5 inst_cell_182_83 (.BL(BL83),.BLN(BLN83),.WL(WL182));
sram_cell_6t_5 inst_cell_182_84 (.BL(BL84),.BLN(BLN84),.WL(WL182));
sram_cell_6t_5 inst_cell_182_85 (.BL(BL85),.BLN(BLN85),.WL(WL182));
sram_cell_6t_5 inst_cell_182_86 (.BL(BL86),.BLN(BLN86),.WL(WL182));
sram_cell_6t_5 inst_cell_182_87 (.BL(BL87),.BLN(BLN87),.WL(WL182));
sram_cell_6t_5 inst_cell_182_88 (.BL(BL88),.BLN(BLN88),.WL(WL182));
sram_cell_6t_5 inst_cell_182_89 (.BL(BL89),.BLN(BLN89),.WL(WL182));
sram_cell_6t_5 inst_cell_182_90 (.BL(BL90),.BLN(BLN90),.WL(WL182));
sram_cell_6t_5 inst_cell_182_91 (.BL(BL91),.BLN(BLN91),.WL(WL182));
sram_cell_6t_5 inst_cell_182_92 (.BL(BL92),.BLN(BLN92),.WL(WL182));
sram_cell_6t_5 inst_cell_182_93 (.BL(BL93),.BLN(BLN93),.WL(WL182));
sram_cell_6t_5 inst_cell_182_94 (.BL(BL94),.BLN(BLN94),.WL(WL182));
sram_cell_6t_5 inst_cell_182_95 (.BL(BL95),.BLN(BLN95),.WL(WL182));
sram_cell_6t_5 inst_cell_182_96 (.BL(BL96),.BLN(BLN96),.WL(WL182));
sram_cell_6t_5 inst_cell_182_97 (.BL(BL97),.BLN(BLN97),.WL(WL182));
sram_cell_6t_5 inst_cell_182_98 (.BL(BL98),.BLN(BLN98),.WL(WL182));
sram_cell_6t_5 inst_cell_182_99 (.BL(BL99),.BLN(BLN99),.WL(WL182));
sram_cell_6t_5 inst_cell_182_100 (.BL(BL100),.BLN(BLN100),.WL(WL182));
sram_cell_6t_5 inst_cell_182_101 (.BL(BL101),.BLN(BLN101),.WL(WL182));
sram_cell_6t_5 inst_cell_182_102 (.BL(BL102),.BLN(BLN102),.WL(WL182));
sram_cell_6t_5 inst_cell_182_103 (.BL(BL103),.BLN(BLN103),.WL(WL182));
sram_cell_6t_5 inst_cell_182_104 (.BL(BL104),.BLN(BLN104),.WL(WL182));
sram_cell_6t_5 inst_cell_182_105 (.BL(BL105),.BLN(BLN105),.WL(WL182));
sram_cell_6t_5 inst_cell_182_106 (.BL(BL106),.BLN(BLN106),.WL(WL182));
sram_cell_6t_5 inst_cell_182_107 (.BL(BL107),.BLN(BLN107),.WL(WL182));
sram_cell_6t_5 inst_cell_182_108 (.BL(BL108),.BLN(BLN108),.WL(WL182));
sram_cell_6t_5 inst_cell_182_109 (.BL(BL109),.BLN(BLN109),.WL(WL182));
sram_cell_6t_5 inst_cell_182_110 (.BL(BL110),.BLN(BLN110),.WL(WL182));
sram_cell_6t_5 inst_cell_182_111 (.BL(BL111),.BLN(BLN111),.WL(WL182));
sram_cell_6t_5 inst_cell_182_112 (.BL(BL112),.BLN(BLN112),.WL(WL182));
sram_cell_6t_5 inst_cell_182_113 (.BL(BL113),.BLN(BLN113),.WL(WL182));
sram_cell_6t_5 inst_cell_182_114 (.BL(BL114),.BLN(BLN114),.WL(WL182));
sram_cell_6t_5 inst_cell_182_115 (.BL(BL115),.BLN(BLN115),.WL(WL182));
sram_cell_6t_5 inst_cell_182_116 (.BL(BL116),.BLN(BLN116),.WL(WL182));
sram_cell_6t_5 inst_cell_182_117 (.BL(BL117),.BLN(BLN117),.WL(WL182));
sram_cell_6t_5 inst_cell_182_118 (.BL(BL118),.BLN(BLN118),.WL(WL182));
sram_cell_6t_5 inst_cell_182_119 (.BL(BL119),.BLN(BLN119),.WL(WL182));
sram_cell_6t_5 inst_cell_182_120 (.BL(BL120),.BLN(BLN120),.WL(WL182));
sram_cell_6t_5 inst_cell_182_121 (.BL(BL121),.BLN(BLN121),.WL(WL182));
sram_cell_6t_5 inst_cell_182_122 (.BL(BL122),.BLN(BLN122),.WL(WL182));
sram_cell_6t_5 inst_cell_182_123 (.BL(BL123),.BLN(BLN123),.WL(WL182));
sram_cell_6t_5 inst_cell_182_124 (.BL(BL124),.BLN(BLN124),.WL(WL182));
sram_cell_6t_5 inst_cell_182_125 (.BL(BL125),.BLN(BLN125),.WL(WL182));
sram_cell_6t_5 inst_cell_182_126 (.BL(BL126),.BLN(BLN126),.WL(WL182));
sram_cell_6t_5 inst_cell_182_127 (.BL(BL127),.BLN(BLN127),.WL(WL182));
sram_cell_6t_5 inst_cell_183_0 (.BL(BL0),.BLN(BLN0),.WL(WL183));
sram_cell_6t_5 inst_cell_183_1 (.BL(BL1),.BLN(BLN1),.WL(WL183));
sram_cell_6t_5 inst_cell_183_2 (.BL(BL2),.BLN(BLN2),.WL(WL183));
sram_cell_6t_5 inst_cell_183_3 (.BL(BL3),.BLN(BLN3),.WL(WL183));
sram_cell_6t_5 inst_cell_183_4 (.BL(BL4),.BLN(BLN4),.WL(WL183));
sram_cell_6t_5 inst_cell_183_5 (.BL(BL5),.BLN(BLN5),.WL(WL183));
sram_cell_6t_5 inst_cell_183_6 (.BL(BL6),.BLN(BLN6),.WL(WL183));
sram_cell_6t_5 inst_cell_183_7 (.BL(BL7),.BLN(BLN7),.WL(WL183));
sram_cell_6t_5 inst_cell_183_8 (.BL(BL8),.BLN(BLN8),.WL(WL183));
sram_cell_6t_5 inst_cell_183_9 (.BL(BL9),.BLN(BLN9),.WL(WL183));
sram_cell_6t_5 inst_cell_183_10 (.BL(BL10),.BLN(BLN10),.WL(WL183));
sram_cell_6t_5 inst_cell_183_11 (.BL(BL11),.BLN(BLN11),.WL(WL183));
sram_cell_6t_5 inst_cell_183_12 (.BL(BL12),.BLN(BLN12),.WL(WL183));
sram_cell_6t_5 inst_cell_183_13 (.BL(BL13),.BLN(BLN13),.WL(WL183));
sram_cell_6t_5 inst_cell_183_14 (.BL(BL14),.BLN(BLN14),.WL(WL183));
sram_cell_6t_5 inst_cell_183_15 (.BL(BL15),.BLN(BLN15),.WL(WL183));
sram_cell_6t_5 inst_cell_183_16 (.BL(BL16),.BLN(BLN16),.WL(WL183));
sram_cell_6t_5 inst_cell_183_17 (.BL(BL17),.BLN(BLN17),.WL(WL183));
sram_cell_6t_5 inst_cell_183_18 (.BL(BL18),.BLN(BLN18),.WL(WL183));
sram_cell_6t_5 inst_cell_183_19 (.BL(BL19),.BLN(BLN19),.WL(WL183));
sram_cell_6t_5 inst_cell_183_20 (.BL(BL20),.BLN(BLN20),.WL(WL183));
sram_cell_6t_5 inst_cell_183_21 (.BL(BL21),.BLN(BLN21),.WL(WL183));
sram_cell_6t_5 inst_cell_183_22 (.BL(BL22),.BLN(BLN22),.WL(WL183));
sram_cell_6t_5 inst_cell_183_23 (.BL(BL23),.BLN(BLN23),.WL(WL183));
sram_cell_6t_5 inst_cell_183_24 (.BL(BL24),.BLN(BLN24),.WL(WL183));
sram_cell_6t_5 inst_cell_183_25 (.BL(BL25),.BLN(BLN25),.WL(WL183));
sram_cell_6t_5 inst_cell_183_26 (.BL(BL26),.BLN(BLN26),.WL(WL183));
sram_cell_6t_5 inst_cell_183_27 (.BL(BL27),.BLN(BLN27),.WL(WL183));
sram_cell_6t_5 inst_cell_183_28 (.BL(BL28),.BLN(BLN28),.WL(WL183));
sram_cell_6t_5 inst_cell_183_29 (.BL(BL29),.BLN(BLN29),.WL(WL183));
sram_cell_6t_5 inst_cell_183_30 (.BL(BL30),.BLN(BLN30),.WL(WL183));
sram_cell_6t_5 inst_cell_183_31 (.BL(BL31),.BLN(BLN31),.WL(WL183));
sram_cell_6t_5 inst_cell_183_32 (.BL(BL32),.BLN(BLN32),.WL(WL183));
sram_cell_6t_5 inst_cell_183_33 (.BL(BL33),.BLN(BLN33),.WL(WL183));
sram_cell_6t_5 inst_cell_183_34 (.BL(BL34),.BLN(BLN34),.WL(WL183));
sram_cell_6t_5 inst_cell_183_35 (.BL(BL35),.BLN(BLN35),.WL(WL183));
sram_cell_6t_5 inst_cell_183_36 (.BL(BL36),.BLN(BLN36),.WL(WL183));
sram_cell_6t_5 inst_cell_183_37 (.BL(BL37),.BLN(BLN37),.WL(WL183));
sram_cell_6t_5 inst_cell_183_38 (.BL(BL38),.BLN(BLN38),.WL(WL183));
sram_cell_6t_5 inst_cell_183_39 (.BL(BL39),.BLN(BLN39),.WL(WL183));
sram_cell_6t_5 inst_cell_183_40 (.BL(BL40),.BLN(BLN40),.WL(WL183));
sram_cell_6t_5 inst_cell_183_41 (.BL(BL41),.BLN(BLN41),.WL(WL183));
sram_cell_6t_5 inst_cell_183_42 (.BL(BL42),.BLN(BLN42),.WL(WL183));
sram_cell_6t_5 inst_cell_183_43 (.BL(BL43),.BLN(BLN43),.WL(WL183));
sram_cell_6t_5 inst_cell_183_44 (.BL(BL44),.BLN(BLN44),.WL(WL183));
sram_cell_6t_5 inst_cell_183_45 (.BL(BL45),.BLN(BLN45),.WL(WL183));
sram_cell_6t_5 inst_cell_183_46 (.BL(BL46),.BLN(BLN46),.WL(WL183));
sram_cell_6t_5 inst_cell_183_47 (.BL(BL47),.BLN(BLN47),.WL(WL183));
sram_cell_6t_5 inst_cell_183_48 (.BL(BL48),.BLN(BLN48),.WL(WL183));
sram_cell_6t_5 inst_cell_183_49 (.BL(BL49),.BLN(BLN49),.WL(WL183));
sram_cell_6t_5 inst_cell_183_50 (.BL(BL50),.BLN(BLN50),.WL(WL183));
sram_cell_6t_5 inst_cell_183_51 (.BL(BL51),.BLN(BLN51),.WL(WL183));
sram_cell_6t_5 inst_cell_183_52 (.BL(BL52),.BLN(BLN52),.WL(WL183));
sram_cell_6t_5 inst_cell_183_53 (.BL(BL53),.BLN(BLN53),.WL(WL183));
sram_cell_6t_5 inst_cell_183_54 (.BL(BL54),.BLN(BLN54),.WL(WL183));
sram_cell_6t_5 inst_cell_183_55 (.BL(BL55),.BLN(BLN55),.WL(WL183));
sram_cell_6t_5 inst_cell_183_56 (.BL(BL56),.BLN(BLN56),.WL(WL183));
sram_cell_6t_5 inst_cell_183_57 (.BL(BL57),.BLN(BLN57),.WL(WL183));
sram_cell_6t_5 inst_cell_183_58 (.BL(BL58),.BLN(BLN58),.WL(WL183));
sram_cell_6t_5 inst_cell_183_59 (.BL(BL59),.BLN(BLN59),.WL(WL183));
sram_cell_6t_5 inst_cell_183_60 (.BL(BL60),.BLN(BLN60),.WL(WL183));
sram_cell_6t_5 inst_cell_183_61 (.BL(BL61),.BLN(BLN61),.WL(WL183));
sram_cell_6t_5 inst_cell_183_62 (.BL(BL62),.BLN(BLN62),.WL(WL183));
sram_cell_6t_5 inst_cell_183_63 (.BL(BL63),.BLN(BLN63),.WL(WL183));
sram_cell_6t_5 inst_cell_183_64 (.BL(BL64),.BLN(BLN64),.WL(WL183));
sram_cell_6t_5 inst_cell_183_65 (.BL(BL65),.BLN(BLN65),.WL(WL183));
sram_cell_6t_5 inst_cell_183_66 (.BL(BL66),.BLN(BLN66),.WL(WL183));
sram_cell_6t_5 inst_cell_183_67 (.BL(BL67),.BLN(BLN67),.WL(WL183));
sram_cell_6t_5 inst_cell_183_68 (.BL(BL68),.BLN(BLN68),.WL(WL183));
sram_cell_6t_5 inst_cell_183_69 (.BL(BL69),.BLN(BLN69),.WL(WL183));
sram_cell_6t_5 inst_cell_183_70 (.BL(BL70),.BLN(BLN70),.WL(WL183));
sram_cell_6t_5 inst_cell_183_71 (.BL(BL71),.BLN(BLN71),.WL(WL183));
sram_cell_6t_5 inst_cell_183_72 (.BL(BL72),.BLN(BLN72),.WL(WL183));
sram_cell_6t_5 inst_cell_183_73 (.BL(BL73),.BLN(BLN73),.WL(WL183));
sram_cell_6t_5 inst_cell_183_74 (.BL(BL74),.BLN(BLN74),.WL(WL183));
sram_cell_6t_5 inst_cell_183_75 (.BL(BL75),.BLN(BLN75),.WL(WL183));
sram_cell_6t_5 inst_cell_183_76 (.BL(BL76),.BLN(BLN76),.WL(WL183));
sram_cell_6t_5 inst_cell_183_77 (.BL(BL77),.BLN(BLN77),.WL(WL183));
sram_cell_6t_5 inst_cell_183_78 (.BL(BL78),.BLN(BLN78),.WL(WL183));
sram_cell_6t_5 inst_cell_183_79 (.BL(BL79),.BLN(BLN79),.WL(WL183));
sram_cell_6t_5 inst_cell_183_80 (.BL(BL80),.BLN(BLN80),.WL(WL183));
sram_cell_6t_5 inst_cell_183_81 (.BL(BL81),.BLN(BLN81),.WL(WL183));
sram_cell_6t_5 inst_cell_183_82 (.BL(BL82),.BLN(BLN82),.WL(WL183));
sram_cell_6t_5 inst_cell_183_83 (.BL(BL83),.BLN(BLN83),.WL(WL183));
sram_cell_6t_5 inst_cell_183_84 (.BL(BL84),.BLN(BLN84),.WL(WL183));
sram_cell_6t_5 inst_cell_183_85 (.BL(BL85),.BLN(BLN85),.WL(WL183));
sram_cell_6t_5 inst_cell_183_86 (.BL(BL86),.BLN(BLN86),.WL(WL183));
sram_cell_6t_5 inst_cell_183_87 (.BL(BL87),.BLN(BLN87),.WL(WL183));
sram_cell_6t_5 inst_cell_183_88 (.BL(BL88),.BLN(BLN88),.WL(WL183));
sram_cell_6t_5 inst_cell_183_89 (.BL(BL89),.BLN(BLN89),.WL(WL183));
sram_cell_6t_5 inst_cell_183_90 (.BL(BL90),.BLN(BLN90),.WL(WL183));
sram_cell_6t_5 inst_cell_183_91 (.BL(BL91),.BLN(BLN91),.WL(WL183));
sram_cell_6t_5 inst_cell_183_92 (.BL(BL92),.BLN(BLN92),.WL(WL183));
sram_cell_6t_5 inst_cell_183_93 (.BL(BL93),.BLN(BLN93),.WL(WL183));
sram_cell_6t_5 inst_cell_183_94 (.BL(BL94),.BLN(BLN94),.WL(WL183));
sram_cell_6t_5 inst_cell_183_95 (.BL(BL95),.BLN(BLN95),.WL(WL183));
sram_cell_6t_5 inst_cell_183_96 (.BL(BL96),.BLN(BLN96),.WL(WL183));
sram_cell_6t_5 inst_cell_183_97 (.BL(BL97),.BLN(BLN97),.WL(WL183));
sram_cell_6t_5 inst_cell_183_98 (.BL(BL98),.BLN(BLN98),.WL(WL183));
sram_cell_6t_5 inst_cell_183_99 (.BL(BL99),.BLN(BLN99),.WL(WL183));
sram_cell_6t_5 inst_cell_183_100 (.BL(BL100),.BLN(BLN100),.WL(WL183));
sram_cell_6t_5 inst_cell_183_101 (.BL(BL101),.BLN(BLN101),.WL(WL183));
sram_cell_6t_5 inst_cell_183_102 (.BL(BL102),.BLN(BLN102),.WL(WL183));
sram_cell_6t_5 inst_cell_183_103 (.BL(BL103),.BLN(BLN103),.WL(WL183));
sram_cell_6t_5 inst_cell_183_104 (.BL(BL104),.BLN(BLN104),.WL(WL183));
sram_cell_6t_5 inst_cell_183_105 (.BL(BL105),.BLN(BLN105),.WL(WL183));
sram_cell_6t_5 inst_cell_183_106 (.BL(BL106),.BLN(BLN106),.WL(WL183));
sram_cell_6t_5 inst_cell_183_107 (.BL(BL107),.BLN(BLN107),.WL(WL183));
sram_cell_6t_5 inst_cell_183_108 (.BL(BL108),.BLN(BLN108),.WL(WL183));
sram_cell_6t_5 inst_cell_183_109 (.BL(BL109),.BLN(BLN109),.WL(WL183));
sram_cell_6t_5 inst_cell_183_110 (.BL(BL110),.BLN(BLN110),.WL(WL183));
sram_cell_6t_5 inst_cell_183_111 (.BL(BL111),.BLN(BLN111),.WL(WL183));
sram_cell_6t_5 inst_cell_183_112 (.BL(BL112),.BLN(BLN112),.WL(WL183));
sram_cell_6t_5 inst_cell_183_113 (.BL(BL113),.BLN(BLN113),.WL(WL183));
sram_cell_6t_5 inst_cell_183_114 (.BL(BL114),.BLN(BLN114),.WL(WL183));
sram_cell_6t_5 inst_cell_183_115 (.BL(BL115),.BLN(BLN115),.WL(WL183));
sram_cell_6t_5 inst_cell_183_116 (.BL(BL116),.BLN(BLN116),.WL(WL183));
sram_cell_6t_5 inst_cell_183_117 (.BL(BL117),.BLN(BLN117),.WL(WL183));
sram_cell_6t_5 inst_cell_183_118 (.BL(BL118),.BLN(BLN118),.WL(WL183));
sram_cell_6t_5 inst_cell_183_119 (.BL(BL119),.BLN(BLN119),.WL(WL183));
sram_cell_6t_5 inst_cell_183_120 (.BL(BL120),.BLN(BLN120),.WL(WL183));
sram_cell_6t_5 inst_cell_183_121 (.BL(BL121),.BLN(BLN121),.WL(WL183));
sram_cell_6t_5 inst_cell_183_122 (.BL(BL122),.BLN(BLN122),.WL(WL183));
sram_cell_6t_5 inst_cell_183_123 (.BL(BL123),.BLN(BLN123),.WL(WL183));
sram_cell_6t_5 inst_cell_183_124 (.BL(BL124),.BLN(BLN124),.WL(WL183));
sram_cell_6t_5 inst_cell_183_125 (.BL(BL125),.BLN(BLN125),.WL(WL183));
sram_cell_6t_5 inst_cell_183_126 (.BL(BL126),.BLN(BLN126),.WL(WL183));
sram_cell_6t_5 inst_cell_183_127 (.BL(BL127),.BLN(BLN127),.WL(WL183));
sram_cell_6t_5 inst_cell_184_0 (.BL(BL0),.BLN(BLN0),.WL(WL184));
sram_cell_6t_5 inst_cell_184_1 (.BL(BL1),.BLN(BLN1),.WL(WL184));
sram_cell_6t_5 inst_cell_184_2 (.BL(BL2),.BLN(BLN2),.WL(WL184));
sram_cell_6t_5 inst_cell_184_3 (.BL(BL3),.BLN(BLN3),.WL(WL184));
sram_cell_6t_5 inst_cell_184_4 (.BL(BL4),.BLN(BLN4),.WL(WL184));
sram_cell_6t_5 inst_cell_184_5 (.BL(BL5),.BLN(BLN5),.WL(WL184));
sram_cell_6t_5 inst_cell_184_6 (.BL(BL6),.BLN(BLN6),.WL(WL184));
sram_cell_6t_5 inst_cell_184_7 (.BL(BL7),.BLN(BLN7),.WL(WL184));
sram_cell_6t_5 inst_cell_184_8 (.BL(BL8),.BLN(BLN8),.WL(WL184));
sram_cell_6t_5 inst_cell_184_9 (.BL(BL9),.BLN(BLN9),.WL(WL184));
sram_cell_6t_5 inst_cell_184_10 (.BL(BL10),.BLN(BLN10),.WL(WL184));
sram_cell_6t_5 inst_cell_184_11 (.BL(BL11),.BLN(BLN11),.WL(WL184));
sram_cell_6t_5 inst_cell_184_12 (.BL(BL12),.BLN(BLN12),.WL(WL184));
sram_cell_6t_5 inst_cell_184_13 (.BL(BL13),.BLN(BLN13),.WL(WL184));
sram_cell_6t_5 inst_cell_184_14 (.BL(BL14),.BLN(BLN14),.WL(WL184));
sram_cell_6t_5 inst_cell_184_15 (.BL(BL15),.BLN(BLN15),.WL(WL184));
sram_cell_6t_5 inst_cell_184_16 (.BL(BL16),.BLN(BLN16),.WL(WL184));
sram_cell_6t_5 inst_cell_184_17 (.BL(BL17),.BLN(BLN17),.WL(WL184));
sram_cell_6t_5 inst_cell_184_18 (.BL(BL18),.BLN(BLN18),.WL(WL184));
sram_cell_6t_5 inst_cell_184_19 (.BL(BL19),.BLN(BLN19),.WL(WL184));
sram_cell_6t_5 inst_cell_184_20 (.BL(BL20),.BLN(BLN20),.WL(WL184));
sram_cell_6t_5 inst_cell_184_21 (.BL(BL21),.BLN(BLN21),.WL(WL184));
sram_cell_6t_5 inst_cell_184_22 (.BL(BL22),.BLN(BLN22),.WL(WL184));
sram_cell_6t_5 inst_cell_184_23 (.BL(BL23),.BLN(BLN23),.WL(WL184));
sram_cell_6t_5 inst_cell_184_24 (.BL(BL24),.BLN(BLN24),.WL(WL184));
sram_cell_6t_5 inst_cell_184_25 (.BL(BL25),.BLN(BLN25),.WL(WL184));
sram_cell_6t_5 inst_cell_184_26 (.BL(BL26),.BLN(BLN26),.WL(WL184));
sram_cell_6t_5 inst_cell_184_27 (.BL(BL27),.BLN(BLN27),.WL(WL184));
sram_cell_6t_5 inst_cell_184_28 (.BL(BL28),.BLN(BLN28),.WL(WL184));
sram_cell_6t_5 inst_cell_184_29 (.BL(BL29),.BLN(BLN29),.WL(WL184));
sram_cell_6t_5 inst_cell_184_30 (.BL(BL30),.BLN(BLN30),.WL(WL184));
sram_cell_6t_5 inst_cell_184_31 (.BL(BL31),.BLN(BLN31),.WL(WL184));
sram_cell_6t_5 inst_cell_184_32 (.BL(BL32),.BLN(BLN32),.WL(WL184));
sram_cell_6t_5 inst_cell_184_33 (.BL(BL33),.BLN(BLN33),.WL(WL184));
sram_cell_6t_5 inst_cell_184_34 (.BL(BL34),.BLN(BLN34),.WL(WL184));
sram_cell_6t_5 inst_cell_184_35 (.BL(BL35),.BLN(BLN35),.WL(WL184));
sram_cell_6t_5 inst_cell_184_36 (.BL(BL36),.BLN(BLN36),.WL(WL184));
sram_cell_6t_5 inst_cell_184_37 (.BL(BL37),.BLN(BLN37),.WL(WL184));
sram_cell_6t_5 inst_cell_184_38 (.BL(BL38),.BLN(BLN38),.WL(WL184));
sram_cell_6t_5 inst_cell_184_39 (.BL(BL39),.BLN(BLN39),.WL(WL184));
sram_cell_6t_5 inst_cell_184_40 (.BL(BL40),.BLN(BLN40),.WL(WL184));
sram_cell_6t_5 inst_cell_184_41 (.BL(BL41),.BLN(BLN41),.WL(WL184));
sram_cell_6t_5 inst_cell_184_42 (.BL(BL42),.BLN(BLN42),.WL(WL184));
sram_cell_6t_5 inst_cell_184_43 (.BL(BL43),.BLN(BLN43),.WL(WL184));
sram_cell_6t_5 inst_cell_184_44 (.BL(BL44),.BLN(BLN44),.WL(WL184));
sram_cell_6t_5 inst_cell_184_45 (.BL(BL45),.BLN(BLN45),.WL(WL184));
sram_cell_6t_5 inst_cell_184_46 (.BL(BL46),.BLN(BLN46),.WL(WL184));
sram_cell_6t_5 inst_cell_184_47 (.BL(BL47),.BLN(BLN47),.WL(WL184));
sram_cell_6t_5 inst_cell_184_48 (.BL(BL48),.BLN(BLN48),.WL(WL184));
sram_cell_6t_5 inst_cell_184_49 (.BL(BL49),.BLN(BLN49),.WL(WL184));
sram_cell_6t_5 inst_cell_184_50 (.BL(BL50),.BLN(BLN50),.WL(WL184));
sram_cell_6t_5 inst_cell_184_51 (.BL(BL51),.BLN(BLN51),.WL(WL184));
sram_cell_6t_5 inst_cell_184_52 (.BL(BL52),.BLN(BLN52),.WL(WL184));
sram_cell_6t_5 inst_cell_184_53 (.BL(BL53),.BLN(BLN53),.WL(WL184));
sram_cell_6t_5 inst_cell_184_54 (.BL(BL54),.BLN(BLN54),.WL(WL184));
sram_cell_6t_5 inst_cell_184_55 (.BL(BL55),.BLN(BLN55),.WL(WL184));
sram_cell_6t_5 inst_cell_184_56 (.BL(BL56),.BLN(BLN56),.WL(WL184));
sram_cell_6t_5 inst_cell_184_57 (.BL(BL57),.BLN(BLN57),.WL(WL184));
sram_cell_6t_5 inst_cell_184_58 (.BL(BL58),.BLN(BLN58),.WL(WL184));
sram_cell_6t_5 inst_cell_184_59 (.BL(BL59),.BLN(BLN59),.WL(WL184));
sram_cell_6t_5 inst_cell_184_60 (.BL(BL60),.BLN(BLN60),.WL(WL184));
sram_cell_6t_5 inst_cell_184_61 (.BL(BL61),.BLN(BLN61),.WL(WL184));
sram_cell_6t_5 inst_cell_184_62 (.BL(BL62),.BLN(BLN62),.WL(WL184));
sram_cell_6t_5 inst_cell_184_63 (.BL(BL63),.BLN(BLN63),.WL(WL184));
sram_cell_6t_5 inst_cell_184_64 (.BL(BL64),.BLN(BLN64),.WL(WL184));
sram_cell_6t_5 inst_cell_184_65 (.BL(BL65),.BLN(BLN65),.WL(WL184));
sram_cell_6t_5 inst_cell_184_66 (.BL(BL66),.BLN(BLN66),.WL(WL184));
sram_cell_6t_5 inst_cell_184_67 (.BL(BL67),.BLN(BLN67),.WL(WL184));
sram_cell_6t_5 inst_cell_184_68 (.BL(BL68),.BLN(BLN68),.WL(WL184));
sram_cell_6t_5 inst_cell_184_69 (.BL(BL69),.BLN(BLN69),.WL(WL184));
sram_cell_6t_5 inst_cell_184_70 (.BL(BL70),.BLN(BLN70),.WL(WL184));
sram_cell_6t_5 inst_cell_184_71 (.BL(BL71),.BLN(BLN71),.WL(WL184));
sram_cell_6t_5 inst_cell_184_72 (.BL(BL72),.BLN(BLN72),.WL(WL184));
sram_cell_6t_5 inst_cell_184_73 (.BL(BL73),.BLN(BLN73),.WL(WL184));
sram_cell_6t_5 inst_cell_184_74 (.BL(BL74),.BLN(BLN74),.WL(WL184));
sram_cell_6t_5 inst_cell_184_75 (.BL(BL75),.BLN(BLN75),.WL(WL184));
sram_cell_6t_5 inst_cell_184_76 (.BL(BL76),.BLN(BLN76),.WL(WL184));
sram_cell_6t_5 inst_cell_184_77 (.BL(BL77),.BLN(BLN77),.WL(WL184));
sram_cell_6t_5 inst_cell_184_78 (.BL(BL78),.BLN(BLN78),.WL(WL184));
sram_cell_6t_5 inst_cell_184_79 (.BL(BL79),.BLN(BLN79),.WL(WL184));
sram_cell_6t_5 inst_cell_184_80 (.BL(BL80),.BLN(BLN80),.WL(WL184));
sram_cell_6t_5 inst_cell_184_81 (.BL(BL81),.BLN(BLN81),.WL(WL184));
sram_cell_6t_5 inst_cell_184_82 (.BL(BL82),.BLN(BLN82),.WL(WL184));
sram_cell_6t_5 inst_cell_184_83 (.BL(BL83),.BLN(BLN83),.WL(WL184));
sram_cell_6t_5 inst_cell_184_84 (.BL(BL84),.BLN(BLN84),.WL(WL184));
sram_cell_6t_5 inst_cell_184_85 (.BL(BL85),.BLN(BLN85),.WL(WL184));
sram_cell_6t_5 inst_cell_184_86 (.BL(BL86),.BLN(BLN86),.WL(WL184));
sram_cell_6t_5 inst_cell_184_87 (.BL(BL87),.BLN(BLN87),.WL(WL184));
sram_cell_6t_5 inst_cell_184_88 (.BL(BL88),.BLN(BLN88),.WL(WL184));
sram_cell_6t_5 inst_cell_184_89 (.BL(BL89),.BLN(BLN89),.WL(WL184));
sram_cell_6t_5 inst_cell_184_90 (.BL(BL90),.BLN(BLN90),.WL(WL184));
sram_cell_6t_5 inst_cell_184_91 (.BL(BL91),.BLN(BLN91),.WL(WL184));
sram_cell_6t_5 inst_cell_184_92 (.BL(BL92),.BLN(BLN92),.WL(WL184));
sram_cell_6t_5 inst_cell_184_93 (.BL(BL93),.BLN(BLN93),.WL(WL184));
sram_cell_6t_5 inst_cell_184_94 (.BL(BL94),.BLN(BLN94),.WL(WL184));
sram_cell_6t_5 inst_cell_184_95 (.BL(BL95),.BLN(BLN95),.WL(WL184));
sram_cell_6t_5 inst_cell_184_96 (.BL(BL96),.BLN(BLN96),.WL(WL184));
sram_cell_6t_5 inst_cell_184_97 (.BL(BL97),.BLN(BLN97),.WL(WL184));
sram_cell_6t_5 inst_cell_184_98 (.BL(BL98),.BLN(BLN98),.WL(WL184));
sram_cell_6t_5 inst_cell_184_99 (.BL(BL99),.BLN(BLN99),.WL(WL184));
sram_cell_6t_5 inst_cell_184_100 (.BL(BL100),.BLN(BLN100),.WL(WL184));
sram_cell_6t_5 inst_cell_184_101 (.BL(BL101),.BLN(BLN101),.WL(WL184));
sram_cell_6t_5 inst_cell_184_102 (.BL(BL102),.BLN(BLN102),.WL(WL184));
sram_cell_6t_5 inst_cell_184_103 (.BL(BL103),.BLN(BLN103),.WL(WL184));
sram_cell_6t_5 inst_cell_184_104 (.BL(BL104),.BLN(BLN104),.WL(WL184));
sram_cell_6t_5 inst_cell_184_105 (.BL(BL105),.BLN(BLN105),.WL(WL184));
sram_cell_6t_5 inst_cell_184_106 (.BL(BL106),.BLN(BLN106),.WL(WL184));
sram_cell_6t_5 inst_cell_184_107 (.BL(BL107),.BLN(BLN107),.WL(WL184));
sram_cell_6t_5 inst_cell_184_108 (.BL(BL108),.BLN(BLN108),.WL(WL184));
sram_cell_6t_5 inst_cell_184_109 (.BL(BL109),.BLN(BLN109),.WL(WL184));
sram_cell_6t_5 inst_cell_184_110 (.BL(BL110),.BLN(BLN110),.WL(WL184));
sram_cell_6t_5 inst_cell_184_111 (.BL(BL111),.BLN(BLN111),.WL(WL184));
sram_cell_6t_5 inst_cell_184_112 (.BL(BL112),.BLN(BLN112),.WL(WL184));
sram_cell_6t_5 inst_cell_184_113 (.BL(BL113),.BLN(BLN113),.WL(WL184));
sram_cell_6t_5 inst_cell_184_114 (.BL(BL114),.BLN(BLN114),.WL(WL184));
sram_cell_6t_5 inst_cell_184_115 (.BL(BL115),.BLN(BLN115),.WL(WL184));
sram_cell_6t_5 inst_cell_184_116 (.BL(BL116),.BLN(BLN116),.WL(WL184));
sram_cell_6t_5 inst_cell_184_117 (.BL(BL117),.BLN(BLN117),.WL(WL184));
sram_cell_6t_5 inst_cell_184_118 (.BL(BL118),.BLN(BLN118),.WL(WL184));
sram_cell_6t_5 inst_cell_184_119 (.BL(BL119),.BLN(BLN119),.WL(WL184));
sram_cell_6t_5 inst_cell_184_120 (.BL(BL120),.BLN(BLN120),.WL(WL184));
sram_cell_6t_5 inst_cell_184_121 (.BL(BL121),.BLN(BLN121),.WL(WL184));
sram_cell_6t_5 inst_cell_184_122 (.BL(BL122),.BLN(BLN122),.WL(WL184));
sram_cell_6t_5 inst_cell_184_123 (.BL(BL123),.BLN(BLN123),.WL(WL184));
sram_cell_6t_5 inst_cell_184_124 (.BL(BL124),.BLN(BLN124),.WL(WL184));
sram_cell_6t_5 inst_cell_184_125 (.BL(BL125),.BLN(BLN125),.WL(WL184));
sram_cell_6t_5 inst_cell_184_126 (.BL(BL126),.BLN(BLN126),.WL(WL184));
sram_cell_6t_5 inst_cell_184_127 (.BL(BL127),.BLN(BLN127),.WL(WL184));
sram_cell_6t_5 inst_cell_185_0 (.BL(BL0),.BLN(BLN0),.WL(WL185));
sram_cell_6t_5 inst_cell_185_1 (.BL(BL1),.BLN(BLN1),.WL(WL185));
sram_cell_6t_5 inst_cell_185_2 (.BL(BL2),.BLN(BLN2),.WL(WL185));
sram_cell_6t_5 inst_cell_185_3 (.BL(BL3),.BLN(BLN3),.WL(WL185));
sram_cell_6t_5 inst_cell_185_4 (.BL(BL4),.BLN(BLN4),.WL(WL185));
sram_cell_6t_5 inst_cell_185_5 (.BL(BL5),.BLN(BLN5),.WL(WL185));
sram_cell_6t_5 inst_cell_185_6 (.BL(BL6),.BLN(BLN6),.WL(WL185));
sram_cell_6t_5 inst_cell_185_7 (.BL(BL7),.BLN(BLN7),.WL(WL185));
sram_cell_6t_5 inst_cell_185_8 (.BL(BL8),.BLN(BLN8),.WL(WL185));
sram_cell_6t_5 inst_cell_185_9 (.BL(BL9),.BLN(BLN9),.WL(WL185));
sram_cell_6t_5 inst_cell_185_10 (.BL(BL10),.BLN(BLN10),.WL(WL185));
sram_cell_6t_5 inst_cell_185_11 (.BL(BL11),.BLN(BLN11),.WL(WL185));
sram_cell_6t_5 inst_cell_185_12 (.BL(BL12),.BLN(BLN12),.WL(WL185));
sram_cell_6t_5 inst_cell_185_13 (.BL(BL13),.BLN(BLN13),.WL(WL185));
sram_cell_6t_5 inst_cell_185_14 (.BL(BL14),.BLN(BLN14),.WL(WL185));
sram_cell_6t_5 inst_cell_185_15 (.BL(BL15),.BLN(BLN15),.WL(WL185));
sram_cell_6t_5 inst_cell_185_16 (.BL(BL16),.BLN(BLN16),.WL(WL185));
sram_cell_6t_5 inst_cell_185_17 (.BL(BL17),.BLN(BLN17),.WL(WL185));
sram_cell_6t_5 inst_cell_185_18 (.BL(BL18),.BLN(BLN18),.WL(WL185));
sram_cell_6t_5 inst_cell_185_19 (.BL(BL19),.BLN(BLN19),.WL(WL185));
sram_cell_6t_5 inst_cell_185_20 (.BL(BL20),.BLN(BLN20),.WL(WL185));
sram_cell_6t_5 inst_cell_185_21 (.BL(BL21),.BLN(BLN21),.WL(WL185));
sram_cell_6t_5 inst_cell_185_22 (.BL(BL22),.BLN(BLN22),.WL(WL185));
sram_cell_6t_5 inst_cell_185_23 (.BL(BL23),.BLN(BLN23),.WL(WL185));
sram_cell_6t_5 inst_cell_185_24 (.BL(BL24),.BLN(BLN24),.WL(WL185));
sram_cell_6t_5 inst_cell_185_25 (.BL(BL25),.BLN(BLN25),.WL(WL185));
sram_cell_6t_5 inst_cell_185_26 (.BL(BL26),.BLN(BLN26),.WL(WL185));
sram_cell_6t_5 inst_cell_185_27 (.BL(BL27),.BLN(BLN27),.WL(WL185));
sram_cell_6t_5 inst_cell_185_28 (.BL(BL28),.BLN(BLN28),.WL(WL185));
sram_cell_6t_5 inst_cell_185_29 (.BL(BL29),.BLN(BLN29),.WL(WL185));
sram_cell_6t_5 inst_cell_185_30 (.BL(BL30),.BLN(BLN30),.WL(WL185));
sram_cell_6t_5 inst_cell_185_31 (.BL(BL31),.BLN(BLN31),.WL(WL185));
sram_cell_6t_5 inst_cell_185_32 (.BL(BL32),.BLN(BLN32),.WL(WL185));
sram_cell_6t_5 inst_cell_185_33 (.BL(BL33),.BLN(BLN33),.WL(WL185));
sram_cell_6t_5 inst_cell_185_34 (.BL(BL34),.BLN(BLN34),.WL(WL185));
sram_cell_6t_5 inst_cell_185_35 (.BL(BL35),.BLN(BLN35),.WL(WL185));
sram_cell_6t_5 inst_cell_185_36 (.BL(BL36),.BLN(BLN36),.WL(WL185));
sram_cell_6t_5 inst_cell_185_37 (.BL(BL37),.BLN(BLN37),.WL(WL185));
sram_cell_6t_5 inst_cell_185_38 (.BL(BL38),.BLN(BLN38),.WL(WL185));
sram_cell_6t_5 inst_cell_185_39 (.BL(BL39),.BLN(BLN39),.WL(WL185));
sram_cell_6t_5 inst_cell_185_40 (.BL(BL40),.BLN(BLN40),.WL(WL185));
sram_cell_6t_5 inst_cell_185_41 (.BL(BL41),.BLN(BLN41),.WL(WL185));
sram_cell_6t_5 inst_cell_185_42 (.BL(BL42),.BLN(BLN42),.WL(WL185));
sram_cell_6t_5 inst_cell_185_43 (.BL(BL43),.BLN(BLN43),.WL(WL185));
sram_cell_6t_5 inst_cell_185_44 (.BL(BL44),.BLN(BLN44),.WL(WL185));
sram_cell_6t_5 inst_cell_185_45 (.BL(BL45),.BLN(BLN45),.WL(WL185));
sram_cell_6t_5 inst_cell_185_46 (.BL(BL46),.BLN(BLN46),.WL(WL185));
sram_cell_6t_5 inst_cell_185_47 (.BL(BL47),.BLN(BLN47),.WL(WL185));
sram_cell_6t_5 inst_cell_185_48 (.BL(BL48),.BLN(BLN48),.WL(WL185));
sram_cell_6t_5 inst_cell_185_49 (.BL(BL49),.BLN(BLN49),.WL(WL185));
sram_cell_6t_5 inst_cell_185_50 (.BL(BL50),.BLN(BLN50),.WL(WL185));
sram_cell_6t_5 inst_cell_185_51 (.BL(BL51),.BLN(BLN51),.WL(WL185));
sram_cell_6t_5 inst_cell_185_52 (.BL(BL52),.BLN(BLN52),.WL(WL185));
sram_cell_6t_5 inst_cell_185_53 (.BL(BL53),.BLN(BLN53),.WL(WL185));
sram_cell_6t_5 inst_cell_185_54 (.BL(BL54),.BLN(BLN54),.WL(WL185));
sram_cell_6t_5 inst_cell_185_55 (.BL(BL55),.BLN(BLN55),.WL(WL185));
sram_cell_6t_5 inst_cell_185_56 (.BL(BL56),.BLN(BLN56),.WL(WL185));
sram_cell_6t_5 inst_cell_185_57 (.BL(BL57),.BLN(BLN57),.WL(WL185));
sram_cell_6t_5 inst_cell_185_58 (.BL(BL58),.BLN(BLN58),.WL(WL185));
sram_cell_6t_5 inst_cell_185_59 (.BL(BL59),.BLN(BLN59),.WL(WL185));
sram_cell_6t_5 inst_cell_185_60 (.BL(BL60),.BLN(BLN60),.WL(WL185));
sram_cell_6t_5 inst_cell_185_61 (.BL(BL61),.BLN(BLN61),.WL(WL185));
sram_cell_6t_5 inst_cell_185_62 (.BL(BL62),.BLN(BLN62),.WL(WL185));
sram_cell_6t_5 inst_cell_185_63 (.BL(BL63),.BLN(BLN63),.WL(WL185));
sram_cell_6t_5 inst_cell_185_64 (.BL(BL64),.BLN(BLN64),.WL(WL185));
sram_cell_6t_5 inst_cell_185_65 (.BL(BL65),.BLN(BLN65),.WL(WL185));
sram_cell_6t_5 inst_cell_185_66 (.BL(BL66),.BLN(BLN66),.WL(WL185));
sram_cell_6t_5 inst_cell_185_67 (.BL(BL67),.BLN(BLN67),.WL(WL185));
sram_cell_6t_5 inst_cell_185_68 (.BL(BL68),.BLN(BLN68),.WL(WL185));
sram_cell_6t_5 inst_cell_185_69 (.BL(BL69),.BLN(BLN69),.WL(WL185));
sram_cell_6t_5 inst_cell_185_70 (.BL(BL70),.BLN(BLN70),.WL(WL185));
sram_cell_6t_5 inst_cell_185_71 (.BL(BL71),.BLN(BLN71),.WL(WL185));
sram_cell_6t_5 inst_cell_185_72 (.BL(BL72),.BLN(BLN72),.WL(WL185));
sram_cell_6t_5 inst_cell_185_73 (.BL(BL73),.BLN(BLN73),.WL(WL185));
sram_cell_6t_5 inst_cell_185_74 (.BL(BL74),.BLN(BLN74),.WL(WL185));
sram_cell_6t_5 inst_cell_185_75 (.BL(BL75),.BLN(BLN75),.WL(WL185));
sram_cell_6t_5 inst_cell_185_76 (.BL(BL76),.BLN(BLN76),.WL(WL185));
sram_cell_6t_5 inst_cell_185_77 (.BL(BL77),.BLN(BLN77),.WL(WL185));
sram_cell_6t_5 inst_cell_185_78 (.BL(BL78),.BLN(BLN78),.WL(WL185));
sram_cell_6t_5 inst_cell_185_79 (.BL(BL79),.BLN(BLN79),.WL(WL185));
sram_cell_6t_5 inst_cell_185_80 (.BL(BL80),.BLN(BLN80),.WL(WL185));
sram_cell_6t_5 inst_cell_185_81 (.BL(BL81),.BLN(BLN81),.WL(WL185));
sram_cell_6t_5 inst_cell_185_82 (.BL(BL82),.BLN(BLN82),.WL(WL185));
sram_cell_6t_5 inst_cell_185_83 (.BL(BL83),.BLN(BLN83),.WL(WL185));
sram_cell_6t_5 inst_cell_185_84 (.BL(BL84),.BLN(BLN84),.WL(WL185));
sram_cell_6t_5 inst_cell_185_85 (.BL(BL85),.BLN(BLN85),.WL(WL185));
sram_cell_6t_5 inst_cell_185_86 (.BL(BL86),.BLN(BLN86),.WL(WL185));
sram_cell_6t_5 inst_cell_185_87 (.BL(BL87),.BLN(BLN87),.WL(WL185));
sram_cell_6t_5 inst_cell_185_88 (.BL(BL88),.BLN(BLN88),.WL(WL185));
sram_cell_6t_5 inst_cell_185_89 (.BL(BL89),.BLN(BLN89),.WL(WL185));
sram_cell_6t_5 inst_cell_185_90 (.BL(BL90),.BLN(BLN90),.WL(WL185));
sram_cell_6t_5 inst_cell_185_91 (.BL(BL91),.BLN(BLN91),.WL(WL185));
sram_cell_6t_5 inst_cell_185_92 (.BL(BL92),.BLN(BLN92),.WL(WL185));
sram_cell_6t_5 inst_cell_185_93 (.BL(BL93),.BLN(BLN93),.WL(WL185));
sram_cell_6t_5 inst_cell_185_94 (.BL(BL94),.BLN(BLN94),.WL(WL185));
sram_cell_6t_5 inst_cell_185_95 (.BL(BL95),.BLN(BLN95),.WL(WL185));
sram_cell_6t_5 inst_cell_185_96 (.BL(BL96),.BLN(BLN96),.WL(WL185));
sram_cell_6t_5 inst_cell_185_97 (.BL(BL97),.BLN(BLN97),.WL(WL185));
sram_cell_6t_5 inst_cell_185_98 (.BL(BL98),.BLN(BLN98),.WL(WL185));
sram_cell_6t_5 inst_cell_185_99 (.BL(BL99),.BLN(BLN99),.WL(WL185));
sram_cell_6t_5 inst_cell_185_100 (.BL(BL100),.BLN(BLN100),.WL(WL185));
sram_cell_6t_5 inst_cell_185_101 (.BL(BL101),.BLN(BLN101),.WL(WL185));
sram_cell_6t_5 inst_cell_185_102 (.BL(BL102),.BLN(BLN102),.WL(WL185));
sram_cell_6t_5 inst_cell_185_103 (.BL(BL103),.BLN(BLN103),.WL(WL185));
sram_cell_6t_5 inst_cell_185_104 (.BL(BL104),.BLN(BLN104),.WL(WL185));
sram_cell_6t_5 inst_cell_185_105 (.BL(BL105),.BLN(BLN105),.WL(WL185));
sram_cell_6t_5 inst_cell_185_106 (.BL(BL106),.BLN(BLN106),.WL(WL185));
sram_cell_6t_5 inst_cell_185_107 (.BL(BL107),.BLN(BLN107),.WL(WL185));
sram_cell_6t_5 inst_cell_185_108 (.BL(BL108),.BLN(BLN108),.WL(WL185));
sram_cell_6t_5 inst_cell_185_109 (.BL(BL109),.BLN(BLN109),.WL(WL185));
sram_cell_6t_5 inst_cell_185_110 (.BL(BL110),.BLN(BLN110),.WL(WL185));
sram_cell_6t_5 inst_cell_185_111 (.BL(BL111),.BLN(BLN111),.WL(WL185));
sram_cell_6t_5 inst_cell_185_112 (.BL(BL112),.BLN(BLN112),.WL(WL185));
sram_cell_6t_5 inst_cell_185_113 (.BL(BL113),.BLN(BLN113),.WL(WL185));
sram_cell_6t_5 inst_cell_185_114 (.BL(BL114),.BLN(BLN114),.WL(WL185));
sram_cell_6t_5 inst_cell_185_115 (.BL(BL115),.BLN(BLN115),.WL(WL185));
sram_cell_6t_5 inst_cell_185_116 (.BL(BL116),.BLN(BLN116),.WL(WL185));
sram_cell_6t_5 inst_cell_185_117 (.BL(BL117),.BLN(BLN117),.WL(WL185));
sram_cell_6t_5 inst_cell_185_118 (.BL(BL118),.BLN(BLN118),.WL(WL185));
sram_cell_6t_5 inst_cell_185_119 (.BL(BL119),.BLN(BLN119),.WL(WL185));
sram_cell_6t_5 inst_cell_185_120 (.BL(BL120),.BLN(BLN120),.WL(WL185));
sram_cell_6t_5 inst_cell_185_121 (.BL(BL121),.BLN(BLN121),.WL(WL185));
sram_cell_6t_5 inst_cell_185_122 (.BL(BL122),.BLN(BLN122),.WL(WL185));
sram_cell_6t_5 inst_cell_185_123 (.BL(BL123),.BLN(BLN123),.WL(WL185));
sram_cell_6t_5 inst_cell_185_124 (.BL(BL124),.BLN(BLN124),.WL(WL185));
sram_cell_6t_5 inst_cell_185_125 (.BL(BL125),.BLN(BLN125),.WL(WL185));
sram_cell_6t_5 inst_cell_185_126 (.BL(BL126),.BLN(BLN126),.WL(WL185));
sram_cell_6t_5 inst_cell_185_127 (.BL(BL127),.BLN(BLN127),.WL(WL185));
sram_cell_6t_5 inst_cell_186_0 (.BL(BL0),.BLN(BLN0),.WL(WL186));
sram_cell_6t_5 inst_cell_186_1 (.BL(BL1),.BLN(BLN1),.WL(WL186));
sram_cell_6t_5 inst_cell_186_2 (.BL(BL2),.BLN(BLN2),.WL(WL186));
sram_cell_6t_5 inst_cell_186_3 (.BL(BL3),.BLN(BLN3),.WL(WL186));
sram_cell_6t_5 inst_cell_186_4 (.BL(BL4),.BLN(BLN4),.WL(WL186));
sram_cell_6t_5 inst_cell_186_5 (.BL(BL5),.BLN(BLN5),.WL(WL186));
sram_cell_6t_5 inst_cell_186_6 (.BL(BL6),.BLN(BLN6),.WL(WL186));
sram_cell_6t_5 inst_cell_186_7 (.BL(BL7),.BLN(BLN7),.WL(WL186));
sram_cell_6t_5 inst_cell_186_8 (.BL(BL8),.BLN(BLN8),.WL(WL186));
sram_cell_6t_5 inst_cell_186_9 (.BL(BL9),.BLN(BLN9),.WL(WL186));
sram_cell_6t_5 inst_cell_186_10 (.BL(BL10),.BLN(BLN10),.WL(WL186));
sram_cell_6t_5 inst_cell_186_11 (.BL(BL11),.BLN(BLN11),.WL(WL186));
sram_cell_6t_5 inst_cell_186_12 (.BL(BL12),.BLN(BLN12),.WL(WL186));
sram_cell_6t_5 inst_cell_186_13 (.BL(BL13),.BLN(BLN13),.WL(WL186));
sram_cell_6t_5 inst_cell_186_14 (.BL(BL14),.BLN(BLN14),.WL(WL186));
sram_cell_6t_5 inst_cell_186_15 (.BL(BL15),.BLN(BLN15),.WL(WL186));
sram_cell_6t_5 inst_cell_186_16 (.BL(BL16),.BLN(BLN16),.WL(WL186));
sram_cell_6t_5 inst_cell_186_17 (.BL(BL17),.BLN(BLN17),.WL(WL186));
sram_cell_6t_5 inst_cell_186_18 (.BL(BL18),.BLN(BLN18),.WL(WL186));
sram_cell_6t_5 inst_cell_186_19 (.BL(BL19),.BLN(BLN19),.WL(WL186));
sram_cell_6t_5 inst_cell_186_20 (.BL(BL20),.BLN(BLN20),.WL(WL186));
sram_cell_6t_5 inst_cell_186_21 (.BL(BL21),.BLN(BLN21),.WL(WL186));
sram_cell_6t_5 inst_cell_186_22 (.BL(BL22),.BLN(BLN22),.WL(WL186));
sram_cell_6t_5 inst_cell_186_23 (.BL(BL23),.BLN(BLN23),.WL(WL186));
sram_cell_6t_5 inst_cell_186_24 (.BL(BL24),.BLN(BLN24),.WL(WL186));
sram_cell_6t_5 inst_cell_186_25 (.BL(BL25),.BLN(BLN25),.WL(WL186));
sram_cell_6t_5 inst_cell_186_26 (.BL(BL26),.BLN(BLN26),.WL(WL186));
sram_cell_6t_5 inst_cell_186_27 (.BL(BL27),.BLN(BLN27),.WL(WL186));
sram_cell_6t_5 inst_cell_186_28 (.BL(BL28),.BLN(BLN28),.WL(WL186));
sram_cell_6t_5 inst_cell_186_29 (.BL(BL29),.BLN(BLN29),.WL(WL186));
sram_cell_6t_5 inst_cell_186_30 (.BL(BL30),.BLN(BLN30),.WL(WL186));
sram_cell_6t_5 inst_cell_186_31 (.BL(BL31),.BLN(BLN31),.WL(WL186));
sram_cell_6t_5 inst_cell_186_32 (.BL(BL32),.BLN(BLN32),.WL(WL186));
sram_cell_6t_5 inst_cell_186_33 (.BL(BL33),.BLN(BLN33),.WL(WL186));
sram_cell_6t_5 inst_cell_186_34 (.BL(BL34),.BLN(BLN34),.WL(WL186));
sram_cell_6t_5 inst_cell_186_35 (.BL(BL35),.BLN(BLN35),.WL(WL186));
sram_cell_6t_5 inst_cell_186_36 (.BL(BL36),.BLN(BLN36),.WL(WL186));
sram_cell_6t_5 inst_cell_186_37 (.BL(BL37),.BLN(BLN37),.WL(WL186));
sram_cell_6t_5 inst_cell_186_38 (.BL(BL38),.BLN(BLN38),.WL(WL186));
sram_cell_6t_5 inst_cell_186_39 (.BL(BL39),.BLN(BLN39),.WL(WL186));
sram_cell_6t_5 inst_cell_186_40 (.BL(BL40),.BLN(BLN40),.WL(WL186));
sram_cell_6t_5 inst_cell_186_41 (.BL(BL41),.BLN(BLN41),.WL(WL186));
sram_cell_6t_5 inst_cell_186_42 (.BL(BL42),.BLN(BLN42),.WL(WL186));
sram_cell_6t_5 inst_cell_186_43 (.BL(BL43),.BLN(BLN43),.WL(WL186));
sram_cell_6t_5 inst_cell_186_44 (.BL(BL44),.BLN(BLN44),.WL(WL186));
sram_cell_6t_5 inst_cell_186_45 (.BL(BL45),.BLN(BLN45),.WL(WL186));
sram_cell_6t_5 inst_cell_186_46 (.BL(BL46),.BLN(BLN46),.WL(WL186));
sram_cell_6t_5 inst_cell_186_47 (.BL(BL47),.BLN(BLN47),.WL(WL186));
sram_cell_6t_5 inst_cell_186_48 (.BL(BL48),.BLN(BLN48),.WL(WL186));
sram_cell_6t_5 inst_cell_186_49 (.BL(BL49),.BLN(BLN49),.WL(WL186));
sram_cell_6t_5 inst_cell_186_50 (.BL(BL50),.BLN(BLN50),.WL(WL186));
sram_cell_6t_5 inst_cell_186_51 (.BL(BL51),.BLN(BLN51),.WL(WL186));
sram_cell_6t_5 inst_cell_186_52 (.BL(BL52),.BLN(BLN52),.WL(WL186));
sram_cell_6t_5 inst_cell_186_53 (.BL(BL53),.BLN(BLN53),.WL(WL186));
sram_cell_6t_5 inst_cell_186_54 (.BL(BL54),.BLN(BLN54),.WL(WL186));
sram_cell_6t_5 inst_cell_186_55 (.BL(BL55),.BLN(BLN55),.WL(WL186));
sram_cell_6t_5 inst_cell_186_56 (.BL(BL56),.BLN(BLN56),.WL(WL186));
sram_cell_6t_5 inst_cell_186_57 (.BL(BL57),.BLN(BLN57),.WL(WL186));
sram_cell_6t_5 inst_cell_186_58 (.BL(BL58),.BLN(BLN58),.WL(WL186));
sram_cell_6t_5 inst_cell_186_59 (.BL(BL59),.BLN(BLN59),.WL(WL186));
sram_cell_6t_5 inst_cell_186_60 (.BL(BL60),.BLN(BLN60),.WL(WL186));
sram_cell_6t_5 inst_cell_186_61 (.BL(BL61),.BLN(BLN61),.WL(WL186));
sram_cell_6t_5 inst_cell_186_62 (.BL(BL62),.BLN(BLN62),.WL(WL186));
sram_cell_6t_5 inst_cell_186_63 (.BL(BL63),.BLN(BLN63),.WL(WL186));
sram_cell_6t_5 inst_cell_186_64 (.BL(BL64),.BLN(BLN64),.WL(WL186));
sram_cell_6t_5 inst_cell_186_65 (.BL(BL65),.BLN(BLN65),.WL(WL186));
sram_cell_6t_5 inst_cell_186_66 (.BL(BL66),.BLN(BLN66),.WL(WL186));
sram_cell_6t_5 inst_cell_186_67 (.BL(BL67),.BLN(BLN67),.WL(WL186));
sram_cell_6t_5 inst_cell_186_68 (.BL(BL68),.BLN(BLN68),.WL(WL186));
sram_cell_6t_5 inst_cell_186_69 (.BL(BL69),.BLN(BLN69),.WL(WL186));
sram_cell_6t_5 inst_cell_186_70 (.BL(BL70),.BLN(BLN70),.WL(WL186));
sram_cell_6t_5 inst_cell_186_71 (.BL(BL71),.BLN(BLN71),.WL(WL186));
sram_cell_6t_5 inst_cell_186_72 (.BL(BL72),.BLN(BLN72),.WL(WL186));
sram_cell_6t_5 inst_cell_186_73 (.BL(BL73),.BLN(BLN73),.WL(WL186));
sram_cell_6t_5 inst_cell_186_74 (.BL(BL74),.BLN(BLN74),.WL(WL186));
sram_cell_6t_5 inst_cell_186_75 (.BL(BL75),.BLN(BLN75),.WL(WL186));
sram_cell_6t_5 inst_cell_186_76 (.BL(BL76),.BLN(BLN76),.WL(WL186));
sram_cell_6t_5 inst_cell_186_77 (.BL(BL77),.BLN(BLN77),.WL(WL186));
sram_cell_6t_5 inst_cell_186_78 (.BL(BL78),.BLN(BLN78),.WL(WL186));
sram_cell_6t_5 inst_cell_186_79 (.BL(BL79),.BLN(BLN79),.WL(WL186));
sram_cell_6t_5 inst_cell_186_80 (.BL(BL80),.BLN(BLN80),.WL(WL186));
sram_cell_6t_5 inst_cell_186_81 (.BL(BL81),.BLN(BLN81),.WL(WL186));
sram_cell_6t_5 inst_cell_186_82 (.BL(BL82),.BLN(BLN82),.WL(WL186));
sram_cell_6t_5 inst_cell_186_83 (.BL(BL83),.BLN(BLN83),.WL(WL186));
sram_cell_6t_5 inst_cell_186_84 (.BL(BL84),.BLN(BLN84),.WL(WL186));
sram_cell_6t_5 inst_cell_186_85 (.BL(BL85),.BLN(BLN85),.WL(WL186));
sram_cell_6t_5 inst_cell_186_86 (.BL(BL86),.BLN(BLN86),.WL(WL186));
sram_cell_6t_5 inst_cell_186_87 (.BL(BL87),.BLN(BLN87),.WL(WL186));
sram_cell_6t_5 inst_cell_186_88 (.BL(BL88),.BLN(BLN88),.WL(WL186));
sram_cell_6t_5 inst_cell_186_89 (.BL(BL89),.BLN(BLN89),.WL(WL186));
sram_cell_6t_5 inst_cell_186_90 (.BL(BL90),.BLN(BLN90),.WL(WL186));
sram_cell_6t_5 inst_cell_186_91 (.BL(BL91),.BLN(BLN91),.WL(WL186));
sram_cell_6t_5 inst_cell_186_92 (.BL(BL92),.BLN(BLN92),.WL(WL186));
sram_cell_6t_5 inst_cell_186_93 (.BL(BL93),.BLN(BLN93),.WL(WL186));
sram_cell_6t_5 inst_cell_186_94 (.BL(BL94),.BLN(BLN94),.WL(WL186));
sram_cell_6t_5 inst_cell_186_95 (.BL(BL95),.BLN(BLN95),.WL(WL186));
sram_cell_6t_5 inst_cell_186_96 (.BL(BL96),.BLN(BLN96),.WL(WL186));
sram_cell_6t_5 inst_cell_186_97 (.BL(BL97),.BLN(BLN97),.WL(WL186));
sram_cell_6t_5 inst_cell_186_98 (.BL(BL98),.BLN(BLN98),.WL(WL186));
sram_cell_6t_5 inst_cell_186_99 (.BL(BL99),.BLN(BLN99),.WL(WL186));
sram_cell_6t_5 inst_cell_186_100 (.BL(BL100),.BLN(BLN100),.WL(WL186));
sram_cell_6t_5 inst_cell_186_101 (.BL(BL101),.BLN(BLN101),.WL(WL186));
sram_cell_6t_5 inst_cell_186_102 (.BL(BL102),.BLN(BLN102),.WL(WL186));
sram_cell_6t_5 inst_cell_186_103 (.BL(BL103),.BLN(BLN103),.WL(WL186));
sram_cell_6t_5 inst_cell_186_104 (.BL(BL104),.BLN(BLN104),.WL(WL186));
sram_cell_6t_5 inst_cell_186_105 (.BL(BL105),.BLN(BLN105),.WL(WL186));
sram_cell_6t_5 inst_cell_186_106 (.BL(BL106),.BLN(BLN106),.WL(WL186));
sram_cell_6t_5 inst_cell_186_107 (.BL(BL107),.BLN(BLN107),.WL(WL186));
sram_cell_6t_5 inst_cell_186_108 (.BL(BL108),.BLN(BLN108),.WL(WL186));
sram_cell_6t_5 inst_cell_186_109 (.BL(BL109),.BLN(BLN109),.WL(WL186));
sram_cell_6t_5 inst_cell_186_110 (.BL(BL110),.BLN(BLN110),.WL(WL186));
sram_cell_6t_5 inst_cell_186_111 (.BL(BL111),.BLN(BLN111),.WL(WL186));
sram_cell_6t_5 inst_cell_186_112 (.BL(BL112),.BLN(BLN112),.WL(WL186));
sram_cell_6t_5 inst_cell_186_113 (.BL(BL113),.BLN(BLN113),.WL(WL186));
sram_cell_6t_5 inst_cell_186_114 (.BL(BL114),.BLN(BLN114),.WL(WL186));
sram_cell_6t_5 inst_cell_186_115 (.BL(BL115),.BLN(BLN115),.WL(WL186));
sram_cell_6t_5 inst_cell_186_116 (.BL(BL116),.BLN(BLN116),.WL(WL186));
sram_cell_6t_5 inst_cell_186_117 (.BL(BL117),.BLN(BLN117),.WL(WL186));
sram_cell_6t_5 inst_cell_186_118 (.BL(BL118),.BLN(BLN118),.WL(WL186));
sram_cell_6t_5 inst_cell_186_119 (.BL(BL119),.BLN(BLN119),.WL(WL186));
sram_cell_6t_5 inst_cell_186_120 (.BL(BL120),.BLN(BLN120),.WL(WL186));
sram_cell_6t_5 inst_cell_186_121 (.BL(BL121),.BLN(BLN121),.WL(WL186));
sram_cell_6t_5 inst_cell_186_122 (.BL(BL122),.BLN(BLN122),.WL(WL186));
sram_cell_6t_5 inst_cell_186_123 (.BL(BL123),.BLN(BLN123),.WL(WL186));
sram_cell_6t_5 inst_cell_186_124 (.BL(BL124),.BLN(BLN124),.WL(WL186));
sram_cell_6t_5 inst_cell_186_125 (.BL(BL125),.BLN(BLN125),.WL(WL186));
sram_cell_6t_5 inst_cell_186_126 (.BL(BL126),.BLN(BLN126),.WL(WL186));
sram_cell_6t_5 inst_cell_186_127 (.BL(BL127),.BLN(BLN127),.WL(WL186));
sram_cell_6t_5 inst_cell_187_0 (.BL(BL0),.BLN(BLN0),.WL(WL187));
sram_cell_6t_5 inst_cell_187_1 (.BL(BL1),.BLN(BLN1),.WL(WL187));
sram_cell_6t_5 inst_cell_187_2 (.BL(BL2),.BLN(BLN2),.WL(WL187));
sram_cell_6t_5 inst_cell_187_3 (.BL(BL3),.BLN(BLN3),.WL(WL187));
sram_cell_6t_5 inst_cell_187_4 (.BL(BL4),.BLN(BLN4),.WL(WL187));
sram_cell_6t_5 inst_cell_187_5 (.BL(BL5),.BLN(BLN5),.WL(WL187));
sram_cell_6t_5 inst_cell_187_6 (.BL(BL6),.BLN(BLN6),.WL(WL187));
sram_cell_6t_5 inst_cell_187_7 (.BL(BL7),.BLN(BLN7),.WL(WL187));
sram_cell_6t_5 inst_cell_187_8 (.BL(BL8),.BLN(BLN8),.WL(WL187));
sram_cell_6t_5 inst_cell_187_9 (.BL(BL9),.BLN(BLN9),.WL(WL187));
sram_cell_6t_5 inst_cell_187_10 (.BL(BL10),.BLN(BLN10),.WL(WL187));
sram_cell_6t_5 inst_cell_187_11 (.BL(BL11),.BLN(BLN11),.WL(WL187));
sram_cell_6t_5 inst_cell_187_12 (.BL(BL12),.BLN(BLN12),.WL(WL187));
sram_cell_6t_5 inst_cell_187_13 (.BL(BL13),.BLN(BLN13),.WL(WL187));
sram_cell_6t_5 inst_cell_187_14 (.BL(BL14),.BLN(BLN14),.WL(WL187));
sram_cell_6t_5 inst_cell_187_15 (.BL(BL15),.BLN(BLN15),.WL(WL187));
sram_cell_6t_5 inst_cell_187_16 (.BL(BL16),.BLN(BLN16),.WL(WL187));
sram_cell_6t_5 inst_cell_187_17 (.BL(BL17),.BLN(BLN17),.WL(WL187));
sram_cell_6t_5 inst_cell_187_18 (.BL(BL18),.BLN(BLN18),.WL(WL187));
sram_cell_6t_5 inst_cell_187_19 (.BL(BL19),.BLN(BLN19),.WL(WL187));
sram_cell_6t_5 inst_cell_187_20 (.BL(BL20),.BLN(BLN20),.WL(WL187));
sram_cell_6t_5 inst_cell_187_21 (.BL(BL21),.BLN(BLN21),.WL(WL187));
sram_cell_6t_5 inst_cell_187_22 (.BL(BL22),.BLN(BLN22),.WL(WL187));
sram_cell_6t_5 inst_cell_187_23 (.BL(BL23),.BLN(BLN23),.WL(WL187));
sram_cell_6t_5 inst_cell_187_24 (.BL(BL24),.BLN(BLN24),.WL(WL187));
sram_cell_6t_5 inst_cell_187_25 (.BL(BL25),.BLN(BLN25),.WL(WL187));
sram_cell_6t_5 inst_cell_187_26 (.BL(BL26),.BLN(BLN26),.WL(WL187));
sram_cell_6t_5 inst_cell_187_27 (.BL(BL27),.BLN(BLN27),.WL(WL187));
sram_cell_6t_5 inst_cell_187_28 (.BL(BL28),.BLN(BLN28),.WL(WL187));
sram_cell_6t_5 inst_cell_187_29 (.BL(BL29),.BLN(BLN29),.WL(WL187));
sram_cell_6t_5 inst_cell_187_30 (.BL(BL30),.BLN(BLN30),.WL(WL187));
sram_cell_6t_5 inst_cell_187_31 (.BL(BL31),.BLN(BLN31),.WL(WL187));
sram_cell_6t_5 inst_cell_187_32 (.BL(BL32),.BLN(BLN32),.WL(WL187));
sram_cell_6t_5 inst_cell_187_33 (.BL(BL33),.BLN(BLN33),.WL(WL187));
sram_cell_6t_5 inst_cell_187_34 (.BL(BL34),.BLN(BLN34),.WL(WL187));
sram_cell_6t_5 inst_cell_187_35 (.BL(BL35),.BLN(BLN35),.WL(WL187));
sram_cell_6t_5 inst_cell_187_36 (.BL(BL36),.BLN(BLN36),.WL(WL187));
sram_cell_6t_5 inst_cell_187_37 (.BL(BL37),.BLN(BLN37),.WL(WL187));
sram_cell_6t_5 inst_cell_187_38 (.BL(BL38),.BLN(BLN38),.WL(WL187));
sram_cell_6t_5 inst_cell_187_39 (.BL(BL39),.BLN(BLN39),.WL(WL187));
sram_cell_6t_5 inst_cell_187_40 (.BL(BL40),.BLN(BLN40),.WL(WL187));
sram_cell_6t_5 inst_cell_187_41 (.BL(BL41),.BLN(BLN41),.WL(WL187));
sram_cell_6t_5 inst_cell_187_42 (.BL(BL42),.BLN(BLN42),.WL(WL187));
sram_cell_6t_5 inst_cell_187_43 (.BL(BL43),.BLN(BLN43),.WL(WL187));
sram_cell_6t_5 inst_cell_187_44 (.BL(BL44),.BLN(BLN44),.WL(WL187));
sram_cell_6t_5 inst_cell_187_45 (.BL(BL45),.BLN(BLN45),.WL(WL187));
sram_cell_6t_5 inst_cell_187_46 (.BL(BL46),.BLN(BLN46),.WL(WL187));
sram_cell_6t_5 inst_cell_187_47 (.BL(BL47),.BLN(BLN47),.WL(WL187));
sram_cell_6t_5 inst_cell_187_48 (.BL(BL48),.BLN(BLN48),.WL(WL187));
sram_cell_6t_5 inst_cell_187_49 (.BL(BL49),.BLN(BLN49),.WL(WL187));
sram_cell_6t_5 inst_cell_187_50 (.BL(BL50),.BLN(BLN50),.WL(WL187));
sram_cell_6t_5 inst_cell_187_51 (.BL(BL51),.BLN(BLN51),.WL(WL187));
sram_cell_6t_5 inst_cell_187_52 (.BL(BL52),.BLN(BLN52),.WL(WL187));
sram_cell_6t_5 inst_cell_187_53 (.BL(BL53),.BLN(BLN53),.WL(WL187));
sram_cell_6t_5 inst_cell_187_54 (.BL(BL54),.BLN(BLN54),.WL(WL187));
sram_cell_6t_5 inst_cell_187_55 (.BL(BL55),.BLN(BLN55),.WL(WL187));
sram_cell_6t_5 inst_cell_187_56 (.BL(BL56),.BLN(BLN56),.WL(WL187));
sram_cell_6t_5 inst_cell_187_57 (.BL(BL57),.BLN(BLN57),.WL(WL187));
sram_cell_6t_5 inst_cell_187_58 (.BL(BL58),.BLN(BLN58),.WL(WL187));
sram_cell_6t_5 inst_cell_187_59 (.BL(BL59),.BLN(BLN59),.WL(WL187));
sram_cell_6t_5 inst_cell_187_60 (.BL(BL60),.BLN(BLN60),.WL(WL187));
sram_cell_6t_5 inst_cell_187_61 (.BL(BL61),.BLN(BLN61),.WL(WL187));
sram_cell_6t_5 inst_cell_187_62 (.BL(BL62),.BLN(BLN62),.WL(WL187));
sram_cell_6t_5 inst_cell_187_63 (.BL(BL63),.BLN(BLN63),.WL(WL187));
sram_cell_6t_5 inst_cell_187_64 (.BL(BL64),.BLN(BLN64),.WL(WL187));
sram_cell_6t_5 inst_cell_187_65 (.BL(BL65),.BLN(BLN65),.WL(WL187));
sram_cell_6t_5 inst_cell_187_66 (.BL(BL66),.BLN(BLN66),.WL(WL187));
sram_cell_6t_5 inst_cell_187_67 (.BL(BL67),.BLN(BLN67),.WL(WL187));
sram_cell_6t_5 inst_cell_187_68 (.BL(BL68),.BLN(BLN68),.WL(WL187));
sram_cell_6t_5 inst_cell_187_69 (.BL(BL69),.BLN(BLN69),.WL(WL187));
sram_cell_6t_5 inst_cell_187_70 (.BL(BL70),.BLN(BLN70),.WL(WL187));
sram_cell_6t_5 inst_cell_187_71 (.BL(BL71),.BLN(BLN71),.WL(WL187));
sram_cell_6t_5 inst_cell_187_72 (.BL(BL72),.BLN(BLN72),.WL(WL187));
sram_cell_6t_5 inst_cell_187_73 (.BL(BL73),.BLN(BLN73),.WL(WL187));
sram_cell_6t_5 inst_cell_187_74 (.BL(BL74),.BLN(BLN74),.WL(WL187));
sram_cell_6t_5 inst_cell_187_75 (.BL(BL75),.BLN(BLN75),.WL(WL187));
sram_cell_6t_5 inst_cell_187_76 (.BL(BL76),.BLN(BLN76),.WL(WL187));
sram_cell_6t_5 inst_cell_187_77 (.BL(BL77),.BLN(BLN77),.WL(WL187));
sram_cell_6t_5 inst_cell_187_78 (.BL(BL78),.BLN(BLN78),.WL(WL187));
sram_cell_6t_5 inst_cell_187_79 (.BL(BL79),.BLN(BLN79),.WL(WL187));
sram_cell_6t_5 inst_cell_187_80 (.BL(BL80),.BLN(BLN80),.WL(WL187));
sram_cell_6t_5 inst_cell_187_81 (.BL(BL81),.BLN(BLN81),.WL(WL187));
sram_cell_6t_5 inst_cell_187_82 (.BL(BL82),.BLN(BLN82),.WL(WL187));
sram_cell_6t_5 inst_cell_187_83 (.BL(BL83),.BLN(BLN83),.WL(WL187));
sram_cell_6t_5 inst_cell_187_84 (.BL(BL84),.BLN(BLN84),.WL(WL187));
sram_cell_6t_5 inst_cell_187_85 (.BL(BL85),.BLN(BLN85),.WL(WL187));
sram_cell_6t_5 inst_cell_187_86 (.BL(BL86),.BLN(BLN86),.WL(WL187));
sram_cell_6t_5 inst_cell_187_87 (.BL(BL87),.BLN(BLN87),.WL(WL187));
sram_cell_6t_5 inst_cell_187_88 (.BL(BL88),.BLN(BLN88),.WL(WL187));
sram_cell_6t_5 inst_cell_187_89 (.BL(BL89),.BLN(BLN89),.WL(WL187));
sram_cell_6t_5 inst_cell_187_90 (.BL(BL90),.BLN(BLN90),.WL(WL187));
sram_cell_6t_5 inst_cell_187_91 (.BL(BL91),.BLN(BLN91),.WL(WL187));
sram_cell_6t_5 inst_cell_187_92 (.BL(BL92),.BLN(BLN92),.WL(WL187));
sram_cell_6t_5 inst_cell_187_93 (.BL(BL93),.BLN(BLN93),.WL(WL187));
sram_cell_6t_5 inst_cell_187_94 (.BL(BL94),.BLN(BLN94),.WL(WL187));
sram_cell_6t_5 inst_cell_187_95 (.BL(BL95),.BLN(BLN95),.WL(WL187));
sram_cell_6t_5 inst_cell_187_96 (.BL(BL96),.BLN(BLN96),.WL(WL187));
sram_cell_6t_5 inst_cell_187_97 (.BL(BL97),.BLN(BLN97),.WL(WL187));
sram_cell_6t_5 inst_cell_187_98 (.BL(BL98),.BLN(BLN98),.WL(WL187));
sram_cell_6t_5 inst_cell_187_99 (.BL(BL99),.BLN(BLN99),.WL(WL187));
sram_cell_6t_5 inst_cell_187_100 (.BL(BL100),.BLN(BLN100),.WL(WL187));
sram_cell_6t_5 inst_cell_187_101 (.BL(BL101),.BLN(BLN101),.WL(WL187));
sram_cell_6t_5 inst_cell_187_102 (.BL(BL102),.BLN(BLN102),.WL(WL187));
sram_cell_6t_5 inst_cell_187_103 (.BL(BL103),.BLN(BLN103),.WL(WL187));
sram_cell_6t_5 inst_cell_187_104 (.BL(BL104),.BLN(BLN104),.WL(WL187));
sram_cell_6t_5 inst_cell_187_105 (.BL(BL105),.BLN(BLN105),.WL(WL187));
sram_cell_6t_5 inst_cell_187_106 (.BL(BL106),.BLN(BLN106),.WL(WL187));
sram_cell_6t_5 inst_cell_187_107 (.BL(BL107),.BLN(BLN107),.WL(WL187));
sram_cell_6t_5 inst_cell_187_108 (.BL(BL108),.BLN(BLN108),.WL(WL187));
sram_cell_6t_5 inst_cell_187_109 (.BL(BL109),.BLN(BLN109),.WL(WL187));
sram_cell_6t_5 inst_cell_187_110 (.BL(BL110),.BLN(BLN110),.WL(WL187));
sram_cell_6t_5 inst_cell_187_111 (.BL(BL111),.BLN(BLN111),.WL(WL187));
sram_cell_6t_5 inst_cell_187_112 (.BL(BL112),.BLN(BLN112),.WL(WL187));
sram_cell_6t_5 inst_cell_187_113 (.BL(BL113),.BLN(BLN113),.WL(WL187));
sram_cell_6t_5 inst_cell_187_114 (.BL(BL114),.BLN(BLN114),.WL(WL187));
sram_cell_6t_5 inst_cell_187_115 (.BL(BL115),.BLN(BLN115),.WL(WL187));
sram_cell_6t_5 inst_cell_187_116 (.BL(BL116),.BLN(BLN116),.WL(WL187));
sram_cell_6t_5 inst_cell_187_117 (.BL(BL117),.BLN(BLN117),.WL(WL187));
sram_cell_6t_5 inst_cell_187_118 (.BL(BL118),.BLN(BLN118),.WL(WL187));
sram_cell_6t_5 inst_cell_187_119 (.BL(BL119),.BLN(BLN119),.WL(WL187));
sram_cell_6t_5 inst_cell_187_120 (.BL(BL120),.BLN(BLN120),.WL(WL187));
sram_cell_6t_5 inst_cell_187_121 (.BL(BL121),.BLN(BLN121),.WL(WL187));
sram_cell_6t_5 inst_cell_187_122 (.BL(BL122),.BLN(BLN122),.WL(WL187));
sram_cell_6t_5 inst_cell_187_123 (.BL(BL123),.BLN(BLN123),.WL(WL187));
sram_cell_6t_5 inst_cell_187_124 (.BL(BL124),.BLN(BLN124),.WL(WL187));
sram_cell_6t_5 inst_cell_187_125 (.BL(BL125),.BLN(BLN125),.WL(WL187));
sram_cell_6t_5 inst_cell_187_126 (.BL(BL126),.BLN(BLN126),.WL(WL187));
sram_cell_6t_5 inst_cell_187_127 (.BL(BL127),.BLN(BLN127),.WL(WL187));
sram_cell_6t_5 inst_cell_188_0 (.BL(BL0),.BLN(BLN0),.WL(WL188));
sram_cell_6t_5 inst_cell_188_1 (.BL(BL1),.BLN(BLN1),.WL(WL188));
sram_cell_6t_5 inst_cell_188_2 (.BL(BL2),.BLN(BLN2),.WL(WL188));
sram_cell_6t_5 inst_cell_188_3 (.BL(BL3),.BLN(BLN3),.WL(WL188));
sram_cell_6t_5 inst_cell_188_4 (.BL(BL4),.BLN(BLN4),.WL(WL188));
sram_cell_6t_5 inst_cell_188_5 (.BL(BL5),.BLN(BLN5),.WL(WL188));
sram_cell_6t_5 inst_cell_188_6 (.BL(BL6),.BLN(BLN6),.WL(WL188));
sram_cell_6t_5 inst_cell_188_7 (.BL(BL7),.BLN(BLN7),.WL(WL188));
sram_cell_6t_5 inst_cell_188_8 (.BL(BL8),.BLN(BLN8),.WL(WL188));
sram_cell_6t_5 inst_cell_188_9 (.BL(BL9),.BLN(BLN9),.WL(WL188));
sram_cell_6t_5 inst_cell_188_10 (.BL(BL10),.BLN(BLN10),.WL(WL188));
sram_cell_6t_5 inst_cell_188_11 (.BL(BL11),.BLN(BLN11),.WL(WL188));
sram_cell_6t_5 inst_cell_188_12 (.BL(BL12),.BLN(BLN12),.WL(WL188));
sram_cell_6t_5 inst_cell_188_13 (.BL(BL13),.BLN(BLN13),.WL(WL188));
sram_cell_6t_5 inst_cell_188_14 (.BL(BL14),.BLN(BLN14),.WL(WL188));
sram_cell_6t_5 inst_cell_188_15 (.BL(BL15),.BLN(BLN15),.WL(WL188));
sram_cell_6t_5 inst_cell_188_16 (.BL(BL16),.BLN(BLN16),.WL(WL188));
sram_cell_6t_5 inst_cell_188_17 (.BL(BL17),.BLN(BLN17),.WL(WL188));
sram_cell_6t_5 inst_cell_188_18 (.BL(BL18),.BLN(BLN18),.WL(WL188));
sram_cell_6t_5 inst_cell_188_19 (.BL(BL19),.BLN(BLN19),.WL(WL188));
sram_cell_6t_5 inst_cell_188_20 (.BL(BL20),.BLN(BLN20),.WL(WL188));
sram_cell_6t_5 inst_cell_188_21 (.BL(BL21),.BLN(BLN21),.WL(WL188));
sram_cell_6t_5 inst_cell_188_22 (.BL(BL22),.BLN(BLN22),.WL(WL188));
sram_cell_6t_5 inst_cell_188_23 (.BL(BL23),.BLN(BLN23),.WL(WL188));
sram_cell_6t_5 inst_cell_188_24 (.BL(BL24),.BLN(BLN24),.WL(WL188));
sram_cell_6t_5 inst_cell_188_25 (.BL(BL25),.BLN(BLN25),.WL(WL188));
sram_cell_6t_5 inst_cell_188_26 (.BL(BL26),.BLN(BLN26),.WL(WL188));
sram_cell_6t_5 inst_cell_188_27 (.BL(BL27),.BLN(BLN27),.WL(WL188));
sram_cell_6t_5 inst_cell_188_28 (.BL(BL28),.BLN(BLN28),.WL(WL188));
sram_cell_6t_5 inst_cell_188_29 (.BL(BL29),.BLN(BLN29),.WL(WL188));
sram_cell_6t_5 inst_cell_188_30 (.BL(BL30),.BLN(BLN30),.WL(WL188));
sram_cell_6t_5 inst_cell_188_31 (.BL(BL31),.BLN(BLN31),.WL(WL188));
sram_cell_6t_5 inst_cell_188_32 (.BL(BL32),.BLN(BLN32),.WL(WL188));
sram_cell_6t_5 inst_cell_188_33 (.BL(BL33),.BLN(BLN33),.WL(WL188));
sram_cell_6t_5 inst_cell_188_34 (.BL(BL34),.BLN(BLN34),.WL(WL188));
sram_cell_6t_5 inst_cell_188_35 (.BL(BL35),.BLN(BLN35),.WL(WL188));
sram_cell_6t_5 inst_cell_188_36 (.BL(BL36),.BLN(BLN36),.WL(WL188));
sram_cell_6t_5 inst_cell_188_37 (.BL(BL37),.BLN(BLN37),.WL(WL188));
sram_cell_6t_5 inst_cell_188_38 (.BL(BL38),.BLN(BLN38),.WL(WL188));
sram_cell_6t_5 inst_cell_188_39 (.BL(BL39),.BLN(BLN39),.WL(WL188));
sram_cell_6t_5 inst_cell_188_40 (.BL(BL40),.BLN(BLN40),.WL(WL188));
sram_cell_6t_5 inst_cell_188_41 (.BL(BL41),.BLN(BLN41),.WL(WL188));
sram_cell_6t_5 inst_cell_188_42 (.BL(BL42),.BLN(BLN42),.WL(WL188));
sram_cell_6t_5 inst_cell_188_43 (.BL(BL43),.BLN(BLN43),.WL(WL188));
sram_cell_6t_5 inst_cell_188_44 (.BL(BL44),.BLN(BLN44),.WL(WL188));
sram_cell_6t_5 inst_cell_188_45 (.BL(BL45),.BLN(BLN45),.WL(WL188));
sram_cell_6t_5 inst_cell_188_46 (.BL(BL46),.BLN(BLN46),.WL(WL188));
sram_cell_6t_5 inst_cell_188_47 (.BL(BL47),.BLN(BLN47),.WL(WL188));
sram_cell_6t_5 inst_cell_188_48 (.BL(BL48),.BLN(BLN48),.WL(WL188));
sram_cell_6t_5 inst_cell_188_49 (.BL(BL49),.BLN(BLN49),.WL(WL188));
sram_cell_6t_5 inst_cell_188_50 (.BL(BL50),.BLN(BLN50),.WL(WL188));
sram_cell_6t_5 inst_cell_188_51 (.BL(BL51),.BLN(BLN51),.WL(WL188));
sram_cell_6t_5 inst_cell_188_52 (.BL(BL52),.BLN(BLN52),.WL(WL188));
sram_cell_6t_5 inst_cell_188_53 (.BL(BL53),.BLN(BLN53),.WL(WL188));
sram_cell_6t_5 inst_cell_188_54 (.BL(BL54),.BLN(BLN54),.WL(WL188));
sram_cell_6t_5 inst_cell_188_55 (.BL(BL55),.BLN(BLN55),.WL(WL188));
sram_cell_6t_5 inst_cell_188_56 (.BL(BL56),.BLN(BLN56),.WL(WL188));
sram_cell_6t_5 inst_cell_188_57 (.BL(BL57),.BLN(BLN57),.WL(WL188));
sram_cell_6t_5 inst_cell_188_58 (.BL(BL58),.BLN(BLN58),.WL(WL188));
sram_cell_6t_5 inst_cell_188_59 (.BL(BL59),.BLN(BLN59),.WL(WL188));
sram_cell_6t_5 inst_cell_188_60 (.BL(BL60),.BLN(BLN60),.WL(WL188));
sram_cell_6t_5 inst_cell_188_61 (.BL(BL61),.BLN(BLN61),.WL(WL188));
sram_cell_6t_5 inst_cell_188_62 (.BL(BL62),.BLN(BLN62),.WL(WL188));
sram_cell_6t_5 inst_cell_188_63 (.BL(BL63),.BLN(BLN63),.WL(WL188));
sram_cell_6t_5 inst_cell_188_64 (.BL(BL64),.BLN(BLN64),.WL(WL188));
sram_cell_6t_5 inst_cell_188_65 (.BL(BL65),.BLN(BLN65),.WL(WL188));
sram_cell_6t_5 inst_cell_188_66 (.BL(BL66),.BLN(BLN66),.WL(WL188));
sram_cell_6t_5 inst_cell_188_67 (.BL(BL67),.BLN(BLN67),.WL(WL188));
sram_cell_6t_5 inst_cell_188_68 (.BL(BL68),.BLN(BLN68),.WL(WL188));
sram_cell_6t_5 inst_cell_188_69 (.BL(BL69),.BLN(BLN69),.WL(WL188));
sram_cell_6t_5 inst_cell_188_70 (.BL(BL70),.BLN(BLN70),.WL(WL188));
sram_cell_6t_5 inst_cell_188_71 (.BL(BL71),.BLN(BLN71),.WL(WL188));
sram_cell_6t_5 inst_cell_188_72 (.BL(BL72),.BLN(BLN72),.WL(WL188));
sram_cell_6t_5 inst_cell_188_73 (.BL(BL73),.BLN(BLN73),.WL(WL188));
sram_cell_6t_5 inst_cell_188_74 (.BL(BL74),.BLN(BLN74),.WL(WL188));
sram_cell_6t_5 inst_cell_188_75 (.BL(BL75),.BLN(BLN75),.WL(WL188));
sram_cell_6t_5 inst_cell_188_76 (.BL(BL76),.BLN(BLN76),.WL(WL188));
sram_cell_6t_5 inst_cell_188_77 (.BL(BL77),.BLN(BLN77),.WL(WL188));
sram_cell_6t_5 inst_cell_188_78 (.BL(BL78),.BLN(BLN78),.WL(WL188));
sram_cell_6t_5 inst_cell_188_79 (.BL(BL79),.BLN(BLN79),.WL(WL188));
sram_cell_6t_5 inst_cell_188_80 (.BL(BL80),.BLN(BLN80),.WL(WL188));
sram_cell_6t_5 inst_cell_188_81 (.BL(BL81),.BLN(BLN81),.WL(WL188));
sram_cell_6t_5 inst_cell_188_82 (.BL(BL82),.BLN(BLN82),.WL(WL188));
sram_cell_6t_5 inst_cell_188_83 (.BL(BL83),.BLN(BLN83),.WL(WL188));
sram_cell_6t_5 inst_cell_188_84 (.BL(BL84),.BLN(BLN84),.WL(WL188));
sram_cell_6t_5 inst_cell_188_85 (.BL(BL85),.BLN(BLN85),.WL(WL188));
sram_cell_6t_5 inst_cell_188_86 (.BL(BL86),.BLN(BLN86),.WL(WL188));
sram_cell_6t_5 inst_cell_188_87 (.BL(BL87),.BLN(BLN87),.WL(WL188));
sram_cell_6t_5 inst_cell_188_88 (.BL(BL88),.BLN(BLN88),.WL(WL188));
sram_cell_6t_5 inst_cell_188_89 (.BL(BL89),.BLN(BLN89),.WL(WL188));
sram_cell_6t_5 inst_cell_188_90 (.BL(BL90),.BLN(BLN90),.WL(WL188));
sram_cell_6t_5 inst_cell_188_91 (.BL(BL91),.BLN(BLN91),.WL(WL188));
sram_cell_6t_5 inst_cell_188_92 (.BL(BL92),.BLN(BLN92),.WL(WL188));
sram_cell_6t_5 inst_cell_188_93 (.BL(BL93),.BLN(BLN93),.WL(WL188));
sram_cell_6t_5 inst_cell_188_94 (.BL(BL94),.BLN(BLN94),.WL(WL188));
sram_cell_6t_5 inst_cell_188_95 (.BL(BL95),.BLN(BLN95),.WL(WL188));
sram_cell_6t_5 inst_cell_188_96 (.BL(BL96),.BLN(BLN96),.WL(WL188));
sram_cell_6t_5 inst_cell_188_97 (.BL(BL97),.BLN(BLN97),.WL(WL188));
sram_cell_6t_5 inst_cell_188_98 (.BL(BL98),.BLN(BLN98),.WL(WL188));
sram_cell_6t_5 inst_cell_188_99 (.BL(BL99),.BLN(BLN99),.WL(WL188));
sram_cell_6t_5 inst_cell_188_100 (.BL(BL100),.BLN(BLN100),.WL(WL188));
sram_cell_6t_5 inst_cell_188_101 (.BL(BL101),.BLN(BLN101),.WL(WL188));
sram_cell_6t_5 inst_cell_188_102 (.BL(BL102),.BLN(BLN102),.WL(WL188));
sram_cell_6t_5 inst_cell_188_103 (.BL(BL103),.BLN(BLN103),.WL(WL188));
sram_cell_6t_5 inst_cell_188_104 (.BL(BL104),.BLN(BLN104),.WL(WL188));
sram_cell_6t_5 inst_cell_188_105 (.BL(BL105),.BLN(BLN105),.WL(WL188));
sram_cell_6t_5 inst_cell_188_106 (.BL(BL106),.BLN(BLN106),.WL(WL188));
sram_cell_6t_5 inst_cell_188_107 (.BL(BL107),.BLN(BLN107),.WL(WL188));
sram_cell_6t_5 inst_cell_188_108 (.BL(BL108),.BLN(BLN108),.WL(WL188));
sram_cell_6t_5 inst_cell_188_109 (.BL(BL109),.BLN(BLN109),.WL(WL188));
sram_cell_6t_5 inst_cell_188_110 (.BL(BL110),.BLN(BLN110),.WL(WL188));
sram_cell_6t_5 inst_cell_188_111 (.BL(BL111),.BLN(BLN111),.WL(WL188));
sram_cell_6t_5 inst_cell_188_112 (.BL(BL112),.BLN(BLN112),.WL(WL188));
sram_cell_6t_5 inst_cell_188_113 (.BL(BL113),.BLN(BLN113),.WL(WL188));
sram_cell_6t_5 inst_cell_188_114 (.BL(BL114),.BLN(BLN114),.WL(WL188));
sram_cell_6t_5 inst_cell_188_115 (.BL(BL115),.BLN(BLN115),.WL(WL188));
sram_cell_6t_5 inst_cell_188_116 (.BL(BL116),.BLN(BLN116),.WL(WL188));
sram_cell_6t_5 inst_cell_188_117 (.BL(BL117),.BLN(BLN117),.WL(WL188));
sram_cell_6t_5 inst_cell_188_118 (.BL(BL118),.BLN(BLN118),.WL(WL188));
sram_cell_6t_5 inst_cell_188_119 (.BL(BL119),.BLN(BLN119),.WL(WL188));
sram_cell_6t_5 inst_cell_188_120 (.BL(BL120),.BLN(BLN120),.WL(WL188));
sram_cell_6t_5 inst_cell_188_121 (.BL(BL121),.BLN(BLN121),.WL(WL188));
sram_cell_6t_5 inst_cell_188_122 (.BL(BL122),.BLN(BLN122),.WL(WL188));
sram_cell_6t_5 inst_cell_188_123 (.BL(BL123),.BLN(BLN123),.WL(WL188));
sram_cell_6t_5 inst_cell_188_124 (.BL(BL124),.BLN(BLN124),.WL(WL188));
sram_cell_6t_5 inst_cell_188_125 (.BL(BL125),.BLN(BLN125),.WL(WL188));
sram_cell_6t_5 inst_cell_188_126 (.BL(BL126),.BLN(BLN126),.WL(WL188));
sram_cell_6t_5 inst_cell_188_127 (.BL(BL127),.BLN(BLN127),.WL(WL188));
sram_cell_6t_5 inst_cell_189_0 (.BL(BL0),.BLN(BLN0),.WL(WL189));
sram_cell_6t_5 inst_cell_189_1 (.BL(BL1),.BLN(BLN1),.WL(WL189));
sram_cell_6t_5 inst_cell_189_2 (.BL(BL2),.BLN(BLN2),.WL(WL189));
sram_cell_6t_5 inst_cell_189_3 (.BL(BL3),.BLN(BLN3),.WL(WL189));
sram_cell_6t_5 inst_cell_189_4 (.BL(BL4),.BLN(BLN4),.WL(WL189));
sram_cell_6t_5 inst_cell_189_5 (.BL(BL5),.BLN(BLN5),.WL(WL189));
sram_cell_6t_5 inst_cell_189_6 (.BL(BL6),.BLN(BLN6),.WL(WL189));
sram_cell_6t_5 inst_cell_189_7 (.BL(BL7),.BLN(BLN7),.WL(WL189));
sram_cell_6t_5 inst_cell_189_8 (.BL(BL8),.BLN(BLN8),.WL(WL189));
sram_cell_6t_5 inst_cell_189_9 (.BL(BL9),.BLN(BLN9),.WL(WL189));
sram_cell_6t_5 inst_cell_189_10 (.BL(BL10),.BLN(BLN10),.WL(WL189));
sram_cell_6t_5 inst_cell_189_11 (.BL(BL11),.BLN(BLN11),.WL(WL189));
sram_cell_6t_5 inst_cell_189_12 (.BL(BL12),.BLN(BLN12),.WL(WL189));
sram_cell_6t_5 inst_cell_189_13 (.BL(BL13),.BLN(BLN13),.WL(WL189));
sram_cell_6t_5 inst_cell_189_14 (.BL(BL14),.BLN(BLN14),.WL(WL189));
sram_cell_6t_5 inst_cell_189_15 (.BL(BL15),.BLN(BLN15),.WL(WL189));
sram_cell_6t_5 inst_cell_189_16 (.BL(BL16),.BLN(BLN16),.WL(WL189));
sram_cell_6t_5 inst_cell_189_17 (.BL(BL17),.BLN(BLN17),.WL(WL189));
sram_cell_6t_5 inst_cell_189_18 (.BL(BL18),.BLN(BLN18),.WL(WL189));
sram_cell_6t_5 inst_cell_189_19 (.BL(BL19),.BLN(BLN19),.WL(WL189));
sram_cell_6t_5 inst_cell_189_20 (.BL(BL20),.BLN(BLN20),.WL(WL189));
sram_cell_6t_5 inst_cell_189_21 (.BL(BL21),.BLN(BLN21),.WL(WL189));
sram_cell_6t_5 inst_cell_189_22 (.BL(BL22),.BLN(BLN22),.WL(WL189));
sram_cell_6t_5 inst_cell_189_23 (.BL(BL23),.BLN(BLN23),.WL(WL189));
sram_cell_6t_5 inst_cell_189_24 (.BL(BL24),.BLN(BLN24),.WL(WL189));
sram_cell_6t_5 inst_cell_189_25 (.BL(BL25),.BLN(BLN25),.WL(WL189));
sram_cell_6t_5 inst_cell_189_26 (.BL(BL26),.BLN(BLN26),.WL(WL189));
sram_cell_6t_5 inst_cell_189_27 (.BL(BL27),.BLN(BLN27),.WL(WL189));
sram_cell_6t_5 inst_cell_189_28 (.BL(BL28),.BLN(BLN28),.WL(WL189));
sram_cell_6t_5 inst_cell_189_29 (.BL(BL29),.BLN(BLN29),.WL(WL189));
sram_cell_6t_5 inst_cell_189_30 (.BL(BL30),.BLN(BLN30),.WL(WL189));
sram_cell_6t_5 inst_cell_189_31 (.BL(BL31),.BLN(BLN31),.WL(WL189));
sram_cell_6t_5 inst_cell_189_32 (.BL(BL32),.BLN(BLN32),.WL(WL189));
sram_cell_6t_5 inst_cell_189_33 (.BL(BL33),.BLN(BLN33),.WL(WL189));
sram_cell_6t_5 inst_cell_189_34 (.BL(BL34),.BLN(BLN34),.WL(WL189));
sram_cell_6t_5 inst_cell_189_35 (.BL(BL35),.BLN(BLN35),.WL(WL189));
sram_cell_6t_5 inst_cell_189_36 (.BL(BL36),.BLN(BLN36),.WL(WL189));
sram_cell_6t_5 inst_cell_189_37 (.BL(BL37),.BLN(BLN37),.WL(WL189));
sram_cell_6t_5 inst_cell_189_38 (.BL(BL38),.BLN(BLN38),.WL(WL189));
sram_cell_6t_5 inst_cell_189_39 (.BL(BL39),.BLN(BLN39),.WL(WL189));
sram_cell_6t_5 inst_cell_189_40 (.BL(BL40),.BLN(BLN40),.WL(WL189));
sram_cell_6t_5 inst_cell_189_41 (.BL(BL41),.BLN(BLN41),.WL(WL189));
sram_cell_6t_5 inst_cell_189_42 (.BL(BL42),.BLN(BLN42),.WL(WL189));
sram_cell_6t_5 inst_cell_189_43 (.BL(BL43),.BLN(BLN43),.WL(WL189));
sram_cell_6t_5 inst_cell_189_44 (.BL(BL44),.BLN(BLN44),.WL(WL189));
sram_cell_6t_5 inst_cell_189_45 (.BL(BL45),.BLN(BLN45),.WL(WL189));
sram_cell_6t_5 inst_cell_189_46 (.BL(BL46),.BLN(BLN46),.WL(WL189));
sram_cell_6t_5 inst_cell_189_47 (.BL(BL47),.BLN(BLN47),.WL(WL189));
sram_cell_6t_5 inst_cell_189_48 (.BL(BL48),.BLN(BLN48),.WL(WL189));
sram_cell_6t_5 inst_cell_189_49 (.BL(BL49),.BLN(BLN49),.WL(WL189));
sram_cell_6t_5 inst_cell_189_50 (.BL(BL50),.BLN(BLN50),.WL(WL189));
sram_cell_6t_5 inst_cell_189_51 (.BL(BL51),.BLN(BLN51),.WL(WL189));
sram_cell_6t_5 inst_cell_189_52 (.BL(BL52),.BLN(BLN52),.WL(WL189));
sram_cell_6t_5 inst_cell_189_53 (.BL(BL53),.BLN(BLN53),.WL(WL189));
sram_cell_6t_5 inst_cell_189_54 (.BL(BL54),.BLN(BLN54),.WL(WL189));
sram_cell_6t_5 inst_cell_189_55 (.BL(BL55),.BLN(BLN55),.WL(WL189));
sram_cell_6t_5 inst_cell_189_56 (.BL(BL56),.BLN(BLN56),.WL(WL189));
sram_cell_6t_5 inst_cell_189_57 (.BL(BL57),.BLN(BLN57),.WL(WL189));
sram_cell_6t_5 inst_cell_189_58 (.BL(BL58),.BLN(BLN58),.WL(WL189));
sram_cell_6t_5 inst_cell_189_59 (.BL(BL59),.BLN(BLN59),.WL(WL189));
sram_cell_6t_5 inst_cell_189_60 (.BL(BL60),.BLN(BLN60),.WL(WL189));
sram_cell_6t_5 inst_cell_189_61 (.BL(BL61),.BLN(BLN61),.WL(WL189));
sram_cell_6t_5 inst_cell_189_62 (.BL(BL62),.BLN(BLN62),.WL(WL189));
sram_cell_6t_5 inst_cell_189_63 (.BL(BL63),.BLN(BLN63),.WL(WL189));
sram_cell_6t_5 inst_cell_189_64 (.BL(BL64),.BLN(BLN64),.WL(WL189));
sram_cell_6t_5 inst_cell_189_65 (.BL(BL65),.BLN(BLN65),.WL(WL189));
sram_cell_6t_5 inst_cell_189_66 (.BL(BL66),.BLN(BLN66),.WL(WL189));
sram_cell_6t_5 inst_cell_189_67 (.BL(BL67),.BLN(BLN67),.WL(WL189));
sram_cell_6t_5 inst_cell_189_68 (.BL(BL68),.BLN(BLN68),.WL(WL189));
sram_cell_6t_5 inst_cell_189_69 (.BL(BL69),.BLN(BLN69),.WL(WL189));
sram_cell_6t_5 inst_cell_189_70 (.BL(BL70),.BLN(BLN70),.WL(WL189));
sram_cell_6t_5 inst_cell_189_71 (.BL(BL71),.BLN(BLN71),.WL(WL189));
sram_cell_6t_5 inst_cell_189_72 (.BL(BL72),.BLN(BLN72),.WL(WL189));
sram_cell_6t_5 inst_cell_189_73 (.BL(BL73),.BLN(BLN73),.WL(WL189));
sram_cell_6t_5 inst_cell_189_74 (.BL(BL74),.BLN(BLN74),.WL(WL189));
sram_cell_6t_5 inst_cell_189_75 (.BL(BL75),.BLN(BLN75),.WL(WL189));
sram_cell_6t_5 inst_cell_189_76 (.BL(BL76),.BLN(BLN76),.WL(WL189));
sram_cell_6t_5 inst_cell_189_77 (.BL(BL77),.BLN(BLN77),.WL(WL189));
sram_cell_6t_5 inst_cell_189_78 (.BL(BL78),.BLN(BLN78),.WL(WL189));
sram_cell_6t_5 inst_cell_189_79 (.BL(BL79),.BLN(BLN79),.WL(WL189));
sram_cell_6t_5 inst_cell_189_80 (.BL(BL80),.BLN(BLN80),.WL(WL189));
sram_cell_6t_5 inst_cell_189_81 (.BL(BL81),.BLN(BLN81),.WL(WL189));
sram_cell_6t_5 inst_cell_189_82 (.BL(BL82),.BLN(BLN82),.WL(WL189));
sram_cell_6t_5 inst_cell_189_83 (.BL(BL83),.BLN(BLN83),.WL(WL189));
sram_cell_6t_5 inst_cell_189_84 (.BL(BL84),.BLN(BLN84),.WL(WL189));
sram_cell_6t_5 inst_cell_189_85 (.BL(BL85),.BLN(BLN85),.WL(WL189));
sram_cell_6t_5 inst_cell_189_86 (.BL(BL86),.BLN(BLN86),.WL(WL189));
sram_cell_6t_5 inst_cell_189_87 (.BL(BL87),.BLN(BLN87),.WL(WL189));
sram_cell_6t_5 inst_cell_189_88 (.BL(BL88),.BLN(BLN88),.WL(WL189));
sram_cell_6t_5 inst_cell_189_89 (.BL(BL89),.BLN(BLN89),.WL(WL189));
sram_cell_6t_5 inst_cell_189_90 (.BL(BL90),.BLN(BLN90),.WL(WL189));
sram_cell_6t_5 inst_cell_189_91 (.BL(BL91),.BLN(BLN91),.WL(WL189));
sram_cell_6t_5 inst_cell_189_92 (.BL(BL92),.BLN(BLN92),.WL(WL189));
sram_cell_6t_5 inst_cell_189_93 (.BL(BL93),.BLN(BLN93),.WL(WL189));
sram_cell_6t_5 inst_cell_189_94 (.BL(BL94),.BLN(BLN94),.WL(WL189));
sram_cell_6t_5 inst_cell_189_95 (.BL(BL95),.BLN(BLN95),.WL(WL189));
sram_cell_6t_5 inst_cell_189_96 (.BL(BL96),.BLN(BLN96),.WL(WL189));
sram_cell_6t_5 inst_cell_189_97 (.BL(BL97),.BLN(BLN97),.WL(WL189));
sram_cell_6t_5 inst_cell_189_98 (.BL(BL98),.BLN(BLN98),.WL(WL189));
sram_cell_6t_5 inst_cell_189_99 (.BL(BL99),.BLN(BLN99),.WL(WL189));
sram_cell_6t_5 inst_cell_189_100 (.BL(BL100),.BLN(BLN100),.WL(WL189));
sram_cell_6t_5 inst_cell_189_101 (.BL(BL101),.BLN(BLN101),.WL(WL189));
sram_cell_6t_5 inst_cell_189_102 (.BL(BL102),.BLN(BLN102),.WL(WL189));
sram_cell_6t_5 inst_cell_189_103 (.BL(BL103),.BLN(BLN103),.WL(WL189));
sram_cell_6t_5 inst_cell_189_104 (.BL(BL104),.BLN(BLN104),.WL(WL189));
sram_cell_6t_5 inst_cell_189_105 (.BL(BL105),.BLN(BLN105),.WL(WL189));
sram_cell_6t_5 inst_cell_189_106 (.BL(BL106),.BLN(BLN106),.WL(WL189));
sram_cell_6t_5 inst_cell_189_107 (.BL(BL107),.BLN(BLN107),.WL(WL189));
sram_cell_6t_5 inst_cell_189_108 (.BL(BL108),.BLN(BLN108),.WL(WL189));
sram_cell_6t_5 inst_cell_189_109 (.BL(BL109),.BLN(BLN109),.WL(WL189));
sram_cell_6t_5 inst_cell_189_110 (.BL(BL110),.BLN(BLN110),.WL(WL189));
sram_cell_6t_5 inst_cell_189_111 (.BL(BL111),.BLN(BLN111),.WL(WL189));
sram_cell_6t_5 inst_cell_189_112 (.BL(BL112),.BLN(BLN112),.WL(WL189));
sram_cell_6t_5 inst_cell_189_113 (.BL(BL113),.BLN(BLN113),.WL(WL189));
sram_cell_6t_5 inst_cell_189_114 (.BL(BL114),.BLN(BLN114),.WL(WL189));
sram_cell_6t_5 inst_cell_189_115 (.BL(BL115),.BLN(BLN115),.WL(WL189));
sram_cell_6t_5 inst_cell_189_116 (.BL(BL116),.BLN(BLN116),.WL(WL189));
sram_cell_6t_5 inst_cell_189_117 (.BL(BL117),.BLN(BLN117),.WL(WL189));
sram_cell_6t_5 inst_cell_189_118 (.BL(BL118),.BLN(BLN118),.WL(WL189));
sram_cell_6t_5 inst_cell_189_119 (.BL(BL119),.BLN(BLN119),.WL(WL189));
sram_cell_6t_5 inst_cell_189_120 (.BL(BL120),.BLN(BLN120),.WL(WL189));
sram_cell_6t_5 inst_cell_189_121 (.BL(BL121),.BLN(BLN121),.WL(WL189));
sram_cell_6t_5 inst_cell_189_122 (.BL(BL122),.BLN(BLN122),.WL(WL189));
sram_cell_6t_5 inst_cell_189_123 (.BL(BL123),.BLN(BLN123),.WL(WL189));
sram_cell_6t_5 inst_cell_189_124 (.BL(BL124),.BLN(BLN124),.WL(WL189));
sram_cell_6t_5 inst_cell_189_125 (.BL(BL125),.BLN(BLN125),.WL(WL189));
sram_cell_6t_5 inst_cell_189_126 (.BL(BL126),.BLN(BLN126),.WL(WL189));
sram_cell_6t_5 inst_cell_189_127 (.BL(BL127),.BLN(BLN127),.WL(WL189));
sram_cell_6t_5 inst_cell_190_0 (.BL(BL0),.BLN(BLN0),.WL(WL190));
sram_cell_6t_5 inst_cell_190_1 (.BL(BL1),.BLN(BLN1),.WL(WL190));
sram_cell_6t_5 inst_cell_190_2 (.BL(BL2),.BLN(BLN2),.WL(WL190));
sram_cell_6t_5 inst_cell_190_3 (.BL(BL3),.BLN(BLN3),.WL(WL190));
sram_cell_6t_5 inst_cell_190_4 (.BL(BL4),.BLN(BLN4),.WL(WL190));
sram_cell_6t_5 inst_cell_190_5 (.BL(BL5),.BLN(BLN5),.WL(WL190));
sram_cell_6t_5 inst_cell_190_6 (.BL(BL6),.BLN(BLN6),.WL(WL190));
sram_cell_6t_5 inst_cell_190_7 (.BL(BL7),.BLN(BLN7),.WL(WL190));
sram_cell_6t_5 inst_cell_190_8 (.BL(BL8),.BLN(BLN8),.WL(WL190));
sram_cell_6t_5 inst_cell_190_9 (.BL(BL9),.BLN(BLN9),.WL(WL190));
sram_cell_6t_5 inst_cell_190_10 (.BL(BL10),.BLN(BLN10),.WL(WL190));
sram_cell_6t_5 inst_cell_190_11 (.BL(BL11),.BLN(BLN11),.WL(WL190));
sram_cell_6t_5 inst_cell_190_12 (.BL(BL12),.BLN(BLN12),.WL(WL190));
sram_cell_6t_5 inst_cell_190_13 (.BL(BL13),.BLN(BLN13),.WL(WL190));
sram_cell_6t_5 inst_cell_190_14 (.BL(BL14),.BLN(BLN14),.WL(WL190));
sram_cell_6t_5 inst_cell_190_15 (.BL(BL15),.BLN(BLN15),.WL(WL190));
sram_cell_6t_5 inst_cell_190_16 (.BL(BL16),.BLN(BLN16),.WL(WL190));
sram_cell_6t_5 inst_cell_190_17 (.BL(BL17),.BLN(BLN17),.WL(WL190));
sram_cell_6t_5 inst_cell_190_18 (.BL(BL18),.BLN(BLN18),.WL(WL190));
sram_cell_6t_5 inst_cell_190_19 (.BL(BL19),.BLN(BLN19),.WL(WL190));
sram_cell_6t_5 inst_cell_190_20 (.BL(BL20),.BLN(BLN20),.WL(WL190));
sram_cell_6t_5 inst_cell_190_21 (.BL(BL21),.BLN(BLN21),.WL(WL190));
sram_cell_6t_5 inst_cell_190_22 (.BL(BL22),.BLN(BLN22),.WL(WL190));
sram_cell_6t_5 inst_cell_190_23 (.BL(BL23),.BLN(BLN23),.WL(WL190));
sram_cell_6t_5 inst_cell_190_24 (.BL(BL24),.BLN(BLN24),.WL(WL190));
sram_cell_6t_5 inst_cell_190_25 (.BL(BL25),.BLN(BLN25),.WL(WL190));
sram_cell_6t_5 inst_cell_190_26 (.BL(BL26),.BLN(BLN26),.WL(WL190));
sram_cell_6t_5 inst_cell_190_27 (.BL(BL27),.BLN(BLN27),.WL(WL190));
sram_cell_6t_5 inst_cell_190_28 (.BL(BL28),.BLN(BLN28),.WL(WL190));
sram_cell_6t_5 inst_cell_190_29 (.BL(BL29),.BLN(BLN29),.WL(WL190));
sram_cell_6t_5 inst_cell_190_30 (.BL(BL30),.BLN(BLN30),.WL(WL190));
sram_cell_6t_5 inst_cell_190_31 (.BL(BL31),.BLN(BLN31),.WL(WL190));
sram_cell_6t_5 inst_cell_190_32 (.BL(BL32),.BLN(BLN32),.WL(WL190));
sram_cell_6t_5 inst_cell_190_33 (.BL(BL33),.BLN(BLN33),.WL(WL190));
sram_cell_6t_5 inst_cell_190_34 (.BL(BL34),.BLN(BLN34),.WL(WL190));
sram_cell_6t_5 inst_cell_190_35 (.BL(BL35),.BLN(BLN35),.WL(WL190));
sram_cell_6t_5 inst_cell_190_36 (.BL(BL36),.BLN(BLN36),.WL(WL190));
sram_cell_6t_5 inst_cell_190_37 (.BL(BL37),.BLN(BLN37),.WL(WL190));
sram_cell_6t_5 inst_cell_190_38 (.BL(BL38),.BLN(BLN38),.WL(WL190));
sram_cell_6t_5 inst_cell_190_39 (.BL(BL39),.BLN(BLN39),.WL(WL190));
sram_cell_6t_5 inst_cell_190_40 (.BL(BL40),.BLN(BLN40),.WL(WL190));
sram_cell_6t_5 inst_cell_190_41 (.BL(BL41),.BLN(BLN41),.WL(WL190));
sram_cell_6t_5 inst_cell_190_42 (.BL(BL42),.BLN(BLN42),.WL(WL190));
sram_cell_6t_5 inst_cell_190_43 (.BL(BL43),.BLN(BLN43),.WL(WL190));
sram_cell_6t_5 inst_cell_190_44 (.BL(BL44),.BLN(BLN44),.WL(WL190));
sram_cell_6t_5 inst_cell_190_45 (.BL(BL45),.BLN(BLN45),.WL(WL190));
sram_cell_6t_5 inst_cell_190_46 (.BL(BL46),.BLN(BLN46),.WL(WL190));
sram_cell_6t_5 inst_cell_190_47 (.BL(BL47),.BLN(BLN47),.WL(WL190));
sram_cell_6t_5 inst_cell_190_48 (.BL(BL48),.BLN(BLN48),.WL(WL190));
sram_cell_6t_5 inst_cell_190_49 (.BL(BL49),.BLN(BLN49),.WL(WL190));
sram_cell_6t_5 inst_cell_190_50 (.BL(BL50),.BLN(BLN50),.WL(WL190));
sram_cell_6t_5 inst_cell_190_51 (.BL(BL51),.BLN(BLN51),.WL(WL190));
sram_cell_6t_5 inst_cell_190_52 (.BL(BL52),.BLN(BLN52),.WL(WL190));
sram_cell_6t_5 inst_cell_190_53 (.BL(BL53),.BLN(BLN53),.WL(WL190));
sram_cell_6t_5 inst_cell_190_54 (.BL(BL54),.BLN(BLN54),.WL(WL190));
sram_cell_6t_5 inst_cell_190_55 (.BL(BL55),.BLN(BLN55),.WL(WL190));
sram_cell_6t_5 inst_cell_190_56 (.BL(BL56),.BLN(BLN56),.WL(WL190));
sram_cell_6t_5 inst_cell_190_57 (.BL(BL57),.BLN(BLN57),.WL(WL190));
sram_cell_6t_5 inst_cell_190_58 (.BL(BL58),.BLN(BLN58),.WL(WL190));
sram_cell_6t_5 inst_cell_190_59 (.BL(BL59),.BLN(BLN59),.WL(WL190));
sram_cell_6t_5 inst_cell_190_60 (.BL(BL60),.BLN(BLN60),.WL(WL190));
sram_cell_6t_5 inst_cell_190_61 (.BL(BL61),.BLN(BLN61),.WL(WL190));
sram_cell_6t_5 inst_cell_190_62 (.BL(BL62),.BLN(BLN62),.WL(WL190));
sram_cell_6t_5 inst_cell_190_63 (.BL(BL63),.BLN(BLN63),.WL(WL190));
sram_cell_6t_5 inst_cell_190_64 (.BL(BL64),.BLN(BLN64),.WL(WL190));
sram_cell_6t_5 inst_cell_190_65 (.BL(BL65),.BLN(BLN65),.WL(WL190));
sram_cell_6t_5 inst_cell_190_66 (.BL(BL66),.BLN(BLN66),.WL(WL190));
sram_cell_6t_5 inst_cell_190_67 (.BL(BL67),.BLN(BLN67),.WL(WL190));
sram_cell_6t_5 inst_cell_190_68 (.BL(BL68),.BLN(BLN68),.WL(WL190));
sram_cell_6t_5 inst_cell_190_69 (.BL(BL69),.BLN(BLN69),.WL(WL190));
sram_cell_6t_5 inst_cell_190_70 (.BL(BL70),.BLN(BLN70),.WL(WL190));
sram_cell_6t_5 inst_cell_190_71 (.BL(BL71),.BLN(BLN71),.WL(WL190));
sram_cell_6t_5 inst_cell_190_72 (.BL(BL72),.BLN(BLN72),.WL(WL190));
sram_cell_6t_5 inst_cell_190_73 (.BL(BL73),.BLN(BLN73),.WL(WL190));
sram_cell_6t_5 inst_cell_190_74 (.BL(BL74),.BLN(BLN74),.WL(WL190));
sram_cell_6t_5 inst_cell_190_75 (.BL(BL75),.BLN(BLN75),.WL(WL190));
sram_cell_6t_5 inst_cell_190_76 (.BL(BL76),.BLN(BLN76),.WL(WL190));
sram_cell_6t_5 inst_cell_190_77 (.BL(BL77),.BLN(BLN77),.WL(WL190));
sram_cell_6t_5 inst_cell_190_78 (.BL(BL78),.BLN(BLN78),.WL(WL190));
sram_cell_6t_5 inst_cell_190_79 (.BL(BL79),.BLN(BLN79),.WL(WL190));
sram_cell_6t_5 inst_cell_190_80 (.BL(BL80),.BLN(BLN80),.WL(WL190));
sram_cell_6t_5 inst_cell_190_81 (.BL(BL81),.BLN(BLN81),.WL(WL190));
sram_cell_6t_5 inst_cell_190_82 (.BL(BL82),.BLN(BLN82),.WL(WL190));
sram_cell_6t_5 inst_cell_190_83 (.BL(BL83),.BLN(BLN83),.WL(WL190));
sram_cell_6t_5 inst_cell_190_84 (.BL(BL84),.BLN(BLN84),.WL(WL190));
sram_cell_6t_5 inst_cell_190_85 (.BL(BL85),.BLN(BLN85),.WL(WL190));
sram_cell_6t_5 inst_cell_190_86 (.BL(BL86),.BLN(BLN86),.WL(WL190));
sram_cell_6t_5 inst_cell_190_87 (.BL(BL87),.BLN(BLN87),.WL(WL190));
sram_cell_6t_5 inst_cell_190_88 (.BL(BL88),.BLN(BLN88),.WL(WL190));
sram_cell_6t_5 inst_cell_190_89 (.BL(BL89),.BLN(BLN89),.WL(WL190));
sram_cell_6t_5 inst_cell_190_90 (.BL(BL90),.BLN(BLN90),.WL(WL190));
sram_cell_6t_5 inst_cell_190_91 (.BL(BL91),.BLN(BLN91),.WL(WL190));
sram_cell_6t_5 inst_cell_190_92 (.BL(BL92),.BLN(BLN92),.WL(WL190));
sram_cell_6t_5 inst_cell_190_93 (.BL(BL93),.BLN(BLN93),.WL(WL190));
sram_cell_6t_5 inst_cell_190_94 (.BL(BL94),.BLN(BLN94),.WL(WL190));
sram_cell_6t_5 inst_cell_190_95 (.BL(BL95),.BLN(BLN95),.WL(WL190));
sram_cell_6t_5 inst_cell_190_96 (.BL(BL96),.BLN(BLN96),.WL(WL190));
sram_cell_6t_5 inst_cell_190_97 (.BL(BL97),.BLN(BLN97),.WL(WL190));
sram_cell_6t_5 inst_cell_190_98 (.BL(BL98),.BLN(BLN98),.WL(WL190));
sram_cell_6t_5 inst_cell_190_99 (.BL(BL99),.BLN(BLN99),.WL(WL190));
sram_cell_6t_5 inst_cell_190_100 (.BL(BL100),.BLN(BLN100),.WL(WL190));
sram_cell_6t_5 inst_cell_190_101 (.BL(BL101),.BLN(BLN101),.WL(WL190));
sram_cell_6t_5 inst_cell_190_102 (.BL(BL102),.BLN(BLN102),.WL(WL190));
sram_cell_6t_5 inst_cell_190_103 (.BL(BL103),.BLN(BLN103),.WL(WL190));
sram_cell_6t_5 inst_cell_190_104 (.BL(BL104),.BLN(BLN104),.WL(WL190));
sram_cell_6t_5 inst_cell_190_105 (.BL(BL105),.BLN(BLN105),.WL(WL190));
sram_cell_6t_5 inst_cell_190_106 (.BL(BL106),.BLN(BLN106),.WL(WL190));
sram_cell_6t_5 inst_cell_190_107 (.BL(BL107),.BLN(BLN107),.WL(WL190));
sram_cell_6t_5 inst_cell_190_108 (.BL(BL108),.BLN(BLN108),.WL(WL190));
sram_cell_6t_5 inst_cell_190_109 (.BL(BL109),.BLN(BLN109),.WL(WL190));
sram_cell_6t_5 inst_cell_190_110 (.BL(BL110),.BLN(BLN110),.WL(WL190));
sram_cell_6t_5 inst_cell_190_111 (.BL(BL111),.BLN(BLN111),.WL(WL190));
sram_cell_6t_5 inst_cell_190_112 (.BL(BL112),.BLN(BLN112),.WL(WL190));
sram_cell_6t_5 inst_cell_190_113 (.BL(BL113),.BLN(BLN113),.WL(WL190));
sram_cell_6t_5 inst_cell_190_114 (.BL(BL114),.BLN(BLN114),.WL(WL190));
sram_cell_6t_5 inst_cell_190_115 (.BL(BL115),.BLN(BLN115),.WL(WL190));
sram_cell_6t_5 inst_cell_190_116 (.BL(BL116),.BLN(BLN116),.WL(WL190));
sram_cell_6t_5 inst_cell_190_117 (.BL(BL117),.BLN(BLN117),.WL(WL190));
sram_cell_6t_5 inst_cell_190_118 (.BL(BL118),.BLN(BLN118),.WL(WL190));
sram_cell_6t_5 inst_cell_190_119 (.BL(BL119),.BLN(BLN119),.WL(WL190));
sram_cell_6t_5 inst_cell_190_120 (.BL(BL120),.BLN(BLN120),.WL(WL190));
sram_cell_6t_5 inst_cell_190_121 (.BL(BL121),.BLN(BLN121),.WL(WL190));
sram_cell_6t_5 inst_cell_190_122 (.BL(BL122),.BLN(BLN122),.WL(WL190));
sram_cell_6t_5 inst_cell_190_123 (.BL(BL123),.BLN(BLN123),.WL(WL190));
sram_cell_6t_5 inst_cell_190_124 (.BL(BL124),.BLN(BLN124),.WL(WL190));
sram_cell_6t_5 inst_cell_190_125 (.BL(BL125),.BLN(BLN125),.WL(WL190));
sram_cell_6t_5 inst_cell_190_126 (.BL(BL126),.BLN(BLN126),.WL(WL190));
sram_cell_6t_5 inst_cell_190_127 (.BL(BL127),.BLN(BLN127),.WL(WL190));
sram_cell_6t_5 inst_cell_191_0 (.BL(BL0),.BLN(BLN0),.WL(WL191));
sram_cell_6t_5 inst_cell_191_1 (.BL(BL1),.BLN(BLN1),.WL(WL191));
sram_cell_6t_5 inst_cell_191_2 (.BL(BL2),.BLN(BLN2),.WL(WL191));
sram_cell_6t_5 inst_cell_191_3 (.BL(BL3),.BLN(BLN3),.WL(WL191));
sram_cell_6t_5 inst_cell_191_4 (.BL(BL4),.BLN(BLN4),.WL(WL191));
sram_cell_6t_5 inst_cell_191_5 (.BL(BL5),.BLN(BLN5),.WL(WL191));
sram_cell_6t_5 inst_cell_191_6 (.BL(BL6),.BLN(BLN6),.WL(WL191));
sram_cell_6t_5 inst_cell_191_7 (.BL(BL7),.BLN(BLN7),.WL(WL191));
sram_cell_6t_5 inst_cell_191_8 (.BL(BL8),.BLN(BLN8),.WL(WL191));
sram_cell_6t_5 inst_cell_191_9 (.BL(BL9),.BLN(BLN9),.WL(WL191));
sram_cell_6t_5 inst_cell_191_10 (.BL(BL10),.BLN(BLN10),.WL(WL191));
sram_cell_6t_5 inst_cell_191_11 (.BL(BL11),.BLN(BLN11),.WL(WL191));
sram_cell_6t_5 inst_cell_191_12 (.BL(BL12),.BLN(BLN12),.WL(WL191));
sram_cell_6t_5 inst_cell_191_13 (.BL(BL13),.BLN(BLN13),.WL(WL191));
sram_cell_6t_5 inst_cell_191_14 (.BL(BL14),.BLN(BLN14),.WL(WL191));
sram_cell_6t_5 inst_cell_191_15 (.BL(BL15),.BLN(BLN15),.WL(WL191));
sram_cell_6t_5 inst_cell_191_16 (.BL(BL16),.BLN(BLN16),.WL(WL191));
sram_cell_6t_5 inst_cell_191_17 (.BL(BL17),.BLN(BLN17),.WL(WL191));
sram_cell_6t_5 inst_cell_191_18 (.BL(BL18),.BLN(BLN18),.WL(WL191));
sram_cell_6t_5 inst_cell_191_19 (.BL(BL19),.BLN(BLN19),.WL(WL191));
sram_cell_6t_5 inst_cell_191_20 (.BL(BL20),.BLN(BLN20),.WL(WL191));
sram_cell_6t_5 inst_cell_191_21 (.BL(BL21),.BLN(BLN21),.WL(WL191));
sram_cell_6t_5 inst_cell_191_22 (.BL(BL22),.BLN(BLN22),.WL(WL191));
sram_cell_6t_5 inst_cell_191_23 (.BL(BL23),.BLN(BLN23),.WL(WL191));
sram_cell_6t_5 inst_cell_191_24 (.BL(BL24),.BLN(BLN24),.WL(WL191));
sram_cell_6t_5 inst_cell_191_25 (.BL(BL25),.BLN(BLN25),.WL(WL191));
sram_cell_6t_5 inst_cell_191_26 (.BL(BL26),.BLN(BLN26),.WL(WL191));
sram_cell_6t_5 inst_cell_191_27 (.BL(BL27),.BLN(BLN27),.WL(WL191));
sram_cell_6t_5 inst_cell_191_28 (.BL(BL28),.BLN(BLN28),.WL(WL191));
sram_cell_6t_5 inst_cell_191_29 (.BL(BL29),.BLN(BLN29),.WL(WL191));
sram_cell_6t_5 inst_cell_191_30 (.BL(BL30),.BLN(BLN30),.WL(WL191));
sram_cell_6t_5 inst_cell_191_31 (.BL(BL31),.BLN(BLN31),.WL(WL191));
sram_cell_6t_5 inst_cell_191_32 (.BL(BL32),.BLN(BLN32),.WL(WL191));
sram_cell_6t_5 inst_cell_191_33 (.BL(BL33),.BLN(BLN33),.WL(WL191));
sram_cell_6t_5 inst_cell_191_34 (.BL(BL34),.BLN(BLN34),.WL(WL191));
sram_cell_6t_5 inst_cell_191_35 (.BL(BL35),.BLN(BLN35),.WL(WL191));
sram_cell_6t_5 inst_cell_191_36 (.BL(BL36),.BLN(BLN36),.WL(WL191));
sram_cell_6t_5 inst_cell_191_37 (.BL(BL37),.BLN(BLN37),.WL(WL191));
sram_cell_6t_5 inst_cell_191_38 (.BL(BL38),.BLN(BLN38),.WL(WL191));
sram_cell_6t_5 inst_cell_191_39 (.BL(BL39),.BLN(BLN39),.WL(WL191));
sram_cell_6t_5 inst_cell_191_40 (.BL(BL40),.BLN(BLN40),.WL(WL191));
sram_cell_6t_5 inst_cell_191_41 (.BL(BL41),.BLN(BLN41),.WL(WL191));
sram_cell_6t_5 inst_cell_191_42 (.BL(BL42),.BLN(BLN42),.WL(WL191));
sram_cell_6t_5 inst_cell_191_43 (.BL(BL43),.BLN(BLN43),.WL(WL191));
sram_cell_6t_5 inst_cell_191_44 (.BL(BL44),.BLN(BLN44),.WL(WL191));
sram_cell_6t_5 inst_cell_191_45 (.BL(BL45),.BLN(BLN45),.WL(WL191));
sram_cell_6t_5 inst_cell_191_46 (.BL(BL46),.BLN(BLN46),.WL(WL191));
sram_cell_6t_5 inst_cell_191_47 (.BL(BL47),.BLN(BLN47),.WL(WL191));
sram_cell_6t_5 inst_cell_191_48 (.BL(BL48),.BLN(BLN48),.WL(WL191));
sram_cell_6t_5 inst_cell_191_49 (.BL(BL49),.BLN(BLN49),.WL(WL191));
sram_cell_6t_5 inst_cell_191_50 (.BL(BL50),.BLN(BLN50),.WL(WL191));
sram_cell_6t_5 inst_cell_191_51 (.BL(BL51),.BLN(BLN51),.WL(WL191));
sram_cell_6t_5 inst_cell_191_52 (.BL(BL52),.BLN(BLN52),.WL(WL191));
sram_cell_6t_5 inst_cell_191_53 (.BL(BL53),.BLN(BLN53),.WL(WL191));
sram_cell_6t_5 inst_cell_191_54 (.BL(BL54),.BLN(BLN54),.WL(WL191));
sram_cell_6t_5 inst_cell_191_55 (.BL(BL55),.BLN(BLN55),.WL(WL191));
sram_cell_6t_5 inst_cell_191_56 (.BL(BL56),.BLN(BLN56),.WL(WL191));
sram_cell_6t_5 inst_cell_191_57 (.BL(BL57),.BLN(BLN57),.WL(WL191));
sram_cell_6t_5 inst_cell_191_58 (.BL(BL58),.BLN(BLN58),.WL(WL191));
sram_cell_6t_5 inst_cell_191_59 (.BL(BL59),.BLN(BLN59),.WL(WL191));
sram_cell_6t_5 inst_cell_191_60 (.BL(BL60),.BLN(BLN60),.WL(WL191));
sram_cell_6t_5 inst_cell_191_61 (.BL(BL61),.BLN(BLN61),.WL(WL191));
sram_cell_6t_5 inst_cell_191_62 (.BL(BL62),.BLN(BLN62),.WL(WL191));
sram_cell_6t_5 inst_cell_191_63 (.BL(BL63),.BLN(BLN63),.WL(WL191));
sram_cell_6t_5 inst_cell_191_64 (.BL(BL64),.BLN(BLN64),.WL(WL191));
sram_cell_6t_5 inst_cell_191_65 (.BL(BL65),.BLN(BLN65),.WL(WL191));
sram_cell_6t_5 inst_cell_191_66 (.BL(BL66),.BLN(BLN66),.WL(WL191));
sram_cell_6t_5 inst_cell_191_67 (.BL(BL67),.BLN(BLN67),.WL(WL191));
sram_cell_6t_5 inst_cell_191_68 (.BL(BL68),.BLN(BLN68),.WL(WL191));
sram_cell_6t_5 inst_cell_191_69 (.BL(BL69),.BLN(BLN69),.WL(WL191));
sram_cell_6t_5 inst_cell_191_70 (.BL(BL70),.BLN(BLN70),.WL(WL191));
sram_cell_6t_5 inst_cell_191_71 (.BL(BL71),.BLN(BLN71),.WL(WL191));
sram_cell_6t_5 inst_cell_191_72 (.BL(BL72),.BLN(BLN72),.WL(WL191));
sram_cell_6t_5 inst_cell_191_73 (.BL(BL73),.BLN(BLN73),.WL(WL191));
sram_cell_6t_5 inst_cell_191_74 (.BL(BL74),.BLN(BLN74),.WL(WL191));
sram_cell_6t_5 inst_cell_191_75 (.BL(BL75),.BLN(BLN75),.WL(WL191));
sram_cell_6t_5 inst_cell_191_76 (.BL(BL76),.BLN(BLN76),.WL(WL191));
sram_cell_6t_5 inst_cell_191_77 (.BL(BL77),.BLN(BLN77),.WL(WL191));
sram_cell_6t_5 inst_cell_191_78 (.BL(BL78),.BLN(BLN78),.WL(WL191));
sram_cell_6t_5 inst_cell_191_79 (.BL(BL79),.BLN(BLN79),.WL(WL191));
sram_cell_6t_5 inst_cell_191_80 (.BL(BL80),.BLN(BLN80),.WL(WL191));
sram_cell_6t_5 inst_cell_191_81 (.BL(BL81),.BLN(BLN81),.WL(WL191));
sram_cell_6t_5 inst_cell_191_82 (.BL(BL82),.BLN(BLN82),.WL(WL191));
sram_cell_6t_5 inst_cell_191_83 (.BL(BL83),.BLN(BLN83),.WL(WL191));
sram_cell_6t_5 inst_cell_191_84 (.BL(BL84),.BLN(BLN84),.WL(WL191));
sram_cell_6t_5 inst_cell_191_85 (.BL(BL85),.BLN(BLN85),.WL(WL191));
sram_cell_6t_5 inst_cell_191_86 (.BL(BL86),.BLN(BLN86),.WL(WL191));
sram_cell_6t_5 inst_cell_191_87 (.BL(BL87),.BLN(BLN87),.WL(WL191));
sram_cell_6t_5 inst_cell_191_88 (.BL(BL88),.BLN(BLN88),.WL(WL191));
sram_cell_6t_5 inst_cell_191_89 (.BL(BL89),.BLN(BLN89),.WL(WL191));
sram_cell_6t_5 inst_cell_191_90 (.BL(BL90),.BLN(BLN90),.WL(WL191));
sram_cell_6t_5 inst_cell_191_91 (.BL(BL91),.BLN(BLN91),.WL(WL191));
sram_cell_6t_5 inst_cell_191_92 (.BL(BL92),.BLN(BLN92),.WL(WL191));
sram_cell_6t_5 inst_cell_191_93 (.BL(BL93),.BLN(BLN93),.WL(WL191));
sram_cell_6t_5 inst_cell_191_94 (.BL(BL94),.BLN(BLN94),.WL(WL191));
sram_cell_6t_5 inst_cell_191_95 (.BL(BL95),.BLN(BLN95),.WL(WL191));
sram_cell_6t_5 inst_cell_191_96 (.BL(BL96),.BLN(BLN96),.WL(WL191));
sram_cell_6t_5 inst_cell_191_97 (.BL(BL97),.BLN(BLN97),.WL(WL191));
sram_cell_6t_5 inst_cell_191_98 (.BL(BL98),.BLN(BLN98),.WL(WL191));
sram_cell_6t_5 inst_cell_191_99 (.BL(BL99),.BLN(BLN99),.WL(WL191));
sram_cell_6t_5 inst_cell_191_100 (.BL(BL100),.BLN(BLN100),.WL(WL191));
sram_cell_6t_5 inst_cell_191_101 (.BL(BL101),.BLN(BLN101),.WL(WL191));
sram_cell_6t_5 inst_cell_191_102 (.BL(BL102),.BLN(BLN102),.WL(WL191));
sram_cell_6t_5 inst_cell_191_103 (.BL(BL103),.BLN(BLN103),.WL(WL191));
sram_cell_6t_5 inst_cell_191_104 (.BL(BL104),.BLN(BLN104),.WL(WL191));
sram_cell_6t_5 inst_cell_191_105 (.BL(BL105),.BLN(BLN105),.WL(WL191));
sram_cell_6t_5 inst_cell_191_106 (.BL(BL106),.BLN(BLN106),.WL(WL191));
sram_cell_6t_5 inst_cell_191_107 (.BL(BL107),.BLN(BLN107),.WL(WL191));
sram_cell_6t_5 inst_cell_191_108 (.BL(BL108),.BLN(BLN108),.WL(WL191));
sram_cell_6t_5 inst_cell_191_109 (.BL(BL109),.BLN(BLN109),.WL(WL191));
sram_cell_6t_5 inst_cell_191_110 (.BL(BL110),.BLN(BLN110),.WL(WL191));
sram_cell_6t_5 inst_cell_191_111 (.BL(BL111),.BLN(BLN111),.WL(WL191));
sram_cell_6t_5 inst_cell_191_112 (.BL(BL112),.BLN(BLN112),.WL(WL191));
sram_cell_6t_5 inst_cell_191_113 (.BL(BL113),.BLN(BLN113),.WL(WL191));
sram_cell_6t_5 inst_cell_191_114 (.BL(BL114),.BLN(BLN114),.WL(WL191));
sram_cell_6t_5 inst_cell_191_115 (.BL(BL115),.BLN(BLN115),.WL(WL191));
sram_cell_6t_5 inst_cell_191_116 (.BL(BL116),.BLN(BLN116),.WL(WL191));
sram_cell_6t_5 inst_cell_191_117 (.BL(BL117),.BLN(BLN117),.WL(WL191));
sram_cell_6t_5 inst_cell_191_118 (.BL(BL118),.BLN(BLN118),.WL(WL191));
sram_cell_6t_5 inst_cell_191_119 (.BL(BL119),.BLN(BLN119),.WL(WL191));
sram_cell_6t_5 inst_cell_191_120 (.BL(BL120),.BLN(BLN120),.WL(WL191));
sram_cell_6t_5 inst_cell_191_121 (.BL(BL121),.BLN(BLN121),.WL(WL191));
sram_cell_6t_5 inst_cell_191_122 (.BL(BL122),.BLN(BLN122),.WL(WL191));
sram_cell_6t_5 inst_cell_191_123 (.BL(BL123),.BLN(BLN123),.WL(WL191));
sram_cell_6t_5 inst_cell_191_124 (.BL(BL124),.BLN(BLN124),.WL(WL191));
sram_cell_6t_5 inst_cell_191_125 (.BL(BL125),.BLN(BLN125),.WL(WL191));
sram_cell_6t_5 inst_cell_191_126 (.BL(BL126),.BLN(BLN126),.WL(WL191));
sram_cell_6t_5 inst_cell_191_127 (.BL(BL127),.BLN(BLN127),.WL(WL191));
sram_cell_6t_5 inst_cell_192_0 (.BL(BL0),.BLN(BLN0),.WL(WL192));
sram_cell_6t_5 inst_cell_192_1 (.BL(BL1),.BLN(BLN1),.WL(WL192));
sram_cell_6t_5 inst_cell_192_2 (.BL(BL2),.BLN(BLN2),.WL(WL192));
sram_cell_6t_5 inst_cell_192_3 (.BL(BL3),.BLN(BLN3),.WL(WL192));
sram_cell_6t_5 inst_cell_192_4 (.BL(BL4),.BLN(BLN4),.WL(WL192));
sram_cell_6t_5 inst_cell_192_5 (.BL(BL5),.BLN(BLN5),.WL(WL192));
sram_cell_6t_5 inst_cell_192_6 (.BL(BL6),.BLN(BLN6),.WL(WL192));
sram_cell_6t_5 inst_cell_192_7 (.BL(BL7),.BLN(BLN7),.WL(WL192));
sram_cell_6t_5 inst_cell_192_8 (.BL(BL8),.BLN(BLN8),.WL(WL192));
sram_cell_6t_5 inst_cell_192_9 (.BL(BL9),.BLN(BLN9),.WL(WL192));
sram_cell_6t_5 inst_cell_192_10 (.BL(BL10),.BLN(BLN10),.WL(WL192));
sram_cell_6t_5 inst_cell_192_11 (.BL(BL11),.BLN(BLN11),.WL(WL192));
sram_cell_6t_5 inst_cell_192_12 (.BL(BL12),.BLN(BLN12),.WL(WL192));
sram_cell_6t_5 inst_cell_192_13 (.BL(BL13),.BLN(BLN13),.WL(WL192));
sram_cell_6t_5 inst_cell_192_14 (.BL(BL14),.BLN(BLN14),.WL(WL192));
sram_cell_6t_5 inst_cell_192_15 (.BL(BL15),.BLN(BLN15),.WL(WL192));
sram_cell_6t_5 inst_cell_192_16 (.BL(BL16),.BLN(BLN16),.WL(WL192));
sram_cell_6t_5 inst_cell_192_17 (.BL(BL17),.BLN(BLN17),.WL(WL192));
sram_cell_6t_5 inst_cell_192_18 (.BL(BL18),.BLN(BLN18),.WL(WL192));
sram_cell_6t_5 inst_cell_192_19 (.BL(BL19),.BLN(BLN19),.WL(WL192));
sram_cell_6t_5 inst_cell_192_20 (.BL(BL20),.BLN(BLN20),.WL(WL192));
sram_cell_6t_5 inst_cell_192_21 (.BL(BL21),.BLN(BLN21),.WL(WL192));
sram_cell_6t_5 inst_cell_192_22 (.BL(BL22),.BLN(BLN22),.WL(WL192));
sram_cell_6t_5 inst_cell_192_23 (.BL(BL23),.BLN(BLN23),.WL(WL192));
sram_cell_6t_5 inst_cell_192_24 (.BL(BL24),.BLN(BLN24),.WL(WL192));
sram_cell_6t_5 inst_cell_192_25 (.BL(BL25),.BLN(BLN25),.WL(WL192));
sram_cell_6t_5 inst_cell_192_26 (.BL(BL26),.BLN(BLN26),.WL(WL192));
sram_cell_6t_5 inst_cell_192_27 (.BL(BL27),.BLN(BLN27),.WL(WL192));
sram_cell_6t_5 inst_cell_192_28 (.BL(BL28),.BLN(BLN28),.WL(WL192));
sram_cell_6t_5 inst_cell_192_29 (.BL(BL29),.BLN(BLN29),.WL(WL192));
sram_cell_6t_5 inst_cell_192_30 (.BL(BL30),.BLN(BLN30),.WL(WL192));
sram_cell_6t_5 inst_cell_192_31 (.BL(BL31),.BLN(BLN31),.WL(WL192));
sram_cell_6t_5 inst_cell_192_32 (.BL(BL32),.BLN(BLN32),.WL(WL192));
sram_cell_6t_5 inst_cell_192_33 (.BL(BL33),.BLN(BLN33),.WL(WL192));
sram_cell_6t_5 inst_cell_192_34 (.BL(BL34),.BLN(BLN34),.WL(WL192));
sram_cell_6t_5 inst_cell_192_35 (.BL(BL35),.BLN(BLN35),.WL(WL192));
sram_cell_6t_5 inst_cell_192_36 (.BL(BL36),.BLN(BLN36),.WL(WL192));
sram_cell_6t_5 inst_cell_192_37 (.BL(BL37),.BLN(BLN37),.WL(WL192));
sram_cell_6t_5 inst_cell_192_38 (.BL(BL38),.BLN(BLN38),.WL(WL192));
sram_cell_6t_5 inst_cell_192_39 (.BL(BL39),.BLN(BLN39),.WL(WL192));
sram_cell_6t_5 inst_cell_192_40 (.BL(BL40),.BLN(BLN40),.WL(WL192));
sram_cell_6t_5 inst_cell_192_41 (.BL(BL41),.BLN(BLN41),.WL(WL192));
sram_cell_6t_5 inst_cell_192_42 (.BL(BL42),.BLN(BLN42),.WL(WL192));
sram_cell_6t_5 inst_cell_192_43 (.BL(BL43),.BLN(BLN43),.WL(WL192));
sram_cell_6t_5 inst_cell_192_44 (.BL(BL44),.BLN(BLN44),.WL(WL192));
sram_cell_6t_5 inst_cell_192_45 (.BL(BL45),.BLN(BLN45),.WL(WL192));
sram_cell_6t_5 inst_cell_192_46 (.BL(BL46),.BLN(BLN46),.WL(WL192));
sram_cell_6t_5 inst_cell_192_47 (.BL(BL47),.BLN(BLN47),.WL(WL192));
sram_cell_6t_5 inst_cell_192_48 (.BL(BL48),.BLN(BLN48),.WL(WL192));
sram_cell_6t_5 inst_cell_192_49 (.BL(BL49),.BLN(BLN49),.WL(WL192));
sram_cell_6t_5 inst_cell_192_50 (.BL(BL50),.BLN(BLN50),.WL(WL192));
sram_cell_6t_5 inst_cell_192_51 (.BL(BL51),.BLN(BLN51),.WL(WL192));
sram_cell_6t_5 inst_cell_192_52 (.BL(BL52),.BLN(BLN52),.WL(WL192));
sram_cell_6t_5 inst_cell_192_53 (.BL(BL53),.BLN(BLN53),.WL(WL192));
sram_cell_6t_5 inst_cell_192_54 (.BL(BL54),.BLN(BLN54),.WL(WL192));
sram_cell_6t_5 inst_cell_192_55 (.BL(BL55),.BLN(BLN55),.WL(WL192));
sram_cell_6t_5 inst_cell_192_56 (.BL(BL56),.BLN(BLN56),.WL(WL192));
sram_cell_6t_5 inst_cell_192_57 (.BL(BL57),.BLN(BLN57),.WL(WL192));
sram_cell_6t_5 inst_cell_192_58 (.BL(BL58),.BLN(BLN58),.WL(WL192));
sram_cell_6t_5 inst_cell_192_59 (.BL(BL59),.BLN(BLN59),.WL(WL192));
sram_cell_6t_5 inst_cell_192_60 (.BL(BL60),.BLN(BLN60),.WL(WL192));
sram_cell_6t_5 inst_cell_192_61 (.BL(BL61),.BLN(BLN61),.WL(WL192));
sram_cell_6t_5 inst_cell_192_62 (.BL(BL62),.BLN(BLN62),.WL(WL192));
sram_cell_6t_5 inst_cell_192_63 (.BL(BL63),.BLN(BLN63),.WL(WL192));
sram_cell_6t_5 inst_cell_192_64 (.BL(BL64),.BLN(BLN64),.WL(WL192));
sram_cell_6t_5 inst_cell_192_65 (.BL(BL65),.BLN(BLN65),.WL(WL192));
sram_cell_6t_5 inst_cell_192_66 (.BL(BL66),.BLN(BLN66),.WL(WL192));
sram_cell_6t_5 inst_cell_192_67 (.BL(BL67),.BLN(BLN67),.WL(WL192));
sram_cell_6t_5 inst_cell_192_68 (.BL(BL68),.BLN(BLN68),.WL(WL192));
sram_cell_6t_5 inst_cell_192_69 (.BL(BL69),.BLN(BLN69),.WL(WL192));
sram_cell_6t_5 inst_cell_192_70 (.BL(BL70),.BLN(BLN70),.WL(WL192));
sram_cell_6t_5 inst_cell_192_71 (.BL(BL71),.BLN(BLN71),.WL(WL192));
sram_cell_6t_5 inst_cell_192_72 (.BL(BL72),.BLN(BLN72),.WL(WL192));
sram_cell_6t_5 inst_cell_192_73 (.BL(BL73),.BLN(BLN73),.WL(WL192));
sram_cell_6t_5 inst_cell_192_74 (.BL(BL74),.BLN(BLN74),.WL(WL192));
sram_cell_6t_5 inst_cell_192_75 (.BL(BL75),.BLN(BLN75),.WL(WL192));
sram_cell_6t_5 inst_cell_192_76 (.BL(BL76),.BLN(BLN76),.WL(WL192));
sram_cell_6t_5 inst_cell_192_77 (.BL(BL77),.BLN(BLN77),.WL(WL192));
sram_cell_6t_5 inst_cell_192_78 (.BL(BL78),.BLN(BLN78),.WL(WL192));
sram_cell_6t_5 inst_cell_192_79 (.BL(BL79),.BLN(BLN79),.WL(WL192));
sram_cell_6t_5 inst_cell_192_80 (.BL(BL80),.BLN(BLN80),.WL(WL192));
sram_cell_6t_5 inst_cell_192_81 (.BL(BL81),.BLN(BLN81),.WL(WL192));
sram_cell_6t_5 inst_cell_192_82 (.BL(BL82),.BLN(BLN82),.WL(WL192));
sram_cell_6t_5 inst_cell_192_83 (.BL(BL83),.BLN(BLN83),.WL(WL192));
sram_cell_6t_5 inst_cell_192_84 (.BL(BL84),.BLN(BLN84),.WL(WL192));
sram_cell_6t_5 inst_cell_192_85 (.BL(BL85),.BLN(BLN85),.WL(WL192));
sram_cell_6t_5 inst_cell_192_86 (.BL(BL86),.BLN(BLN86),.WL(WL192));
sram_cell_6t_5 inst_cell_192_87 (.BL(BL87),.BLN(BLN87),.WL(WL192));
sram_cell_6t_5 inst_cell_192_88 (.BL(BL88),.BLN(BLN88),.WL(WL192));
sram_cell_6t_5 inst_cell_192_89 (.BL(BL89),.BLN(BLN89),.WL(WL192));
sram_cell_6t_5 inst_cell_192_90 (.BL(BL90),.BLN(BLN90),.WL(WL192));
sram_cell_6t_5 inst_cell_192_91 (.BL(BL91),.BLN(BLN91),.WL(WL192));
sram_cell_6t_5 inst_cell_192_92 (.BL(BL92),.BLN(BLN92),.WL(WL192));
sram_cell_6t_5 inst_cell_192_93 (.BL(BL93),.BLN(BLN93),.WL(WL192));
sram_cell_6t_5 inst_cell_192_94 (.BL(BL94),.BLN(BLN94),.WL(WL192));
sram_cell_6t_5 inst_cell_192_95 (.BL(BL95),.BLN(BLN95),.WL(WL192));
sram_cell_6t_5 inst_cell_192_96 (.BL(BL96),.BLN(BLN96),.WL(WL192));
sram_cell_6t_5 inst_cell_192_97 (.BL(BL97),.BLN(BLN97),.WL(WL192));
sram_cell_6t_5 inst_cell_192_98 (.BL(BL98),.BLN(BLN98),.WL(WL192));
sram_cell_6t_5 inst_cell_192_99 (.BL(BL99),.BLN(BLN99),.WL(WL192));
sram_cell_6t_5 inst_cell_192_100 (.BL(BL100),.BLN(BLN100),.WL(WL192));
sram_cell_6t_5 inst_cell_192_101 (.BL(BL101),.BLN(BLN101),.WL(WL192));
sram_cell_6t_5 inst_cell_192_102 (.BL(BL102),.BLN(BLN102),.WL(WL192));
sram_cell_6t_5 inst_cell_192_103 (.BL(BL103),.BLN(BLN103),.WL(WL192));
sram_cell_6t_5 inst_cell_192_104 (.BL(BL104),.BLN(BLN104),.WL(WL192));
sram_cell_6t_5 inst_cell_192_105 (.BL(BL105),.BLN(BLN105),.WL(WL192));
sram_cell_6t_5 inst_cell_192_106 (.BL(BL106),.BLN(BLN106),.WL(WL192));
sram_cell_6t_5 inst_cell_192_107 (.BL(BL107),.BLN(BLN107),.WL(WL192));
sram_cell_6t_5 inst_cell_192_108 (.BL(BL108),.BLN(BLN108),.WL(WL192));
sram_cell_6t_5 inst_cell_192_109 (.BL(BL109),.BLN(BLN109),.WL(WL192));
sram_cell_6t_5 inst_cell_192_110 (.BL(BL110),.BLN(BLN110),.WL(WL192));
sram_cell_6t_5 inst_cell_192_111 (.BL(BL111),.BLN(BLN111),.WL(WL192));
sram_cell_6t_5 inst_cell_192_112 (.BL(BL112),.BLN(BLN112),.WL(WL192));
sram_cell_6t_5 inst_cell_192_113 (.BL(BL113),.BLN(BLN113),.WL(WL192));
sram_cell_6t_5 inst_cell_192_114 (.BL(BL114),.BLN(BLN114),.WL(WL192));
sram_cell_6t_5 inst_cell_192_115 (.BL(BL115),.BLN(BLN115),.WL(WL192));
sram_cell_6t_5 inst_cell_192_116 (.BL(BL116),.BLN(BLN116),.WL(WL192));
sram_cell_6t_5 inst_cell_192_117 (.BL(BL117),.BLN(BLN117),.WL(WL192));
sram_cell_6t_5 inst_cell_192_118 (.BL(BL118),.BLN(BLN118),.WL(WL192));
sram_cell_6t_5 inst_cell_192_119 (.BL(BL119),.BLN(BLN119),.WL(WL192));
sram_cell_6t_5 inst_cell_192_120 (.BL(BL120),.BLN(BLN120),.WL(WL192));
sram_cell_6t_5 inst_cell_192_121 (.BL(BL121),.BLN(BLN121),.WL(WL192));
sram_cell_6t_5 inst_cell_192_122 (.BL(BL122),.BLN(BLN122),.WL(WL192));
sram_cell_6t_5 inst_cell_192_123 (.BL(BL123),.BLN(BLN123),.WL(WL192));
sram_cell_6t_5 inst_cell_192_124 (.BL(BL124),.BLN(BLN124),.WL(WL192));
sram_cell_6t_5 inst_cell_192_125 (.BL(BL125),.BLN(BLN125),.WL(WL192));
sram_cell_6t_5 inst_cell_192_126 (.BL(BL126),.BLN(BLN126),.WL(WL192));
sram_cell_6t_5 inst_cell_192_127 (.BL(BL127),.BLN(BLN127),.WL(WL192));
sram_cell_6t_5 inst_cell_193_0 (.BL(BL0),.BLN(BLN0),.WL(WL193));
sram_cell_6t_5 inst_cell_193_1 (.BL(BL1),.BLN(BLN1),.WL(WL193));
sram_cell_6t_5 inst_cell_193_2 (.BL(BL2),.BLN(BLN2),.WL(WL193));
sram_cell_6t_5 inst_cell_193_3 (.BL(BL3),.BLN(BLN3),.WL(WL193));
sram_cell_6t_5 inst_cell_193_4 (.BL(BL4),.BLN(BLN4),.WL(WL193));
sram_cell_6t_5 inst_cell_193_5 (.BL(BL5),.BLN(BLN5),.WL(WL193));
sram_cell_6t_5 inst_cell_193_6 (.BL(BL6),.BLN(BLN6),.WL(WL193));
sram_cell_6t_5 inst_cell_193_7 (.BL(BL7),.BLN(BLN7),.WL(WL193));
sram_cell_6t_5 inst_cell_193_8 (.BL(BL8),.BLN(BLN8),.WL(WL193));
sram_cell_6t_5 inst_cell_193_9 (.BL(BL9),.BLN(BLN9),.WL(WL193));
sram_cell_6t_5 inst_cell_193_10 (.BL(BL10),.BLN(BLN10),.WL(WL193));
sram_cell_6t_5 inst_cell_193_11 (.BL(BL11),.BLN(BLN11),.WL(WL193));
sram_cell_6t_5 inst_cell_193_12 (.BL(BL12),.BLN(BLN12),.WL(WL193));
sram_cell_6t_5 inst_cell_193_13 (.BL(BL13),.BLN(BLN13),.WL(WL193));
sram_cell_6t_5 inst_cell_193_14 (.BL(BL14),.BLN(BLN14),.WL(WL193));
sram_cell_6t_5 inst_cell_193_15 (.BL(BL15),.BLN(BLN15),.WL(WL193));
sram_cell_6t_5 inst_cell_193_16 (.BL(BL16),.BLN(BLN16),.WL(WL193));
sram_cell_6t_5 inst_cell_193_17 (.BL(BL17),.BLN(BLN17),.WL(WL193));
sram_cell_6t_5 inst_cell_193_18 (.BL(BL18),.BLN(BLN18),.WL(WL193));
sram_cell_6t_5 inst_cell_193_19 (.BL(BL19),.BLN(BLN19),.WL(WL193));
sram_cell_6t_5 inst_cell_193_20 (.BL(BL20),.BLN(BLN20),.WL(WL193));
sram_cell_6t_5 inst_cell_193_21 (.BL(BL21),.BLN(BLN21),.WL(WL193));
sram_cell_6t_5 inst_cell_193_22 (.BL(BL22),.BLN(BLN22),.WL(WL193));
sram_cell_6t_5 inst_cell_193_23 (.BL(BL23),.BLN(BLN23),.WL(WL193));
sram_cell_6t_5 inst_cell_193_24 (.BL(BL24),.BLN(BLN24),.WL(WL193));
sram_cell_6t_5 inst_cell_193_25 (.BL(BL25),.BLN(BLN25),.WL(WL193));
sram_cell_6t_5 inst_cell_193_26 (.BL(BL26),.BLN(BLN26),.WL(WL193));
sram_cell_6t_5 inst_cell_193_27 (.BL(BL27),.BLN(BLN27),.WL(WL193));
sram_cell_6t_5 inst_cell_193_28 (.BL(BL28),.BLN(BLN28),.WL(WL193));
sram_cell_6t_5 inst_cell_193_29 (.BL(BL29),.BLN(BLN29),.WL(WL193));
sram_cell_6t_5 inst_cell_193_30 (.BL(BL30),.BLN(BLN30),.WL(WL193));
sram_cell_6t_5 inst_cell_193_31 (.BL(BL31),.BLN(BLN31),.WL(WL193));
sram_cell_6t_5 inst_cell_193_32 (.BL(BL32),.BLN(BLN32),.WL(WL193));
sram_cell_6t_5 inst_cell_193_33 (.BL(BL33),.BLN(BLN33),.WL(WL193));
sram_cell_6t_5 inst_cell_193_34 (.BL(BL34),.BLN(BLN34),.WL(WL193));
sram_cell_6t_5 inst_cell_193_35 (.BL(BL35),.BLN(BLN35),.WL(WL193));
sram_cell_6t_5 inst_cell_193_36 (.BL(BL36),.BLN(BLN36),.WL(WL193));
sram_cell_6t_5 inst_cell_193_37 (.BL(BL37),.BLN(BLN37),.WL(WL193));
sram_cell_6t_5 inst_cell_193_38 (.BL(BL38),.BLN(BLN38),.WL(WL193));
sram_cell_6t_5 inst_cell_193_39 (.BL(BL39),.BLN(BLN39),.WL(WL193));
sram_cell_6t_5 inst_cell_193_40 (.BL(BL40),.BLN(BLN40),.WL(WL193));
sram_cell_6t_5 inst_cell_193_41 (.BL(BL41),.BLN(BLN41),.WL(WL193));
sram_cell_6t_5 inst_cell_193_42 (.BL(BL42),.BLN(BLN42),.WL(WL193));
sram_cell_6t_5 inst_cell_193_43 (.BL(BL43),.BLN(BLN43),.WL(WL193));
sram_cell_6t_5 inst_cell_193_44 (.BL(BL44),.BLN(BLN44),.WL(WL193));
sram_cell_6t_5 inst_cell_193_45 (.BL(BL45),.BLN(BLN45),.WL(WL193));
sram_cell_6t_5 inst_cell_193_46 (.BL(BL46),.BLN(BLN46),.WL(WL193));
sram_cell_6t_5 inst_cell_193_47 (.BL(BL47),.BLN(BLN47),.WL(WL193));
sram_cell_6t_5 inst_cell_193_48 (.BL(BL48),.BLN(BLN48),.WL(WL193));
sram_cell_6t_5 inst_cell_193_49 (.BL(BL49),.BLN(BLN49),.WL(WL193));
sram_cell_6t_5 inst_cell_193_50 (.BL(BL50),.BLN(BLN50),.WL(WL193));
sram_cell_6t_5 inst_cell_193_51 (.BL(BL51),.BLN(BLN51),.WL(WL193));
sram_cell_6t_5 inst_cell_193_52 (.BL(BL52),.BLN(BLN52),.WL(WL193));
sram_cell_6t_5 inst_cell_193_53 (.BL(BL53),.BLN(BLN53),.WL(WL193));
sram_cell_6t_5 inst_cell_193_54 (.BL(BL54),.BLN(BLN54),.WL(WL193));
sram_cell_6t_5 inst_cell_193_55 (.BL(BL55),.BLN(BLN55),.WL(WL193));
sram_cell_6t_5 inst_cell_193_56 (.BL(BL56),.BLN(BLN56),.WL(WL193));
sram_cell_6t_5 inst_cell_193_57 (.BL(BL57),.BLN(BLN57),.WL(WL193));
sram_cell_6t_5 inst_cell_193_58 (.BL(BL58),.BLN(BLN58),.WL(WL193));
sram_cell_6t_5 inst_cell_193_59 (.BL(BL59),.BLN(BLN59),.WL(WL193));
sram_cell_6t_5 inst_cell_193_60 (.BL(BL60),.BLN(BLN60),.WL(WL193));
sram_cell_6t_5 inst_cell_193_61 (.BL(BL61),.BLN(BLN61),.WL(WL193));
sram_cell_6t_5 inst_cell_193_62 (.BL(BL62),.BLN(BLN62),.WL(WL193));
sram_cell_6t_5 inst_cell_193_63 (.BL(BL63),.BLN(BLN63),.WL(WL193));
sram_cell_6t_5 inst_cell_193_64 (.BL(BL64),.BLN(BLN64),.WL(WL193));
sram_cell_6t_5 inst_cell_193_65 (.BL(BL65),.BLN(BLN65),.WL(WL193));
sram_cell_6t_5 inst_cell_193_66 (.BL(BL66),.BLN(BLN66),.WL(WL193));
sram_cell_6t_5 inst_cell_193_67 (.BL(BL67),.BLN(BLN67),.WL(WL193));
sram_cell_6t_5 inst_cell_193_68 (.BL(BL68),.BLN(BLN68),.WL(WL193));
sram_cell_6t_5 inst_cell_193_69 (.BL(BL69),.BLN(BLN69),.WL(WL193));
sram_cell_6t_5 inst_cell_193_70 (.BL(BL70),.BLN(BLN70),.WL(WL193));
sram_cell_6t_5 inst_cell_193_71 (.BL(BL71),.BLN(BLN71),.WL(WL193));
sram_cell_6t_5 inst_cell_193_72 (.BL(BL72),.BLN(BLN72),.WL(WL193));
sram_cell_6t_5 inst_cell_193_73 (.BL(BL73),.BLN(BLN73),.WL(WL193));
sram_cell_6t_5 inst_cell_193_74 (.BL(BL74),.BLN(BLN74),.WL(WL193));
sram_cell_6t_5 inst_cell_193_75 (.BL(BL75),.BLN(BLN75),.WL(WL193));
sram_cell_6t_5 inst_cell_193_76 (.BL(BL76),.BLN(BLN76),.WL(WL193));
sram_cell_6t_5 inst_cell_193_77 (.BL(BL77),.BLN(BLN77),.WL(WL193));
sram_cell_6t_5 inst_cell_193_78 (.BL(BL78),.BLN(BLN78),.WL(WL193));
sram_cell_6t_5 inst_cell_193_79 (.BL(BL79),.BLN(BLN79),.WL(WL193));
sram_cell_6t_5 inst_cell_193_80 (.BL(BL80),.BLN(BLN80),.WL(WL193));
sram_cell_6t_5 inst_cell_193_81 (.BL(BL81),.BLN(BLN81),.WL(WL193));
sram_cell_6t_5 inst_cell_193_82 (.BL(BL82),.BLN(BLN82),.WL(WL193));
sram_cell_6t_5 inst_cell_193_83 (.BL(BL83),.BLN(BLN83),.WL(WL193));
sram_cell_6t_5 inst_cell_193_84 (.BL(BL84),.BLN(BLN84),.WL(WL193));
sram_cell_6t_5 inst_cell_193_85 (.BL(BL85),.BLN(BLN85),.WL(WL193));
sram_cell_6t_5 inst_cell_193_86 (.BL(BL86),.BLN(BLN86),.WL(WL193));
sram_cell_6t_5 inst_cell_193_87 (.BL(BL87),.BLN(BLN87),.WL(WL193));
sram_cell_6t_5 inst_cell_193_88 (.BL(BL88),.BLN(BLN88),.WL(WL193));
sram_cell_6t_5 inst_cell_193_89 (.BL(BL89),.BLN(BLN89),.WL(WL193));
sram_cell_6t_5 inst_cell_193_90 (.BL(BL90),.BLN(BLN90),.WL(WL193));
sram_cell_6t_5 inst_cell_193_91 (.BL(BL91),.BLN(BLN91),.WL(WL193));
sram_cell_6t_5 inst_cell_193_92 (.BL(BL92),.BLN(BLN92),.WL(WL193));
sram_cell_6t_5 inst_cell_193_93 (.BL(BL93),.BLN(BLN93),.WL(WL193));
sram_cell_6t_5 inst_cell_193_94 (.BL(BL94),.BLN(BLN94),.WL(WL193));
sram_cell_6t_5 inst_cell_193_95 (.BL(BL95),.BLN(BLN95),.WL(WL193));
sram_cell_6t_5 inst_cell_193_96 (.BL(BL96),.BLN(BLN96),.WL(WL193));
sram_cell_6t_5 inst_cell_193_97 (.BL(BL97),.BLN(BLN97),.WL(WL193));
sram_cell_6t_5 inst_cell_193_98 (.BL(BL98),.BLN(BLN98),.WL(WL193));
sram_cell_6t_5 inst_cell_193_99 (.BL(BL99),.BLN(BLN99),.WL(WL193));
sram_cell_6t_5 inst_cell_193_100 (.BL(BL100),.BLN(BLN100),.WL(WL193));
sram_cell_6t_5 inst_cell_193_101 (.BL(BL101),.BLN(BLN101),.WL(WL193));
sram_cell_6t_5 inst_cell_193_102 (.BL(BL102),.BLN(BLN102),.WL(WL193));
sram_cell_6t_5 inst_cell_193_103 (.BL(BL103),.BLN(BLN103),.WL(WL193));
sram_cell_6t_5 inst_cell_193_104 (.BL(BL104),.BLN(BLN104),.WL(WL193));
sram_cell_6t_5 inst_cell_193_105 (.BL(BL105),.BLN(BLN105),.WL(WL193));
sram_cell_6t_5 inst_cell_193_106 (.BL(BL106),.BLN(BLN106),.WL(WL193));
sram_cell_6t_5 inst_cell_193_107 (.BL(BL107),.BLN(BLN107),.WL(WL193));
sram_cell_6t_5 inst_cell_193_108 (.BL(BL108),.BLN(BLN108),.WL(WL193));
sram_cell_6t_5 inst_cell_193_109 (.BL(BL109),.BLN(BLN109),.WL(WL193));
sram_cell_6t_5 inst_cell_193_110 (.BL(BL110),.BLN(BLN110),.WL(WL193));
sram_cell_6t_5 inst_cell_193_111 (.BL(BL111),.BLN(BLN111),.WL(WL193));
sram_cell_6t_5 inst_cell_193_112 (.BL(BL112),.BLN(BLN112),.WL(WL193));
sram_cell_6t_5 inst_cell_193_113 (.BL(BL113),.BLN(BLN113),.WL(WL193));
sram_cell_6t_5 inst_cell_193_114 (.BL(BL114),.BLN(BLN114),.WL(WL193));
sram_cell_6t_5 inst_cell_193_115 (.BL(BL115),.BLN(BLN115),.WL(WL193));
sram_cell_6t_5 inst_cell_193_116 (.BL(BL116),.BLN(BLN116),.WL(WL193));
sram_cell_6t_5 inst_cell_193_117 (.BL(BL117),.BLN(BLN117),.WL(WL193));
sram_cell_6t_5 inst_cell_193_118 (.BL(BL118),.BLN(BLN118),.WL(WL193));
sram_cell_6t_5 inst_cell_193_119 (.BL(BL119),.BLN(BLN119),.WL(WL193));
sram_cell_6t_5 inst_cell_193_120 (.BL(BL120),.BLN(BLN120),.WL(WL193));
sram_cell_6t_5 inst_cell_193_121 (.BL(BL121),.BLN(BLN121),.WL(WL193));
sram_cell_6t_5 inst_cell_193_122 (.BL(BL122),.BLN(BLN122),.WL(WL193));
sram_cell_6t_5 inst_cell_193_123 (.BL(BL123),.BLN(BLN123),.WL(WL193));
sram_cell_6t_5 inst_cell_193_124 (.BL(BL124),.BLN(BLN124),.WL(WL193));
sram_cell_6t_5 inst_cell_193_125 (.BL(BL125),.BLN(BLN125),.WL(WL193));
sram_cell_6t_5 inst_cell_193_126 (.BL(BL126),.BLN(BLN126),.WL(WL193));
sram_cell_6t_5 inst_cell_193_127 (.BL(BL127),.BLN(BLN127),.WL(WL193));
sram_cell_6t_5 inst_cell_194_0 (.BL(BL0),.BLN(BLN0),.WL(WL194));
sram_cell_6t_5 inst_cell_194_1 (.BL(BL1),.BLN(BLN1),.WL(WL194));
sram_cell_6t_5 inst_cell_194_2 (.BL(BL2),.BLN(BLN2),.WL(WL194));
sram_cell_6t_5 inst_cell_194_3 (.BL(BL3),.BLN(BLN3),.WL(WL194));
sram_cell_6t_5 inst_cell_194_4 (.BL(BL4),.BLN(BLN4),.WL(WL194));
sram_cell_6t_5 inst_cell_194_5 (.BL(BL5),.BLN(BLN5),.WL(WL194));
sram_cell_6t_5 inst_cell_194_6 (.BL(BL6),.BLN(BLN6),.WL(WL194));
sram_cell_6t_5 inst_cell_194_7 (.BL(BL7),.BLN(BLN7),.WL(WL194));
sram_cell_6t_5 inst_cell_194_8 (.BL(BL8),.BLN(BLN8),.WL(WL194));
sram_cell_6t_5 inst_cell_194_9 (.BL(BL9),.BLN(BLN9),.WL(WL194));
sram_cell_6t_5 inst_cell_194_10 (.BL(BL10),.BLN(BLN10),.WL(WL194));
sram_cell_6t_5 inst_cell_194_11 (.BL(BL11),.BLN(BLN11),.WL(WL194));
sram_cell_6t_5 inst_cell_194_12 (.BL(BL12),.BLN(BLN12),.WL(WL194));
sram_cell_6t_5 inst_cell_194_13 (.BL(BL13),.BLN(BLN13),.WL(WL194));
sram_cell_6t_5 inst_cell_194_14 (.BL(BL14),.BLN(BLN14),.WL(WL194));
sram_cell_6t_5 inst_cell_194_15 (.BL(BL15),.BLN(BLN15),.WL(WL194));
sram_cell_6t_5 inst_cell_194_16 (.BL(BL16),.BLN(BLN16),.WL(WL194));
sram_cell_6t_5 inst_cell_194_17 (.BL(BL17),.BLN(BLN17),.WL(WL194));
sram_cell_6t_5 inst_cell_194_18 (.BL(BL18),.BLN(BLN18),.WL(WL194));
sram_cell_6t_5 inst_cell_194_19 (.BL(BL19),.BLN(BLN19),.WL(WL194));
sram_cell_6t_5 inst_cell_194_20 (.BL(BL20),.BLN(BLN20),.WL(WL194));
sram_cell_6t_5 inst_cell_194_21 (.BL(BL21),.BLN(BLN21),.WL(WL194));
sram_cell_6t_5 inst_cell_194_22 (.BL(BL22),.BLN(BLN22),.WL(WL194));
sram_cell_6t_5 inst_cell_194_23 (.BL(BL23),.BLN(BLN23),.WL(WL194));
sram_cell_6t_5 inst_cell_194_24 (.BL(BL24),.BLN(BLN24),.WL(WL194));
sram_cell_6t_5 inst_cell_194_25 (.BL(BL25),.BLN(BLN25),.WL(WL194));
sram_cell_6t_5 inst_cell_194_26 (.BL(BL26),.BLN(BLN26),.WL(WL194));
sram_cell_6t_5 inst_cell_194_27 (.BL(BL27),.BLN(BLN27),.WL(WL194));
sram_cell_6t_5 inst_cell_194_28 (.BL(BL28),.BLN(BLN28),.WL(WL194));
sram_cell_6t_5 inst_cell_194_29 (.BL(BL29),.BLN(BLN29),.WL(WL194));
sram_cell_6t_5 inst_cell_194_30 (.BL(BL30),.BLN(BLN30),.WL(WL194));
sram_cell_6t_5 inst_cell_194_31 (.BL(BL31),.BLN(BLN31),.WL(WL194));
sram_cell_6t_5 inst_cell_194_32 (.BL(BL32),.BLN(BLN32),.WL(WL194));
sram_cell_6t_5 inst_cell_194_33 (.BL(BL33),.BLN(BLN33),.WL(WL194));
sram_cell_6t_5 inst_cell_194_34 (.BL(BL34),.BLN(BLN34),.WL(WL194));
sram_cell_6t_5 inst_cell_194_35 (.BL(BL35),.BLN(BLN35),.WL(WL194));
sram_cell_6t_5 inst_cell_194_36 (.BL(BL36),.BLN(BLN36),.WL(WL194));
sram_cell_6t_5 inst_cell_194_37 (.BL(BL37),.BLN(BLN37),.WL(WL194));
sram_cell_6t_5 inst_cell_194_38 (.BL(BL38),.BLN(BLN38),.WL(WL194));
sram_cell_6t_5 inst_cell_194_39 (.BL(BL39),.BLN(BLN39),.WL(WL194));
sram_cell_6t_5 inst_cell_194_40 (.BL(BL40),.BLN(BLN40),.WL(WL194));
sram_cell_6t_5 inst_cell_194_41 (.BL(BL41),.BLN(BLN41),.WL(WL194));
sram_cell_6t_5 inst_cell_194_42 (.BL(BL42),.BLN(BLN42),.WL(WL194));
sram_cell_6t_5 inst_cell_194_43 (.BL(BL43),.BLN(BLN43),.WL(WL194));
sram_cell_6t_5 inst_cell_194_44 (.BL(BL44),.BLN(BLN44),.WL(WL194));
sram_cell_6t_5 inst_cell_194_45 (.BL(BL45),.BLN(BLN45),.WL(WL194));
sram_cell_6t_5 inst_cell_194_46 (.BL(BL46),.BLN(BLN46),.WL(WL194));
sram_cell_6t_5 inst_cell_194_47 (.BL(BL47),.BLN(BLN47),.WL(WL194));
sram_cell_6t_5 inst_cell_194_48 (.BL(BL48),.BLN(BLN48),.WL(WL194));
sram_cell_6t_5 inst_cell_194_49 (.BL(BL49),.BLN(BLN49),.WL(WL194));
sram_cell_6t_5 inst_cell_194_50 (.BL(BL50),.BLN(BLN50),.WL(WL194));
sram_cell_6t_5 inst_cell_194_51 (.BL(BL51),.BLN(BLN51),.WL(WL194));
sram_cell_6t_5 inst_cell_194_52 (.BL(BL52),.BLN(BLN52),.WL(WL194));
sram_cell_6t_5 inst_cell_194_53 (.BL(BL53),.BLN(BLN53),.WL(WL194));
sram_cell_6t_5 inst_cell_194_54 (.BL(BL54),.BLN(BLN54),.WL(WL194));
sram_cell_6t_5 inst_cell_194_55 (.BL(BL55),.BLN(BLN55),.WL(WL194));
sram_cell_6t_5 inst_cell_194_56 (.BL(BL56),.BLN(BLN56),.WL(WL194));
sram_cell_6t_5 inst_cell_194_57 (.BL(BL57),.BLN(BLN57),.WL(WL194));
sram_cell_6t_5 inst_cell_194_58 (.BL(BL58),.BLN(BLN58),.WL(WL194));
sram_cell_6t_5 inst_cell_194_59 (.BL(BL59),.BLN(BLN59),.WL(WL194));
sram_cell_6t_5 inst_cell_194_60 (.BL(BL60),.BLN(BLN60),.WL(WL194));
sram_cell_6t_5 inst_cell_194_61 (.BL(BL61),.BLN(BLN61),.WL(WL194));
sram_cell_6t_5 inst_cell_194_62 (.BL(BL62),.BLN(BLN62),.WL(WL194));
sram_cell_6t_5 inst_cell_194_63 (.BL(BL63),.BLN(BLN63),.WL(WL194));
sram_cell_6t_5 inst_cell_194_64 (.BL(BL64),.BLN(BLN64),.WL(WL194));
sram_cell_6t_5 inst_cell_194_65 (.BL(BL65),.BLN(BLN65),.WL(WL194));
sram_cell_6t_5 inst_cell_194_66 (.BL(BL66),.BLN(BLN66),.WL(WL194));
sram_cell_6t_5 inst_cell_194_67 (.BL(BL67),.BLN(BLN67),.WL(WL194));
sram_cell_6t_5 inst_cell_194_68 (.BL(BL68),.BLN(BLN68),.WL(WL194));
sram_cell_6t_5 inst_cell_194_69 (.BL(BL69),.BLN(BLN69),.WL(WL194));
sram_cell_6t_5 inst_cell_194_70 (.BL(BL70),.BLN(BLN70),.WL(WL194));
sram_cell_6t_5 inst_cell_194_71 (.BL(BL71),.BLN(BLN71),.WL(WL194));
sram_cell_6t_5 inst_cell_194_72 (.BL(BL72),.BLN(BLN72),.WL(WL194));
sram_cell_6t_5 inst_cell_194_73 (.BL(BL73),.BLN(BLN73),.WL(WL194));
sram_cell_6t_5 inst_cell_194_74 (.BL(BL74),.BLN(BLN74),.WL(WL194));
sram_cell_6t_5 inst_cell_194_75 (.BL(BL75),.BLN(BLN75),.WL(WL194));
sram_cell_6t_5 inst_cell_194_76 (.BL(BL76),.BLN(BLN76),.WL(WL194));
sram_cell_6t_5 inst_cell_194_77 (.BL(BL77),.BLN(BLN77),.WL(WL194));
sram_cell_6t_5 inst_cell_194_78 (.BL(BL78),.BLN(BLN78),.WL(WL194));
sram_cell_6t_5 inst_cell_194_79 (.BL(BL79),.BLN(BLN79),.WL(WL194));
sram_cell_6t_5 inst_cell_194_80 (.BL(BL80),.BLN(BLN80),.WL(WL194));
sram_cell_6t_5 inst_cell_194_81 (.BL(BL81),.BLN(BLN81),.WL(WL194));
sram_cell_6t_5 inst_cell_194_82 (.BL(BL82),.BLN(BLN82),.WL(WL194));
sram_cell_6t_5 inst_cell_194_83 (.BL(BL83),.BLN(BLN83),.WL(WL194));
sram_cell_6t_5 inst_cell_194_84 (.BL(BL84),.BLN(BLN84),.WL(WL194));
sram_cell_6t_5 inst_cell_194_85 (.BL(BL85),.BLN(BLN85),.WL(WL194));
sram_cell_6t_5 inst_cell_194_86 (.BL(BL86),.BLN(BLN86),.WL(WL194));
sram_cell_6t_5 inst_cell_194_87 (.BL(BL87),.BLN(BLN87),.WL(WL194));
sram_cell_6t_5 inst_cell_194_88 (.BL(BL88),.BLN(BLN88),.WL(WL194));
sram_cell_6t_5 inst_cell_194_89 (.BL(BL89),.BLN(BLN89),.WL(WL194));
sram_cell_6t_5 inst_cell_194_90 (.BL(BL90),.BLN(BLN90),.WL(WL194));
sram_cell_6t_5 inst_cell_194_91 (.BL(BL91),.BLN(BLN91),.WL(WL194));
sram_cell_6t_5 inst_cell_194_92 (.BL(BL92),.BLN(BLN92),.WL(WL194));
sram_cell_6t_5 inst_cell_194_93 (.BL(BL93),.BLN(BLN93),.WL(WL194));
sram_cell_6t_5 inst_cell_194_94 (.BL(BL94),.BLN(BLN94),.WL(WL194));
sram_cell_6t_5 inst_cell_194_95 (.BL(BL95),.BLN(BLN95),.WL(WL194));
sram_cell_6t_5 inst_cell_194_96 (.BL(BL96),.BLN(BLN96),.WL(WL194));
sram_cell_6t_5 inst_cell_194_97 (.BL(BL97),.BLN(BLN97),.WL(WL194));
sram_cell_6t_5 inst_cell_194_98 (.BL(BL98),.BLN(BLN98),.WL(WL194));
sram_cell_6t_5 inst_cell_194_99 (.BL(BL99),.BLN(BLN99),.WL(WL194));
sram_cell_6t_5 inst_cell_194_100 (.BL(BL100),.BLN(BLN100),.WL(WL194));
sram_cell_6t_5 inst_cell_194_101 (.BL(BL101),.BLN(BLN101),.WL(WL194));
sram_cell_6t_5 inst_cell_194_102 (.BL(BL102),.BLN(BLN102),.WL(WL194));
sram_cell_6t_5 inst_cell_194_103 (.BL(BL103),.BLN(BLN103),.WL(WL194));
sram_cell_6t_5 inst_cell_194_104 (.BL(BL104),.BLN(BLN104),.WL(WL194));
sram_cell_6t_5 inst_cell_194_105 (.BL(BL105),.BLN(BLN105),.WL(WL194));
sram_cell_6t_5 inst_cell_194_106 (.BL(BL106),.BLN(BLN106),.WL(WL194));
sram_cell_6t_5 inst_cell_194_107 (.BL(BL107),.BLN(BLN107),.WL(WL194));
sram_cell_6t_5 inst_cell_194_108 (.BL(BL108),.BLN(BLN108),.WL(WL194));
sram_cell_6t_5 inst_cell_194_109 (.BL(BL109),.BLN(BLN109),.WL(WL194));
sram_cell_6t_5 inst_cell_194_110 (.BL(BL110),.BLN(BLN110),.WL(WL194));
sram_cell_6t_5 inst_cell_194_111 (.BL(BL111),.BLN(BLN111),.WL(WL194));
sram_cell_6t_5 inst_cell_194_112 (.BL(BL112),.BLN(BLN112),.WL(WL194));
sram_cell_6t_5 inst_cell_194_113 (.BL(BL113),.BLN(BLN113),.WL(WL194));
sram_cell_6t_5 inst_cell_194_114 (.BL(BL114),.BLN(BLN114),.WL(WL194));
sram_cell_6t_5 inst_cell_194_115 (.BL(BL115),.BLN(BLN115),.WL(WL194));
sram_cell_6t_5 inst_cell_194_116 (.BL(BL116),.BLN(BLN116),.WL(WL194));
sram_cell_6t_5 inst_cell_194_117 (.BL(BL117),.BLN(BLN117),.WL(WL194));
sram_cell_6t_5 inst_cell_194_118 (.BL(BL118),.BLN(BLN118),.WL(WL194));
sram_cell_6t_5 inst_cell_194_119 (.BL(BL119),.BLN(BLN119),.WL(WL194));
sram_cell_6t_5 inst_cell_194_120 (.BL(BL120),.BLN(BLN120),.WL(WL194));
sram_cell_6t_5 inst_cell_194_121 (.BL(BL121),.BLN(BLN121),.WL(WL194));
sram_cell_6t_5 inst_cell_194_122 (.BL(BL122),.BLN(BLN122),.WL(WL194));
sram_cell_6t_5 inst_cell_194_123 (.BL(BL123),.BLN(BLN123),.WL(WL194));
sram_cell_6t_5 inst_cell_194_124 (.BL(BL124),.BLN(BLN124),.WL(WL194));
sram_cell_6t_5 inst_cell_194_125 (.BL(BL125),.BLN(BLN125),.WL(WL194));
sram_cell_6t_5 inst_cell_194_126 (.BL(BL126),.BLN(BLN126),.WL(WL194));
sram_cell_6t_5 inst_cell_194_127 (.BL(BL127),.BLN(BLN127),.WL(WL194));
sram_cell_6t_5 inst_cell_195_0 (.BL(BL0),.BLN(BLN0),.WL(WL195));
sram_cell_6t_5 inst_cell_195_1 (.BL(BL1),.BLN(BLN1),.WL(WL195));
sram_cell_6t_5 inst_cell_195_2 (.BL(BL2),.BLN(BLN2),.WL(WL195));
sram_cell_6t_5 inst_cell_195_3 (.BL(BL3),.BLN(BLN3),.WL(WL195));
sram_cell_6t_5 inst_cell_195_4 (.BL(BL4),.BLN(BLN4),.WL(WL195));
sram_cell_6t_5 inst_cell_195_5 (.BL(BL5),.BLN(BLN5),.WL(WL195));
sram_cell_6t_5 inst_cell_195_6 (.BL(BL6),.BLN(BLN6),.WL(WL195));
sram_cell_6t_5 inst_cell_195_7 (.BL(BL7),.BLN(BLN7),.WL(WL195));
sram_cell_6t_5 inst_cell_195_8 (.BL(BL8),.BLN(BLN8),.WL(WL195));
sram_cell_6t_5 inst_cell_195_9 (.BL(BL9),.BLN(BLN9),.WL(WL195));
sram_cell_6t_5 inst_cell_195_10 (.BL(BL10),.BLN(BLN10),.WL(WL195));
sram_cell_6t_5 inst_cell_195_11 (.BL(BL11),.BLN(BLN11),.WL(WL195));
sram_cell_6t_5 inst_cell_195_12 (.BL(BL12),.BLN(BLN12),.WL(WL195));
sram_cell_6t_5 inst_cell_195_13 (.BL(BL13),.BLN(BLN13),.WL(WL195));
sram_cell_6t_5 inst_cell_195_14 (.BL(BL14),.BLN(BLN14),.WL(WL195));
sram_cell_6t_5 inst_cell_195_15 (.BL(BL15),.BLN(BLN15),.WL(WL195));
sram_cell_6t_5 inst_cell_195_16 (.BL(BL16),.BLN(BLN16),.WL(WL195));
sram_cell_6t_5 inst_cell_195_17 (.BL(BL17),.BLN(BLN17),.WL(WL195));
sram_cell_6t_5 inst_cell_195_18 (.BL(BL18),.BLN(BLN18),.WL(WL195));
sram_cell_6t_5 inst_cell_195_19 (.BL(BL19),.BLN(BLN19),.WL(WL195));
sram_cell_6t_5 inst_cell_195_20 (.BL(BL20),.BLN(BLN20),.WL(WL195));
sram_cell_6t_5 inst_cell_195_21 (.BL(BL21),.BLN(BLN21),.WL(WL195));
sram_cell_6t_5 inst_cell_195_22 (.BL(BL22),.BLN(BLN22),.WL(WL195));
sram_cell_6t_5 inst_cell_195_23 (.BL(BL23),.BLN(BLN23),.WL(WL195));
sram_cell_6t_5 inst_cell_195_24 (.BL(BL24),.BLN(BLN24),.WL(WL195));
sram_cell_6t_5 inst_cell_195_25 (.BL(BL25),.BLN(BLN25),.WL(WL195));
sram_cell_6t_5 inst_cell_195_26 (.BL(BL26),.BLN(BLN26),.WL(WL195));
sram_cell_6t_5 inst_cell_195_27 (.BL(BL27),.BLN(BLN27),.WL(WL195));
sram_cell_6t_5 inst_cell_195_28 (.BL(BL28),.BLN(BLN28),.WL(WL195));
sram_cell_6t_5 inst_cell_195_29 (.BL(BL29),.BLN(BLN29),.WL(WL195));
sram_cell_6t_5 inst_cell_195_30 (.BL(BL30),.BLN(BLN30),.WL(WL195));
sram_cell_6t_5 inst_cell_195_31 (.BL(BL31),.BLN(BLN31),.WL(WL195));
sram_cell_6t_5 inst_cell_195_32 (.BL(BL32),.BLN(BLN32),.WL(WL195));
sram_cell_6t_5 inst_cell_195_33 (.BL(BL33),.BLN(BLN33),.WL(WL195));
sram_cell_6t_5 inst_cell_195_34 (.BL(BL34),.BLN(BLN34),.WL(WL195));
sram_cell_6t_5 inst_cell_195_35 (.BL(BL35),.BLN(BLN35),.WL(WL195));
sram_cell_6t_5 inst_cell_195_36 (.BL(BL36),.BLN(BLN36),.WL(WL195));
sram_cell_6t_5 inst_cell_195_37 (.BL(BL37),.BLN(BLN37),.WL(WL195));
sram_cell_6t_5 inst_cell_195_38 (.BL(BL38),.BLN(BLN38),.WL(WL195));
sram_cell_6t_5 inst_cell_195_39 (.BL(BL39),.BLN(BLN39),.WL(WL195));
sram_cell_6t_5 inst_cell_195_40 (.BL(BL40),.BLN(BLN40),.WL(WL195));
sram_cell_6t_5 inst_cell_195_41 (.BL(BL41),.BLN(BLN41),.WL(WL195));
sram_cell_6t_5 inst_cell_195_42 (.BL(BL42),.BLN(BLN42),.WL(WL195));
sram_cell_6t_5 inst_cell_195_43 (.BL(BL43),.BLN(BLN43),.WL(WL195));
sram_cell_6t_5 inst_cell_195_44 (.BL(BL44),.BLN(BLN44),.WL(WL195));
sram_cell_6t_5 inst_cell_195_45 (.BL(BL45),.BLN(BLN45),.WL(WL195));
sram_cell_6t_5 inst_cell_195_46 (.BL(BL46),.BLN(BLN46),.WL(WL195));
sram_cell_6t_5 inst_cell_195_47 (.BL(BL47),.BLN(BLN47),.WL(WL195));
sram_cell_6t_5 inst_cell_195_48 (.BL(BL48),.BLN(BLN48),.WL(WL195));
sram_cell_6t_5 inst_cell_195_49 (.BL(BL49),.BLN(BLN49),.WL(WL195));
sram_cell_6t_5 inst_cell_195_50 (.BL(BL50),.BLN(BLN50),.WL(WL195));
sram_cell_6t_5 inst_cell_195_51 (.BL(BL51),.BLN(BLN51),.WL(WL195));
sram_cell_6t_5 inst_cell_195_52 (.BL(BL52),.BLN(BLN52),.WL(WL195));
sram_cell_6t_5 inst_cell_195_53 (.BL(BL53),.BLN(BLN53),.WL(WL195));
sram_cell_6t_5 inst_cell_195_54 (.BL(BL54),.BLN(BLN54),.WL(WL195));
sram_cell_6t_5 inst_cell_195_55 (.BL(BL55),.BLN(BLN55),.WL(WL195));
sram_cell_6t_5 inst_cell_195_56 (.BL(BL56),.BLN(BLN56),.WL(WL195));
sram_cell_6t_5 inst_cell_195_57 (.BL(BL57),.BLN(BLN57),.WL(WL195));
sram_cell_6t_5 inst_cell_195_58 (.BL(BL58),.BLN(BLN58),.WL(WL195));
sram_cell_6t_5 inst_cell_195_59 (.BL(BL59),.BLN(BLN59),.WL(WL195));
sram_cell_6t_5 inst_cell_195_60 (.BL(BL60),.BLN(BLN60),.WL(WL195));
sram_cell_6t_5 inst_cell_195_61 (.BL(BL61),.BLN(BLN61),.WL(WL195));
sram_cell_6t_5 inst_cell_195_62 (.BL(BL62),.BLN(BLN62),.WL(WL195));
sram_cell_6t_5 inst_cell_195_63 (.BL(BL63),.BLN(BLN63),.WL(WL195));
sram_cell_6t_5 inst_cell_195_64 (.BL(BL64),.BLN(BLN64),.WL(WL195));
sram_cell_6t_5 inst_cell_195_65 (.BL(BL65),.BLN(BLN65),.WL(WL195));
sram_cell_6t_5 inst_cell_195_66 (.BL(BL66),.BLN(BLN66),.WL(WL195));
sram_cell_6t_5 inst_cell_195_67 (.BL(BL67),.BLN(BLN67),.WL(WL195));
sram_cell_6t_5 inst_cell_195_68 (.BL(BL68),.BLN(BLN68),.WL(WL195));
sram_cell_6t_5 inst_cell_195_69 (.BL(BL69),.BLN(BLN69),.WL(WL195));
sram_cell_6t_5 inst_cell_195_70 (.BL(BL70),.BLN(BLN70),.WL(WL195));
sram_cell_6t_5 inst_cell_195_71 (.BL(BL71),.BLN(BLN71),.WL(WL195));
sram_cell_6t_5 inst_cell_195_72 (.BL(BL72),.BLN(BLN72),.WL(WL195));
sram_cell_6t_5 inst_cell_195_73 (.BL(BL73),.BLN(BLN73),.WL(WL195));
sram_cell_6t_5 inst_cell_195_74 (.BL(BL74),.BLN(BLN74),.WL(WL195));
sram_cell_6t_5 inst_cell_195_75 (.BL(BL75),.BLN(BLN75),.WL(WL195));
sram_cell_6t_5 inst_cell_195_76 (.BL(BL76),.BLN(BLN76),.WL(WL195));
sram_cell_6t_5 inst_cell_195_77 (.BL(BL77),.BLN(BLN77),.WL(WL195));
sram_cell_6t_5 inst_cell_195_78 (.BL(BL78),.BLN(BLN78),.WL(WL195));
sram_cell_6t_5 inst_cell_195_79 (.BL(BL79),.BLN(BLN79),.WL(WL195));
sram_cell_6t_5 inst_cell_195_80 (.BL(BL80),.BLN(BLN80),.WL(WL195));
sram_cell_6t_5 inst_cell_195_81 (.BL(BL81),.BLN(BLN81),.WL(WL195));
sram_cell_6t_5 inst_cell_195_82 (.BL(BL82),.BLN(BLN82),.WL(WL195));
sram_cell_6t_5 inst_cell_195_83 (.BL(BL83),.BLN(BLN83),.WL(WL195));
sram_cell_6t_5 inst_cell_195_84 (.BL(BL84),.BLN(BLN84),.WL(WL195));
sram_cell_6t_5 inst_cell_195_85 (.BL(BL85),.BLN(BLN85),.WL(WL195));
sram_cell_6t_5 inst_cell_195_86 (.BL(BL86),.BLN(BLN86),.WL(WL195));
sram_cell_6t_5 inst_cell_195_87 (.BL(BL87),.BLN(BLN87),.WL(WL195));
sram_cell_6t_5 inst_cell_195_88 (.BL(BL88),.BLN(BLN88),.WL(WL195));
sram_cell_6t_5 inst_cell_195_89 (.BL(BL89),.BLN(BLN89),.WL(WL195));
sram_cell_6t_5 inst_cell_195_90 (.BL(BL90),.BLN(BLN90),.WL(WL195));
sram_cell_6t_5 inst_cell_195_91 (.BL(BL91),.BLN(BLN91),.WL(WL195));
sram_cell_6t_5 inst_cell_195_92 (.BL(BL92),.BLN(BLN92),.WL(WL195));
sram_cell_6t_5 inst_cell_195_93 (.BL(BL93),.BLN(BLN93),.WL(WL195));
sram_cell_6t_5 inst_cell_195_94 (.BL(BL94),.BLN(BLN94),.WL(WL195));
sram_cell_6t_5 inst_cell_195_95 (.BL(BL95),.BLN(BLN95),.WL(WL195));
sram_cell_6t_5 inst_cell_195_96 (.BL(BL96),.BLN(BLN96),.WL(WL195));
sram_cell_6t_5 inst_cell_195_97 (.BL(BL97),.BLN(BLN97),.WL(WL195));
sram_cell_6t_5 inst_cell_195_98 (.BL(BL98),.BLN(BLN98),.WL(WL195));
sram_cell_6t_5 inst_cell_195_99 (.BL(BL99),.BLN(BLN99),.WL(WL195));
sram_cell_6t_5 inst_cell_195_100 (.BL(BL100),.BLN(BLN100),.WL(WL195));
sram_cell_6t_5 inst_cell_195_101 (.BL(BL101),.BLN(BLN101),.WL(WL195));
sram_cell_6t_5 inst_cell_195_102 (.BL(BL102),.BLN(BLN102),.WL(WL195));
sram_cell_6t_5 inst_cell_195_103 (.BL(BL103),.BLN(BLN103),.WL(WL195));
sram_cell_6t_5 inst_cell_195_104 (.BL(BL104),.BLN(BLN104),.WL(WL195));
sram_cell_6t_5 inst_cell_195_105 (.BL(BL105),.BLN(BLN105),.WL(WL195));
sram_cell_6t_5 inst_cell_195_106 (.BL(BL106),.BLN(BLN106),.WL(WL195));
sram_cell_6t_5 inst_cell_195_107 (.BL(BL107),.BLN(BLN107),.WL(WL195));
sram_cell_6t_5 inst_cell_195_108 (.BL(BL108),.BLN(BLN108),.WL(WL195));
sram_cell_6t_5 inst_cell_195_109 (.BL(BL109),.BLN(BLN109),.WL(WL195));
sram_cell_6t_5 inst_cell_195_110 (.BL(BL110),.BLN(BLN110),.WL(WL195));
sram_cell_6t_5 inst_cell_195_111 (.BL(BL111),.BLN(BLN111),.WL(WL195));
sram_cell_6t_5 inst_cell_195_112 (.BL(BL112),.BLN(BLN112),.WL(WL195));
sram_cell_6t_5 inst_cell_195_113 (.BL(BL113),.BLN(BLN113),.WL(WL195));
sram_cell_6t_5 inst_cell_195_114 (.BL(BL114),.BLN(BLN114),.WL(WL195));
sram_cell_6t_5 inst_cell_195_115 (.BL(BL115),.BLN(BLN115),.WL(WL195));
sram_cell_6t_5 inst_cell_195_116 (.BL(BL116),.BLN(BLN116),.WL(WL195));
sram_cell_6t_5 inst_cell_195_117 (.BL(BL117),.BLN(BLN117),.WL(WL195));
sram_cell_6t_5 inst_cell_195_118 (.BL(BL118),.BLN(BLN118),.WL(WL195));
sram_cell_6t_5 inst_cell_195_119 (.BL(BL119),.BLN(BLN119),.WL(WL195));
sram_cell_6t_5 inst_cell_195_120 (.BL(BL120),.BLN(BLN120),.WL(WL195));
sram_cell_6t_5 inst_cell_195_121 (.BL(BL121),.BLN(BLN121),.WL(WL195));
sram_cell_6t_5 inst_cell_195_122 (.BL(BL122),.BLN(BLN122),.WL(WL195));
sram_cell_6t_5 inst_cell_195_123 (.BL(BL123),.BLN(BLN123),.WL(WL195));
sram_cell_6t_5 inst_cell_195_124 (.BL(BL124),.BLN(BLN124),.WL(WL195));
sram_cell_6t_5 inst_cell_195_125 (.BL(BL125),.BLN(BLN125),.WL(WL195));
sram_cell_6t_5 inst_cell_195_126 (.BL(BL126),.BLN(BLN126),.WL(WL195));
sram_cell_6t_5 inst_cell_195_127 (.BL(BL127),.BLN(BLN127),.WL(WL195));
sram_cell_6t_5 inst_cell_196_0 (.BL(BL0),.BLN(BLN0),.WL(WL196));
sram_cell_6t_5 inst_cell_196_1 (.BL(BL1),.BLN(BLN1),.WL(WL196));
sram_cell_6t_5 inst_cell_196_2 (.BL(BL2),.BLN(BLN2),.WL(WL196));
sram_cell_6t_5 inst_cell_196_3 (.BL(BL3),.BLN(BLN3),.WL(WL196));
sram_cell_6t_5 inst_cell_196_4 (.BL(BL4),.BLN(BLN4),.WL(WL196));
sram_cell_6t_5 inst_cell_196_5 (.BL(BL5),.BLN(BLN5),.WL(WL196));
sram_cell_6t_5 inst_cell_196_6 (.BL(BL6),.BLN(BLN6),.WL(WL196));
sram_cell_6t_5 inst_cell_196_7 (.BL(BL7),.BLN(BLN7),.WL(WL196));
sram_cell_6t_5 inst_cell_196_8 (.BL(BL8),.BLN(BLN8),.WL(WL196));
sram_cell_6t_5 inst_cell_196_9 (.BL(BL9),.BLN(BLN9),.WL(WL196));
sram_cell_6t_5 inst_cell_196_10 (.BL(BL10),.BLN(BLN10),.WL(WL196));
sram_cell_6t_5 inst_cell_196_11 (.BL(BL11),.BLN(BLN11),.WL(WL196));
sram_cell_6t_5 inst_cell_196_12 (.BL(BL12),.BLN(BLN12),.WL(WL196));
sram_cell_6t_5 inst_cell_196_13 (.BL(BL13),.BLN(BLN13),.WL(WL196));
sram_cell_6t_5 inst_cell_196_14 (.BL(BL14),.BLN(BLN14),.WL(WL196));
sram_cell_6t_5 inst_cell_196_15 (.BL(BL15),.BLN(BLN15),.WL(WL196));
sram_cell_6t_5 inst_cell_196_16 (.BL(BL16),.BLN(BLN16),.WL(WL196));
sram_cell_6t_5 inst_cell_196_17 (.BL(BL17),.BLN(BLN17),.WL(WL196));
sram_cell_6t_5 inst_cell_196_18 (.BL(BL18),.BLN(BLN18),.WL(WL196));
sram_cell_6t_5 inst_cell_196_19 (.BL(BL19),.BLN(BLN19),.WL(WL196));
sram_cell_6t_5 inst_cell_196_20 (.BL(BL20),.BLN(BLN20),.WL(WL196));
sram_cell_6t_5 inst_cell_196_21 (.BL(BL21),.BLN(BLN21),.WL(WL196));
sram_cell_6t_5 inst_cell_196_22 (.BL(BL22),.BLN(BLN22),.WL(WL196));
sram_cell_6t_5 inst_cell_196_23 (.BL(BL23),.BLN(BLN23),.WL(WL196));
sram_cell_6t_5 inst_cell_196_24 (.BL(BL24),.BLN(BLN24),.WL(WL196));
sram_cell_6t_5 inst_cell_196_25 (.BL(BL25),.BLN(BLN25),.WL(WL196));
sram_cell_6t_5 inst_cell_196_26 (.BL(BL26),.BLN(BLN26),.WL(WL196));
sram_cell_6t_5 inst_cell_196_27 (.BL(BL27),.BLN(BLN27),.WL(WL196));
sram_cell_6t_5 inst_cell_196_28 (.BL(BL28),.BLN(BLN28),.WL(WL196));
sram_cell_6t_5 inst_cell_196_29 (.BL(BL29),.BLN(BLN29),.WL(WL196));
sram_cell_6t_5 inst_cell_196_30 (.BL(BL30),.BLN(BLN30),.WL(WL196));
sram_cell_6t_5 inst_cell_196_31 (.BL(BL31),.BLN(BLN31),.WL(WL196));
sram_cell_6t_5 inst_cell_196_32 (.BL(BL32),.BLN(BLN32),.WL(WL196));
sram_cell_6t_5 inst_cell_196_33 (.BL(BL33),.BLN(BLN33),.WL(WL196));
sram_cell_6t_5 inst_cell_196_34 (.BL(BL34),.BLN(BLN34),.WL(WL196));
sram_cell_6t_5 inst_cell_196_35 (.BL(BL35),.BLN(BLN35),.WL(WL196));
sram_cell_6t_5 inst_cell_196_36 (.BL(BL36),.BLN(BLN36),.WL(WL196));
sram_cell_6t_5 inst_cell_196_37 (.BL(BL37),.BLN(BLN37),.WL(WL196));
sram_cell_6t_5 inst_cell_196_38 (.BL(BL38),.BLN(BLN38),.WL(WL196));
sram_cell_6t_5 inst_cell_196_39 (.BL(BL39),.BLN(BLN39),.WL(WL196));
sram_cell_6t_5 inst_cell_196_40 (.BL(BL40),.BLN(BLN40),.WL(WL196));
sram_cell_6t_5 inst_cell_196_41 (.BL(BL41),.BLN(BLN41),.WL(WL196));
sram_cell_6t_5 inst_cell_196_42 (.BL(BL42),.BLN(BLN42),.WL(WL196));
sram_cell_6t_5 inst_cell_196_43 (.BL(BL43),.BLN(BLN43),.WL(WL196));
sram_cell_6t_5 inst_cell_196_44 (.BL(BL44),.BLN(BLN44),.WL(WL196));
sram_cell_6t_5 inst_cell_196_45 (.BL(BL45),.BLN(BLN45),.WL(WL196));
sram_cell_6t_5 inst_cell_196_46 (.BL(BL46),.BLN(BLN46),.WL(WL196));
sram_cell_6t_5 inst_cell_196_47 (.BL(BL47),.BLN(BLN47),.WL(WL196));
sram_cell_6t_5 inst_cell_196_48 (.BL(BL48),.BLN(BLN48),.WL(WL196));
sram_cell_6t_5 inst_cell_196_49 (.BL(BL49),.BLN(BLN49),.WL(WL196));
sram_cell_6t_5 inst_cell_196_50 (.BL(BL50),.BLN(BLN50),.WL(WL196));
sram_cell_6t_5 inst_cell_196_51 (.BL(BL51),.BLN(BLN51),.WL(WL196));
sram_cell_6t_5 inst_cell_196_52 (.BL(BL52),.BLN(BLN52),.WL(WL196));
sram_cell_6t_5 inst_cell_196_53 (.BL(BL53),.BLN(BLN53),.WL(WL196));
sram_cell_6t_5 inst_cell_196_54 (.BL(BL54),.BLN(BLN54),.WL(WL196));
sram_cell_6t_5 inst_cell_196_55 (.BL(BL55),.BLN(BLN55),.WL(WL196));
sram_cell_6t_5 inst_cell_196_56 (.BL(BL56),.BLN(BLN56),.WL(WL196));
sram_cell_6t_5 inst_cell_196_57 (.BL(BL57),.BLN(BLN57),.WL(WL196));
sram_cell_6t_5 inst_cell_196_58 (.BL(BL58),.BLN(BLN58),.WL(WL196));
sram_cell_6t_5 inst_cell_196_59 (.BL(BL59),.BLN(BLN59),.WL(WL196));
sram_cell_6t_5 inst_cell_196_60 (.BL(BL60),.BLN(BLN60),.WL(WL196));
sram_cell_6t_5 inst_cell_196_61 (.BL(BL61),.BLN(BLN61),.WL(WL196));
sram_cell_6t_5 inst_cell_196_62 (.BL(BL62),.BLN(BLN62),.WL(WL196));
sram_cell_6t_5 inst_cell_196_63 (.BL(BL63),.BLN(BLN63),.WL(WL196));
sram_cell_6t_5 inst_cell_196_64 (.BL(BL64),.BLN(BLN64),.WL(WL196));
sram_cell_6t_5 inst_cell_196_65 (.BL(BL65),.BLN(BLN65),.WL(WL196));
sram_cell_6t_5 inst_cell_196_66 (.BL(BL66),.BLN(BLN66),.WL(WL196));
sram_cell_6t_5 inst_cell_196_67 (.BL(BL67),.BLN(BLN67),.WL(WL196));
sram_cell_6t_5 inst_cell_196_68 (.BL(BL68),.BLN(BLN68),.WL(WL196));
sram_cell_6t_5 inst_cell_196_69 (.BL(BL69),.BLN(BLN69),.WL(WL196));
sram_cell_6t_5 inst_cell_196_70 (.BL(BL70),.BLN(BLN70),.WL(WL196));
sram_cell_6t_5 inst_cell_196_71 (.BL(BL71),.BLN(BLN71),.WL(WL196));
sram_cell_6t_5 inst_cell_196_72 (.BL(BL72),.BLN(BLN72),.WL(WL196));
sram_cell_6t_5 inst_cell_196_73 (.BL(BL73),.BLN(BLN73),.WL(WL196));
sram_cell_6t_5 inst_cell_196_74 (.BL(BL74),.BLN(BLN74),.WL(WL196));
sram_cell_6t_5 inst_cell_196_75 (.BL(BL75),.BLN(BLN75),.WL(WL196));
sram_cell_6t_5 inst_cell_196_76 (.BL(BL76),.BLN(BLN76),.WL(WL196));
sram_cell_6t_5 inst_cell_196_77 (.BL(BL77),.BLN(BLN77),.WL(WL196));
sram_cell_6t_5 inst_cell_196_78 (.BL(BL78),.BLN(BLN78),.WL(WL196));
sram_cell_6t_5 inst_cell_196_79 (.BL(BL79),.BLN(BLN79),.WL(WL196));
sram_cell_6t_5 inst_cell_196_80 (.BL(BL80),.BLN(BLN80),.WL(WL196));
sram_cell_6t_5 inst_cell_196_81 (.BL(BL81),.BLN(BLN81),.WL(WL196));
sram_cell_6t_5 inst_cell_196_82 (.BL(BL82),.BLN(BLN82),.WL(WL196));
sram_cell_6t_5 inst_cell_196_83 (.BL(BL83),.BLN(BLN83),.WL(WL196));
sram_cell_6t_5 inst_cell_196_84 (.BL(BL84),.BLN(BLN84),.WL(WL196));
sram_cell_6t_5 inst_cell_196_85 (.BL(BL85),.BLN(BLN85),.WL(WL196));
sram_cell_6t_5 inst_cell_196_86 (.BL(BL86),.BLN(BLN86),.WL(WL196));
sram_cell_6t_5 inst_cell_196_87 (.BL(BL87),.BLN(BLN87),.WL(WL196));
sram_cell_6t_5 inst_cell_196_88 (.BL(BL88),.BLN(BLN88),.WL(WL196));
sram_cell_6t_5 inst_cell_196_89 (.BL(BL89),.BLN(BLN89),.WL(WL196));
sram_cell_6t_5 inst_cell_196_90 (.BL(BL90),.BLN(BLN90),.WL(WL196));
sram_cell_6t_5 inst_cell_196_91 (.BL(BL91),.BLN(BLN91),.WL(WL196));
sram_cell_6t_5 inst_cell_196_92 (.BL(BL92),.BLN(BLN92),.WL(WL196));
sram_cell_6t_5 inst_cell_196_93 (.BL(BL93),.BLN(BLN93),.WL(WL196));
sram_cell_6t_5 inst_cell_196_94 (.BL(BL94),.BLN(BLN94),.WL(WL196));
sram_cell_6t_5 inst_cell_196_95 (.BL(BL95),.BLN(BLN95),.WL(WL196));
sram_cell_6t_5 inst_cell_196_96 (.BL(BL96),.BLN(BLN96),.WL(WL196));
sram_cell_6t_5 inst_cell_196_97 (.BL(BL97),.BLN(BLN97),.WL(WL196));
sram_cell_6t_5 inst_cell_196_98 (.BL(BL98),.BLN(BLN98),.WL(WL196));
sram_cell_6t_5 inst_cell_196_99 (.BL(BL99),.BLN(BLN99),.WL(WL196));
sram_cell_6t_5 inst_cell_196_100 (.BL(BL100),.BLN(BLN100),.WL(WL196));
sram_cell_6t_5 inst_cell_196_101 (.BL(BL101),.BLN(BLN101),.WL(WL196));
sram_cell_6t_5 inst_cell_196_102 (.BL(BL102),.BLN(BLN102),.WL(WL196));
sram_cell_6t_5 inst_cell_196_103 (.BL(BL103),.BLN(BLN103),.WL(WL196));
sram_cell_6t_5 inst_cell_196_104 (.BL(BL104),.BLN(BLN104),.WL(WL196));
sram_cell_6t_5 inst_cell_196_105 (.BL(BL105),.BLN(BLN105),.WL(WL196));
sram_cell_6t_5 inst_cell_196_106 (.BL(BL106),.BLN(BLN106),.WL(WL196));
sram_cell_6t_5 inst_cell_196_107 (.BL(BL107),.BLN(BLN107),.WL(WL196));
sram_cell_6t_5 inst_cell_196_108 (.BL(BL108),.BLN(BLN108),.WL(WL196));
sram_cell_6t_5 inst_cell_196_109 (.BL(BL109),.BLN(BLN109),.WL(WL196));
sram_cell_6t_5 inst_cell_196_110 (.BL(BL110),.BLN(BLN110),.WL(WL196));
sram_cell_6t_5 inst_cell_196_111 (.BL(BL111),.BLN(BLN111),.WL(WL196));
sram_cell_6t_5 inst_cell_196_112 (.BL(BL112),.BLN(BLN112),.WL(WL196));
sram_cell_6t_5 inst_cell_196_113 (.BL(BL113),.BLN(BLN113),.WL(WL196));
sram_cell_6t_5 inst_cell_196_114 (.BL(BL114),.BLN(BLN114),.WL(WL196));
sram_cell_6t_5 inst_cell_196_115 (.BL(BL115),.BLN(BLN115),.WL(WL196));
sram_cell_6t_5 inst_cell_196_116 (.BL(BL116),.BLN(BLN116),.WL(WL196));
sram_cell_6t_5 inst_cell_196_117 (.BL(BL117),.BLN(BLN117),.WL(WL196));
sram_cell_6t_5 inst_cell_196_118 (.BL(BL118),.BLN(BLN118),.WL(WL196));
sram_cell_6t_5 inst_cell_196_119 (.BL(BL119),.BLN(BLN119),.WL(WL196));
sram_cell_6t_5 inst_cell_196_120 (.BL(BL120),.BLN(BLN120),.WL(WL196));
sram_cell_6t_5 inst_cell_196_121 (.BL(BL121),.BLN(BLN121),.WL(WL196));
sram_cell_6t_5 inst_cell_196_122 (.BL(BL122),.BLN(BLN122),.WL(WL196));
sram_cell_6t_5 inst_cell_196_123 (.BL(BL123),.BLN(BLN123),.WL(WL196));
sram_cell_6t_5 inst_cell_196_124 (.BL(BL124),.BLN(BLN124),.WL(WL196));
sram_cell_6t_5 inst_cell_196_125 (.BL(BL125),.BLN(BLN125),.WL(WL196));
sram_cell_6t_5 inst_cell_196_126 (.BL(BL126),.BLN(BLN126),.WL(WL196));
sram_cell_6t_5 inst_cell_196_127 (.BL(BL127),.BLN(BLN127),.WL(WL196));
sram_cell_6t_5 inst_cell_197_0 (.BL(BL0),.BLN(BLN0),.WL(WL197));
sram_cell_6t_5 inst_cell_197_1 (.BL(BL1),.BLN(BLN1),.WL(WL197));
sram_cell_6t_5 inst_cell_197_2 (.BL(BL2),.BLN(BLN2),.WL(WL197));
sram_cell_6t_5 inst_cell_197_3 (.BL(BL3),.BLN(BLN3),.WL(WL197));
sram_cell_6t_5 inst_cell_197_4 (.BL(BL4),.BLN(BLN4),.WL(WL197));
sram_cell_6t_5 inst_cell_197_5 (.BL(BL5),.BLN(BLN5),.WL(WL197));
sram_cell_6t_5 inst_cell_197_6 (.BL(BL6),.BLN(BLN6),.WL(WL197));
sram_cell_6t_5 inst_cell_197_7 (.BL(BL7),.BLN(BLN7),.WL(WL197));
sram_cell_6t_5 inst_cell_197_8 (.BL(BL8),.BLN(BLN8),.WL(WL197));
sram_cell_6t_5 inst_cell_197_9 (.BL(BL9),.BLN(BLN9),.WL(WL197));
sram_cell_6t_5 inst_cell_197_10 (.BL(BL10),.BLN(BLN10),.WL(WL197));
sram_cell_6t_5 inst_cell_197_11 (.BL(BL11),.BLN(BLN11),.WL(WL197));
sram_cell_6t_5 inst_cell_197_12 (.BL(BL12),.BLN(BLN12),.WL(WL197));
sram_cell_6t_5 inst_cell_197_13 (.BL(BL13),.BLN(BLN13),.WL(WL197));
sram_cell_6t_5 inst_cell_197_14 (.BL(BL14),.BLN(BLN14),.WL(WL197));
sram_cell_6t_5 inst_cell_197_15 (.BL(BL15),.BLN(BLN15),.WL(WL197));
sram_cell_6t_5 inst_cell_197_16 (.BL(BL16),.BLN(BLN16),.WL(WL197));
sram_cell_6t_5 inst_cell_197_17 (.BL(BL17),.BLN(BLN17),.WL(WL197));
sram_cell_6t_5 inst_cell_197_18 (.BL(BL18),.BLN(BLN18),.WL(WL197));
sram_cell_6t_5 inst_cell_197_19 (.BL(BL19),.BLN(BLN19),.WL(WL197));
sram_cell_6t_5 inst_cell_197_20 (.BL(BL20),.BLN(BLN20),.WL(WL197));
sram_cell_6t_5 inst_cell_197_21 (.BL(BL21),.BLN(BLN21),.WL(WL197));
sram_cell_6t_5 inst_cell_197_22 (.BL(BL22),.BLN(BLN22),.WL(WL197));
sram_cell_6t_5 inst_cell_197_23 (.BL(BL23),.BLN(BLN23),.WL(WL197));
sram_cell_6t_5 inst_cell_197_24 (.BL(BL24),.BLN(BLN24),.WL(WL197));
sram_cell_6t_5 inst_cell_197_25 (.BL(BL25),.BLN(BLN25),.WL(WL197));
sram_cell_6t_5 inst_cell_197_26 (.BL(BL26),.BLN(BLN26),.WL(WL197));
sram_cell_6t_5 inst_cell_197_27 (.BL(BL27),.BLN(BLN27),.WL(WL197));
sram_cell_6t_5 inst_cell_197_28 (.BL(BL28),.BLN(BLN28),.WL(WL197));
sram_cell_6t_5 inst_cell_197_29 (.BL(BL29),.BLN(BLN29),.WL(WL197));
sram_cell_6t_5 inst_cell_197_30 (.BL(BL30),.BLN(BLN30),.WL(WL197));
sram_cell_6t_5 inst_cell_197_31 (.BL(BL31),.BLN(BLN31),.WL(WL197));
sram_cell_6t_5 inst_cell_197_32 (.BL(BL32),.BLN(BLN32),.WL(WL197));
sram_cell_6t_5 inst_cell_197_33 (.BL(BL33),.BLN(BLN33),.WL(WL197));
sram_cell_6t_5 inst_cell_197_34 (.BL(BL34),.BLN(BLN34),.WL(WL197));
sram_cell_6t_5 inst_cell_197_35 (.BL(BL35),.BLN(BLN35),.WL(WL197));
sram_cell_6t_5 inst_cell_197_36 (.BL(BL36),.BLN(BLN36),.WL(WL197));
sram_cell_6t_5 inst_cell_197_37 (.BL(BL37),.BLN(BLN37),.WL(WL197));
sram_cell_6t_5 inst_cell_197_38 (.BL(BL38),.BLN(BLN38),.WL(WL197));
sram_cell_6t_5 inst_cell_197_39 (.BL(BL39),.BLN(BLN39),.WL(WL197));
sram_cell_6t_5 inst_cell_197_40 (.BL(BL40),.BLN(BLN40),.WL(WL197));
sram_cell_6t_5 inst_cell_197_41 (.BL(BL41),.BLN(BLN41),.WL(WL197));
sram_cell_6t_5 inst_cell_197_42 (.BL(BL42),.BLN(BLN42),.WL(WL197));
sram_cell_6t_5 inst_cell_197_43 (.BL(BL43),.BLN(BLN43),.WL(WL197));
sram_cell_6t_5 inst_cell_197_44 (.BL(BL44),.BLN(BLN44),.WL(WL197));
sram_cell_6t_5 inst_cell_197_45 (.BL(BL45),.BLN(BLN45),.WL(WL197));
sram_cell_6t_5 inst_cell_197_46 (.BL(BL46),.BLN(BLN46),.WL(WL197));
sram_cell_6t_5 inst_cell_197_47 (.BL(BL47),.BLN(BLN47),.WL(WL197));
sram_cell_6t_5 inst_cell_197_48 (.BL(BL48),.BLN(BLN48),.WL(WL197));
sram_cell_6t_5 inst_cell_197_49 (.BL(BL49),.BLN(BLN49),.WL(WL197));
sram_cell_6t_5 inst_cell_197_50 (.BL(BL50),.BLN(BLN50),.WL(WL197));
sram_cell_6t_5 inst_cell_197_51 (.BL(BL51),.BLN(BLN51),.WL(WL197));
sram_cell_6t_5 inst_cell_197_52 (.BL(BL52),.BLN(BLN52),.WL(WL197));
sram_cell_6t_5 inst_cell_197_53 (.BL(BL53),.BLN(BLN53),.WL(WL197));
sram_cell_6t_5 inst_cell_197_54 (.BL(BL54),.BLN(BLN54),.WL(WL197));
sram_cell_6t_5 inst_cell_197_55 (.BL(BL55),.BLN(BLN55),.WL(WL197));
sram_cell_6t_5 inst_cell_197_56 (.BL(BL56),.BLN(BLN56),.WL(WL197));
sram_cell_6t_5 inst_cell_197_57 (.BL(BL57),.BLN(BLN57),.WL(WL197));
sram_cell_6t_5 inst_cell_197_58 (.BL(BL58),.BLN(BLN58),.WL(WL197));
sram_cell_6t_5 inst_cell_197_59 (.BL(BL59),.BLN(BLN59),.WL(WL197));
sram_cell_6t_5 inst_cell_197_60 (.BL(BL60),.BLN(BLN60),.WL(WL197));
sram_cell_6t_5 inst_cell_197_61 (.BL(BL61),.BLN(BLN61),.WL(WL197));
sram_cell_6t_5 inst_cell_197_62 (.BL(BL62),.BLN(BLN62),.WL(WL197));
sram_cell_6t_5 inst_cell_197_63 (.BL(BL63),.BLN(BLN63),.WL(WL197));
sram_cell_6t_5 inst_cell_197_64 (.BL(BL64),.BLN(BLN64),.WL(WL197));
sram_cell_6t_5 inst_cell_197_65 (.BL(BL65),.BLN(BLN65),.WL(WL197));
sram_cell_6t_5 inst_cell_197_66 (.BL(BL66),.BLN(BLN66),.WL(WL197));
sram_cell_6t_5 inst_cell_197_67 (.BL(BL67),.BLN(BLN67),.WL(WL197));
sram_cell_6t_5 inst_cell_197_68 (.BL(BL68),.BLN(BLN68),.WL(WL197));
sram_cell_6t_5 inst_cell_197_69 (.BL(BL69),.BLN(BLN69),.WL(WL197));
sram_cell_6t_5 inst_cell_197_70 (.BL(BL70),.BLN(BLN70),.WL(WL197));
sram_cell_6t_5 inst_cell_197_71 (.BL(BL71),.BLN(BLN71),.WL(WL197));
sram_cell_6t_5 inst_cell_197_72 (.BL(BL72),.BLN(BLN72),.WL(WL197));
sram_cell_6t_5 inst_cell_197_73 (.BL(BL73),.BLN(BLN73),.WL(WL197));
sram_cell_6t_5 inst_cell_197_74 (.BL(BL74),.BLN(BLN74),.WL(WL197));
sram_cell_6t_5 inst_cell_197_75 (.BL(BL75),.BLN(BLN75),.WL(WL197));
sram_cell_6t_5 inst_cell_197_76 (.BL(BL76),.BLN(BLN76),.WL(WL197));
sram_cell_6t_5 inst_cell_197_77 (.BL(BL77),.BLN(BLN77),.WL(WL197));
sram_cell_6t_5 inst_cell_197_78 (.BL(BL78),.BLN(BLN78),.WL(WL197));
sram_cell_6t_5 inst_cell_197_79 (.BL(BL79),.BLN(BLN79),.WL(WL197));
sram_cell_6t_5 inst_cell_197_80 (.BL(BL80),.BLN(BLN80),.WL(WL197));
sram_cell_6t_5 inst_cell_197_81 (.BL(BL81),.BLN(BLN81),.WL(WL197));
sram_cell_6t_5 inst_cell_197_82 (.BL(BL82),.BLN(BLN82),.WL(WL197));
sram_cell_6t_5 inst_cell_197_83 (.BL(BL83),.BLN(BLN83),.WL(WL197));
sram_cell_6t_5 inst_cell_197_84 (.BL(BL84),.BLN(BLN84),.WL(WL197));
sram_cell_6t_5 inst_cell_197_85 (.BL(BL85),.BLN(BLN85),.WL(WL197));
sram_cell_6t_5 inst_cell_197_86 (.BL(BL86),.BLN(BLN86),.WL(WL197));
sram_cell_6t_5 inst_cell_197_87 (.BL(BL87),.BLN(BLN87),.WL(WL197));
sram_cell_6t_5 inst_cell_197_88 (.BL(BL88),.BLN(BLN88),.WL(WL197));
sram_cell_6t_5 inst_cell_197_89 (.BL(BL89),.BLN(BLN89),.WL(WL197));
sram_cell_6t_5 inst_cell_197_90 (.BL(BL90),.BLN(BLN90),.WL(WL197));
sram_cell_6t_5 inst_cell_197_91 (.BL(BL91),.BLN(BLN91),.WL(WL197));
sram_cell_6t_5 inst_cell_197_92 (.BL(BL92),.BLN(BLN92),.WL(WL197));
sram_cell_6t_5 inst_cell_197_93 (.BL(BL93),.BLN(BLN93),.WL(WL197));
sram_cell_6t_5 inst_cell_197_94 (.BL(BL94),.BLN(BLN94),.WL(WL197));
sram_cell_6t_5 inst_cell_197_95 (.BL(BL95),.BLN(BLN95),.WL(WL197));
sram_cell_6t_5 inst_cell_197_96 (.BL(BL96),.BLN(BLN96),.WL(WL197));
sram_cell_6t_5 inst_cell_197_97 (.BL(BL97),.BLN(BLN97),.WL(WL197));
sram_cell_6t_5 inst_cell_197_98 (.BL(BL98),.BLN(BLN98),.WL(WL197));
sram_cell_6t_5 inst_cell_197_99 (.BL(BL99),.BLN(BLN99),.WL(WL197));
sram_cell_6t_5 inst_cell_197_100 (.BL(BL100),.BLN(BLN100),.WL(WL197));
sram_cell_6t_5 inst_cell_197_101 (.BL(BL101),.BLN(BLN101),.WL(WL197));
sram_cell_6t_5 inst_cell_197_102 (.BL(BL102),.BLN(BLN102),.WL(WL197));
sram_cell_6t_5 inst_cell_197_103 (.BL(BL103),.BLN(BLN103),.WL(WL197));
sram_cell_6t_5 inst_cell_197_104 (.BL(BL104),.BLN(BLN104),.WL(WL197));
sram_cell_6t_5 inst_cell_197_105 (.BL(BL105),.BLN(BLN105),.WL(WL197));
sram_cell_6t_5 inst_cell_197_106 (.BL(BL106),.BLN(BLN106),.WL(WL197));
sram_cell_6t_5 inst_cell_197_107 (.BL(BL107),.BLN(BLN107),.WL(WL197));
sram_cell_6t_5 inst_cell_197_108 (.BL(BL108),.BLN(BLN108),.WL(WL197));
sram_cell_6t_5 inst_cell_197_109 (.BL(BL109),.BLN(BLN109),.WL(WL197));
sram_cell_6t_5 inst_cell_197_110 (.BL(BL110),.BLN(BLN110),.WL(WL197));
sram_cell_6t_5 inst_cell_197_111 (.BL(BL111),.BLN(BLN111),.WL(WL197));
sram_cell_6t_5 inst_cell_197_112 (.BL(BL112),.BLN(BLN112),.WL(WL197));
sram_cell_6t_5 inst_cell_197_113 (.BL(BL113),.BLN(BLN113),.WL(WL197));
sram_cell_6t_5 inst_cell_197_114 (.BL(BL114),.BLN(BLN114),.WL(WL197));
sram_cell_6t_5 inst_cell_197_115 (.BL(BL115),.BLN(BLN115),.WL(WL197));
sram_cell_6t_5 inst_cell_197_116 (.BL(BL116),.BLN(BLN116),.WL(WL197));
sram_cell_6t_5 inst_cell_197_117 (.BL(BL117),.BLN(BLN117),.WL(WL197));
sram_cell_6t_5 inst_cell_197_118 (.BL(BL118),.BLN(BLN118),.WL(WL197));
sram_cell_6t_5 inst_cell_197_119 (.BL(BL119),.BLN(BLN119),.WL(WL197));
sram_cell_6t_5 inst_cell_197_120 (.BL(BL120),.BLN(BLN120),.WL(WL197));
sram_cell_6t_5 inst_cell_197_121 (.BL(BL121),.BLN(BLN121),.WL(WL197));
sram_cell_6t_5 inst_cell_197_122 (.BL(BL122),.BLN(BLN122),.WL(WL197));
sram_cell_6t_5 inst_cell_197_123 (.BL(BL123),.BLN(BLN123),.WL(WL197));
sram_cell_6t_5 inst_cell_197_124 (.BL(BL124),.BLN(BLN124),.WL(WL197));
sram_cell_6t_5 inst_cell_197_125 (.BL(BL125),.BLN(BLN125),.WL(WL197));
sram_cell_6t_5 inst_cell_197_126 (.BL(BL126),.BLN(BLN126),.WL(WL197));
sram_cell_6t_5 inst_cell_197_127 (.BL(BL127),.BLN(BLN127),.WL(WL197));
sram_cell_6t_5 inst_cell_198_0 (.BL(BL0),.BLN(BLN0),.WL(WL198));
sram_cell_6t_5 inst_cell_198_1 (.BL(BL1),.BLN(BLN1),.WL(WL198));
sram_cell_6t_5 inst_cell_198_2 (.BL(BL2),.BLN(BLN2),.WL(WL198));
sram_cell_6t_5 inst_cell_198_3 (.BL(BL3),.BLN(BLN3),.WL(WL198));
sram_cell_6t_5 inst_cell_198_4 (.BL(BL4),.BLN(BLN4),.WL(WL198));
sram_cell_6t_5 inst_cell_198_5 (.BL(BL5),.BLN(BLN5),.WL(WL198));
sram_cell_6t_5 inst_cell_198_6 (.BL(BL6),.BLN(BLN6),.WL(WL198));
sram_cell_6t_5 inst_cell_198_7 (.BL(BL7),.BLN(BLN7),.WL(WL198));
sram_cell_6t_5 inst_cell_198_8 (.BL(BL8),.BLN(BLN8),.WL(WL198));
sram_cell_6t_5 inst_cell_198_9 (.BL(BL9),.BLN(BLN9),.WL(WL198));
sram_cell_6t_5 inst_cell_198_10 (.BL(BL10),.BLN(BLN10),.WL(WL198));
sram_cell_6t_5 inst_cell_198_11 (.BL(BL11),.BLN(BLN11),.WL(WL198));
sram_cell_6t_5 inst_cell_198_12 (.BL(BL12),.BLN(BLN12),.WL(WL198));
sram_cell_6t_5 inst_cell_198_13 (.BL(BL13),.BLN(BLN13),.WL(WL198));
sram_cell_6t_5 inst_cell_198_14 (.BL(BL14),.BLN(BLN14),.WL(WL198));
sram_cell_6t_5 inst_cell_198_15 (.BL(BL15),.BLN(BLN15),.WL(WL198));
sram_cell_6t_5 inst_cell_198_16 (.BL(BL16),.BLN(BLN16),.WL(WL198));
sram_cell_6t_5 inst_cell_198_17 (.BL(BL17),.BLN(BLN17),.WL(WL198));
sram_cell_6t_5 inst_cell_198_18 (.BL(BL18),.BLN(BLN18),.WL(WL198));
sram_cell_6t_5 inst_cell_198_19 (.BL(BL19),.BLN(BLN19),.WL(WL198));
sram_cell_6t_5 inst_cell_198_20 (.BL(BL20),.BLN(BLN20),.WL(WL198));
sram_cell_6t_5 inst_cell_198_21 (.BL(BL21),.BLN(BLN21),.WL(WL198));
sram_cell_6t_5 inst_cell_198_22 (.BL(BL22),.BLN(BLN22),.WL(WL198));
sram_cell_6t_5 inst_cell_198_23 (.BL(BL23),.BLN(BLN23),.WL(WL198));
sram_cell_6t_5 inst_cell_198_24 (.BL(BL24),.BLN(BLN24),.WL(WL198));
sram_cell_6t_5 inst_cell_198_25 (.BL(BL25),.BLN(BLN25),.WL(WL198));
sram_cell_6t_5 inst_cell_198_26 (.BL(BL26),.BLN(BLN26),.WL(WL198));
sram_cell_6t_5 inst_cell_198_27 (.BL(BL27),.BLN(BLN27),.WL(WL198));
sram_cell_6t_5 inst_cell_198_28 (.BL(BL28),.BLN(BLN28),.WL(WL198));
sram_cell_6t_5 inst_cell_198_29 (.BL(BL29),.BLN(BLN29),.WL(WL198));
sram_cell_6t_5 inst_cell_198_30 (.BL(BL30),.BLN(BLN30),.WL(WL198));
sram_cell_6t_5 inst_cell_198_31 (.BL(BL31),.BLN(BLN31),.WL(WL198));
sram_cell_6t_5 inst_cell_198_32 (.BL(BL32),.BLN(BLN32),.WL(WL198));
sram_cell_6t_5 inst_cell_198_33 (.BL(BL33),.BLN(BLN33),.WL(WL198));
sram_cell_6t_5 inst_cell_198_34 (.BL(BL34),.BLN(BLN34),.WL(WL198));
sram_cell_6t_5 inst_cell_198_35 (.BL(BL35),.BLN(BLN35),.WL(WL198));
sram_cell_6t_5 inst_cell_198_36 (.BL(BL36),.BLN(BLN36),.WL(WL198));
sram_cell_6t_5 inst_cell_198_37 (.BL(BL37),.BLN(BLN37),.WL(WL198));
sram_cell_6t_5 inst_cell_198_38 (.BL(BL38),.BLN(BLN38),.WL(WL198));
sram_cell_6t_5 inst_cell_198_39 (.BL(BL39),.BLN(BLN39),.WL(WL198));
sram_cell_6t_5 inst_cell_198_40 (.BL(BL40),.BLN(BLN40),.WL(WL198));
sram_cell_6t_5 inst_cell_198_41 (.BL(BL41),.BLN(BLN41),.WL(WL198));
sram_cell_6t_5 inst_cell_198_42 (.BL(BL42),.BLN(BLN42),.WL(WL198));
sram_cell_6t_5 inst_cell_198_43 (.BL(BL43),.BLN(BLN43),.WL(WL198));
sram_cell_6t_5 inst_cell_198_44 (.BL(BL44),.BLN(BLN44),.WL(WL198));
sram_cell_6t_5 inst_cell_198_45 (.BL(BL45),.BLN(BLN45),.WL(WL198));
sram_cell_6t_5 inst_cell_198_46 (.BL(BL46),.BLN(BLN46),.WL(WL198));
sram_cell_6t_5 inst_cell_198_47 (.BL(BL47),.BLN(BLN47),.WL(WL198));
sram_cell_6t_5 inst_cell_198_48 (.BL(BL48),.BLN(BLN48),.WL(WL198));
sram_cell_6t_5 inst_cell_198_49 (.BL(BL49),.BLN(BLN49),.WL(WL198));
sram_cell_6t_5 inst_cell_198_50 (.BL(BL50),.BLN(BLN50),.WL(WL198));
sram_cell_6t_5 inst_cell_198_51 (.BL(BL51),.BLN(BLN51),.WL(WL198));
sram_cell_6t_5 inst_cell_198_52 (.BL(BL52),.BLN(BLN52),.WL(WL198));
sram_cell_6t_5 inst_cell_198_53 (.BL(BL53),.BLN(BLN53),.WL(WL198));
sram_cell_6t_5 inst_cell_198_54 (.BL(BL54),.BLN(BLN54),.WL(WL198));
sram_cell_6t_5 inst_cell_198_55 (.BL(BL55),.BLN(BLN55),.WL(WL198));
sram_cell_6t_5 inst_cell_198_56 (.BL(BL56),.BLN(BLN56),.WL(WL198));
sram_cell_6t_5 inst_cell_198_57 (.BL(BL57),.BLN(BLN57),.WL(WL198));
sram_cell_6t_5 inst_cell_198_58 (.BL(BL58),.BLN(BLN58),.WL(WL198));
sram_cell_6t_5 inst_cell_198_59 (.BL(BL59),.BLN(BLN59),.WL(WL198));
sram_cell_6t_5 inst_cell_198_60 (.BL(BL60),.BLN(BLN60),.WL(WL198));
sram_cell_6t_5 inst_cell_198_61 (.BL(BL61),.BLN(BLN61),.WL(WL198));
sram_cell_6t_5 inst_cell_198_62 (.BL(BL62),.BLN(BLN62),.WL(WL198));
sram_cell_6t_5 inst_cell_198_63 (.BL(BL63),.BLN(BLN63),.WL(WL198));
sram_cell_6t_5 inst_cell_198_64 (.BL(BL64),.BLN(BLN64),.WL(WL198));
sram_cell_6t_5 inst_cell_198_65 (.BL(BL65),.BLN(BLN65),.WL(WL198));
sram_cell_6t_5 inst_cell_198_66 (.BL(BL66),.BLN(BLN66),.WL(WL198));
sram_cell_6t_5 inst_cell_198_67 (.BL(BL67),.BLN(BLN67),.WL(WL198));
sram_cell_6t_5 inst_cell_198_68 (.BL(BL68),.BLN(BLN68),.WL(WL198));
sram_cell_6t_5 inst_cell_198_69 (.BL(BL69),.BLN(BLN69),.WL(WL198));
sram_cell_6t_5 inst_cell_198_70 (.BL(BL70),.BLN(BLN70),.WL(WL198));
sram_cell_6t_5 inst_cell_198_71 (.BL(BL71),.BLN(BLN71),.WL(WL198));
sram_cell_6t_5 inst_cell_198_72 (.BL(BL72),.BLN(BLN72),.WL(WL198));
sram_cell_6t_5 inst_cell_198_73 (.BL(BL73),.BLN(BLN73),.WL(WL198));
sram_cell_6t_5 inst_cell_198_74 (.BL(BL74),.BLN(BLN74),.WL(WL198));
sram_cell_6t_5 inst_cell_198_75 (.BL(BL75),.BLN(BLN75),.WL(WL198));
sram_cell_6t_5 inst_cell_198_76 (.BL(BL76),.BLN(BLN76),.WL(WL198));
sram_cell_6t_5 inst_cell_198_77 (.BL(BL77),.BLN(BLN77),.WL(WL198));
sram_cell_6t_5 inst_cell_198_78 (.BL(BL78),.BLN(BLN78),.WL(WL198));
sram_cell_6t_5 inst_cell_198_79 (.BL(BL79),.BLN(BLN79),.WL(WL198));
sram_cell_6t_5 inst_cell_198_80 (.BL(BL80),.BLN(BLN80),.WL(WL198));
sram_cell_6t_5 inst_cell_198_81 (.BL(BL81),.BLN(BLN81),.WL(WL198));
sram_cell_6t_5 inst_cell_198_82 (.BL(BL82),.BLN(BLN82),.WL(WL198));
sram_cell_6t_5 inst_cell_198_83 (.BL(BL83),.BLN(BLN83),.WL(WL198));
sram_cell_6t_5 inst_cell_198_84 (.BL(BL84),.BLN(BLN84),.WL(WL198));
sram_cell_6t_5 inst_cell_198_85 (.BL(BL85),.BLN(BLN85),.WL(WL198));
sram_cell_6t_5 inst_cell_198_86 (.BL(BL86),.BLN(BLN86),.WL(WL198));
sram_cell_6t_5 inst_cell_198_87 (.BL(BL87),.BLN(BLN87),.WL(WL198));
sram_cell_6t_5 inst_cell_198_88 (.BL(BL88),.BLN(BLN88),.WL(WL198));
sram_cell_6t_5 inst_cell_198_89 (.BL(BL89),.BLN(BLN89),.WL(WL198));
sram_cell_6t_5 inst_cell_198_90 (.BL(BL90),.BLN(BLN90),.WL(WL198));
sram_cell_6t_5 inst_cell_198_91 (.BL(BL91),.BLN(BLN91),.WL(WL198));
sram_cell_6t_5 inst_cell_198_92 (.BL(BL92),.BLN(BLN92),.WL(WL198));
sram_cell_6t_5 inst_cell_198_93 (.BL(BL93),.BLN(BLN93),.WL(WL198));
sram_cell_6t_5 inst_cell_198_94 (.BL(BL94),.BLN(BLN94),.WL(WL198));
sram_cell_6t_5 inst_cell_198_95 (.BL(BL95),.BLN(BLN95),.WL(WL198));
sram_cell_6t_5 inst_cell_198_96 (.BL(BL96),.BLN(BLN96),.WL(WL198));
sram_cell_6t_5 inst_cell_198_97 (.BL(BL97),.BLN(BLN97),.WL(WL198));
sram_cell_6t_5 inst_cell_198_98 (.BL(BL98),.BLN(BLN98),.WL(WL198));
sram_cell_6t_5 inst_cell_198_99 (.BL(BL99),.BLN(BLN99),.WL(WL198));
sram_cell_6t_5 inst_cell_198_100 (.BL(BL100),.BLN(BLN100),.WL(WL198));
sram_cell_6t_5 inst_cell_198_101 (.BL(BL101),.BLN(BLN101),.WL(WL198));
sram_cell_6t_5 inst_cell_198_102 (.BL(BL102),.BLN(BLN102),.WL(WL198));
sram_cell_6t_5 inst_cell_198_103 (.BL(BL103),.BLN(BLN103),.WL(WL198));
sram_cell_6t_5 inst_cell_198_104 (.BL(BL104),.BLN(BLN104),.WL(WL198));
sram_cell_6t_5 inst_cell_198_105 (.BL(BL105),.BLN(BLN105),.WL(WL198));
sram_cell_6t_5 inst_cell_198_106 (.BL(BL106),.BLN(BLN106),.WL(WL198));
sram_cell_6t_5 inst_cell_198_107 (.BL(BL107),.BLN(BLN107),.WL(WL198));
sram_cell_6t_5 inst_cell_198_108 (.BL(BL108),.BLN(BLN108),.WL(WL198));
sram_cell_6t_5 inst_cell_198_109 (.BL(BL109),.BLN(BLN109),.WL(WL198));
sram_cell_6t_5 inst_cell_198_110 (.BL(BL110),.BLN(BLN110),.WL(WL198));
sram_cell_6t_5 inst_cell_198_111 (.BL(BL111),.BLN(BLN111),.WL(WL198));
sram_cell_6t_5 inst_cell_198_112 (.BL(BL112),.BLN(BLN112),.WL(WL198));
sram_cell_6t_5 inst_cell_198_113 (.BL(BL113),.BLN(BLN113),.WL(WL198));
sram_cell_6t_5 inst_cell_198_114 (.BL(BL114),.BLN(BLN114),.WL(WL198));
sram_cell_6t_5 inst_cell_198_115 (.BL(BL115),.BLN(BLN115),.WL(WL198));
sram_cell_6t_5 inst_cell_198_116 (.BL(BL116),.BLN(BLN116),.WL(WL198));
sram_cell_6t_5 inst_cell_198_117 (.BL(BL117),.BLN(BLN117),.WL(WL198));
sram_cell_6t_5 inst_cell_198_118 (.BL(BL118),.BLN(BLN118),.WL(WL198));
sram_cell_6t_5 inst_cell_198_119 (.BL(BL119),.BLN(BLN119),.WL(WL198));
sram_cell_6t_5 inst_cell_198_120 (.BL(BL120),.BLN(BLN120),.WL(WL198));
sram_cell_6t_5 inst_cell_198_121 (.BL(BL121),.BLN(BLN121),.WL(WL198));
sram_cell_6t_5 inst_cell_198_122 (.BL(BL122),.BLN(BLN122),.WL(WL198));
sram_cell_6t_5 inst_cell_198_123 (.BL(BL123),.BLN(BLN123),.WL(WL198));
sram_cell_6t_5 inst_cell_198_124 (.BL(BL124),.BLN(BLN124),.WL(WL198));
sram_cell_6t_5 inst_cell_198_125 (.BL(BL125),.BLN(BLN125),.WL(WL198));
sram_cell_6t_5 inst_cell_198_126 (.BL(BL126),.BLN(BLN126),.WL(WL198));
sram_cell_6t_5 inst_cell_198_127 (.BL(BL127),.BLN(BLN127),.WL(WL198));
sram_cell_6t_5 inst_cell_199_0 (.BL(BL0),.BLN(BLN0),.WL(WL199));
sram_cell_6t_5 inst_cell_199_1 (.BL(BL1),.BLN(BLN1),.WL(WL199));
sram_cell_6t_5 inst_cell_199_2 (.BL(BL2),.BLN(BLN2),.WL(WL199));
sram_cell_6t_5 inst_cell_199_3 (.BL(BL3),.BLN(BLN3),.WL(WL199));
sram_cell_6t_5 inst_cell_199_4 (.BL(BL4),.BLN(BLN4),.WL(WL199));
sram_cell_6t_5 inst_cell_199_5 (.BL(BL5),.BLN(BLN5),.WL(WL199));
sram_cell_6t_5 inst_cell_199_6 (.BL(BL6),.BLN(BLN6),.WL(WL199));
sram_cell_6t_5 inst_cell_199_7 (.BL(BL7),.BLN(BLN7),.WL(WL199));
sram_cell_6t_5 inst_cell_199_8 (.BL(BL8),.BLN(BLN8),.WL(WL199));
sram_cell_6t_5 inst_cell_199_9 (.BL(BL9),.BLN(BLN9),.WL(WL199));
sram_cell_6t_5 inst_cell_199_10 (.BL(BL10),.BLN(BLN10),.WL(WL199));
sram_cell_6t_5 inst_cell_199_11 (.BL(BL11),.BLN(BLN11),.WL(WL199));
sram_cell_6t_5 inst_cell_199_12 (.BL(BL12),.BLN(BLN12),.WL(WL199));
sram_cell_6t_5 inst_cell_199_13 (.BL(BL13),.BLN(BLN13),.WL(WL199));
sram_cell_6t_5 inst_cell_199_14 (.BL(BL14),.BLN(BLN14),.WL(WL199));
sram_cell_6t_5 inst_cell_199_15 (.BL(BL15),.BLN(BLN15),.WL(WL199));
sram_cell_6t_5 inst_cell_199_16 (.BL(BL16),.BLN(BLN16),.WL(WL199));
sram_cell_6t_5 inst_cell_199_17 (.BL(BL17),.BLN(BLN17),.WL(WL199));
sram_cell_6t_5 inst_cell_199_18 (.BL(BL18),.BLN(BLN18),.WL(WL199));
sram_cell_6t_5 inst_cell_199_19 (.BL(BL19),.BLN(BLN19),.WL(WL199));
sram_cell_6t_5 inst_cell_199_20 (.BL(BL20),.BLN(BLN20),.WL(WL199));
sram_cell_6t_5 inst_cell_199_21 (.BL(BL21),.BLN(BLN21),.WL(WL199));
sram_cell_6t_5 inst_cell_199_22 (.BL(BL22),.BLN(BLN22),.WL(WL199));
sram_cell_6t_5 inst_cell_199_23 (.BL(BL23),.BLN(BLN23),.WL(WL199));
sram_cell_6t_5 inst_cell_199_24 (.BL(BL24),.BLN(BLN24),.WL(WL199));
sram_cell_6t_5 inst_cell_199_25 (.BL(BL25),.BLN(BLN25),.WL(WL199));
sram_cell_6t_5 inst_cell_199_26 (.BL(BL26),.BLN(BLN26),.WL(WL199));
sram_cell_6t_5 inst_cell_199_27 (.BL(BL27),.BLN(BLN27),.WL(WL199));
sram_cell_6t_5 inst_cell_199_28 (.BL(BL28),.BLN(BLN28),.WL(WL199));
sram_cell_6t_5 inst_cell_199_29 (.BL(BL29),.BLN(BLN29),.WL(WL199));
sram_cell_6t_5 inst_cell_199_30 (.BL(BL30),.BLN(BLN30),.WL(WL199));
sram_cell_6t_5 inst_cell_199_31 (.BL(BL31),.BLN(BLN31),.WL(WL199));
sram_cell_6t_5 inst_cell_199_32 (.BL(BL32),.BLN(BLN32),.WL(WL199));
sram_cell_6t_5 inst_cell_199_33 (.BL(BL33),.BLN(BLN33),.WL(WL199));
sram_cell_6t_5 inst_cell_199_34 (.BL(BL34),.BLN(BLN34),.WL(WL199));
sram_cell_6t_5 inst_cell_199_35 (.BL(BL35),.BLN(BLN35),.WL(WL199));
sram_cell_6t_5 inst_cell_199_36 (.BL(BL36),.BLN(BLN36),.WL(WL199));
sram_cell_6t_5 inst_cell_199_37 (.BL(BL37),.BLN(BLN37),.WL(WL199));
sram_cell_6t_5 inst_cell_199_38 (.BL(BL38),.BLN(BLN38),.WL(WL199));
sram_cell_6t_5 inst_cell_199_39 (.BL(BL39),.BLN(BLN39),.WL(WL199));
sram_cell_6t_5 inst_cell_199_40 (.BL(BL40),.BLN(BLN40),.WL(WL199));
sram_cell_6t_5 inst_cell_199_41 (.BL(BL41),.BLN(BLN41),.WL(WL199));
sram_cell_6t_5 inst_cell_199_42 (.BL(BL42),.BLN(BLN42),.WL(WL199));
sram_cell_6t_5 inst_cell_199_43 (.BL(BL43),.BLN(BLN43),.WL(WL199));
sram_cell_6t_5 inst_cell_199_44 (.BL(BL44),.BLN(BLN44),.WL(WL199));
sram_cell_6t_5 inst_cell_199_45 (.BL(BL45),.BLN(BLN45),.WL(WL199));
sram_cell_6t_5 inst_cell_199_46 (.BL(BL46),.BLN(BLN46),.WL(WL199));
sram_cell_6t_5 inst_cell_199_47 (.BL(BL47),.BLN(BLN47),.WL(WL199));
sram_cell_6t_5 inst_cell_199_48 (.BL(BL48),.BLN(BLN48),.WL(WL199));
sram_cell_6t_5 inst_cell_199_49 (.BL(BL49),.BLN(BLN49),.WL(WL199));
sram_cell_6t_5 inst_cell_199_50 (.BL(BL50),.BLN(BLN50),.WL(WL199));
sram_cell_6t_5 inst_cell_199_51 (.BL(BL51),.BLN(BLN51),.WL(WL199));
sram_cell_6t_5 inst_cell_199_52 (.BL(BL52),.BLN(BLN52),.WL(WL199));
sram_cell_6t_5 inst_cell_199_53 (.BL(BL53),.BLN(BLN53),.WL(WL199));
sram_cell_6t_5 inst_cell_199_54 (.BL(BL54),.BLN(BLN54),.WL(WL199));
sram_cell_6t_5 inst_cell_199_55 (.BL(BL55),.BLN(BLN55),.WL(WL199));
sram_cell_6t_5 inst_cell_199_56 (.BL(BL56),.BLN(BLN56),.WL(WL199));
sram_cell_6t_5 inst_cell_199_57 (.BL(BL57),.BLN(BLN57),.WL(WL199));
sram_cell_6t_5 inst_cell_199_58 (.BL(BL58),.BLN(BLN58),.WL(WL199));
sram_cell_6t_5 inst_cell_199_59 (.BL(BL59),.BLN(BLN59),.WL(WL199));
sram_cell_6t_5 inst_cell_199_60 (.BL(BL60),.BLN(BLN60),.WL(WL199));
sram_cell_6t_5 inst_cell_199_61 (.BL(BL61),.BLN(BLN61),.WL(WL199));
sram_cell_6t_5 inst_cell_199_62 (.BL(BL62),.BLN(BLN62),.WL(WL199));
sram_cell_6t_5 inst_cell_199_63 (.BL(BL63),.BLN(BLN63),.WL(WL199));
sram_cell_6t_5 inst_cell_199_64 (.BL(BL64),.BLN(BLN64),.WL(WL199));
sram_cell_6t_5 inst_cell_199_65 (.BL(BL65),.BLN(BLN65),.WL(WL199));
sram_cell_6t_5 inst_cell_199_66 (.BL(BL66),.BLN(BLN66),.WL(WL199));
sram_cell_6t_5 inst_cell_199_67 (.BL(BL67),.BLN(BLN67),.WL(WL199));
sram_cell_6t_5 inst_cell_199_68 (.BL(BL68),.BLN(BLN68),.WL(WL199));
sram_cell_6t_5 inst_cell_199_69 (.BL(BL69),.BLN(BLN69),.WL(WL199));
sram_cell_6t_5 inst_cell_199_70 (.BL(BL70),.BLN(BLN70),.WL(WL199));
sram_cell_6t_5 inst_cell_199_71 (.BL(BL71),.BLN(BLN71),.WL(WL199));
sram_cell_6t_5 inst_cell_199_72 (.BL(BL72),.BLN(BLN72),.WL(WL199));
sram_cell_6t_5 inst_cell_199_73 (.BL(BL73),.BLN(BLN73),.WL(WL199));
sram_cell_6t_5 inst_cell_199_74 (.BL(BL74),.BLN(BLN74),.WL(WL199));
sram_cell_6t_5 inst_cell_199_75 (.BL(BL75),.BLN(BLN75),.WL(WL199));
sram_cell_6t_5 inst_cell_199_76 (.BL(BL76),.BLN(BLN76),.WL(WL199));
sram_cell_6t_5 inst_cell_199_77 (.BL(BL77),.BLN(BLN77),.WL(WL199));
sram_cell_6t_5 inst_cell_199_78 (.BL(BL78),.BLN(BLN78),.WL(WL199));
sram_cell_6t_5 inst_cell_199_79 (.BL(BL79),.BLN(BLN79),.WL(WL199));
sram_cell_6t_5 inst_cell_199_80 (.BL(BL80),.BLN(BLN80),.WL(WL199));
sram_cell_6t_5 inst_cell_199_81 (.BL(BL81),.BLN(BLN81),.WL(WL199));
sram_cell_6t_5 inst_cell_199_82 (.BL(BL82),.BLN(BLN82),.WL(WL199));
sram_cell_6t_5 inst_cell_199_83 (.BL(BL83),.BLN(BLN83),.WL(WL199));
sram_cell_6t_5 inst_cell_199_84 (.BL(BL84),.BLN(BLN84),.WL(WL199));
sram_cell_6t_5 inst_cell_199_85 (.BL(BL85),.BLN(BLN85),.WL(WL199));
sram_cell_6t_5 inst_cell_199_86 (.BL(BL86),.BLN(BLN86),.WL(WL199));
sram_cell_6t_5 inst_cell_199_87 (.BL(BL87),.BLN(BLN87),.WL(WL199));
sram_cell_6t_5 inst_cell_199_88 (.BL(BL88),.BLN(BLN88),.WL(WL199));
sram_cell_6t_5 inst_cell_199_89 (.BL(BL89),.BLN(BLN89),.WL(WL199));
sram_cell_6t_5 inst_cell_199_90 (.BL(BL90),.BLN(BLN90),.WL(WL199));
sram_cell_6t_5 inst_cell_199_91 (.BL(BL91),.BLN(BLN91),.WL(WL199));
sram_cell_6t_5 inst_cell_199_92 (.BL(BL92),.BLN(BLN92),.WL(WL199));
sram_cell_6t_5 inst_cell_199_93 (.BL(BL93),.BLN(BLN93),.WL(WL199));
sram_cell_6t_5 inst_cell_199_94 (.BL(BL94),.BLN(BLN94),.WL(WL199));
sram_cell_6t_5 inst_cell_199_95 (.BL(BL95),.BLN(BLN95),.WL(WL199));
sram_cell_6t_5 inst_cell_199_96 (.BL(BL96),.BLN(BLN96),.WL(WL199));
sram_cell_6t_5 inst_cell_199_97 (.BL(BL97),.BLN(BLN97),.WL(WL199));
sram_cell_6t_5 inst_cell_199_98 (.BL(BL98),.BLN(BLN98),.WL(WL199));
sram_cell_6t_5 inst_cell_199_99 (.BL(BL99),.BLN(BLN99),.WL(WL199));
sram_cell_6t_5 inst_cell_199_100 (.BL(BL100),.BLN(BLN100),.WL(WL199));
sram_cell_6t_5 inst_cell_199_101 (.BL(BL101),.BLN(BLN101),.WL(WL199));
sram_cell_6t_5 inst_cell_199_102 (.BL(BL102),.BLN(BLN102),.WL(WL199));
sram_cell_6t_5 inst_cell_199_103 (.BL(BL103),.BLN(BLN103),.WL(WL199));
sram_cell_6t_5 inst_cell_199_104 (.BL(BL104),.BLN(BLN104),.WL(WL199));
sram_cell_6t_5 inst_cell_199_105 (.BL(BL105),.BLN(BLN105),.WL(WL199));
sram_cell_6t_5 inst_cell_199_106 (.BL(BL106),.BLN(BLN106),.WL(WL199));
sram_cell_6t_5 inst_cell_199_107 (.BL(BL107),.BLN(BLN107),.WL(WL199));
sram_cell_6t_5 inst_cell_199_108 (.BL(BL108),.BLN(BLN108),.WL(WL199));
sram_cell_6t_5 inst_cell_199_109 (.BL(BL109),.BLN(BLN109),.WL(WL199));
sram_cell_6t_5 inst_cell_199_110 (.BL(BL110),.BLN(BLN110),.WL(WL199));
sram_cell_6t_5 inst_cell_199_111 (.BL(BL111),.BLN(BLN111),.WL(WL199));
sram_cell_6t_5 inst_cell_199_112 (.BL(BL112),.BLN(BLN112),.WL(WL199));
sram_cell_6t_5 inst_cell_199_113 (.BL(BL113),.BLN(BLN113),.WL(WL199));
sram_cell_6t_5 inst_cell_199_114 (.BL(BL114),.BLN(BLN114),.WL(WL199));
sram_cell_6t_5 inst_cell_199_115 (.BL(BL115),.BLN(BLN115),.WL(WL199));
sram_cell_6t_5 inst_cell_199_116 (.BL(BL116),.BLN(BLN116),.WL(WL199));
sram_cell_6t_5 inst_cell_199_117 (.BL(BL117),.BLN(BLN117),.WL(WL199));
sram_cell_6t_5 inst_cell_199_118 (.BL(BL118),.BLN(BLN118),.WL(WL199));
sram_cell_6t_5 inst_cell_199_119 (.BL(BL119),.BLN(BLN119),.WL(WL199));
sram_cell_6t_5 inst_cell_199_120 (.BL(BL120),.BLN(BLN120),.WL(WL199));
sram_cell_6t_5 inst_cell_199_121 (.BL(BL121),.BLN(BLN121),.WL(WL199));
sram_cell_6t_5 inst_cell_199_122 (.BL(BL122),.BLN(BLN122),.WL(WL199));
sram_cell_6t_5 inst_cell_199_123 (.BL(BL123),.BLN(BLN123),.WL(WL199));
sram_cell_6t_5 inst_cell_199_124 (.BL(BL124),.BLN(BLN124),.WL(WL199));
sram_cell_6t_5 inst_cell_199_125 (.BL(BL125),.BLN(BLN125),.WL(WL199));
sram_cell_6t_5 inst_cell_199_126 (.BL(BL126),.BLN(BLN126),.WL(WL199));
sram_cell_6t_5 inst_cell_199_127 (.BL(BL127),.BLN(BLN127),.WL(WL199));
sram_cell_6t_5 inst_cell_200_0 (.BL(BL0),.BLN(BLN0),.WL(WL200));
sram_cell_6t_5 inst_cell_200_1 (.BL(BL1),.BLN(BLN1),.WL(WL200));
sram_cell_6t_5 inst_cell_200_2 (.BL(BL2),.BLN(BLN2),.WL(WL200));
sram_cell_6t_5 inst_cell_200_3 (.BL(BL3),.BLN(BLN3),.WL(WL200));
sram_cell_6t_5 inst_cell_200_4 (.BL(BL4),.BLN(BLN4),.WL(WL200));
sram_cell_6t_5 inst_cell_200_5 (.BL(BL5),.BLN(BLN5),.WL(WL200));
sram_cell_6t_5 inst_cell_200_6 (.BL(BL6),.BLN(BLN6),.WL(WL200));
sram_cell_6t_5 inst_cell_200_7 (.BL(BL7),.BLN(BLN7),.WL(WL200));
sram_cell_6t_5 inst_cell_200_8 (.BL(BL8),.BLN(BLN8),.WL(WL200));
sram_cell_6t_5 inst_cell_200_9 (.BL(BL9),.BLN(BLN9),.WL(WL200));
sram_cell_6t_5 inst_cell_200_10 (.BL(BL10),.BLN(BLN10),.WL(WL200));
sram_cell_6t_5 inst_cell_200_11 (.BL(BL11),.BLN(BLN11),.WL(WL200));
sram_cell_6t_5 inst_cell_200_12 (.BL(BL12),.BLN(BLN12),.WL(WL200));
sram_cell_6t_5 inst_cell_200_13 (.BL(BL13),.BLN(BLN13),.WL(WL200));
sram_cell_6t_5 inst_cell_200_14 (.BL(BL14),.BLN(BLN14),.WL(WL200));
sram_cell_6t_5 inst_cell_200_15 (.BL(BL15),.BLN(BLN15),.WL(WL200));
sram_cell_6t_5 inst_cell_200_16 (.BL(BL16),.BLN(BLN16),.WL(WL200));
sram_cell_6t_5 inst_cell_200_17 (.BL(BL17),.BLN(BLN17),.WL(WL200));
sram_cell_6t_5 inst_cell_200_18 (.BL(BL18),.BLN(BLN18),.WL(WL200));
sram_cell_6t_5 inst_cell_200_19 (.BL(BL19),.BLN(BLN19),.WL(WL200));
sram_cell_6t_5 inst_cell_200_20 (.BL(BL20),.BLN(BLN20),.WL(WL200));
sram_cell_6t_5 inst_cell_200_21 (.BL(BL21),.BLN(BLN21),.WL(WL200));
sram_cell_6t_5 inst_cell_200_22 (.BL(BL22),.BLN(BLN22),.WL(WL200));
sram_cell_6t_5 inst_cell_200_23 (.BL(BL23),.BLN(BLN23),.WL(WL200));
sram_cell_6t_5 inst_cell_200_24 (.BL(BL24),.BLN(BLN24),.WL(WL200));
sram_cell_6t_5 inst_cell_200_25 (.BL(BL25),.BLN(BLN25),.WL(WL200));
sram_cell_6t_5 inst_cell_200_26 (.BL(BL26),.BLN(BLN26),.WL(WL200));
sram_cell_6t_5 inst_cell_200_27 (.BL(BL27),.BLN(BLN27),.WL(WL200));
sram_cell_6t_5 inst_cell_200_28 (.BL(BL28),.BLN(BLN28),.WL(WL200));
sram_cell_6t_5 inst_cell_200_29 (.BL(BL29),.BLN(BLN29),.WL(WL200));
sram_cell_6t_5 inst_cell_200_30 (.BL(BL30),.BLN(BLN30),.WL(WL200));
sram_cell_6t_5 inst_cell_200_31 (.BL(BL31),.BLN(BLN31),.WL(WL200));
sram_cell_6t_5 inst_cell_200_32 (.BL(BL32),.BLN(BLN32),.WL(WL200));
sram_cell_6t_5 inst_cell_200_33 (.BL(BL33),.BLN(BLN33),.WL(WL200));
sram_cell_6t_5 inst_cell_200_34 (.BL(BL34),.BLN(BLN34),.WL(WL200));
sram_cell_6t_5 inst_cell_200_35 (.BL(BL35),.BLN(BLN35),.WL(WL200));
sram_cell_6t_5 inst_cell_200_36 (.BL(BL36),.BLN(BLN36),.WL(WL200));
sram_cell_6t_5 inst_cell_200_37 (.BL(BL37),.BLN(BLN37),.WL(WL200));
sram_cell_6t_5 inst_cell_200_38 (.BL(BL38),.BLN(BLN38),.WL(WL200));
sram_cell_6t_5 inst_cell_200_39 (.BL(BL39),.BLN(BLN39),.WL(WL200));
sram_cell_6t_5 inst_cell_200_40 (.BL(BL40),.BLN(BLN40),.WL(WL200));
sram_cell_6t_5 inst_cell_200_41 (.BL(BL41),.BLN(BLN41),.WL(WL200));
sram_cell_6t_5 inst_cell_200_42 (.BL(BL42),.BLN(BLN42),.WL(WL200));
sram_cell_6t_5 inst_cell_200_43 (.BL(BL43),.BLN(BLN43),.WL(WL200));
sram_cell_6t_5 inst_cell_200_44 (.BL(BL44),.BLN(BLN44),.WL(WL200));
sram_cell_6t_5 inst_cell_200_45 (.BL(BL45),.BLN(BLN45),.WL(WL200));
sram_cell_6t_5 inst_cell_200_46 (.BL(BL46),.BLN(BLN46),.WL(WL200));
sram_cell_6t_5 inst_cell_200_47 (.BL(BL47),.BLN(BLN47),.WL(WL200));
sram_cell_6t_5 inst_cell_200_48 (.BL(BL48),.BLN(BLN48),.WL(WL200));
sram_cell_6t_5 inst_cell_200_49 (.BL(BL49),.BLN(BLN49),.WL(WL200));
sram_cell_6t_5 inst_cell_200_50 (.BL(BL50),.BLN(BLN50),.WL(WL200));
sram_cell_6t_5 inst_cell_200_51 (.BL(BL51),.BLN(BLN51),.WL(WL200));
sram_cell_6t_5 inst_cell_200_52 (.BL(BL52),.BLN(BLN52),.WL(WL200));
sram_cell_6t_5 inst_cell_200_53 (.BL(BL53),.BLN(BLN53),.WL(WL200));
sram_cell_6t_5 inst_cell_200_54 (.BL(BL54),.BLN(BLN54),.WL(WL200));
sram_cell_6t_5 inst_cell_200_55 (.BL(BL55),.BLN(BLN55),.WL(WL200));
sram_cell_6t_5 inst_cell_200_56 (.BL(BL56),.BLN(BLN56),.WL(WL200));
sram_cell_6t_5 inst_cell_200_57 (.BL(BL57),.BLN(BLN57),.WL(WL200));
sram_cell_6t_5 inst_cell_200_58 (.BL(BL58),.BLN(BLN58),.WL(WL200));
sram_cell_6t_5 inst_cell_200_59 (.BL(BL59),.BLN(BLN59),.WL(WL200));
sram_cell_6t_5 inst_cell_200_60 (.BL(BL60),.BLN(BLN60),.WL(WL200));
sram_cell_6t_5 inst_cell_200_61 (.BL(BL61),.BLN(BLN61),.WL(WL200));
sram_cell_6t_5 inst_cell_200_62 (.BL(BL62),.BLN(BLN62),.WL(WL200));
sram_cell_6t_5 inst_cell_200_63 (.BL(BL63),.BLN(BLN63),.WL(WL200));
sram_cell_6t_5 inst_cell_200_64 (.BL(BL64),.BLN(BLN64),.WL(WL200));
sram_cell_6t_5 inst_cell_200_65 (.BL(BL65),.BLN(BLN65),.WL(WL200));
sram_cell_6t_5 inst_cell_200_66 (.BL(BL66),.BLN(BLN66),.WL(WL200));
sram_cell_6t_5 inst_cell_200_67 (.BL(BL67),.BLN(BLN67),.WL(WL200));
sram_cell_6t_5 inst_cell_200_68 (.BL(BL68),.BLN(BLN68),.WL(WL200));
sram_cell_6t_5 inst_cell_200_69 (.BL(BL69),.BLN(BLN69),.WL(WL200));
sram_cell_6t_5 inst_cell_200_70 (.BL(BL70),.BLN(BLN70),.WL(WL200));
sram_cell_6t_5 inst_cell_200_71 (.BL(BL71),.BLN(BLN71),.WL(WL200));
sram_cell_6t_5 inst_cell_200_72 (.BL(BL72),.BLN(BLN72),.WL(WL200));
sram_cell_6t_5 inst_cell_200_73 (.BL(BL73),.BLN(BLN73),.WL(WL200));
sram_cell_6t_5 inst_cell_200_74 (.BL(BL74),.BLN(BLN74),.WL(WL200));
sram_cell_6t_5 inst_cell_200_75 (.BL(BL75),.BLN(BLN75),.WL(WL200));
sram_cell_6t_5 inst_cell_200_76 (.BL(BL76),.BLN(BLN76),.WL(WL200));
sram_cell_6t_5 inst_cell_200_77 (.BL(BL77),.BLN(BLN77),.WL(WL200));
sram_cell_6t_5 inst_cell_200_78 (.BL(BL78),.BLN(BLN78),.WL(WL200));
sram_cell_6t_5 inst_cell_200_79 (.BL(BL79),.BLN(BLN79),.WL(WL200));
sram_cell_6t_5 inst_cell_200_80 (.BL(BL80),.BLN(BLN80),.WL(WL200));
sram_cell_6t_5 inst_cell_200_81 (.BL(BL81),.BLN(BLN81),.WL(WL200));
sram_cell_6t_5 inst_cell_200_82 (.BL(BL82),.BLN(BLN82),.WL(WL200));
sram_cell_6t_5 inst_cell_200_83 (.BL(BL83),.BLN(BLN83),.WL(WL200));
sram_cell_6t_5 inst_cell_200_84 (.BL(BL84),.BLN(BLN84),.WL(WL200));
sram_cell_6t_5 inst_cell_200_85 (.BL(BL85),.BLN(BLN85),.WL(WL200));
sram_cell_6t_5 inst_cell_200_86 (.BL(BL86),.BLN(BLN86),.WL(WL200));
sram_cell_6t_5 inst_cell_200_87 (.BL(BL87),.BLN(BLN87),.WL(WL200));
sram_cell_6t_5 inst_cell_200_88 (.BL(BL88),.BLN(BLN88),.WL(WL200));
sram_cell_6t_5 inst_cell_200_89 (.BL(BL89),.BLN(BLN89),.WL(WL200));
sram_cell_6t_5 inst_cell_200_90 (.BL(BL90),.BLN(BLN90),.WL(WL200));
sram_cell_6t_5 inst_cell_200_91 (.BL(BL91),.BLN(BLN91),.WL(WL200));
sram_cell_6t_5 inst_cell_200_92 (.BL(BL92),.BLN(BLN92),.WL(WL200));
sram_cell_6t_5 inst_cell_200_93 (.BL(BL93),.BLN(BLN93),.WL(WL200));
sram_cell_6t_5 inst_cell_200_94 (.BL(BL94),.BLN(BLN94),.WL(WL200));
sram_cell_6t_5 inst_cell_200_95 (.BL(BL95),.BLN(BLN95),.WL(WL200));
sram_cell_6t_5 inst_cell_200_96 (.BL(BL96),.BLN(BLN96),.WL(WL200));
sram_cell_6t_5 inst_cell_200_97 (.BL(BL97),.BLN(BLN97),.WL(WL200));
sram_cell_6t_5 inst_cell_200_98 (.BL(BL98),.BLN(BLN98),.WL(WL200));
sram_cell_6t_5 inst_cell_200_99 (.BL(BL99),.BLN(BLN99),.WL(WL200));
sram_cell_6t_5 inst_cell_200_100 (.BL(BL100),.BLN(BLN100),.WL(WL200));
sram_cell_6t_5 inst_cell_200_101 (.BL(BL101),.BLN(BLN101),.WL(WL200));
sram_cell_6t_5 inst_cell_200_102 (.BL(BL102),.BLN(BLN102),.WL(WL200));
sram_cell_6t_5 inst_cell_200_103 (.BL(BL103),.BLN(BLN103),.WL(WL200));
sram_cell_6t_5 inst_cell_200_104 (.BL(BL104),.BLN(BLN104),.WL(WL200));
sram_cell_6t_5 inst_cell_200_105 (.BL(BL105),.BLN(BLN105),.WL(WL200));
sram_cell_6t_5 inst_cell_200_106 (.BL(BL106),.BLN(BLN106),.WL(WL200));
sram_cell_6t_5 inst_cell_200_107 (.BL(BL107),.BLN(BLN107),.WL(WL200));
sram_cell_6t_5 inst_cell_200_108 (.BL(BL108),.BLN(BLN108),.WL(WL200));
sram_cell_6t_5 inst_cell_200_109 (.BL(BL109),.BLN(BLN109),.WL(WL200));
sram_cell_6t_5 inst_cell_200_110 (.BL(BL110),.BLN(BLN110),.WL(WL200));
sram_cell_6t_5 inst_cell_200_111 (.BL(BL111),.BLN(BLN111),.WL(WL200));
sram_cell_6t_5 inst_cell_200_112 (.BL(BL112),.BLN(BLN112),.WL(WL200));
sram_cell_6t_5 inst_cell_200_113 (.BL(BL113),.BLN(BLN113),.WL(WL200));
sram_cell_6t_5 inst_cell_200_114 (.BL(BL114),.BLN(BLN114),.WL(WL200));
sram_cell_6t_5 inst_cell_200_115 (.BL(BL115),.BLN(BLN115),.WL(WL200));
sram_cell_6t_5 inst_cell_200_116 (.BL(BL116),.BLN(BLN116),.WL(WL200));
sram_cell_6t_5 inst_cell_200_117 (.BL(BL117),.BLN(BLN117),.WL(WL200));
sram_cell_6t_5 inst_cell_200_118 (.BL(BL118),.BLN(BLN118),.WL(WL200));
sram_cell_6t_5 inst_cell_200_119 (.BL(BL119),.BLN(BLN119),.WL(WL200));
sram_cell_6t_5 inst_cell_200_120 (.BL(BL120),.BLN(BLN120),.WL(WL200));
sram_cell_6t_5 inst_cell_200_121 (.BL(BL121),.BLN(BLN121),.WL(WL200));
sram_cell_6t_5 inst_cell_200_122 (.BL(BL122),.BLN(BLN122),.WL(WL200));
sram_cell_6t_5 inst_cell_200_123 (.BL(BL123),.BLN(BLN123),.WL(WL200));
sram_cell_6t_5 inst_cell_200_124 (.BL(BL124),.BLN(BLN124),.WL(WL200));
sram_cell_6t_5 inst_cell_200_125 (.BL(BL125),.BLN(BLN125),.WL(WL200));
sram_cell_6t_5 inst_cell_200_126 (.BL(BL126),.BLN(BLN126),.WL(WL200));
sram_cell_6t_5 inst_cell_200_127 (.BL(BL127),.BLN(BLN127),.WL(WL200));
sram_cell_6t_5 inst_cell_201_0 (.BL(BL0),.BLN(BLN0),.WL(WL201));
sram_cell_6t_5 inst_cell_201_1 (.BL(BL1),.BLN(BLN1),.WL(WL201));
sram_cell_6t_5 inst_cell_201_2 (.BL(BL2),.BLN(BLN2),.WL(WL201));
sram_cell_6t_5 inst_cell_201_3 (.BL(BL3),.BLN(BLN3),.WL(WL201));
sram_cell_6t_5 inst_cell_201_4 (.BL(BL4),.BLN(BLN4),.WL(WL201));
sram_cell_6t_5 inst_cell_201_5 (.BL(BL5),.BLN(BLN5),.WL(WL201));
sram_cell_6t_5 inst_cell_201_6 (.BL(BL6),.BLN(BLN6),.WL(WL201));
sram_cell_6t_5 inst_cell_201_7 (.BL(BL7),.BLN(BLN7),.WL(WL201));
sram_cell_6t_5 inst_cell_201_8 (.BL(BL8),.BLN(BLN8),.WL(WL201));
sram_cell_6t_5 inst_cell_201_9 (.BL(BL9),.BLN(BLN9),.WL(WL201));
sram_cell_6t_5 inst_cell_201_10 (.BL(BL10),.BLN(BLN10),.WL(WL201));
sram_cell_6t_5 inst_cell_201_11 (.BL(BL11),.BLN(BLN11),.WL(WL201));
sram_cell_6t_5 inst_cell_201_12 (.BL(BL12),.BLN(BLN12),.WL(WL201));
sram_cell_6t_5 inst_cell_201_13 (.BL(BL13),.BLN(BLN13),.WL(WL201));
sram_cell_6t_5 inst_cell_201_14 (.BL(BL14),.BLN(BLN14),.WL(WL201));
sram_cell_6t_5 inst_cell_201_15 (.BL(BL15),.BLN(BLN15),.WL(WL201));
sram_cell_6t_5 inst_cell_201_16 (.BL(BL16),.BLN(BLN16),.WL(WL201));
sram_cell_6t_5 inst_cell_201_17 (.BL(BL17),.BLN(BLN17),.WL(WL201));
sram_cell_6t_5 inst_cell_201_18 (.BL(BL18),.BLN(BLN18),.WL(WL201));
sram_cell_6t_5 inst_cell_201_19 (.BL(BL19),.BLN(BLN19),.WL(WL201));
sram_cell_6t_5 inst_cell_201_20 (.BL(BL20),.BLN(BLN20),.WL(WL201));
sram_cell_6t_5 inst_cell_201_21 (.BL(BL21),.BLN(BLN21),.WL(WL201));
sram_cell_6t_5 inst_cell_201_22 (.BL(BL22),.BLN(BLN22),.WL(WL201));
sram_cell_6t_5 inst_cell_201_23 (.BL(BL23),.BLN(BLN23),.WL(WL201));
sram_cell_6t_5 inst_cell_201_24 (.BL(BL24),.BLN(BLN24),.WL(WL201));
sram_cell_6t_5 inst_cell_201_25 (.BL(BL25),.BLN(BLN25),.WL(WL201));
sram_cell_6t_5 inst_cell_201_26 (.BL(BL26),.BLN(BLN26),.WL(WL201));
sram_cell_6t_5 inst_cell_201_27 (.BL(BL27),.BLN(BLN27),.WL(WL201));
sram_cell_6t_5 inst_cell_201_28 (.BL(BL28),.BLN(BLN28),.WL(WL201));
sram_cell_6t_5 inst_cell_201_29 (.BL(BL29),.BLN(BLN29),.WL(WL201));
sram_cell_6t_5 inst_cell_201_30 (.BL(BL30),.BLN(BLN30),.WL(WL201));
sram_cell_6t_5 inst_cell_201_31 (.BL(BL31),.BLN(BLN31),.WL(WL201));
sram_cell_6t_5 inst_cell_201_32 (.BL(BL32),.BLN(BLN32),.WL(WL201));
sram_cell_6t_5 inst_cell_201_33 (.BL(BL33),.BLN(BLN33),.WL(WL201));
sram_cell_6t_5 inst_cell_201_34 (.BL(BL34),.BLN(BLN34),.WL(WL201));
sram_cell_6t_5 inst_cell_201_35 (.BL(BL35),.BLN(BLN35),.WL(WL201));
sram_cell_6t_5 inst_cell_201_36 (.BL(BL36),.BLN(BLN36),.WL(WL201));
sram_cell_6t_5 inst_cell_201_37 (.BL(BL37),.BLN(BLN37),.WL(WL201));
sram_cell_6t_5 inst_cell_201_38 (.BL(BL38),.BLN(BLN38),.WL(WL201));
sram_cell_6t_5 inst_cell_201_39 (.BL(BL39),.BLN(BLN39),.WL(WL201));
sram_cell_6t_5 inst_cell_201_40 (.BL(BL40),.BLN(BLN40),.WL(WL201));
sram_cell_6t_5 inst_cell_201_41 (.BL(BL41),.BLN(BLN41),.WL(WL201));
sram_cell_6t_5 inst_cell_201_42 (.BL(BL42),.BLN(BLN42),.WL(WL201));
sram_cell_6t_5 inst_cell_201_43 (.BL(BL43),.BLN(BLN43),.WL(WL201));
sram_cell_6t_5 inst_cell_201_44 (.BL(BL44),.BLN(BLN44),.WL(WL201));
sram_cell_6t_5 inst_cell_201_45 (.BL(BL45),.BLN(BLN45),.WL(WL201));
sram_cell_6t_5 inst_cell_201_46 (.BL(BL46),.BLN(BLN46),.WL(WL201));
sram_cell_6t_5 inst_cell_201_47 (.BL(BL47),.BLN(BLN47),.WL(WL201));
sram_cell_6t_5 inst_cell_201_48 (.BL(BL48),.BLN(BLN48),.WL(WL201));
sram_cell_6t_5 inst_cell_201_49 (.BL(BL49),.BLN(BLN49),.WL(WL201));
sram_cell_6t_5 inst_cell_201_50 (.BL(BL50),.BLN(BLN50),.WL(WL201));
sram_cell_6t_5 inst_cell_201_51 (.BL(BL51),.BLN(BLN51),.WL(WL201));
sram_cell_6t_5 inst_cell_201_52 (.BL(BL52),.BLN(BLN52),.WL(WL201));
sram_cell_6t_5 inst_cell_201_53 (.BL(BL53),.BLN(BLN53),.WL(WL201));
sram_cell_6t_5 inst_cell_201_54 (.BL(BL54),.BLN(BLN54),.WL(WL201));
sram_cell_6t_5 inst_cell_201_55 (.BL(BL55),.BLN(BLN55),.WL(WL201));
sram_cell_6t_5 inst_cell_201_56 (.BL(BL56),.BLN(BLN56),.WL(WL201));
sram_cell_6t_5 inst_cell_201_57 (.BL(BL57),.BLN(BLN57),.WL(WL201));
sram_cell_6t_5 inst_cell_201_58 (.BL(BL58),.BLN(BLN58),.WL(WL201));
sram_cell_6t_5 inst_cell_201_59 (.BL(BL59),.BLN(BLN59),.WL(WL201));
sram_cell_6t_5 inst_cell_201_60 (.BL(BL60),.BLN(BLN60),.WL(WL201));
sram_cell_6t_5 inst_cell_201_61 (.BL(BL61),.BLN(BLN61),.WL(WL201));
sram_cell_6t_5 inst_cell_201_62 (.BL(BL62),.BLN(BLN62),.WL(WL201));
sram_cell_6t_5 inst_cell_201_63 (.BL(BL63),.BLN(BLN63),.WL(WL201));
sram_cell_6t_5 inst_cell_201_64 (.BL(BL64),.BLN(BLN64),.WL(WL201));
sram_cell_6t_5 inst_cell_201_65 (.BL(BL65),.BLN(BLN65),.WL(WL201));
sram_cell_6t_5 inst_cell_201_66 (.BL(BL66),.BLN(BLN66),.WL(WL201));
sram_cell_6t_5 inst_cell_201_67 (.BL(BL67),.BLN(BLN67),.WL(WL201));
sram_cell_6t_5 inst_cell_201_68 (.BL(BL68),.BLN(BLN68),.WL(WL201));
sram_cell_6t_5 inst_cell_201_69 (.BL(BL69),.BLN(BLN69),.WL(WL201));
sram_cell_6t_5 inst_cell_201_70 (.BL(BL70),.BLN(BLN70),.WL(WL201));
sram_cell_6t_5 inst_cell_201_71 (.BL(BL71),.BLN(BLN71),.WL(WL201));
sram_cell_6t_5 inst_cell_201_72 (.BL(BL72),.BLN(BLN72),.WL(WL201));
sram_cell_6t_5 inst_cell_201_73 (.BL(BL73),.BLN(BLN73),.WL(WL201));
sram_cell_6t_5 inst_cell_201_74 (.BL(BL74),.BLN(BLN74),.WL(WL201));
sram_cell_6t_5 inst_cell_201_75 (.BL(BL75),.BLN(BLN75),.WL(WL201));
sram_cell_6t_5 inst_cell_201_76 (.BL(BL76),.BLN(BLN76),.WL(WL201));
sram_cell_6t_5 inst_cell_201_77 (.BL(BL77),.BLN(BLN77),.WL(WL201));
sram_cell_6t_5 inst_cell_201_78 (.BL(BL78),.BLN(BLN78),.WL(WL201));
sram_cell_6t_5 inst_cell_201_79 (.BL(BL79),.BLN(BLN79),.WL(WL201));
sram_cell_6t_5 inst_cell_201_80 (.BL(BL80),.BLN(BLN80),.WL(WL201));
sram_cell_6t_5 inst_cell_201_81 (.BL(BL81),.BLN(BLN81),.WL(WL201));
sram_cell_6t_5 inst_cell_201_82 (.BL(BL82),.BLN(BLN82),.WL(WL201));
sram_cell_6t_5 inst_cell_201_83 (.BL(BL83),.BLN(BLN83),.WL(WL201));
sram_cell_6t_5 inst_cell_201_84 (.BL(BL84),.BLN(BLN84),.WL(WL201));
sram_cell_6t_5 inst_cell_201_85 (.BL(BL85),.BLN(BLN85),.WL(WL201));
sram_cell_6t_5 inst_cell_201_86 (.BL(BL86),.BLN(BLN86),.WL(WL201));
sram_cell_6t_5 inst_cell_201_87 (.BL(BL87),.BLN(BLN87),.WL(WL201));
sram_cell_6t_5 inst_cell_201_88 (.BL(BL88),.BLN(BLN88),.WL(WL201));
sram_cell_6t_5 inst_cell_201_89 (.BL(BL89),.BLN(BLN89),.WL(WL201));
sram_cell_6t_5 inst_cell_201_90 (.BL(BL90),.BLN(BLN90),.WL(WL201));
sram_cell_6t_5 inst_cell_201_91 (.BL(BL91),.BLN(BLN91),.WL(WL201));
sram_cell_6t_5 inst_cell_201_92 (.BL(BL92),.BLN(BLN92),.WL(WL201));
sram_cell_6t_5 inst_cell_201_93 (.BL(BL93),.BLN(BLN93),.WL(WL201));
sram_cell_6t_5 inst_cell_201_94 (.BL(BL94),.BLN(BLN94),.WL(WL201));
sram_cell_6t_5 inst_cell_201_95 (.BL(BL95),.BLN(BLN95),.WL(WL201));
sram_cell_6t_5 inst_cell_201_96 (.BL(BL96),.BLN(BLN96),.WL(WL201));
sram_cell_6t_5 inst_cell_201_97 (.BL(BL97),.BLN(BLN97),.WL(WL201));
sram_cell_6t_5 inst_cell_201_98 (.BL(BL98),.BLN(BLN98),.WL(WL201));
sram_cell_6t_5 inst_cell_201_99 (.BL(BL99),.BLN(BLN99),.WL(WL201));
sram_cell_6t_5 inst_cell_201_100 (.BL(BL100),.BLN(BLN100),.WL(WL201));
sram_cell_6t_5 inst_cell_201_101 (.BL(BL101),.BLN(BLN101),.WL(WL201));
sram_cell_6t_5 inst_cell_201_102 (.BL(BL102),.BLN(BLN102),.WL(WL201));
sram_cell_6t_5 inst_cell_201_103 (.BL(BL103),.BLN(BLN103),.WL(WL201));
sram_cell_6t_5 inst_cell_201_104 (.BL(BL104),.BLN(BLN104),.WL(WL201));
sram_cell_6t_5 inst_cell_201_105 (.BL(BL105),.BLN(BLN105),.WL(WL201));
sram_cell_6t_5 inst_cell_201_106 (.BL(BL106),.BLN(BLN106),.WL(WL201));
sram_cell_6t_5 inst_cell_201_107 (.BL(BL107),.BLN(BLN107),.WL(WL201));
sram_cell_6t_5 inst_cell_201_108 (.BL(BL108),.BLN(BLN108),.WL(WL201));
sram_cell_6t_5 inst_cell_201_109 (.BL(BL109),.BLN(BLN109),.WL(WL201));
sram_cell_6t_5 inst_cell_201_110 (.BL(BL110),.BLN(BLN110),.WL(WL201));
sram_cell_6t_5 inst_cell_201_111 (.BL(BL111),.BLN(BLN111),.WL(WL201));
sram_cell_6t_5 inst_cell_201_112 (.BL(BL112),.BLN(BLN112),.WL(WL201));
sram_cell_6t_5 inst_cell_201_113 (.BL(BL113),.BLN(BLN113),.WL(WL201));
sram_cell_6t_5 inst_cell_201_114 (.BL(BL114),.BLN(BLN114),.WL(WL201));
sram_cell_6t_5 inst_cell_201_115 (.BL(BL115),.BLN(BLN115),.WL(WL201));
sram_cell_6t_5 inst_cell_201_116 (.BL(BL116),.BLN(BLN116),.WL(WL201));
sram_cell_6t_5 inst_cell_201_117 (.BL(BL117),.BLN(BLN117),.WL(WL201));
sram_cell_6t_5 inst_cell_201_118 (.BL(BL118),.BLN(BLN118),.WL(WL201));
sram_cell_6t_5 inst_cell_201_119 (.BL(BL119),.BLN(BLN119),.WL(WL201));
sram_cell_6t_5 inst_cell_201_120 (.BL(BL120),.BLN(BLN120),.WL(WL201));
sram_cell_6t_5 inst_cell_201_121 (.BL(BL121),.BLN(BLN121),.WL(WL201));
sram_cell_6t_5 inst_cell_201_122 (.BL(BL122),.BLN(BLN122),.WL(WL201));
sram_cell_6t_5 inst_cell_201_123 (.BL(BL123),.BLN(BLN123),.WL(WL201));
sram_cell_6t_5 inst_cell_201_124 (.BL(BL124),.BLN(BLN124),.WL(WL201));
sram_cell_6t_5 inst_cell_201_125 (.BL(BL125),.BLN(BLN125),.WL(WL201));
sram_cell_6t_5 inst_cell_201_126 (.BL(BL126),.BLN(BLN126),.WL(WL201));
sram_cell_6t_5 inst_cell_201_127 (.BL(BL127),.BLN(BLN127),.WL(WL201));
sram_cell_6t_5 inst_cell_202_0 (.BL(BL0),.BLN(BLN0),.WL(WL202));
sram_cell_6t_5 inst_cell_202_1 (.BL(BL1),.BLN(BLN1),.WL(WL202));
sram_cell_6t_5 inst_cell_202_2 (.BL(BL2),.BLN(BLN2),.WL(WL202));
sram_cell_6t_5 inst_cell_202_3 (.BL(BL3),.BLN(BLN3),.WL(WL202));
sram_cell_6t_5 inst_cell_202_4 (.BL(BL4),.BLN(BLN4),.WL(WL202));
sram_cell_6t_5 inst_cell_202_5 (.BL(BL5),.BLN(BLN5),.WL(WL202));
sram_cell_6t_5 inst_cell_202_6 (.BL(BL6),.BLN(BLN6),.WL(WL202));
sram_cell_6t_5 inst_cell_202_7 (.BL(BL7),.BLN(BLN7),.WL(WL202));
sram_cell_6t_5 inst_cell_202_8 (.BL(BL8),.BLN(BLN8),.WL(WL202));
sram_cell_6t_5 inst_cell_202_9 (.BL(BL9),.BLN(BLN9),.WL(WL202));
sram_cell_6t_5 inst_cell_202_10 (.BL(BL10),.BLN(BLN10),.WL(WL202));
sram_cell_6t_5 inst_cell_202_11 (.BL(BL11),.BLN(BLN11),.WL(WL202));
sram_cell_6t_5 inst_cell_202_12 (.BL(BL12),.BLN(BLN12),.WL(WL202));
sram_cell_6t_5 inst_cell_202_13 (.BL(BL13),.BLN(BLN13),.WL(WL202));
sram_cell_6t_5 inst_cell_202_14 (.BL(BL14),.BLN(BLN14),.WL(WL202));
sram_cell_6t_5 inst_cell_202_15 (.BL(BL15),.BLN(BLN15),.WL(WL202));
sram_cell_6t_5 inst_cell_202_16 (.BL(BL16),.BLN(BLN16),.WL(WL202));
sram_cell_6t_5 inst_cell_202_17 (.BL(BL17),.BLN(BLN17),.WL(WL202));
sram_cell_6t_5 inst_cell_202_18 (.BL(BL18),.BLN(BLN18),.WL(WL202));
sram_cell_6t_5 inst_cell_202_19 (.BL(BL19),.BLN(BLN19),.WL(WL202));
sram_cell_6t_5 inst_cell_202_20 (.BL(BL20),.BLN(BLN20),.WL(WL202));
sram_cell_6t_5 inst_cell_202_21 (.BL(BL21),.BLN(BLN21),.WL(WL202));
sram_cell_6t_5 inst_cell_202_22 (.BL(BL22),.BLN(BLN22),.WL(WL202));
sram_cell_6t_5 inst_cell_202_23 (.BL(BL23),.BLN(BLN23),.WL(WL202));
sram_cell_6t_5 inst_cell_202_24 (.BL(BL24),.BLN(BLN24),.WL(WL202));
sram_cell_6t_5 inst_cell_202_25 (.BL(BL25),.BLN(BLN25),.WL(WL202));
sram_cell_6t_5 inst_cell_202_26 (.BL(BL26),.BLN(BLN26),.WL(WL202));
sram_cell_6t_5 inst_cell_202_27 (.BL(BL27),.BLN(BLN27),.WL(WL202));
sram_cell_6t_5 inst_cell_202_28 (.BL(BL28),.BLN(BLN28),.WL(WL202));
sram_cell_6t_5 inst_cell_202_29 (.BL(BL29),.BLN(BLN29),.WL(WL202));
sram_cell_6t_5 inst_cell_202_30 (.BL(BL30),.BLN(BLN30),.WL(WL202));
sram_cell_6t_5 inst_cell_202_31 (.BL(BL31),.BLN(BLN31),.WL(WL202));
sram_cell_6t_5 inst_cell_202_32 (.BL(BL32),.BLN(BLN32),.WL(WL202));
sram_cell_6t_5 inst_cell_202_33 (.BL(BL33),.BLN(BLN33),.WL(WL202));
sram_cell_6t_5 inst_cell_202_34 (.BL(BL34),.BLN(BLN34),.WL(WL202));
sram_cell_6t_5 inst_cell_202_35 (.BL(BL35),.BLN(BLN35),.WL(WL202));
sram_cell_6t_5 inst_cell_202_36 (.BL(BL36),.BLN(BLN36),.WL(WL202));
sram_cell_6t_5 inst_cell_202_37 (.BL(BL37),.BLN(BLN37),.WL(WL202));
sram_cell_6t_5 inst_cell_202_38 (.BL(BL38),.BLN(BLN38),.WL(WL202));
sram_cell_6t_5 inst_cell_202_39 (.BL(BL39),.BLN(BLN39),.WL(WL202));
sram_cell_6t_5 inst_cell_202_40 (.BL(BL40),.BLN(BLN40),.WL(WL202));
sram_cell_6t_5 inst_cell_202_41 (.BL(BL41),.BLN(BLN41),.WL(WL202));
sram_cell_6t_5 inst_cell_202_42 (.BL(BL42),.BLN(BLN42),.WL(WL202));
sram_cell_6t_5 inst_cell_202_43 (.BL(BL43),.BLN(BLN43),.WL(WL202));
sram_cell_6t_5 inst_cell_202_44 (.BL(BL44),.BLN(BLN44),.WL(WL202));
sram_cell_6t_5 inst_cell_202_45 (.BL(BL45),.BLN(BLN45),.WL(WL202));
sram_cell_6t_5 inst_cell_202_46 (.BL(BL46),.BLN(BLN46),.WL(WL202));
sram_cell_6t_5 inst_cell_202_47 (.BL(BL47),.BLN(BLN47),.WL(WL202));
sram_cell_6t_5 inst_cell_202_48 (.BL(BL48),.BLN(BLN48),.WL(WL202));
sram_cell_6t_5 inst_cell_202_49 (.BL(BL49),.BLN(BLN49),.WL(WL202));
sram_cell_6t_5 inst_cell_202_50 (.BL(BL50),.BLN(BLN50),.WL(WL202));
sram_cell_6t_5 inst_cell_202_51 (.BL(BL51),.BLN(BLN51),.WL(WL202));
sram_cell_6t_5 inst_cell_202_52 (.BL(BL52),.BLN(BLN52),.WL(WL202));
sram_cell_6t_5 inst_cell_202_53 (.BL(BL53),.BLN(BLN53),.WL(WL202));
sram_cell_6t_5 inst_cell_202_54 (.BL(BL54),.BLN(BLN54),.WL(WL202));
sram_cell_6t_5 inst_cell_202_55 (.BL(BL55),.BLN(BLN55),.WL(WL202));
sram_cell_6t_5 inst_cell_202_56 (.BL(BL56),.BLN(BLN56),.WL(WL202));
sram_cell_6t_5 inst_cell_202_57 (.BL(BL57),.BLN(BLN57),.WL(WL202));
sram_cell_6t_5 inst_cell_202_58 (.BL(BL58),.BLN(BLN58),.WL(WL202));
sram_cell_6t_5 inst_cell_202_59 (.BL(BL59),.BLN(BLN59),.WL(WL202));
sram_cell_6t_5 inst_cell_202_60 (.BL(BL60),.BLN(BLN60),.WL(WL202));
sram_cell_6t_5 inst_cell_202_61 (.BL(BL61),.BLN(BLN61),.WL(WL202));
sram_cell_6t_5 inst_cell_202_62 (.BL(BL62),.BLN(BLN62),.WL(WL202));
sram_cell_6t_5 inst_cell_202_63 (.BL(BL63),.BLN(BLN63),.WL(WL202));
sram_cell_6t_5 inst_cell_202_64 (.BL(BL64),.BLN(BLN64),.WL(WL202));
sram_cell_6t_5 inst_cell_202_65 (.BL(BL65),.BLN(BLN65),.WL(WL202));
sram_cell_6t_5 inst_cell_202_66 (.BL(BL66),.BLN(BLN66),.WL(WL202));
sram_cell_6t_5 inst_cell_202_67 (.BL(BL67),.BLN(BLN67),.WL(WL202));
sram_cell_6t_5 inst_cell_202_68 (.BL(BL68),.BLN(BLN68),.WL(WL202));
sram_cell_6t_5 inst_cell_202_69 (.BL(BL69),.BLN(BLN69),.WL(WL202));
sram_cell_6t_5 inst_cell_202_70 (.BL(BL70),.BLN(BLN70),.WL(WL202));
sram_cell_6t_5 inst_cell_202_71 (.BL(BL71),.BLN(BLN71),.WL(WL202));
sram_cell_6t_5 inst_cell_202_72 (.BL(BL72),.BLN(BLN72),.WL(WL202));
sram_cell_6t_5 inst_cell_202_73 (.BL(BL73),.BLN(BLN73),.WL(WL202));
sram_cell_6t_5 inst_cell_202_74 (.BL(BL74),.BLN(BLN74),.WL(WL202));
sram_cell_6t_5 inst_cell_202_75 (.BL(BL75),.BLN(BLN75),.WL(WL202));
sram_cell_6t_5 inst_cell_202_76 (.BL(BL76),.BLN(BLN76),.WL(WL202));
sram_cell_6t_5 inst_cell_202_77 (.BL(BL77),.BLN(BLN77),.WL(WL202));
sram_cell_6t_5 inst_cell_202_78 (.BL(BL78),.BLN(BLN78),.WL(WL202));
sram_cell_6t_5 inst_cell_202_79 (.BL(BL79),.BLN(BLN79),.WL(WL202));
sram_cell_6t_5 inst_cell_202_80 (.BL(BL80),.BLN(BLN80),.WL(WL202));
sram_cell_6t_5 inst_cell_202_81 (.BL(BL81),.BLN(BLN81),.WL(WL202));
sram_cell_6t_5 inst_cell_202_82 (.BL(BL82),.BLN(BLN82),.WL(WL202));
sram_cell_6t_5 inst_cell_202_83 (.BL(BL83),.BLN(BLN83),.WL(WL202));
sram_cell_6t_5 inst_cell_202_84 (.BL(BL84),.BLN(BLN84),.WL(WL202));
sram_cell_6t_5 inst_cell_202_85 (.BL(BL85),.BLN(BLN85),.WL(WL202));
sram_cell_6t_5 inst_cell_202_86 (.BL(BL86),.BLN(BLN86),.WL(WL202));
sram_cell_6t_5 inst_cell_202_87 (.BL(BL87),.BLN(BLN87),.WL(WL202));
sram_cell_6t_5 inst_cell_202_88 (.BL(BL88),.BLN(BLN88),.WL(WL202));
sram_cell_6t_5 inst_cell_202_89 (.BL(BL89),.BLN(BLN89),.WL(WL202));
sram_cell_6t_5 inst_cell_202_90 (.BL(BL90),.BLN(BLN90),.WL(WL202));
sram_cell_6t_5 inst_cell_202_91 (.BL(BL91),.BLN(BLN91),.WL(WL202));
sram_cell_6t_5 inst_cell_202_92 (.BL(BL92),.BLN(BLN92),.WL(WL202));
sram_cell_6t_5 inst_cell_202_93 (.BL(BL93),.BLN(BLN93),.WL(WL202));
sram_cell_6t_5 inst_cell_202_94 (.BL(BL94),.BLN(BLN94),.WL(WL202));
sram_cell_6t_5 inst_cell_202_95 (.BL(BL95),.BLN(BLN95),.WL(WL202));
sram_cell_6t_5 inst_cell_202_96 (.BL(BL96),.BLN(BLN96),.WL(WL202));
sram_cell_6t_5 inst_cell_202_97 (.BL(BL97),.BLN(BLN97),.WL(WL202));
sram_cell_6t_5 inst_cell_202_98 (.BL(BL98),.BLN(BLN98),.WL(WL202));
sram_cell_6t_5 inst_cell_202_99 (.BL(BL99),.BLN(BLN99),.WL(WL202));
sram_cell_6t_5 inst_cell_202_100 (.BL(BL100),.BLN(BLN100),.WL(WL202));
sram_cell_6t_5 inst_cell_202_101 (.BL(BL101),.BLN(BLN101),.WL(WL202));
sram_cell_6t_5 inst_cell_202_102 (.BL(BL102),.BLN(BLN102),.WL(WL202));
sram_cell_6t_5 inst_cell_202_103 (.BL(BL103),.BLN(BLN103),.WL(WL202));
sram_cell_6t_5 inst_cell_202_104 (.BL(BL104),.BLN(BLN104),.WL(WL202));
sram_cell_6t_5 inst_cell_202_105 (.BL(BL105),.BLN(BLN105),.WL(WL202));
sram_cell_6t_5 inst_cell_202_106 (.BL(BL106),.BLN(BLN106),.WL(WL202));
sram_cell_6t_5 inst_cell_202_107 (.BL(BL107),.BLN(BLN107),.WL(WL202));
sram_cell_6t_5 inst_cell_202_108 (.BL(BL108),.BLN(BLN108),.WL(WL202));
sram_cell_6t_5 inst_cell_202_109 (.BL(BL109),.BLN(BLN109),.WL(WL202));
sram_cell_6t_5 inst_cell_202_110 (.BL(BL110),.BLN(BLN110),.WL(WL202));
sram_cell_6t_5 inst_cell_202_111 (.BL(BL111),.BLN(BLN111),.WL(WL202));
sram_cell_6t_5 inst_cell_202_112 (.BL(BL112),.BLN(BLN112),.WL(WL202));
sram_cell_6t_5 inst_cell_202_113 (.BL(BL113),.BLN(BLN113),.WL(WL202));
sram_cell_6t_5 inst_cell_202_114 (.BL(BL114),.BLN(BLN114),.WL(WL202));
sram_cell_6t_5 inst_cell_202_115 (.BL(BL115),.BLN(BLN115),.WL(WL202));
sram_cell_6t_5 inst_cell_202_116 (.BL(BL116),.BLN(BLN116),.WL(WL202));
sram_cell_6t_5 inst_cell_202_117 (.BL(BL117),.BLN(BLN117),.WL(WL202));
sram_cell_6t_5 inst_cell_202_118 (.BL(BL118),.BLN(BLN118),.WL(WL202));
sram_cell_6t_5 inst_cell_202_119 (.BL(BL119),.BLN(BLN119),.WL(WL202));
sram_cell_6t_5 inst_cell_202_120 (.BL(BL120),.BLN(BLN120),.WL(WL202));
sram_cell_6t_5 inst_cell_202_121 (.BL(BL121),.BLN(BLN121),.WL(WL202));
sram_cell_6t_5 inst_cell_202_122 (.BL(BL122),.BLN(BLN122),.WL(WL202));
sram_cell_6t_5 inst_cell_202_123 (.BL(BL123),.BLN(BLN123),.WL(WL202));
sram_cell_6t_5 inst_cell_202_124 (.BL(BL124),.BLN(BLN124),.WL(WL202));
sram_cell_6t_5 inst_cell_202_125 (.BL(BL125),.BLN(BLN125),.WL(WL202));
sram_cell_6t_5 inst_cell_202_126 (.BL(BL126),.BLN(BLN126),.WL(WL202));
sram_cell_6t_5 inst_cell_202_127 (.BL(BL127),.BLN(BLN127),.WL(WL202));
sram_cell_6t_5 inst_cell_203_0 (.BL(BL0),.BLN(BLN0),.WL(WL203));
sram_cell_6t_5 inst_cell_203_1 (.BL(BL1),.BLN(BLN1),.WL(WL203));
sram_cell_6t_5 inst_cell_203_2 (.BL(BL2),.BLN(BLN2),.WL(WL203));
sram_cell_6t_5 inst_cell_203_3 (.BL(BL3),.BLN(BLN3),.WL(WL203));
sram_cell_6t_5 inst_cell_203_4 (.BL(BL4),.BLN(BLN4),.WL(WL203));
sram_cell_6t_5 inst_cell_203_5 (.BL(BL5),.BLN(BLN5),.WL(WL203));
sram_cell_6t_5 inst_cell_203_6 (.BL(BL6),.BLN(BLN6),.WL(WL203));
sram_cell_6t_5 inst_cell_203_7 (.BL(BL7),.BLN(BLN7),.WL(WL203));
sram_cell_6t_5 inst_cell_203_8 (.BL(BL8),.BLN(BLN8),.WL(WL203));
sram_cell_6t_5 inst_cell_203_9 (.BL(BL9),.BLN(BLN9),.WL(WL203));
sram_cell_6t_5 inst_cell_203_10 (.BL(BL10),.BLN(BLN10),.WL(WL203));
sram_cell_6t_5 inst_cell_203_11 (.BL(BL11),.BLN(BLN11),.WL(WL203));
sram_cell_6t_5 inst_cell_203_12 (.BL(BL12),.BLN(BLN12),.WL(WL203));
sram_cell_6t_5 inst_cell_203_13 (.BL(BL13),.BLN(BLN13),.WL(WL203));
sram_cell_6t_5 inst_cell_203_14 (.BL(BL14),.BLN(BLN14),.WL(WL203));
sram_cell_6t_5 inst_cell_203_15 (.BL(BL15),.BLN(BLN15),.WL(WL203));
sram_cell_6t_5 inst_cell_203_16 (.BL(BL16),.BLN(BLN16),.WL(WL203));
sram_cell_6t_5 inst_cell_203_17 (.BL(BL17),.BLN(BLN17),.WL(WL203));
sram_cell_6t_5 inst_cell_203_18 (.BL(BL18),.BLN(BLN18),.WL(WL203));
sram_cell_6t_5 inst_cell_203_19 (.BL(BL19),.BLN(BLN19),.WL(WL203));
sram_cell_6t_5 inst_cell_203_20 (.BL(BL20),.BLN(BLN20),.WL(WL203));
sram_cell_6t_5 inst_cell_203_21 (.BL(BL21),.BLN(BLN21),.WL(WL203));
sram_cell_6t_5 inst_cell_203_22 (.BL(BL22),.BLN(BLN22),.WL(WL203));
sram_cell_6t_5 inst_cell_203_23 (.BL(BL23),.BLN(BLN23),.WL(WL203));
sram_cell_6t_5 inst_cell_203_24 (.BL(BL24),.BLN(BLN24),.WL(WL203));
sram_cell_6t_5 inst_cell_203_25 (.BL(BL25),.BLN(BLN25),.WL(WL203));
sram_cell_6t_5 inst_cell_203_26 (.BL(BL26),.BLN(BLN26),.WL(WL203));
sram_cell_6t_5 inst_cell_203_27 (.BL(BL27),.BLN(BLN27),.WL(WL203));
sram_cell_6t_5 inst_cell_203_28 (.BL(BL28),.BLN(BLN28),.WL(WL203));
sram_cell_6t_5 inst_cell_203_29 (.BL(BL29),.BLN(BLN29),.WL(WL203));
sram_cell_6t_5 inst_cell_203_30 (.BL(BL30),.BLN(BLN30),.WL(WL203));
sram_cell_6t_5 inst_cell_203_31 (.BL(BL31),.BLN(BLN31),.WL(WL203));
sram_cell_6t_5 inst_cell_203_32 (.BL(BL32),.BLN(BLN32),.WL(WL203));
sram_cell_6t_5 inst_cell_203_33 (.BL(BL33),.BLN(BLN33),.WL(WL203));
sram_cell_6t_5 inst_cell_203_34 (.BL(BL34),.BLN(BLN34),.WL(WL203));
sram_cell_6t_5 inst_cell_203_35 (.BL(BL35),.BLN(BLN35),.WL(WL203));
sram_cell_6t_5 inst_cell_203_36 (.BL(BL36),.BLN(BLN36),.WL(WL203));
sram_cell_6t_5 inst_cell_203_37 (.BL(BL37),.BLN(BLN37),.WL(WL203));
sram_cell_6t_5 inst_cell_203_38 (.BL(BL38),.BLN(BLN38),.WL(WL203));
sram_cell_6t_5 inst_cell_203_39 (.BL(BL39),.BLN(BLN39),.WL(WL203));
sram_cell_6t_5 inst_cell_203_40 (.BL(BL40),.BLN(BLN40),.WL(WL203));
sram_cell_6t_5 inst_cell_203_41 (.BL(BL41),.BLN(BLN41),.WL(WL203));
sram_cell_6t_5 inst_cell_203_42 (.BL(BL42),.BLN(BLN42),.WL(WL203));
sram_cell_6t_5 inst_cell_203_43 (.BL(BL43),.BLN(BLN43),.WL(WL203));
sram_cell_6t_5 inst_cell_203_44 (.BL(BL44),.BLN(BLN44),.WL(WL203));
sram_cell_6t_5 inst_cell_203_45 (.BL(BL45),.BLN(BLN45),.WL(WL203));
sram_cell_6t_5 inst_cell_203_46 (.BL(BL46),.BLN(BLN46),.WL(WL203));
sram_cell_6t_5 inst_cell_203_47 (.BL(BL47),.BLN(BLN47),.WL(WL203));
sram_cell_6t_5 inst_cell_203_48 (.BL(BL48),.BLN(BLN48),.WL(WL203));
sram_cell_6t_5 inst_cell_203_49 (.BL(BL49),.BLN(BLN49),.WL(WL203));
sram_cell_6t_5 inst_cell_203_50 (.BL(BL50),.BLN(BLN50),.WL(WL203));
sram_cell_6t_5 inst_cell_203_51 (.BL(BL51),.BLN(BLN51),.WL(WL203));
sram_cell_6t_5 inst_cell_203_52 (.BL(BL52),.BLN(BLN52),.WL(WL203));
sram_cell_6t_5 inst_cell_203_53 (.BL(BL53),.BLN(BLN53),.WL(WL203));
sram_cell_6t_5 inst_cell_203_54 (.BL(BL54),.BLN(BLN54),.WL(WL203));
sram_cell_6t_5 inst_cell_203_55 (.BL(BL55),.BLN(BLN55),.WL(WL203));
sram_cell_6t_5 inst_cell_203_56 (.BL(BL56),.BLN(BLN56),.WL(WL203));
sram_cell_6t_5 inst_cell_203_57 (.BL(BL57),.BLN(BLN57),.WL(WL203));
sram_cell_6t_5 inst_cell_203_58 (.BL(BL58),.BLN(BLN58),.WL(WL203));
sram_cell_6t_5 inst_cell_203_59 (.BL(BL59),.BLN(BLN59),.WL(WL203));
sram_cell_6t_5 inst_cell_203_60 (.BL(BL60),.BLN(BLN60),.WL(WL203));
sram_cell_6t_5 inst_cell_203_61 (.BL(BL61),.BLN(BLN61),.WL(WL203));
sram_cell_6t_5 inst_cell_203_62 (.BL(BL62),.BLN(BLN62),.WL(WL203));
sram_cell_6t_5 inst_cell_203_63 (.BL(BL63),.BLN(BLN63),.WL(WL203));
sram_cell_6t_5 inst_cell_203_64 (.BL(BL64),.BLN(BLN64),.WL(WL203));
sram_cell_6t_5 inst_cell_203_65 (.BL(BL65),.BLN(BLN65),.WL(WL203));
sram_cell_6t_5 inst_cell_203_66 (.BL(BL66),.BLN(BLN66),.WL(WL203));
sram_cell_6t_5 inst_cell_203_67 (.BL(BL67),.BLN(BLN67),.WL(WL203));
sram_cell_6t_5 inst_cell_203_68 (.BL(BL68),.BLN(BLN68),.WL(WL203));
sram_cell_6t_5 inst_cell_203_69 (.BL(BL69),.BLN(BLN69),.WL(WL203));
sram_cell_6t_5 inst_cell_203_70 (.BL(BL70),.BLN(BLN70),.WL(WL203));
sram_cell_6t_5 inst_cell_203_71 (.BL(BL71),.BLN(BLN71),.WL(WL203));
sram_cell_6t_5 inst_cell_203_72 (.BL(BL72),.BLN(BLN72),.WL(WL203));
sram_cell_6t_5 inst_cell_203_73 (.BL(BL73),.BLN(BLN73),.WL(WL203));
sram_cell_6t_5 inst_cell_203_74 (.BL(BL74),.BLN(BLN74),.WL(WL203));
sram_cell_6t_5 inst_cell_203_75 (.BL(BL75),.BLN(BLN75),.WL(WL203));
sram_cell_6t_5 inst_cell_203_76 (.BL(BL76),.BLN(BLN76),.WL(WL203));
sram_cell_6t_5 inst_cell_203_77 (.BL(BL77),.BLN(BLN77),.WL(WL203));
sram_cell_6t_5 inst_cell_203_78 (.BL(BL78),.BLN(BLN78),.WL(WL203));
sram_cell_6t_5 inst_cell_203_79 (.BL(BL79),.BLN(BLN79),.WL(WL203));
sram_cell_6t_5 inst_cell_203_80 (.BL(BL80),.BLN(BLN80),.WL(WL203));
sram_cell_6t_5 inst_cell_203_81 (.BL(BL81),.BLN(BLN81),.WL(WL203));
sram_cell_6t_5 inst_cell_203_82 (.BL(BL82),.BLN(BLN82),.WL(WL203));
sram_cell_6t_5 inst_cell_203_83 (.BL(BL83),.BLN(BLN83),.WL(WL203));
sram_cell_6t_5 inst_cell_203_84 (.BL(BL84),.BLN(BLN84),.WL(WL203));
sram_cell_6t_5 inst_cell_203_85 (.BL(BL85),.BLN(BLN85),.WL(WL203));
sram_cell_6t_5 inst_cell_203_86 (.BL(BL86),.BLN(BLN86),.WL(WL203));
sram_cell_6t_5 inst_cell_203_87 (.BL(BL87),.BLN(BLN87),.WL(WL203));
sram_cell_6t_5 inst_cell_203_88 (.BL(BL88),.BLN(BLN88),.WL(WL203));
sram_cell_6t_5 inst_cell_203_89 (.BL(BL89),.BLN(BLN89),.WL(WL203));
sram_cell_6t_5 inst_cell_203_90 (.BL(BL90),.BLN(BLN90),.WL(WL203));
sram_cell_6t_5 inst_cell_203_91 (.BL(BL91),.BLN(BLN91),.WL(WL203));
sram_cell_6t_5 inst_cell_203_92 (.BL(BL92),.BLN(BLN92),.WL(WL203));
sram_cell_6t_5 inst_cell_203_93 (.BL(BL93),.BLN(BLN93),.WL(WL203));
sram_cell_6t_5 inst_cell_203_94 (.BL(BL94),.BLN(BLN94),.WL(WL203));
sram_cell_6t_5 inst_cell_203_95 (.BL(BL95),.BLN(BLN95),.WL(WL203));
sram_cell_6t_5 inst_cell_203_96 (.BL(BL96),.BLN(BLN96),.WL(WL203));
sram_cell_6t_5 inst_cell_203_97 (.BL(BL97),.BLN(BLN97),.WL(WL203));
sram_cell_6t_5 inst_cell_203_98 (.BL(BL98),.BLN(BLN98),.WL(WL203));
sram_cell_6t_5 inst_cell_203_99 (.BL(BL99),.BLN(BLN99),.WL(WL203));
sram_cell_6t_5 inst_cell_203_100 (.BL(BL100),.BLN(BLN100),.WL(WL203));
sram_cell_6t_5 inst_cell_203_101 (.BL(BL101),.BLN(BLN101),.WL(WL203));
sram_cell_6t_5 inst_cell_203_102 (.BL(BL102),.BLN(BLN102),.WL(WL203));
sram_cell_6t_5 inst_cell_203_103 (.BL(BL103),.BLN(BLN103),.WL(WL203));
sram_cell_6t_5 inst_cell_203_104 (.BL(BL104),.BLN(BLN104),.WL(WL203));
sram_cell_6t_5 inst_cell_203_105 (.BL(BL105),.BLN(BLN105),.WL(WL203));
sram_cell_6t_5 inst_cell_203_106 (.BL(BL106),.BLN(BLN106),.WL(WL203));
sram_cell_6t_5 inst_cell_203_107 (.BL(BL107),.BLN(BLN107),.WL(WL203));
sram_cell_6t_5 inst_cell_203_108 (.BL(BL108),.BLN(BLN108),.WL(WL203));
sram_cell_6t_5 inst_cell_203_109 (.BL(BL109),.BLN(BLN109),.WL(WL203));
sram_cell_6t_5 inst_cell_203_110 (.BL(BL110),.BLN(BLN110),.WL(WL203));
sram_cell_6t_5 inst_cell_203_111 (.BL(BL111),.BLN(BLN111),.WL(WL203));
sram_cell_6t_5 inst_cell_203_112 (.BL(BL112),.BLN(BLN112),.WL(WL203));
sram_cell_6t_5 inst_cell_203_113 (.BL(BL113),.BLN(BLN113),.WL(WL203));
sram_cell_6t_5 inst_cell_203_114 (.BL(BL114),.BLN(BLN114),.WL(WL203));
sram_cell_6t_5 inst_cell_203_115 (.BL(BL115),.BLN(BLN115),.WL(WL203));
sram_cell_6t_5 inst_cell_203_116 (.BL(BL116),.BLN(BLN116),.WL(WL203));
sram_cell_6t_5 inst_cell_203_117 (.BL(BL117),.BLN(BLN117),.WL(WL203));
sram_cell_6t_5 inst_cell_203_118 (.BL(BL118),.BLN(BLN118),.WL(WL203));
sram_cell_6t_5 inst_cell_203_119 (.BL(BL119),.BLN(BLN119),.WL(WL203));
sram_cell_6t_5 inst_cell_203_120 (.BL(BL120),.BLN(BLN120),.WL(WL203));
sram_cell_6t_5 inst_cell_203_121 (.BL(BL121),.BLN(BLN121),.WL(WL203));
sram_cell_6t_5 inst_cell_203_122 (.BL(BL122),.BLN(BLN122),.WL(WL203));
sram_cell_6t_5 inst_cell_203_123 (.BL(BL123),.BLN(BLN123),.WL(WL203));
sram_cell_6t_5 inst_cell_203_124 (.BL(BL124),.BLN(BLN124),.WL(WL203));
sram_cell_6t_5 inst_cell_203_125 (.BL(BL125),.BLN(BLN125),.WL(WL203));
sram_cell_6t_5 inst_cell_203_126 (.BL(BL126),.BLN(BLN126),.WL(WL203));
sram_cell_6t_5 inst_cell_203_127 (.BL(BL127),.BLN(BLN127),.WL(WL203));
sram_cell_6t_5 inst_cell_204_0 (.BL(BL0),.BLN(BLN0),.WL(WL204));
sram_cell_6t_5 inst_cell_204_1 (.BL(BL1),.BLN(BLN1),.WL(WL204));
sram_cell_6t_5 inst_cell_204_2 (.BL(BL2),.BLN(BLN2),.WL(WL204));
sram_cell_6t_5 inst_cell_204_3 (.BL(BL3),.BLN(BLN3),.WL(WL204));
sram_cell_6t_5 inst_cell_204_4 (.BL(BL4),.BLN(BLN4),.WL(WL204));
sram_cell_6t_5 inst_cell_204_5 (.BL(BL5),.BLN(BLN5),.WL(WL204));
sram_cell_6t_5 inst_cell_204_6 (.BL(BL6),.BLN(BLN6),.WL(WL204));
sram_cell_6t_5 inst_cell_204_7 (.BL(BL7),.BLN(BLN7),.WL(WL204));
sram_cell_6t_5 inst_cell_204_8 (.BL(BL8),.BLN(BLN8),.WL(WL204));
sram_cell_6t_5 inst_cell_204_9 (.BL(BL9),.BLN(BLN9),.WL(WL204));
sram_cell_6t_5 inst_cell_204_10 (.BL(BL10),.BLN(BLN10),.WL(WL204));
sram_cell_6t_5 inst_cell_204_11 (.BL(BL11),.BLN(BLN11),.WL(WL204));
sram_cell_6t_5 inst_cell_204_12 (.BL(BL12),.BLN(BLN12),.WL(WL204));
sram_cell_6t_5 inst_cell_204_13 (.BL(BL13),.BLN(BLN13),.WL(WL204));
sram_cell_6t_5 inst_cell_204_14 (.BL(BL14),.BLN(BLN14),.WL(WL204));
sram_cell_6t_5 inst_cell_204_15 (.BL(BL15),.BLN(BLN15),.WL(WL204));
sram_cell_6t_5 inst_cell_204_16 (.BL(BL16),.BLN(BLN16),.WL(WL204));
sram_cell_6t_5 inst_cell_204_17 (.BL(BL17),.BLN(BLN17),.WL(WL204));
sram_cell_6t_5 inst_cell_204_18 (.BL(BL18),.BLN(BLN18),.WL(WL204));
sram_cell_6t_5 inst_cell_204_19 (.BL(BL19),.BLN(BLN19),.WL(WL204));
sram_cell_6t_5 inst_cell_204_20 (.BL(BL20),.BLN(BLN20),.WL(WL204));
sram_cell_6t_5 inst_cell_204_21 (.BL(BL21),.BLN(BLN21),.WL(WL204));
sram_cell_6t_5 inst_cell_204_22 (.BL(BL22),.BLN(BLN22),.WL(WL204));
sram_cell_6t_5 inst_cell_204_23 (.BL(BL23),.BLN(BLN23),.WL(WL204));
sram_cell_6t_5 inst_cell_204_24 (.BL(BL24),.BLN(BLN24),.WL(WL204));
sram_cell_6t_5 inst_cell_204_25 (.BL(BL25),.BLN(BLN25),.WL(WL204));
sram_cell_6t_5 inst_cell_204_26 (.BL(BL26),.BLN(BLN26),.WL(WL204));
sram_cell_6t_5 inst_cell_204_27 (.BL(BL27),.BLN(BLN27),.WL(WL204));
sram_cell_6t_5 inst_cell_204_28 (.BL(BL28),.BLN(BLN28),.WL(WL204));
sram_cell_6t_5 inst_cell_204_29 (.BL(BL29),.BLN(BLN29),.WL(WL204));
sram_cell_6t_5 inst_cell_204_30 (.BL(BL30),.BLN(BLN30),.WL(WL204));
sram_cell_6t_5 inst_cell_204_31 (.BL(BL31),.BLN(BLN31),.WL(WL204));
sram_cell_6t_5 inst_cell_204_32 (.BL(BL32),.BLN(BLN32),.WL(WL204));
sram_cell_6t_5 inst_cell_204_33 (.BL(BL33),.BLN(BLN33),.WL(WL204));
sram_cell_6t_5 inst_cell_204_34 (.BL(BL34),.BLN(BLN34),.WL(WL204));
sram_cell_6t_5 inst_cell_204_35 (.BL(BL35),.BLN(BLN35),.WL(WL204));
sram_cell_6t_5 inst_cell_204_36 (.BL(BL36),.BLN(BLN36),.WL(WL204));
sram_cell_6t_5 inst_cell_204_37 (.BL(BL37),.BLN(BLN37),.WL(WL204));
sram_cell_6t_5 inst_cell_204_38 (.BL(BL38),.BLN(BLN38),.WL(WL204));
sram_cell_6t_5 inst_cell_204_39 (.BL(BL39),.BLN(BLN39),.WL(WL204));
sram_cell_6t_5 inst_cell_204_40 (.BL(BL40),.BLN(BLN40),.WL(WL204));
sram_cell_6t_5 inst_cell_204_41 (.BL(BL41),.BLN(BLN41),.WL(WL204));
sram_cell_6t_5 inst_cell_204_42 (.BL(BL42),.BLN(BLN42),.WL(WL204));
sram_cell_6t_5 inst_cell_204_43 (.BL(BL43),.BLN(BLN43),.WL(WL204));
sram_cell_6t_5 inst_cell_204_44 (.BL(BL44),.BLN(BLN44),.WL(WL204));
sram_cell_6t_5 inst_cell_204_45 (.BL(BL45),.BLN(BLN45),.WL(WL204));
sram_cell_6t_5 inst_cell_204_46 (.BL(BL46),.BLN(BLN46),.WL(WL204));
sram_cell_6t_5 inst_cell_204_47 (.BL(BL47),.BLN(BLN47),.WL(WL204));
sram_cell_6t_5 inst_cell_204_48 (.BL(BL48),.BLN(BLN48),.WL(WL204));
sram_cell_6t_5 inst_cell_204_49 (.BL(BL49),.BLN(BLN49),.WL(WL204));
sram_cell_6t_5 inst_cell_204_50 (.BL(BL50),.BLN(BLN50),.WL(WL204));
sram_cell_6t_5 inst_cell_204_51 (.BL(BL51),.BLN(BLN51),.WL(WL204));
sram_cell_6t_5 inst_cell_204_52 (.BL(BL52),.BLN(BLN52),.WL(WL204));
sram_cell_6t_5 inst_cell_204_53 (.BL(BL53),.BLN(BLN53),.WL(WL204));
sram_cell_6t_5 inst_cell_204_54 (.BL(BL54),.BLN(BLN54),.WL(WL204));
sram_cell_6t_5 inst_cell_204_55 (.BL(BL55),.BLN(BLN55),.WL(WL204));
sram_cell_6t_5 inst_cell_204_56 (.BL(BL56),.BLN(BLN56),.WL(WL204));
sram_cell_6t_5 inst_cell_204_57 (.BL(BL57),.BLN(BLN57),.WL(WL204));
sram_cell_6t_5 inst_cell_204_58 (.BL(BL58),.BLN(BLN58),.WL(WL204));
sram_cell_6t_5 inst_cell_204_59 (.BL(BL59),.BLN(BLN59),.WL(WL204));
sram_cell_6t_5 inst_cell_204_60 (.BL(BL60),.BLN(BLN60),.WL(WL204));
sram_cell_6t_5 inst_cell_204_61 (.BL(BL61),.BLN(BLN61),.WL(WL204));
sram_cell_6t_5 inst_cell_204_62 (.BL(BL62),.BLN(BLN62),.WL(WL204));
sram_cell_6t_5 inst_cell_204_63 (.BL(BL63),.BLN(BLN63),.WL(WL204));
sram_cell_6t_5 inst_cell_204_64 (.BL(BL64),.BLN(BLN64),.WL(WL204));
sram_cell_6t_5 inst_cell_204_65 (.BL(BL65),.BLN(BLN65),.WL(WL204));
sram_cell_6t_5 inst_cell_204_66 (.BL(BL66),.BLN(BLN66),.WL(WL204));
sram_cell_6t_5 inst_cell_204_67 (.BL(BL67),.BLN(BLN67),.WL(WL204));
sram_cell_6t_5 inst_cell_204_68 (.BL(BL68),.BLN(BLN68),.WL(WL204));
sram_cell_6t_5 inst_cell_204_69 (.BL(BL69),.BLN(BLN69),.WL(WL204));
sram_cell_6t_5 inst_cell_204_70 (.BL(BL70),.BLN(BLN70),.WL(WL204));
sram_cell_6t_5 inst_cell_204_71 (.BL(BL71),.BLN(BLN71),.WL(WL204));
sram_cell_6t_5 inst_cell_204_72 (.BL(BL72),.BLN(BLN72),.WL(WL204));
sram_cell_6t_5 inst_cell_204_73 (.BL(BL73),.BLN(BLN73),.WL(WL204));
sram_cell_6t_5 inst_cell_204_74 (.BL(BL74),.BLN(BLN74),.WL(WL204));
sram_cell_6t_5 inst_cell_204_75 (.BL(BL75),.BLN(BLN75),.WL(WL204));
sram_cell_6t_5 inst_cell_204_76 (.BL(BL76),.BLN(BLN76),.WL(WL204));
sram_cell_6t_5 inst_cell_204_77 (.BL(BL77),.BLN(BLN77),.WL(WL204));
sram_cell_6t_5 inst_cell_204_78 (.BL(BL78),.BLN(BLN78),.WL(WL204));
sram_cell_6t_5 inst_cell_204_79 (.BL(BL79),.BLN(BLN79),.WL(WL204));
sram_cell_6t_5 inst_cell_204_80 (.BL(BL80),.BLN(BLN80),.WL(WL204));
sram_cell_6t_5 inst_cell_204_81 (.BL(BL81),.BLN(BLN81),.WL(WL204));
sram_cell_6t_5 inst_cell_204_82 (.BL(BL82),.BLN(BLN82),.WL(WL204));
sram_cell_6t_5 inst_cell_204_83 (.BL(BL83),.BLN(BLN83),.WL(WL204));
sram_cell_6t_5 inst_cell_204_84 (.BL(BL84),.BLN(BLN84),.WL(WL204));
sram_cell_6t_5 inst_cell_204_85 (.BL(BL85),.BLN(BLN85),.WL(WL204));
sram_cell_6t_5 inst_cell_204_86 (.BL(BL86),.BLN(BLN86),.WL(WL204));
sram_cell_6t_5 inst_cell_204_87 (.BL(BL87),.BLN(BLN87),.WL(WL204));
sram_cell_6t_5 inst_cell_204_88 (.BL(BL88),.BLN(BLN88),.WL(WL204));
sram_cell_6t_5 inst_cell_204_89 (.BL(BL89),.BLN(BLN89),.WL(WL204));
sram_cell_6t_5 inst_cell_204_90 (.BL(BL90),.BLN(BLN90),.WL(WL204));
sram_cell_6t_5 inst_cell_204_91 (.BL(BL91),.BLN(BLN91),.WL(WL204));
sram_cell_6t_5 inst_cell_204_92 (.BL(BL92),.BLN(BLN92),.WL(WL204));
sram_cell_6t_5 inst_cell_204_93 (.BL(BL93),.BLN(BLN93),.WL(WL204));
sram_cell_6t_5 inst_cell_204_94 (.BL(BL94),.BLN(BLN94),.WL(WL204));
sram_cell_6t_5 inst_cell_204_95 (.BL(BL95),.BLN(BLN95),.WL(WL204));
sram_cell_6t_5 inst_cell_204_96 (.BL(BL96),.BLN(BLN96),.WL(WL204));
sram_cell_6t_5 inst_cell_204_97 (.BL(BL97),.BLN(BLN97),.WL(WL204));
sram_cell_6t_5 inst_cell_204_98 (.BL(BL98),.BLN(BLN98),.WL(WL204));
sram_cell_6t_5 inst_cell_204_99 (.BL(BL99),.BLN(BLN99),.WL(WL204));
sram_cell_6t_5 inst_cell_204_100 (.BL(BL100),.BLN(BLN100),.WL(WL204));
sram_cell_6t_5 inst_cell_204_101 (.BL(BL101),.BLN(BLN101),.WL(WL204));
sram_cell_6t_5 inst_cell_204_102 (.BL(BL102),.BLN(BLN102),.WL(WL204));
sram_cell_6t_5 inst_cell_204_103 (.BL(BL103),.BLN(BLN103),.WL(WL204));
sram_cell_6t_5 inst_cell_204_104 (.BL(BL104),.BLN(BLN104),.WL(WL204));
sram_cell_6t_5 inst_cell_204_105 (.BL(BL105),.BLN(BLN105),.WL(WL204));
sram_cell_6t_5 inst_cell_204_106 (.BL(BL106),.BLN(BLN106),.WL(WL204));
sram_cell_6t_5 inst_cell_204_107 (.BL(BL107),.BLN(BLN107),.WL(WL204));
sram_cell_6t_5 inst_cell_204_108 (.BL(BL108),.BLN(BLN108),.WL(WL204));
sram_cell_6t_5 inst_cell_204_109 (.BL(BL109),.BLN(BLN109),.WL(WL204));
sram_cell_6t_5 inst_cell_204_110 (.BL(BL110),.BLN(BLN110),.WL(WL204));
sram_cell_6t_5 inst_cell_204_111 (.BL(BL111),.BLN(BLN111),.WL(WL204));
sram_cell_6t_5 inst_cell_204_112 (.BL(BL112),.BLN(BLN112),.WL(WL204));
sram_cell_6t_5 inst_cell_204_113 (.BL(BL113),.BLN(BLN113),.WL(WL204));
sram_cell_6t_5 inst_cell_204_114 (.BL(BL114),.BLN(BLN114),.WL(WL204));
sram_cell_6t_5 inst_cell_204_115 (.BL(BL115),.BLN(BLN115),.WL(WL204));
sram_cell_6t_5 inst_cell_204_116 (.BL(BL116),.BLN(BLN116),.WL(WL204));
sram_cell_6t_5 inst_cell_204_117 (.BL(BL117),.BLN(BLN117),.WL(WL204));
sram_cell_6t_5 inst_cell_204_118 (.BL(BL118),.BLN(BLN118),.WL(WL204));
sram_cell_6t_5 inst_cell_204_119 (.BL(BL119),.BLN(BLN119),.WL(WL204));
sram_cell_6t_5 inst_cell_204_120 (.BL(BL120),.BLN(BLN120),.WL(WL204));
sram_cell_6t_5 inst_cell_204_121 (.BL(BL121),.BLN(BLN121),.WL(WL204));
sram_cell_6t_5 inst_cell_204_122 (.BL(BL122),.BLN(BLN122),.WL(WL204));
sram_cell_6t_5 inst_cell_204_123 (.BL(BL123),.BLN(BLN123),.WL(WL204));
sram_cell_6t_5 inst_cell_204_124 (.BL(BL124),.BLN(BLN124),.WL(WL204));
sram_cell_6t_5 inst_cell_204_125 (.BL(BL125),.BLN(BLN125),.WL(WL204));
sram_cell_6t_5 inst_cell_204_126 (.BL(BL126),.BLN(BLN126),.WL(WL204));
sram_cell_6t_5 inst_cell_204_127 (.BL(BL127),.BLN(BLN127),.WL(WL204));
sram_cell_6t_5 inst_cell_205_0 (.BL(BL0),.BLN(BLN0),.WL(WL205));
sram_cell_6t_5 inst_cell_205_1 (.BL(BL1),.BLN(BLN1),.WL(WL205));
sram_cell_6t_5 inst_cell_205_2 (.BL(BL2),.BLN(BLN2),.WL(WL205));
sram_cell_6t_5 inst_cell_205_3 (.BL(BL3),.BLN(BLN3),.WL(WL205));
sram_cell_6t_5 inst_cell_205_4 (.BL(BL4),.BLN(BLN4),.WL(WL205));
sram_cell_6t_5 inst_cell_205_5 (.BL(BL5),.BLN(BLN5),.WL(WL205));
sram_cell_6t_5 inst_cell_205_6 (.BL(BL6),.BLN(BLN6),.WL(WL205));
sram_cell_6t_5 inst_cell_205_7 (.BL(BL7),.BLN(BLN7),.WL(WL205));
sram_cell_6t_5 inst_cell_205_8 (.BL(BL8),.BLN(BLN8),.WL(WL205));
sram_cell_6t_5 inst_cell_205_9 (.BL(BL9),.BLN(BLN9),.WL(WL205));
sram_cell_6t_5 inst_cell_205_10 (.BL(BL10),.BLN(BLN10),.WL(WL205));
sram_cell_6t_5 inst_cell_205_11 (.BL(BL11),.BLN(BLN11),.WL(WL205));
sram_cell_6t_5 inst_cell_205_12 (.BL(BL12),.BLN(BLN12),.WL(WL205));
sram_cell_6t_5 inst_cell_205_13 (.BL(BL13),.BLN(BLN13),.WL(WL205));
sram_cell_6t_5 inst_cell_205_14 (.BL(BL14),.BLN(BLN14),.WL(WL205));
sram_cell_6t_5 inst_cell_205_15 (.BL(BL15),.BLN(BLN15),.WL(WL205));
sram_cell_6t_5 inst_cell_205_16 (.BL(BL16),.BLN(BLN16),.WL(WL205));
sram_cell_6t_5 inst_cell_205_17 (.BL(BL17),.BLN(BLN17),.WL(WL205));
sram_cell_6t_5 inst_cell_205_18 (.BL(BL18),.BLN(BLN18),.WL(WL205));
sram_cell_6t_5 inst_cell_205_19 (.BL(BL19),.BLN(BLN19),.WL(WL205));
sram_cell_6t_5 inst_cell_205_20 (.BL(BL20),.BLN(BLN20),.WL(WL205));
sram_cell_6t_5 inst_cell_205_21 (.BL(BL21),.BLN(BLN21),.WL(WL205));
sram_cell_6t_5 inst_cell_205_22 (.BL(BL22),.BLN(BLN22),.WL(WL205));
sram_cell_6t_5 inst_cell_205_23 (.BL(BL23),.BLN(BLN23),.WL(WL205));
sram_cell_6t_5 inst_cell_205_24 (.BL(BL24),.BLN(BLN24),.WL(WL205));
sram_cell_6t_5 inst_cell_205_25 (.BL(BL25),.BLN(BLN25),.WL(WL205));
sram_cell_6t_5 inst_cell_205_26 (.BL(BL26),.BLN(BLN26),.WL(WL205));
sram_cell_6t_5 inst_cell_205_27 (.BL(BL27),.BLN(BLN27),.WL(WL205));
sram_cell_6t_5 inst_cell_205_28 (.BL(BL28),.BLN(BLN28),.WL(WL205));
sram_cell_6t_5 inst_cell_205_29 (.BL(BL29),.BLN(BLN29),.WL(WL205));
sram_cell_6t_5 inst_cell_205_30 (.BL(BL30),.BLN(BLN30),.WL(WL205));
sram_cell_6t_5 inst_cell_205_31 (.BL(BL31),.BLN(BLN31),.WL(WL205));
sram_cell_6t_5 inst_cell_205_32 (.BL(BL32),.BLN(BLN32),.WL(WL205));
sram_cell_6t_5 inst_cell_205_33 (.BL(BL33),.BLN(BLN33),.WL(WL205));
sram_cell_6t_5 inst_cell_205_34 (.BL(BL34),.BLN(BLN34),.WL(WL205));
sram_cell_6t_5 inst_cell_205_35 (.BL(BL35),.BLN(BLN35),.WL(WL205));
sram_cell_6t_5 inst_cell_205_36 (.BL(BL36),.BLN(BLN36),.WL(WL205));
sram_cell_6t_5 inst_cell_205_37 (.BL(BL37),.BLN(BLN37),.WL(WL205));
sram_cell_6t_5 inst_cell_205_38 (.BL(BL38),.BLN(BLN38),.WL(WL205));
sram_cell_6t_5 inst_cell_205_39 (.BL(BL39),.BLN(BLN39),.WL(WL205));
sram_cell_6t_5 inst_cell_205_40 (.BL(BL40),.BLN(BLN40),.WL(WL205));
sram_cell_6t_5 inst_cell_205_41 (.BL(BL41),.BLN(BLN41),.WL(WL205));
sram_cell_6t_5 inst_cell_205_42 (.BL(BL42),.BLN(BLN42),.WL(WL205));
sram_cell_6t_5 inst_cell_205_43 (.BL(BL43),.BLN(BLN43),.WL(WL205));
sram_cell_6t_5 inst_cell_205_44 (.BL(BL44),.BLN(BLN44),.WL(WL205));
sram_cell_6t_5 inst_cell_205_45 (.BL(BL45),.BLN(BLN45),.WL(WL205));
sram_cell_6t_5 inst_cell_205_46 (.BL(BL46),.BLN(BLN46),.WL(WL205));
sram_cell_6t_5 inst_cell_205_47 (.BL(BL47),.BLN(BLN47),.WL(WL205));
sram_cell_6t_5 inst_cell_205_48 (.BL(BL48),.BLN(BLN48),.WL(WL205));
sram_cell_6t_5 inst_cell_205_49 (.BL(BL49),.BLN(BLN49),.WL(WL205));
sram_cell_6t_5 inst_cell_205_50 (.BL(BL50),.BLN(BLN50),.WL(WL205));
sram_cell_6t_5 inst_cell_205_51 (.BL(BL51),.BLN(BLN51),.WL(WL205));
sram_cell_6t_5 inst_cell_205_52 (.BL(BL52),.BLN(BLN52),.WL(WL205));
sram_cell_6t_5 inst_cell_205_53 (.BL(BL53),.BLN(BLN53),.WL(WL205));
sram_cell_6t_5 inst_cell_205_54 (.BL(BL54),.BLN(BLN54),.WL(WL205));
sram_cell_6t_5 inst_cell_205_55 (.BL(BL55),.BLN(BLN55),.WL(WL205));
sram_cell_6t_5 inst_cell_205_56 (.BL(BL56),.BLN(BLN56),.WL(WL205));
sram_cell_6t_5 inst_cell_205_57 (.BL(BL57),.BLN(BLN57),.WL(WL205));
sram_cell_6t_5 inst_cell_205_58 (.BL(BL58),.BLN(BLN58),.WL(WL205));
sram_cell_6t_5 inst_cell_205_59 (.BL(BL59),.BLN(BLN59),.WL(WL205));
sram_cell_6t_5 inst_cell_205_60 (.BL(BL60),.BLN(BLN60),.WL(WL205));
sram_cell_6t_5 inst_cell_205_61 (.BL(BL61),.BLN(BLN61),.WL(WL205));
sram_cell_6t_5 inst_cell_205_62 (.BL(BL62),.BLN(BLN62),.WL(WL205));
sram_cell_6t_5 inst_cell_205_63 (.BL(BL63),.BLN(BLN63),.WL(WL205));
sram_cell_6t_5 inst_cell_205_64 (.BL(BL64),.BLN(BLN64),.WL(WL205));
sram_cell_6t_5 inst_cell_205_65 (.BL(BL65),.BLN(BLN65),.WL(WL205));
sram_cell_6t_5 inst_cell_205_66 (.BL(BL66),.BLN(BLN66),.WL(WL205));
sram_cell_6t_5 inst_cell_205_67 (.BL(BL67),.BLN(BLN67),.WL(WL205));
sram_cell_6t_5 inst_cell_205_68 (.BL(BL68),.BLN(BLN68),.WL(WL205));
sram_cell_6t_5 inst_cell_205_69 (.BL(BL69),.BLN(BLN69),.WL(WL205));
sram_cell_6t_5 inst_cell_205_70 (.BL(BL70),.BLN(BLN70),.WL(WL205));
sram_cell_6t_5 inst_cell_205_71 (.BL(BL71),.BLN(BLN71),.WL(WL205));
sram_cell_6t_5 inst_cell_205_72 (.BL(BL72),.BLN(BLN72),.WL(WL205));
sram_cell_6t_5 inst_cell_205_73 (.BL(BL73),.BLN(BLN73),.WL(WL205));
sram_cell_6t_5 inst_cell_205_74 (.BL(BL74),.BLN(BLN74),.WL(WL205));
sram_cell_6t_5 inst_cell_205_75 (.BL(BL75),.BLN(BLN75),.WL(WL205));
sram_cell_6t_5 inst_cell_205_76 (.BL(BL76),.BLN(BLN76),.WL(WL205));
sram_cell_6t_5 inst_cell_205_77 (.BL(BL77),.BLN(BLN77),.WL(WL205));
sram_cell_6t_5 inst_cell_205_78 (.BL(BL78),.BLN(BLN78),.WL(WL205));
sram_cell_6t_5 inst_cell_205_79 (.BL(BL79),.BLN(BLN79),.WL(WL205));
sram_cell_6t_5 inst_cell_205_80 (.BL(BL80),.BLN(BLN80),.WL(WL205));
sram_cell_6t_5 inst_cell_205_81 (.BL(BL81),.BLN(BLN81),.WL(WL205));
sram_cell_6t_5 inst_cell_205_82 (.BL(BL82),.BLN(BLN82),.WL(WL205));
sram_cell_6t_5 inst_cell_205_83 (.BL(BL83),.BLN(BLN83),.WL(WL205));
sram_cell_6t_5 inst_cell_205_84 (.BL(BL84),.BLN(BLN84),.WL(WL205));
sram_cell_6t_5 inst_cell_205_85 (.BL(BL85),.BLN(BLN85),.WL(WL205));
sram_cell_6t_5 inst_cell_205_86 (.BL(BL86),.BLN(BLN86),.WL(WL205));
sram_cell_6t_5 inst_cell_205_87 (.BL(BL87),.BLN(BLN87),.WL(WL205));
sram_cell_6t_5 inst_cell_205_88 (.BL(BL88),.BLN(BLN88),.WL(WL205));
sram_cell_6t_5 inst_cell_205_89 (.BL(BL89),.BLN(BLN89),.WL(WL205));
sram_cell_6t_5 inst_cell_205_90 (.BL(BL90),.BLN(BLN90),.WL(WL205));
sram_cell_6t_5 inst_cell_205_91 (.BL(BL91),.BLN(BLN91),.WL(WL205));
sram_cell_6t_5 inst_cell_205_92 (.BL(BL92),.BLN(BLN92),.WL(WL205));
sram_cell_6t_5 inst_cell_205_93 (.BL(BL93),.BLN(BLN93),.WL(WL205));
sram_cell_6t_5 inst_cell_205_94 (.BL(BL94),.BLN(BLN94),.WL(WL205));
sram_cell_6t_5 inst_cell_205_95 (.BL(BL95),.BLN(BLN95),.WL(WL205));
sram_cell_6t_5 inst_cell_205_96 (.BL(BL96),.BLN(BLN96),.WL(WL205));
sram_cell_6t_5 inst_cell_205_97 (.BL(BL97),.BLN(BLN97),.WL(WL205));
sram_cell_6t_5 inst_cell_205_98 (.BL(BL98),.BLN(BLN98),.WL(WL205));
sram_cell_6t_5 inst_cell_205_99 (.BL(BL99),.BLN(BLN99),.WL(WL205));
sram_cell_6t_5 inst_cell_205_100 (.BL(BL100),.BLN(BLN100),.WL(WL205));
sram_cell_6t_5 inst_cell_205_101 (.BL(BL101),.BLN(BLN101),.WL(WL205));
sram_cell_6t_5 inst_cell_205_102 (.BL(BL102),.BLN(BLN102),.WL(WL205));
sram_cell_6t_5 inst_cell_205_103 (.BL(BL103),.BLN(BLN103),.WL(WL205));
sram_cell_6t_5 inst_cell_205_104 (.BL(BL104),.BLN(BLN104),.WL(WL205));
sram_cell_6t_5 inst_cell_205_105 (.BL(BL105),.BLN(BLN105),.WL(WL205));
sram_cell_6t_5 inst_cell_205_106 (.BL(BL106),.BLN(BLN106),.WL(WL205));
sram_cell_6t_5 inst_cell_205_107 (.BL(BL107),.BLN(BLN107),.WL(WL205));
sram_cell_6t_5 inst_cell_205_108 (.BL(BL108),.BLN(BLN108),.WL(WL205));
sram_cell_6t_5 inst_cell_205_109 (.BL(BL109),.BLN(BLN109),.WL(WL205));
sram_cell_6t_5 inst_cell_205_110 (.BL(BL110),.BLN(BLN110),.WL(WL205));
sram_cell_6t_5 inst_cell_205_111 (.BL(BL111),.BLN(BLN111),.WL(WL205));
sram_cell_6t_5 inst_cell_205_112 (.BL(BL112),.BLN(BLN112),.WL(WL205));
sram_cell_6t_5 inst_cell_205_113 (.BL(BL113),.BLN(BLN113),.WL(WL205));
sram_cell_6t_5 inst_cell_205_114 (.BL(BL114),.BLN(BLN114),.WL(WL205));
sram_cell_6t_5 inst_cell_205_115 (.BL(BL115),.BLN(BLN115),.WL(WL205));
sram_cell_6t_5 inst_cell_205_116 (.BL(BL116),.BLN(BLN116),.WL(WL205));
sram_cell_6t_5 inst_cell_205_117 (.BL(BL117),.BLN(BLN117),.WL(WL205));
sram_cell_6t_5 inst_cell_205_118 (.BL(BL118),.BLN(BLN118),.WL(WL205));
sram_cell_6t_5 inst_cell_205_119 (.BL(BL119),.BLN(BLN119),.WL(WL205));
sram_cell_6t_5 inst_cell_205_120 (.BL(BL120),.BLN(BLN120),.WL(WL205));
sram_cell_6t_5 inst_cell_205_121 (.BL(BL121),.BLN(BLN121),.WL(WL205));
sram_cell_6t_5 inst_cell_205_122 (.BL(BL122),.BLN(BLN122),.WL(WL205));
sram_cell_6t_5 inst_cell_205_123 (.BL(BL123),.BLN(BLN123),.WL(WL205));
sram_cell_6t_5 inst_cell_205_124 (.BL(BL124),.BLN(BLN124),.WL(WL205));
sram_cell_6t_5 inst_cell_205_125 (.BL(BL125),.BLN(BLN125),.WL(WL205));
sram_cell_6t_5 inst_cell_205_126 (.BL(BL126),.BLN(BLN126),.WL(WL205));
sram_cell_6t_5 inst_cell_205_127 (.BL(BL127),.BLN(BLN127),.WL(WL205));
sram_cell_6t_5 inst_cell_206_0 (.BL(BL0),.BLN(BLN0),.WL(WL206));
sram_cell_6t_5 inst_cell_206_1 (.BL(BL1),.BLN(BLN1),.WL(WL206));
sram_cell_6t_5 inst_cell_206_2 (.BL(BL2),.BLN(BLN2),.WL(WL206));
sram_cell_6t_5 inst_cell_206_3 (.BL(BL3),.BLN(BLN3),.WL(WL206));
sram_cell_6t_5 inst_cell_206_4 (.BL(BL4),.BLN(BLN4),.WL(WL206));
sram_cell_6t_5 inst_cell_206_5 (.BL(BL5),.BLN(BLN5),.WL(WL206));
sram_cell_6t_5 inst_cell_206_6 (.BL(BL6),.BLN(BLN6),.WL(WL206));
sram_cell_6t_5 inst_cell_206_7 (.BL(BL7),.BLN(BLN7),.WL(WL206));
sram_cell_6t_5 inst_cell_206_8 (.BL(BL8),.BLN(BLN8),.WL(WL206));
sram_cell_6t_5 inst_cell_206_9 (.BL(BL9),.BLN(BLN9),.WL(WL206));
sram_cell_6t_5 inst_cell_206_10 (.BL(BL10),.BLN(BLN10),.WL(WL206));
sram_cell_6t_5 inst_cell_206_11 (.BL(BL11),.BLN(BLN11),.WL(WL206));
sram_cell_6t_5 inst_cell_206_12 (.BL(BL12),.BLN(BLN12),.WL(WL206));
sram_cell_6t_5 inst_cell_206_13 (.BL(BL13),.BLN(BLN13),.WL(WL206));
sram_cell_6t_5 inst_cell_206_14 (.BL(BL14),.BLN(BLN14),.WL(WL206));
sram_cell_6t_5 inst_cell_206_15 (.BL(BL15),.BLN(BLN15),.WL(WL206));
sram_cell_6t_5 inst_cell_206_16 (.BL(BL16),.BLN(BLN16),.WL(WL206));
sram_cell_6t_5 inst_cell_206_17 (.BL(BL17),.BLN(BLN17),.WL(WL206));
sram_cell_6t_5 inst_cell_206_18 (.BL(BL18),.BLN(BLN18),.WL(WL206));
sram_cell_6t_5 inst_cell_206_19 (.BL(BL19),.BLN(BLN19),.WL(WL206));
sram_cell_6t_5 inst_cell_206_20 (.BL(BL20),.BLN(BLN20),.WL(WL206));
sram_cell_6t_5 inst_cell_206_21 (.BL(BL21),.BLN(BLN21),.WL(WL206));
sram_cell_6t_5 inst_cell_206_22 (.BL(BL22),.BLN(BLN22),.WL(WL206));
sram_cell_6t_5 inst_cell_206_23 (.BL(BL23),.BLN(BLN23),.WL(WL206));
sram_cell_6t_5 inst_cell_206_24 (.BL(BL24),.BLN(BLN24),.WL(WL206));
sram_cell_6t_5 inst_cell_206_25 (.BL(BL25),.BLN(BLN25),.WL(WL206));
sram_cell_6t_5 inst_cell_206_26 (.BL(BL26),.BLN(BLN26),.WL(WL206));
sram_cell_6t_5 inst_cell_206_27 (.BL(BL27),.BLN(BLN27),.WL(WL206));
sram_cell_6t_5 inst_cell_206_28 (.BL(BL28),.BLN(BLN28),.WL(WL206));
sram_cell_6t_5 inst_cell_206_29 (.BL(BL29),.BLN(BLN29),.WL(WL206));
sram_cell_6t_5 inst_cell_206_30 (.BL(BL30),.BLN(BLN30),.WL(WL206));
sram_cell_6t_5 inst_cell_206_31 (.BL(BL31),.BLN(BLN31),.WL(WL206));
sram_cell_6t_5 inst_cell_206_32 (.BL(BL32),.BLN(BLN32),.WL(WL206));
sram_cell_6t_5 inst_cell_206_33 (.BL(BL33),.BLN(BLN33),.WL(WL206));
sram_cell_6t_5 inst_cell_206_34 (.BL(BL34),.BLN(BLN34),.WL(WL206));
sram_cell_6t_5 inst_cell_206_35 (.BL(BL35),.BLN(BLN35),.WL(WL206));
sram_cell_6t_5 inst_cell_206_36 (.BL(BL36),.BLN(BLN36),.WL(WL206));
sram_cell_6t_5 inst_cell_206_37 (.BL(BL37),.BLN(BLN37),.WL(WL206));
sram_cell_6t_5 inst_cell_206_38 (.BL(BL38),.BLN(BLN38),.WL(WL206));
sram_cell_6t_5 inst_cell_206_39 (.BL(BL39),.BLN(BLN39),.WL(WL206));
sram_cell_6t_5 inst_cell_206_40 (.BL(BL40),.BLN(BLN40),.WL(WL206));
sram_cell_6t_5 inst_cell_206_41 (.BL(BL41),.BLN(BLN41),.WL(WL206));
sram_cell_6t_5 inst_cell_206_42 (.BL(BL42),.BLN(BLN42),.WL(WL206));
sram_cell_6t_5 inst_cell_206_43 (.BL(BL43),.BLN(BLN43),.WL(WL206));
sram_cell_6t_5 inst_cell_206_44 (.BL(BL44),.BLN(BLN44),.WL(WL206));
sram_cell_6t_5 inst_cell_206_45 (.BL(BL45),.BLN(BLN45),.WL(WL206));
sram_cell_6t_5 inst_cell_206_46 (.BL(BL46),.BLN(BLN46),.WL(WL206));
sram_cell_6t_5 inst_cell_206_47 (.BL(BL47),.BLN(BLN47),.WL(WL206));
sram_cell_6t_5 inst_cell_206_48 (.BL(BL48),.BLN(BLN48),.WL(WL206));
sram_cell_6t_5 inst_cell_206_49 (.BL(BL49),.BLN(BLN49),.WL(WL206));
sram_cell_6t_5 inst_cell_206_50 (.BL(BL50),.BLN(BLN50),.WL(WL206));
sram_cell_6t_5 inst_cell_206_51 (.BL(BL51),.BLN(BLN51),.WL(WL206));
sram_cell_6t_5 inst_cell_206_52 (.BL(BL52),.BLN(BLN52),.WL(WL206));
sram_cell_6t_5 inst_cell_206_53 (.BL(BL53),.BLN(BLN53),.WL(WL206));
sram_cell_6t_5 inst_cell_206_54 (.BL(BL54),.BLN(BLN54),.WL(WL206));
sram_cell_6t_5 inst_cell_206_55 (.BL(BL55),.BLN(BLN55),.WL(WL206));
sram_cell_6t_5 inst_cell_206_56 (.BL(BL56),.BLN(BLN56),.WL(WL206));
sram_cell_6t_5 inst_cell_206_57 (.BL(BL57),.BLN(BLN57),.WL(WL206));
sram_cell_6t_5 inst_cell_206_58 (.BL(BL58),.BLN(BLN58),.WL(WL206));
sram_cell_6t_5 inst_cell_206_59 (.BL(BL59),.BLN(BLN59),.WL(WL206));
sram_cell_6t_5 inst_cell_206_60 (.BL(BL60),.BLN(BLN60),.WL(WL206));
sram_cell_6t_5 inst_cell_206_61 (.BL(BL61),.BLN(BLN61),.WL(WL206));
sram_cell_6t_5 inst_cell_206_62 (.BL(BL62),.BLN(BLN62),.WL(WL206));
sram_cell_6t_5 inst_cell_206_63 (.BL(BL63),.BLN(BLN63),.WL(WL206));
sram_cell_6t_5 inst_cell_206_64 (.BL(BL64),.BLN(BLN64),.WL(WL206));
sram_cell_6t_5 inst_cell_206_65 (.BL(BL65),.BLN(BLN65),.WL(WL206));
sram_cell_6t_5 inst_cell_206_66 (.BL(BL66),.BLN(BLN66),.WL(WL206));
sram_cell_6t_5 inst_cell_206_67 (.BL(BL67),.BLN(BLN67),.WL(WL206));
sram_cell_6t_5 inst_cell_206_68 (.BL(BL68),.BLN(BLN68),.WL(WL206));
sram_cell_6t_5 inst_cell_206_69 (.BL(BL69),.BLN(BLN69),.WL(WL206));
sram_cell_6t_5 inst_cell_206_70 (.BL(BL70),.BLN(BLN70),.WL(WL206));
sram_cell_6t_5 inst_cell_206_71 (.BL(BL71),.BLN(BLN71),.WL(WL206));
sram_cell_6t_5 inst_cell_206_72 (.BL(BL72),.BLN(BLN72),.WL(WL206));
sram_cell_6t_5 inst_cell_206_73 (.BL(BL73),.BLN(BLN73),.WL(WL206));
sram_cell_6t_5 inst_cell_206_74 (.BL(BL74),.BLN(BLN74),.WL(WL206));
sram_cell_6t_5 inst_cell_206_75 (.BL(BL75),.BLN(BLN75),.WL(WL206));
sram_cell_6t_5 inst_cell_206_76 (.BL(BL76),.BLN(BLN76),.WL(WL206));
sram_cell_6t_5 inst_cell_206_77 (.BL(BL77),.BLN(BLN77),.WL(WL206));
sram_cell_6t_5 inst_cell_206_78 (.BL(BL78),.BLN(BLN78),.WL(WL206));
sram_cell_6t_5 inst_cell_206_79 (.BL(BL79),.BLN(BLN79),.WL(WL206));
sram_cell_6t_5 inst_cell_206_80 (.BL(BL80),.BLN(BLN80),.WL(WL206));
sram_cell_6t_5 inst_cell_206_81 (.BL(BL81),.BLN(BLN81),.WL(WL206));
sram_cell_6t_5 inst_cell_206_82 (.BL(BL82),.BLN(BLN82),.WL(WL206));
sram_cell_6t_5 inst_cell_206_83 (.BL(BL83),.BLN(BLN83),.WL(WL206));
sram_cell_6t_5 inst_cell_206_84 (.BL(BL84),.BLN(BLN84),.WL(WL206));
sram_cell_6t_5 inst_cell_206_85 (.BL(BL85),.BLN(BLN85),.WL(WL206));
sram_cell_6t_5 inst_cell_206_86 (.BL(BL86),.BLN(BLN86),.WL(WL206));
sram_cell_6t_5 inst_cell_206_87 (.BL(BL87),.BLN(BLN87),.WL(WL206));
sram_cell_6t_5 inst_cell_206_88 (.BL(BL88),.BLN(BLN88),.WL(WL206));
sram_cell_6t_5 inst_cell_206_89 (.BL(BL89),.BLN(BLN89),.WL(WL206));
sram_cell_6t_5 inst_cell_206_90 (.BL(BL90),.BLN(BLN90),.WL(WL206));
sram_cell_6t_5 inst_cell_206_91 (.BL(BL91),.BLN(BLN91),.WL(WL206));
sram_cell_6t_5 inst_cell_206_92 (.BL(BL92),.BLN(BLN92),.WL(WL206));
sram_cell_6t_5 inst_cell_206_93 (.BL(BL93),.BLN(BLN93),.WL(WL206));
sram_cell_6t_5 inst_cell_206_94 (.BL(BL94),.BLN(BLN94),.WL(WL206));
sram_cell_6t_5 inst_cell_206_95 (.BL(BL95),.BLN(BLN95),.WL(WL206));
sram_cell_6t_5 inst_cell_206_96 (.BL(BL96),.BLN(BLN96),.WL(WL206));
sram_cell_6t_5 inst_cell_206_97 (.BL(BL97),.BLN(BLN97),.WL(WL206));
sram_cell_6t_5 inst_cell_206_98 (.BL(BL98),.BLN(BLN98),.WL(WL206));
sram_cell_6t_5 inst_cell_206_99 (.BL(BL99),.BLN(BLN99),.WL(WL206));
sram_cell_6t_5 inst_cell_206_100 (.BL(BL100),.BLN(BLN100),.WL(WL206));
sram_cell_6t_5 inst_cell_206_101 (.BL(BL101),.BLN(BLN101),.WL(WL206));
sram_cell_6t_5 inst_cell_206_102 (.BL(BL102),.BLN(BLN102),.WL(WL206));
sram_cell_6t_5 inst_cell_206_103 (.BL(BL103),.BLN(BLN103),.WL(WL206));
sram_cell_6t_5 inst_cell_206_104 (.BL(BL104),.BLN(BLN104),.WL(WL206));
sram_cell_6t_5 inst_cell_206_105 (.BL(BL105),.BLN(BLN105),.WL(WL206));
sram_cell_6t_5 inst_cell_206_106 (.BL(BL106),.BLN(BLN106),.WL(WL206));
sram_cell_6t_5 inst_cell_206_107 (.BL(BL107),.BLN(BLN107),.WL(WL206));
sram_cell_6t_5 inst_cell_206_108 (.BL(BL108),.BLN(BLN108),.WL(WL206));
sram_cell_6t_5 inst_cell_206_109 (.BL(BL109),.BLN(BLN109),.WL(WL206));
sram_cell_6t_5 inst_cell_206_110 (.BL(BL110),.BLN(BLN110),.WL(WL206));
sram_cell_6t_5 inst_cell_206_111 (.BL(BL111),.BLN(BLN111),.WL(WL206));
sram_cell_6t_5 inst_cell_206_112 (.BL(BL112),.BLN(BLN112),.WL(WL206));
sram_cell_6t_5 inst_cell_206_113 (.BL(BL113),.BLN(BLN113),.WL(WL206));
sram_cell_6t_5 inst_cell_206_114 (.BL(BL114),.BLN(BLN114),.WL(WL206));
sram_cell_6t_5 inst_cell_206_115 (.BL(BL115),.BLN(BLN115),.WL(WL206));
sram_cell_6t_5 inst_cell_206_116 (.BL(BL116),.BLN(BLN116),.WL(WL206));
sram_cell_6t_5 inst_cell_206_117 (.BL(BL117),.BLN(BLN117),.WL(WL206));
sram_cell_6t_5 inst_cell_206_118 (.BL(BL118),.BLN(BLN118),.WL(WL206));
sram_cell_6t_5 inst_cell_206_119 (.BL(BL119),.BLN(BLN119),.WL(WL206));
sram_cell_6t_5 inst_cell_206_120 (.BL(BL120),.BLN(BLN120),.WL(WL206));
sram_cell_6t_5 inst_cell_206_121 (.BL(BL121),.BLN(BLN121),.WL(WL206));
sram_cell_6t_5 inst_cell_206_122 (.BL(BL122),.BLN(BLN122),.WL(WL206));
sram_cell_6t_5 inst_cell_206_123 (.BL(BL123),.BLN(BLN123),.WL(WL206));
sram_cell_6t_5 inst_cell_206_124 (.BL(BL124),.BLN(BLN124),.WL(WL206));
sram_cell_6t_5 inst_cell_206_125 (.BL(BL125),.BLN(BLN125),.WL(WL206));
sram_cell_6t_5 inst_cell_206_126 (.BL(BL126),.BLN(BLN126),.WL(WL206));
sram_cell_6t_5 inst_cell_206_127 (.BL(BL127),.BLN(BLN127),.WL(WL206));
sram_cell_6t_5 inst_cell_207_0 (.BL(BL0),.BLN(BLN0),.WL(WL207));
sram_cell_6t_5 inst_cell_207_1 (.BL(BL1),.BLN(BLN1),.WL(WL207));
sram_cell_6t_5 inst_cell_207_2 (.BL(BL2),.BLN(BLN2),.WL(WL207));
sram_cell_6t_5 inst_cell_207_3 (.BL(BL3),.BLN(BLN3),.WL(WL207));
sram_cell_6t_5 inst_cell_207_4 (.BL(BL4),.BLN(BLN4),.WL(WL207));
sram_cell_6t_5 inst_cell_207_5 (.BL(BL5),.BLN(BLN5),.WL(WL207));
sram_cell_6t_5 inst_cell_207_6 (.BL(BL6),.BLN(BLN6),.WL(WL207));
sram_cell_6t_5 inst_cell_207_7 (.BL(BL7),.BLN(BLN7),.WL(WL207));
sram_cell_6t_5 inst_cell_207_8 (.BL(BL8),.BLN(BLN8),.WL(WL207));
sram_cell_6t_5 inst_cell_207_9 (.BL(BL9),.BLN(BLN9),.WL(WL207));
sram_cell_6t_5 inst_cell_207_10 (.BL(BL10),.BLN(BLN10),.WL(WL207));
sram_cell_6t_5 inst_cell_207_11 (.BL(BL11),.BLN(BLN11),.WL(WL207));
sram_cell_6t_5 inst_cell_207_12 (.BL(BL12),.BLN(BLN12),.WL(WL207));
sram_cell_6t_5 inst_cell_207_13 (.BL(BL13),.BLN(BLN13),.WL(WL207));
sram_cell_6t_5 inst_cell_207_14 (.BL(BL14),.BLN(BLN14),.WL(WL207));
sram_cell_6t_5 inst_cell_207_15 (.BL(BL15),.BLN(BLN15),.WL(WL207));
sram_cell_6t_5 inst_cell_207_16 (.BL(BL16),.BLN(BLN16),.WL(WL207));
sram_cell_6t_5 inst_cell_207_17 (.BL(BL17),.BLN(BLN17),.WL(WL207));
sram_cell_6t_5 inst_cell_207_18 (.BL(BL18),.BLN(BLN18),.WL(WL207));
sram_cell_6t_5 inst_cell_207_19 (.BL(BL19),.BLN(BLN19),.WL(WL207));
sram_cell_6t_5 inst_cell_207_20 (.BL(BL20),.BLN(BLN20),.WL(WL207));
sram_cell_6t_5 inst_cell_207_21 (.BL(BL21),.BLN(BLN21),.WL(WL207));
sram_cell_6t_5 inst_cell_207_22 (.BL(BL22),.BLN(BLN22),.WL(WL207));
sram_cell_6t_5 inst_cell_207_23 (.BL(BL23),.BLN(BLN23),.WL(WL207));
sram_cell_6t_5 inst_cell_207_24 (.BL(BL24),.BLN(BLN24),.WL(WL207));
sram_cell_6t_5 inst_cell_207_25 (.BL(BL25),.BLN(BLN25),.WL(WL207));
sram_cell_6t_5 inst_cell_207_26 (.BL(BL26),.BLN(BLN26),.WL(WL207));
sram_cell_6t_5 inst_cell_207_27 (.BL(BL27),.BLN(BLN27),.WL(WL207));
sram_cell_6t_5 inst_cell_207_28 (.BL(BL28),.BLN(BLN28),.WL(WL207));
sram_cell_6t_5 inst_cell_207_29 (.BL(BL29),.BLN(BLN29),.WL(WL207));
sram_cell_6t_5 inst_cell_207_30 (.BL(BL30),.BLN(BLN30),.WL(WL207));
sram_cell_6t_5 inst_cell_207_31 (.BL(BL31),.BLN(BLN31),.WL(WL207));
sram_cell_6t_5 inst_cell_207_32 (.BL(BL32),.BLN(BLN32),.WL(WL207));
sram_cell_6t_5 inst_cell_207_33 (.BL(BL33),.BLN(BLN33),.WL(WL207));
sram_cell_6t_5 inst_cell_207_34 (.BL(BL34),.BLN(BLN34),.WL(WL207));
sram_cell_6t_5 inst_cell_207_35 (.BL(BL35),.BLN(BLN35),.WL(WL207));
sram_cell_6t_5 inst_cell_207_36 (.BL(BL36),.BLN(BLN36),.WL(WL207));
sram_cell_6t_5 inst_cell_207_37 (.BL(BL37),.BLN(BLN37),.WL(WL207));
sram_cell_6t_5 inst_cell_207_38 (.BL(BL38),.BLN(BLN38),.WL(WL207));
sram_cell_6t_5 inst_cell_207_39 (.BL(BL39),.BLN(BLN39),.WL(WL207));
sram_cell_6t_5 inst_cell_207_40 (.BL(BL40),.BLN(BLN40),.WL(WL207));
sram_cell_6t_5 inst_cell_207_41 (.BL(BL41),.BLN(BLN41),.WL(WL207));
sram_cell_6t_5 inst_cell_207_42 (.BL(BL42),.BLN(BLN42),.WL(WL207));
sram_cell_6t_5 inst_cell_207_43 (.BL(BL43),.BLN(BLN43),.WL(WL207));
sram_cell_6t_5 inst_cell_207_44 (.BL(BL44),.BLN(BLN44),.WL(WL207));
sram_cell_6t_5 inst_cell_207_45 (.BL(BL45),.BLN(BLN45),.WL(WL207));
sram_cell_6t_5 inst_cell_207_46 (.BL(BL46),.BLN(BLN46),.WL(WL207));
sram_cell_6t_5 inst_cell_207_47 (.BL(BL47),.BLN(BLN47),.WL(WL207));
sram_cell_6t_5 inst_cell_207_48 (.BL(BL48),.BLN(BLN48),.WL(WL207));
sram_cell_6t_5 inst_cell_207_49 (.BL(BL49),.BLN(BLN49),.WL(WL207));
sram_cell_6t_5 inst_cell_207_50 (.BL(BL50),.BLN(BLN50),.WL(WL207));
sram_cell_6t_5 inst_cell_207_51 (.BL(BL51),.BLN(BLN51),.WL(WL207));
sram_cell_6t_5 inst_cell_207_52 (.BL(BL52),.BLN(BLN52),.WL(WL207));
sram_cell_6t_5 inst_cell_207_53 (.BL(BL53),.BLN(BLN53),.WL(WL207));
sram_cell_6t_5 inst_cell_207_54 (.BL(BL54),.BLN(BLN54),.WL(WL207));
sram_cell_6t_5 inst_cell_207_55 (.BL(BL55),.BLN(BLN55),.WL(WL207));
sram_cell_6t_5 inst_cell_207_56 (.BL(BL56),.BLN(BLN56),.WL(WL207));
sram_cell_6t_5 inst_cell_207_57 (.BL(BL57),.BLN(BLN57),.WL(WL207));
sram_cell_6t_5 inst_cell_207_58 (.BL(BL58),.BLN(BLN58),.WL(WL207));
sram_cell_6t_5 inst_cell_207_59 (.BL(BL59),.BLN(BLN59),.WL(WL207));
sram_cell_6t_5 inst_cell_207_60 (.BL(BL60),.BLN(BLN60),.WL(WL207));
sram_cell_6t_5 inst_cell_207_61 (.BL(BL61),.BLN(BLN61),.WL(WL207));
sram_cell_6t_5 inst_cell_207_62 (.BL(BL62),.BLN(BLN62),.WL(WL207));
sram_cell_6t_5 inst_cell_207_63 (.BL(BL63),.BLN(BLN63),.WL(WL207));
sram_cell_6t_5 inst_cell_207_64 (.BL(BL64),.BLN(BLN64),.WL(WL207));
sram_cell_6t_5 inst_cell_207_65 (.BL(BL65),.BLN(BLN65),.WL(WL207));
sram_cell_6t_5 inst_cell_207_66 (.BL(BL66),.BLN(BLN66),.WL(WL207));
sram_cell_6t_5 inst_cell_207_67 (.BL(BL67),.BLN(BLN67),.WL(WL207));
sram_cell_6t_5 inst_cell_207_68 (.BL(BL68),.BLN(BLN68),.WL(WL207));
sram_cell_6t_5 inst_cell_207_69 (.BL(BL69),.BLN(BLN69),.WL(WL207));
sram_cell_6t_5 inst_cell_207_70 (.BL(BL70),.BLN(BLN70),.WL(WL207));
sram_cell_6t_5 inst_cell_207_71 (.BL(BL71),.BLN(BLN71),.WL(WL207));
sram_cell_6t_5 inst_cell_207_72 (.BL(BL72),.BLN(BLN72),.WL(WL207));
sram_cell_6t_5 inst_cell_207_73 (.BL(BL73),.BLN(BLN73),.WL(WL207));
sram_cell_6t_5 inst_cell_207_74 (.BL(BL74),.BLN(BLN74),.WL(WL207));
sram_cell_6t_5 inst_cell_207_75 (.BL(BL75),.BLN(BLN75),.WL(WL207));
sram_cell_6t_5 inst_cell_207_76 (.BL(BL76),.BLN(BLN76),.WL(WL207));
sram_cell_6t_5 inst_cell_207_77 (.BL(BL77),.BLN(BLN77),.WL(WL207));
sram_cell_6t_5 inst_cell_207_78 (.BL(BL78),.BLN(BLN78),.WL(WL207));
sram_cell_6t_5 inst_cell_207_79 (.BL(BL79),.BLN(BLN79),.WL(WL207));
sram_cell_6t_5 inst_cell_207_80 (.BL(BL80),.BLN(BLN80),.WL(WL207));
sram_cell_6t_5 inst_cell_207_81 (.BL(BL81),.BLN(BLN81),.WL(WL207));
sram_cell_6t_5 inst_cell_207_82 (.BL(BL82),.BLN(BLN82),.WL(WL207));
sram_cell_6t_5 inst_cell_207_83 (.BL(BL83),.BLN(BLN83),.WL(WL207));
sram_cell_6t_5 inst_cell_207_84 (.BL(BL84),.BLN(BLN84),.WL(WL207));
sram_cell_6t_5 inst_cell_207_85 (.BL(BL85),.BLN(BLN85),.WL(WL207));
sram_cell_6t_5 inst_cell_207_86 (.BL(BL86),.BLN(BLN86),.WL(WL207));
sram_cell_6t_5 inst_cell_207_87 (.BL(BL87),.BLN(BLN87),.WL(WL207));
sram_cell_6t_5 inst_cell_207_88 (.BL(BL88),.BLN(BLN88),.WL(WL207));
sram_cell_6t_5 inst_cell_207_89 (.BL(BL89),.BLN(BLN89),.WL(WL207));
sram_cell_6t_5 inst_cell_207_90 (.BL(BL90),.BLN(BLN90),.WL(WL207));
sram_cell_6t_5 inst_cell_207_91 (.BL(BL91),.BLN(BLN91),.WL(WL207));
sram_cell_6t_5 inst_cell_207_92 (.BL(BL92),.BLN(BLN92),.WL(WL207));
sram_cell_6t_5 inst_cell_207_93 (.BL(BL93),.BLN(BLN93),.WL(WL207));
sram_cell_6t_5 inst_cell_207_94 (.BL(BL94),.BLN(BLN94),.WL(WL207));
sram_cell_6t_5 inst_cell_207_95 (.BL(BL95),.BLN(BLN95),.WL(WL207));
sram_cell_6t_5 inst_cell_207_96 (.BL(BL96),.BLN(BLN96),.WL(WL207));
sram_cell_6t_5 inst_cell_207_97 (.BL(BL97),.BLN(BLN97),.WL(WL207));
sram_cell_6t_5 inst_cell_207_98 (.BL(BL98),.BLN(BLN98),.WL(WL207));
sram_cell_6t_5 inst_cell_207_99 (.BL(BL99),.BLN(BLN99),.WL(WL207));
sram_cell_6t_5 inst_cell_207_100 (.BL(BL100),.BLN(BLN100),.WL(WL207));
sram_cell_6t_5 inst_cell_207_101 (.BL(BL101),.BLN(BLN101),.WL(WL207));
sram_cell_6t_5 inst_cell_207_102 (.BL(BL102),.BLN(BLN102),.WL(WL207));
sram_cell_6t_5 inst_cell_207_103 (.BL(BL103),.BLN(BLN103),.WL(WL207));
sram_cell_6t_5 inst_cell_207_104 (.BL(BL104),.BLN(BLN104),.WL(WL207));
sram_cell_6t_5 inst_cell_207_105 (.BL(BL105),.BLN(BLN105),.WL(WL207));
sram_cell_6t_5 inst_cell_207_106 (.BL(BL106),.BLN(BLN106),.WL(WL207));
sram_cell_6t_5 inst_cell_207_107 (.BL(BL107),.BLN(BLN107),.WL(WL207));
sram_cell_6t_5 inst_cell_207_108 (.BL(BL108),.BLN(BLN108),.WL(WL207));
sram_cell_6t_5 inst_cell_207_109 (.BL(BL109),.BLN(BLN109),.WL(WL207));
sram_cell_6t_5 inst_cell_207_110 (.BL(BL110),.BLN(BLN110),.WL(WL207));
sram_cell_6t_5 inst_cell_207_111 (.BL(BL111),.BLN(BLN111),.WL(WL207));
sram_cell_6t_5 inst_cell_207_112 (.BL(BL112),.BLN(BLN112),.WL(WL207));
sram_cell_6t_5 inst_cell_207_113 (.BL(BL113),.BLN(BLN113),.WL(WL207));
sram_cell_6t_5 inst_cell_207_114 (.BL(BL114),.BLN(BLN114),.WL(WL207));
sram_cell_6t_5 inst_cell_207_115 (.BL(BL115),.BLN(BLN115),.WL(WL207));
sram_cell_6t_5 inst_cell_207_116 (.BL(BL116),.BLN(BLN116),.WL(WL207));
sram_cell_6t_5 inst_cell_207_117 (.BL(BL117),.BLN(BLN117),.WL(WL207));
sram_cell_6t_5 inst_cell_207_118 (.BL(BL118),.BLN(BLN118),.WL(WL207));
sram_cell_6t_5 inst_cell_207_119 (.BL(BL119),.BLN(BLN119),.WL(WL207));
sram_cell_6t_5 inst_cell_207_120 (.BL(BL120),.BLN(BLN120),.WL(WL207));
sram_cell_6t_5 inst_cell_207_121 (.BL(BL121),.BLN(BLN121),.WL(WL207));
sram_cell_6t_5 inst_cell_207_122 (.BL(BL122),.BLN(BLN122),.WL(WL207));
sram_cell_6t_5 inst_cell_207_123 (.BL(BL123),.BLN(BLN123),.WL(WL207));
sram_cell_6t_5 inst_cell_207_124 (.BL(BL124),.BLN(BLN124),.WL(WL207));
sram_cell_6t_5 inst_cell_207_125 (.BL(BL125),.BLN(BLN125),.WL(WL207));
sram_cell_6t_5 inst_cell_207_126 (.BL(BL126),.BLN(BLN126),.WL(WL207));
sram_cell_6t_5 inst_cell_207_127 (.BL(BL127),.BLN(BLN127),.WL(WL207));
sram_cell_6t_5 inst_cell_208_0 (.BL(BL0),.BLN(BLN0),.WL(WL208));
sram_cell_6t_5 inst_cell_208_1 (.BL(BL1),.BLN(BLN1),.WL(WL208));
sram_cell_6t_5 inst_cell_208_2 (.BL(BL2),.BLN(BLN2),.WL(WL208));
sram_cell_6t_5 inst_cell_208_3 (.BL(BL3),.BLN(BLN3),.WL(WL208));
sram_cell_6t_5 inst_cell_208_4 (.BL(BL4),.BLN(BLN4),.WL(WL208));
sram_cell_6t_5 inst_cell_208_5 (.BL(BL5),.BLN(BLN5),.WL(WL208));
sram_cell_6t_5 inst_cell_208_6 (.BL(BL6),.BLN(BLN6),.WL(WL208));
sram_cell_6t_5 inst_cell_208_7 (.BL(BL7),.BLN(BLN7),.WL(WL208));
sram_cell_6t_5 inst_cell_208_8 (.BL(BL8),.BLN(BLN8),.WL(WL208));
sram_cell_6t_5 inst_cell_208_9 (.BL(BL9),.BLN(BLN9),.WL(WL208));
sram_cell_6t_5 inst_cell_208_10 (.BL(BL10),.BLN(BLN10),.WL(WL208));
sram_cell_6t_5 inst_cell_208_11 (.BL(BL11),.BLN(BLN11),.WL(WL208));
sram_cell_6t_5 inst_cell_208_12 (.BL(BL12),.BLN(BLN12),.WL(WL208));
sram_cell_6t_5 inst_cell_208_13 (.BL(BL13),.BLN(BLN13),.WL(WL208));
sram_cell_6t_5 inst_cell_208_14 (.BL(BL14),.BLN(BLN14),.WL(WL208));
sram_cell_6t_5 inst_cell_208_15 (.BL(BL15),.BLN(BLN15),.WL(WL208));
sram_cell_6t_5 inst_cell_208_16 (.BL(BL16),.BLN(BLN16),.WL(WL208));
sram_cell_6t_5 inst_cell_208_17 (.BL(BL17),.BLN(BLN17),.WL(WL208));
sram_cell_6t_5 inst_cell_208_18 (.BL(BL18),.BLN(BLN18),.WL(WL208));
sram_cell_6t_5 inst_cell_208_19 (.BL(BL19),.BLN(BLN19),.WL(WL208));
sram_cell_6t_5 inst_cell_208_20 (.BL(BL20),.BLN(BLN20),.WL(WL208));
sram_cell_6t_5 inst_cell_208_21 (.BL(BL21),.BLN(BLN21),.WL(WL208));
sram_cell_6t_5 inst_cell_208_22 (.BL(BL22),.BLN(BLN22),.WL(WL208));
sram_cell_6t_5 inst_cell_208_23 (.BL(BL23),.BLN(BLN23),.WL(WL208));
sram_cell_6t_5 inst_cell_208_24 (.BL(BL24),.BLN(BLN24),.WL(WL208));
sram_cell_6t_5 inst_cell_208_25 (.BL(BL25),.BLN(BLN25),.WL(WL208));
sram_cell_6t_5 inst_cell_208_26 (.BL(BL26),.BLN(BLN26),.WL(WL208));
sram_cell_6t_5 inst_cell_208_27 (.BL(BL27),.BLN(BLN27),.WL(WL208));
sram_cell_6t_5 inst_cell_208_28 (.BL(BL28),.BLN(BLN28),.WL(WL208));
sram_cell_6t_5 inst_cell_208_29 (.BL(BL29),.BLN(BLN29),.WL(WL208));
sram_cell_6t_5 inst_cell_208_30 (.BL(BL30),.BLN(BLN30),.WL(WL208));
sram_cell_6t_5 inst_cell_208_31 (.BL(BL31),.BLN(BLN31),.WL(WL208));
sram_cell_6t_5 inst_cell_208_32 (.BL(BL32),.BLN(BLN32),.WL(WL208));
sram_cell_6t_5 inst_cell_208_33 (.BL(BL33),.BLN(BLN33),.WL(WL208));
sram_cell_6t_5 inst_cell_208_34 (.BL(BL34),.BLN(BLN34),.WL(WL208));
sram_cell_6t_5 inst_cell_208_35 (.BL(BL35),.BLN(BLN35),.WL(WL208));
sram_cell_6t_5 inst_cell_208_36 (.BL(BL36),.BLN(BLN36),.WL(WL208));
sram_cell_6t_5 inst_cell_208_37 (.BL(BL37),.BLN(BLN37),.WL(WL208));
sram_cell_6t_5 inst_cell_208_38 (.BL(BL38),.BLN(BLN38),.WL(WL208));
sram_cell_6t_5 inst_cell_208_39 (.BL(BL39),.BLN(BLN39),.WL(WL208));
sram_cell_6t_5 inst_cell_208_40 (.BL(BL40),.BLN(BLN40),.WL(WL208));
sram_cell_6t_5 inst_cell_208_41 (.BL(BL41),.BLN(BLN41),.WL(WL208));
sram_cell_6t_5 inst_cell_208_42 (.BL(BL42),.BLN(BLN42),.WL(WL208));
sram_cell_6t_5 inst_cell_208_43 (.BL(BL43),.BLN(BLN43),.WL(WL208));
sram_cell_6t_5 inst_cell_208_44 (.BL(BL44),.BLN(BLN44),.WL(WL208));
sram_cell_6t_5 inst_cell_208_45 (.BL(BL45),.BLN(BLN45),.WL(WL208));
sram_cell_6t_5 inst_cell_208_46 (.BL(BL46),.BLN(BLN46),.WL(WL208));
sram_cell_6t_5 inst_cell_208_47 (.BL(BL47),.BLN(BLN47),.WL(WL208));
sram_cell_6t_5 inst_cell_208_48 (.BL(BL48),.BLN(BLN48),.WL(WL208));
sram_cell_6t_5 inst_cell_208_49 (.BL(BL49),.BLN(BLN49),.WL(WL208));
sram_cell_6t_5 inst_cell_208_50 (.BL(BL50),.BLN(BLN50),.WL(WL208));
sram_cell_6t_5 inst_cell_208_51 (.BL(BL51),.BLN(BLN51),.WL(WL208));
sram_cell_6t_5 inst_cell_208_52 (.BL(BL52),.BLN(BLN52),.WL(WL208));
sram_cell_6t_5 inst_cell_208_53 (.BL(BL53),.BLN(BLN53),.WL(WL208));
sram_cell_6t_5 inst_cell_208_54 (.BL(BL54),.BLN(BLN54),.WL(WL208));
sram_cell_6t_5 inst_cell_208_55 (.BL(BL55),.BLN(BLN55),.WL(WL208));
sram_cell_6t_5 inst_cell_208_56 (.BL(BL56),.BLN(BLN56),.WL(WL208));
sram_cell_6t_5 inst_cell_208_57 (.BL(BL57),.BLN(BLN57),.WL(WL208));
sram_cell_6t_5 inst_cell_208_58 (.BL(BL58),.BLN(BLN58),.WL(WL208));
sram_cell_6t_5 inst_cell_208_59 (.BL(BL59),.BLN(BLN59),.WL(WL208));
sram_cell_6t_5 inst_cell_208_60 (.BL(BL60),.BLN(BLN60),.WL(WL208));
sram_cell_6t_5 inst_cell_208_61 (.BL(BL61),.BLN(BLN61),.WL(WL208));
sram_cell_6t_5 inst_cell_208_62 (.BL(BL62),.BLN(BLN62),.WL(WL208));
sram_cell_6t_5 inst_cell_208_63 (.BL(BL63),.BLN(BLN63),.WL(WL208));
sram_cell_6t_5 inst_cell_208_64 (.BL(BL64),.BLN(BLN64),.WL(WL208));
sram_cell_6t_5 inst_cell_208_65 (.BL(BL65),.BLN(BLN65),.WL(WL208));
sram_cell_6t_5 inst_cell_208_66 (.BL(BL66),.BLN(BLN66),.WL(WL208));
sram_cell_6t_5 inst_cell_208_67 (.BL(BL67),.BLN(BLN67),.WL(WL208));
sram_cell_6t_5 inst_cell_208_68 (.BL(BL68),.BLN(BLN68),.WL(WL208));
sram_cell_6t_5 inst_cell_208_69 (.BL(BL69),.BLN(BLN69),.WL(WL208));
sram_cell_6t_5 inst_cell_208_70 (.BL(BL70),.BLN(BLN70),.WL(WL208));
sram_cell_6t_5 inst_cell_208_71 (.BL(BL71),.BLN(BLN71),.WL(WL208));
sram_cell_6t_5 inst_cell_208_72 (.BL(BL72),.BLN(BLN72),.WL(WL208));
sram_cell_6t_5 inst_cell_208_73 (.BL(BL73),.BLN(BLN73),.WL(WL208));
sram_cell_6t_5 inst_cell_208_74 (.BL(BL74),.BLN(BLN74),.WL(WL208));
sram_cell_6t_5 inst_cell_208_75 (.BL(BL75),.BLN(BLN75),.WL(WL208));
sram_cell_6t_5 inst_cell_208_76 (.BL(BL76),.BLN(BLN76),.WL(WL208));
sram_cell_6t_5 inst_cell_208_77 (.BL(BL77),.BLN(BLN77),.WL(WL208));
sram_cell_6t_5 inst_cell_208_78 (.BL(BL78),.BLN(BLN78),.WL(WL208));
sram_cell_6t_5 inst_cell_208_79 (.BL(BL79),.BLN(BLN79),.WL(WL208));
sram_cell_6t_5 inst_cell_208_80 (.BL(BL80),.BLN(BLN80),.WL(WL208));
sram_cell_6t_5 inst_cell_208_81 (.BL(BL81),.BLN(BLN81),.WL(WL208));
sram_cell_6t_5 inst_cell_208_82 (.BL(BL82),.BLN(BLN82),.WL(WL208));
sram_cell_6t_5 inst_cell_208_83 (.BL(BL83),.BLN(BLN83),.WL(WL208));
sram_cell_6t_5 inst_cell_208_84 (.BL(BL84),.BLN(BLN84),.WL(WL208));
sram_cell_6t_5 inst_cell_208_85 (.BL(BL85),.BLN(BLN85),.WL(WL208));
sram_cell_6t_5 inst_cell_208_86 (.BL(BL86),.BLN(BLN86),.WL(WL208));
sram_cell_6t_5 inst_cell_208_87 (.BL(BL87),.BLN(BLN87),.WL(WL208));
sram_cell_6t_5 inst_cell_208_88 (.BL(BL88),.BLN(BLN88),.WL(WL208));
sram_cell_6t_5 inst_cell_208_89 (.BL(BL89),.BLN(BLN89),.WL(WL208));
sram_cell_6t_5 inst_cell_208_90 (.BL(BL90),.BLN(BLN90),.WL(WL208));
sram_cell_6t_5 inst_cell_208_91 (.BL(BL91),.BLN(BLN91),.WL(WL208));
sram_cell_6t_5 inst_cell_208_92 (.BL(BL92),.BLN(BLN92),.WL(WL208));
sram_cell_6t_5 inst_cell_208_93 (.BL(BL93),.BLN(BLN93),.WL(WL208));
sram_cell_6t_5 inst_cell_208_94 (.BL(BL94),.BLN(BLN94),.WL(WL208));
sram_cell_6t_5 inst_cell_208_95 (.BL(BL95),.BLN(BLN95),.WL(WL208));
sram_cell_6t_5 inst_cell_208_96 (.BL(BL96),.BLN(BLN96),.WL(WL208));
sram_cell_6t_5 inst_cell_208_97 (.BL(BL97),.BLN(BLN97),.WL(WL208));
sram_cell_6t_5 inst_cell_208_98 (.BL(BL98),.BLN(BLN98),.WL(WL208));
sram_cell_6t_5 inst_cell_208_99 (.BL(BL99),.BLN(BLN99),.WL(WL208));
sram_cell_6t_5 inst_cell_208_100 (.BL(BL100),.BLN(BLN100),.WL(WL208));
sram_cell_6t_5 inst_cell_208_101 (.BL(BL101),.BLN(BLN101),.WL(WL208));
sram_cell_6t_5 inst_cell_208_102 (.BL(BL102),.BLN(BLN102),.WL(WL208));
sram_cell_6t_5 inst_cell_208_103 (.BL(BL103),.BLN(BLN103),.WL(WL208));
sram_cell_6t_5 inst_cell_208_104 (.BL(BL104),.BLN(BLN104),.WL(WL208));
sram_cell_6t_5 inst_cell_208_105 (.BL(BL105),.BLN(BLN105),.WL(WL208));
sram_cell_6t_5 inst_cell_208_106 (.BL(BL106),.BLN(BLN106),.WL(WL208));
sram_cell_6t_5 inst_cell_208_107 (.BL(BL107),.BLN(BLN107),.WL(WL208));
sram_cell_6t_5 inst_cell_208_108 (.BL(BL108),.BLN(BLN108),.WL(WL208));
sram_cell_6t_5 inst_cell_208_109 (.BL(BL109),.BLN(BLN109),.WL(WL208));
sram_cell_6t_5 inst_cell_208_110 (.BL(BL110),.BLN(BLN110),.WL(WL208));
sram_cell_6t_5 inst_cell_208_111 (.BL(BL111),.BLN(BLN111),.WL(WL208));
sram_cell_6t_5 inst_cell_208_112 (.BL(BL112),.BLN(BLN112),.WL(WL208));
sram_cell_6t_5 inst_cell_208_113 (.BL(BL113),.BLN(BLN113),.WL(WL208));
sram_cell_6t_5 inst_cell_208_114 (.BL(BL114),.BLN(BLN114),.WL(WL208));
sram_cell_6t_5 inst_cell_208_115 (.BL(BL115),.BLN(BLN115),.WL(WL208));
sram_cell_6t_5 inst_cell_208_116 (.BL(BL116),.BLN(BLN116),.WL(WL208));
sram_cell_6t_5 inst_cell_208_117 (.BL(BL117),.BLN(BLN117),.WL(WL208));
sram_cell_6t_5 inst_cell_208_118 (.BL(BL118),.BLN(BLN118),.WL(WL208));
sram_cell_6t_5 inst_cell_208_119 (.BL(BL119),.BLN(BLN119),.WL(WL208));
sram_cell_6t_5 inst_cell_208_120 (.BL(BL120),.BLN(BLN120),.WL(WL208));
sram_cell_6t_5 inst_cell_208_121 (.BL(BL121),.BLN(BLN121),.WL(WL208));
sram_cell_6t_5 inst_cell_208_122 (.BL(BL122),.BLN(BLN122),.WL(WL208));
sram_cell_6t_5 inst_cell_208_123 (.BL(BL123),.BLN(BLN123),.WL(WL208));
sram_cell_6t_5 inst_cell_208_124 (.BL(BL124),.BLN(BLN124),.WL(WL208));
sram_cell_6t_5 inst_cell_208_125 (.BL(BL125),.BLN(BLN125),.WL(WL208));
sram_cell_6t_5 inst_cell_208_126 (.BL(BL126),.BLN(BLN126),.WL(WL208));
sram_cell_6t_5 inst_cell_208_127 (.BL(BL127),.BLN(BLN127),.WL(WL208));
sram_cell_6t_5 inst_cell_209_0 (.BL(BL0),.BLN(BLN0),.WL(WL209));
sram_cell_6t_5 inst_cell_209_1 (.BL(BL1),.BLN(BLN1),.WL(WL209));
sram_cell_6t_5 inst_cell_209_2 (.BL(BL2),.BLN(BLN2),.WL(WL209));
sram_cell_6t_5 inst_cell_209_3 (.BL(BL3),.BLN(BLN3),.WL(WL209));
sram_cell_6t_5 inst_cell_209_4 (.BL(BL4),.BLN(BLN4),.WL(WL209));
sram_cell_6t_5 inst_cell_209_5 (.BL(BL5),.BLN(BLN5),.WL(WL209));
sram_cell_6t_5 inst_cell_209_6 (.BL(BL6),.BLN(BLN6),.WL(WL209));
sram_cell_6t_5 inst_cell_209_7 (.BL(BL7),.BLN(BLN7),.WL(WL209));
sram_cell_6t_5 inst_cell_209_8 (.BL(BL8),.BLN(BLN8),.WL(WL209));
sram_cell_6t_5 inst_cell_209_9 (.BL(BL9),.BLN(BLN9),.WL(WL209));
sram_cell_6t_5 inst_cell_209_10 (.BL(BL10),.BLN(BLN10),.WL(WL209));
sram_cell_6t_5 inst_cell_209_11 (.BL(BL11),.BLN(BLN11),.WL(WL209));
sram_cell_6t_5 inst_cell_209_12 (.BL(BL12),.BLN(BLN12),.WL(WL209));
sram_cell_6t_5 inst_cell_209_13 (.BL(BL13),.BLN(BLN13),.WL(WL209));
sram_cell_6t_5 inst_cell_209_14 (.BL(BL14),.BLN(BLN14),.WL(WL209));
sram_cell_6t_5 inst_cell_209_15 (.BL(BL15),.BLN(BLN15),.WL(WL209));
sram_cell_6t_5 inst_cell_209_16 (.BL(BL16),.BLN(BLN16),.WL(WL209));
sram_cell_6t_5 inst_cell_209_17 (.BL(BL17),.BLN(BLN17),.WL(WL209));
sram_cell_6t_5 inst_cell_209_18 (.BL(BL18),.BLN(BLN18),.WL(WL209));
sram_cell_6t_5 inst_cell_209_19 (.BL(BL19),.BLN(BLN19),.WL(WL209));
sram_cell_6t_5 inst_cell_209_20 (.BL(BL20),.BLN(BLN20),.WL(WL209));
sram_cell_6t_5 inst_cell_209_21 (.BL(BL21),.BLN(BLN21),.WL(WL209));
sram_cell_6t_5 inst_cell_209_22 (.BL(BL22),.BLN(BLN22),.WL(WL209));
sram_cell_6t_5 inst_cell_209_23 (.BL(BL23),.BLN(BLN23),.WL(WL209));
sram_cell_6t_5 inst_cell_209_24 (.BL(BL24),.BLN(BLN24),.WL(WL209));
sram_cell_6t_5 inst_cell_209_25 (.BL(BL25),.BLN(BLN25),.WL(WL209));
sram_cell_6t_5 inst_cell_209_26 (.BL(BL26),.BLN(BLN26),.WL(WL209));
sram_cell_6t_5 inst_cell_209_27 (.BL(BL27),.BLN(BLN27),.WL(WL209));
sram_cell_6t_5 inst_cell_209_28 (.BL(BL28),.BLN(BLN28),.WL(WL209));
sram_cell_6t_5 inst_cell_209_29 (.BL(BL29),.BLN(BLN29),.WL(WL209));
sram_cell_6t_5 inst_cell_209_30 (.BL(BL30),.BLN(BLN30),.WL(WL209));
sram_cell_6t_5 inst_cell_209_31 (.BL(BL31),.BLN(BLN31),.WL(WL209));
sram_cell_6t_5 inst_cell_209_32 (.BL(BL32),.BLN(BLN32),.WL(WL209));
sram_cell_6t_5 inst_cell_209_33 (.BL(BL33),.BLN(BLN33),.WL(WL209));
sram_cell_6t_5 inst_cell_209_34 (.BL(BL34),.BLN(BLN34),.WL(WL209));
sram_cell_6t_5 inst_cell_209_35 (.BL(BL35),.BLN(BLN35),.WL(WL209));
sram_cell_6t_5 inst_cell_209_36 (.BL(BL36),.BLN(BLN36),.WL(WL209));
sram_cell_6t_5 inst_cell_209_37 (.BL(BL37),.BLN(BLN37),.WL(WL209));
sram_cell_6t_5 inst_cell_209_38 (.BL(BL38),.BLN(BLN38),.WL(WL209));
sram_cell_6t_5 inst_cell_209_39 (.BL(BL39),.BLN(BLN39),.WL(WL209));
sram_cell_6t_5 inst_cell_209_40 (.BL(BL40),.BLN(BLN40),.WL(WL209));
sram_cell_6t_5 inst_cell_209_41 (.BL(BL41),.BLN(BLN41),.WL(WL209));
sram_cell_6t_5 inst_cell_209_42 (.BL(BL42),.BLN(BLN42),.WL(WL209));
sram_cell_6t_5 inst_cell_209_43 (.BL(BL43),.BLN(BLN43),.WL(WL209));
sram_cell_6t_5 inst_cell_209_44 (.BL(BL44),.BLN(BLN44),.WL(WL209));
sram_cell_6t_5 inst_cell_209_45 (.BL(BL45),.BLN(BLN45),.WL(WL209));
sram_cell_6t_5 inst_cell_209_46 (.BL(BL46),.BLN(BLN46),.WL(WL209));
sram_cell_6t_5 inst_cell_209_47 (.BL(BL47),.BLN(BLN47),.WL(WL209));
sram_cell_6t_5 inst_cell_209_48 (.BL(BL48),.BLN(BLN48),.WL(WL209));
sram_cell_6t_5 inst_cell_209_49 (.BL(BL49),.BLN(BLN49),.WL(WL209));
sram_cell_6t_5 inst_cell_209_50 (.BL(BL50),.BLN(BLN50),.WL(WL209));
sram_cell_6t_5 inst_cell_209_51 (.BL(BL51),.BLN(BLN51),.WL(WL209));
sram_cell_6t_5 inst_cell_209_52 (.BL(BL52),.BLN(BLN52),.WL(WL209));
sram_cell_6t_5 inst_cell_209_53 (.BL(BL53),.BLN(BLN53),.WL(WL209));
sram_cell_6t_5 inst_cell_209_54 (.BL(BL54),.BLN(BLN54),.WL(WL209));
sram_cell_6t_5 inst_cell_209_55 (.BL(BL55),.BLN(BLN55),.WL(WL209));
sram_cell_6t_5 inst_cell_209_56 (.BL(BL56),.BLN(BLN56),.WL(WL209));
sram_cell_6t_5 inst_cell_209_57 (.BL(BL57),.BLN(BLN57),.WL(WL209));
sram_cell_6t_5 inst_cell_209_58 (.BL(BL58),.BLN(BLN58),.WL(WL209));
sram_cell_6t_5 inst_cell_209_59 (.BL(BL59),.BLN(BLN59),.WL(WL209));
sram_cell_6t_5 inst_cell_209_60 (.BL(BL60),.BLN(BLN60),.WL(WL209));
sram_cell_6t_5 inst_cell_209_61 (.BL(BL61),.BLN(BLN61),.WL(WL209));
sram_cell_6t_5 inst_cell_209_62 (.BL(BL62),.BLN(BLN62),.WL(WL209));
sram_cell_6t_5 inst_cell_209_63 (.BL(BL63),.BLN(BLN63),.WL(WL209));
sram_cell_6t_5 inst_cell_209_64 (.BL(BL64),.BLN(BLN64),.WL(WL209));
sram_cell_6t_5 inst_cell_209_65 (.BL(BL65),.BLN(BLN65),.WL(WL209));
sram_cell_6t_5 inst_cell_209_66 (.BL(BL66),.BLN(BLN66),.WL(WL209));
sram_cell_6t_5 inst_cell_209_67 (.BL(BL67),.BLN(BLN67),.WL(WL209));
sram_cell_6t_5 inst_cell_209_68 (.BL(BL68),.BLN(BLN68),.WL(WL209));
sram_cell_6t_5 inst_cell_209_69 (.BL(BL69),.BLN(BLN69),.WL(WL209));
sram_cell_6t_5 inst_cell_209_70 (.BL(BL70),.BLN(BLN70),.WL(WL209));
sram_cell_6t_5 inst_cell_209_71 (.BL(BL71),.BLN(BLN71),.WL(WL209));
sram_cell_6t_5 inst_cell_209_72 (.BL(BL72),.BLN(BLN72),.WL(WL209));
sram_cell_6t_5 inst_cell_209_73 (.BL(BL73),.BLN(BLN73),.WL(WL209));
sram_cell_6t_5 inst_cell_209_74 (.BL(BL74),.BLN(BLN74),.WL(WL209));
sram_cell_6t_5 inst_cell_209_75 (.BL(BL75),.BLN(BLN75),.WL(WL209));
sram_cell_6t_5 inst_cell_209_76 (.BL(BL76),.BLN(BLN76),.WL(WL209));
sram_cell_6t_5 inst_cell_209_77 (.BL(BL77),.BLN(BLN77),.WL(WL209));
sram_cell_6t_5 inst_cell_209_78 (.BL(BL78),.BLN(BLN78),.WL(WL209));
sram_cell_6t_5 inst_cell_209_79 (.BL(BL79),.BLN(BLN79),.WL(WL209));
sram_cell_6t_5 inst_cell_209_80 (.BL(BL80),.BLN(BLN80),.WL(WL209));
sram_cell_6t_5 inst_cell_209_81 (.BL(BL81),.BLN(BLN81),.WL(WL209));
sram_cell_6t_5 inst_cell_209_82 (.BL(BL82),.BLN(BLN82),.WL(WL209));
sram_cell_6t_5 inst_cell_209_83 (.BL(BL83),.BLN(BLN83),.WL(WL209));
sram_cell_6t_5 inst_cell_209_84 (.BL(BL84),.BLN(BLN84),.WL(WL209));
sram_cell_6t_5 inst_cell_209_85 (.BL(BL85),.BLN(BLN85),.WL(WL209));
sram_cell_6t_5 inst_cell_209_86 (.BL(BL86),.BLN(BLN86),.WL(WL209));
sram_cell_6t_5 inst_cell_209_87 (.BL(BL87),.BLN(BLN87),.WL(WL209));
sram_cell_6t_5 inst_cell_209_88 (.BL(BL88),.BLN(BLN88),.WL(WL209));
sram_cell_6t_5 inst_cell_209_89 (.BL(BL89),.BLN(BLN89),.WL(WL209));
sram_cell_6t_5 inst_cell_209_90 (.BL(BL90),.BLN(BLN90),.WL(WL209));
sram_cell_6t_5 inst_cell_209_91 (.BL(BL91),.BLN(BLN91),.WL(WL209));
sram_cell_6t_5 inst_cell_209_92 (.BL(BL92),.BLN(BLN92),.WL(WL209));
sram_cell_6t_5 inst_cell_209_93 (.BL(BL93),.BLN(BLN93),.WL(WL209));
sram_cell_6t_5 inst_cell_209_94 (.BL(BL94),.BLN(BLN94),.WL(WL209));
sram_cell_6t_5 inst_cell_209_95 (.BL(BL95),.BLN(BLN95),.WL(WL209));
sram_cell_6t_5 inst_cell_209_96 (.BL(BL96),.BLN(BLN96),.WL(WL209));
sram_cell_6t_5 inst_cell_209_97 (.BL(BL97),.BLN(BLN97),.WL(WL209));
sram_cell_6t_5 inst_cell_209_98 (.BL(BL98),.BLN(BLN98),.WL(WL209));
sram_cell_6t_5 inst_cell_209_99 (.BL(BL99),.BLN(BLN99),.WL(WL209));
sram_cell_6t_5 inst_cell_209_100 (.BL(BL100),.BLN(BLN100),.WL(WL209));
sram_cell_6t_5 inst_cell_209_101 (.BL(BL101),.BLN(BLN101),.WL(WL209));
sram_cell_6t_5 inst_cell_209_102 (.BL(BL102),.BLN(BLN102),.WL(WL209));
sram_cell_6t_5 inst_cell_209_103 (.BL(BL103),.BLN(BLN103),.WL(WL209));
sram_cell_6t_5 inst_cell_209_104 (.BL(BL104),.BLN(BLN104),.WL(WL209));
sram_cell_6t_5 inst_cell_209_105 (.BL(BL105),.BLN(BLN105),.WL(WL209));
sram_cell_6t_5 inst_cell_209_106 (.BL(BL106),.BLN(BLN106),.WL(WL209));
sram_cell_6t_5 inst_cell_209_107 (.BL(BL107),.BLN(BLN107),.WL(WL209));
sram_cell_6t_5 inst_cell_209_108 (.BL(BL108),.BLN(BLN108),.WL(WL209));
sram_cell_6t_5 inst_cell_209_109 (.BL(BL109),.BLN(BLN109),.WL(WL209));
sram_cell_6t_5 inst_cell_209_110 (.BL(BL110),.BLN(BLN110),.WL(WL209));
sram_cell_6t_5 inst_cell_209_111 (.BL(BL111),.BLN(BLN111),.WL(WL209));
sram_cell_6t_5 inst_cell_209_112 (.BL(BL112),.BLN(BLN112),.WL(WL209));
sram_cell_6t_5 inst_cell_209_113 (.BL(BL113),.BLN(BLN113),.WL(WL209));
sram_cell_6t_5 inst_cell_209_114 (.BL(BL114),.BLN(BLN114),.WL(WL209));
sram_cell_6t_5 inst_cell_209_115 (.BL(BL115),.BLN(BLN115),.WL(WL209));
sram_cell_6t_5 inst_cell_209_116 (.BL(BL116),.BLN(BLN116),.WL(WL209));
sram_cell_6t_5 inst_cell_209_117 (.BL(BL117),.BLN(BLN117),.WL(WL209));
sram_cell_6t_5 inst_cell_209_118 (.BL(BL118),.BLN(BLN118),.WL(WL209));
sram_cell_6t_5 inst_cell_209_119 (.BL(BL119),.BLN(BLN119),.WL(WL209));
sram_cell_6t_5 inst_cell_209_120 (.BL(BL120),.BLN(BLN120),.WL(WL209));
sram_cell_6t_5 inst_cell_209_121 (.BL(BL121),.BLN(BLN121),.WL(WL209));
sram_cell_6t_5 inst_cell_209_122 (.BL(BL122),.BLN(BLN122),.WL(WL209));
sram_cell_6t_5 inst_cell_209_123 (.BL(BL123),.BLN(BLN123),.WL(WL209));
sram_cell_6t_5 inst_cell_209_124 (.BL(BL124),.BLN(BLN124),.WL(WL209));
sram_cell_6t_5 inst_cell_209_125 (.BL(BL125),.BLN(BLN125),.WL(WL209));
sram_cell_6t_5 inst_cell_209_126 (.BL(BL126),.BLN(BLN126),.WL(WL209));
sram_cell_6t_5 inst_cell_209_127 (.BL(BL127),.BLN(BLN127),.WL(WL209));
sram_cell_6t_5 inst_cell_210_0 (.BL(BL0),.BLN(BLN0),.WL(WL210));
sram_cell_6t_5 inst_cell_210_1 (.BL(BL1),.BLN(BLN1),.WL(WL210));
sram_cell_6t_5 inst_cell_210_2 (.BL(BL2),.BLN(BLN2),.WL(WL210));
sram_cell_6t_5 inst_cell_210_3 (.BL(BL3),.BLN(BLN3),.WL(WL210));
sram_cell_6t_5 inst_cell_210_4 (.BL(BL4),.BLN(BLN4),.WL(WL210));
sram_cell_6t_5 inst_cell_210_5 (.BL(BL5),.BLN(BLN5),.WL(WL210));
sram_cell_6t_5 inst_cell_210_6 (.BL(BL6),.BLN(BLN6),.WL(WL210));
sram_cell_6t_5 inst_cell_210_7 (.BL(BL7),.BLN(BLN7),.WL(WL210));
sram_cell_6t_5 inst_cell_210_8 (.BL(BL8),.BLN(BLN8),.WL(WL210));
sram_cell_6t_5 inst_cell_210_9 (.BL(BL9),.BLN(BLN9),.WL(WL210));
sram_cell_6t_5 inst_cell_210_10 (.BL(BL10),.BLN(BLN10),.WL(WL210));
sram_cell_6t_5 inst_cell_210_11 (.BL(BL11),.BLN(BLN11),.WL(WL210));
sram_cell_6t_5 inst_cell_210_12 (.BL(BL12),.BLN(BLN12),.WL(WL210));
sram_cell_6t_5 inst_cell_210_13 (.BL(BL13),.BLN(BLN13),.WL(WL210));
sram_cell_6t_5 inst_cell_210_14 (.BL(BL14),.BLN(BLN14),.WL(WL210));
sram_cell_6t_5 inst_cell_210_15 (.BL(BL15),.BLN(BLN15),.WL(WL210));
sram_cell_6t_5 inst_cell_210_16 (.BL(BL16),.BLN(BLN16),.WL(WL210));
sram_cell_6t_5 inst_cell_210_17 (.BL(BL17),.BLN(BLN17),.WL(WL210));
sram_cell_6t_5 inst_cell_210_18 (.BL(BL18),.BLN(BLN18),.WL(WL210));
sram_cell_6t_5 inst_cell_210_19 (.BL(BL19),.BLN(BLN19),.WL(WL210));
sram_cell_6t_5 inst_cell_210_20 (.BL(BL20),.BLN(BLN20),.WL(WL210));
sram_cell_6t_5 inst_cell_210_21 (.BL(BL21),.BLN(BLN21),.WL(WL210));
sram_cell_6t_5 inst_cell_210_22 (.BL(BL22),.BLN(BLN22),.WL(WL210));
sram_cell_6t_5 inst_cell_210_23 (.BL(BL23),.BLN(BLN23),.WL(WL210));
sram_cell_6t_5 inst_cell_210_24 (.BL(BL24),.BLN(BLN24),.WL(WL210));
sram_cell_6t_5 inst_cell_210_25 (.BL(BL25),.BLN(BLN25),.WL(WL210));
sram_cell_6t_5 inst_cell_210_26 (.BL(BL26),.BLN(BLN26),.WL(WL210));
sram_cell_6t_5 inst_cell_210_27 (.BL(BL27),.BLN(BLN27),.WL(WL210));
sram_cell_6t_5 inst_cell_210_28 (.BL(BL28),.BLN(BLN28),.WL(WL210));
sram_cell_6t_5 inst_cell_210_29 (.BL(BL29),.BLN(BLN29),.WL(WL210));
sram_cell_6t_5 inst_cell_210_30 (.BL(BL30),.BLN(BLN30),.WL(WL210));
sram_cell_6t_5 inst_cell_210_31 (.BL(BL31),.BLN(BLN31),.WL(WL210));
sram_cell_6t_5 inst_cell_210_32 (.BL(BL32),.BLN(BLN32),.WL(WL210));
sram_cell_6t_5 inst_cell_210_33 (.BL(BL33),.BLN(BLN33),.WL(WL210));
sram_cell_6t_5 inst_cell_210_34 (.BL(BL34),.BLN(BLN34),.WL(WL210));
sram_cell_6t_5 inst_cell_210_35 (.BL(BL35),.BLN(BLN35),.WL(WL210));
sram_cell_6t_5 inst_cell_210_36 (.BL(BL36),.BLN(BLN36),.WL(WL210));
sram_cell_6t_5 inst_cell_210_37 (.BL(BL37),.BLN(BLN37),.WL(WL210));
sram_cell_6t_5 inst_cell_210_38 (.BL(BL38),.BLN(BLN38),.WL(WL210));
sram_cell_6t_5 inst_cell_210_39 (.BL(BL39),.BLN(BLN39),.WL(WL210));
sram_cell_6t_5 inst_cell_210_40 (.BL(BL40),.BLN(BLN40),.WL(WL210));
sram_cell_6t_5 inst_cell_210_41 (.BL(BL41),.BLN(BLN41),.WL(WL210));
sram_cell_6t_5 inst_cell_210_42 (.BL(BL42),.BLN(BLN42),.WL(WL210));
sram_cell_6t_5 inst_cell_210_43 (.BL(BL43),.BLN(BLN43),.WL(WL210));
sram_cell_6t_5 inst_cell_210_44 (.BL(BL44),.BLN(BLN44),.WL(WL210));
sram_cell_6t_5 inst_cell_210_45 (.BL(BL45),.BLN(BLN45),.WL(WL210));
sram_cell_6t_5 inst_cell_210_46 (.BL(BL46),.BLN(BLN46),.WL(WL210));
sram_cell_6t_5 inst_cell_210_47 (.BL(BL47),.BLN(BLN47),.WL(WL210));
sram_cell_6t_5 inst_cell_210_48 (.BL(BL48),.BLN(BLN48),.WL(WL210));
sram_cell_6t_5 inst_cell_210_49 (.BL(BL49),.BLN(BLN49),.WL(WL210));
sram_cell_6t_5 inst_cell_210_50 (.BL(BL50),.BLN(BLN50),.WL(WL210));
sram_cell_6t_5 inst_cell_210_51 (.BL(BL51),.BLN(BLN51),.WL(WL210));
sram_cell_6t_5 inst_cell_210_52 (.BL(BL52),.BLN(BLN52),.WL(WL210));
sram_cell_6t_5 inst_cell_210_53 (.BL(BL53),.BLN(BLN53),.WL(WL210));
sram_cell_6t_5 inst_cell_210_54 (.BL(BL54),.BLN(BLN54),.WL(WL210));
sram_cell_6t_5 inst_cell_210_55 (.BL(BL55),.BLN(BLN55),.WL(WL210));
sram_cell_6t_5 inst_cell_210_56 (.BL(BL56),.BLN(BLN56),.WL(WL210));
sram_cell_6t_5 inst_cell_210_57 (.BL(BL57),.BLN(BLN57),.WL(WL210));
sram_cell_6t_5 inst_cell_210_58 (.BL(BL58),.BLN(BLN58),.WL(WL210));
sram_cell_6t_5 inst_cell_210_59 (.BL(BL59),.BLN(BLN59),.WL(WL210));
sram_cell_6t_5 inst_cell_210_60 (.BL(BL60),.BLN(BLN60),.WL(WL210));
sram_cell_6t_5 inst_cell_210_61 (.BL(BL61),.BLN(BLN61),.WL(WL210));
sram_cell_6t_5 inst_cell_210_62 (.BL(BL62),.BLN(BLN62),.WL(WL210));
sram_cell_6t_5 inst_cell_210_63 (.BL(BL63),.BLN(BLN63),.WL(WL210));
sram_cell_6t_5 inst_cell_210_64 (.BL(BL64),.BLN(BLN64),.WL(WL210));
sram_cell_6t_5 inst_cell_210_65 (.BL(BL65),.BLN(BLN65),.WL(WL210));
sram_cell_6t_5 inst_cell_210_66 (.BL(BL66),.BLN(BLN66),.WL(WL210));
sram_cell_6t_5 inst_cell_210_67 (.BL(BL67),.BLN(BLN67),.WL(WL210));
sram_cell_6t_5 inst_cell_210_68 (.BL(BL68),.BLN(BLN68),.WL(WL210));
sram_cell_6t_5 inst_cell_210_69 (.BL(BL69),.BLN(BLN69),.WL(WL210));
sram_cell_6t_5 inst_cell_210_70 (.BL(BL70),.BLN(BLN70),.WL(WL210));
sram_cell_6t_5 inst_cell_210_71 (.BL(BL71),.BLN(BLN71),.WL(WL210));
sram_cell_6t_5 inst_cell_210_72 (.BL(BL72),.BLN(BLN72),.WL(WL210));
sram_cell_6t_5 inst_cell_210_73 (.BL(BL73),.BLN(BLN73),.WL(WL210));
sram_cell_6t_5 inst_cell_210_74 (.BL(BL74),.BLN(BLN74),.WL(WL210));
sram_cell_6t_5 inst_cell_210_75 (.BL(BL75),.BLN(BLN75),.WL(WL210));
sram_cell_6t_5 inst_cell_210_76 (.BL(BL76),.BLN(BLN76),.WL(WL210));
sram_cell_6t_5 inst_cell_210_77 (.BL(BL77),.BLN(BLN77),.WL(WL210));
sram_cell_6t_5 inst_cell_210_78 (.BL(BL78),.BLN(BLN78),.WL(WL210));
sram_cell_6t_5 inst_cell_210_79 (.BL(BL79),.BLN(BLN79),.WL(WL210));
sram_cell_6t_5 inst_cell_210_80 (.BL(BL80),.BLN(BLN80),.WL(WL210));
sram_cell_6t_5 inst_cell_210_81 (.BL(BL81),.BLN(BLN81),.WL(WL210));
sram_cell_6t_5 inst_cell_210_82 (.BL(BL82),.BLN(BLN82),.WL(WL210));
sram_cell_6t_5 inst_cell_210_83 (.BL(BL83),.BLN(BLN83),.WL(WL210));
sram_cell_6t_5 inst_cell_210_84 (.BL(BL84),.BLN(BLN84),.WL(WL210));
sram_cell_6t_5 inst_cell_210_85 (.BL(BL85),.BLN(BLN85),.WL(WL210));
sram_cell_6t_5 inst_cell_210_86 (.BL(BL86),.BLN(BLN86),.WL(WL210));
sram_cell_6t_5 inst_cell_210_87 (.BL(BL87),.BLN(BLN87),.WL(WL210));
sram_cell_6t_5 inst_cell_210_88 (.BL(BL88),.BLN(BLN88),.WL(WL210));
sram_cell_6t_5 inst_cell_210_89 (.BL(BL89),.BLN(BLN89),.WL(WL210));
sram_cell_6t_5 inst_cell_210_90 (.BL(BL90),.BLN(BLN90),.WL(WL210));
sram_cell_6t_5 inst_cell_210_91 (.BL(BL91),.BLN(BLN91),.WL(WL210));
sram_cell_6t_5 inst_cell_210_92 (.BL(BL92),.BLN(BLN92),.WL(WL210));
sram_cell_6t_5 inst_cell_210_93 (.BL(BL93),.BLN(BLN93),.WL(WL210));
sram_cell_6t_5 inst_cell_210_94 (.BL(BL94),.BLN(BLN94),.WL(WL210));
sram_cell_6t_5 inst_cell_210_95 (.BL(BL95),.BLN(BLN95),.WL(WL210));
sram_cell_6t_5 inst_cell_210_96 (.BL(BL96),.BLN(BLN96),.WL(WL210));
sram_cell_6t_5 inst_cell_210_97 (.BL(BL97),.BLN(BLN97),.WL(WL210));
sram_cell_6t_5 inst_cell_210_98 (.BL(BL98),.BLN(BLN98),.WL(WL210));
sram_cell_6t_5 inst_cell_210_99 (.BL(BL99),.BLN(BLN99),.WL(WL210));
sram_cell_6t_5 inst_cell_210_100 (.BL(BL100),.BLN(BLN100),.WL(WL210));
sram_cell_6t_5 inst_cell_210_101 (.BL(BL101),.BLN(BLN101),.WL(WL210));
sram_cell_6t_5 inst_cell_210_102 (.BL(BL102),.BLN(BLN102),.WL(WL210));
sram_cell_6t_5 inst_cell_210_103 (.BL(BL103),.BLN(BLN103),.WL(WL210));
sram_cell_6t_5 inst_cell_210_104 (.BL(BL104),.BLN(BLN104),.WL(WL210));
sram_cell_6t_5 inst_cell_210_105 (.BL(BL105),.BLN(BLN105),.WL(WL210));
sram_cell_6t_5 inst_cell_210_106 (.BL(BL106),.BLN(BLN106),.WL(WL210));
sram_cell_6t_5 inst_cell_210_107 (.BL(BL107),.BLN(BLN107),.WL(WL210));
sram_cell_6t_5 inst_cell_210_108 (.BL(BL108),.BLN(BLN108),.WL(WL210));
sram_cell_6t_5 inst_cell_210_109 (.BL(BL109),.BLN(BLN109),.WL(WL210));
sram_cell_6t_5 inst_cell_210_110 (.BL(BL110),.BLN(BLN110),.WL(WL210));
sram_cell_6t_5 inst_cell_210_111 (.BL(BL111),.BLN(BLN111),.WL(WL210));
sram_cell_6t_5 inst_cell_210_112 (.BL(BL112),.BLN(BLN112),.WL(WL210));
sram_cell_6t_5 inst_cell_210_113 (.BL(BL113),.BLN(BLN113),.WL(WL210));
sram_cell_6t_5 inst_cell_210_114 (.BL(BL114),.BLN(BLN114),.WL(WL210));
sram_cell_6t_5 inst_cell_210_115 (.BL(BL115),.BLN(BLN115),.WL(WL210));
sram_cell_6t_5 inst_cell_210_116 (.BL(BL116),.BLN(BLN116),.WL(WL210));
sram_cell_6t_5 inst_cell_210_117 (.BL(BL117),.BLN(BLN117),.WL(WL210));
sram_cell_6t_5 inst_cell_210_118 (.BL(BL118),.BLN(BLN118),.WL(WL210));
sram_cell_6t_5 inst_cell_210_119 (.BL(BL119),.BLN(BLN119),.WL(WL210));
sram_cell_6t_5 inst_cell_210_120 (.BL(BL120),.BLN(BLN120),.WL(WL210));
sram_cell_6t_5 inst_cell_210_121 (.BL(BL121),.BLN(BLN121),.WL(WL210));
sram_cell_6t_5 inst_cell_210_122 (.BL(BL122),.BLN(BLN122),.WL(WL210));
sram_cell_6t_5 inst_cell_210_123 (.BL(BL123),.BLN(BLN123),.WL(WL210));
sram_cell_6t_5 inst_cell_210_124 (.BL(BL124),.BLN(BLN124),.WL(WL210));
sram_cell_6t_5 inst_cell_210_125 (.BL(BL125),.BLN(BLN125),.WL(WL210));
sram_cell_6t_5 inst_cell_210_126 (.BL(BL126),.BLN(BLN126),.WL(WL210));
sram_cell_6t_5 inst_cell_210_127 (.BL(BL127),.BLN(BLN127),.WL(WL210));
sram_cell_6t_5 inst_cell_211_0 (.BL(BL0),.BLN(BLN0),.WL(WL211));
sram_cell_6t_5 inst_cell_211_1 (.BL(BL1),.BLN(BLN1),.WL(WL211));
sram_cell_6t_5 inst_cell_211_2 (.BL(BL2),.BLN(BLN2),.WL(WL211));
sram_cell_6t_5 inst_cell_211_3 (.BL(BL3),.BLN(BLN3),.WL(WL211));
sram_cell_6t_5 inst_cell_211_4 (.BL(BL4),.BLN(BLN4),.WL(WL211));
sram_cell_6t_5 inst_cell_211_5 (.BL(BL5),.BLN(BLN5),.WL(WL211));
sram_cell_6t_5 inst_cell_211_6 (.BL(BL6),.BLN(BLN6),.WL(WL211));
sram_cell_6t_5 inst_cell_211_7 (.BL(BL7),.BLN(BLN7),.WL(WL211));
sram_cell_6t_5 inst_cell_211_8 (.BL(BL8),.BLN(BLN8),.WL(WL211));
sram_cell_6t_5 inst_cell_211_9 (.BL(BL9),.BLN(BLN9),.WL(WL211));
sram_cell_6t_5 inst_cell_211_10 (.BL(BL10),.BLN(BLN10),.WL(WL211));
sram_cell_6t_5 inst_cell_211_11 (.BL(BL11),.BLN(BLN11),.WL(WL211));
sram_cell_6t_5 inst_cell_211_12 (.BL(BL12),.BLN(BLN12),.WL(WL211));
sram_cell_6t_5 inst_cell_211_13 (.BL(BL13),.BLN(BLN13),.WL(WL211));
sram_cell_6t_5 inst_cell_211_14 (.BL(BL14),.BLN(BLN14),.WL(WL211));
sram_cell_6t_5 inst_cell_211_15 (.BL(BL15),.BLN(BLN15),.WL(WL211));
sram_cell_6t_5 inst_cell_211_16 (.BL(BL16),.BLN(BLN16),.WL(WL211));
sram_cell_6t_5 inst_cell_211_17 (.BL(BL17),.BLN(BLN17),.WL(WL211));
sram_cell_6t_5 inst_cell_211_18 (.BL(BL18),.BLN(BLN18),.WL(WL211));
sram_cell_6t_5 inst_cell_211_19 (.BL(BL19),.BLN(BLN19),.WL(WL211));
sram_cell_6t_5 inst_cell_211_20 (.BL(BL20),.BLN(BLN20),.WL(WL211));
sram_cell_6t_5 inst_cell_211_21 (.BL(BL21),.BLN(BLN21),.WL(WL211));
sram_cell_6t_5 inst_cell_211_22 (.BL(BL22),.BLN(BLN22),.WL(WL211));
sram_cell_6t_5 inst_cell_211_23 (.BL(BL23),.BLN(BLN23),.WL(WL211));
sram_cell_6t_5 inst_cell_211_24 (.BL(BL24),.BLN(BLN24),.WL(WL211));
sram_cell_6t_5 inst_cell_211_25 (.BL(BL25),.BLN(BLN25),.WL(WL211));
sram_cell_6t_5 inst_cell_211_26 (.BL(BL26),.BLN(BLN26),.WL(WL211));
sram_cell_6t_5 inst_cell_211_27 (.BL(BL27),.BLN(BLN27),.WL(WL211));
sram_cell_6t_5 inst_cell_211_28 (.BL(BL28),.BLN(BLN28),.WL(WL211));
sram_cell_6t_5 inst_cell_211_29 (.BL(BL29),.BLN(BLN29),.WL(WL211));
sram_cell_6t_5 inst_cell_211_30 (.BL(BL30),.BLN(BLN30),.WL(WL211));
sram_cell_6t_5 inst_cell_211_31 (.BL(BL31),.BLN(BLN31),.WL(WL211));
sram_cell_6t_5 inst_cell_211_32 (.BL(BL32),.BLN(BLN32),.WL(WL211));
sram_cell_6t_5 inst_cell_211_33 (.BL(BL33),.BLN(BLN33),.WL(WL211));
sram_cell_6t_5 inst_cell_211_34 (.BL(BL34),.BLN(BLN34),.WL(WL211));
sram_cell_6t_5 inst_cell_211_35 (.BL(BL35),.BLN(BLN35),.WL(WL211));
sram_cell_6t_5 inst_cell_211_36 (.BL(BL36),.BLN(BLN36),.WL(WL211));
sram_cell_6t_5 inst_cell_211_37 (.BL(BL37),.BLN(BLN37),.WL(WL211));
sram_cell_6t_5 inst_cell_211_38 (.BL(BL38),.BLN(BLN38),.WL(WL211));
sram_cell_6t_5 inst_cell_211_39 (.BL(BL39),.BLN(BLN39),.WL(WL211));
sram_cell_6t_5 inst_cell_211_40 (.BL(BL40),.BLN(BLN40),.WL(WL211));
sram_cell_6t_5 inst_cell_211_41 (.BL(BL41),.BLN(BLN41),.WL(WL211));
sram_cell_6t_5 inst_cell_211_42 (.BL(BL42),.BLN(BLN42),.WL(WL211));
sram_cell_6t_5 inst_cell_211_43 (.BL(BL43),.BLN(BLN43),.WL(WL211));
sram_cell_6t_5 inst_cell_211_44 (.BL(BL44),.BLN(BLN44),.WL(WL211));
sram_cell_6t_5 inst_cell_211_45 (.BL(BL45),.BLN(BLN45),.WL(WL211));
sram_cell_6t_5 inst_cell_211_46 (.BL(BL46),.BLN(BLN46),.WL(WL211));
sram_cell_6t_5 inst_cell_211_47 (.BL(BL47),.BLN(BLN47),.WL(WL211));
sram_cell_6t_5 inst_cell_211_48 (.BL(BL48),.BLN(BLN48),.WL(WL211));
sram_cell_6t_5 inst_cell_211_49 (.BL(BL49),.BLN(BLN49),.WL(WL211));
sram_cell_6t_5 inst_cell_211_50 (.BL(BL50),.BLN(BLN50),.WL(WL211));
sram_cell_6t_5 inst_cell_211_51 (.BL(BL51),.BLN(BLN51),.WL(WL211));
sram_cell_6t_5 inst_cell_211_52 (.BL(BL52),.BLN(BLN52),.WL(WL211));
sram_cell_6t_5 inst_cell_211_53 (.BL(BL53),.BLN(BLN53),.WL(WL211));
sram_cell_6t_5 inst_cell_211_54 (.BL(BL54),.BLN(BLN54),.WL(WL211));
sram_cell_6t_5 inst_cell_211_55 (.BL(BL55),.BLN(BLN55),.WL(WL211));
sram_cell_6t_5 inst_cell_211_56 (.BL(BL56),.BLN(BLN56),.WL(WL211));
sram_cell_6t_5 inst_cell_211_57 (.BL(BL57),.BLN(BLN57),.WL(WL211));
sram_cell_6t_5 inst_cell_211_58 (.BL(BL58),.BLN(BLN58),.WL(WL211));
sram_cell_6t_5 inst_cell_211_59 (.BL(BL59),.BLN(BLN59),.WL(WL211));
sram_cell_6t_5 inst_cell_211_60 (.BL(BL60),.BLN(BLN60),.WL(WL211));
sram_cell_6t_5 inst_cell_211_61 (.BL(BL61),.BLN(BLN61),.WL(WL211));
sram_cell_6t_5 inst_cell_211_62 (.BL(BL62),.BLN(BLN62),.WL(WL211));
sram_cell_6t_5 inst_cell_211_63 (.BL(BL63),.BLN(BLN63),.WL(WL211));
sram_cell_6t_5 inst_cell_211_64 (.BL(BL64),.BLN(BLN64),.WL(WL211));
sram_cell_6t_5 inst_cell_211_65 (.BL(BL65),.BLN(BLN65),.WL(WL211));
sram_cell_6t_5 inst_cell_211_66 (.BL(BL66),.BLN(BLN66),.WL(WL211));
sram_cell_6t_5 inst_cell_211_67 (.BL(BL67),.BLN(BLN67),.WL(WL211));
sram_cell_6t_5 inst_cell_211_68 (.BL(BL68),.BLN(BLN68),.WL(WL211));
sram_cell_6t_5 inst_cell_211_69 (.BL(BL69),.BLN(BLN69),.WL(WL211));
sram_cell_6t_5 inst_cell_211_70 (.BL(BL70),.BLN(BLN70),.WL(WL211));
sram_cell_6t_5 inst_cell_211_71 (.BL(BL71),.BLN(BLN71),.WL(WL211));
sram_cell_6t_5 inst_cell_211_72 (.BL(BL72),.BLN(BLN72),.WL(WL211));
sram_cell_6t_5 inst_cell_211_73 (.BL(BL73),.BLN(BLN73),.WL(WL211));
sram_cell_6t_5 inst_cell_211_74 (.BL(BL74),.BLN(BLN74),.WL(WL211));
sram_cell_6t_5 inst_cell_211_75 (.BL(BL75),.BLN(BLN75),.WL(WL211));
sram_cell_6t_5 inst_cell_211_76 (.BL(BL76),.BLN(BLN76),.WL(WL211));
sram_cell_6t_5 inst_cell_211_77 (.BL(BL77),.BLN(BLN77),.WL(WL211));
sram_cell_6t_5 inst_cell_211_78 (.BL(BL78),.BLN(BLN78),.WL(WL211));
sram_cell_6t_5 inst_cell_211_79 (.BL(BL79),.BLN(BLN79),.WL(WL211));
sram_cell_6t_5 inst_cell_211_80 (.BL(BL80),.BLN(BLN80),.WL(WL211));
sram_cell_6t_5 inst_cell_211_81 (.BL(BL81),.BLN(BLN81),.WL(WL211));
sram_cell_6t_5 inst_cell_211_82 (.BL(BL82),.BLN(BLN82),.WL(WL211));
sram_cell_6t_5 inst_cell_211_83 (.BL(BL83),.BLN(BLN83),.WL(WL211));
sram_cell_6t_5 inst_cell_211_84 (.BL(BL84),.BLN(BLN84),.WL(WL211));
sram_cell_6t_5 inst_cell_211_85 (.BL(BL85),.BLN(BLN85),.WL(WL211));
sram_cell_6t_5 inst_cell_211_86 (.BL(BL86),.BLN(BLN86),.WL(WL211));
sram_cell_6t_5 inst_cell_211_87 (.BL(BL87),.BLN(BLN87),.WL(WL211));
sram_cell_6t_5 inst_cell_211_88 (.BL(BL88),.BLN(BLN88),.WL(WL211));
sram_cell_6t_5 inst_cell_211_89 (.BL(BL89),.BLN(BLN89),.WL(WL211));
sram_cell_6t_5 inst_cell_211_90 (.BL(BL90),.BLN(BLN90),.WL(WL211));
sram_cell_6t_5 inst_cell_211_91 (.BL(BL91),.BLN(BLN91),.WL(WL211));
sram_cell_6t_5 inst_cell_211_92 (.BL(BL92),.BLN(BLN92),.WL(WL211));
sram_cell_6t_5 inst_cell_211_93 (.BL(BL93),.BLN(BLN93),.WL(WL211));
sram_cell_6t_5 inst_cell_211_94 (.BL(BL94),.BLN(BLN94),.WL(WL211));
sram_cell_6t_5 inst_cell_211_95 (.BL(BL95),.BLN(BLN95),.WL(WL211));
sram_cell_6t_5 inst_cell_211_96 (.BL(BL96),.BLN(BLN96),.WL(WL211));
sram_cell_6t_5 inst_cell_211_97 (.BL(BL97),.BLN(BLN97),.WL(WL211));
sram_cell_6t_5 inst_cell_211_98 (.BL(BL98),.BLN(BLN98),.WL(WL211));
sram_cell_6t_5 inst_cell_211_99 (.BL(BL99),.BLN(BLN99),.WL(WL211));
sram_cell_6t_5 inst_cell_211_100 (.BL(BL100),.BLN(BLN100),.WL(WL211));
sram_cell_6t_5 inst_cell_211_101 (.BL(BL101),.BLN(BLN101),.WL(WL211));
sram_cell_6t_5 inst_cell_211_102 (.BL(BL102),.BLN(BLN102),.WL(WL211));
sram_cell_6t_5 inst_cell_211_103 (.BL(BL103),.BLN(BLN103),.WL(WL211));
sram_cell_6t_5 inst_cell_211_104 (.BL(BL104),.BLN(BLN104),.WL(WL211));
sram_cell_6t_5 inst_cell_211_105 (.BL(BL105),.BLN(BLN105),.WL(WL211));
sram_cell_6t_5 inst_cell_211_106 (.BL(BL106),.BLN(BLN106),.WL(WL211));
sram_cell_6t_5 inst_cell_211_107 (.BL(BL107),.BLN(BLN107),.WL(WL211));
sram_cell_6t_5 inst_cell_211_108 (.BL(BL108),.BLN(BLN108),.WL(WL211));
sram_cell_6t_5 inst_cell_211_109 (.BL(BL109),.BLN(BLN109),.WL(WL211));
sram_cell_6t_5 inst_cell_211_110 (.BL(BL110),.BLN(BLN110),.WL(WL211));
sram_cell_6t_5 inst_cell_211_111 (.BL(BL111),.BLN(BLN111),.WL(WL211));
sram_cell_6t_5 inst_cell_211_112 (.BL(BL112),.BLN(BLN112),.WL(WL211));
sram_cell_6t_5 inst_cell_211_113 (.BL(BL113),.BLN(BLN113),.WL(WL211));
sram_cell_6t_5 inst_cell_211_114 (.BL(BL114),.BLN(BLN114),.WL(WL211));
sram_cell_6t_5 inst_cell_211_115 (.BL(BL115),.BLN(BLN115),.WL(WL211));
sram_cell_6t_5 inst_cell_211_116 (.BL(BL116),.BLN(BLN116),.WL(WL211));
sram_cell_6t_5 inst_cell_211_117 (.BL(BL117),.BLN(BLN117),.WL(WL211));
sram_cell_6t_5 inst_cell_211_118 (.BL(BL118),.BLN(BLN118),.WL(WL211));
sram_cell_6t_5 inst_cell_211_119 (.BL(BL119),.BLN(BLN119),.WL(WL211));
sram_cell_6t_5 inst_cell_211_120 (.BL(BL120),.BLN(BLN120),.WL(WL211));
sram_cell_6t_5 inst_cell_211_121 (.BL(BL121),.BLN(BLN121),.WL(WL211));
sram_cell_6t_5 inst_cell_211_122 (.BL(BL122),.BLN(BLN122),.WL(WL211));
sram_cell_6t_5 inst_cell_211_123 (.BL(BL123),.BLN(BLN123),.WL(WL211));
sram_cell_6t_5 inst_cell_211_124 (.BL(BL124),.BLN(BLN124),.WL(WL211));
sram_cell_6t_5 inst_cell_211_125 (.BL(BL125),.BLN(BLN125),.WL(WL211));
sram_cell_6t_5 inst_cell_211_126 (.BL(BL126),.BLN(BLN126),.WL(WL211));
sram_cell_6t_5 inst_cell_211_127 (.BL(BL127),.BLN(BLN127),.WL(WL211));
sram_cell_6t_5 inst_cell_212_0 (.BL(BL0),.BLN(BLN0),.WL(WL212));
sram_cell_6t_5 inst_cell_212_1 (.BL(BL1),.BLN(BLN1),.WL(WL212));
sram_cell_6t_5 inst_cell_212_2 (.BL(BL2),.BLN(BLN2),.WL(WL212));
sram_cell_6t_5 inst_cell_212_3 (.BL(BL3),.BLN(BLN3),.WL(WL212));
sram_cell_6t_5 inst_cell_212_4 (.BL(BL4),.BLN(BLN4),.WL(WL212));
sram_cell_6t_5 inst_cell_212_5 (.BL(BL5),.BLN(BLN5),.WL(WL212));
sram_cell_6t_5 inst_cell_212_6 (.BL(BL6),.BLN(BLN6),.WL(WL212));
sram_cell_6t_5 inst_cell_212_7 (.BL(BL7),.BLN(BLN7),.WL(WL212));
sram_cell_6t_5 inst_cell_212_8 (.BL(BL8),.BLN(BLN8),.WL(WL212));
sram_cell_6t_5 inst_cell_212_9 (.BL(BL9),.BLN(BLN9),.WL(WL212));
sram_cell_6t_5 inst_cell_212_10 (.BL(BL10),.BLN(BLN10),.WL(WL212));
sram_cell_6t_5 inst_cell_212_11 (.BL(BL11),.BLN(BLN11),.WL(WL212));
sram_cell_6t_5 inst_cell_212_12 (.BL(BL12),.BLN(BLN12),.WL(WL212));
sram_cell_6t_5 inst_cell_212_13 (.BL(BL13),.BLN(BLN13),.WL(WL212));
sram_cell_6t_5 inst_cell_212_14 (.BL(BL14),.BLN(BLN14),.WL(WL212));
sram_cell_6t_5 inst_cell_212_15 (.BL(BL15),.BLN(BLN15),.WL(WL212));
sram_cell_6t_5 inst_cell_212_16 (.BL(BL16),.BLN(BLN16),.WL(WL212));
sram_cell_6t_5 inst_cell_212_17 (.BL(BL17),.BLN(BLN17),.WL(WL212));
sram_cell_6t_5 inst_cell_212_18 (.BL(BL18),.BLN(BLN18),.WL(WL212));
sram_cell_6t_5 inst_cell_212_19 (.BL(BL19),.BLN(BLN19),.WL(WL212));
sram_cell_6t_5 inst_cell_212_20 (.BL(BL20),.BLN(BLN20),.WL(WL212));
sram_cell_6t_5 inst_cell_212_21 (.BL(BL21),.BLN(BLN21),.WL(WL212));
sram_cell_6t_5 inst_cell_212_22 (.BL(BL22),.BLN(BLN22),.WL(WL212));
sram_cell_6t_5 inst_cell_212_23 (.BL(BL23),.BLN(BLN23),.WL(WL212));
sram_cell_6t_5 inst_cell_212_24 (.BL(BL24),.BLN(BLN24),.WL(WL212));
sram_cell_6t_5 inst_cell_212_25 (.BL(BL25),.BLN(BLN25),.WL(WL212));
sram_cell_6t_5 inst_cell_212_26 (.BL(BL26),.BLN(BLN26),.WL(WL212));
sram_cell_6t_5 inst_cell_212_27 (.BL(BL27),.BLN(BLN27),.WL(WL212));
sram_cell_6t_5 inst_cell_212_28 (.BL(BL28),.BLN(BLN28),.WL(WL212));
sram_cell_6t_5 inst_cell_212_29 (.BL(BL29),.BLN(BLN29),.WL(WL212));
sram_cell_6t_5 inst_cell_212_30 (.BL(BL30),.BLN(BLN30),.WL(WL212));
sram_cell_6t_5 inst_cell_212_31 (.BL(BL31),.BLN(BLN31),.WL(WL212));
sram_cell_6t_5 inst_cell_212_32 (.BL(BL32),.BLN(BLN32),.WL(WL212));
sram_cell_6t_5 inst_cell_212_33 (.BL(BL33),.BLN(BLN33),.WL(WL212));
sram_cell_6t_5 inst_cell_212_34 (.BL(BL34),.BLN(BLN34),.WL(WL212));
sram_cell_6t_5 inst_cell_212_35 (.BL(BL35),.BLN(BLN35),.WL(WL212));
sram_cell_6t_5 inst_cell_212_36 (.BL(BL36),.BLN(BLN36),.WL(WL212));
sram_cell_6t_5 inst_cell_212_37 (.BL(BL37),.BLN(BLN37),.WL(WL212));
sram_cell_6t_5 inst_cell_212_38 (.BL(BL38),.BLN(BLN38),.WL(WL212));
sram_cell_6t_5 inst_cell_212_39 (.BL(BL39),.BLN(BLN39),.WL(WL212));
sram_cell_6t_5 inst_cell_212_40 (.BL(BL40),.BLN(BLN40),.WL(WL212));
sram_cell_6t_5 inst_cell_212_41 (.BL(BL41),.BLN(BLN41),.WL(WL212));
sram_cell_6t_5 inst_cell_212_42 (.BL(BL42),.BLN(BLN42),.WL(WL212));
sram_cell_6t_5 inst_cell_212_43 (.BL(BL43),.BLN(BLN43),.WL(WL212));
sram_cell_6t_5 inst_cell_212_44 (.BL(BL44),.BLN(BLN44),.WL(WL212));
sram_cell_6t_5 inst_cell_212_45 (.BL(BL45),.BLN(BLN45),.WL(WL212));
sram_cell_6t_5 inst_cell_212_46 (.BL(BL46),.BLN(BLN46),.WL(WL212));
sram_cell_6t_5 inst_cell_212_47 (.BL(BL47),.BLN(BLN47),.WL(WL212));
sram_cell_6t_5 inst_cell_212_48 (.BL(BL48),.BLN(BLN48),.WL(WL212));
sram_cell_6t_5 inst_cell_212_49 (.BL(BL49),.BLN(BLN49),.WL(WL212));
sram_cell_6t_5 inst_cell_212_50 (.BL(BL50),.BLN(BLN50),.WL(WL212));
sram_cell_6t_5 inst_cell_212_51 (.BL(BL51),.BLN(BLN51),.WL(WL212));
sram_cell_6t_5 inst_cell_212_52 (.BL(BL52),.BLN(BLN52),.WL(WL212));
sram_cell_6t_5 inst_cell_212_53 (.BL(BL53),.BLN(BLN53),.WL(WL212));
sram_cell_6t_5 inst_cell_212_54 (.BL(BL54),.BLN(BLN54),.WL(WL212));
sram_cell_6t_5 inst_cell_212_55 (.BL(BL55),.BLN(BLN55),.WL(WL212));
sram_cell_6t_5 inst_cell_212_56 (.BL(BL56),.BLN(BLN56),.WL(WL212));
sram_cell_6t_5 inst_cell_212_57 (.BL(BL57),.BLN(BLN57),.WL(WL212));
sram_cell_6t_5 inst_cell_212_58 (.BL(BL58),.BLN(BLN58),.WL(WL212));
sram_cell_6t_5 inst_cell_212_59 (.BL(BL59),.BLN(BLN59),.WL(WL212));
sram_cell_6t_5 inst_cell_212_60 (.BL(BL60),.BLN(BLN60),.WL(WL212));
sram_cell_6t_5 inst_cell_212_61 (.BL(BL61),.BLN(BLN61),.WL(WL212));
sram_cell_6t_5 inst_cell_212_62 (.BL(BL62),.BLN(BLN62),.WL(WL212));
sram_cell_6t_5 inst_cell_212_63 (.BL(BL63),.BLN(BLN63),.WL(WL212));
sram_cell_6t_5 inst_cell_212_64 (.BL(BL64),.BLN(BLN64),.WL(WL212));
sram_cell_6t_5 inst_cell_212_65 (.BL(BL65),.BLN(BLN65),.WL(WL212));
sram_cell_6t_5 inst_cell_212_66 (.BL(BL66),.BLN(BLN66),.WL(WL212));
sram_cell_6t_5 inst_cell_212_67 (.BL(BL67),.BLN(BLN67),.WL(WL212));
sram_cell_6t_5 inst_cell_212_68 (.BL(BL68),.BLN(BLN68),.WL(WL212));
sram_cell_6t_5 inst_cell_212_69 (.BL(BL69),.BLN(BLN69),.WL(WL212));
sram_cell_6t_5 inst_cell_212_70 (.BL(BL70),.BLN(BLN70),.WL(WL212));
sram_cell_6t_5 inst_cell_212_71 (.BL(BL71),.BLN(BLN71),.WL(WL212));
sram_cell_6t_5 inst_cell_212_72 (.BL(BL72),.BLN(BLN72),.WL(WL212));
sram_cell_6t_5 inst_cell_212_73 (.BL(BL73),.BLN(BLN73),.WL(WL212));
sram_cell_6t_5 inst_cell_212_74 (.BL(BL74),.BLN(BLN74),.WL(WL212));
sram_cell_6t_5 inst_cell_212_75 (.BL(BL75),.BLN(BLN75),.WL(WL212));
sram_cell_6t_5 inst_cell_212_76 (.BL(BL76),.BLN(BLN76),.WL(WL212));
sram_cell_6t_5 inst_cell_212_77 (.BL(BL77),.BLN(BLN77),.WL(WL212));
sram_cell_6t_5 inst_cell_212_78 (.BL(BL78),.BLN(BLN78),.WL(WL212));
sram_cell_6t_5 inst_cell_212_79 (.BL(BL79),.BLN(BLN79),.WL(WL212));
sram_cell_6t_5 inst_cell_212_80 (.BL(BL80),.BLN(BLN80),.WL(WL212));
sram_cell_6t_5 inst_cell_212_81 (.BL(BL81),.BLN(BLN81),.WL(WL212));
sram_cell_6t_5 inst_cell_212_82 (.BL(BL82),.BLN(BLN82),.WL(WL212));
sram_cell_6t_5 inst_cell_212_83 (.BL(BL83),.BLN(BLN83),.WL(WL212));
sram_cell_6t_5 inst_cell_212_84 (.BL(BL84),.BLN(BLN84),.WL(WL212));
sram_cell_6t_5 inst_cell_212_85 (.BL(BL85),.BLN(BLN85),.WL(WL212));
sram_cell_6t_5 inst_cell_212_86 (.BL(BL86),.BLN(BLN86),.WL(WL212));
sram_cell_6t_5 inst_cell_212_87 (.BL(BL87),.BLN(BLN87),.WL(WL212));
sram_cell_6t_5 inst_cell_212_88 (.BL(BL88),.BLN(BLN88),.WL(WL212));
sram_cell_6t_5 inst_cell_212_89 (.BL(BL89),.BLN(BLN89),.WL(WL212));
sram_cell_6t_5 inst_cell_212_90 (.BL(BL90),.BLN(BLN90),.WL(WL212));
sram_cell_6t_5 inst_cell_212_91 (.BL(BL91),.BLN(BLN91),.WL(WL212));
sram_cell_6t_5 inst_cell_212_92 (.BL(BL92),.BLN(BLN92),.WL(WL212));
sram_cell_6t_5 inst_cell_212_93 (.BL(BL93),.BLN(BLN93),.WL(WL212));
sram_cell_6t_5 inst_cell_212_94 (.BL(BL94),.BLN(BLN94),.WL(WL212));
sram_cell_6t_5 inst_cell_212_95 (.BL(BL95),.BLN(BLN95),.WL(WL212));
sram_cell_6t_5 inst_cell_212_96 (.BL(BL96),.BLN(BLN96),.WL(WL212));
sram_cell_6t_5 inst_cell_212_97 (.BL(BL97),.BLN(BLN97),.WL(WL212));
sram_cell_6t_5 inst_cell_212_98 (.BL(BL98),.BLN(BLN98),.WL(WL212));
sram_cell_6t_5 inst_cell_212_99 (.BL(BL99),.BLN(BLN99),.WL(WL212));
sram_cell_6t_5 inst_cell_212_100 (.BL(BL100),.BLN(BLN100),.WL(WL212));
sram_cell_6t_5 inst_cell_212_101 (.BL(BL101),.BLN(BLN101),.WL(WL212));
sram_cell_6t_5 inst_cell_212_102 (.BL(BL102),.BLN(BLN102),.WL(WL212));
sram_cell_6t_5 inst_cell_212_103 (.BL(BL103),.BLN(BLN103),.WL(WL212));
sram_cell_6t_5 inst_cell_212_104 (.BL(BL104),.BLN(BLN104),.WL(WL212));
sram_cell_6t_5 inst_cell_212_105 (.BL(BL105),.BLN(BLN105),.WL(WL212));
sram_cell_6t_5 inst_cell_212_106 (.BL(BL106),.BLN(BLN106),.WL(WL212));
sram_cell_6t_5 inst_cell_212_107 (.BL(BL107),.BLN(BLN107),.WL(WL212));
sram_cell_6t_5 inst_cell_212_108 (.BL(BL108),.BLN(BLN108),.WL(WL212));
sram_cell_6t_5 inst_cell_212_109 (.BL(BL109),.BLN(BLN109),.WL(WL212));
sram_cell_6t_5 inst_cell_212_110 (.BL(BL110),.BLN(BLN110),.WL(WL212));
sram_cell_6t_5 inst_cell_212_111 (.BL(BL111),.BLN(BLN111),.WL(WL212));
sram_cell_6t_5 inst_cell_212_112 (.BL(BL112),.BLN(BLN112),.WL(WL212));
sram_cell_6t_5 inst_cell_212_113 (.BL(BL113),.BLN(BLN113),.WL(WL212));
sram_cell_6t_5 inst_cell_212_114 (.BL(BL114),.BLN(BLN114),.WL(WL212));
sram_cell_6t_5 inst_cell_212_115 (.BL(BL115),.BLN(BLN115),.WL(WL212));
sram_cell_6t_5 inst_cell_212_116 (.BL(BL116),.BLN(BLN116),.WL(WL212));
sram_cell_6t_5 inst_cell_212_117 (.BL(BL117),.BLN(BLN117),.WL(WL212));
sram_cell_6t_5 inst_cell_212_118 (.BL(BL118),.BLN(BLN118),.WL(WL212));
sram_cell_6t_5 inst_cell_212_119 (.BL(BL119),.BLN(BLN119),.WL(WL212));
sram_cell_6t_5 inst_cell_212_120 (.BL(BL120),.BLN(BLN120),.WL(WL212));
sram_cell_6t_5 inst_cell_212_121 (.BL(BL121),.BLN(BLN121),.WL(WL212));
sram_cell_6t_5 inst_cell_212_122 (.BL(BL122),.BLN(BLN122),.WL(WL212));
sram_cell_6t_5 inst_cell_212_123 (.BL(BL123),.BLN(BLN123),.WL(WL212));
sram_cell_6t_5 inst_cell_212_124 (.BL(BL124),.BLN(BLN124),.WL(WL212));
sram_cell_6t_5 inst_cell_212_125 (.BL(BL125),.BLN(BLN125),.WL(WL212));
sram_cell_6t_5 inst_cell_212_126 (.BL(BL126),.BLN(BLN126),.WL(WL212));
sram_cell_6t_5 inst_cell_212_127 (.BL(BL127),.BLN(BLN127),.WL(WL212));
sram_cell_6t_5 inst_cell_213_0 (.BL(BL0),.BLN(BLN0),.WL(WL213));
sram_cell_6t_5 inst_cell_213_1 (.BL(BL1),.BLN(BLN1),.WL(WL213));
sram_cell_6t_5 inst_cell_213_2 (.BL(BL2),.BLN(BLN2),.WL(WL213));
sram_cell_6t_5 inst_cell_213_3 (.BL(BL3),.BLN(BLN3),.WL(WL213));
sram_cell_6t_5 inst_cell_213_4 (.BL(BL4),.BLN(BLN4),.WL(WL213));
sram_cell_6t_5 inst_cell_213_5 (.BL(BL5),.BLN(BLN5),.WL(WL213));
sram_cell_6t_5 inst_cell_213_6 (.BL(BL6),.BLN(BLN6),.WL(WL213));
sram_cell_6t_5 inst_cell_213_7 (.BL(BL7),.BLN(BLN7),.WL(WL213));
sram_cell_6t_5 inst_cell_213_8 (.BL(BL8),.BLN(BLN8),.WL(WL213));
sram_cell_6t_5 inst_cell_213_9 (.BL(BL9),.BLN(BLN9),.WL(WL213));
sram_cell_6t_5 inst_cell_213_10 (.BL(BL10),.BLN(BLN10),.WL(WL213));
sram_cell_6t_5 inst_cell_213_11 (.BL(BL11),.BLN(BLN11),.WL(WL213));
sram_cell_6t_5 inst_cell_213_12 (.BL(BL12),.BLN(BLN12),.WL(WL213));
sram_cell_6t_5 inst_cell_213_13 (.BL(BL13),.BLN(BLN13),.WL(WL213));
sram_cell_6t_5 inst_cell_213_14 (.BL(BL14),.BLN(BLN14),.WL(WL213));
sram_cell_6t_5 inst_cell_213_15 (.BL(BL15),.BLN(BLN15),.WL(WL213));
sram_cell_6t_5 inst_cell_213_16 (.BL(BL16),.BLN(BLN16),.WL(WL213));
sram_cell_6t_5 inst_cell_213_17 (.BL(BL17),.BLN(BLN17),.WL(WL213));
sram_cell_6t_5 inst_cell_213_18 (.BL(BL18),.BLN(BLN18),.WL(WL213));
sram_cell_6t_5 inst_cell_213_19 (.BL(BL19),.BLN(BLN19),.WL(WL213));
sram_cell_6t_5 inst_cell_213_20 (.BL(BL20),.BLN(BLN20),.WL(WL213));
sram_cell_6t_5 inst_cell_213_21 (.BL(BL21),.BLN(BLN21),.WL(WL213));
sram_cell_6t_5 inst_cell_213_22 (.BL(BL22),.BLN(BLN22),.WL(WL213));
sram_cell_6t_5 inst_cell_213_23 (.BL(BL23),.BLN(BLN23),.WL(WL213));
sram_cell_6t_5 inst_cell_213_24 (.BL(BL24),.BLN(BLN24),.WL(WL213));
sram_cell_6t_5 inst_cell_213_25 (.BL(BL25),.BLN(BLN25),.WL(WL213));
sram_cell_6t_5 inst_cell_213_26 (.BL(BL26),.BLN(BLN26),.WL(WL213));
sram_cell_6t_5 inst_cell_213_27 (.BL(BL27),.BLN(BLN27),.WL(WL213));
sram_cell_6t_5 inst_cell_213_28 (.BL(BL28),.BLN(BLN28),.WL(WL213));
sram_cell_6t_5 inst_cell_213_29 (.BL(BL29),.BLN(BLN29),.WL(WL213));
sram_cell_6t_5 inst_cell_213_30 (.BL(BL30),.BLN(BLN30),.WL(WL213));
sram_cell_6t_5 inst_cell_213_31 (.BL(BL31),.BLN(BLN31),.WL(WL213));
sram_cell_6t_5 inst_cell_213_32 (.BL(BL32),.BLN(BLN32),.WL(WL213));
sram_cell_6t_5 inst_cell_213_33 (.BL(BL33),.BLN(BLN33),.WL(WL213));
sram_cell_6t_5 inst_cell_213_34 (.BL(BL34),.BLN(BLN34),.WL(WL213));
sram_cell_6t_5 inst_cell_213_35 (.BL(BL35),.BLN(BLN35),.WL(WL213));
sram_cell_6t_5 inst_cell_213_36 (.BL(BL36),.BLN(BLN36),.WL(WL213));
sram_cell_6t_5 inst_cell_213_37 (.BL(BL37),.BLN(BLN37),.WL(WL213));
sram_cell_6t_5 inst_cell_213_38 (.BL(BL38),.BLN(BLN38),.WL(WL213));
sram_cell_6t_5 inst_cell_213_39 (.BL(BL39),.BLN(BLN39),.WL(WL213));
sram_cell_6t_5 inst_cell_213_40 (.BL(BL40),.BLN(BLN40),.WL(WL213));
sram_cell_6t_5 inst_cell_213_41 (.BL(BL41),.BLN(BLN41),.WL(WL213));
sram_cell_6t_5 inst_cell_213_42 (.BL(BL42),.BLN(BLN42),.WL(WL213));
sram_cell_6t_5 inst_cell_213_43 (.BL(BL43),.BLN(BLN43),.WL(WL213));
sram_cell_6t_5 inst_cell_213_44 (.BL(BL44),.BLN(BLN44),.WL(WL213));
sram_cell_6t_5 inst_cell_213_45 (.BL(BL45),.BLN(BLN45),.WL(WL213));
sram_cell_6t_5 inst_cell_213_46 (.BL(BL46),.BLN(BLN46),.WL(WL213));
sram_cell_6t_5 inst_cell_213_47 (.BL(BL47),.BLN(BLN47),.WL(WL213));
sram_cell_6t_5 inst_cell_213_48 (.BL(BL48),.BLN(BLN48),.WL(WL213));
sram_cell_6t_5 inst_cell_213_49 (.BL(BL49),.BLN(BLN49),.WL(WL213));
sram_cell_6t_5 inst_cell_213_50 (.BL(BL50),.BLN(BLN50),.WL(WL213));
sram_cell_6t_5 inst_cell_213_51 (.BL(BL51),.BLN(BLN51),.WL(WL213));
sram_cell_6t_5 inst_cell_213_52 (.BL(BL52),.BLN(BLN52),.WL(WL213));
sram_cell_6t_5 inst_cell_213_53 (.BL(BL53),.BLN(BLN53),.WL(WL213));
sram_cell_6t_5 inst_cell_213_54 (.BL(BL54),.BLN(BLN54),.WL(WL213));
sram_cell_6t_5 inst_cell_213_55 (.BL(BL55),.BLN(BLN55),.WL(WL213));
sram_cell_6t_5 inst_cell_213_56 (.BL(BL56),.BLN(BLN56),.WL(WL213));
sram_cell_6t_5 inst_cell_213_57 (.BL(BL57),.BLN(BLN57),.WL(WL213));
sram_cell_6t_5 inst_cell_213_58 (.BL(BL58),.BLN(BLN58),.WL(WL213));
sram_cell_6t_5 inst_cell_213_59 (.BL(BL59),.BLN(BLN59),.WL(WL213));
sram_cell_6t_5 inst_cell_213_60 (.BL(BL60),.BLN(BLN60),.WL(WL213));
sram_cell_6t_5 inst_cell_213_61 (.BL(BL61),.BLN(BLN61),.WL(WL213));
sram_cell_6t_5 inst_cell_213_62 (.BL(BL62),.BLN(BLN62),.WL(WL213));
sram_cell_6t_5 inst_cell_213_63 (.BL(BL63),.BLN(BLN63),.WL(WL213));
sram_cell_6t_5 inst_cell_213_64 (.BL(BL64),.BLN(BLN64),.WL(WL213));
sram_cell_6t_5 inst_cell_213_65 (.BL(BL65),.BLN(BLN65),.WL(WL213));
sram_cell_6t_5 inst_cell_213_66 (.BL(BL66),.BLN(BLN66),.WL(WL213));
sram_cell_6t_5 inst_cell_213_67 (.BL(BL67),.BLN(BLN67),.WL(WL213));
sram_cell_6t_5 inst_cell_213_68 (.BL(BL68),.BLN(BLN68),.WL(WL213));
sram_cell_6t_5 inst_cell_213_69 (.BL(BL69),.BLN(BLN69),.WL(WL213));
sram_cell_6t_5 inst_cell_213_70 (.BL(BL70),.BLN(BLN70),.WL(WL213));
sram_cell_6t_5 inst_cell_213_71 (.BL(BL71),.BLN(BLN71),.WL(WL213));
sram_cell_6t_5 inst_cell_213_72 (.BL(BL72),.BLN(BLN72),.WL(WL213));
sram_cell_6t_5 inst_cell_213_73 (.BL(BL73),.BLN(BLN73),.WL(WL213));
sram_cell_6t_5 inst_cell_213_74 (.BL(BL74),.BLN(BLN74),.WL(WL213));
sram_cell_6t_5 inst_cell_213_75 (.BL(BL75),.BLN(BLN75),.WL(WL213));
sram_cell_6t_5 inst_cell_213_76 (.BL(BL76),.BLN(BLN76),.WL(WL213));
sram_cell_6t_5 inst_cell_213_77 (.BL(BL77),.BLN(BLN77),.WL(WL213));
sram_cell_6t_5 inst_cell_213_78 (.BL(BL78),.BLN(BLN78),.WL(WL213));
sram_cell_6t_5 inst_cell_213_79 (.BL(BL79),.BLN(BLN79),.WL(WL213));
sram_cell_6t_5 inst_cell_213_80 (.BL(BL80),.BLN(BLN80),.WL(WL213));
sram_cell_6t_5 inst_cell_213_81 (.BL(BL81),.BLN(BLN81),.WL(WL213));
sram_cell_6t_5 inst_cell_213_82 (.BL(BL82),.BLN(BLN82),.WL(WL213));
sram_cell_6t_5 inst_cell_213_83 (.BL(BL83),.BLN(BLN83),.WL(WL213));
sram_cell_6t_5 inst_cell_213_84 (.BL(BL84),.BLN(BLN84),.WL(WL213));
sram_cell_6t_5 inst_cell_213_85 (.BL(BL85),.BLN(BLN85),.WL(WL213));
sram_cell_6t_5 inst_cell_213_86 (.BL(BL86),.BLN(BLN86),.WL(WL213));
sram_cell_6t_5 inst_cell_213_87 (.BL(BL87),.BLN(BLN87),.WL(WL213));
sram_cell_6t_5 inst_cell_213_88 (.BL(BL88),.BLN(BLN88),.WL(WL213));
sram_cell_6t_5 inst_cell_213_89 (.BL(BL89),.BLN(BLN89),.WL(WL213));
sram_cell_6t_5 inst_cell_213_90 (.BL(BL90),.BLN(BLN90),.WL(WL213));
sram_cell_6t_5 inst_cell_213_91 (.BL(BL91),.BLN(BLN91),.WL(WL213));
sram_cell_6t_5 inst_cell_213_92 (.BL(BL92),.BLN(BLN92),.WL(WL213));
sram_cell_6t_5 inst_cell_213_93 (.BL(BL93),.BLN(BLN93),.WL(WL213));
sram_cell_6t_5 inst_cell_213_94 (.BL(BL94),.BLN(BLN94),.WL(WL213));
sram_cell_6t_5 inst_cell_213_95 (.BL(BL95),.BLN(BLN95),.WL(WL213));
sram_cell_6t_5 inst_cell_213_96 (.BL(BL96),.BLN(BLN96),.WL(WL213));
sram_cell_6t_5 inst_cell_213_97 (.BL(BL97),.BLN(BLN97),.WL(WL213));
sram_cell_6t_5 inst_cell_213_98 (.BL(BL98),.BLN(BLN98),.WL(WL213));
sram_cell_6t_5 inst_cell_213_99 (.BL(BL99),.BLN(BLN99),.WL(WL213));
sram_cell_6t_5 inst_cell_213_100 (.BL(BL100),.BLN(BLN100),.WL(WL213));
sram_cell_6t_5 inst_cell_213_101 (.BL(BL101),.BLN(BLN101),.WL(WL213));
sram_cell_6t_5 inst_cell_213_102 (.BL(BL102),.BLN(BLN102),.WL(WL213));
sram_cell_6t_5 inst_cell_213_103 (.BL(BL103),.BLN(BLN103),.WL(WL213));
sram_cell_6t_5 inst_cell_213_104 (.BL(BL104),.BLN(BLN104),.WL(WL213));
sram_cell_6t_5 inst_cell_213_105 (.BL(BL105),.BLN(BLN105),.WL(WL213));
sram_cell_6t_5 inst_cell_213_106 (.BL(BL106),.BLN(BLN106),.WL(WL213));
sram_cell_6t_5 inst_cell_213_107 (.BL(BL107),.BLN(BLN107),.WL(WL213));
sram_cell_6t_5 inst_cell_213_108 (.BL(BL108),.BLN(BLN108),.WL(WL213));
sram_cell_6t_5 inst_cell_213_109 (.BL(BL109),.BLN(BLN109),.WL(WL213));
sram_cell_6t_5 inst_cell_213_110 (.BL(BL110),.BLN(BLN110),.WL(WL213));
sram_cell_6t_5 inst_cell_213_111 (.BL(BL111),.BLN(BLN111),.WL(WL213));
sram_cell_6t_5 inst_cell_213_112 (.BL(BL112),.BLN(BLN112),.WL(WL213));
sram_cell_6t_5 inst_cell_213_113 (.BL(BL113),.BLN(BLN113),.WL(WL213));
sram_cell_6t_5 inst_cell_213_114 (.BL(BL114),.BLN(BLN114),.WL(WL213));
sram_cell_6t_5 inst_cell_213_115 (.BL(BL115),.BLN(BLN115),.WL(WL213));
sram_cell_6t_5 inst_cell_213_116 (.BL(BL116),.BLN(BLN116),.WL(WL213));
sram_cell_6t_5 inst_cell_213_117 (.BL(BL117),.BLN(BLN117),.WL(WL213));
sram_cell_6t_5 inst_cell_213_118 (.BL(BL118),.BLN(BLN118),.WL(WL213));
sram_cell_6t_5 inst_cell_213_119 (.BL(BL119),.BLN(BLN119),.WL(WL213));
sram_cell_6t_5 inst_cell_213_120 (.BL(BL120),.BLN(BLN120),.WL(WL213));
sram_cell_6t_5 inst_cell_213_121 (.BL(BL121),.BLN(BLN121),.WL(WL213));
sram_cell_6t_5 inst_cell_213_122 (.BL(BL122),.BLN(BLN122),.WL(WL213));
sram_cell_6t_5 inst_cell_213_123 (.BL(BL123),.BLN(BLN123),.WL(WL213));
sram_cell_6t_5 inst_cell_213_124 (.BL(BL124),.BLN(BLN124),.WL(WL213));
sram_cell_6t_5 inst_cell_213_125 (.BL(BL125),.BLN(BLN125),.WL(WL213));
sram_cell_6t_5 inst_cell_213_126 (.BL(BL126),.BLN(BLN126),.WL(WL213));
sram_cell_6t_5 inst_cell_213_127 (.BL(BL127),.BLN(BLN127),.WL(WL213));
sram_cell_6t_5 inst_cell_214_0 (.BL(BL0),.BLN(BLN0),.WL(WL214));
sram_cell_6t_5 inst_cell_214_1 (.BL(BL1),.BLN(BLN1),.WL(WL214));
sram_cell_6t_5 inst_cell_214_2 (.BL(BL2),.BLN(BLN2),.WL(WL214));
sram_cell_6t_5 inst_cell_214_3 (.BL(BL3),.BLN(BLN3),.WL(WL214));
sram_cell_6t_5 inst_cell_214_4 (.BL(BL4),.BLN(BLN4),.WL(WL214));
sram_cell_6t_5 inst_cell_214_5 (.BL(BL5),.BLN(BLN5),.WL(WL214));
sram_cell_6t_5 inst_cell_214_6 (.BL(BL6),.BLN(BLN6),.WL(WL214));
sram_cell_6t_5 inst_cell_214_7 (.BL(BL7),.BLN(BLN7),.WL(WL214));
sram_cell_6t_5 inst_cell_214_8 (.BL(BL8),.BLN(BLN8),.WL(WL214));
sram_cell_6t_5 inst_cell_214_9 (.BL(BL9),.BLN(BLN9),.WL(WL214));
sram_cell_6t_5 inst_cell_214_10 (.BL(BL10),.BLN(BLN10),.WL(WL214));
sram_cell_6t_5 inst_cell_214_11 (.BL(BL11),.BLN(BLN11),.WL(WL214));
sram_cell_6t_5 inst_cell_214_12 (.BL(BL12),.BLN(BLN12),.WL(WL214));
sram_cell_6t_5 inst_cell_214_13 (.BL(BL13),.BLN(BLN13),.WL(WL214));
sram_cell_6t_5 inst_cell_214_14 (.BL(BL14),.BLN(BLN14),.WL(WL214));
sram_cell_6t_5 inst_cell_214_15 (.BL(BL15),.BLN(BLN15),.WL(WL214));
sram_cell_6t_5 inst_cell_214_16 (.BL(BL16),.BLN(BLN16),.WL(WL214));
sram_cell_6t_5 inst_cell_214_17 (.BL(BL17),.BLN(BLN17),.WL(WL214));
sram_cell_6t_5 inst_cell_214_18 (.BL(BL18),.BLN(BLN18),.WL(WL214));
sram_cell_6t_5 inst_cell_214_19 (.BL(BL19),.BLN(BLN19),.WL(WL214));
sram_cell_6t_5 inst_cell_214_20 (.BL(BL20),.BLN(BLN20),.WL(WL214));
sram_cell_6t_5 inst_cell_214_21 (.BL(BL21),.BLN(BLN21),.WL(WL214));
sram_cell_6t_5 inst_cell_214_22 (.BL(BL22),.BLN(BLN22),.WL(WL214));
sram_cell_6t_5 inst_cell_214_23 (.BL(BL23),.BLN(BLN23),.WL(WL214));
sram_cell_6t_5 inst_cell_214_24 (.BL(BL24),.BLN(BLN24),.WL(WL214));
sram_cell_6t_5 inst_cell_214_25 (.BL(BL25),.BLN(BLN25),.WL(WL214));
sram_cell_6t_5 inst_cell_214_26 (.BL(BL26),.BLN(BLN26),.WL(WL214));
sram_cell_6t_5 inst_cell_214_27 (.BL(BL27),.BLN(BLN27),.WL(WL214));
sram_cell_6t_5 inst_cell_214_28 (.BL(BL28),.BLN(BLN28),.WL(WL214));
sram_cell_6t_5 inst_cell_214_29 (.BL(BL29),.BLN(BLN29),.WL(WL214));
sram_cell_6t_5 inst_cell_214_30 (.BL(BL30),.BLN(BLN30),.WL(WL214));
sram_cell_6t_5 inst_cell_214_31 (.BL(BL31),.BLN(BLN31),.WL(WL214));
sram_cell_6t_5 inst_cell_214_32 (.BL(BL32),.BLN(BLN32),.WL(WL214));
sram_cell_6t_5 inst_cell_214_33 (.BL(BL33),.BLN(BLN33),.WL(WL214));
sram_cell_6t_5 inst_cell_214_34 (.BL(BL34),.BLN(BLN34),.WL(WL214));
sram_cell_6t_5 inst_cell_214_35 (.BL(BL35),.BLN(BLN35),.WL(WL214));
sram_cell_6t_5 inst_cell_214_36 (.BL(BL36),.BLN(BLN36),.WL(WL214));
sram_cell_6t_5 inst_cell_214_37 (.BL(BL37),.BLN(BLN37),.WL(WL214));
sram_cell_6t_5 inst_cell_214_38 (.BL(BL38),.BLN(BLN38),.WL(WL214));
sram_cell_6t_5 inst_cell_214_39 (.BL(BL39),.BLN(BLN39),.WL(WL214));
sram_cell_6t_5 inst_cell_214_40 (.BL(BL40),.BLN(BLN40),.WL(WL214));
sram_cell_6t_5 inst_cell_214_41 (.BL(BL41),.BLN(BLN41),.WL(WL214));
sram_cell_6t_5 inst_cell_214_42 (.BL(BL42),.BLN(BLN42),.WL(WL214));
sram_cell_6t_5 inst_cell_214_43 (.BL(BL43),.BLN(BLN43),.WL(WL214));
sram_cell_6t_5 inst_cell_214_44 (.BL(BL44),.BLN(BLN44),.WL(WL214));
sram_cell_6t_5 inst_cell_214_45 (.BL(BL45),.BLN(BLN45),.WL(WL214));
sram_cell_6t_5 inst_cell_214_46 (.BL(BL46),.BLN(BLN46),.WL(WL214));
sram_cell_6t_5 inst_cell_214_47 (.BL(BL47),.BLN(BLN47),.WL(WL214));
sram_cell_6t_5 inst_cell_214_48 (.BL(BL48),.BLN(BLN48),.WL(WL214));
sram_cell_6t_5 inst_cell_214_49 (.BL(BL49),.BLN(BLN49),.WL(WL214));
sram_cell_6t_5 inst_cell_214_50 (.BL(BL50),.BLN(BLN50),.WL(WL214));
sram_cell_6t_5 inst_cell_214_51 (.BL(BL51),.BLN(BLN51),.WL(WL214));
sram_cell_6t_5 inst_cell_214_52 (.BL(BL52),.BLN(BLN52),.WL(WL214));
sram_cell_6t_5 inst_cell_214_53 (.BL(BL53),.BLN(BLN53),.WL(WL214));
sram_cell_6t_5 inst_cell_214_54 (.BL(BL54),.BLN(BLN54),.WL(WL214));
sram_cell_6t_5 inst_cell_214_55 (.BL(BL55),.BLN(BLN55),.WL(WL214));
sram_cell_6t_5 inst_cell_214_56 (.BL(BL56),.BLN(BLN56),.WL(WL214));
sram_cell_6t_5 inst_cell_214_57 (.BL(BL57),.BLN(BLN57),.WL(WL214));
sram_cell_6t_5 inst_cell_214_58 (.BL(BL58),.BLN(BLN58),.WL(WL214));
sram_cell_6t_5 inst_cell_214_59 (.BL(BL59),.BLN(BLN59),.WL(WL214));
sram_cell_6t_5 inst_cell_214_60 (.BL(BL60),.BLN(BLN60),.WL(WL214));
sram_cell_6t_5 inst_cell_214_61 (.BL(BL61),.BLN(BLN61),.WL(WL214));
sram_cell_6t_5 inst_cell_214_62 (.BL(BL62),.BLN(BLN62),.WL(WL214));
sram_cell_6t_5 inst_cell_214_63 (.BL(BL63),.BLN(BLN63),.WL(WL214));
sram_cell_6t_5 inst_cell_214_64 (.BL(BL64),.BLN(BLN64),.WL(WL214));
sram_cell_6t_5 inst_cell_214_65 (.BL(BL65),.BLN(BLN65),.WL(WL214));
sram_cell_6t_5 inst_cell_214_66 (.BL(BL66),.BLN(BLN66),.WL(WL214));
sram_cell_6t_5 inst_cell_214_67 (.BL(BL67),.BLN(BLN67),.WL(WL214));
sram_cell_6t_5 inst_cell_214_68 (.BL(BL68),.BLN(BLN68),.WL(WL214));
sram_cell_6t_5 inst_cell_214_69 (.BL(BL69),.BLN(BLN69),.WL(WL214));
sram_cell_6t_5 inst_cell_214_70 (.BL(BL70),.BLN(BLN70),.WL(WL214));
sram_cell_6t_5 inst_cell_214_71 (.BL(BL71),.BLN(BLN71),.WL(WL214));
sram_cell_6t_5 inst_cell_214_72 (.BL(BL72),.BLN(BLN72),.WL(WL214));
sram_cell_6t_5 inst_cell_214_73 (.BL(BL73),.BLN(BLN73),.WL(WL214));
sram_cell_6t_5 inst_cell_214_74 (.BL(BL74),.BLN(BLN74),.WL(WL214));
sram_cell_6t_5 inst_cell_214_75 (.BL(BL75),.BLN(BLN75),.WL(WL214));
sram_cell_6t_5 inst_cell_214_76 (.BL(BL76),.BLN(BLN76),.WL(WL214));
sram_cell_6t_5 inst_cell_214_77 (.BL(BL77),.BLN(BLN77),.WL(WL214));
sram_cell_6t_5 inst_cell_214_78 (.BL(BL78),.BLN(BLN78),.WL(WL214));
sram_cell_6t_5 inst_cell_214_79 (.BL(BL79),.BLN(BLN79),.WL(WL214));
sram_cell_6t_5 inst_cell_214_80 (.BL(BL80),.BLN(BLN80),.WL(WL214));
sram_cell_6t_5 inst_cell_214_81 (.BL(BL81),.BLN(BLN81),.WL(WL214));
sram_cell_6t_5 inst_cell_214_82 (.BL(BL82),.BLN(BLN82),.WL(WL214));
sram_cell_6t_5 inst_cell_214_83 (.BL(BL83),.BLN(BLN83),.WL(WL214));
sram_cell_6t_5 inst_cell_214_84 (.BL(BL84),.BLN(BLN84),.WL(WL214));
sram_cell_6t_5 inst_cell_214_85 (.BL(BL85),.BLN(BLN85),.WL(WL214));
sram_cell_6t_5 inst_cell_214_86 (.BL(BL86),.BLN(BLN86),.WL(WL214));
sram_cell_6t_5 inst_cell_214_87 (.BL(BL87),.BLN(BLN87),.WL(WL214));
sram_cell_6t_5 inst_cell_214_88 (.BL(BL88),.BLN(BLN88),.WL(WL214));
sram_cell_6t_5 inst_cell_214_89 (.BL(BL89),.BLN(BLN89),.WL(WL214));
sram_cell_6t_5 inst_cell_214_90 (.BL(BL90),.BLN(BLN90),.WL(WL214));
sram_cell_6t_5 inst_cell_214_91 (.BL(BL91),.BLN(BLN91),.WL(WL214));
sram_cell_6t_5 inst_cell_214_92 (.BL(BL92),.BLN(BLN92),.WL(WL214));
sram_cell_6t_5 inst_cell_214_93 (.BL(BL93),.BLN(BLN93),.WL(WL214));
sram_cell_6t_5 inst_cell_214_94 (.BL(BL94),.BLN(BLN94),.WL(WL214));
sram_cell_6t_5 inst_cell_214_95 (.BL(BL95),.BLN(BLN95),.WL(WL214));
sram_cell_6t_5 inst_cell_214_96 (.BL(BL96),.BLN(BLN96),.WL(WL214));
sram_cell_6t_5 inst_cell_214_97 (.BL(BL97),.BLN(BLN97),.WL(WL214));
sram_cell_6t_5 inst_cell_214_98 (.BL(BL98),.BLN(BLN98),.WL(WL214));
sram_cell_6t_5 inst_cell_214_99 (.BL(BL99),.BLN(BLN99),.WL(WL214));
sram_cell_6t_5 inst_cell_214_100 (.BL(BL100),.BLN(BLN100),.WL(WL214));
sram_cell_6t_5 inst_cell_214_101 (.BL(BL101),.BLN(BLN101),.WL(WL214));
sram_cell_6t_5 inst_cell_214_102 (.BL(BL102),.BLN(BLN102),.WL(WL214));
sram_cell_6t_5 inst_cell_214_103 (.BL(BL103),.BLN(BLN103),.WL(WL214));
sram_cell_6t_5 inst_cell_214_104 (.BL(BL104),.BLN(BLN104),.WL(WL214));
sram_cell_6t_5 inst_cell_214_105 (.BL(BL105),.BLN(BLN105),.WL(WL214));
sram_cell_6t_5 inst_cell_214_106 (.BL(BL106),.BLN(BLN106),.WL(WL214));
sram_cell_6t_5 inst_cell_214_107 (.BL(BL107),.BLN(BLN107),.WL(WL214));
sram_cell_6t_5 inst_cell_214_108 (.BL(BL108),.BLN(BLN108),.WL(WL214));
sram_cell_6t_5 inst_cell_214_109 (.BL(BL109),.BLN(BLN109),.WL(WL214));
sram_cell_6t_5 inst_cell_214_110 (.BL(BL110),.BLN(BLN110),.WL(WL214));
sram_cell_6t_5 inst_cell_214_111 (.BL(BL111),.BLN(BLN111),.WL(WL214));
sram_cell_6t_5 inst_cell_214_112 (.BL(BL112),.BLN(BLN112),.WL(WL214));
sram_cell_6t_5 inst_cell_214_113 (.BL(BL113),.BLN(BLN113),.WL(WL214));
sram_cell_6t_5 inst_cell_214_114 (.BL(BL114),.BLN(BLN114),.WL(WL214));
sram_cell_6t_5 inst_cell_214_115 (.BL(BL115),.BLN(BLN115),.WL(WL214));
sram_cell_6t_5 inst_cell_214_116 (.BL(BL116),.BLN(BLN116),.WL(WL214));
sram_cell_6t_5 inst_cell_214_117 (.BL(BL117),.BLN(BLN117),.WL(WL214));
sram_cell_6t_5 inst_cell_214_118 (.BL(BL118),.BLN(BLN118),.WL(WL214));
sram_cell_6t_5 inst_cell_214_119 (.BL(BL119),.BLN(BLN119),.WL(WL214));
sram_cell_6t_5 inst_cell_214_120 (.BL(BL120),.BLN(BLN120),.WL(WL214));
sram_cell_6t_5 inst_cell_214_121 (.BL(BL121),.BLN(BLN121),.WL(WL214));
sram_cell_6t_5 inst_cell_214_122 (.BL(BL122),.BLN(BLN122),.WL(WL214));
sram_cell_6t_5 inst_cell_214_123 (.BL(BL123),.BLN(BLN123),.WL(WL214));
sram_cell_6t_5 inst_cell_214_124 (.BL(BL124),.BLN(BLN124),.WL(WL214));
sram_cell_6t_5 inst_cell_214_125 (.BL(BL125),.BLN(BLN125),.WL(WL214));
sram_cell_6t_5 inst_cell_214_126 (.BL(BL126),.BLN(BLN126),.WL(WL214));
sram_cell_6t_5 inst_cell_214_127 (.BL(BL127),.BLN(BLN127),.WL(WL214));
sram_cell_6t_5 inst_cell_215_0 (.BL(BL0),.BLN(BLN0),.WL(WL215));
sram_cell_6t_5 inst_cell_215_1 (.BL(BL1),.BLN(BLN1),.WL(WL215));
sram_cell_6t_5 inst_cell_215_2 (.BL(BL2),.BLN(BLN2),.WL(WL215));
sram_cell_6t_5 inst_cell_215_3 (.BL(BL3),.BLN(BLN3),.WL(WL215));
sram_cell_6t_5 inst_cell_215_4 (.BL(BL4),.BLN(BLN4),.WL(WL215));
sram_cell_6t_5 inst_cell_215_5 (.BL(BL5),.BLN(BLN5),.WL(WL215));
sram_cell_6t_5 inst_cell_215_6 (.BL(BL6),.BLN(BLN6),.WL(WL215));
sram_cell_6t_5 inst_cell_215_7 (.BL(BL7),.BLN(BLN7),.WL(WL215));
sram_cell_6t_5 inst_cell_215_8 (.BL(BL8),.BLN(BLN8),.WL(WL215));
sram_cell_6t_5 inst_cell_215_9 (.BL(BL9),.BLN(BLN9),.WL(WL215));
sram_cell_6t_5 inst_cell_215_10 (.BL(BL10),.BLN(BLN10),.WL(WL215));
sram_cell_6t_5 inst_cell_215_11 (.BL(BL11),.BLN(BLN11),.WL(WL215));
sram_cell_6t_5 inst_cell_215_12 (.BL(BL12),.BLN(BLN12),.WL(WL215));
sram_cell_6t_5 inst_cell_215_13 (.BL(BL13),.BLN(BLN13),.WL(WL215));
sram_cell_6t_5 inst_cell_215_14 (.BL(BL14),.BLN(BLN14),.WL(WL215));
sram_cell_6t_5 inst_cell_215_15 (.BL(BL15),.BLN(BLN15),.WL(WL215));
sram_cell_6t_5 inst_cell_215_16 (.BL(BL16),.BLN(BLN16),.WL(WL215));
sram_cell_6t_5 inst_cell_215_17 (.BL(BL17),.BLN(BLN17),.WL(WL215));
sram_cell_6t_5 inst_cell_215_18 (.BL(BL18),.BLN(BLN18),.WL(WL215));
sram_cell_6t_5 inst_cell_215_19 (.BL(BL19),.BLN(BLN19),.WL(WL215));
sram_cell_6t_5 inst_cell_215_20 (.BL(BL20),.BLN(BLN20),.WL(WL215));
sram_cell_6t_5 inst_cell_215_21 (.BL(BL21),.BLN(BLN21),.WL(WL215));
sram_cell_6t_5 inst_cell_215_22 (.BL(BL22),.BLN(BLN22),.WL(WL215));
sram_cell_6t_5 inst_cell_215_23 (.BL(BL23),.BLN(BLN23),.WL(WL215));
sram_cell_6t_5 inst_cell_215_24 (.BL(BL24),.BLN(BLN24),.WL(WL215));
sram_cell_6t_5 inst_cell_215_25 (.BL(BL25),.BLN(BLN25),.WL(WL215));
sram_cell_6t_5 inst_cell_215_26 (.BL(BL26),.BLN(BLN26),.WL(WL215));
sram_cell_6t_5 inst_cell_215_27 (.BL(BL27),.BLN(BLN27),.WL(WL215));
sram_cell_6t_5 inst_cell_215_28 (.BL(BL28),.BLN(BLN28),.WL(WL215));
sram_cell_6t_5 inst_cell_215_29 (.BL(BL29),.BLN(BLN29),.WL(WL215));
sram_cell_6t_5 inst_cell_215_30 (.BL(BL30),.BLN(BLN30),.WL(WL215));
sram_cell_6t_5 inst_cell_215_31 (.BL(BL31),.BLN(BLN31),.WL(WL215));
sram_cell_6t_5 inst_cell_215_32 (.BL(BL32),.BLN(BLN32),.WL(WL215));
sram_cell_6t_5 inst_cell_215_33 (.BL(BL33),.BLN(BLN33),.WL(WL215));
sram_cell_6t_5 inst_cell_215_34 (.BL(BL34),.BLN(BLN34),.WL(WL215));
sram_cell_6t_5 inst_cell_215_35 (.BL(BL35),.BLN(BLN35),.WL(WL215));
sram_cell_6t_5 inst_cell_215_36 (.BL(BL36),.BLN(BLN36),.WL(WL215));
sram_cell_6t_5 inst_cell_215_37 (.BL(BL37),.BLN(BLN37),.WL(WL215));
sram_cell_6t_5 inst_cell_215_38 (.BL(BL38),.BLN(BLN38),.WL(WL215));
sram_cell_6t_5 inst_cell_215_39 (.BL(BL39),.BLN(BLN39),.WL(WL215));
sram_cell_6t_5 inst_cell_215_40 (.BL(BL40),.BLN(BLN40),.WL(WL215));
sram_cell_6t_5 inst_cell_215_41 (.BL(BL41),.BLN(BLN41),.WL(WL215));
sram_cell_6t_5 inst_cell_215_42 (.BL(BL42),.BLN(BLN42),.WL(WL215));
sram_cell_6t_5 inst_cell_215_43 (.BL(BL43),.BLN(BLN43),.WL(WL215));
sram_cell_6t_5 inst_cell_215_44 (.BL(BL44),.BLN(BLN44),.WL(WL215));
sram_cell_6t_5 inst_cell_215_45 (.BL(BL45),.BLN(BLN45),.WL(WL215));
sram_cell_6t_5 inst_cell_215_46 (.BL(BL46),.BLN(BLN46),.WL(WL215));
sram_cell_6t_5 inst_cell_215_47 (.BL(BL47),.BLN(BLN47),.WL(WL215));
sram_cell_6t_5 inst_cell_215_48 (.BL(BL48),.BLN(BLN48),.WL(WL215));
sram_cell_6t_5 inst_cell_215_49 (.BL(BL49),.BLN(BLN49),.WL(WL215));
sram_cell_6t_5 inst_cell_215_50 (.BL(BL50),.BLN(BLN50),.WL(WL215));
sram_cell_6t_5 inst_cell_215_51 (.BL(BL51),.BLN(BLN51),.WL(WL215));
sram_cell_6t_5 inst_cell_215_52 (.BL(BL52),.BLN(BLN52),.WL(WL215));
sram_cell_6t_5 inst_cell_215_53 (.BL(BL53),.BLN(BLN53),.WL(WL215));
sram_cell_6t_5 inst_cell_215_54 (.BL(BL54),.BLN(BLN54),.WL(WL215));
sram_cell_6t_5 inst_cell_215_55 (.BL(BL55),.BLN(BLN55),.WL(WL215));
sram_cell_6t_5 inst_cell_215_56 (.BL(BL56),.BLN(BLN56),.WL(WL215));
sram_cell_6t_5 inst_cell_215_57 (.BL(BL57),.BLN(BLN57),.WL(WL215));
sram_cell_6t_5 inst_cell_215_58 (.BL(BL58),.BLN(BLN58),.WL(WL215));
sram_cell_6t_5 inst_cell_215_59 (.BL(BL59),.BLN(BLN59),.WL(WL215));
sram_cell_6t_5 inst_cell_215_60 (.BL(BL60),.BLN(BLN60),.WL(WL215));
sram_cell_6t_5 inst_cell_215_61 (.BL(BL61),.BLN(BLN61),.WL(WL215));
sram_cell_6t_5 inst_cell_215_62 (.BL(BL62),.BLN(BLN62),.WL(WL215));
sram_cell_6t_5 inst_cell_215_63 (.BL(BL63),.BLN(BLN63),.WL(WL215));
sram_cell_6t_5 inst_cell_215_64 (.BL(BL64),.BLN(BLN64),.WL(WL215));
sram_cell_6t_5 inst_cell_215_65 (.BL(BL65),.BLN(BLN65),.WL(WL215));
sram_cell_6t_5 inst_cell_215_66 (.BL(BL66),.BLN(BLN66),.WL(WL215));
sram_cell_6t_5 inst_cell_215_67 (.BL(BL67),.BLN(BLN67),.WL(WL215));
sram_cell_6t_5 inst_cell_215_68 (.BL(BL68),.BLN(BLN68),.WL(WL215));
sram_cell_6t_5 inst_cell_215_69 (.BL(BL69),.BLN(BLN69),.WL(WL215));
sram_cell_6t_5 inst_cell_215_70 (.BL(BL70),.BLN(BLN70),.WL(WL215));
sram_cell_6t_5 inst_cell_215_71 (.BL(BL71),.BLN(BLN71),.WL(WL215));
sram_cell_6t_5 inst_cell_215_72 (.BL(BL72),.BLN(BLN72),.WL(WL215));
sram_cell_6t_5 inst_cell_215_73 (.BL(BL73),.BLN(BLN73),.WL(WL215));
sram_cell_6t_5 inst_cell_215_74 (.BL(BL74),.BLN(BLN74),.WL(WL215));
sram_cell_6t_5 inst_cell_215_75 (.BL(BL75),.BLN(BLN75),.WL(WL215));
sram_cell_6t_5 inst_cell_215_76 (.BL(BL76),.BLN(BLN76),.WL(WL215));
sram_cell_6t_5 inst_cell_215_77 (.BL(BL77),.BLN(BLN77),.WL(WL215));
sram_cell_6t_5 inst_cell_215_78 (.BL(BL78),.BLN(BLN78),.WL(WL215));
sram_cell_6t_5 inst_cell_215_79 (.BL(BL79),.BLN(BLN79),.WL(WL215));
sram_cell_6t_5 inst_cell_215_80 (.BL(BL80),.BLN(BLN80),.WL(WL215));
sram_cell_6t_5 inst_cell_215_81 (.BL(BL81),.BLN(BLN81),.WL(WL215));
sram_cell_6t_5 inst_cell_215_82 (.BL(BL82),.BLN(BLN82),.WL(WL215));
sram_cell_6t_5 inst_cell_215_83 (.BL(BL83),.BLN(BLN83),.WL(WL215));
sram_cell_6t_5 inst_cell_215_84 (.BL(BL84),.BLN(BLN84),.WL(WL215));
sram_cell_6t_5 inst_cell_215_85 (.BL(BL85),.BLN(BLN85),.WL(WL215));
sram_cell_6t_5 inst_cell_215_86 (.BL(BL86),.BLN(BLN86),.WL(WL215));
sram_cell_6t_5 inst_cell_215_87 (.BL(BL87),.BLN(BLN87),.WL(WL215));
sram_cell_6t_5 inst_cell_215_88 (.BL(BL88),.BLN(BLN88),.WL(WL215));
sram_cell_6t_5 inst_cell_215_89 (.BL(BL89),.BLN(BLN89),.WL(WL215));
sram_cell_6t_5 inst_cell_215_90 (.BL(BL90),.BLN(BLN90),.WL(WL215));
sram_cell_6t_5 inst_cell_215_91 (.BL(BL91),.BLN(BLN91),.WL(WL215));
sram_cell_6t_5 inst_cell_215_92 (.BL(BL92),.BLN(BLN92),.WL(WL215));
sram_cell_6t_5 inst_cell_215_93 (.BL(BL93),.BLN(BLN93),.WL(WL215));
sram_cell_6t_5 inst_cell_215_94 (.BL(BL94),.BLN(BLN94),.WL(WL215));
sram_cell_6t_5 inst_cell_215_95 (.BL(BL95),.BLN(BLN95),.WL(WL215));
sram_cell_6t_5 inst_cell_215_96 (.BL(BL96),.BLN(BLN96),.WL(WL215));
sram_cell_6t_5 inst_cell_215_97 (.BL(BL97),.BLN(BLN97),.WL(WL215));
sram_cell_6t_5 inst_cell_215_98 (.BL(BL98),.BLN(BLN98),.WL(WL215));
sram_cell_6t_5 inst_cell_215_99 (.BL(BL99),.BLN(BLN99),.WL(WL215));
sram_cell_6t_5 inst_cell_215_100 (.BL(BL100),.BLN(BLN100),.WL(WL215));
sram_cell_6t_5 inst_cell_215_101 (.BL(BL101),.BLN(BLN101),.WL(WL215));
sram_cell_6t_5 inst_cell_215_102 (.BL(BL102),.BLN(BLN102),.WL(WL215));
sram_cell_6t_5 inst_cell_215_103 (.BL(BL103),.BLN(BLN103),.WL(WL215));
sram_cell_6t_5 inst_cell_215_104 (.BL(BL104),.BLN(BLN104),.WL(WL215));
sram_cell_6t_5 inst_cell_215_105 (.BL(BL105),.BLN(BLN105),.WL(WL215));
sram_cell_6t_5 inst_cell_215_106 (.BL(BL106),.BLN(BLN106),.WL(WL215));
sram_cell_6t_5 inst_cell_215_107 (.BL(BL107),.BLN(BLN107),.WL(WL215));
sram_cell_6t_5 inst_cell_215_108 (.BL(BL108),.BLN(BLN108),.WL(WL215));
sram_cell_6t_5 inst_cell_215_109 (.BL(BL109),.BLN(BLN109),.WL(WL215));
sram_cell_6t_5 inst_cell_215_110 (.BL(BL110),.BLN(BLN110),.WL(WL215));
sram_cell_6t_5 inst_cell_215_111 (.BL(BL111),.BLN(BLN111),.WL(WL215));
sram_cell_6t_5 inst_cell_215_112 (.BL(BL112),.BLN(BLN112),.WL(WL215));
sram_cell_6t_5 inst_cell_215_113 (.BL(BL113),.BLN(BLN113),.WL(WL215));
sram_cell_6t_5 inst_cell_215_114 (.BL(BL114),.BLN(BLN114),.WL(WL215));
sram_cell_6t_5 inst_cell_215_115 (.BL(BL115),.BLN(BLN115),.WL(WL215));
sram_cell_6t_5 inst_cell_215_116 (.BL(BL116),.BLN(BLN116),.WL(WL215));
sram_cell_6t_5 inst_cell_215_117 (.BL(BL117),.BLN(BLN117),.WL(WL215));
sram_cell_6t_5 inst_cell_215_118 (.BL(BL118),.BLN(BLN118),.WL(WL215));
sram_cell_6t_5 inst_cell_215_119 (.BL(BL119),.BLN(BLN119),.WL(WL215));
sram_cell_6t_5 inst_cell_215_120 (.BL(BL120),.BLN(BLN120),.WL(WL215));
sram_cell_6t_5 inst_cell_215_121 (.BL(BL121),.BLN(BLN121),.WL(WL215));
sram_cell_6t_5 inst_cell_215_122 (.BL(BL122),.BLN(BLN122),.WL(WL215));
sram_cell_6t_5 inst_cell_215_123 (.BL(BL123),.BLN(BLN123),.WL(WL215));
sram_cell_6t_5 inst_cell_215_124 (.BL(BL124),.BLN(BLN124),.WL(WL215));
sram_cell_6t_5 inst_cell_215_125 (.BL(BL125),.BLN(BLN125),.WL(WL215));
sram_cell_6t_5 inst_cell_215_126 (.BL(BL126),.BLN(BLN126),.WL(WL215));
sram_cell_6t_5 inst_cell_215_127 (.BL(BL127),.BLN(BLN127),.WL(WL215));
sram_cell_6t_5 inst_cell_216_0 (.BL(BL0),.BLN(BLN0),.WL(WL216));
sram_cell_6t_5 inst_cell_216_1 (.BL(BL1),.BLN(BLN1),.WL(WL216));
sram_cell_6t_5 inst_cell_216_2 (.BL(BL2),.BLN(BLN2),.WL(WL216));
sram_cell_6t_5 inst_cell_216_3 (.BL(BL3),.BLN(BLN3),.WL(WL216));
sram_cell_6t_5 inst_cell_216_4 (.BL(BL4),.BLN(BLN4),.WL(WL216));
sram_cell_6t_5 inst_cell_216_5 (.BL(BL5),.BLN(BLN5),.WL(WL216));
sram_cell_6t_5 inst_cell_216_6 (.BL(BL6),.BLN(BLN6),.WL(WL216));
sram_cell_6t_5 inst_cell_216_7 (.BL(BL7),.BLN(BLN7),.WL(WL216));
sram_cell_6t_5 inst_cell_216_8 (.BL(BL8),.BLN(BLN8),.WL(WL216));
sram_cell_6t_5 inst_cell_216_9 (.BL(BL9),.BLN(BLN9),.WL(WL216));
sram_cell_6t_5 inst_cell_216_10 (.BL(BL10),.BLN(BLN10),.WL(WL216));
sram_cell_6t_5 inst_cell_216_11 (.BL(BL11),.BLN(BLN11),.WL(WL216));
sram_cell_6t_5 inst_cell_216_12 (.BL(BL12),.BLN(BLN12),.WL(WL216));
sram_cell_6t_5 inst_cell_216_13 (.BL(BL13),.BLN(BLN13),.WL(WL216));
sram_cell_6t_5 inst_cell_216_14 (.BL(BL14),.BLN(BLN14),.WL(WL216));
sram_cell_6t_5 inst_cell_216_15 (.BL(BL15),.BLN(BLN15),.WL(WL216));
sram_cell_6t_5 inst_cell_216_16 (.BL(BL16),.BLN(BLN16),.WL(WL216));
sram_cell_6t_5 inst_cell_216_17 (.BL(BL17),.BLN(BLN17),.WL(WL216));
sram_cell_6t_5 inst_cell_216_18 (.BL(BL18),.BLN(BLN18),.WL(WL216));
sram_cell_6t_5 inst_cell_216_19 (.BL(BL19),.BLN(BLN19),.WL(WL216));
sram_cell_6t_5 inst_cell_216_20 (.BL(BL20),.BLN(BLN20),.WL(WL216));
sram_cell_6t_5 inst_cell_216_21 (.BL(BL21),.BLN(BLN21),.WL(WL216));
sram_cell_6t_5 inst_cell_216_22 (.BL(BL22),.BLN(BLN22),.WL(WL216));
sram_cell_6t_5 inst_cell_216_23 (.BL(BL23),.BLN(BLN23),.WL(WL216));
sram_cell_6t_5 inst_cell_216_24 (.BL(BL24),.BLN(BLN24),.WL(WL216));
sram_cell_6t_5 inst_cell_216_25 (.BL(BL25),.BLN(BLN25),.WL(WL216));
sram_cell_6t_5 inst_cell_216_26 (.BL(BL26),.BLN(BLN26),.WL(WL216));
sram_cell_6t_5 inst_cell_216_27 (.BL(BL27),.BLN(BLN27),.WL(WL216));
sram_cell_6t_5 inst_cell_216_28 (.BL(BL28),.BLN(BLN28),.WL(WL216));
sram_cell_6t_5 inst_cell_216_29 (.BL(BL29),.BLN(BLN29),.WL(WL216));
sram_cell_6t_5 inst_cell_216_30 (.BL(BL30),.BLN(BLN30),.WL(WL216));
sram_cell_6t_5 inst_cell_216_31 (.BL(BL31),.BLN(BLN31),.WL(WL216));
sram_cell_6t_5 inst_cell_216_32 (.BL(BL32),.BLN(BLN32),.WL(WL216));
sram_cell_6t_5 inst_cell_216_33 (.BL(BL33),.BLN(BLN33),.WL(WL216));
sram_cell_6t_5 inst_cell_216_34 (.BL(BL34),.BLN(BLN34),.WL(WL216));
sram_cell_6t_5 inst_cell_216_35 (.BL(BL35),.BLN(BLN35),.WL(WL216));
sram_cell_6t_5 inst_cell_216_36 (.BL(BL36),.BLN(BLN36),.WL(WL216));
sram_cell_6t_5 inst_cell_216_37 (.BL(BL37),.BLN(BLN37),.WL(WL216));
sram_cell_6t_5 inst_cell_216_38 (.BL(BL38),.BLN(BLN38),.WL(WL216));
sram_cell_6t_5 inst_cell_216_39 (.BL(BL39),.BLN(BLN39),.WL(WL216));
sram_cell_6t_5 inst_cell_216_40 (.BL(BL40),.BLN(BLN40),.WL(WL216));
sram_cell_6t_5 inst_cell_216_41 (.BL(BL41),.BLN(BLN41),.WL(WL216));
sram_cell_6t_5 inst_cell_216_42 (.BL(BL42),.BLN(BLN42),.WL(WL216));
sram_cell_6t_5 inst_cell_216_43 (.BL(BL43),.BLN(BLN43),.WL(WL216));
sram_cell_6t_5 inst_cell_216_44 (.BL(BL44),.BLN(BLN44),.WL(WL216));
sram_cell_6t_5 inst_cell_216_45 (.BL(BL45),.BLN(BLN45),.WL(WL216));
sram_cell_6t_5 inst_cell_216_46 (.BL(BL46),.BLN(BLN46),.WL(WL216));
sram_cell_6t_5 inst_cell_216_47 (.BL(BL47),.BLN(BLN47),.WL(WL216));
sram_cell_6t_5 inst_cell_216_48 (.BL(BL48),.BLN(BLN48),.WL(WL216));
sram_cell_6t_5 inst_cell_216_49 (.BL(BL49),.BLN(BLN49),.WL(WL216));
sram_cell_6t_5 inst_cell_216_50 (.BL(BL50),.BLN(BLN50),.WL(WL216));
sram_cell_6t_5 inst_cell_216_51 (.BL(BL51),.BLN(BLN51),.WL(WL216));
sram_cell_6t_5 inst_cell_216_52 (.BL(BL52),.BLN(BLN52),.WL(WL216));
sram_cell_6t_5 inst_cell_216_53 (.BL(BL53),.BLN(BLN53),.WL(WL216));
sram_cell_6t_5 inst_cell_216_54 (.BL(BL54),.BLN(BLN54),.WL(WL216));
sram_cell_6t_5 inst_cell_216_55 (.BL(BL55),.BLN(BLN55),.WL(WL216));
sram_cell_6t_5 inst_cell_216_56 (.BL(BL56),.BLN(BLN56),.WL(WL216));
sram_cell_6t_5 inst_cell_216_57 (.BL(BL57),.BLN(BLN57),.WL(WL216));
sram_cell_6t_5 inst_cell_216_58 (.BL(BL58),.BLN(BLN58),.WL(WL216));
sram_cell_6t_5 inst_cell_216_59 (.BL(BL59),.BLN(BLN59),.WL(WL216));
sram_cell_6t_5 inst_cell_216_60 (.BL(BL60),.BLN(BLN60),.WL(WL216));
sram_cell_6t_5 inst_cell_216_61 (.BL(BL61),.BLN(BLN61),.WL(WL216));
sram_cell_6t_5 inst_cell_216_62 (.BL(BL62),.BLN(BLN62),.WL(WL216));
sram_cell_6t_5 inst_cell_216_63 (.BL(BL63),.BLN(BLN63),.WL(WL216));
sram_cell_6t_5 inst_cell_216_64 (.BL(BL64),.BLN(BLN64),.WL(WL216));
sram_cell_6t_5 inst_cell_216_65 (.BL(BL65),.BLN(BLN65),.WL(WL216));
sram_cell_6t_5 inst_cell_216_66 (.BL(BL66),.BLN(BLN66),.WL(WL216));
sram_cell_6t_5 inst_cell_216_67 (.BL(BL67),.BLN(BLN67),.WL(WL216));
sram_cell_6t_5 inst_cell_216_68 (.BL(BL68),.BLN(BLN68),.WL(WL216));
sram_cell_6t_5 inst_cell_216_69 (.BL(BL69),.BLN(BLN69),.WL(WL216));
sram_cell_6t_5 inst_cell_216_70 (.BL(BL70),.BLN(BLN70),.WL(WL216));
sram_cell_6t_5 inst_cell_216_71 (.BL(BL71),.BLN(BLN71),.WL(WL216));
sram_cell_6t_5 inst_cell_216_72 (.BL(BL72),.BLN(BLN72),.WL(WL216));
sram_cell_6t_5 inst_cell_216_73 (.BL(BL73),.BLN(BLN73),.WL(WL216));
sram_cell_6t_5 inst_cell_216_74 (.BL(BL74),.BLN(BLN74),.WL(WL216));
sram_cell_6t_5 inst_cell_216_75 (.BL(BL75),.BLN(BLN75),.WL(WL216));
sram_cell_6t_5 inst_cell_216_76 (.BL(BL76),.BLN(BLN76),.WL(WL216));
sram_cell_6t_5 inst_cell_216_77 (.BL(BL77),.BLN(BLN77),.WL(WL216));
sram_cell_6t_5 inst_cell_216_78 (.BL(BL78),.BLN(BLN78),.WL(WL216));
sram_cell_6t_5 inst_cell_216_79 (.BL(BL79),.BLN(BLN79),.WL(WL216));
sram_cell_6t_5 inst_cell_216_80 (.BL(BL80),.BLN(BLN80),.WL(WL216));
sram_cell_6t_5 inst_cell_216_81 (.BL(BL81),.BLN(BLN81),.WL(WL216));
sram_cell_6t_5 inst_cell_216_82 (.BL(BL82),.BLN(BLN82),.WL(WL216));
sram_cell_6t_5 inst_cell_216_83 (.BL(BL83),.BLN(BLN83),.WL(WL216));
sram_cell_6t_5 inst_cell_216_84 (.BL(BL84),.BLN(BLN84),.WL(WL216));
sram_cell_6t_5 inst_cell_216_85 (.BL(BL85),.BLN(BLN85),.WL(WL216));
sram_cell_6t_5 inst_cell_216_86 (.BL(BL86),.BLN(BLN86),.WL(WL216));
sram_cell_6t_5 inst_cell_216_87 (.BL(BL87),.BLN(BLN87),.WL(WL216));
sram_cell_6t_5 inst_cell_216_88 (.BL(BL88),.BLN(BLN88),.WL(WL216));
sram_cell_6t_5 inst_cell_216_89 (.BL(BL89),.BLN(BLN89),.WL(WL216));
sram_cell_6t_5 inst_cell_216_90 (.BL(BL90),.BLN(BLN90),.WL(WL216));
sram_cell_6t_5 inst_cell_216_91 (.BL(BL91),.BLN(BLN91),.WL(WL216));
sram_cell_6t_5 inst_cell_216_92 (.BL(BL92),.BLN(BLN92),.WL(WL216));
sram_cell_6t_5 inst_cell_216_93 (.BL(BL93),.BLN(BLN93),.WL(WL216));
sram_cell_6t_5 inst_cell_216_94 (.BL(BL94),.BLN(BLN94),.WL(WL216));
sram_cell_6t_5 inst_cell_216_95 (.BL(BL95),.BLN(BLN95),.WL(WL216));
sram_cell_6t_5 inst_cell_216_96 (.BL(BL96),.BLN(BLN96),.WL(WL216));
sram_cell_6t_5 inst_cell_216_97 (.BL(BL97),.BLN(BLN97),.WL(WL216));
sram_cell_6t_5 inst_cell_216_98 (.BL(BL98),.BLN(BLN98),.WL(WL216));
sram_cell_6t_5 inst_cell_216_99 (.BL(BL99),.BLN(BLN99),.WL(WL216));
sram_cell_6t_5 inst_cell_216_100 (.BL(BL100),.BLN(BLN100),.WL(WL216));
sram_cell_6t_5 inst_cell_216_101 (.BL(BL101),.BLN(BLN101),.WL(WL216));
sram_cell_6t_5 inst_cell_216_102 (.BL(BL102),.BLN(BLN102),.WL(WL216));
sram_cell_6t_5 inst_cell_216_103 (.BL(BL103),.BLN(BLN103),.WL(WL216));
sram_cell_6t_5 inst_cell_216_104 (.BL(BL104),.BLN(BLN104),.WL(WL216));
sram_cell_6t_5 inst_cell_216_105 (.BL(BL105),.BLN(BLN105),.WL(WL216));
sram_cell_6t_5 inst_cell_216_106 (.BL(BL106),.BLN(BLN106),.WL(WL216));
sram_cell_6t_5 inst_cell_216_107 (.BL(BL107),.BLN(BLN107),.WL(WL216));
sram_cell_6t_5 inst_cell_216_108 (.BL(BL108),.BLN(BLN108),.WL(WL216));
sram_cell_6t_5 inst_cell_216_109 (.BL(BL109),.BLN(BLN109),.WL(WL216));
sram_cell_6t_5 inst_cell_216_110 (.BL(BL110),.BLN(BLN110),.WL(WL216));
sram_cell_6t_5 inst_cell_216_111 (.BL(BL111),.BLN(BLN111),.WL(WL216));
sram_cell_6t_5 inst_cell_216_112 (.BL(BL112),.BLN(BLN112),.WL(WL216));
sram_cell_6t_5 inst_cell_216_113 (.BL(BL113),.BLN(BLN113),.WL(WL216));
sram_cell_6t_5 inst_cell_216_114 (.BL(BL114),.BLN(BLN114),.WL(WL216));
sram_cell_6t_5 inst_cell_216_115 (.BL(BL115),.BLN(BLN115),.WL(WL216));
sram_cell_6t_5 inst_cell_216_116 (.BL(BL116),.BLN(BLN116),.WL(WL216));
sram_cell_6t_5 inst_cell_216_117 (.BL(BL117),.BLN(BLN117),.WL(WL216));
sram_cell_6t_5 inst_cell_216_118 (.BL(BL118),.BLN(BLN118),.WL(WL216));
sram_cell_6t_5 inst_cell_216_119 (.BL(BL119),.BLN(BLN119),.WL(WL216));
sram_cell_6t_5 inst_cell_216_120 (.BL(BL120),.BLN(BLN120),.WL(WL216));
sram_cell_6t_5 inst_cell_216_121 (.BL(BL121),.BLN(BLN121),.WL(WL216));
sram_cell_6t_5 inst_cell_216_122 (.BL(BL122),.BLN(BLN122),.WL(WL216));
sram_cell_6t_5 inst_cell_216_123 (.BL(BL123),.BLN(BLN123),.WL(WL216));
sram_cell_6t_5 inst_cell_216_124 (.BL(BL124),.BLN(BLN124),.WL(WL216));
sram_cell_6t_5 inst_cell_216_125 (.BL(BL125),.BLN(BLN125),.WL(WL216));
sram_cell_6t_5 inst_cell_216_126 (.BL(BL126),.BLN(BLN126),.WL(WL216));
sram_cell_6t_5 inst_cell_216_127 (.BL(BL127),.BLN(BLN127),.WL(WL216));
sram_cell_6t_5 inst_cell_217_0 (.BL(BL0),.BLN(BLN0),.WL(WL217));
sram_cell_6t_5 inst_cell_217_1 (.BL(BL1),.BLN(BLN1),.WL(WL217));
sram_cell_6t_5 inst_cell_217_2 (.BL(BL2),.BLN(BLN2),.WL(WL217));
sram_cell_6t_5 inst_cell_217_3 (.BL(BL3),.BLN(BLN3),.WL(WL217));
sram_cell_6t_5 inst_cell_217_4 (.BL(BL4),.BLN(BLN4),.WL(WL217));
sram_cell_6t_5 inst_cell_217_5 (.BL(BL5),.BLN(BLN5),.WL(WL217));
sram_cell_6t_5 inst_cell_217_6 (.BL(BL6),.BLN(BLN6),.WL(WL217));
sram_cell_6t_5 inst_cell_217_7 (.BL(BL7),.BLN(BLN7),.WL(WL217));
sram_cell_6t_5 inst_cell_217_8 (.BL(BL8),.BLN(BLN8),.WL(WL217));
sram_cell_6t_5 inst_cell_217_9 (.BL(BL9),.BLN(BLN9),.WL(WL217));
sram_cell_6t_5 inst_cell_217_10 (.BL(BL10),.BLN(BLN10),.WL(WL217));
sram_cell_6t_5 inst_cell_217_11 (.BL(BL11),.BLN(BLN11),.WL(WL217));
sram_cell_6t_5 inst_cell_217_12 (.BL(BL12),.BLN(BLN12),.WL(WL217));
sram_cell_6t_5 inst_cell_217_13 (.BL(BL13),.BLN(BLN13),.WL(WL217));
sram_cell_6t_5 inst_cell_217_14 (.BL(BL14),.BLN(BLN14),.WL(WL217));
sram_cell_6t_5 inst_cell_217_15 (.BL(BL15),.BLN(BLN15),.WL(WL217));
sram_cell_6t_5 inst_cell_217_16 (.BL(BL16),.BLN(BLN16),.WL(WL217));
sram_cell_6t_5 inst_cell_217_17 (.BL(BL17),.BLN(BLN17),.WL(WL217));
sram_cell_6t_5 inst_cell_217_18 (.BL(BL18),.BLN(BLN18),.WL(WL217));
sram_cell_6t_5 inst_cell_217_19 (.BL(BL19),.BLN(BLN19),.WL(WL217));
sram_cell_6t_5 inst_cell_217_20 (.BL(BL20),.BLN(BLN20),.WL(WL217));
sram_cell_6t_5 inst_cell_217_21 (.BL(BL21),.BLN(BLN21),.WL(WL217));
sram_cell_6t_5 inst_cell_217_22 (.BL(BL22),.BLN(BLN22),.WL(WL217));
sram_cell_6t_5 inst_cell_217_23 (.BL(BL23),.BLN(BLN23),.WL(WL217));
sram_cell_6t_5 inst_cell_217_24 (.BL(BL24),.BLN(BLN24),.WL(WL217));
sram_cell_6t_5 inst_cell_217_25 (.BL(BL25),.BLN(BLN25),.WL(WL217));
sram_cell_6t_5 inst_cell_217_26 (.BL(BL26),.BLN(BLN26),.WL(WL217));
sram_cell_6t_5 inst_cell_217_27 (.BL(BL27),.BLN(BLN27),.WL(WL217));
sram_cell_6t_5 inst_cell_217_28 (.BL(BL28),.BLN(BLN28),.WL(WL217));
sram_cell_6t_5 inst_cell_217_29 (.BL(BL29),.BLN(BLN29),.WL(WL217));
sram_cell_6t_5 inst_cell_217_30 (.BL(BL30),.BLN(BLN30),.WL(WL217));
sram_cell_6t_5 inst_cell_217_31 (.BL(BL31),.BLN(BLN31),.WL(WL217));
sram_cell_6t_5 inst_cell_217_32 (.BL(BL32),.BLN(BLN32),.WL(WL217));
sram_cell_6t_5 inst_cell_217_33 (.BL(BL33),.BLN(BLN33),.WL(WL217));
sram_cell_6t_5 inst_cell_217_34 (.BL(BL34),.BLN(BLN34),.WL(WL217));
sram_cell_6t_5 inst_cell_217_35 (.BL(BL35),.BLN(BLN35),.WL(WL217));
sram_cell_6t_5 inst_cell_217_36 (.BL(BL36),.BLN(BLN36),.WL(WL217));
sram_cell_6t_5 inst_cell_217_37 (.BL(BL37),.BLN(BLN37),.WL(WL217));
sram_cell_6t_5 inst_cell_217_38 (.BL(BL38),.BLN(BLN38),.WL(WL217));
sram_cell_6t_5 inst_cell_217_39 (.BL(BL39),.BLN(BLN39),.WL(WL217));
sram_cell_6t_5 inst_cell_217_40 (.BL(BL40),.BLN(BLN40),.WL(WL217));
sram_cell_6t_5 inst_cell_217_41 (.BL(BL41),.BLN(BLN41),.WL(WL217));
sram_cell_6t_5 inst_cell_217_42 (.BL(BL42),.BLN(BLN42),.WL(WL217));
sram_cell_6t_5 inst_cell_217_43 (.BL(BL43),.BLN(BLN43),.WL(WL217));
sram_cell_6t_5 inst_cell_217_44 (.BL(BL44),.BLN(BLN44),.WL(WL217));
sram_cell_6t_5 inst_cell_217_45 (.BL(BL45),.BLN(BLN45),.WL(WL217));
sram_cell_6t_5 inst_cell_217_46 (.BL(BL46),.BLN(BLN46),.WL(WL217));
sram_cell_6t_5 inst_cell_217_47 (.BL(BL47),.BLN(BLN47),.WL(WL217));
sram_cell_6t_5 inst_cell_217_48 (.BL(BL48),.BLN(BLN48),.WL(WL217));
sram_cell_6t_5 inst_cell_217_49 (.BL(BL49),.BLN(BLN49),.WL(WL217));
sram_cell_6t_5 inst_cell_217_50 (.BL(BL50),.BLN(BLN50),.WL(WL217));
sram_cell_6t_5 inst_cell_217_51 (.BL(BL51),.BLN(BLN51),.WL(WL217));
sram_cell_6t_5 inst_cell_217_52 (.BL(BL52),.BLN(BLN52),.WL(WL217));
sram_cell_6t_5 inst_cell_217_53 (.BL(BL53),.BLN(BLN53),.WL(WL217));
sram_cell_6t_5 inst_cell_217_54 (.BL(BL54),.BLN(BLN54),.WL(WL217));
sram_cell_6t_5 inst_cell_217_55 (.BL(BL55),.BLN(BLN55),.WL(WL217));
sram_cell_6t_5 inst_cell_217_56 (.BL(BL56),.BLN(BLN56),.WL(WL217));
sram_cell_6t_5 inst_cell_217_57 (.BL(BL57),.BLN(BLN57),.WL(WL217));
sram_cell_6t_5 inst_cell_217_58 (.BL(BL58),.BLN(BLN58),.WL(WL217));
sram_cell_6t_5 inst_cell_217_59 (.BL(BL59),.BLN(BLN59),.WL(WL217));
sram_cell_6t_5 inst_cell_217_60 (.BL(BL60),.BLN(BLN60),.WL(WL217));
sram_cell_6t_5 inst_cell_217_61 (.BL(BL61),.BLN(BLN61),.WL(WL217));
sram_cell_6t_5 inst_cell_217_62 (.BL(BL62),.BLN(BLN62),.WL(WL217));
sram_cell_6t_5 inst_cell_217_63 (.BL(BL63),.BLN(BLN63),.WL(WL217));
sram_cell_6t_5 inst_cell_217_64 (.BL(BL64),.BLN(BLN64),.WL(WL217));
sram_cell_6t_5 inst_cell_217_65 (.BL(BL65),.BLN(BLN65),.WL(WL217));
sram_cell_6t_5 inst_cell_217_66 (.BL(BL66),.BLN(BLN66),.WL(WL217));
sram_cell_6t_5 inst_cell_217_67 (.BL(BL67),.BLN(BLN67),.WL(WL217));
sram_cell_6t_5 inst_cell_217_68 (.BL(BL68),.BLN(BLN68),.WL(WL217));
sram_cell_6t_5 inst_cell_217_69 (.BL(BL69),.BLN(BLN69),.WL(WL217));
sram_cell_6t_5 inst_cell_217_70 (.BL(BL70),.BLN(BLN70),.WL(WL217));
sram_cell_6t_5 inst_cell_217_71 (.BL(BL71),.BLN(BLN71),.WL(WL217));
sram_cell_6t_5 inst_cell_217_72 (.BL(BL72),.BLN(BLN72),.WL(WL217));
sram_cell_6t_5 inst_cell_217_73 (.BL(BL73),.BLN(BLN73),.WL(WL217));
sram_cell_6t_5 inst_cell_217_74 (.BL(BL74),.BLN(BLN74),.WL(WL217));
sram_cell_6t_5 inst_cell_217_75 (.BL(BL75),.BLN(BLN75),.WL(WL217));
sram_cell_6t_5 inst_cell_217_76 (.BL(BL76),.BLN(BLN76),.WL(WL217));
sram_cell_6t_5 inst_cell_217_77 (.BL(BL77),.BLN(BLN77),.WL(WL217));
sram_cell_6t_5 inst_cell_217_78 (.BL(BL78),.BLN(BLN78),.WL(WL217));
sram_cell_6t_5 inst_cell_217_79 (.BL(BL79),.BLN(BLN79),.WL(WL217));
sram_cell_6t_5 inst_cell_217_80 (.BL(BL80),.BLN(BLN80),.WL(WL217));
sram_cell_6t_5 inst_cell_217_81 (.BL(BL81),.BLN(BLN81),.WL(WL217));
sram_cell_6t_5 inst_cell_217_82 (.BL(BL82),.BLN(BLN82),.WL(WL217));
sram_cell_6t_5 inst_cell_217_83 (.BL(BL83),.BLN(BLN83),.WL(WL217));
sram_cell_6t_5 inst_cell_217_84 (.BL(BL84),.BLN(BLN84),.WL(WL217));
sram_cell_6t_5 inst_cell_217_85 (.BL(BL85),.BLN(BLN85),.WL(WL217));
sram_cell_6t_5 inst_cell_217_86 (.BL(BL86),.BLN(BLN86),.WL(WL217));
sram_cell_6t_5 inst_cell_217_87 (.BL(BL87),.BLN(BLN87),.WL(WL217));
sram_cell_6t_5 inst_cell_217_88 (.BL(BL88),.BLN(BLN88),.WL(WL217));
sram_cell_6t_5 inst_cell_217_89 (.BL(BL89),.BLN(BLN89),.WL(WL217));
sram_cell_6t_5 inst_cell_217_90 (.BL(BL90),.BLN(BLN90),.WL(WL217));
sram_cell_6t_5 inst_cell_217_91 (.BL(BL91),.BLN(BLN91),.WL(WL217));
sram_cell_6t_5 inst_cell_217_92 (.BL(BL92),.BLN(BLN92),.WL(WL217));
sram_cell_6t_5 inst_cell_217_93 (.BL(BL93),.BLN(BLN93),.WL(WL217));
sram_cell_6t_5 inst_cell_217_94 (.BL(BL94),.BLN(BLN94),.WL(WL217));
sram_cell_6t_5 inst_cell_217_95 (.BL(BL95),.BLN(BLN95),.WL(WL217));
sram_cell_6t_5 inst_cell_217_96 (.BL(BL96),.BLN(BLN96),.WL(WL217));
sram_cell_6t_5 inst_cell_217_97 (.BL(BL97),.BLN(BLN97),.WL(WL217));
sram_cell_6t_5 inst_cell_217_98 (.BL(BL98),.BLN(BLN98),.WL(WL217));
sram_cell_6t_5 inst_cell_217_99 (.BL(BL99),.BLN(BLN99),.WL(WL217));
sram_cell_6t_5 inst_cell_217_100 (.BL(BL100),.BLN(BLN100),.WL(WL217));
sram_cell_6t_5 inst_cell_217_101 (.BL(BL101),.BLN(BLN101),.WL(WL217));
sram_cell_6t_5 inst_cell_217_102 (.BL(BL102),.BLN(BLN102),.WL(WL217));
sram_cell_6t_5 inst_cell_217_103 (.BL(BL103),.BLN(BLN103),.WL(WL217));
sram_cell_6t_5 inst_cell_217_104 (.BL(BL104),.BLN(BLN104),.WL(WL217));
sram_cell_6t_5 inst_cell_217_105 (.BL(BL105),.BLN(BLN105),.WL(WL217));
sram_cell_6t_5 inst_cell_217_106 (.BL(BL106),.BLN(BLN106),.WL(WL217));
sram_cell_6t_5 inst_cell_217_107 (.BL(BL107),.BLN(BLN107),.WL(WL217));
sram_cell_6t_5 inst_cell_217_108 (.BL(BL108),.BLN(BLN108),.WL(WL217));
sram_cell_6t_5 inst_cell_217_109 (.BL(BL109),.BLN(BLN109),.WL(WL217));
sram_cell_6t_5 inst_cell_217_110 (.BL(BL110),.BLN(BLN110),.WL(WL217));
sram_cell_6t_5 inst_cell_217_111 (.BL(BL111),.BLN(BLN111),.WL(WL217));
sram_cell_6t_5 inst_cell_217_112 (.BL(BL112),.BLN(BLN112),.WL(WL217));
sram_cell_6t_5 inst_cell_217_113 (.BL(BL113),.BLN(BLN113),.WL(WL217));
sram_cell_6t_5 inst_cell_217_114 (.BL(BL114),.BLN(BLN114),.WL(WL217));
sram_cell_6t_5 inst_cell_217_115 (.BL(BL115),.BLN(BLN115),.WL(WL217));
sram_cell_6t_5 inst_cell_217_116 (.BL(BL116),.BLN(BLN116),.WL(WL217));
sram_cell_6t_5 inst_cell_217_117 (.BL(BL117),.BLN(BLN117),.WL(WL217));
sram_cell_6t_5 inst_cell_217_118 (.BL(BL118),.BLN(BLN118),.WL(WL217));
sram_cell_6t_5 inst_cell_217_119 (.BL(BL119),.BLN(BLN119),.WL(WL217));
sram_cell_6t_5 inst_cell_217_120 (.BL(BL120),.BLN(BLN120),.WL(WL217));
sram_cell_6t_5 inst_cell_217_121 (.BL(BL121),.BLN(BLN121),.WL(WL217));
sram_cell_6t_5 inst_cell_217_122 (.BL(BL122),.BLN(BLN122),.WL(WL217));
sram_cell_6t_5 inst_cell_217_123 (.BL(BL123),.BLN(BLN123),.WL(WL217));
sram_cell_6t_5 inst_cell_217_124 (.BL(BL124),.BLN(BLN124),.WL(WL217));
sram_cell_6t_5 inst_cell_217_125 (.BL(BL125),.BLN(BLN125),.WL(WL217));
sram_cell_6t_5 inst_cell_217_126 (.BL(BL126),.BLN(BLN126),.WL(WL217));
sram_cell_6t_5 inst_cell_217_127 (.BL(BL127),.BLN(BLN127),.WL(WL217));
sram_cell_6t_5 inst_cell_218_0 (.BL(BL0),.BLN(BLN0),.WL(WL218));
sram_cell_6t_5 inst_cell_218_1 (.BL(BL1),.BLN(BLN1),.WL(WL218));
sram_cell_6t_5 inst_cell_218_2 (.BL(BL2),.BLN(BLN2),.WL(WL218));
sram_cell_6t_5 inst_cell_218_3 (.BL(BL3),.BLN(BLN3),.WL(WL218));
sram_cell_6t_5 inst_cell_218_4 (.BL(BL4),.BLN(BLN4),.WL(WL218));
sram_cell_6t_5 inst_cell_218_5 (.BL(BL5),.BLN(BLN5),.WL(WL218));
sram_cell_6t_5 inst_cell_218_6 (.BL(BL6),.BLN(BLN6),.WL(WL218));
sram_cell_6t_5 inst_cell_218_7 (.BL(BL7),.BLN(BLN7),.WL(WL218));
sram_cell_6t_5 inst_cell_218_8 (.BL(BL8),.BLN(BLN8),.WL(WL218));
sram_cell_6t_5 inst_cell_218_9 (.BL(BL9),.BLN(BLN9),.WL(WL218));
sram_cell_6t_5 inst_cell_218_10 (.BL(BL10),.BLN(BLN10),.WL(WL218));
sram_cell_6t_5 inst_cell_218_11 (.BL(BL11),.BLN(BLN11),.WL(WL218));
sram_cell_6t_5 inst_cell_218_12 (.BL(BL12),.BLN(BLN12),.WL(WL218));
sram_cell_6t_5 inst_cell_218_13 (.BL(BL13),.BLN(BLN13),.WL(WL218));
sram_cell_6t_5 inst_cell_218_14 (.BL(BL14),.BLN(BLN14),.WL(WL218));
sram_cell_6t_5 inst_cell_218_15 (.BL(BL15),.BLN(BLN15),.WL(WL218));
sram_cell_6t_5 inst_cell_218_16 (.BL(BL16),.BLN(BLN16),.WL(WL218));
sram_cell_6t_5 inst_cell_218_17 (.BL(BL17),.BLN(BLN17),.WL(WL218));
sram_cell_6t_5 inst_cell_218_18 (.BL(BL18),.BLN(BLN18),.WL(WL218));
sram_cell_6t_5 inst_cell_218_19 (.BL(BL19),.BLN(BLN19),.WL(WL218));
sram_cell_6t_5 inst_cell_218_20 (.BL(BL20),.BLN(BLN20),.WL(WL218));
sram_cell_6t_5 inst_cell_218_21 (.BL(BL21),.BLN(BLN21),.WL(WL218));
sram_cell_6t_5 inst_cell_218_22 (.BL(BL22),.BLN(BLN22),.WL(WL218));
sram_cell_6t_5 inst_cell_218_23 (.BL(BL23),.BLN(BLN23),.WL(WL218));
sram_cell_6t_5 inst_cell_218_24 (.BL(BL24),.BLN(BLN24),.WL(WL218));
sram_cell_6t_5 inst_cell_218_25 (.BL(BL25),.BLN(BLN25),.WL(WL218));
sram_cell_6t_5 inst_cell_218_26 (.BL(BL26),.BLN(BLN26),.WL(WL218));
sram_cell_6t_5 inst_cell_218_27 (.BL(BL27),.BLN(BLN27),.WL(WL218));
sram_cell_6t_5 inst_cell_218_28 (.BL(BL28),.BLN(BLN28),.WL(WL218));
sram_cell_6t_5 inst_cell_218_29 (.BL(BL29),.BLN(BLN29),.WL(WL218));
sram_cell_6t_5 inst_cell_218_30 (.BL(BL30),.BLN(BLN30),.WL(WL218));
sram_cell_6t_5 inst_cell_218_31 (.BL(BL31),.BLN(BLN31),.WL(WL218));
sram_cell_6t_5 inst_cell_218_32 (.BL(BL32),.BLN(BLN32),.WL(WL218));
sram_cell_6t_5 inst_cell_218_33 (.BL(BL33),.BLN(BLN33),.WL(WL218));
sram_cell_6t_5 inst_cell_218_34 (.BL(BL34),.BLN(BLN34),.WL(WL218));
sram_cell_6t_5 inst_cell_218_35 (.BL(BL35),.BLN(BLN35),.WL(WL218));
sram_cell_6t_5 inst_cell_218_36 (.BL(BL36),.BLN(BLN36),.WL(WL218));
sram_cell_6t_5 inst_cell_218_37 (.BL(BL37),.BLN(BLN37),.WL(WL218));
sram_cell_6t_5 inst_cell_218_38 (.BL(BL38),.BLN(BLN38),.WL(WL218));
sram_cell_6t_5 inst_cell_218_39 (.BL(BL39),.BLN(BLN39),.WL(WL218));
sram_cell_6t_5 inst_cell_218_40 (.BL(BL40),.BLN(BLN40),.WL(WL218));
sram_cell_6t_5 inst_cell_218_41 (.BL(BL41),.BLN(BLN41),.WL(WL218));
sram_cell_6t_5 inst_cell_218_42 (.BL(BL42),.BLN(BLN42),.WL(WL218));
sram_cell_6t_5 inst_cell_218_43 (.BL(BL43),.BLN(BLN43),.WL(WL218));
sram_cell_6t_5 inst_cell_218_44 (.BL(BL44),.BLN(BLN44),.WL(WL218));
sram_cell_6t_5 inst_cell_218_45 (.BL(BL45),.BLN(BLN45),.WL(WL218));
sram_cell_6t_5 inst_cell_218_46 (.BL(BL46),.BLN(BLN46),.WL(WL218));
sram_cell_6t_5 inst_cell_218_47 (.BL(BL47),.BLN(BLN47),.WL(WL218));
sram_cell_6t_5 inst_cell_218_48 (.BL(BL48),.BLN(BLN48),.WL(WL218));
sram_cell_6t_5 inst_cell_218_49 (.BL(BL49),.BLN(BLN49),.WL(WL218));
sram_cell_6t_5 inst_cell_218_50 (.BL(BL50),.BLN(BLN50),.WL(WL218));
sram_cell_6t_5 inst_cell_218_51 (.BL(BL51),.BLN(BLN51),.WL(WL218));
sram_cell_6t_5 inst_cell_218_52 (.BL(BL52),.BLN(BLN52),.WL(WL218));
sram_cell_6t_5 inst_cell_218_53 (.BL(BL53),.BLN(BLN53),.WL(WL218));
sram_cell_6t_5 inst_cell_218_54 (.BL(BL54),.BLN(BLN54),.WL(WL218));
sram_cell_6t_5 inst_cell_218_55 (.BL(BL55),.BLN(BLN55),.WL(WL218));
sram_cell_6t_5 inst_cell_218_56 (.BL(BL56),.BLN(BLN56),.WL(WL218));
sram_cell_6t_5 inst_cell_218_57 (.BL(BL57),.BLN(BLN57),.WL(WL218));
sram_cell_6t_5 inst_cell_218_58 (.BL(BL58),.BLN(BLN58),.WL(WL218));
sram_cell_6t_5 inst_cell_218_59 (.BL(BL59),.BLN(BLN59),.WL(WL218));
sram_cell_6t_5 inst_cell_218_60 (.BL(BL60),.BLN(BLN60),.WL(WL218));
sram_cell_6t_5 inst_cell_218_61 (.BL(BL61),.BLN(BLN61),.WL(WL218));
sram_cell_6t_5 inst_cell_218_62 (.BL(BL62),.BLN(BLN62),.WL(WL218));
sram_cell_6t_5 inst_cell_218_63 (.BL(BL63),.BLN(BLN63),.WL(WL218));
sram_cell_6t_5 inst_cell_218_64 (.BL(BL64),.BLN(BLN64),.WL(WL218));
sram_cell_6t_5 inst_cell_218_65 (.BL(BL65),.BLN(BLN65),.WL(WL218));
sram_cell_6t_5 inst_cell_218_66 (.BL(BL66),.BLN(BLN66),.WL(WL218));
sram_cell_6t_5 inst_cell_218_67 (.BL(BL67),.BLN(BLN67),.WL(WL218));
sram_cell_6t_5 inst_cell_218_68 (.BL(BL68),.BLN(BLN68),.WL(WL218));
sram_cell_6t_5 inst_cell_218_69 (.BL(BL69),.BLN(BLN69),.WL(WL218));
sram_cell_6t_5 inst_cell_218_70 (.BL(BL70),.BLN(BLN70),.WL(WL218));
sram_cell_6t_5 inst_cell_218_71 (.BL(BL71),.BLN(BLN71),.WL(WL218));
sram_cell_6t_5 inst_cell_218_72 (.BL(BL72),.BLN(BLN72),.WL(WL218));
sram_cell_6t_5 inst_cell_218_73 (.BL(BL73),.BLN(BLN73),.WL(WL218));
sram_cell_6t_5 inst_cell_218_74 (.BL(BL74),.BLN(BLN74),.WL(WL218));
sram_cell_6t_5 inst_cell_218_75 (.BL(BL75),.BLN(BLN75),.WL(WL218));
sram_cell_6t_5 inst_cell_218_76 (.BL(BL76),.BLN(BLN76),.WL(WL218));
sram_cell_6t_5 inst_cell_218_77 (.BL(BL77),.BLN(BLN77),.WL(WL218));
sram_cell_6t_5 inst_cell_218_78 (.BL(BL78),.BLN(BLN78),.WL(WL218));
sram_cell_6t_5 inst_cell_218_79 (.BL(BL79),.BLN(BLN79),.WL(WL218));
sram_cell_6t_5 inst_cell_218_80 (.BL(BL80),.BLN(BLN80),.WL(WL218));
sram_cell_6t_5 inst_cell_218_81 (.BL(BL81),.BLN(BLN81),.WL(WL218));
sram_cell_6t_5 inst_cell_218_82 (.BL(BL82),.BLN(BLN82),.WL(WL218));
sram_cell_6t_5 inst_cell_218_83 (.BL(BL83),.BLN(BLN83),.WL(WL218));
sram_cell_6t_5 inst_cell_218_84 (.BL(BL84),.BLN(BLN84),.WL(WL218));
sram_cell_6t_5 inst_cell_218_85 (.BL(BL85),.BLN(BLN85),.WL(WL218));
sram_cell_6t_5 inst_cell_218_86 (.BL(BL86),.BLN(BLN86),.WL(WL218));
sram_cell_6t_5 inst_cell_218_87 (.BL(BL87),.BLN(BLN87),.WL(WL218));
sram_cell_6t_5 inst_cell_218_88 (.BL(BL88),.BLN(BLN88),.WL(WL218));
sram_cell_6t_5 inst_cell_218_89 (.BL(BL89),.BLN(BLN89),.WL(WL218));
sram_cell_6t_5 inst_cell_218_90 (.BL(BL90),.BLN(BLN90),.WL(WL218));
sram_cell_6t_5 inst_cell_218_91 (.BL(BL91),.BLN(BLN91),.WL(WL218));
sram_cell_6t_5 inst_cell_218_92 (.BL(BL92),.BLN(BLN92),.WL(WL218));
sram_cell_6t_5 inst_cell_218_93 (.BL(BL93),.BLN(BLN93),.WL(WL218));
sram_cell_6t_5 inst_cell_218_94 (.BL(BL94),.BLN(BLN94),.WL(WL218));
sram_cell_6t_5 inst_cell_218_95 (.BL(BL95),.BLN(BLN95),.WL(WL218));
sram_cell_6t_5 inst_cell_218_96 (.BL(BL96),.BLN(BLN96),.WL(WL218));
sram_cell_6t_5 inst_cell_218_97 (.BL(BL97),.BLN(BLN97),.WL(WL218));
sram_cell_6t_5 inst_cell_218_98 (.BL(BL98),.BLN(BLN98),.WL(WL218));
sram_cell_6t_5 inst_cell_218_99 (.BL(BL99),.BLN(BLN99),.WL(WL218));
sram_cell_6t_5 inst_cell_218_100 (.BL(BL100),.BLN(BLN100),.WL(WL218));
sram_cell_6t_5 inst_cell_218_101 (.BL(BL101),.BLN(BLN101),.WL(WL218));
sram_cell_6t_5 inst_cell_218_102 (.BL(BL102),.BLN(BLN102),.WL(WL218));
sram_cell_6t_5 inst_cell_218_103 (.BL(BL103),.BLN(BLN103),.WL(WL218));
sram_cell_6t_5 inst_cell_218_104 (.BL(BL104),.BLN(BLN104),.WL(WL218));
sram_cell_6t_5 inst_cell_218_105 (.BL(BL105),.BLN(BLN105),.WL(WL218));
sram_cell_6t_5 inst_cell_218_106 (.BL(BL106),.BLN(BLN106),.WL(WL218));
sram_cell_6t_5 inst_cell_218_107 (.BL(BL107),.BLN(BLN107),.WL(WL218));
sram_cell_6t_5 inst_cell_218_108 (.BL(BL108),.BLN(BLN108),.WL(WL218));
sram_cell_6t_5 inst_cell_218_109 (.BL(BL109),.BLN(BLN109),.WL(WL218));
sram_cell_6t_5 inst_cell_218_110 (.BL(BL110),.BLN(BLN110),.WL(WL218));
sram_cell_6t_5 inst_cell_218_111 (.BL(BL111),.BLN(BLN111),.WL(WL218));
sram_cell_6t_5 inst_cell_218_112 (.BL(BL112),.BLN(BLN112),.WL(WL218));
sram_cell_6t_5 inst_cell_218_113 (.BL(BL113),.BLN(BLN113),.WL(WL218));
sram_cell_6t_5 inst_cell_218_114 (.BL(BL114),.BLN(BLN114),.WL(WL218));
sram_cell_6t_5 inst_cell_218_115 (.BL(BL115),.BLN(BLN115),.WL(WL218));
sram_cell_6t_5 inst_cell_218_116 (.BL(BL116),.BLN(BLN116),.WL(WL218));
sram_cell_6t_5 inst_cell_218_117 (.BL(BL117),.BLN(BLN117),.WL(WL218));
sram_cell_6t_5 inst_cell_218_118 (.BL(BL118),.BLN(BLN118),.WL(WL218));
sram_cell_6t_5 inst_cell_218_119 (.BL(BL119),.BLN(BLN119),.WL(WL218));
sram_cell_6t_5 inst_cell_218_120 (.BL(BL120),.BLN(BLN120),.WL(WL218));
sram_cell_6t_5 inst_cell_218_121 (.BL(BL121),.BLN(BLN121),.WL(WL218));
sram_cell_6t_5 inst_cell_218_122 (.BL(BL122),.BLN(BLN122),.WL(WL218));
sram_cell_6t_5 inst_cell_218_123 (.BL(BL123),.BLN(BLN123),.WL(WL218));
sram_cell_6t_5 inst_cell_218_124 (.BL(BL124),.BLN(BLN124),.WL(WL218));
sram_cell_6t_5 inst_cell_218_125 (.BL(BL125),.BLN(BLN125),.WL(WL218));
sram_cell_6t_5 inst_cell_218_126 (.BL(BL126),.BLN(BLN126),.WL(WL218));
sram_cell_6t_5 inst_cell_218_127 (.BL(BL127),.BLN(BLN127),.WL(WL218));
sram_cell_6t_5 inst_cell_219_0 (.BL(BL0),.BLN(BLN0),.WL(WL219));
sram_cell_6t_5 inst_cell_219_1 (.BL(BL1),.BLN(BLN1),.WL(WL219));
sram_cell_6t_5 inst_cell_219_2 (.BL(BL2),.BLN(BLN2),.WL(WL219));
sram_cell_6t_5 inst_cell_219_3 (.BL(BL3),.BLN(BLN3),.WL(WL219));
sram_cell_6t_5 inst_cell_219_4 (.BL(BL4),.BLN(BLN4),.WL(WL219));
sram_cell_6t_5 inst_cell_219_5 (.BL(BL5),.BLN(BLN5),.WL(WL219));
sram_cell_6t_5 inst_cell_219_6 (.BL(BL6),.BLN(BLN6),.WL(WL219));
sram_cell_6t_5 inst_cell_219_7 (.BL(BL7),.BLN(BLN7),.WL(WL219));
sram_cell_6t_5 inst_cell_219_8 (.BL(BL8),.BLN(BLN8),.WL(WL219));
sram_cell_6t_5 inst_cell_219_9 (.BL(BL9),.BLN(BLN9),.WL(WL219));
sram_cell_6t_5 inst_cell_219_10 (.BL(BL10),.BLN(BLN10),.WL(WL219));
sram_cell_6t_5 inst_cell_219_11 (.BL(BL11),.BLN(BLN11),.WL(WL219));
sram_cell_6t_5 inst_cell_219_12 (.BL(BL12),.BLN(BLN12),.WL(WL219));
sram_cell_6t_5 inst_cell_219_13 (.BL(BL13),.BLN(BLN13),.WL(WL219));
sram_cell_6t_5 inst_cell_219_14 (.BL(BL14),.BLN(BLN14),.WL(WL219));
sram_cell_6t_5 inst_cell_219_15 (.BL(BL15),.BLN(BLN15),.WL(WL219));
sram_cell_6t_5 inst_cell_219_16 (.BL(BL16),.BLN(BLN16),.WL(WL219));
sram_cell_6t_5 inst_cell_219_17 (.BL(BL17),.BLN(BLN17),.WL(WL219));
sram_cell_6t_5 inst_cell_219_18 (.BL(BL18),.BLN(BLN18),.WL(WL219));
sram_cell_6t_5 inst_cell_219_19 (.BL(BL19),.BLN(BLN19),.WL(WL219));
sram_cell_6t_5 inst_cell_219_20 (.BL(BL20),.BLN(BLN20),.WL(WL219));
sram_cell_6t_5 inst_cell_219_21 (.BL(BL21),.BLN(BLN21),.WL(WL219));
sram_cell_6t_5 inst_cell_219_22 (.BL(BL22),.BLN(BLN22),.WL(WL219));
sram_cell_6t_5 inst_cell_219_23 (.BL(BL23),.BLN(BLN23),.WL(WL219));
sram_cell_6t_5 inst_cell_219_24 (.BL(BL24),.BLN(BLN24),.WL(WL219));
sram_cell_6t_5 inst_cell_219_25 (.BL(BL25),.BLN(BLN25),.WL(WL219));
sram_cell_6t_5 inst_cell_219_26 (.BL(BL26),.BLN(BLN26),.WL(WL219));
sram_cell_6t_5 inst_cell_219_27 (.BL(BL27),.BLN(BLN27),.WL(WL219));
sram_cell_6t_5 inst_cell_219_28 (.BL(BL28),.BLN(BLN28),.WL(WL219));
sram_cell_6t_5 inst_cell_219_29 (.BL(BL29),.BLN(BLN29),.WL(WL219));
sram_cell_6t_5 inst_cell_219_30 (.BL(BL30),.BLN(BLN30),.WL(WL219));
sram_cell_6t_5 inst_cell_219_31 (.BL(BL31),.BLN(BLN31),.WL(WL219));
sram_cell_6t_5 inst_cell_219_32 (.BL(BL32),.BLN(BLN32),.WL(WL219));
sram_cell_6t_5 inst_cell_219_33 (.BL(BL33),.BLN(BLN33),.WL(WL219));
sram_cell_6t_5 inst_cell_219_34 (.BL(BL34),.BLN(BLN34),.WL(WL219));
sram_cell_6t_5 inst_cell_219_35 (.BL(BL35),.BLN(BLN35),.WL(WL219));
sram_cell_6t_5 inst_cell_219_36 (.BL(BL36),.BLN(BLN36),.WL(WL219));
sram_cell_6t_5 inst_cell_219_37 (.BL(BL37),.BLN(BLN37),.WL(WL219));
sram_cell_6t_5 inst_cell_219_38 (.BL(BL38),.BLN(BLN38),.WL(WL219));
sram_cell_6t_5 inst_cell_219_39 (.BL(BL39),.BLN(BLN39),.WL(WL219));
sram_cell_6t_5 inst_cell_219_40 (.BL(BL40),.BLN(BLN40),.WL(WL219));
sram_cell_6t_5 inst_cell_219_41 (.BL(BL41),.BLN(BLN41),.WL(WL219));
sram_cell_6t_5 inst_cell_219_42 (.BL(BL42),.BLN(BLN42),.WL(WL219));
sram_cell_6t_5 inst_cell_219_43 (.BL(BL43),.BLN(BLN43),.WL(WL219));
sram_cell_6t_5 inst_cell_219_44 (.BL(BL44),.BLN(BLN44),.WL(WL219));
sram_cell_6t_5 inst_cell_219_45 (.BL(BL45),.BLN(BLN45),.WL(WL219));
sram_cell_6t_5 inst_cell_219_46 (.BL(BL46),.BLN(BLN46),.WL(WL219));
sram_cell_6t_5 inst_cell_219_47 (.BL(BL47),.BLN(BLN47),.WL(WL219));
sram_cell_6t_5 inst_cell_219_48 (.BL(BL48),.BLN(BLN48),.WL(WL219));
sram_cell_6t_5 inst_cell_219_49 (.BL(BL49),.BLN(BLN49),.WL(WL219));
sram_cell_6t_5 inst_cell_219_50 (.BL(BL50),.BLN(BLN50),.WL(WL219));
sram_cell_6t_5 inst_cell_219_51 (.BL(BL51),.BLN(BLN51),.WL(WL219));
sram_cell_6t_5 inst_cell_219_52 (.BL(BL52),.BLN(BLN52),.WL(WL219));
sram_cell_6t_5 inst_cell_219_53 (.BL(BL53),.BLN(BLN53),.WL(WL219));
sram_cell_6t_5 inst_cell_219_54 (.BL(BL54),.BLN(BLN54),.WL(WL219));
sram_cell_6t_5 inst_cell_219_55 (.BL(BL55),.BLN(BLN55),.WL(WL219));
sram_cell_6t_5 inst_cell_219_56 (.BL(BL56),.BLN(BLN56),.WL(WL219));
sram_cell_6t_5 inst_cell_219_57 (.BL(BL57),.BLN(BLN57),.WL(WL219));
sram_cell_6t_5 inst_cell_219_58 (.BL(BL58),.BLN(BLN58),.WL(WL219));
sram_cell_6t_5 inst_cell_219_59 (.BL(BL59),.BLN(BLN59),.WL(WL219));
sram_cell_6t_5 inst_cell_219_60 (.BL(BL60),.BLN(BLN60),.WL(WL219));
sram_cell_6t_5 inst_cell_219_61 (.BL(BL61),.BLN(BLN61),.WL(WL219));
sram_cell_6t_5 inst_cell_219_62 (.BL(BL62),.BLN(BLN62),.WL(WL219));
sram_cell_6t_5 inst_cell_219_63 (.BL(BL63),.BLN(BLN63),.WL(WL219));
sram_cell_6t_5 inst_cell_219_64 (.BL(BL64),.BLN(BLN64),.WL(WL219));
sram_cell_6t_5 inst_cell_219_65 (.BL(BL65),.BLN(BLN65),.WL(WL219));
sram_cell_6t_5 inst_cell_219_66 (.BL(BL66),.BLN(BLN66),.WL(WL219));
sram_cell_6t_5 inst_cell_219_67 (.BL(BL67),.BLN(BLN67),.WL(WL219));
sram_cell_6t_5 inst_cell_219_68 (.BL(BL68),.BLN(BLN68),.WL(WL219));
sram_cell_6t_5 inst_cell_219_69 (.BL(BL69),.BLN(BLN69),.WL(WL219));
sram_cell_6t_5 inst_cell_219_70 (.BL(BL70),.BLN(BLN70),.WL(WL219));
sram_cell_6t_5 inst_cell_219_71 (.BL(BL71),.BLN(BLN71),.WL(WL219));
sram_cell_6t_5 inst_cell_219_72 (.BL(BL72),.BLN(BLN72),.WL(WL219));
sram_cell_6t_5 inst_cell_219_73 (.BL(BL73),.BLN(BLN73),.WL(WL219));
sram_cell_6t_5 inst_cell_219_74 (.BL(BL74),.BLN(BLN74),.WL(WL219));
sram_cell_6t_5 inst_cell_219_75 (.BL(BL75),.BLN(BLN75),.WL(WL219));
sram_cell_6t_5 inst_cell_219_76 (.BL(BL76),.BLN(BLN76),.WL(WL219));
sram_cell_6t_5 inst_cell_219_77 (.BL(BL77),.BLN(BLN77),.WL(WL219));
sram_cell_6t_5 inst_cell_219_78 (.BL(BL78),.BLN(BLN78),.WL(WL219));
sram_cell_6t_5 inst_cell_219_79 (.BL(BL79),.BLN(BLN79),.WL(WL219));
sram_cell_6t_5 inst_cell_219_80 (.BL(BL80),.BLN(BLN80),.WL(WL219));
sram_cell_6t_5 inst_cell_219_81 (.BL(BL81),.BLN(BLN81),.WL(WL219));
sram_cell_6t_5 inst_cell_219_82 (.BL(BL82),.BLN(BLN82),.WL(WL219));
sram_cell_6t_5 inst_cell_219_83 (.BL(BL83),.BLN(BLN83),.WL(WL219));
sram_cell_6t_5 inst_cell_219_84 (.BL(BL84),.BLN(BLN84),.WL(WL219));
sram_cell_6t_5 inst_cell_219_85 (.BL(BL85),.BLN(BLN85),.WL(WL219));
sram_cell_6t_5 inst_cell_219_86 (.BL(BL86),.BLN(BLN86),.WL(WL219));
sram_cell_6t_5 inst_cell_219_87 (.BL(BL87),.BLN(BLN87),.WL(WL219));
sram_cell_6t_5 inst_cell_219_88 (.BL(BL88),.BLN(BLN88),.WL(WL219));
sram_cell_6t_5 inst_cell_219_89 (.BL(BL89),.BLN(BLN89),.WL(WL219));
sram_cell_6t_5 inst_cell_219_90 (.BL(BL90),.BLN(BLN90),.WL(WL219));
sram_cell_6t_5 inst_cell_219_91 (.BL(BL91),.BLN(BLN91),.WL(WL219));
sram_cell_6t_5 inst_cell_219_92 (.BL(BL92),.BLN(BLN92),.WL(WL219));
sram_cell_6t_5 inst_cell_219_93 (.BL(BL93),.BLN(BLN93),.WL(WL219));
sram_cell_6t_5 inst_cell_219_94 (.BL(BL94),.BLN(BLN94),.WL(WL219));
sram_cell_6t_5 inst_cell_219_95 (.BL(BL95),.BLN(BLN95),.WL(WL219));
sram_cell_6t_5 inst_cell_219_96 (.BL(BL96),.BLN(BLN96),.WL(WL219));
sram_cell_6t_5 inst_cell_219_97 (.BL(BL97),.BLN(BLN97),.WL(WL219));
sram_cell_6t_5 inst_cell_219_98 (.BL(BL98),.BLN(BLN98),.WL(WL219));
sram_cell_6t_5 inst_cell_219_99 (.BL(BL99),.BLN(BLN99),.WL(WL219));
sram_cell_6t_5 inst_cell_219_100 (.BL(BL100),.BLN(BLN100),.WL(WL219));
sram_cell_6t_5 inst_cell_219_101 (.BL(BL101),.BLN(BLN101),.WL(WL219));
sram_cell_6t_5 inst_cell_219_102 (.BL(BL102),.BLN(BLN102),.WL(WL219));
sram_cell_6t_5 inst_cell_219_103 (.BL(BL103),.BLN(BLN103),.WL(WL219));
sram_cell_6t_5 inst_cell_219_104 (.BL(BL104),.BLN(BLN104),.WL(WL219));
sram_cell_6t_5 inst_cell_219_105 (.BL(BL105),.BLN(BLN105),.WL(WL219));
sram_cell_6t_5 inst_cell_219_106 (.BL(BL106),.BLN(BLN106),.WL(WL219));
sram_cell_6t_5 inst_cell_219_107 (.BL(BL107),.BLN(BLN107),.WL(WL219));
sram_cell_6t_5 inst_cell_219_108 (.BL(BL108),.BLN(BLN108),.WL(WL219));
sram_cell_6t_5 inst_cell_219_109 (.BL(BL109),.BLN(BLN109),.WL(WL219));
sram_cell_6t_5 inst_cell_219_110 (.BL(BL110),.BLN(BLN110),.WL(WL219));
sram_cell_6t_5 inst_cell_219_111 (.BL(BL111),.BLN(BLN111),.WL(WL219));
sram_cell_6t_5 inst_cell_219_112 (.BL(BL112),.BLN(BLN112),.WL(WL219));
sram_cell_6t_5 inst_cell_219_113 (.BL(BL113),.BLN(BLN113),.WL(WL219));
sram_cell_6t_5 inst_cell_219_114 (.BL(BL114),.BLN(BLN114),.WL(WL219));
sram_cell_6t_5 inst_cell_219_115 (.BL(BL115),.BLN(BLN115),.WL(WL219));
sram_cell_6t_5 inst_cell_219_116 (.BL(BL116),.BLN(BLN116),.WL(WL219));
sram_cell_6t_5 inst_cell_219_117 (.BL(BL117),.BLN(BLN117),.WL(WL219));
sram_cell_6t_5 inst_cell_219_118 (.BL(BL118),.BLN(BLN118),.WL(WL219));
sram_cell_6t_5 inst_cell_219_119 (.BL(BL119),.BLN(BLN119),.WL(WL219));
sram_cell_6t_5 inst_cell_219_120 (.BL(BL120),.BLN(BLN120),.WL(WL219));
sram_cell_6t_5 inst_cell_219_121 (.BL(BL121),.BLN(BLN121),.WL(WL219));
sram_cell_6t_5 inst_cell_219_122 (.BL(BL122),.BLN(BLN122),.WL(WL219));
sram_cell_6t_5 inst_cell_219_123 (.BL(BL123),.BLN(BLN123),.WL(WL219));
sram_cell_6t_5 inst_cell_219_124 (.BL(BL124),.BLN(BLN124),.WL(WL219));
sram_cell_6t_5 inst_cell_219_125 (.BL(BL125),.BLN(BLN125),.WL(WL219));
sram_cell_6t_5 inst_cell_219_126 (.BL(BL126),.BLN(BLN126),.WL(WL219));
sram_cell_6t_5 inst_cell_219_127 (.BL(BL127),.BLN(BLN127),.WL(WL219));
sram_cell_6t_5 inst_cell_220_0 (.BL(BL0),.BLN(BLN0),.WL(WL220));
sram_cell_6t_5 inst_cell_220_1 (.BL(BL1),.BLN(BLN1),.WL(WL220));
sram_cell_6t_5 inst_cell_220_2 (.BL(BL2),.BLN(BLN2),.WL(WL220));
sram_cell_6t_5 inst_cell_220_3 (.BL(BL3),.BLN(BLN3),.WL(WL220));
sram_cell_6t_5 inst_cell_220_4 (.BL(BL4),.BLN(BLN4),.WL(WL220));
sram_cell_6t_5 inst_cell_220_5 (.BL(BL5),.BLN(BLN5),.WL(WL220));
sram_cell_6t_5 inst_cell_220_6 (.BL(BL6),.BLN(BLN6),.WL(WL220));
sram_cell_6t_5 inst_cell_220_7 (.BL(BL7),.BLN(BLN7),.WL(WL220));
sram_cell_6t_5 inst_cell_220_8 (.BL(BL8),.BLN(BLN8),.WL(WL220));
sram_cell_6t_5 inst_cell_220_9 (.BL(BL9),.BLN(BLN9),.WL(WL220));
sram_cell_6t_5 inst_cell_220_10 (.BL(BL10),.BLN(BLN10),.WL(WL220));
sram_cell_6t_5 inst_cell_220_11 (.BL(BL11),.BLN(BLN11),.WL(WL220));
sram_cell_6t_5 inst_cell_220_12 (.BL(BL12),.BLN(BLN12),.WL(WL220));
sram_cell_6t_5 inst_cell_220_13 (.BL(BL13),.BLN(BLN13),.WL(WL220));
sram_cell_6t_5 inst_cell_220_14 (.BL(BL14),.BLN(BLN14),.WL(WL220));
sram_cell_6t_5 inst_cell_220_15 (.BL(BL15),.BLN(BLN15),.WL(WL220));
sram_cell_6t_5 inst_cell_220_16 (.BL(BL16),.BLN(BLN16),.WL(WL220));
sram_cell_6t_5 inst_cell_220_17 (.BL(BL17),.BLN(BLN17),.WL(WL220));
sram_cell_6t_5 inst_cell_220_18 (.BL(BL18),.BLN(BLN18),.WL(WL220));
sram_cell_6t_5 inst_cell_220_19 (.BL(BL19),.BLN(BLN19),.WL(WL220));
sram_cell_6t_5 inst_cell_220_20 (.BL(BL20),.BLN(BLN20),.WL(WL220));
sram_cell_6t_5 inst_cell_220_21 (.BL(BL21),.BLN(BLN21),.WL(WL220));
sram_cell_6t_5 inst_cell_220_22 (.BL(BL22),.BLN(BLN22),.WL(WL220));
sram_cell_6t_5 inst_cell_220_23 (.BL(BL23),.BLN(BLN23),.WL(WL220));
sram_cell_6t_5 inst_cell_220_24 (.BL(BL24),.BLN(BLN24),.WL(WL220));
sram_cell_6t_5 inst_cell_220_25 (.BL(BL25),.BLN(BLN25),.WL(WL220));
sram_cell_6t_5 inst_cell_220_26 (.BL(BL26),.BLN(BLN26),.WL(WL220));
sram_cell_6t_5 inst_cell_220_27 (.BL(BL27),.BLN(BLN27),.WL(WL220));
sram_cell_6t_5 inst_cell_220_28 (.BL(BL28),.BLN(BLN28),.WL(WL220));
sram_cell_6t_5 inst_cell_220_29 (.BL(BL29),.BLN(BLN29),.WL(WL220));
sram_cell_6t_5 inst_cell_220_30 (.BL(BL30),.BLN(BLN30),.WL(WL220));
sram_cell_6t_5 inst_cell_220_31 (.BL(BL31),.BLN(BLN31),.WL(WL220));
sram_cell_6t_5 inst_cell_220_32 (.BL(BL32),.BLN(BLN32),.WL(WL220));
sram_cell_6t_5 inst_cell_220_33 (.BL(BL33),.BLN(BLN33),.WL(WL220));
sram_cell_6t_5 inst_cell_220_34 (.BL(BL34),.BLN(BLN34),.WL(WL220));
sram_cell_6t_5 inst_cell_220_35 (.BL(BL35),.BLN(BLN35),.WL(WL220));
sram_cell_6t_5 inst_cell_220_36 (.BL(BL36),.BLN(BLN36),.WL(WL220));
sram_cell_6t_5 inst_cell_220_37 (.BL(BL37),.BLN(BLN37),.WL(WL220));
sram_cell_6t_5 inst_cell_220_38 (.BL(BL38),.BLN(BLN38),.WL(WL220));
sram_cell_6t_5 inst_cell_220_39 (.BL(BL39),.BLN(BLN39),.WL(WL220));
sram_cell_6t_5 inst_cell_220_40 (.BL(BL40),.BLN(BLN40),.WL(WL220));
sram_cell_6t_5 inst_cell_220_41 (.BL(BL41),.BLN(BLN41),.WL(WL220));
sram_cell_6t_5 inst_cell_220_42 (.BL(BL42),.BLN(BLN42),.WL(WL220));
sram_cell_6t_5 inst_cell_220_43 (.BL(BL43),.BLN(BLN43),.WL(WL220));
sram_cell_6t_5 inst_cell_220_44 (.BL(BL44),.BLN(BLN44),.WL(WL220));
sram_cell_6t_5 inst_cell_220_45 (.BL(BL45),.BLN(BLN45),.WL(WL220));
sram_cell_6t_5 inst_cell_220_46 (.BL(BL46),.BLN(BLN46),.WL(WL220));
sram_cell_6t_5 inst_cell_220_47 (.BL(BL47),.BLN(BLN47),.WL(WL220));
sram_cell_6t_5 inst_cell_220_48 (.BL(BL48),.BLN(BLN48),.WL(WL220));
sram_cell_6t_5 inst_cell_220_49 (.BL(BL49),.BLN(BLN49),.WL(WL220));
sram_cell_6t_5 inst_cell_220_50 (.BL(BL50),.BLN(BLN50),.WL(WL220));
sram_cell_6t_5 inst_cell_220_51 (.BL(BL51),.BLN(BLN51),.WL(WL220));
sram_cell_6t_5 inst_cell_220_52 (.BL(BL52),.BLN(BLN52),.WL(WL220));
sram_cell_6t_5 inst_cell_220_53 (.BL(BL53),.BLN(BLN53),.WL(WL220));
sram_cell_6t_5 inst_cell_220_54 (.BL(BL54),.BLN(BLN54),.WL(WL220));
sram_cell_6t_5 inst_cell_220_55 (.BL(BL55),.BLN(BLN55),.WL(WL220));
sram_cell_6t_5 inst_cell_220_56 (.BL(BL56),.BLN(BLN56),.WL(WL220));
sram_cell_6t_5 inst_cell_220_57 (.BL(BL57),.BLN(BLN57),.WL(WL220));
sram_cell_6t_5 inst_cell_220_58 (.BL(BL58),.BLN(BLN58),.WL(WL220));
sram_cell_6t_5 inst_cell_220_59 (.BL(BL59),.BLN(BLN59),.WL(WL220));
sram_cell_6t_5 inst_cell_220_60 (.BL(BL60),.BLN(BLN60),.WL(WL220));
sram_cell_6t_5 inst_cell_220_61 (.BL(BL61),.BLN(BLN61),.WL(WL220));
sram_cell_6t_5 inst_cell_220_62 (.BL(BL62),.BLN(BLN62),.WL(WL220));
sram_cell_6t_5 inst_cell_220_63 (.BL(BL63),.BLN(BLN63),.WL(WL220));
sram_cell_6t_5 inst_cell_220_64 (.BL(BL64),.BLN(BLN64),.WL(WL220));
sram_cell_6t_5 inst_cell_220_65 (.BL(BL65),.BLN(BLN65),.WL(WL220));
sram_cell_6t_5 inst_cell_220_66 (.BL(BL66),.BLN(BLN66),.WL(WL220));
sram_cell_6t_5 inst_cell_220_67 (.BL(BL67),.BLN(BLN67),.WL(WL220));
sram_cell_6t_5 inst_cell_220_68 (.BL(BL68),.BLN(BLN68),.WL(WL220));
sram_cell_6t_5 inst_cell_220_69 (.BL(BL69),.BLN(BLN69),.WL(WL220));
sram_cell_6t_5 inst_cell_220_70 (.BL(BL70),.BLN(BLN70),.WL(WL220));
sram_cell_6t_5 inst_cell_220_71 (.BL(BL71),.BLN(BLN71),.WL(WL220));
sram_cell_6t_5 inst_cell_220_72 (.BL(BL72),.BLN(BLN72),.WL(WL220));
sram_cell_6t_5 inst_cell_220_73 (.BL(BL73),.BLN(BLN73),.WL(WL220));
sram_cell_6t_5 inst_cell_220_74 (.BL(BL74),.BLN(BLN74),.WL(WL220));
sram_cell_6t_5 inst_cell_220_75 (.BL(BL75),.BLN(BLN75),.WL(WL220));
sram_cell_6t_5 inst_cell_220_76 (.BL(BL76),.BLN(BLN76),.WL(WL220));
sram_cell_6t_5 inst_cell_220_77 (.BL(BL77),.BLN(BLN77),.WL(WL220));
sram_cell_6t_5 inst_cell_220_78 (.BL(BL78),.BLN(BLN78),.WL(WL220));
sram_cell_6t_5 inst_cell_220_79 (.BL(BL79),.BLN(BLN79),.WL(WL220));
sram_cell_6t_5 inst_cell_220_80 (.BL(BL80),.BLN(BLN80),.WL(WL220));
sram_cell_6t_5 inst_cell_220_81 (.BL(BL81),.BLN(BLN81),.WL(WL220));
sram_cell_6t_5 inst_cell_220_82 (.BL(BL82),.BLN(BLN82),.WL(WL220));
sram_cell_6t_5 inst_cell_220_83 (.BL(BL83),.BLN(BLN83),.WL(WL220));
sram_cell_6t_5 inst_cell_220_84 (.BL(BL84),.BLN(BLN84),.WL(WL220));
sram_cell_6t_5 inst_cell_220_85 (.BL(BL85),.BLN(BLN85),.WL(WL220));
sram_cell_6t_5 inst_cell_220_86 (.BL(BL86),.BLN(BLN86),.WL(WL220));
sram_cell_6t_5 inst_cell_220_87 (.BL(BL87),.BLN(BLN87),.WL(WL220));
sram_cell_6t_5 inst_cell_220_88 (.BL(BL88),.BLN(BLN88),.WL(WL220));
sram_cell_6t_5 inst_cell_220_89 (.BL(BL89),.BLN(BLN89),.WL(WL220));
sram_cell_6t_5 inst_cell_220_90 (.BL(BL90),.BLN(BLN90),.WL(WL220));
sram_cell_6t_5 inst_cell_220_91 (.BL(BL91),.BLN(BLN91),.WL(WL220));
sram_cell_6t_5 inst_cell_220_92 (.BL(BL92),.BLN(BLN92),.WL(WL220));
sram_cell_6t_5 inst_cell_220_93 (.BL(BL93),.BLN(BLN93),.WL(WL220));
sram_cell_6t_5 inst_cell_220_94 (.BL(BL94),.BLN(BLN94),.WL(WL220));
sram_cell_6t_5 inst_cell_220_95 (.BL(BL95),.BLN(BLN95),.WL(WL220));
sram_cell_6t_5 inst_cell_220_96 (.BL(BL96),.BLN(BLN96),.WL(WL220));
sram_cell_6t_5 inst_cell_220_97 (.BL(BL97),.BLN(BLN97),.WL(WL220));
sram_cell_6t_5 inst_cell_220_98 (.BL(BL98),.BLN(BLN98),.WL(WL220));
sram_cell_6t_5 inst_cell_220_99 (.BL(BL99),.BLN(BLN99),.WL(WL220));
sram_cell_6t_5 inst_cell_220_100 (.BL(BL100),.BLN(BLN100),.WL(WL220));
sram_cell_6t_5 inst_cell_220_101 (.BL(BL101),.BLN(BLN101),.WL(WL220));
sram_cell_6t_5 inst_cell_220_102 (.BL(BL102),.BLN(BLN102),.WL(WL220));
sram_cell_6t_5 inst_cell_220_103 (.BL(BL103),.BLN(BLN103),.WL(WL220));
sram_cell_6t_5 inst_cell_220_104 (.BL(BL104),.BLN(BLN104),.WL(WL220));
sram_cell_6t_5 inst_cell_220_105 (.BL(BL105),.BLN(BLN105),.WL(WL220));
sram_cell_6t_5 inst_cell_220_106 (.BL(BL106),.BLN(BLN106),.WL(WL220));
sram_cell_6t_5 inst_cell_220_107 (.BL(BL107),.BLN(BLN107),.WL(WL220));
sram_cell_6t_5 inst_cell_220_108 (.BL(BL108),.BLN(BLN108),.WL(WL220));
sram_cell_6t_5 inst_cell_220_109 (.BL(BL109),.BLN(BLN109),.WL(WL220));
sram_cell_6t_5 inst_cell_220_110 (.BL(BL110),.BLN(BLN110),.WL(WL220));
sram_cell_6t_5 inst_cell_220_111 (.BL(BL111),.BLN(BLN111),.WL(WL220));
sram_cell_6t_5 inst_cell_220_112 (.BL(BL112),.BLN(BLN112),.WL(WL220));
sram_cell_6t_5 inst_cell_220_113 (.BL(BL113),.BLN(BLN113),.WL(WL220));
sram_cell_6t_5 inst_cell_220_114 (.BL(BL114),.BLN(BLN114),.WL(WL220));
sram_cell_6t_5 inst_cell_220_115 (.BL(BL115),.BLN(BLN115),.WL(WL220));
sram_cell_6t_5 inst_cell_220_116 (.BL(BL116),.BLN(BLN116),.WL(WL220));
sram_cell_6t_5 inst_cell_220_117 (.BL(BL117),.BLN(BLN117),.WL(WL220));
sram_cell_6t_5 inst_cell_220_118 (.BL(BL118),.BLN(BLN118),.WL(WL220));
sram_cell_6t_5 inst_cell_220_119 (.BL(BL119),.BLN(BLN119),.WL(WL220));
sram_cell_6t_5 inst_cell_220_120 (.BL(BL120),.BLN(BLN120),.WL(WL220));
sram_cell_6t_5 inst_cell_220_121 (.BL(BL121),.BLN(BLN121),.WL(WL220));
sram_cell_6t_5 inst_cell_220_122 (.BL(BL122),.BLN(BLN122),.WL(WL220));
sram_cell_6t_5 inst_cell_220_123 (.BL(BL123),.BLN(BLN123),.WL(WL220));
sram_cell_6t_5 inst_cell_220_124 (.BL(BL124),.BLN(BLN124),.WL(WL220));
sram_cell_6t_5 inst_cell_220_125 (.BL(BL125),.BLN(BLN125),.WL(WL220));
sram_cell_6t_5 inst_cell_220_126 (.BL(BL126),.BLN(BLN126),.WL(WL220));
sram_cell_6t_5 inst_cell_220_127 (.BL(BL127),.BLN(BLN127),.WL(WL220));
sram_cell_6t_5 inst_cell_221_0 (.BL(BL0),.BLN(BLN0),.WL(WL221));
sram_cell_6t_5 inst_cell_221_1 (.BL(BL1),.BLN(BLN1),.WL(WL221));
sram_cell_6t_5 inst_cell_221_2 (.BL(BL2),.BLN(BLN2),.WL(WL221));
sram_cell_6t_5 inst_cell_221_3 (.BL(BL3),.BLN(BLN3),.WL(WL221));
sram_cell_6t_5 inst_cell_221_4 (.BL(BL4),.BLN(BLN4),.WL(WL221));
sram_cell_6t_5 inst_cell_221_5 (.BL(BL5),.BLN(BLN5),.WL(WL221));
sram_cell_6t_5 inst_cell_221_6 (.BL(BL6),.BLN(BLN6),.WL(WL221));
sram_cell_6t_5 inst_cell_221_7 (.BL(BL7),.BLN(BLN7),.WL(WL221));
sram_cell_6t_5 inst_cell_221_8 (.BL(BL8),.BLN(BLN8),.WL(WL221));
sram_cell_6t_5 inst_cell_221_9 (.BL(BL9),.BLN(BLN9),.WL(WL221));
sram_cell_6t_5 inst_cell_221_10 (.BL(BL10),.BLN(BLN10),.WL(WL221));
sram_cell_6t_5 inst_cell_221_11 (.BL(BL11),.BLN(BLN11),.WL(WL221));
sram_cell_6t_5 inst_cell_221_12 (.BL(BL12),.BLN(BLN12),.WL(WL221));
sram_cell_6t_5 inst_cell_221_13 (.BL(BL13),.BLN(BLN13),.WL(WL221));
sram_cell_6t_5 inst_cell_221_14 (.BL(BL14),.BLN(BLN14),.WL(WL221));
sram_cell_6t_5 inst_cell_221_15 (.BL(BL15),.BLN(BLN15),.WL(WL221));
sram_cell_6t_5 inst_cell_221_16 (.BL(BL16),.BLN(BLN16),.WL(WL221));
sram_cell_6t_5 inst_cell_221_17 (.BL(BL17),.BLN(BLN17),.WL(WL221));
sram_cell_6t_5 inst_cell_221_18 (.BL(BL18),.BLN(BLN18),.WL(WL221));
sram_cell_6t_5 inst_cell_221_19 (.BL(BL19),.BLN(BLN19),.WL(WL221));
sram_cell_6t_5 inst_cell_221_20 (.BL(BL20),.BLN(BLN20),.WL(WL221));
sram_cell_6t_5 inst_cell_221_21 (.BL(BL21),.BLN(BLN21),.WL(WL221));
sram_cell_6t_5 inst_cell_221_22 (.BL(BL22),.BLN(BLN22),.WL(WL221));
sram_cell_6t_5 inst_cell_221_23 (.BL(BL23),.BLN(BLN23),.WL(WL221));
sram_cell_6t_5 inst_cell_221_24 (.BL(BL24),.BLN(BLN24),.WL(WL221));
sram_cell_6t_5 inst_cell_221_25 (.BL(BL25),.BLN(BLN25),.WL(WL221));
sram_cell_6t_5 inst_cell_221_26 (.BL(BL26),.BLN(BLN26),.WL(WL221));
sram_cell_6t_5 inst_cell_221_27 (.BL(BL27),.BLN(BLN27),.WL(WL221));
sram_cell_6t_5 inst_cell_221_28 (.BL(BL28),.BLN(BLN28),.WL(WL221));
sram_cell_6t_5 inst_cell_221_29 (.BL(BL29),.BLN(BLN29),.WL(WL221));
sram_cell_6t_5 inst_cell_221_30 (.BL(BL30),.BLN(BLN30),.WL(WL221));
sram_cell_6t_5 inst_cell_221_31 (.BL(BL31),.BLN(BLN31),.WL(WL221));
sram_cell_6t_5 inst_cell_221_32 (.BL(BL32),.BLN(BLN32),.WL(WL221));
sram_cell_6t_5 inst_cell_221_33 (.BL(BL33),.BLN(BLN33),.WL(WL221));
sram_cell_6t_5 inst_cell_221_34 (.BL(BL34),.BLN(BLN34),.WL(WL221));
sram_cell_6t_5 inst_cell_221_35 (.BL(BL35),.BLN(BLN35),.WL(WL221));
sram_cell_6t_5 inst_cell_221_36 (.BL(BL36),.BLN(BLN36),.WL(WL221));
sram_cell_6t_5 inst_cell_221_37 (.BL(BL37),.BLN(BLN37),.WL(WL221));
sram_cell_6t_5 inst_cell_221_38 (.BL(BL38),.BLN(BLN38),.WL(WL221));
sram_cell_6t_5 inst_cell_221_39 (.BL(BL39),.BLN(BLN39),.WL(WL221));
sram_cell_6t_5 inst_cell_221_40 (.BL(BL40),.BLN(BLN40),.WL(WL221));
sram_cell_6t_5 inst_cell_221_41 (.BL(BL41),.BLN(BLN41),.WL(WL221));
sram_cell_6t_5 inst_cell_221_42 (.BL(BL42),.BLN(BLN42),.WL(WL221));
sram_cell_6t_5 inst_cell_221_43 (.BL(BL43),.BLN(BLN43),.WL(WL221));
sram_cell_6t_5 inst_cell_221_44 (.BL(BL44),.BLN(BLN44),.WL(WL221));
sram_cell_6t_5 inst_cell_221_45 (.BL(BL45),.BLN(BLN45),.WL(WL221));
sram_cell_6t_5 inst_cell_221_46 (.BL(BL46),.BLN(BLN46),.WL(WL221));
sram_cell_6t_5 inst_cell_221_47 (.BL(BL47),.BLN(BLN47),.WL(WL221));
sram_cell_6t_5 inst_cell_221_48 (.BL(BL48),.BLN(BLN48),.WL(WL221));
sram_cell_6t_5 inst_cell_221_49 (.BL(BL49),.BLN(BLN49),.WL(WL221));
sram_cell_6t_5 inst_cell_221_50 (.BL(BL50),.BLN(BLN50),.WL(WL221));
sram_cell_6t_5 inst_cell_221_51 (.BL(BL51),.BLN(BLN51),.WL(WL221));
sram_cell_6t_5 inst_cell_221_52 (.BL(BL52),.BLN(BLN52),.WL(WL221));
sram_cell_6t_5 inst_cell_221_53 (.BL(BL53),.BLN(BLN53),.WL(WL221));
sram_cell_6t_5 inst_cell_221_54 (.BL(BL54),.BLN(BLN54),.WL(WL221));
sram_cell_6t_5 inst_cell_221_55 (.BL(BL55),.BLN(BLN55),.WL(WL221));
sram_cell_6t_5 inst_cell_221_56 (.BL(BL56),.BLN(BLN56),.WL(WL221));
sram_cell_6t_5 inst_cell_221_57 (.BL(BL57),.BLN(BLN57),.WL(WL221));
sram_cell_6t_5 inst_cell_221_58 (.BL(BL58),.BLN(BLN58),.WL(WL221));
sram_cell_6t_5 inst_cell_221_59 (.BL(BL59),.BLN(BLN59),.WL(WL221));
sram_cell_6t_5 inst_cell_221_60 (.BL(BL60),.BLN(BLN60),.WL(WL221));
sram_cell_6t_5 inst_cell_221_61 (.BL(BL61),.BLN(BLN61),.WL(WL221));
sram_cell_6t_5 inst_cell_221_62 (.BL(BL62),.BLN(BLN62),.WL(WL221));
sram_cell_6t_5 inst_cell_221_63 (.BL(BL63),.BLN(BLN63),.WL(WL221));
sram_cell_6t_5 inst_cell_221_64 (.BL(BL64),.BLN(BLN64),.WL(WL221));
sram_cell_6t_5 inst_cell_221_65 (.BL(BL65),.BLN(BLN65),.WL(WL221));
sram_cell_6t_5 inst_cell_221_66 (.BL(BL66),.BLN(BLN66),.WL(WL221));
sram_cell_6t_5 inst_cell_221_67 (.BL(BL67),.BLN(BLN67),.WL(WL221));
sram_cell_6t_5 inst_cell_221_68 (.BL(BL68),.BLN(BLN68),.WL(WL221));
sram_cell_6t_5 inst_cell_221_69 (.BL(BL69),.BLN(BLN69),.WL(WL221));
sram_cell_6t_5 inst_cell_221_70 (.BL(BL70),.BLN(BLN70),.WL(WL221));
sram_cell_6t_5 inst_cell_221_71 (.BL(BL71),.BLN(BLN71),.WL(WL221));
sram_cell_6t_5 inst_cell_221_72 (.BL(BL72),.BLN(BLN72),.WL(WL221));
sram_cell_6t_5 inst_cell_221_73 (.BL(BL73),.BLN(BLN73),.WL(WL221));
sram_cell_6t_5 inst_cell_221_74 (.BL(BL74),.BLN(BLN74),.WL(WL221));
sram_cell_6t_5 inst_cell_221_75 (.BL(BL75),.BLN(BLN75),.WL(WL221));
sram_cell_6t_5 inst_cell_221_76 (.BL(BL76),.BLN(BLN76),.WL(WL221));
sram_cell_6t_5 inst_cell_221_77 (.BL(BL77),.BLN(BLN77),.WL(WL221));
sram_cell_6t_5 inst_cell_221_78 (.BL(BL78),.BLN(BLN78),.WL(WL221));
sram_cell_6t_5 inst_cell_221_79 (.BL(BL79),.BLN(BLN79),.WL(WL221));
sram_cell_6t_5 inst_cell_221_80 (.BL(BL80),.BLN(BLN80),.WL(WL221));
sram_cell_6t_5 inst_cell_221_81 (.BL(BL81),.BLN(BLN81),.WL(WL221));
sram_cell_6t_5 inst_cell_221_82 (.BL(BL82),.BLN(BLN82),.WL(WL221));
sram_cell_6t_5 inst_cell_221_83 (.BL(BL83),.BLN(BLN83),.WL(WL221));
sram_cell_6t_5 inst_cell_221_84 (.BL(BL84),.BLN(BLN84),.WL(WL221));
sram_cell_6t_5 inst_cell_221_85 (.BL(BL85),.BLN(BLN85),.WL(WL221));
sram_cell_6t_5 inst_cell_221_86 (.BL(BL86),.BLN(BLN86),.WL(WL221));
sram_cell_6t_5 inst_cell_221_87 (.BL(BL87),.BLN(BLN87),.WL(WL221));
sram_cell_6t_5 inst_cell_221_88 (.BL(BL88),.BLN(BLN88),.WL(WL221));
sram_cell_6t_5 inst_cell_221_89 (.BL(BL89),.BLN(BLN89),.WL(WL221));
sram_cell_6t_5 inst_cell_221_90 (.BL(BL90),.BLN(BLN90),.WL(WL221));
sram_cell_6t_5 inst_cell_221_91 (.BL(BL91),.BLN(BLN91),.WL(WL221));
sram_cell_6t_5 inst_cell_221_92 (.BL(BL92),.BLN(BLN92),.WL(WL221));
sram_cell_6t_5 inst_cell_221_93 (.BL(BL93),.BLN(BLN93),.WL(WL221));
sram_cell_6t_5 inst_cell_221_94 (.BL(BL94),.BLN(BLN94),.WL(WL221));
sram_cell_6t_5 inst_cell_221_95 (.BL(BL95),.BLN(BLN95),.WL(WL221));
sram_cell_6t_5 inst_cell_221_96 (.BL(BL96),.BLN(BLN96),.WL(WL221));
sram_cell_6t_5 inst_cell_221_97 (.BL(BL97),.BLN(BLN97),.WL(WL221));
sram_cell_6t_5 inst_cell_221_98 (.BL(BL98),.BLN(BLN98),.WL(WL221));
sram_cell_6t_5 inst_cell_221_99 (.BL(BL99),.BLN(BLN99),.WL(WL221));
sram_cell_6t_5 inst_cell_221_100 (.BL(BL100),.BLN(BLN100),.WL(WL221));
sram_cell_6t_5 inst_cell_221_101 (.BL(BL101),.BLN(BLN101),.WL(WL221));
sram_cell_6t_5 inst_cell_221_102 (.BL(BL102),.BLN(BLN102),.WL(WL221));
sram_cell_6t_5 inst_cell_221_103 (.BL(BL103),.BLN(BLN103),.WL(WL221));
sram_cell_6t_5 inst_cell_221_104 (.BL(BL104),.BLN(BLN104),.WL(WL221));
sram_cell_6t_5 inst_cell_221_105 (.BL(BL105),.BLN(BLN105),.WL(WL221));
sram_cell_6t_5 inst_cell_221_106 (.BL(BL106),.BLN(BLN106),.WL(WL221));
sram_cell_6t_5 inst_cell_221_107 (.BL(BL107),.BLN(BLN107),.WL(WL221));
sram_cell_6t_5 inst_cell_221_108 (.BL(BL108),.BLN(BLN108),.WL(WL221));
sram_cell_6t_5 inst_cell_221_109 (.BL(BL109),.BLN(BLN109),.WL(WL221));
sram_cell_6t_5 inst_cell_221_110 (.BL(BL110),.BLN(BLN110),.WL(WL221));
sram_cell_6t_5 inst_cell_221_111 (.BL(BL111),.BLN(BLN111),.WL(WL221));
sram_cell_6t_5 inst_cell_221_112 (.BL(BL112),.BLN(BLN112),.WL(WL221));
sram_cell_6t_5 inst_cell_221_113 (.BL(BL113),.BLN(BLN113),.WL(WL221));
sram_cell_6t_5 inst_cell_221_114 (.BL(BL114),.BLN(BLN114),.WL(WL221));
sram_cell_6t_5 inst_cell_221_115 (.BL(BL115),.BLN(BLN115),.WL(WL221));
sram_cell_6t_5 inst_cell_221_116 (.BL(BL116),.BLN(BLN116),.WL(WL221));
sram_cell_6t_5 inst_cell_221_117 (.BL(BL117),.BLN(BLN117),.WL(WL221));
sram_cell_6t_5 inst_cell_221_118 (.BL(BL118),.BLN(BLN118),.WL(WL221));
sram_cell_6t_5 inst_cell_221_119 (.BL(BL119),.BLN(BLN119),.WL(WL221));
sram_cell_6t_5 inst_cell_221_120 (.BL(BL120),.BLN(BLN120),.WL(WL221));
sram_cell_6t_5 inst_cell_221_121 (.BL(BL121),.BLN(BLN121),.WL(WL221));
sram_cell_6t_5 inst_cell_221_122 (.BL(BL122),.BLN(BLN122),.WL(WL221));
sram_cell_6t_5 inst_cell_221_123 (.BL(BL123),.BLN(BLN123),.WL(WL221));
sram_cell_6t_5 inst_cell_221_124 (.BL(BL124),.BLN(BLN124),.WL(WL221));
sram_cell_6t_5 inst_cell_221_125 (.BL(BL125),.BLN(BLN125),.WL(WL221));
sram_cell_6t_5 inst_cell_221_126 (.BL(BL126),.BLN(BLN126),.WL(WL221));
sram_cell_6t_5 inst_cell_221_127 (.BL(BL127),.BLN(BLN127),.WL(WL221));
sram_cell_6t_5 inst_cell_222_0 (.BL(BL0),.BLN(BLN0),.WL(WL222));
sram_cell_6t_5 inst_cell_222_1 (.BL(BL1),.BLN(BLN1),.WL(WL222));
sram_cell_6t_5 inst_cell_222_2 (.BL(BL2),.BLN(BLN2),.WL(WL222));
sram_cell_6t_5 inst_cell_222_3 (.BL(BL3),.BLN(BLN3),.WL(WL222));
sram_cell_6t_5 inst_cell_222_4 (.BL(BL4),.BLN(BLN4),.WL(WL222));
sram_cell_6t_5 inst_cell_222_5 (.BL(BL5),.BLN(BLN5),.WL(WL222));
sram_cell_6t_5 inst_cell_222_6 (.BL(BL6),.BLN(BLN6),.WL(WL222));
sram_cell_6t_5 inst_cell_222_7 (.BL(BL7),.BLN(BLN7),.WL(WL222));
sram_cell_6t_5 inst_cell_222_8 (.BL(BL8),.BLN(BLN8),.WL(WL222));
sram_cell_6t_5 inst_cell_222_9 (.BL(BL9),.BLN(BLN9),.WL(WL222));
sram_cell_6t_5 inst_cell_222_10 (.BL(BL10),.BLN(BLN10),.WL(WL222));
sram_cell_6t_5 inst_cell_222_11 (.BL(BL11),.BLN(BLN11),.WL(WL222));
sram_cell_6t_5 inst_cell_222_12 (.BL(BL12),.BLN(BLN12),.WL(WL222));
sram_cell_6t_5 inst_cell_222_13 (.BL(BL13),.BLN(BLN13),.WL(WL222));
sram_cell_6t_5 inst_cell_222_14 (.BL(BL14),.BLN(BLN14),.WL(WL222));
sram_cell_6t_5 inst_cell_222_15 (.BL(BL15),.BLN(BLN15),.WL(WL222));
sram_cell_6t_5 inst_cell_222_16 (.BL(BL16),.BLN(BLN16),.WL(WL222));
sram_cell_6t_5 inst_cell_222_17 (.BL(BL17),.BLN(BLN17),.WL(WL222));
sram_cell_6t_5 inst_cell_222_18 (.BL(BL18),.BLN(BLN18),.WL(WL222));
sram_cell_6t_5 inst_cell_222_19 (.BL(BL19),.BLN(BLN19),.WL(WL222));
sram_cell_6t_5 inst_cell_222_20 (.BL(BL20),.BLN(BLN20),.WL(WL222));
sram_cell_6t_5 inst_cell_222_21 (.BL(BL21),.BLN(BLN21),.WL(WL222));
sram_cell_6t_5 inst_cell_222_22 (.BL(BL22),.BLN(BLN22),.WL(WL222));
sram_cell_6t_5 inst_cell_222_23 (.BL(BL23),.BLN(BLN23),.WL(WL222));
sram_cell_6t_5 inst_cell_222_24 (.BL(BL24),.BLN(BLN24),.WL(WL222));
sram_cell_6t_5 inst_cell_222_25 (.BL(BL25),.BLN(BLN25),.WL(WL222));
sram_cell_6t_5 inst_cell_222_26 (.BL(BL26),.BLN(BLN26),.WL(WL222));
sram_cell_6t_5 inst_cell_222_27 (.BL(BL27),.BLN(BLN27),.WL(WL222));
sram_cell_6t_5 inst_cell_222_28 (.BL(BL28),.BLN(BLN28),.WL(WL222));
sram_cell_6t_5 inst_cell_222_29 (.BL(BL29),.BLN(BLN29),.WL(WL222));
sram_cell_6t_5 inst_cell_222_30 (.BL(BL30),.BLN(BLN30),.WL(WL222));
sram_cell_6t_5 inst_cell_222_31 (.BL(BL31),.BLN(BLN31),.WL(WL222));
sram_cell_6t_5 inst_cell_222_32 (.BL(BL32),.BLN(BLN32),.WL(WL222));
sram_cell_6t_5 inst_cell_222_33 (.BL(BL33),.BLN(BLN33),.WL(WL222));
sram_cell_6t_5 inst_cell_222_34 (.BL(BL34),.BLN(BLN34),.WL(WL222));
sram_cell_6t_5 inst_cell_222_35 (.BL(BL35),.BLN(BLN35),.WL(WL222));
sram_cell_6t_5 inst_cell_222_36 (.BL(BL36),.BLN(BLN36),.WL(WL222));
sram_cell_6t_5 inst_cell_222_37 (.BL(BL37),.BLN(BLN37),.WL(WL222));
sram_cell_6t_5 inst_cell_222_38 (.BL(BL38),.BLN(BLN38),.WL(WL222));
sram_cell_6t_5 inst_cell_222_39 (.BL(BL39),.BLN(BLN39),.WL(WL222));
sram_cell_6t_5 inst_cell_222_40 (.BL(BL40),.BLN(BLN40),.WL(WL222));
sram_cell_6t_5 inst_cell_222_41 (.BL(BL41),.BLN(BLN41),.WL(WL222));
sram_cell_6t_5 inst_cell_222_42 (.BL(BL42),.BLN(BLN42),.WL(WL222));
sram_cell_6t_5 inst_cell_222_43 (.BL(BL43),.BLN(BLN43),.WL(WL222));
sram_cell_6t_5 inst_cell_222_44 (.BL(BL44),.BLN(BLN44),.WL(WL222));
sram_cell_6t_5 inst_cell_222_45 (.BL(BL45),.BLN(BLN45),.WL(WL222));
sram_cell_6t_5 inst_cell_222_46 (.BL(BL46),.BLN(BLN46),.WL(WL222));
sram_cell_6t_5 inst_cell_222_47 (.BL(BL47),.BLN(BLN47),.WL(WL222));
sram_cell_6t_5 inst_cell_222_48 (.BL(BL48),.BLN(BLN48),.WL(WL222));
sram_cell_6t_5 inst_cell_222_49 (.BL(BL49),.BLN(BLN49),.WL(WL222));
sram_cell_6t_5 inst_cell_222_50 (.BL(BL50),.BLN(BLN50),.WL(WL222));
sram_cell_6t_5 inst_cell_222_51 (.BL(BL51),.BLN(BLN51),.WL(WL222));
sram_cell_6t_5 inst_cell_222_52 (.BL(BL52),.BLN(BLN52),.WL(WL222));
sram_cell_6t_5 inst_cell_222_53 (.BL(BL53),.BLN(BLN53),.WL(WL222));
sram_cell_6t_5 inst_cell_222_54 (.BL(BL54),.BLN(BLN54),.WL(WL222));
sram_cell_6t_5 inst_cell_222_55 (.BL(BL55),.BLN(BLN55),.WL(WL222));
sram_cell_6t_5 inst_cell_222_56 (.BL(BL56),.BLN(BLN56),.WL(WL222));
sram_cell_6t_5 inst_cell_222_57 (.BL(BL57),.BLN(BLN57),.WL(WL222));
sram_cell_6t_5 inst_cell_222_58 (.BL(BL58),.BLN(BLN58),.WL(WL222));
sram_cell_6t_5 inst_cell_222_59 (.BL(BL59),.BLN(BLN59),.WL(WL222));
sram_cell_6t_5 inst_cell_222_60 (.BL(BL60),.BLN(BLN60),.WL(WL222));
sram_cell_6t_5 inst_cell_222_61 (.BL(BL61),.BLN(BLN61),.WL(WL222));
sram_cell_6t_5 inst_cell_222_62 (.BL(BL62),.BLN(BLN62),.WL(WL222));
sram_cell_6t_5 inst_cell_222_63 (.BL(BL63),.BLN(BLN63),.WL(WL222));
sram_cell_6t_5 inst_cell_222_64 (.BL(BL64),.BLN(BLN64),.WL(WL222));
sram_cell_6t_5 inst_cell_222_65 (.BL(BL65),.BLN(BLN65),.WL(WL222));
sram_cell_6t_5 inst_cell_222_66 (.BL(BL66),.BLN(BLN66),.WL(WL222));
sram_cell_6t_5 inst_cell_222_67 (.BL(BL67),.BLN(BLN67),.WL(WL222));
sram_cell_6t_5 inst_cell_222_68 (.BL(BL68),.BLN(BLN68),.WL(WL222));
sram_cell_6t_5 inst_cell_222_69 (.BL(BL69),.BLN(BLN69),.WL(WL222));
sram_cell_6t_5 inst_cell_222_70 (.BL(BL70),.BLN(BLN70),.WL(WL222));
sram_cell_6t_5 inst_cell_222_71 (.BL(BL71),.BLN(BLN71),.WL(WL222));
sram_cell_6t_5 inst_cell_222_72 (.BL(BL72),.BLN(BLN72),.WL(WL222));
sram_cell_6t_5 inst_cell_222_73 (.BL(BL73),.BLN(BLN73),.WL(WL222));
sram_cell_6t_5 inst_cell_222_74 (.BL(BL74),.BLN(BLN74),.WL(WL222));
sram_cell_6t_5 inst_cell_222_75 (.BL(BL75),.BLN(BLN75),.WL(WL222));
sram_cell_6t_5 inst_cell_222_76 (.BL(BL76),.BLN(BLN76),.WL(WL222));
sram_cell_6t_5 inst_cell_222_77 (.BL(BL77),.BLN(BLN77),.WL(WL222));
sram_cell_6t_5 inst_cell_222_78 (.BL(BL78),.BLN(BLN78),.WL(WL222));
sram_cell_6t_5 inst_cell_222_79 (.BL(BL79),.BLN(BLN79),.WL(WL222));
sram_cell_6t_5 inst_cell_222_80 (.BL(BL80),.BLN(BLN80),.WL(WL222));
sram_cell_6t_5 inst_cell_222_81 (.BL(BL81),.BLN(BLN81),.WL(WL222));
sram_cell_6t_5 inst_cell_222_82 (.BL(BL82),.BLN(BLN82),.WL(WL222));
sram_cell_6t_5 inst_cell_222_83 (.BL(BL83),.BLN(BLN83),.WL(WL222));
sram_cell_6t_5 inst_cell_222_84 (.BL(BL84),.BLN(BLN84),.WL(WL222));
sram_cell_6t_5 inst_cell_222_85 (.BL(BL85),.BLN(BLN85),.WL(WL222));
sram_cell_6t_5 inst_cell_222_86 (.BL(BL86),.BLN(BLN86),.WL(WL222));
sram_cell_6t_5 inst_cell_222_87 (.BL(BL87),.BLN(BLN87),.WL(WL222));
sram_cell_6t_5 inst_cell_222_88 (.BL(BL88),.BLN(BLN88),.WL(WL222));
sram_cell_6t_5 inst_cell_222_89 (.BL(BL89),.BLN(BLN89),.WL(WL222));
sram_cell_6t_5 inst_cell_222_90 (.BL(BL90),.BLN(BLN90),.WL(WL222));
sram_cell_6t_5 inst_cell_222_91 (.BL(BL91),.BLN(BLN91),.WL(WL222));
sram_cell_6t_5 inst_cell_222_92 (.BL(BL92),.BLN(BLN92),.WL(WL222));
sram_cell_6t_5 inst_cell_222_93 (.BL(BL93),.BLN(BLN93),.WL(WL222));
sram_cell_6t_5 inst_cell_222_94 (.BL(BL94),.BLN(BLN94),.WL(WL222));
sram_cell_6t_5 inst_cell_222_95 (.BL(BL95),.BLN(BLN95),.WL(WL222));
sram_cell_6t_5 inst_cell_222_96 (.BL(BL96),.BLN(BLN96),.WL(WL222));
sram_cell_6t_5 inst_cell_222_97 (.BL(BL97),.BLN(BLN97),.WL(WL222));
sram_cell_6t_5 inst_cell_222_98 (.BL(BL98),.BLN(BLN98),.WL(WL222));
sram_cell_6t_5 inst_cell_222_99 (.BL(BL99),.BLN(BLN99),.WL(WL222));
sram_cell_6t_5 inst_cell_222_100 (.BL(BL100),.BLN(BLN100),.WL(WL222));
sram_cell_6t_5 inst_cell_222_101 (.BL(BL101),.BLN(BLN101),.WL(WL222));
sram_cell_6t_5 inst_cell_222_102 (.BL(BL102),.BLN(BLN102),.WL(WL222));
sram_cell_6t_5 inst_cell_222_103 (.BL(BL103),.BLN(BLN103),.WL(WL222));
sram_cell_6t_5 inst_cell_222_104 (.BL(BL104),.BLN(BLN104),.WL(WL222));
sram_cell_6t_5 inst_cell_222_105 (.BL(BL105),.BLN(BLN105),.WL(WL222));
sram_cell_6t_5 inst_cell_222_106 (.BL(BL106),.BLN(BLN106),.WL(WL222));
sram_cell_6t_5 inst_cell_222_107 (.BL(BL107),.BLN(BLN107),.WL(WL222));
sram_cell_6t_5 inst_cell_222_108 (.BL(BL108),.BLN(BLN108),.WL(WL222));
sram_cell_6t_5 inst_cell_222_109 (.BL(BL109),.BLN(BLN109),.WL(WL222));
sram_cell_6t_5 inst_cell_222_110 (.BL(BL110),.BLN(BLN110),.WL(WL222));
sram_cell_6t_5 inst_cell_222_111 (.BL(BL111),.BLN(BLN111),.WL(WL222));
sram_cell_6t_5 inst_cell_222_112 (.BL(BL112),.BLN(BLN112),.WL(WL222));
sram_cell_6t_5 inst_cell_222_113 (.BL(BL113),.BLN(BLN113),.WL(WL222));
sram_cell_6t_5 inst_cell_222_114 (.BL(BL114),.BLN(BLN114),.WL(WL222));
sram_cell_6t_5 inst_cell_222_115 (.BL(BL115),.BLN(BLN115),.WL(WL222));
sram_cell_6t_5 inst_cell_222_116 (.BL(BL116),.BLN(BLN116),.WL(WL222));
sram_cell_6t_5 inst_cell_222_117 (.BL(BL117),.BLN(BLN117),.WL(WL222));
sram_cell_6t_5 inst_cell_222_118 (.BL(BL118),.BLN(BLN118),.WL(WL222));
sram_cell_6t_5 inst_cell_222_119 (.BL(BL119),.BLN(BLN119),.WL(WL222));
sram_cell_6t_5 inst_cell_222_120 (.BL(BL120),.BLN(BLN120),.WL(WL222));
sram_cell_6t_5 inst_cell_222_121 (.BL(BL121),.BLN(BLN121),.WL(WL222));
sram_cell_6t_5 inst_cell_222_122 (.BL(BL122),.BLN(BLN122),.WL(WL222));
sram_cell_6t_5 inst_cell_222_123 (.BL(BL123),.BLN(BLN123),.WL(WL222));
sram_cell_6t_5 inst_cell_222_124 (.BL(BL124),.BLN(BLN124),.WL(WL222));
sram_cell_6t_5 inst_cell_222_125 (.BL(BL125),.BLN(BLN125),.WL(WL222));
sram_cell_6t_5 inst_cell_222_126 (.BL(BL126),.BLN(BLN126),.WL(WL222));
sram_cell_6t_5 inst_cell_222_127 (.BL(BL127),.BLN(BLN127),.WL(WL222));
sram_cell_6t_5 inst_cell_223_0 (.BL(BL0),.BLN(BLN0),.WL(WL223));
sram_cell_6t_5 inst_cell_223_1 (.BL(BL1),.BLN(BLN1),.WL(WL223));
sram_cell_6t_5 inst_cell_223_2 (.BL(BL2),.BLN(BLN2),.WL(WL223));
sram_cell_6t_5 inst_cell_223_3 (.BL(BL3),.BLN(BLN3),.WL(WL223));
sram_cell_6t_5 inst_cell_223_4 (.BL(BL4),.BLN(BLN4),.WL(WL223));
sram_cell_6t_5 inst_cell_223_5 (.BL(BL5),.BLN(BLN5),.WL(WL223));
sram_cell_6t_5 inst_cell_223_6 (.BL(BL6),.BLN(BLN6),.WL(WL223));
sram_cell_6t_5 inst_cell_223_7 (.BL(BL7),.BLN(BLN7),.WL(WL223));
sram_cell_6t_5 inst_cell_223_8 (.BL(BL8),.BLN(BLN8),.WL(WL223));
sram_cell_6t_5 inst_cell_223_9 (.BL(BL9),.BLN(BLN9),.WL(WL223));
sram_cell_6t_5 inst_cell_223_10 (.BL(BL10),.BLN(BLN10),.WL(WL223));
sram_cell_6t_5 inst_cell_223_11 (.BL(BL11),.BLN(BLN11),.WL(WL223));
sram_cell_6t_5 inst_cell_223_12 (.BL(BL12),.BLN(BLN12),.WL(WL223));
sram_cell_6t_5 inst_cell_223_13 (.BL(BL13),.BLN(BLN13),.WL(WL223));
sram_cell_6t_5 inst_cell_223_14 (.BL(BL14),.BLN(BLN14),.WL(WL223));
sram_cell_6t_5 inst_cell_223_15 (.BL(BL15),.BLN(BLN15),.WL(WL223));
sram_cell_6t_5 inst_cell_223_16 (.BL(BL16),.BLN(BLN16),.WL(WL223));
sram_cell_6t_5 inst_cell_223_17 (.BL(BL17),.BLN(BLN17),.WL(WL223));
sram_cell_6t_5 inst_cell_223_18 (.BL(BL18),.BLN(BLN18),.WL(WL223));
sram_cell_6t_5 inst_cell_223_19 (.BL(BL19),.BLN(BLN19),.WL(WL223));
sram_cell_6t_5 inst_cell_223_20 (.BL(BL20),.BLN(BLN20),.WL(WL223));
sram_cell_6t_5 inst_cell_223_21 (.BL(BL21),.BLN(BLN21),.WL(WL223));
sram_cell_6t_5 inst_cell_223_22 (.BL(BL22),.BLN(BLN22),.WL(WL223));
sram_cell_6t_5 inst_cell_223_23 (.BL(BL23),.BLN(BLN23),.WL(WL223));
sram_cell_6t_5 inst_cell_223_24 (.BL(BL24),.BLN(BLN24),.WL(WL223));
sram_cell_6t_5 inst_cell_223_25 (.BL(BL25),.BLN(BLN25),.WL(WL223));
sram_cell_6t_5 inst_cell_223_26 (.BL(BL26),.BLN(BLN26),.WL(WL223));
sram_cell_6t_5 inst_cell_223_27 (.BL(BL27),.BLN(BLN27),.WL(WL223));
sram_cell_6t_5 inst_cell_223_28 (.BL(BL28),.BLN(BLN28),.WL(WL223));
sram_cell_6t_5 inst_cell_223_29 (.BL(BL29),.BLN(BLN29),.WL(WL223));
sram_cell_6t_5 inst_cell_223_30 (.BL(BL30),.BLN(BLN30),.WL(WL223));
sram_cell_6t_5 inst_cell_223_31 (.BL(BL31),.BLN(BLN31),.WL(WL223));
sram_cell_6t_5 inst_cell_223_32 (.BL(BL32),.BLN(BLN32),.WL(WL223));
sram_cell_6t_5 inst_cell_223_33 (.BL(BL33),.BLN(BLN33),.WL(WL223));
sram_cell_6t_5 inst_cell_223_34 (.BL(BL34),.BLN(BLN34),.WL(WL223));
sram_cell_6t_5 inst_cell_223_35 (.BL(BL35),.BLN(BLN35),.WL(WL223));
sram_cell_6t_5 inst_cell_223_36 (.BL(BL36),.BLN(BLN36),.WL(WL223));
sram_cell_6t_5 inst_cell_223_37 (.BL(BL37),.BLN(BLN37),.WL(WL223));
sram_cell_6t_5 inst_cell_223_38 (.BL(BL38),.BLN(BLN38),.WL(WL223));
sram_cell_6t_5 inst_cell_223_39 (.BL(BL39),.BLN(BLN39),.WL(WL223));
sram_cell_6t_5 inst_cell_223_40 (.BL(BL40),.BLN(BLN40),.WL(WL223));
sram_cell_6t_5 inst_cell_223_41 (.BL(BL41),.BLN(BLN41),.WL(WL223));
sram_cell_6t_5 inst_cell_223_42 (.BL(BL42),.BLN(BLN42),.WL(WL223));
sram_cell_6t_5 inst_cell_223_43 (.BL(BL43),.BLN(BLN43),.WL(WL223));
sram_cell_6t_5 inst_cell_223_44 (.BL(BL44),.BLN(BLN44),.WL(WL223));
sram_cell_6t_5 inst_cell_223_45 (.BL(BL45),.BLN(BLN45),.WL(WL223));
sram_cell_6t_5 inst_cell_223_46 (.BL(BL46),.BLN(BLN46),.WL(WL223));
sram_cell_6t_5 inst_cell_223_47 (.BL(BL47),.BLN(BLN47),.WL(WL223));
sram_cell_6t_5 inst_cell_223_48 (.BL(BL48),.BLN(BLN48),.WL(WL223));
sram_cell_6t_5 inst_cell_223_49 (.BL(BL49),.BLN(BLN49),.WL(WL223));
sram_cell_6t_5 inst_cell_223_50 (.BL(BL50),.BLN(BLN50),.WL(WL223));
sram_cell_6t_5 inst_cell_223_51 (.BL(BL51),.BLN(BLN51),.WL(WL223));
sram_cell_6t_5 inst_cell_223_52 (.BL(BL52),.BLN(BLN52),.WL(WL223));
sram_cell_6t_5 inst_cell_223_53 (.BL(BL53),.BLN(BLN53),.WL(WL223));
sram_cell_6t_5 inst_cell_223_54 (.BL(BL54),.BLN(BLN54),.WL(WL223));
sram_cell_6t_5 inst_cell_223_55 (.BL(BL55),.BLN(BLN55),.WL(WL223));
sram_cell_6t_5 inst_cell_223_56 (.BL(BL56),.BLN(BLN56),.WL(WL223));
sram_cell_6t_5 inst_cell_223_57 (.BL(BL57),.BLN(BLN57),.WL(WL223));
sram_cell_6t_5 inst_cell_223_58 (.BL(BL58),.BLN(BLN58),.WL(WL223));
sram_cell_6t_5 inst_cell_223_59 (.BL(BL59),.BLN(BLN59),.WL(WL223));
sram_cell_6t_5 inst_cell_223_60 (.BL(BL60),.BLN(BLN60),.WL(WL223));
sram_cell_6t_5 inst_cell_223_61 (.BL(BL61),.BLN(BLN61),.WL(WL223));
sram_cell_6t_5 inst_cell_223_62 (.BL(BL62),.BLN(BLN62),.WL(WL223));
sram_cell_6t_5 inst_cell_223_63 (.BL(BL63),.BLN(BLN63),.WL(WL223));
sram_cell_6t_5 inst_cell_223_64 (.BL(BL64),.BLN(BLN64),.WL(WL223));
sram_cell_6t_5 inst_cell_223_65 (.BL(BL65),.BLN(BLN65),.WL(WL223));
sram_cell_6t_5 inst_cell_223_66 (.BL(BL66),.BLN(BLN66),.WL(WL223));
sram_cell_6t_5 inst_cell_223_67 (.BL(BL67),.BLN(BLN67),.WL(WL223));
sram_cell_6t_5 inst_cell_223_68 (.BL(BL68),.BLN(BLN68),.WL(WL223));
sram_cell_6t_5 inst_cell_223_69 (.BL(BL69),.BLN(BLN69),.WL(WL223));
sram_cell_6t_5 inst_cell_223_70 (.BL(BL70),.BLN(BLN70),.WL(WL223));
sram_cell_6t_5 inst_cell_223_71 (.BL(BL71),.BLN(BLN71),.WL(WL223));
sram_cell_6t_5 inst_cell_223_72 (.BL(BL72),.BLN(BLN72),.WL(WL223));
sram_cell_6t_5 inst_cell_223_73 (.BL(BL73),.BLN(BLN73),.WL(WL223));
sram_cell_6t_5 inst_cell_223_74 (.BL(BL74),.BLN(BLN74),.WL(WL223));
sram_cell_6t_5 inst_cell_223_75 (.BL(BL75),.BLN(BLN75),.WL(WL223));
sram_cell_6t_5 inst_cell_223_76 (.BL(BL76),.BLN(BLN76),.WL(WL223));
sram_cell_6t_5 inst_cell_223_77 (.BL(BL77),.BLN(BLN77),.WL(WL223));
sram_cell_6t_5 inst_cell_223_78 (.BL(BL78),.BLN(BLN78),.WL(WL223));
sram_cell_6t_5 inst_cell_223_79 (.BL(BL79),.BLN(BLN79),.WL(WL223));
sram_cell_6t_5 inst_cell_223_80 (.BL(BL80),.BLN(BLN80),.WL(WL223));
sram_cell_6t_5 inst_cell_223_81 (.BL(BL81),.BLN(BLN81),.WL(WL223));
sram_cell_6t_5 inst_cell_223_82 (.BL(BL82),.BLN(BLN82),.WL(WL223));
sram_cell_6t_5 inst_cell_223_83 (.BL(BL83),.BLN(BLN83),.WL(WL223));
sram_cell_6t_5 inst_cell_223_84 (.BL(BL84),.BLN(BLN84),.WL(WL223));
sram_cell_6t_5 inst_cell_223_85 (.BL(BL85),.BLN(BLN85),.WL(WL223));
sram_cell_6t_5 inst_cell_223_86 (.BL(BL86),.BLN(BLN86),.WL(WL223));
sram_cell_6t_5 inst_cell_223_87 (.BL(BL87),.BLN(BLN87),.WL(WL223));
sram_cell_6t_5 inst_cell_223_88 (.BL(BL88),.BLN(BLN88),.WL(WL223));
sram_cell_6t_5 inst_cell_223_89 (.BL(BL89),.BLN(BLN89),.WL(WL223));
sram_cell_6t_5 inst_cell_223_90 (.BL(BL90),.BLN(BLN90),.WL(WL223));
sram_cell_6t_5 inst_cell_223_91 (.BL(BL91),.BLN(BLN91),.WL(WL223));
sram_cell_6t_5 inst_cell_223_92 (.BL(BL92),.BLN(BLN92),.WL(WL223));
sram_cell_6t_5 inst_cell_223_93 (.BL(BL93),.BLN(BLN93),.WL(WL223));
sram_cell_6t_5 inst_cell_223_94 (.BL(BL94),.BLN(BLN94),.WL(WL223));
sram_cell_6t_5 inst_cell_223_95 (.BL(BL95),.BLN(BLN95),.WL(WL223));
sram_cell_6t_5 inst_cell_223_96 (.BL(BL96),.BLN(BLN96),.WL(WL223));
sram_cell_6t_5 inst_cell_223_97 (.BL(BL97),.BLN(BLN97),.WL(WL223));
sram_cell_6t_5 inst_cell_223_98 (.BL(BL98),.BLN(BLN98),.WL(WL223));
sram_cell_6t_5 inst_cell_223_99 (.BL(BL99),.BLN(BLN99),.WL(WL223));
sram_cell_6t_5 inst_cell_223_100 (.BL(BL100),.BLN(BLN100),.WL(WL223));
sram_cell_6t_5 inst_cell_223_101 (.BL(BL101),.BLN(BLN101),.WL(WL223));
sram_cell_6t_5 inst_cell_223_102 (.BL(BL102),.BLN(BLN102),.WL(WL223));
sram_cell_6t_5 inst_cell_223_103 (.BL(BL103),.BLN(BLN103),.WL(WL223));
sram_cell_6t_5 inst_cell_223_104 (.BL(BL104),.BLN(BLN104),.WL(WL223));
sram_cell_6t_5 inst_cell_223_105 (.BL(BL105),.BLN(BLN105),.WL(WL223));
sram_cell_6t_5 inst_cell_223_106 (.BL(BL106),.BLN(BLN106),.WL(WL223));
sram_cell_6t_5 inst_cell_223_107 (.BL(BL107),.BLN(BLN107),.WL(WL223));
sram_cell_6t_5 inst_cell_223_108 (.BL(BL108),.BLN(BLN108),.WL(WL223));
sram_cell_6t_5 inst_cell_223_109 (.BL(BL109),.BLN(BLN109),.WL(WL223));
sram_cell_6t_5 inst_cell_223_110 (.BL(BL110),.BLN(BLN110),.WL(WL223));
sram_cell_6t_5 inst_cell_223_111 (.BL(BL111),.BLN(BLN111),.WL(WL223));
sram_cell_6t_5 inst_cell_223_112 (.BL(BL112),.BLN(BLN112),.WL(WL223));
sram_cell_6t_5 inst_cell_223_113 (.BL(BL113),.BLN(BLN113),.WL(WL223));
sram_cell_6t_5 inst_cell_223_114 (.BL(BL114),.BLN(BLN114),.WL(WL223));
sram_cell_6t_5 inst_cell_223_115 (.BL(BL115),.BLN(BLN115),.WL(WL223));
sram_cell_6t_5 inst_cell_223_116 (.BL(BL116),.BLN(BLN116),.WL(WL223));
sram_cell_6t_5 inst_cell_223_117 (.BL(BL117),.BLN(BLN117),.WL(WL223));
sram_cell_6t_5 inst_cell_223_118 (.BL(BL118),.BLN(BLN118),.WL(WL223));
sram_cell_6t_5 inst_cell_223_119 (.BL(BL119),.BLN(BLN119),.WL(WL223));
sram_cell_6t_5 inst_cell_223_120 (.BL(BL120),.BLN(BLN120),.WL(WL223));
sram_cell_6t_5 inst_cell_223_121 (.BL(BL121),.BLN(BLN121),.WL(WL223));
sram_cell_6t_5 inst_cell_223_122 (.BL(BL122),.BLN(BLN122),.WL(WL223));
sram_cell_6t_5 inst_cell_223_123 (.BL(BL123),.BLN(BLN123),.WL(WL223));
sram_cell_6t_5 inst_cell_223_124 (.BL(BL124),.BLN(BLN124),.WL(WL223));
sram_cell_6t_5 inst_cell_223_125 (.BL(BL125),.BLN(BLN125),.WL(WL223));
sram_cell_6t_5 inst_cell_223_126 (.BL(BL126),.BLN(BLN126),.WL(WL223));
sram_cell_6t_5 inst_cell_223_127 (.BL(BL127),.BLN(BLN127),.WL(WL223));
sram_cell_6t_5 inst_cell_224_0 (.BL(BL0),.BLN(BLN0),.WL(WL224));
sram_cell_6t_5 inst_cell_224_1 (.BL(BL1),.BLN(BLN1),.WL(WL224));
sram_cell_6t_5 inst_cell_224_2 (.BL(BL2),.BLN(BLN2),.WL(WL224));
sram_cell_6t_5 inst_cell_224_3 (.BL(BL3),.BLN(BLN3),.WL(WL224));
sram_cell_6t_5 inst_cell_224_4 (.BL(BL4),.BLN(BLN4),.WL(WL224));
sram_cell_6t_5 inst_cell_224_5 (.BL(BL5),.BLN(BLN5),.WL(WL224));
sram_cell_6t_5 inst_cell_224_6 (.BL(BL6),.BLN(BLN6),.WL(WL224));
sram_cell_6t_5 inst_cell_224_7 (.BL(BL7),.BLN(BLN7),.WL(WL224));
sram_cell_6t_5 inst_cell_224_8 (.BL(BL8),.BLN(BLN8),.WL(WL224));
sram_cell_6t_5 inst_cell_224_9 (.BL(BL9),.BLN(BLN9),.WL(WL224));
sram_cell_6t_5 inst_cell_224_10 (.BL(BL10),.BLN(BLN10),.WL(WL224));
sram_cell_6t_5 inst_cell_224_11 (.BL(BL11),.BLN(BLN11),.WL(WL224));
sram_cell_6t_5 inst_cell_224_12 (.BL(BL12),.BLN(BLN12),.WL(WL224));
sram_cell_6t_5 inst_cell_224_13 (.BL(BL13),.BLN(BLN13),.WL(WL224));
sram_cell_6t_5 inst_cell_224_14 (.BL(BL14),.BLN(BLN14),.WL(WL224));
sram_cell_6t_5 inst_cell_224_15 (.BL(BL15),.BLN(BLN15),.WL(WL224));
sram_cell_6t_5 inst_cell_224_16 (.BL(BL16),.BLN(BLN16),.WL(WL224));
sram_cell_6t_5 inst_cell_224_17 (.BL(BL17),.BLN(BLN17),.WL(WL224));
sram_cell_6t_5 inst_cell_224_18 (.BL(BL18),.BLN(BLN18),.WL(WL224));
sram_cell_6t_5 inst_cell_224_19 (.BL(BL19),.BLN(BLN19),.WL(WL224));
sram_cell_6t_5 inst_cell_224_20 (.BL(BL20),.BLN(BLN20),.WL(WL224));
sram_cell_6t_5 inst_cell_224_21 (.BL(BL21),.BLN(BLN21),.WL(WL224));
sram_cell_6t_5 inst_cell_224_22 (.BL(BL22),.BLN(BLN22),.WL(WL224));
sram_cell_6t_5 inst_cell_224_23 (.BL(BL23),.BLN(BLN23),.WL(WL224));
sram_cell_6t_5 inst_cell_224_24 (.BL(BL24),.BLN(BLN24),.WL(WL224));
sram_cell_6t_5 inst_cell_224_25 (.BL(BL25),.BLN(BLN25),.WL(WL224));
sram_cell_6t_5 inst_cell_224_26 (.BL(BL26),.BLN(BLN26),.WL(WL224));
sram_cell_6t_5 inst_cell_224_27 (.BL(BL27),.BLN(BLN27),.WL(WL224));
sram_cell_6t_5 inst_cell_224_28 (.BL(BL28),.BLN(BLN28),.WL(WL224));
sram_cell_6t_5 inst_cell_224_29 (.BL(BL29),.BLN(BLN29),.WL(WL224));
sram_cell_6t_5 inst_cell_224_30 (.BL(BL30),.BLN(BLN30),.WL(WL224));
sram_cell_6t_5 inst_cell_224_31 (.BL(BL31),.BLN(BLN31),.WL(WL224));
sram_cell_6t_5 inst_cell_224_32 (.BL(BL32),.BLN(BLN32),.WL(WL224));
sram_cell_6t_5 inst_cell_224_33 (.BL(BL33),.BLN(BLN33),.WL(WL224));
sram_cell_6t_5 inst_cell_224_34 (.BL(BL34),.BLN(BLN34),.WL(WL224));
sram_cell_6t_5 inst_cell_224_35 (.BL(BL35),.BLN(BLN35),.WL(WL224));
sram_cell_6t_5 inst_cell_224_36 (.BL(BL36),.BLN(BLN36),.WL(WL224));
sram_cell_6t_5 inst_cell_224_37 (.BL(BL37),.BLN(BLN37),.WL(WL224));
sram_cell_6t_5 inst_cell_224_38 (.BL(BL38),.BLN(BLN38),.WL(WL224));
sram_cell_6t_5 inst_cell_224_39 (.BL(BL39),.BLN(BLN39),.WL(WL224));
sram_cell_6t_5 inst_cell_224_40 (.BL(BL40),.BLN(BLN40),.WL(WL224));
sram_cell_6t_5 inst_cell_224_41 (.BL(BL41),.BLN(BLN41),.WL(WL224));
sram_cell_6t_5 inst_cell_224_42 (.BL(BL42),.BLN(BLN42),.WL(WL224));
sram_cell_6t_5 inst_cell_224_43 (.BL(BL43),.BLN(BLN43),.WL(WL224));
sram_cell_6t_5 inst_cell_224_44 (.BL(BL44),.BLN(BLN44),.WL(WL224));
sram_cell_6t_5 inst_cell_224_45 (.BL(BL45),.BLN(BLN45),.WL(WL224));
sram_cell_6t_5 inst_cell_224_46 (.BL(BL46),.BLN(BLN46),.WL(WL224));
sram_cell_6t_5 inst_cell_224_47 (.BL(BL47),.BLN(BLN47),.WL(WL224));
sram_cell_6t_5 inst_cell_224_48 (.BL(BL48),.BLN(BLN48),.WL(WL224));
sram_cell_6t_5 inst_cell_224_49 (.BL(BL49),.BLN(BLN49),.WL(WL224));
sram_cell_6t_5 inst_cell_224_50 (.BL(BL50),.BLN(BLN50),.WL(WL224));
sram_cell_6t_5 inst_cell_224_51 (.BL(BL51),.BLN(BLN51),.WL(WL224));
sram_cell_6t_5 inst_cell_224_52 (.BL(BL52),.BLN(BLN52),.WL(WL224));
sram_cell_6t_5 inst_cell_224_53 (.BL(BL53),.BLN(BLN53),.WL(WL224));
sram_cell_6t_5 inst_cell_224_54 (.BL(BL54),.BLN(BLN54),.WL(WL224));
sram_cell_6t_5 inst_cell_224_55 (.BL(BL55),.BLN(BLN55),.WL(WL224));
sram_cell_6t_5 inst_cell_224_56 (.BL(BL56),.BLN(BLN56),.WL(WL224));
sram_cell_6t_5 inst_cell_224_57 (.BL(BL57),.BLN(BLN57),.WL(WL224));
sram_cell_6t_5 inst_cell_224_58 (.BL(BL58),.BLN(BLN58),.WL(WL224));
sram_cell_6t_5 inst_cell_224_59 (.BL(BL59),.BLN(BLN59),.WL(WL224));
sram_cell_6t_5 inst_cell_224_60 (.BL(BL60),.BLN(BLN60),.WL(WL224));
sram_cell_6t_5 inst_cell_224_61 (.BL(BL61),.BLN(BLN61),.WL(WL224));
sram_cell_6t_5 inst_cell_224_62 (.BL(BL62),.BLN(BLN62),.WL(WL224));
sram_cell_6t_5 inst_cell_224_63 (.BL(BL63),.BLN(BLN63),.WL(WL224));
sram_cell_6t_5 inst_cell_224_64 (.BL(BL64),.BLN(BLN64),.WL(WL224));
sram_cell_6t_5 inst_cell_224_65 (.BL(BL65),.BLN(BLN65),.WL(WL224));
sram_cell_6t_5 inst_cell_224_66 (.BL(BL66),.BLN(BLN66),.WL(WL224));
sram_cell_6t_5 inst_cell_224_67 (.BL(BL67),.BLN(BLN67),.WL(WL224));
sram_cell_6t_5 inst_cell_224_68 (.BL(BL68),.BLN(BLN68),.WL(WL224));
sram_cell_6t_5 inst_cell_224_69 (.BL(BL69),.BLN(BLN69),.WL(WL224));
sram_cell_6t_5 inst_cell_224_70 (.BL(BL70),.BLN(BLN70),.WL(WL224));
sram_cell_6t_5 inst_cell_224_71 (.BL(BL71),.BLN(BLN71),.WL(WL224));
sram_cell_6t_5 inst_cell_224_72 (.BL(BL72),.BLN(BLN72),.WL(WL224));
sram_cell_6t_5 inst_cell_224_73 (.BL(BL73),.BLN(BLN73),.WL(WL224));
sram_cell_6t_5 inst_cell_224_74 (.BL(BL74),.BLN(BLN74),.WL(WL224));
sram_cell_6t_5 inst_cell_224_75 (.BL(BL75),.BLN(BLN75),.WL(WL224));
sram_cell_6t_5 inst_cell_224_76 (.BL(BL76),.BLN(BLN76),.WL(WL224));
sram_cell_6t_5 inst_cell_224_77 (.BL(BL77),.BLN(BLN77),.WL(WL224));
sram_cell_6t_5 inst_cell_224_78 (.BL(BL78),.BLN(BLN78),.WL(WL224));
sram_cell_6t_5 inst_cell_224_79 (.BL(BL79),.BLN(BLN79),.WL(WL224));
sram_cell_6t_5 inst_cell_224_80 (.BL(BL80),.BLN(BLN80),.WL(WL224));
sram_cell_6t_5 inst_cell_224_81 (.BL(BL81),.BLN(BLN81),.WL(WL224));
sram_cell_6t_5 inst_cell_224_82 (.BL(BL82),.BLN(BLN82),.WL(WL224));
sram_cell_6t_5 inst_cell_224_83 (.BL(BL83),.BLN(BLN83),.WL(WL224));
sram_cell_6t_5 inst_cell_224_84 (.BL(BL84),.BLN(BLN84),.WL(WL224));
sram_cell_6t_5 inst_cell_224_85 (.BL(BL85),.BLN(BLN85),.WL(WL224));
sram_cell_6t_5 inst_cell_224_86 (.BL(BL86),.BLN(BLN86),.WL(WL224));
sram_cell_6t_5 inst_cell_224_87 (.BL(BL87),.BLN(BLN87),.WL(WL224));
sram_cell_6t_5 inst_cell_224_88 (.BL(BL88),.BLN(BLN88),.WL(WL224));
sram_cell_6t_5 inst_cell_224_89 (.BL(BL89),.BLN(BLN89),.WL(WL224));
sram_cell_6t_5 inst_cell_224_90 (.BL(BL90),.BLN(BLN90),.WL(WL224));
sram_cell_6t_5 inst_cell_224_91 (.BL(BL91),.BLN(BLN91),.WL(WL224));
sram_cell_6t_5 inst_cell_224_92 (.BL(BL92),.BLN(BLN92),.WL(WL224));
sram_cell_6t_5 inst_cell_224_93 (.BL(BL93),.BLN(BLN93),.WL(WL224));
sram_cell_6t_5 inst_cell_224_94 (.BL(BL94),.BLN(BLN94),.WL(WL224));
sram_cell_6t_5 inst_cell_224_95 (.BL(BL95),.BLN(BLN95),.WL(WL224));
sram_cell_6t_5 inst_cell_224_96 (.BL(BL96),.BLN(BLN96),.WL(WL224));
sram_cell_6t_5 inst_cell_224_97 (.BL(BL97),.BLN(BLN97),.WL(WL224));
sram_cell_6t_5 inst_cell_224_98 (.BL(BL98),.BLN(BLN98),.WL(WL224));
sram_cell_6t_5 inst_cell_224_99 (.BL(BL99),.BLN(BLN99),.WL(WL224));
sram_cell_6t_5 inst_cell_224_100 (.BL(BL100),.BLN(BLN100),.WL(WL224));
sram_cell_6t_5 inst_cell_224_101 (.BL(BL101),.BLN(BLN101),.WL(WL224));
sram_cell_6t_5 inst_cell_224_102 (.BL(BL102),.BLN(BLN102),.WL(WL224));
sram_cell_6t_5 inst_cell_224_103 (.BL(BL103),.BLN(BLN103),.WL(WL224));
sram_cell_6t_5 inst_cell_224_104 (.BL(BL104),.BLN(BLN104),.WL(WL224));
sram_cell_6t_5 inst_cell_224_105 (.BL(BL105),.BLN(BLN105),.WL(WL224));
sram_cell_6t_5 inst_cell_224_106 (.BL(BL106),.BLN(BLN106),.WL(WL224));
sram_cell_6t_5 inst_cell_224_107 (.BL(BL107),.BLN(BLN107),.WL(WL224));
sram_cell_6t_5 inst_cell_224_108 (.BL(BL108),.BLN(BLN108),.WL(WL224));
sram_cell_6t_5 inst_cell_224_109 (.BL(BL109),.BLN(BLN109),.WL(WL224));
sram_cell_6t_5 inst_cell_224_110 (.BL(BL110),.BLN(BLN110),.WL(WL224));
sram_cell_6t_5 inst_cell_224_111 (.BL(BL111),.BLN(BLN111),.WL(WL224));
sram_cell_6t_5 inst_cell_224_112 (.BL(BL112),.BLN(BLN112),.WL(WL224));
sram_cell_6t_5 inst_cell_224_113 (.BL(BL113),.BLN(BLN113),.WL(WL224));
sram_cell_6t_5 inst_cell_224_114 (.BL(BL114),.BLN(BLN114),.WL(WL224));
sram_cell_6t_5 inst_cell_224_115 (.BL(BL115),.BLN(BLN115),.WL(WL224));
sram_cell_6t_5 inst_cell_224_116 (.BL(BL116),.BLN(BLN116),.WL(WL224));
sram_cell_6t_5 inst_cell_224_117 (.BL(BL117),.BLN(BLN117),.WL(WL224));
sram_cell_6t_5 inst_cell_224_118 (.BL(BL118),.BLN(BLN118),.WL(WL224));
sram_cell_6t_5 inst_cell_224_119 (.BL(BL119),.BLN(BLN119),.WL(WL224));
sram_cell_6t_5 inst_cell_224_120 (.BL(BL120),.BLN(BLN120),.WL(WL224));
sram_cell_6t_5 inst_cell_224_121 (.BL(BL121),.BLN(BLN121),.WL(WL224));
sram_cell_6t_5 inst_cell_224_122 (.BL(BL122),.BLN(BLN122),.WL(WL224));
sram_cell_6t_5 inst_cell_224_123 (.BL(BL123),.BLN(BLN123),.WL(WL224));
sram_cell_6t_5 inst_cell_224_124 (.BL(BL124),.BLN(BLN124),.WL(WL224));
sram_cell_6t_5 inst_cell_224_125 (.BL(BL125),.BLN(BLN125),.WL(WL224));
sram_cell_6t_5 inst_cell_224_126 (.BL(BL126),.BLN(BLN126),.WL(WL224));
sram_cell_6t_5 inst_cell_224_127 (.BL(BL127),.BLN(BLN127),.WL(WL224));
sram_cell_6t_5 inst_cell_225_0 (.BL(BL0),.BLN(BLN0),.WL(WL225));
sram_cell_6t_5 inst_cell_225_1 (.BL(BL1),.BLN(BLN1),.WL(WL225));
sram_cell_6t_5 inst_cell_225_2 (.BL(BL2),.BLN(BLN2),.WL(WL225));
sram_cell_6t_5 inst_cell_225_3 (.BL(BL3),.BLN(BLN3),.WL(WL225));
sram_cell_6t_5 inst_cell_225_4 (.BL(BL4),.BLN(BLN4),.WL(WL225));
sram_cell_6t_5 inst_cell_225_5 (.BL(BL5),.BLN(BLN5),.WL(WL225));
sram_cell_6t_5 inst_cell_225_6 (.BL(BL6),.BLN(BLN6),.WL(WL225));
sram_cell_6t_5 inst_cell_225_7 (.BL(BL7),.BLN(BLN7),.WL(WL225));
sram_cell_6t_5 inst_cell_225_8 (.BL(BL8),.BLN(BLN8),.WL(WL225));
sram_cell_6t_5 inst_cell_225_9 (.BL(BL9),.BLN(BLN9),.WL(WL225));
sram_cell_6t_5 inst_cell_225_10 (.BL(BL10),.BLN(BLN10),.WL(WL225));
sram_cell_6t_5 inst_cell_225_11 (.BL(BL11),.BLN(BLN11),.WL(WL225));
sram_cell_6t_5 inst_cell_225_12 (.BL(BL12),.BLN(BLN12),.WL(WL225));
sram_cell_6t_5 inst_cell_225_13 (.BL(BL13),.BLN(BLN13),.WL(WL225));
sram_cell_6t_5 inst_cell_225_14 (.BL(BL14),.BLN(BLN14),.WL(WL225));
sram_cell_6t_5 inst_cell_225_15 (.BL(BL15),.BLN(BLN15),.WL(WL225));
sram_cell_6t_5 inst_cell_225_16 (.BL(BL16),.BLN(BLN16),.WL(WL225));
sram_cell_6t_5 inst_cell_225_17 (.BL(BL17),.BLN(BLN17),.WL(WL225));
sram_cell_6t_5 inst_cell_225_18 (.BL(BL18),.BLN(BLN18),.WL(WL225));
sram_cell_6t_5 inst_cell_225_19 (.BL(BL19),.BLN(BLN19),.WL(WL225));
sram_cell_6t_5 inst_cell_225_20 (.BL(BL20),.BLN(BLN20),.WL(WL225));
sram_cell_6t_5 inst_cell_225_21 (.BL(BL21),.BLN(BLN21),.WL(WL225));
sram_cell_6t_5 inst_cell_225_22 (.BL(BL22),.BLN(BLN22),.WL(WL225));
sram_cell_6t_5 inst_cell_225_23 (.BL(BL23),.BLN(BLN23),.WL(WL225));
sram_cell_6t_5 inst_cell_225_24 (.BL(BL24),.BLN(BLN24),.WL(WL225));
sram_cell_6t_5 inst_cell_225_25 (.BL(BL25),.BLN(BLN25),.WL(WL225));
sram_cell_6t_5 inst_cell_225_26 (.BL(BL26),.BLN(BLN26),.WL(WL225));
sram_cell_6t_5 inst_cell_225_27 (.BL(BL27),.BLN(BLN27),.WL(WL225));
sram_cell_6t_5 inst_cell_225_28 (.BL(BL28),.BLN(BLN28),.WL(WL225));
sram_cell_6t_5 inst_cell_225_29 (.BL(BL29),.BLN(BLN29),.WL(WL225));
sram_cell_6t_5 inst_cell_225_30 (.BL(BL30),.BLN(BLN30),.WL(WL225));
sram_cell_6t_5 inst_cell_225_31 (.BL(BL31),.BLN(BLN31),.WL(WL225));
sram_cell_6t_5 inst_cell_225_32 (.BL(BL32),.BLN(BLN32),.WL(WL225));
sram_cell_6t_5 inst_cell_225_33 (.BL(BL33),.BLN(BLN33),.WL(WL225));
sram_cell_6t_5 inst_cell_225_34 (.BL(BL34),.BLN(BLN34),.WL(WL225));
sram_cell_6t_5 inst_cell_225_35 (.BL(BL35),.BLN(BLN35),.WL(WL225));
sram_cell_6t_5 inst_cell_225_36 (.BL(BL36),.BLN(BLN36),.WL(WL225));
sram_cell_6t_5 inst_cell_225_37 (.BL(BL37),.BLN(BLN37),.WL(WL225));
sram_cell_6t_5 inst_cell_225_38 (.BL(BL38),.BLN(BLN38),.WL(WL225));
sram_cell_6t_5 inst_cell_225_39 (.BL(BL39),.BLN(BLN39),.WL(WL225));
sram_cell_6t_5 inst_cell_225_40 (.BL(BL40),.BLN(BLN40),.WL(WL225));
sram_cell_6t_5 inst_cell_225_41 (.BL(BL41),.BLN(BLN41),.WL(WL225));
sram_cell_6t_5 inst_cell_225_42 (.BL(BL42),.BLN(BLN42),.WL(WL225));
sram_cell_6t_5 inst_cell_225_43 (.BL(BL43),.BLN(BLN43),.WL(WL225));
sram_cell_6t_5 inst_cell_225_44 (.BL(BL44),.BLN(BLN44),.WL(WL225));
sram_cell_6t_5 inst_cell_225_45 (.BL(BL45),.BLN(BLN45),.WL(WL225));
sram_cell_6t_5 inst_cell_225_46 (.BL(BL46),.BLN(BLN46),.WL(WL225));
sram_cell_6t_5 inst_cell_225_47 (.BL(BL47),.BLN(BLN47),.WL(WL225));
sram_cell_6t_5 inst_cell_225_48 (.BL(BL48),.BLN(BLN48),.WL(WL225));
sram_cell_6t_5 inst_cell_225_49 (.BL(BL49),.BLN(BLN49),.WL(WL225));
sram_cell_6t_5 inst_cell_225_50 (.BL(BL50),.BLN(BLN50),.WL(WL225));
sram_cell_6t_5 inst_cell_225_51 (.BL(BL51),.BLN(BLN51),.WL(WL225));
sram_cell_6t_5 inst_cell_225_52 (.BL(BL52),.BLN(BLN52),.WL(WL225));
sram_cell_6t_5 inst_cell_225_53 (.BL(BL53),.BLN(BLN53),.WL(WL225));
sram_cell_6t_5 inst_cell_225_54 (.BL(BL54),.BLN(BLN54),.WL(WL225));
sram_cell_6t_5 inst_cell_225_55 (.BL(BL55),.BLN(BLN55),.WL(WL225));
sram_cell_6t_5 inst_cell_225_56 (.BL(BL56),.BLN(BLN56),.WL(WL225));
sram_cell_6t_5 inst_cell_225_57 (.BL(BL57),.BLN(BLN57),.WL(WL225));
sram_cell_6t_5 inst_cell_225_58 (.BL(BL58),.BLN(BLN58),.WL(WL225));
sram_cell_6t_5 inst_cell_225_59 (.BL(BL59),.BLN(BLN59),.WL(WL225));
sram_cell_6t_5 inst_cell_225_60 (.BL(BL60),.BLN(BLN60),.WL(WL225));
sram_cell_6t_5 inst_cell_225_61 (.BL(BL61),.BLN(BLN61),.WL(WL225));
sram_cell_6t_5 inst_cell_225_62 (.BL(BL62),.BLN(BLN62),.WL(WL225));
sram_cell_6t_5 inst_cell_225_63 (.BL(BL63),.BLN(BLN63),.WL(WL225));
sram_cell_6t_5 inst_cell_225_64 (.BL(BL64),.BLN(BLN64),.WL(WL225));
sram_cell_6t_5 inst_cell_225_65 (.BL(BL65),.BLN(BLN65),.WL(WL225));
sram_cell_6t_5 inst_cell_225_66 (.BL(BL66),.BLN(BLN66),.WL(WL225));
sram_cell_6t_5 inst_cell_225_67 (.BL(BL67),.BLN(BLN67),.WL(WL225));
sram_cell_6t_5 inst_cell_225_68 (.BL(BL68),.BLN(BLN68),.WL(WL225));
sram_cell_6t_5 inst_cell_225_69 (.BL(BL69),.BLN(BLN69),.WL(WL225));
sram_cell_6t_5 inst_cell_225_70 (.BL(BL70),.BLN(BLN70),.WL(WL225));
sram_cell_6t_5 inst_cell_225_71 (.BL(BL71),.BLN(BLN71),.WL(WL225));
sram_cell_6t_5 inst_cell_225_72 (.BL(BL72),.BLN(BLN72),.WL(WL225));
sram_cell_6t_5 inst_cell_225_73 (.BL(BL73),.BLN(BLN73),.WL(WL225));
sram_cell_6t_5 inst_cell_225_74 (.BL(BL74),.BLN(BLN74),.WL(WL225));
sram_cell_6t_5 inst_cell_225_75 (.BL(BL75),.BLN(BLN75),.WL(WL225));
sram_cell_6t_5 inst_cell_225_76 (.BL(BL76),.BLN(BLN76),.WL(WL225));
sram_cell_6t_5 inst_cell_225_77 (.BL(BL77),.BLN(BLN77),.WL(WL225));
sram_cell_6t_5 inst_cell_225_78 (.BL(BL78),.BLN(BLN78),.WL(WL225));
sram_cell_6t_5 inst_cell_225_79 (.BL(BL79),.BLN(BLN79),.WL(WL225));
sram_cell_6t_5 inst_cell_225_80 (.BL(BL80),.BLN(BLN80),.WL(WL225));
sram_cell_6t_5 inst_cell_225_81 (.BL(BL81),.BLN(BLN81),.WL(WL225));
sram_cell_6t_5 inst_cell_225_82 (.BL(BL82),.BLN(BLN82),.WL(WL225));
sram_cell_6t_5 inst_cell_225_83 (.BL(BL83),.BLN(BLN83),.WL(WL225));
sram_cell_6t_5 inst_cell_225_84 (.BL(BL84),.BLN(BLN84),.WL(WL225));
sram_cell_6t_5 inst_cell_225_85 (.BL(BL85),.BLN(BLN85),.WL(WL225));
sram_cell_6t_5 inst_cell_225_86 (.BL(BL86),.BLN(BLN86),.WL(WL225));
sram_cell_6t_5 inst_cell_225_87 (.BL(BL87),.BLN(BLN87),.WL(WL225));
sram_cell_6t_5 inst_cell_225_88 (.BL(BL88),.BLN(BLN88),.WL(WL225));
sram_cell_6t_5 inst_cell_225_89 (.BL(BL89),.BLN(BLN89),.WL(WL225));
sram_cell_6t_5 inst_cell_225_90 (.BL(BL90),.BLN(BLN90),.WL(WL225));
sram_cell_6t_5 inst_cell_225_91 (.BL(BL91),.BLN(BLN91),.WL(WL225));
sram_cell_6t_5 inst_cell_225_92 (.BL(BL92),.BLN(BLN92),.WL(WL225));
sram_cell_6t_5 inst_cell_225_93 (.BL(BL93),.BLN(BLN93),.WL(WL225));
sram_cell_6t_5 inst_cell_225_94 (.BL(BL94),.BLN(BLN94),.WL(WL225));
sram_cell_6t_5 inst_cell_225_95 (.BL(BL95),.BLN(BLN95),.WL(WL225));
sram_cell_6t_5 inst_cell_225_96 (.BL(BL96),.BLN(BLN96),.WL(WL225));
sram_cell_6t_5 inst_cell_225_97 (.BL(BL97),.BLN(BLN97),.WL(WL225));
sram_cell_6t_5 inst_cell_225_98 (.BL(BL98),.BLN(BLN98),.WL(WL225));
sram_cell_6t_5 inst_cell_225_99 (.BL(BL99),.BLN(BLN99),.WL(WL225));
sram_cell_6t_5 inst_cell_225_100 (.BL(BL100),.BLN(BLN100),.WL(WL225));
sram_cell_6t_5 inst_cell_225_101 (.BL(BL101),.BLN(BLN101),.WL(WL225));
sram_cell_6t_5 inst_cell_225_102 (.BL(BL102),.BLN(BLN102),.WL(WL225));
sram_cell_6t_5 inst_cell_225_103 (.BL(BL103),.BLN(BLN103),.WL(WL225));
sram_cell_6t_5 inst_cell_225_104 (.BL(BL104),.BLN(BLN104),.WL(WL225));
sram_cell_6t_5 inst_cell_225_105 (.BL(BL105),.BLN(BLN105),.WL(WL225));
sram_cell_6t_5 inst_cell_225_106 (.BL(BL106),.BLN(BLN106),.WL(WL225));
sram_cell_6t_5 inst_cell_225_107 (.BL(BL107),.BLN(BLN107),.WL(WL225));
sram_cell_6t_5 inst_cell_225_108 (.BL(BL108),.BLN(BLN108),.WL(WL225));
sram_cell_6t_5 inst_cell_225_109 (.BL(BL109),.BLN(BLN109),.WL(WL225));
sram_cell_6t_5 inst_cell_225_110 (.BL(BL110),.BLN(BLN110),.WL(WL225));
sram_cell_6t_5 inst_cell_225_111 (.BL(BL111),.BLN(BLN111),.WL(WL225));
sram_cell_6t_5 inst_cell_225_112 (.BL(BL112),.BLN(BLN112),.WL(WL225));
sram_cell_6t_5 inst_cell_225_113 (.BL(BL113),.BLN(BLN113),.WL(WL225));
sram_cell_6t_5 inst_cell_225_114 (.BL(BL114),.BLN(BLN114),.WL(WL225));
sram_cell_6t_5 inst_cell_225_115 (.BL(BL115),.BLN(BLN115),.WL(WL225));
sram_cell_6t_5 inst_cell_225_116 (.BL(BL116),.BLN(BLN116),.WL(WL225));
sram_cell_6t_5 inst_cell_225_117 (.BL(BL117),.BLN(BLN117),.WL(WL225));
sram_cell_6t_5 inst_cell_225_118 (.BL(BL118),.BLN(BLN118),.WL(WL225));
sram_cell_6t_5 inst_cell_225_119 (.BL(BL119),.BLN(BLN119),.WL(WL225));
sram_cell_6t_5 inst_cell_225_120 (.BL(BL120),.BLN(BLN120),.WL(WL225));
sram_cell_6t_5 inst_cell_225_121 (.BL(BL121),.BLN(BLN121),.WL(WL225));
sram_cell_6t_5 inst_cell_225_122 (.BL(BL122),.BLN(BLN122),.WL(WL225));
sram_cell_6t_5 inst_cell_225_123 (.BL(BL123),.BLN(BLN123),.WL(WL225));
sram_cell_6t_5 inst_cell_225_124 (.BL(BL124),.BLN(BLN124),.WL(WL225));
sram_cell_6t_5 inst_cell_225_125 (.BL(BL125),.BLN(BLN125),.WL(WL225));
sram_cell_6t_5 inst_cell_225_126 (.BL(BL126),.BLN(BLN126),.WL(WL225));
sram_cell_6t_5 inst_cell_225_127 (.BL(BL127),.BLN(BLN127),.WL(WL225));
sram_cell_6t_5 inst_cell_226_0 (.BL(BL0),.BLN(BLN0),.WL(WL226));
sram_cell_6t_5 inst_cell_226_1 (.BL(BL1),.BLN(BLN1),.WL(WL226));
sram_cell_6t_5 inst_cell_226_2 (.BL(BL2),.BLN(BLN2),.WL(WL226));
sram_cell_6t_5 inst_cell_226_3 (.BL(BL3),.BLN(BLN3),.WL(WL226));
sram_cell_6t_5 inst_cell_226_4 (.BL(BL4),.BLN(BLN4),.WL(WL226));
sram_cell_6t_5 inst_cell_226_5 (.BL(BL5),.BLN(BLN5),.WL(WL226));
sram_cell_6t_5 inst_cell_226_6 (.BL(BL6),.BLN(BLN6),.WL(WL226));
sram_cell_6t_5 inst_cell_226_7 (.BL(BL7),.BLN(BLN7),.WL(WL226));
sram_cell_6t_5 inst_cell_226_8 (.BL(BL8),.BLN(BLN8),.WL(WL226));
sram_cell_6t_5 inst_cell_226_9 (.BL(BL9),.BLN(BLN9),.WL(WL226));
sram_cell_6t_5 inst_cell_226_10 (.BL(BL10),.BLN(BLN10),.WL(WL226));
sram_cell_6t_5 inst_cell_226_11 (.BL(BL11),.BLN(BLN11),.WL(WL226));
sram_cell_6t_5 inst_cell_226_12 (.BL(BL12),.BLN(BLN12),.WL(WL226));
sram_cell_6t_5 inst_cell_226_13 (.BL(BL13),.BLN(BLN13),.WL(WL226));
sram_cell_6t_5 inst_cell_226_14 (.BL(BL14),.BLN(BLN14),.WL(WL226));
sram_cell_6t_5 inst_cell_226_15 (.BL(BL15),.BLN(BLN15),.WL(WL226));
sram_cell_6t_5 inst_cell_226_16 (.BL(BL16),.BLN(BLN16),.WL(WL226));
sram_cell_6t_5 inst_cell_226_17 (.BL(BL17),.BLN(BLN17),.WL(WL226));
sram_cell_6t_5 inst_cell_226_18 (.BL(BL18),.BLN(BLN18),.WL(WL226));
sram_cell_6t_5 inst_cell_226_19 (.BL(BL19),.BLN(BLN19),.WL(WL226));
sram_cell_6t_5 inst_cell_226_20 (.BL(BL20),.BLN(BLN20),.WL(WL226));
sram_cell_6t_5 inst_cell_226_21 (.BL(BL21),.BLN(BLN21),.WL(WL226));
sram_cell_6t_5 inst_cell_226_22 (.BL(BL22),.BLN(BLN22),.WL(WL226));
sram_cell_6t_5 inst_cell_226_23 (.BL(BL23),.BLN(BLN23),.WL(WL226));
sram_cell_6t_5 inst_cell_226_24 (.BL(BL24),.BLN(BLN24),.WL(WL226));
sram_cell_6t_5 inst_cell_226_25 (.BL(BL25),.BLN(BLN25),.WL(WL226));
sram_cell_6t_5 inst_cell_226_26 (.BL(BL26),.BLN(BLN26),.WL(WL226));
sram_cell_6t_5 inst_cell_226_27 (.BL(BL27),.BLN(BLN27),.WL(WL226));
sram_cell_6t_5 inst_cell_226_28 (.BL(BL28),.BLN(BLN28),.WL(WL226));
sram_cell_6t_5 inst_cell_226_29 (.BL(BL29),.BLN(BLN29),.WL(WL226));
sram_cell_6t_5 inst_cell_226_30 (.BL(BL30),.BLN(BLN30),.WL(WL226));
sram_cell_6t_5 inst_cell_226_31 (.BL(BL31),.BLN(BLN31),.WL(WL226));
sram_cell_6t_5 inst_cell_226_32 (.BL(BL32),.BLN(BLN32),.WL(WL226));
sram_cell_6t_5 inst_cell_226_33 (.BL(BL33),.BLN(BLN33),.WL(WL226));
sram_cell_6t_5 inst_cell_226_34 (.BL(BL34),.BLN(BLN34),.WL(WL226));
sram_cell_6t_5 inst_cell_226_35 (.BL(BL35),.BLN(BLN35),.WL(WL226));
sram_cell_6t_5 inst_cell_226_36 (.BL(BL36),.BLN(BLN36),.WL(WL226));
sram_cell_6t_5 inst_cell_226_37 (.BL(BL37),.BLN(BLN37),.WL(WL226));
sram_cell_6t_5 inst_cell_226_38 (.BL(BL38),.BLN(BLN38),.WL(WL226));
sram_cell_6t_5 inst_cell_226_39 (.BL(BL39),.BLN(BLN39),.WL(WL226));
sram_cell_6t_5 inst_cell_226_40 (.BL(BL40),.BLN(BLN40),.WL(WL226));
sram_cell_6t_5 inst_cell_226_41 (.BL(BL41),.BLN(BLN41),.WL(WL226));
sram_cell_6t_5 inst_cell_226_42 (.BL(BL42),.BLN(BLN42),.WL(WL226));
sram_cell_6t_5 inst_cell_226_43 (.BL(BL43),.BLN(BLN43),.WL(WL226));
sram_cell_6t_5 inst_cell_226_44 (.BL(BL44),.BLN(BLN44),.WL(WL226));
sram_cell_6t_5 inst_cell_226_45 (.BL(BL45),.BLN(BLN45),.WL(WL226));
sram_cell_6t_5 inst_cell_226_46 (.BL(BL46),.BLN(BLN46),.WL(WL226));
sram_cell_6t_5 inst_cell_226_47 (.BL(BL47),.BLN(BLN47),.WL(WL226));
sram_cell_6t_5 inst_cell_226_48 (.BL(BL48),.BLN(BLN48),.WL(WL226));
sram_cell_6t_5 inst_cell_226_49 (.BL(BL49),.BLN(BLN49),.WL(WL226));
sram_cell_6t_5 inst_cell_226_50 (.BL(BL50),.BLN(BLN50),.WL(WL226));
sram_cell_6t_5 inst_cell_226_51 (.BL(BL51),.BLN(BLN51),.WL(WL226));
sram_cell_6t_5 inst_cell_226_52 (.BL(BL52),.BLN(BLN52),.WL(WL226));
sram_cell_6t_5 inst_cell_226_53 (.BL(BL53),.BLN(BLN53),.WL(WL226));
sram_cell_6t_5 inst_cell_226_54 (.BL(BL54),.BLN(BLN54),.WL(WL226));
sram_cell_6t_5 inst_cell_226_55 (.BL(BL55),.BLN(BLN55),.WL(WL226));
sram_cell_6t_5 inst_cell_226_56 (.BL(BL56),.BLN(BLN56),.WL(WL226));
sram_cell_6t_5 inst_cell_226_57 (.BL(BL57),.BLN(BLN57),.WL(WL226));
sram_cell_6t_5 inst_cell_226_58 (.BL(BL58),.BLN(BLN58),.WL(WL226));
sram_cell_6t_5 inst_cell_226_59 (.BL(BL59),.BLN(BLN59),.WL(WL226));
sram_cell_6t_5 inst_cell_226_60 (.BL(BL60),.BLN(BLN60),.WL(WL226));
sram_cell_6t_5 inst_cell_226_61 (.BL(BL61),.BLN(BLN61),.WL(WL226));
sram_cell_6t_5 inst_cell_226_62 (.BL(BL62),.BLN(BLN62),.WL(WL226));
sram_cell_6t_5 inst_cell_226_63 (.BL(BL63),.BLN(BLN63),.WL(WL226));
sram_cell_6t_5 inst_cell_226_64 (.BL(BL64),.BLN(BLN64),.WL(WL226));
sram_cell_6t_5 inst_cell_226_65 (.BL(BL65),.BLN(BLN65),.WL(WL226));
sram_cell_6t_5 inst_cell_226_66 (.BL(BL66),.BLN(BLN66),.WL(WL226));
sram_cell_6t_5 inst_cell_226_67 (.BL(BL67),.BLN(BLN67),.WL(WL226));
sram_cell_6t_5 inst_cell_226_68 (.BL(BL68),.BLN(BLN68),.WL(WL226));
sram_cell_6t_5 inst_cell_226_69 (.BL(BL69),.BLN(BLN69),.WL(WL226));
sram_cell_6t_5 inst_cell_226_70 (.BL(BL70),.BLN(BLN70),.WL(WL226));
sram_cell_6t_5 inst_cell_226_71 (.BL(BL71),.BLN(BLN71),.WL(WL226));
sram_cell_6t_5 inst_cell_226_72 (.BL(BL72),.BLN(BLN72),.WL(WL226));
sram_cell_6t_5 inst_cell_226_73 (.BL(BL73),.BLN(BLN73),.WL(WL226));
sram_cell_6t_5 inst_cell_226_74 (.BL(BL74),.BLN(BLN74),.WL(WL226));
sram_cell_6t_5 inst_cell_226_75 (.BL(BL75),.BLN(BLN75),.WL(WL226));
sram_cell_6t_5 inst_cell_226_76 (.BL(BL76),.BLN(BLN76),.WL(WL226));
sram_cell_6t_5 inst_cell_226_77 (.BL(BL77),.BLN(BLN77),.WL(WL226));
sram_cell_6t_5 inst_cell_226_78 (.BL(BL78),.BLN(BLN78),.WL(WL226));
sram_cell_6t_5 inst_cell_226_79 (.BL(BL79),.BLN(BLN79),.WL(WL226));
sram_cell_6t_5 inst_cell_226_80 (.BL(BL80),.BLN(BLN80),.WL(WL226));
sram_cell_6t_5 inst_cell_226_81 (.BL(BL81),.BLN(BLN81),.WL(WL226));
sram_cell_6t_5 inst_cell_226_82 (.BL(BL82),.BLN(BLN82),.WL(WL226));
sram_cell_6t_5 inst_cell_226_83 (.BL(BL83),.BLN(BLN83),.WL(WL226));
sram_cell_6t_5 inst_cell_226_84 (.BL(BL84),.BLN(BLN84),.WL(WL226));
sram_cell_6t_5 inst_cell_226_85 (.BL(BL85),.BLN(BLN85),.WL(WL226));
sram_cell_6t_5 inst_cell_226_86 (.BL(BL86),.BLN(BLN86),.WL(WL226));
sram_cell_6t_5 inst_cell_226_87 (.BL(BL87),.BLN(BLN87),.WL(WL226));
sram_cell_6t_5 inst_cell_226_88 (.BL(BL88),.BLN(BLN88),.WL(WL226));
sram_cell_6t_5 inst_cell_226_89 (.BL(BL89),.BLN(BLN89),.WL(WL226));
sram_cell_6t_5 inst_cell_226_90 (.BL(BL90),.BLN(BLN90),.WL(WL226));
sram_cell_6t_5 inst_cell_226_91 (.BL(BL91),.BLN(BLN91),.WL(WL226));
sram_cell_6t_5 inst_cell_226_92 (.BL(BL92),.BLN(BLN92),.WL(WL226));
sram_cell_6t_5 inst_cell_226_93 (.BL(BL93),.BLN(BLN93),.WL(WL226));
sram_cell_6t_5 inst_cell_226_94 (.BL(BL94),.BLN(BLN94),.WL(WL226));
sram_cell_6t_5 inst_cell_226_95 (.BL(BL95),.BLN(BLN95),.WL(WL226));
sram_cell_6t_5 inst_cell_226_96 (.BL(BL96),.BLN(BLN96),.WL(WL226));
sram_cell_6t_5 inst_cell_226_97 (.BL(BL97),.BLN(BLN97),.WL(WL226));
sram_cell_6t_5 inst_cell_226_98 (.BL(BL98),.BLN(BLN98),.WL(WL226));
sram_cell_6t_5 inst_cell_226_99 (.BL(BL99),.BLN(BLN99),.WL(WL226));
sram_cell_6t_5 inst_cell_226_100 (.BL(BL100),.BLN(BLN100),.WL(WL226));
sram_cell_6t_5 inst_cell_226_101 (.BL(BL101),.BLN(BLN101),.WL(WL226));
sram_cell_6t_5 inst_cell_226_102 (.BL(BL102),.BLN(BLN102),.WL(WL226));
sram_cell_6t_5 inst_cell_226_103 (.BL(BL103),.BLN(BLN103),.WL(WL226));
sram_cell_6t_5 inst_cell_226_104 (.BL(BL104),.BLN(BLN104),.WL(WL226));
sram_cell_6t_5 inst_cell_226_105 (.BL(BL105),.BLN(BLN105),.WL(WL226));
sram_cell_6t_5 inst_cell_226_106 (.BL(BL106),.BLN(BLN106),.WL(WL226));
sram_cell_6t_5 inst_cell_226_107 (.BL(BL107),.BLN(BLN107),.WL(WL226));
sram_cell_6t_5 inst_cell_226_108 (.BL(BL108),.BLN(BLN108),.WL(WL226));
sram_cell_6t_5 inst_cell_226_109 (.BL(BL109),.BLN(BLN109),.WL(WL226));
sram_cell_6t_5 inst_cell_226_110 (.BL(BL110),.BLN(BLN110),.WL(WL226));
sram_cell_6t_5 inst_cell_226_111 (.BL(BL111),.BLN(BLN111),.WL(WL226));
sram_cell_6t_5 inst_cell_226_112 (.BL(BL112),.BLN(BLN112),.WL(WL226));
sram_cell_6t_5 inst_cell_226_113 (.BL(BL113),.BLN(BLN113),.WL(WL226));
sram_cell_6t_5 inst_cell_226_114 (.BL(BL114),.BLN(BLN114),.WL(WL226));
sram_cell_6t_5 inst_cell_226_115 (.BL(BL115),.BLN(BLN115),.WL(WL226));
sram_cell_6t_5 inst_cell_226_116 (.BL(BL116),.BLN(BLN116),.WL(WL226));
sram_cell_6t_5 inst_cell_226_117 (.BL(BL117),.BLN(BLN117),.WL(WL226));
sram_cell_6t_5 inst_cell_226_118 (.BL(BL118),.BLN(BLN118),.WL(WL226));
sram_cell_6t_5 inst_cell_226_119 (.BL(BL119),.BLN(BLN119),.WL(WL226));
sram_cell_6t_5 inst_cell_226_120 (.BL(BL120),.BLN(BLN120),.WL(WL226));
sram_cell_6t_5 inst_cell_226_121 (.BL(BL121),.BLN(BLN121),.WL(WL226));
sram_cell_6t_5 inst_cell_226_122 (.BL(BL122),.BLN(BLN122),.WL(WL226));
sram_cell_6t_5 inst_cell_226_123 (.BL(BL123),.BLN(BLN123),.WL(WL226));
sram_cell_6t_5 inst_cell_226_124 (.BL(BL124),.BLN(BLN124),.WL(WL226));
sram_cell_6t_5 inst_cell_226_125 (.BL(BL125),.BLN(BLN125),.WL(WL226));
sram_cell_6t_5 inst_cell_226_126 (.BL(BL126),.BLN(BLN126),.WL(WL226));
sram_cell_6t_5 inst_cell_226_127 (.BL(BL127),.BLN(BLN127),.WL(WL226));
sram_cell_6t_5 inst_cell_227_0 (.BL(BL0),.BLN(BLN0),.WL(WL227));
sram_cell_6t_5 inst_cell_227_1 (.BL(BL1),.BLN(BLN1),.WL(WL227));
sram_cell_6t_5 inst_cell_227_2 (.BL(BL2),.BLN(BLN2),.WL(WL227));
sram_cell_6t_5 inst_cell_227_3 (.BL(BL3),.BLN(BLN3),.WL(WL227));
sram_cell_6t_5 inst_cell_227_4 (.BL(BL4),.BLN(BLN4),.WL(WL227));
sram_cell_6t_5 inst_cell_227_5 (.BL(BL5),.BLN(BLN5),.WL(WL227));
sram_cell_6t_5 inst_cell_227_6 (.BL(BL6),.BLN(BLN6),.WL(WL227));
sram_cell_6t_5 inst_cell_227_7 (.BL(BL7),.BLN(BLN7),.WL(WL227));
sram_cell_6t_5 inst_cell_227_8 (.BL(BL8),.BLN(BLN8),.WL(WL227));
sram_cell_6t_5 inst_cell_227_9 (.BL(BL9),.BLN(BLN9),.WL(WL227));
sram_cell_6t_5 inst_cell_227_10 (.BL(BL10),.BLN(BLN10),.WL(WL227));
sram_cell_6t_5 inst_cell_227_11 (.BL(BL11),.BLN(BLN11),.WL(WL227));
sram_cell_6t_5 inst_cell_227_12 (.BL(BL12),.BLN(BLN12),.WL(WL227));
sram_cell_6t_5 inst_cell_227_13 (.BL(BL13),.BLN(BLN13),.WL(WL227));
sram_cell_6t_5 inst_cell_227_14 (.BL(BL14),.BLN(BLN14),.WL(WL227));
sram_cell_6t_5 inst_cell_227_15 (.BL(BL15),.BLN(BLN15),.WL(WL227));
sram_cell_6t_5 inst_cell_227_16 (.BL(BL16),.BLN(BLN16),.WL(WL227));
sram_cell_6t_5 inst_cell_227_17 (.BL(BL17),.BLN(BLN17),.WL(WL227));
sram_cell_6t_5 inst_cell_227_18 (.BL(BL18),.BLN(BLN18),.WL(WL227));
sram_cell_6t_5 inst_cell_227_19 (.BL(BL19),.BLN(BLN19),.WL(WL227));
sram_cell_6t_5 inst_cell_227_20 (.BL(BL20),.BLN(BLN20),.WL(WL227));
sram_cell_6t_5 inst_cell_227_21 (.BL(BL21),.BLN(BLN21),.WL(WL227));
sram_cell_6t_5 inst_cell_227_22 (.BL(BL22),.BLN(BLN22),.WL(WL227));
sram_cell_6t_5 inst_cell_227_23 (.BL(BL23),.BLN(BLN23),.WL(WL227));
sram_cell_6t_5 inst_cell_227_24 (.BL(BL24),.BLN(BLN24),.WL(WL227));
sram_cell_6t_5 inst_cell_227_25 (.BL(BL25),.BLN(BLN25),.WL(WL227));
sram_cell_6t_5 inst_cell_227_26 (.BL(BL26),.BLN(BLN26),.WL(WL227));
sram_cell_6t_5 inst_cell_227_27 (.BL(BL27),.BLN(BLN27),.WL(WL227));
sram_cell_6t_5 inst_cell_227_28 (.BL(BL28),.BLN(BLN28),.WL(WL227));
sram_cell_6t_5 inst_cell_227_29 (.BL(BL29),.BLN(BLN29),.WL(WL227));
sram_cell_6t_5 inst_cell_227_30 (.BL(BL30),.BLN(BLN30),.WL(WL227));
sram_cell_6t_5 inst_cell_227_31 (.BL(BL31),.BLN(BLN31),.WL(WL227));
sram_cell_6t_5 inst_cell_227_32 (.BL(BL32),.BLN(BLN32),.WL(WL227));
sram_cell_6t_5 inst_cell_227_33 (.BL(BL33),.BLN(BLN33),.WL(WL227));
sram_cell_6t_5 inst_cell_227_34 (.BL(BL34),.BLN(BLN34),.WL(WL227));
sram_cell_6t_5 inst_cell_227_35 (.BL(BL35),.BLN(BLN35),.WL(WL227));
sram_cell_6t_5 inst_cell_227_36 (.BL(BL36),.BLN(BLN36),.WL(WL227));
sram_cell_6t_5 inst_cell_227_37 (.BL(BL37),.BLN(BLN37),.WL(WL227));
sram_cell_6t_5 inst_cell_227_38 (.BL(BL38),.BLN(BLN38),.WL(WL227));
sram_cell_6t_5 inst_cell_227_39 (.BL(BL39),.BLN(BLN39),.WL(WL227));
sram_cell_6t_5 inst_cell_227_40 (.BL(BL40),.BLN(BLN40),.WL(WL227));
sram_cell_6t_5 inst_cell_227_41 (.BL(BL41),.BLN(BLN41),.WL(WL227));
sram_cell_6t_5 inst_cell_227_42 (.BL(BL42),.BLN(BLN42),.WL(WL227));
sram_cell_6t_5 inst_cell_227_43 (.BL(BL43),.BLN(BLN43),.WL(WL227));
sram_cell_6t_5 inst_cell_227_44 (.BL(BL44),.BLN(BLN44),.WL(WL227));
sram_cell_6t_5 inst_cell_227_45 (.BL(BL45),.BLN(BLN45),.WL(WL227));
sram_cell_6t_5 inst_cell_227_46 (.BL(BL46),.BLN(BLN46),.WL(WL227));
sram_cell_6t_5 inst_cell_227_47 (.BL(BL47),.BLN(BLN47),.WL(WL227));
sram_cell_6t_5 inst_cell_227_48 (.BL(BL48),.BLN(BLN48),.WL(WL227));
sram_cell_6t_5 inst_cell_227_49 (.BL(BL49),.BLN(BLN49),.WL(WL227));
sram_cell_6t_5 inst_cell_227_50 (.BL(BL50),.BLN(BLN50),.WL(WL227));
sram_cell_6t_5 inst_cell_227_51 (.BL(BL51),.BLN(BLN51),.WL(WL227));
sram_cell_6t_5 inst_cell_227_52 (.BL(BL52),.BLN(BLN52),.WL(WL227));
sram_cell_6t_5 inst_cell_227_53 (.BL(BL53),.BLN(BLN53),.WL(WL227));
sram_cell_6t_5 inst_cell_227_54 (.BL(BL54),.BLN(BLN54),.WL(WL227));
sram_cell_6t_5 inst_cell_227_55 (.BL(BL55),.BLN(BLN55),.WL(WL227));
sram_cell_6t_5 inst_cell_227_56 (.BL(BL56),.BLN(BLN56),.WL(WL227));
sram_cell_6t_5 inst_cell_227_57 (.BL(BL57),.BLN(BLN57),.WL(WL227));
sram_cell_6t_5 inst_cell_227_58 (.BL(BL58),.BLN(BLN58),.WL(WL227));
sram_cell_6t_5 inst_cell_227_59 (.BL(BL59),.BLN(BLN59),.WL(WL227));
sram_cell_6t_5 inst_cell_227_60 (.BL(BL60),.BLN(BLN60),.WL(WL227));
sram_cell_6t_5 inst_cell_227_61 (.BL(BL61),.BLN(BLN61),.WL(WL227));
sram_cell_6t_5 inst_cell_227_62 (.BL(BL62),.BLN(BLN62),.WL(WL227));
sram_cell_6t_5 inst_cell_227_63 (.BL(BL63),.BLN(BLN63),.WL(WL227));
sram_cell_6t_5 inst_cell_227_64 (.BL(BL64),.BLN(BLN64),.WL(WL227));
sram_cell_6t_5 inst_cell_227_65 (.BL(BL65),.BLN(BLN65),.WL(WL227));
sram_cell_6t_5 inst_cell_227_66 (.BL(BL66),.BLN(BLN66),.WL(WL227));
sram_cell_6t_5 inst_cell_227_67 (.BL(BL67),.BLN(BLN67),.WL(WL227));
sram_cell_6t_5 inst_cell_227_68 (.BL(BL68),.BLN(BLN68),.WL(WL227));
sram_cell_6t_5 inst_cell_227_69 (.BL(BL69),.BLN(BLN69),.WL(WL227));
sram_cell_6t_5 inst_cell_227_70 (.BL(BL70),.BLN(BLN70),.WL(WL227));
sram_cell_6t_5 inst_cell_227_71 (.BL(BL71),.BLN(BLN71),.WL(WL227));
sram_cell_6t_5 inst_cell_227_72 (.BL(BL72),.BLN(BLN72),.WL(WL227));
sram_cell_6t_5 inst_cell_227_73 (.BL(BL73),.BLN(BLN73),.WL(WL227));
sram_cell_6t_5 inst_cell_227_74 (.BL(BL74),.BLN(BLN74),.WL(WL227));
sram_cell_6t_5 inst_cell_227_75 (.BL(BL75),.BLN(BLN75),.WL(WL227));
sram_cell_6t_5 inst_cell_227_76 (.BL(BL76),.BLN(BLN76),.WL(WL227));
sram_cell_6t_5 inst_cell_227_77 (.BL(BL77),.BLN(BLN77),.WL(WL227));
sram_cell_6t_5 inst_cell_227_78 (.BL(BL78),.BLN(BLN78),.WL(WL227));
sram_cell_6t_5 inst_cell_227_79 (.BL(BL79),.BLN(BLN79),.WL(WL227));
sram_cell_6t_5 inst_cell_227_80 (.BL(BL80),.BLN(BLN80),.WL(WL227));
sram_cell_6t_5 inst_cell_227_81 (.BL(BL81),.BLN(BLN81),.WL(WL227));
sram_cell_6t_5 inst_cell_227_82 (.BL(BL82),.BLN(BLN82),.WL(WL227));
sram_cell_6t_5 inst_cell_227_83 (.BL(BL83),.BLN(BLN83),.WL(WL227));
sram_cell_6t_5 inst_cell_227_84 (.BL(BL84),.BLN(BLN84),.WL(WL227));
sram_cell_6t_5 inst_cell_227_85 (.BL(BL85),.BLN(BLN85),.WL(WL227));
sram_cell_6t_5 inst_cell_227_86 (.BL(BL86),.BLN(BLN86),.WL(WL227));
sram_cell_6t_5 inst_cell_227_87 (.BL(BL87),.BLN(BLN87),.WL(WL227));
sram_cell_6t_5 inst_cell_227_88 (.BL(BL88),.BLN(BLN88),.WL(WL227));
sram_cell_6t_5 inst_cell_227_89 (.BL(BL89),.BLN(BLN89),.WL(WL227));
sram_cell_6t_5 inst_cell_227_90 (.BL(BL90),.BLN(BLN90),.WL(WL227));
sram_cell_6t_5 inst_cell_227_91 (.BL(BL91),.BLN(BLN91),.WL(WL227));
sram_cell_6t_5 inst_cell_227_92 (.BL(BL92),.BLN(BLN92),.WL(WL227));
sram_cell_6t_5 inst_cell_227_93 (.BL(BL93),.BLN(BLN93),.WL(WL227));
sram_cell_6t_5 inst_cell_227_94 (.BL(BL94),.BLN(BLN94),.WL(WL227));
sram_cell_6t_5 inst_cell_227_95 (.BL(BL95),.BLN(BLN95),.WL(WL227));
sram_cell_6t_5 inst_cell_227_96 (.BL(BL96),.BLN(BLN96),.WL(WL227));
sram_cell_6t_5 inst_cell_227_97 (.BL(BL97),.BLN(BLN97),.WL(WL227));
sram_cell_6t_5 inst_cell_227_98 (.BL(BL98),.BLN(BLN98),.WL(WL227));
sram_cell_6t_5 inst_cell_227_99 (.BL(BL99),.BLN(BLN99),.WL(WL227));
sram_cell_6t_5 inst_cell_227_100 (.BL(BL100),.BLN(BLN100),.WL(WL227));
sram_cell_6t_5 inst_cell_227_101 (.BL(BL101),.BLN(BLN101),.WL(WL227));
sram_cell_6t_5 inst_cell_227_102 (.BL(BL102),.BLN(BLN102),.WL(WL227));
sram_cell_6t_5 inst_cell_227_103 (.BL(BL103),.BLN(BLN103),.WL(WL227));
sram_cell_6t_5 inst_cell_227_104 (.BL(BL104),.BLN(BLN104),.WL(WL227));
sram_cell_6t_5 inst_cell_227_105 (.BL(BL105),.BLN(BLN105),.WL(WL227));
sram_cell_6t_5 inst_cell_227_106 (.BL(BL106),.BLN(BLN106),.WL(WL227));
sram_cell_6t_5 inst_cell_227_107 (.BL(BL107),.BLN(BLN107),.WL(WL227));
sram_cell_6t_5 inst_cell_227_108 (.BL(BL108),.BLN(BLN108),.WL(WL227));
sram_cell_6t_5 inst_cell_227_109 (.BL(BL109),.BLN(BLN109),.WL(WL227));
sram_cell_6t_5 inst_cell_227_110 (.BL(BL110),.BLN(BLN110),.WL(WL227));
sram_cell_6t_5 inst_cell_227_111 (.BL(BL111),.BLN(BLN111),.WL(WL227));
sram_cell_6t_5 inst_cell_227_112 (.BL(BL112),.BLN(BLN112),.WL(WL227));
sram_cell_6t_5 inst_cell_227_113 (.BL(BL113),.BLN(BLN113),.WL(WL227));
sram_cell_6t_5 inst_cell_227_114 (.BL(BL114),.BLN(BLN114),.WL(WL227));
sram_cell_6t_5 inst_cell_227_115 (.BL(BL115),.BLN(BLN115),.WL(WL227));
sram_cell_6t_5 inst_cell_227_116 (.BL(BL116),.BLN(BLN116),.WL(WL227));
sram_cell_6t_5 inst_cell_227_117 (.BL(BL117),.BLN(BLN117),.WL(WL227));
sram_cell_6t_5 inst_cell_227_118 (.BL(BL118),.BLN(BLN118),.WL(WL227));
sram_cell_6t_5 inst_cell_227_119 (.BL(BL119),.BLN(BLN119),.WL(WL227));
sram_cell_6t_5 inst_cell_227_120 (.BL(BL120),.BLN(BLN120),.WL(WL227));
sram_cell_6t_5 inst_cell_227_121 (.BL(BL121),.BLN(BLN121),.WL(WL227));
sram_cell_6t_5 inst_cell_227_122 (.BL(BL122),.BLN(BLN122),.WL(WL227));
sram_cell_6t_5 inst_cell_227_123 (.BL(BL123),.BLN(BLN123),.WL(WL227));
sram_cell_6t_5 inst_cell_227_124 (.BL(BL124),.BLN(BLN124),.WL(WL227));
sram_cell_6t_5 inst_cell_227_125 (.BL(BL125),.BLN(BLN125),.WL(WL227));
sram_cell_6t_5 inst_cell_227_126 (.BL(BL126),.BLN(BLN126),.WL(WL227));
sram_cell_6t_5 inst_cell_227_127 (.BL(BL127),.BLN(BLN127),.WL(WL227));
sram_cell_6t_5 inst_cell_228_0 (.BL(BL0),.BLN(BLN0),.WL(WL228));
sram_cell_6t_5 inst_cell_228_1 (.BL(BL1),.BLN(BLN1),.WL(WL228));
sram_cell_6t_5 inst_cell_228_2 (.BL(BL2),.BLN(BLN2),.WL(WL228));
sram_cell_6t_5 inst_cell_228_3 (.BL(BL3),.BLN(BLN3),.WL(WL228));
sram_cell_6t_5 inst_cell_228_4 (.BL(BL4),.BLN(BLN4),.WL(WL228));
sram_cell_6t_5 inst_cell_228_5 (.BL(BL5),.BLN(BLN5),.WL(WL228));
sram_cell_6t_5 inst_cell_228_6 (.BL(BL6),.BLN(BLN6),.WL(WL228));
sram_cell_6t_5 inst_cell_228_7 (.BL(BL7),.BLN(BLN7),.WL(WL228));
sram_cell_6t_5 inst_cell_228_8 (.BL(BL8),.BLN(BLN8),.WL(WL228));
sram_cell_6t_5 inst_cell_228_9 (.BL(BL9),.BLN(BLN9),.WL(WL228));
sram_cell_6t_5 inst_cell_228_10 (.BL(BL10),.BLN(BLN10),.WL(WL228));
sram_cell_6t_5 inst_cell_228_11 (.BL(BL11),.BLN(BLN11),.WL(WL228));
sram_cell_6t_5 inst_cell_228_12 (.BL(BL12),.BLN(BLN12),.WL(WL228));
sram_cell_6t_5 inst_cell_228_13 (.BL(BL13),.BLN(BLN13),.WL(WL228));
sram_cell_6t_5 inst_cell_228_14 (.BL(BL14),.BLN(BLN14),.WL(WL228));
sram_cell_6t_5 inst_cell_228_15 (.BL(BL15),.BLN(BLN15),.WL(WL228));
sram_cell_6t_5 inst_cell_228_16 (.BL(BL16),.BLN(BLN16),.WL(WL228));
sram_cell_6t_5 inst_cell_228_17 (.BL(BL17),.BLN(BLN17),.WL(WL228));
sram_cell_6t_5 inst_cell_228_18 (.BL(BL18),.BLN(BLN18),.WL(WL228));
sram_cell_6t_5 inst_cell_228_19 (.BL(BL19),.BLN(BLN19),.WL(WL228));
sram_cell_6t_5 inst_cell_228_20 (.BL(BL20),.BLN(BLN20),.WL(WL228));
sram_cell_6t_5 inst_cell_228_21 (.BL(BL21),.BLN(BLN21),.WL(WL228));
sram_cell_6t_5 inst_cell_228_22 (.BL(BL22),.BLN(BLN22),.WL(WL228));
sram_cell_6t_5 inst_cell_228_23 (.BL(BL23),.BLN(BLN23),.WL(WL228));
sram_cell_6t_5 inst_cell_228_24 (.BL(BL24),.BLN(BLN24),.WL(WL228));
sram_cell_6t_5 inst_cell_228_25 (.BL(BL25),.BLN(BLN25),.WL(WL228));
sram_cell_6t_5 inst_cell_228_26 (.BL(BL26),.BLN(BLN26),.WL(WL228));
sram_cell_6t_5 inst_cell_228_27 (.BL(BL27),.BLN(BLN27),.WL(WL228));
sram_cell_6t_5 inst_cell_228_28 (.BL(BL28),.BLN(BLN28),.WL(WL228));
sram_cell_6t_5 inst_cell_228_29 (.BL(BL29),.BLN(BLN29),.WL(WL228));
sram_cell_6t_5 inst_cell_228_30 (.BL(BL30),.BLN(BLN30),.WL(WL228));
sram_cell_6t_5 inst_cell_228_31 (.BL(BL31),.BLN(BLN31),.WL(WL228));
sram_cell_6t_5 inst_cell_228_32 (.BL(BL32),.BLN(BLN32),.WL(WL228));
sram_cell_6t_5 inst_cell_228_33 (.BL(BL33),.BLN(BLN33),.WL(WL228));
sram_cell_6t_5 inst_cell_228_34 (.BL(BL34),.BLN(BLN34),.WL(WL228));
sram_cell_6t_5 inst_cell_228_35 (.BL(BL35),.BLN(BLN35),.WL(WL228));
sram_cell_6t_5 inst_cell_228_36 (.BL(BL36),.BLN(BLN36),.WL(WL228));
sram_cell_6t_5 inst_cell_228_37 (.BL(BL37),.BLN(BLN37),.WL(WL228));
sram_cell_6t_5 inst_cell_228_38 (.BL(BL38),.BLN(BLN38),.WL(WL228));
sram_cell_6t_5 inst_cell_228_39 (.BL(BL39),.BLN(BLN39),.WL(WL228));
sram_cell_6t_5 inst_cell_228_40 (.BL(BL40),.BLN(BLN40),.WL(WL228));
sram_cell_6t_5 inst_cell_228_41 (.BL(BL41),.BLN(BLN41),.WL(WL228));
sram_cell_6t_5 inst_cell_228_42 (.BL(BL42),.BLN(BLN42),.WL(WL228));
sram_cell_6t_5 inst_cell_228_43 (.BL(BL43),.BLN(BLN43),.WL(WL228));
sram_cell_6t_5 inst_cell_228_44 (.BL(BL44),.BLN(BLN44),.WL(WL228));
sram_cell_6t_5 inst_cell_228_45 (.BL(BL45),.BLN(BLN45),.WL(WL228));
sram_cell_6t_5 inst_cell_228_46 (.BL(BL46),.BLN(BLN46),.WL(WL228));
sram_cell_6t_5 inst_cell_228_47 (.BL(BL47),.BLN(BLN47),.WL(WL228));
sram_cell_6t_5 inst_cell_228_48 (.BL(BL48),.BLN(BLN48),.WL(WL228));
sram_cell_6t_5 inst_cell_228_49 (.BL(BL49),.BLN(BLN49),.WL(WL228));
sram_cell_6t_5 inst_cell_228_50 (.BL(BL50),.BLN(BLN50),.WL(WL228));
sram_cell_6t_5 inst_cell_228_51 (.BL(BL51),.BLN(BLN51),.WL(WL228));
sram_cell_6t_5 inst_cell_228_52 (.BL(BL52),.BLN(BLN52),.WL(WL228));
sram_cell_6t_5 inst_cell_228_53 (.BL(BL53),.BLN(BLN53),.WL(WL228));
sram_cell_6t_5 inst_cell_228_54 (.BL(BL54),.BLN(BLN54),.WL(WL228));
sram_cell_6t_5 inst_cell_228_55 (.BL(BL55),.BLN(BLN55),.WL(WL228));
sram_cell_6t_5 inst_cell_228_56 (.BL(BL56),.BLN(BLN56),.WL(WL228));
sram_cell_6t_5 inst_cell_228_57 (.BL(BL57),.BLN(BLN57),.WL(WL228));
sram_cell_6t_5 inst_cell_228_58 (.BL(BL58),.BLN(BLN58),.WL(WL228));
sram_cell_6t_5 inst_cell_228_59 (.BL(BL59),.BLN(BLN59),.WL(WL228));
sram_cell_6t_5 inst_cell_228_60 (.BL(BL60),.BLN(BLN60),.WL(WL228));
sram_cell_6t_5 inst_cell_228_61 (.BL(BL61),.BLN(BLN61),.WL(WL228));
sram_cell_6t_5 inst_cell_228_62 (.BL(BL62),.BLN(BLN62),.WL(WL228));
sram_cell_6t_5 inst_cell_228_63 (.BL(BL63),.BLN(BLN63),.WL(WL228));
sram_cell_6t_5 inst_cell_228_64 (.BL(BL64),.BLN(BLN64),.WL(WL228));
sram_cell_6t_5 inst_cell_228_65 (.BL(BL65),.BLN(BLN65),.WL(WL228));
sram_cell_6t_5 inst_cell_228_66 (.BL(BL66),.BLN(BLN66),.WL(WL228));
sram_cell_6t_5 inst_cell_228_67 (.BL(BL67),.BLN(BLN67),.WL(WL228));
sram_cell_6t_5 inst_cell_228_68 (.BL(BL68),.BLN(BLN68),.WL(WL228));
sram_cell_6t_5 inst_cell_228_69 (.BL(BL69),.BLN(BLN69),.WL(WL228));
sram_cell_6t_5 inst_cell_228_70 (.BL(BL70),.BLN(BLN70),.WL(WL228));
sram_cell_6t_5 inst_cell_228_71 (.BL(BL71),.BLN(BLN71),.WL(WL228));
sram_cell_6t_5 inst_cell_228_72 (.BL(BL72),.BLN(BLN72),.WL(WL228));
sram_cell_6t_5 inst_cell_228_73 (.BL(BL73),.BLN(BLN73),.WL(WL228));
sram_cell_6t_5 inst_cell_228_74 (.BL(BL74),.BLN(BLN74),.WL(WL228));
sram_cell_6t_5 inst_cell_228_75 (.BL(BL75),.BLN(BLN75),.WL(WL228));
sram_cell_6t_5 inst_cell_228_76 (.BL(BL76),.BLN(BLN76),.WL(WL228));
sram_cell_6t_5 inst_cell_228_77 (.BL(BL77),.BLN(BLN77),.WL(WL228));
sram_cell_6t_5 inst_cell_228_78 (.BL(BL78),.BLN(BLN78),.WL(WL228));
sram_cell_6t_5 inst_cell_228_79 (.BL(BL79),.BLN(BLN79),.WL(WL228));
sram_cell_6t_5 inst_cell_228_80 (.BL(BL80),.BLN(BLN80),.WL(WL228));
sram_cell_6t_5 inst_cell_228_81 (.BL(BL81),.BLN(BLN81),.WL(WL228));
sram_cell_6t_5 inst_cell_228_82 (.BL(BL82),.BLN(BLN82),.WL(WL228));
sram_cell_6t_5 inst_cell_228_83 (.BL(BL83),.BLN(BLN83),.WL(WL228));
sram_cell_6t_5 inst_cell_228_84 (.BL(BL84),.BLN(BLN84),.WL(WL228));
sram_cell_6t_5 inst_cell_228_85 (.BL(BL85),.BLN(BLN85),.WL(WL228));
sram_cell_6t_5 inst_cell_228_86 (.BL(BL86),.BLN(BLN86),.WL(WL228));
sram_cell_6t_5 inst_cell_228_87 (.BL(BL87),.BLN(BLN87),.WL(WL228));
sram_cell_6t_5 inst_cell_228_88 (.BL(BL88),.BLN(BLN88),.WL(WL228));
sram_cell_6t_5 inst_cell_228_89 (.BL(BL89),.BLN(BLN89),.WL(WL228));
sram_cell_6t_5 inst_cell_228_90 (.BL(BL90),.BLN(BLN90),.WL(WL228));
sram_cell_6t_5 inst_cell_228_91 (.BL(BL91),.BLN(BLN91),.WL(WL228));
sram_cell_6t_5 inst_cell_228_92 (.BL(BL92),.BLN(BLN92),.WL(WL228));
sram_cell_6t_5 inst_cell_228_93 (.BL(BL93),.BLN(BLN93),.WL(WL228));
sram_cell_6t_5 inst_cell_228_94 (.BL(BL94),.BLN(BLN94),.WL(WL228));
sram_cell_6t_5 inst_cell_228_95 (.BL(BL95),.BLN(BLN95),.WL(WL228));
sram_cell_6t_5 inst_cell_228_96 (.BL(BL96),.BLN(BLN96),.WL(WL228));
sram_cell_6t_5 inst_cell_228_97 (.BL(BL97),.BLN(BLN97),.WL(WL228));
sram_cell_6t_5 inst_cell_228_98 (.BL(BL98),.BLN(BLN98),.WL(WL228));
sram_cell_6t_5 inst_cell_228_99 (.BL(BL99),.BLN(BLN99),.WL(WL228));
sram_cell_6t_5 inst_cell_228_100 (.BL(BL100),.BLN(BLN100),.WL(WL228));
sram_cell_6t_5 inst_cell_228_101 (.BL(BL101),.BLN(BLN101),.WL(WL228));
sram_cell_6t_5 inst_cell_228_102 (.BL(BL102),.BLN(BLN102),.WL(WL228));
sram_cell_6t_5 inst_cell_228_103 (.BL(BL103),.BLN(BLN103),.WL(WL228));
sram_cell_6t_5 inst_cell_228_104 (.BL(BL104),.BLN(BLN104),.WL(WL228));
sram_cell_6t_5 inst_cell_228_105 (.BL(BL105),.BLN(BLN105),.WL(WL228));
sram_cell_6t_5 inst_cell_228_106 (.BL(BL106),.BLN(BLN106),.WL(WL228));
sram_cell_6t_5 inst_cell_228_107 (.BL(BL107),.BLN(BLN107),.WL(WL228));
sram_cell_6t_5 inst_cell_228_108 (.BL(BL108),.BLN(BLN108),.WL(WL228));
sram_cell_6t_5 inst_cell_228_109 (.BL(BL109),.BLN(BLN109),.WL(WL228));
sram_cell_6t_5 inst_cell_228_110 (.BL(BL110),.BLN(BLN110),.WL(WL228));
sram_cell_6t_5 inst_cell_228_111 (.BL(BL111),.BLN(BLN111),.WL(WL228));
sram_cell_6t_5 inst_cell_228_112 (.BL(BL112),.BLN(BLN112),.WL(WL228));
sram_cell_6t_5 inst_cell_228_113 (.BL(BL113),.BLN(BLN113),.WL(WL228));
sram_cell_6t_5 inst_cell_228_114 (.BL(BL114),.BLN(BLN114),.WL(WL228));
sram_cell_6t_5 inst_cell_228_115 (.BL(BL115),.BLN(BLN115),.WL(WL228));
sram_cell_6t_5 inst_cell_228_116 (.BL(BL116),.BLN(BLN116),.WL(WL228));
sram_cell_6t_5 inst_cell_228_117 (.BL(BL117),.BLN(BLN117),.WL(WL228));
sram_cell_6t_5 inst_cell_228_118 (.BL(BL118),.BLN(BLN118),.WL(WL228));
sram_cell_6t_5 inst_cell_228_119 (.BL(BL119),.BLN(BLN119),.WL(WL228));
sram_cell_6t_5 inst_cell_228_120 (.BL(BL120),.BLN(BLN120),.WL(WL228));
sram_cell_6t_5 inst_cell_228_121 (.BL(BL121),.BLN(BLN121),.WL(WL228));
sram_cell_6t_5 inst_cell_228_122 (.BL(BL122),.BLN(BLN122),.WL(WL228));
sram_cell_6t_5 inst_cell_228_123 (.BL(BL123),.BLN(BLN123),.WL(WL228));
sram_cell_6t_5 inst_cell_228_124 (.BL(BL124),.BLN(BLN124),.WL(WL228));
sram_cell_6t_5 inst_cell_228_125 (.BL(BL125),.BLN(BLN125),.WL(WL228));
sram_cell_6t_5 inst_cell_228_126 (.BL(BL126),.BLN(BLN126),.WL(WL228));
sram_cell_6t_5 inst_cell_228_127 (.BL(BL127),.BLN(BLN127),.WL(WL228));
sram_cell_6t_5 inst_cell_229_0 (.BL(BL0),.BLN(BLN0),.WL(WL229));
sram_cell_6t_5 inst_cell_229_1 (.BL(BL1),.BLN(BLN1),.WL(WL229));
sram_cell_6t_5 inst_cell_229_2 (.BL(BL2),.BLN(BLN2),.WL(WL229));
sram_cell_6t_5 inst_cell_229_3 (.BL(BL3),.BLN(BLN3),.WL(WL229));
sram_cell_6t_5 inst_cell_229_4 (.BL(BL4),.BLN(BLN4),.WL(WL229));
sram_cell_6t_5 inst_cell_229_5 (.BL(BL5),.BLN(BLN5),.WL(WL229));
sram_cell_6t_5 inst_cell_229_6 (.BL(BL6),.BLN(BLN6),.WL(WL229));
sram_cell_6t_5 inst_cell_229_7 (.BL(BL7),.BLN(BLN7),.WL(WL229));
sram_cell_6t_5 inst_cell_229_8 (.BL(BL8),.BLN(BLN8),.WL(WL229));
sram_cell_6t_5 inst_cell_229_9 (.BL(BL9),.BLN(BLN9),.WL(WL229));
sram_cell_6t_5 inst_cell_229_10 (.BL(BL10),.BLN(BLN10),.WL(WL229));
sram_cell_6t_5 inst_cell_229_11 (.BL(BL11),.BLN(BLN11),.WL(WL229));
sram_cell_6t_5 inst_cell_229_12 (.BL(BL12),.BLN(BLN12),.WL(WL229));
sram_cell_6t_5 inst_cell_229_13 (.BL(BL13),.BLN(BLN13),.WL(WL229));
sram_cell_6t_5 inst_cell_229_14 (.BL(BL14),.BLN(BLN14),.WL(WL229));
sram_cell_6t_5 inst_cell_229_15 (.BL(BL15),.BLN(BLN15),.WL(WL229));
sram_cell_6t_5 inst_cell_229_16 (.BL(BL16),.BLN(BLN16),.WL(WL229));
sram_cell_6t_5 inst_cell_229_17 (.BL(BL17),.BLN(BLN17),.WL(WL229));
sram_cell_6t_5 inst_cell_229_18 (.BL(BL18),.BLN(BLN18),.WL(WL229));
sram_cell_6t_5 inst_cell_229_19 (.BL(BL19),.BLN(BLN19),.WL(WL229));
sram_cell_6t_5 inst_cell_229_20 (.BL(BL20),.BLN(BLN20),.WL(WL229));
sram_cell_6t_5 inst_cell_229_21 (.BL(BL21),.BLN(BLN21),.WL(WL229));
sram_cell_6t_5 inst_cell_229_22 (.BL(BL22),.BLN(BLN22),.WL(WL229));
sram_cell_6t_5 inst_cell_229_23 (.BL(BL23),.BLN(BLN23),.WL(WL229));
sram_cell_6t_5 inst_cell_229_24 (.BL(BL24),.BLN(BLN24),.WL(WL229));
sram_cell_6t_5 inst_cell_229_25 (.BL(BL25),.BLN(BLN25),.WL(WL229));
sram_cell_6t_5 inst_cell_229_26 (.BL(BL26),.BLN(BLN26),.WL(WL229));
sram_cell_6t_5 inst_cell_229_27 (.BL(BL27),.BLN(BLN27),.WL(WL229));
sram_cell_6t_5 inst_cell_229_28 (.BL(BL28),.BLN(BLN28),.WL(WL229));
sram_cell_6t_5 inst_cell_229_29 (.BL(BL29),.BLN(BLN29),.WL(WL229));
sram_cell_6t_5 inst_cell_229_30 (.BL(BL30),.BLN(BLN30),.WL(WL229));
sram_cell_6t_5 inst_cell_229_31 (.BL(BL31),.BLN(BLN31),.WL(WL229));
sram_cell_6t_5 inst_cell_229_32 (.BL(BL32),.BLN(BLN32),.WL(WL229));
sram_cell_6t_5 inst_cell_229_33 (.BL(BL33),.BLN(BLN33),.WL(WL229));
sram_cell_6t_5 inst_cell_229_34 (.BL(BL34),.BLN(BLN34),.WL(WL229));
sram_cell_6t_5 inst_cell_229_35 (.BL(BL35),.BLN(BLN35),.WL(WL229));
sram_cell_6t_5 inst_cell_229_36 (.BL(BL36),.BLN(BLN36),.WL(WL229));
sram_cell_6t_5 inst_cell_229_37 (.BL(BL37),.BLN(BLN37),.WL(WL229));
sram_cell_6t_5 inst_cell_229_38 (.BL(BL38),.BLN(BLN38),.WL(WL229));
sram_cell_6t_5 inst_cell_229_39 (.BL(BL39),.BLN(BLN39),.WL(WL229));
sram_cell_6t_5 inst_cell_229_40 (.BL(BL40),.BLN(BLN40),.WL(WL229));
sram_cell_6t_5 inst_cell_229_41 (.BL(BL41),.BLN(BLN41),.WL(WL229));
sram_cell_6t_5 inst_cell_229_42 (.BL(BL42),.BLN(BLN42),.WL(WL229));
sram_cell_6t_5 inst_cell_229_43 (.BL(BL43),.BLN(BLN43),.WL(WL229));
sram_cell_6t_5 inst_cell_229_44 (.BL(BL44),.BLN(BLN44),.WL(WL229));
sram_cell_6t_5 inst_cell_229_45 (.BL(BL45),.BLN(BLN45),.WL(WL229));
sram_cell_6t_5 inst_cell_229_46 (.BL(BL46),.BLN(BLN46),.WL(WL229));
sram_cell_6t_5 inst_cell_229_47 (.BL(BL47),.BLN(BLN47),.WL(WL229));
sram_cell_6t_5 inst_cell_229_48 (.BL(BL48),.BLN(BLN48),.WL(WL229));
sram_cell_6t_5 inst_cell_229_49 (.BL(BL49),.BLN(BLN49),.WL(WL229));
sram_cell_6t_5 inst_cell_229_50 (.BL(BL50),.BLN(BLN50),.WL(WL229));
sram_cell_6t_5 inst_cell_229_51 (.BL(BL51),.BLN(BLN51),.WL(WL229));
sram_cell_6t_5 inst_cell_229_52 (.BL(BL52),.BLN(BLN52),.WL(WL229));
sram_cell_6t_5 inst_cell_229_53 (.BL(BL53),.BLN(BLN53),.WL(WL229));
sram_cell_6t_5 inst_cell_229_54 (.BL(BL54),.BLN(BLN54),.WL(WL229));
sram_cell_6t_5 inst_cell_229_55 (.BL(BL55),.BLN(BLN55),.WL(WL229));
sram_cell_6t_5 inst_cell_229_56 (.BL(BL56),.BLN(BLN56),.WL(WL229));
sram_cell_6t_5 inst_cell_229_57 (.BL(BL57),.BLN(BLN57),.WL(WL229));
sram_cell_6t_5 inst_cell_229_58 (.BL(BL58),.BLN(BLN58),.WL(WL229));
sram_cell_6t_5 inst_cell_229_59 (.BL(BL59),.BLN(BLN59),.WL(WL229));
sram_cell_6t_5 inst_cell_229_60 (.BL(BL60),.BLN(BLN60),.WL(WL229));
sram_cell_6t_5 inst_cell_229_61 (.BL(BL61),.BLN(BLN61),.WL(WL229));
sram_cell_6t_5 inst_cell_229_62 (.BL(BL62),.BLN(BLN62),.WL(WL229));
sram_cell_6t_5 inst_cell_229_63 (.BL(BL63),.BLN(BLN63),.WL(WL229));
sram_cell_6t_5 inst_cell_229_64 (.BL(BL64),.BLN(BLN64),.WL(WL229));
sram_cell_6t_5 inst_cell_229_65 (.BL(BL65),.BLN(BLN65),.WL(WL229));
sram_cell_6t_5 inst_cell_229_66 (.BL(BL66),.BLN(BLN66),.WL(WL229));
sram_cell_6t_5 inst_cell_229_67 (.BL(BL67),.BLN(BLN67),.WL(WL229));
sram_cell_6t_5 inst_cell_229_68 (.BL(BL68),.BLN(BLN68),.WL(WL229));
sram_cell_6t_5 inst_cell_229_69 (.BL(BL69),.BLN(BLN69),.WL(WL229));
sram_cell_6t_5 inst_cell_229_70 (.BL(BL70),.BLN(BLN70),.WL(WL229));
sram_cell_6t_5 inst_cell_229_71 (.BL(BL71),.BLN(BLN71),.WL(WL229));
sram_cell_6t_5 inst_cell_229_72 (.BL(BL72),.BLN(BLN72),.WL(WL229));
sram_cell_6t_5 inst_cell_229_73 (.BL(BL73),.BLN(BLN73),.WL(WL229));
sram_cell_6t_5 inst_cell_229_74 (.BL(BL74),.BLN(BLN74),.WL(WL229));
sram_cell_6t_5 inst_cell_229_75 (.BL(BL75),.BLN(BLN75),.WL(WL229));
sram_cell_6t_5 inst_cell_229_76 (.BL(BL76),.BLN(BLN76),.WL(WL229));
sram_cell_6t_5 inst_cell_229_77 (.BL(BL77),.BLN(BLN77),.WL(WL229));
sram_cell_6t_5 inst_cell_229_78 (.BL(BL78),.BLN(BLN78),.WL(WL229));
sram_cell_6t_5 inst_cell_229_79 (.BL(BL79),.BLN(BLN79),.WL(WL229));
sram_cell_6t_5 inst_cell_229_80 (.BL(BL80),.BLN(BLN80),.WL(WL229));
sram_cell_6t_5 inst_cell_229_81 (.BL(BL81),.BLN(BLN81),.WL(WL229));
sram_cell_6t_5 inst_cell_229_82 (.BL(BL82),.BLN(BLN82),.WL(WL229));
sram_cell_6t_5 inst_cell_229_83 (.BL(BL83),.BLN(BLN83),.WL(WL229));
sram_cell_6t_5 inst_cell_229_84 (.BL(BL84),.BLN(BLN84),.WL(WL229));
sram_cell_6t_5 inst_cell_229_85 (.BL(BL85),.BLN(BLN85),.WL(WL229));
sram_cell_6t_5 inst_cell_229_86 (.BL(BL86),.BLN(BLN86),.WL(WL229));
sram_cell_6t_5 inst_cell_229_87 (.BL(BL87),.BLN(BLN87),.WL(WL229));
sram_cell_6t_5 inst_cell_229_88 (.BL(BL88),.BLN(BLN88),.WL(WL229));
sram_cell_6t_5 inst_cell_229_89 (.BL(BL89),.BLN(BLN89),.WL(WL229));
sram_cell_6t_5 inst_cell_229_90 (.BL(BL90),.BLN(BLN90),.WL(WL229));
sram_cell_6t_5 inst_cell_229_91 (.BL(BL91),.BLN(BLN91),.WL(WL229));
sram_cell_6t_5 inst_cell_229_92 (.BL(BL92),.BLN(BLN92),.WL(WL229));
sram_cell_6t_5 inst_cell_229_93 (.BL(BL93),.BLN(BLN93),.WL(WL229));
sram_cell_6t_5 inst_cell_229_94 (.BL(BL94),.BLN(BLN94),.WL(WL229));
sram_cell_6t_5 inst_cell_229_95 (.BL(BL95),.BLN(BLN95),.WL(WL229));
sram_cell_6t_5 inst_cell_229_96 (.BL(BL96),.BLN(BLN96),.WL(WL229));
sram_cell_6t_5 inst_cell_229_97 (.BL(BL97),.BLN(BLN97),.WL(WL229));
sram_cell_6t_5 inst_cell_229_98 (.BL(BL98),.BLN(BLN98),.WL(WL229));
sram_cell_6t_5 inst_cell_229_99 (.BL(BL99),.BLN(BLN99),.WL(WL229));
sram_cell_6t_5 inst_cell_229_100 (.BL(BL100),.BLN(BLN100),.WL(WL229));
sram_cell_6t_5 inst_cell_229_101 (.BL(BL101),.BLN(BLN101),.WL(WL229));
sram_cell_6t_5 inst_cell_229_102 (.BL(BL102),.BLN(BLN102),.WL(WL229));
sram_cell_6t_5 inst_cell_229_103 (.BL(BL103),.BLN(BLN103),.WL(WL229));
sram_cell_6t_5 inst_cell_229_104 (.BL(BL104),.BLN(BLN104),.WL(WL229));
sram_cell_6t_5 inst_cell_229_105 (.BL(BL105),.BLN(BLN105),.WL(WL229));
sram_cell_6t_5 inst_cell_229_106 (.BL(BL106),.BLN(BLN106),.WL(WL229));
sram_cell_6t_5 inst_cell_229_107 (.BL(BL107),.BLN(BLN107),.WL(WL229));
sram_cell_6t_5 inst_cell_229_108 (.BL(BL108),.BLN(BLN108),.WL(WL229));
sram_cell_6t_5 inst_cell_229_109 (.BL(BL109),.BLN(BLN109),.WL(WL229));
sram_cell_6t_5 inst_cell_229_110 (.BL(BL110),.BLN(BLN110),.WL(WL229));
sram_cell_6t_5 inst_cell_229_111 (.BL(BL111),.BLN(BLN111),.WL(WL229));
sram_cell_6t_5 inst_cell_229_112 (.BL(BL112),.BLN(BLN112),.WL(WL229));
sram_cell_6t_5 inst_cell_229_113 (.BL(BL113),.BLN(BLN113),.WL(WL229));
sram_cell_6t_5 inst_cell_229_114 (.BL(BL114),.BLN(BLN114),.WL(WL229));
sram_cell_6t_5 inst_cell_229_115 (.BL(BL115),.BLN(BLN115),.WL(WL229));
sram_cell_6t_5 inst_cell_229_116 (.BL(BL116),.BLN(BLN116),.WL(WL229));
sram_cell_6t_5 inst_cell_229_117 (.BL(BL117),.BLN(BLN117),.WL(WL229));
sram_cell_6t_5 inst_cell_229_118 (.BL(BL118),.BLN(BLN118),.WL(WL229));
sram_cell_6t_5 inst_cell_229_119 (.BL(BL119),.BLN(BLN119),.WL(WL229));
sram_cell_6t_5 inst_cell_229_120 (.BL(BL120),.BLN(BLN120),.WL(WL229));
sram_cell_6t_5 inst_cell_229_121 (.BL(BL121),.BLN(BLN121),.WL(WL229));
sram_cell_6t_5 inst_cell_229_122 (.BL(BL122),.BLN(BLN122),.WL(WL229));
sram_cell_6t_5 inst_cell_229_123 (.BL(BL123),.BLN(BLN123),.WL(WL229));
sram_cell_6t_5 inst_cell_229_124 (.BL(BL124),.BLN(BLN124),.WL(WL229));
sram_cell_6t_5 inst_cell_229_125 (.BL(BL125),.BLN(BLN125),.WL(WL229));
sram_cell_6t_5 inst_cell_229_126 (.BL(BL126),.BLN(BLN126),.WL(WL229));
sram_cell_6t_5 inst_cell_229_127 (.BL(BL127),.BLN(BLN127),.WL(WL229));
sram_cell_6t_5 inst_cell_230_0 (.BL(BL0),.BLN(BLN0),.WL(WL230));
sram_cell_6t_5 inst_cell_230_1 (.BL(BL1),.BLN(BLN1),.WL(WL230));
sram_cell_6t_5 inst_cell_230_2 (.BL(BL2),.BLN(BLN2),.WL(WL230));
sram_cell_6t_5 inst_cell_230_3 (.BL(BL3),.BLN(BLN3),.WL(WL230));
sram_cell_6t_5 inst_cell_230_4 (.BL(BL4),.BLN(BLN4),.WL(WL230));
sram_cell_6t_5 inst_cell_230_5 (.BL(BL5),.BLN(BLN5),.WL(WL230));
sram_cell_6t_5 inst_cell_230_6 (.BL(BL6),.BLN(BLN6),.WL(WL230));
sram_cell_6t_5 inst_cell_230_7 (.BL(BL7),.BLN(BLN7),.WL(WL230));
sram_cell_6t_5 inst_cell_230_8 (.BL(BL8),.BLN(BLN8),.WL(WL230));
sram_cell_6t_5 inst_cell_230_9 (.BL(BL9),.BLN(BLN9),.WL(WL230));
sram_cell_6t_5 inst_cell_230_10 (.BL(BL10),.BLN(BLN10),.WL(WL230));
sram_cell_6t_5 inst_cell_230_11 (.BL(BL11),.BLN(BLN11),.WL(WL230));
sram_cell_6t_5 inst_cell_230_12 (.BL(BL12),.BLN(BLN12),.WL(WL230));
sram_cell_6t_5 inst_cell_230_13 (.BL(BL13),.BLN(BLN13),.WL(WL230));
sram_cell_6t_5 inst_cell_230_14 (.BL(BL14),.BLN(BLN14),.WL(WL230));
sram_cell_6t_5 inst_cell_230_15 (.BL(BL15),.BLN(BLN15),.WL(WL230));
sram_cell_6t_5 inst_cell_230_16 (.BL(BL16),.BLN(BLN16),.WL(WL230));
sram_cell_6t_5 inst_cell_230_17 (.BL(BL17),.BLN(BLN17),.WL(WL230));
sram_cell_6t_5 inst_cell_230_18 (.BL(BL18),.BLN(BLN18),.WL(WL230));
sram_cell_6t_5 inst_cell_230_19 (.BL(BL19),.BLN(BLN19),.WL(WL230));
sram_cell_6t_5 inst_cell_230_20 (.BL(BL20),.BLN(BLN20),.WL(WL230));
sram_cell_6t_5 inst_cell_230_21 (.BL(BL21),.BLN(BLN21),.WL(WL230));
sram_cell_6t_5 inst_cell_230_22 (.BL(BL22),.BLN(BLN22),.WL(WL230));
sram_cell_6t_5 inst_cell_230_23 (.BL(BL23),.BLN(BLN23),.WL(WL230));
sram_cell_6t_5 inst_cell_230_24 (.BL(BL24),.BLN(BLN24),.WL(WL230));
sram_cell_6t_5 inst_cell_230_25 (.BL(BL25),.BLN(BLN25),.WL(WL230));
sram_cell_6t_5 inst_cell_230_26 (.BL(BL26),.BLN(BLN26),.WL(WL230));
sram_cell_6t_5 inst_cell_230_27 (.BL(BL27),.BLN(BLN27),.WL(WL230));
sram_cell_6t_5 inst_cell_230_28 (.BL(BL28),.BLN(BLN28),.WL(WL230));
sram_cell_6t_5 inst_cell_230_29 (.BL(BL29),.BLN(BLN29),.WL(WL230));
sram_cell_6t_5 inst_cell_230_30 (.BL(BL30),.BLN(BLN30),.WL(WL230));
sram_cell_6t_5 inst_cell_230_31 (.BL(BL31),.BLN(BLN31),.WL(WL230));
sram_cell_6t_5 inst_cell_230_32 (.BL(BL32),.BLN(BLN32),.WL(WL230));
sram_cell_6t_5 inst_cell_230_33 (.BL(BL33),.BLN(BLN33),.WL(WL230));
sram_cell_6t_5 inst_cell_230_34 (.BL(BL34),.BLN(BLN34),.WL(WL230));
sram_cell_6t_5 inst_cell_230_35 (.BL(BL35),.BLN(BLN35),.WL(WL230));
sram_cell_6t_5 inst_cell_230_36 (.BL(BL36),.BLN(BLN36),.WL(WL230));
sram_cell_6t_5 inst_cell_230_37 (.BL(BL37),.BLN(BLN37),.WL(WL230));
sram_cell_6t_5 inst_cell_230_38 (.BL(BL38),.BLN(BLN38),.WL(WL230));
sram_cell_6t_5 inst_cell_230_39 (.BL(BL39),.BLN(BLN39),.WL(WL230));
sram_cell_6t_5 inst_cell_230_40 (.BL(BL40),.BLN(BLN40),.WL(WL230));
sram_cell_6t_5 inst_cell_230_41 (.BL(BL41),.BLN(BLN41),.WL(WL230));
sram_cell_6t_5 inst_cell_230_42 (.BL(BL42),.BLN(BLN42),.WL(WL230));
sram_cell_6t_5 inst_cell_230_43 (.BL(BL43),.BLN(BLN43),.WL(WL230));
sram_cell_6t_5 inst_cell_230_44 (.BL(BL44),.BLN(BLN44),.WL(WL230));
sram_cell_6t_5 inst_cell_230_45 (.BL(BL45),.BLN(BLN45),.WL(WL230));
sram_cell_6t_5 inst_cell_230_46 (.BL(BL46),.BLN(BLN46),.WL(WL230));
sram_cell_6t_5 inst_cell_230_47 (.BL(BL47),.BLN(BLN47),.WL(WL230));
sram_cell_6t_5 inst_cell_230_48 (.BL(BL48),.BLN(BLN48),.WL(WL230));
sram_cell_6t_5 inst_cell_230_49 (.BL(BL49),.BLN(BLN49),.WL(WL230));
sram_cell_6t_5 inst_cell_230_50 (.BL(BL50),.BLN(BLN50),.WL(WL230));
sram_cell_6t_5 inst_cell_230_51 (.BL(BL51),.BLN(BLN51),.WL(WL230));
sram_cell_6t_5 inst_cell_230_52 (.BL(BL52),.BLN(BLN52),.WL(WL230));
sram_cell_6t_5 inst_cell_230_53 (.BL(BL53),.BLN(BLN53),.WL(WL230));
sram_cell_6t_5 inst_cell_230_54 (.BL(BL54),.BLN(BLN54),.WL(WL230));
sram_cell_6t_5 inst_cell_230_55 (.BL(BL55),.BLN(BLN55),.WL(WL230));
sram_cell_6t_5 inst_cell_230_56 (.BL(BL56),.BLN(BLN56),.WL(WL230));
sram_cell_6t_5 inst_cell_230_57 (.BL(BL57),.BLN(BLN57),.WL(WL230));
sram_cell_6t_5 inst_cell_230_58 (.BL(BL58),.BLN(BLN58),.WL(WL230));
sram_cell_6t_5 inst_cell_230_59 (.BL(BL59),.BLN(BLN59),.WL(WL230));
sram_cell_6t_5 inst_cell_230_60 (.BL(BL60),.BLN(BLN60),.WL(WL230));
sram_cell_6t_5 inst_cell_230_61 (.BL(BL61),.BLN(BLN61),.WL(WL230));
sram_cell_6t_5 inst_cell_230_62 (.BL(BL62),.BLN(BLN62),.WL(WL230));
sram_cell_6t_5 inst_cell_230_63 (.BL(BL63),.BLN(BLN63),.WL(WL230));
sram_cell_6t_5 inst_cell_230_64 (.BL(BL64),.BLN(BLN64),.WL(WL230));
sram_cell_6t_5 inst_cell_230_65 (.BL(BL65),.BLN(BLN65),.WL(WL230));
sram_cell_6t_5 inst_cell_230_66 (.BL(BL66),.BLN(BLN66),.WL(WL230));
sram_cell_6t_5 inst_cell_230_67 (.BL(BL67),.BLN(BLN67),.WL(WL230));
sram_cell_6t_5 inst_cell_230_68 (.BL(BL68),.BLN(BLN68),.WL(WL230));
sram_cell_6t_5 inst_cell_230_69 (.BL(BL69),.BLN(BLN69),.WL(WL230));
sram_cell_6t_5 inst_cell_230_70 (.BL(BL70),.BLN(BLN70),.WL(WL230));
sram_cell_6t_5 inst_cell_230_71 (.BL(BL71),.BLN(BLN71),.WL(WL230));
sram_cell_6t_5 inst_cell_230_72 (.BL(BL72),.BLN(BLN72),.WL(WL230));
sram_cell_6t_5 inst_cell_230_73 (.BL(BL73),.BLN(BLN73),.WL(WL230));
sram_cell_6t_5 inst_cell_230_74 (.BL(BL74),.BLN(BLN74),.WL(WL230));
sram_cell_6t_5 inst_cell_230_75 (.BL(BL75),.BLN(BLN75),.WL(WL230));
sram_cell_6t_5 inst_cell_230_76 (.BL(BL76),.BLN(BLN76),.WL(WL230));
sram_cell_6t_5 inst_cell_230_77 (.BL(BL77),.BLN(BLN77),.WL(WL230));
sram_cell_6t_5 inst_cell_230_78 (.BL(BL78),.BLN(BLN78),.WL(WL230));
sram_cell_6t_5 inst_cell_230_79 (.BL(BL79),.BLN(BLN79),.WL(WL230));
sram_cell_6t_5 inst_cell_230_80 (.BL(BL80),.BLN(BLN80),.WL(WL230));
sram_cell_6t_5 inst_cell_230_81 (.BL(BL81),.BLN(BLN81),.WL(WL230));
sram_cell_6t_5 inst_cell_230_82 (.BL(BL82),.BLN(BLN82),.WL(WL230));
sram_cell_6t_5 inst_cell_230_83 (.BL(BL83),.BLN(BLN83),.WL(WL230));
sram_cell_6t_5 inst_cell_230_84 (.BL(BL84),.BLN(BLN84),.WL(WL230));
sram_cell_6t_5 inst_cell_230_85 (.BL(BL85),.BLN(BLN85),.WL(WL230));
sram_cell_6t_5 inst_cell_230_86 (.BL(BL86),.BLN(BLN86),.WL(WL230));
sram_cell_6t_5 inst_cell_230_87 (.BL(BL87),.BLN(BLN87),.WL(WL230));
sram_cell_6t_5 inst_cell_230_88 (.BL(BL88),.BLN(BLN88),.WL(WL230));
sram_cell_6t_5 inst_cell_230_89 (.BL(BL89),.BLN(BLN89),.WL(WL230));
sram_cell_6t_5 inst_cell_230_90 (.BL(BL90),.BLN(BLN90),.WL(WL230));
sram_cell_6t_5 inst_cell_230_91 (.BL(BL91),.BLN(BLN91),.WL(WL230));
sram_cell_6t_5 inst_cell_230_92 (.BL(BL92),.BLN(BLN92),.WL(WL230));
sram_cell_6t_5 inst_cell_230_93 (.BL(BL93),.BLN(BLN93),.WL(WL230));
sram_cell_6t_5 inst_cell_230_94 (.BL(BL94),.BLN(BLN94),.WL(WL230));
sram_cell_6t_5 inst_cell_230_95 (.BL(BL95),.BLN(BLN95),.WL(WL230));
sram_cell_6t_5 inst_cell_230_96 (.BL(BL96),.BLN(BLN96),.WL(WL230));
sram_cell_6t_5 inst_cell_230_97 (.BL(BL97),.BLN(BLN97),.WL(WL230));
sram_cell_6t_5 inst_cell_230_98 (.BL(BL98),.BLN(BLN98),.WL(WL230));
sram_cell_6t_5 inst_cell_230_99 (.BL(BL99),.BLN(BLN99),.WL(WL230));
sram_cell_6t_5 inst_cell_230_100 (.BL(BL100),.BLN(BLN100),.WL(WL230));
sram_cell_6t_5 inst_cell_230_101 (.BL(BL101),.BLN(BLN101),.WL(WL230));
sram_cell_6t_5 inst_cell_230_102 (.BL(BL102),.BLN(BLN102),.WL(WL230));
sram_cell_6t_5 inst_cell_230_103 (.BL(BL103),.BLN(BLN103),.WL(WL230));
sram_cell_6t_5 inst_cell_230_104 (.BL(BL104),.BLN(BLN104),.WL(WL230));
sram_cell_6t_5 inst_cell_230_105 (.BL(BL105),.BLN(BLN105),.WL(WL230));
sram_cell_6t_5 inst_cell_230_106 (.BL(BL106),.BLN(BLN106),.WL(WL230));
sram_cell_6t_5 inst_cell_230_107 (.BL(BL107),.BLN(BLN107),.WL(WL230));
sram_cell_6t_5 inst_cell_230_108 (.BL(BL108),.BLN(BLN108),.WL(WL230));
sram_cell_6t_5 inst_cell_230_109 (.BL(BL109),.BLN(BLN109),.WL(WL230));
sram_cell_6t_5 inst_cell_230_110 (.BL(BL110),.BLN(BLN110),.WL(WL230));
sram_cell_6t_5 inst_cell_230_111 (.BL(BL111),.BLN(BLN111),.WL(WL230));
sram_cell_6t_5 inst_cell_230_112 (.BL(BL112),.BLN(BLN112),.WL(WL230));
sram_cell_6t_5 inst_cell_230_113 (.BL(BL113),.BLN(BLN113),.WL(WL230));
sram_cell_6t_5 inst_cell_230_114 (.BL(BL114),.BLN(BLN114),.WL(WL230));
sram_cell_6t_5 inst_cell_230_115 (.BL(BL115),.BLN(BLN115),.WL(WL230));
sram_cell_6t_5 inst_cell_230_116 (.BL(BL116),.BLN(BLN116),.WL(WL230));
sram_cell_6t_5 inst_cell_230_117 (.BL(BL117),.BLN(BLN117),.WL(WL230));
sram_cell_6t_5 inst_cell_230_118 (.BL(BL118),.BLN(BLN118),.WL(WL230));
sram_cell_6t_5 inst_cell_230_119 (.BL(BL119),.BLN(BLN119),.WL(WL230));
sram_cell_6t_5 inst_cell_230_120 (.BL(BL120),.BLN(BLN120),.WL(WL230));
sram_cell_6t_5 inst_cell_230_121 (.BL(BL121),.BLN(BLN121),.WL(WL230));
sram_cell_6t_5 inst_cell_230_122 (.BL(BL122),.BLN(BLN122),.WL(WL230));
sram_cell_6t_5 inst_cell_230_123 (.BL(BL123),.BLN(BLN123),.WL(WL230));
sram_cell_6t_5 inst_cell_230_124 (.BL(BL124),.BLN(BLN124),.WL(WL230));
sram_cell_6t_5 inst_cell_230_125 (.BL(BL125),.BLN(BLN125),.WL(WL230));
sram_cell_6t_5 inst_cell_230_126 (.BL(BL126),.BLN(BLN126),.WL(WL230));
sram_cell_6t_5 inst_cell_230_127 (.BL(BL127),.BLN(BLN127),.WL(WL230));
sram_cell_6t_5 inst_cell_231_0 (.BL(BL0),.BLN(BLN0),.WL(WL231));
sram_cell_6t_5 inst_cell_231_1 (.BL(BL1),.BLN(BLN1),.WL(WL231));
sram_cell_6t_5 inst_cell_231_2 (.BL(BL2),.BLN(BLN2),.WL(WL231));
sram_cell_6t_5 inst_cell_231_3 (.BL(BL3),.BLN(BLN3),.WL(WL231));
sram_cell_6t_5 inst_cell_231_4 (.BL(BL4),.BLN(BLN4),.WL(WL231));
sram_cell_6t_5 inst_cell_231_5 (.BL(BL5),.BLN(BLN5),.WL(WL231));
sram_cell_6t_5 inst_cell_231_6 (.BL(BL6),.BLN(BLN6),.WL(WL231));
sram_cell_6t_5 inst_cell_231_7 (.BL(BL7),.BLN(BLN7),.WL(WL231));
sram_cell_6t_5 inst_cell_231_8 (.BL(BL8),.BLN(BLN8),.WL(WL231));
sram_cell_6t_5 inst_cell_231_9 (.BL(BL9),.BLN(BLN9),.WL(WL231));
sram_cell_6t_5 inst_cell_231_10 (.BL(BL10),.BLN(BLN10),.WL(WL231));
sram_cell_6t_5 inst_cell_231_11 (.BL(BL11),.BLN(BLN11),.WL(WL231));
sram_cell_6t_5 inst_cell_231_12 (.BL(BL12),.BLN(BLN12),.WL(WL231));
sram_cell_6t_5 inst_cell_231_13 (.BL(BL13),.BLN(BLN13),.WL(WL231));
sram_cell_6t_5 inst_cell_231_14 (.BL(BL14),.BLN(BLN14),.WL(WL231));
sram_cell_6t_5 inst_cell_231_15 (.BL(BL15),.BLN(BLN15),.WL(WL231));
sram_cell_6t_5 inst_cell_231_16 (.BL(BL16),.BLN(BLN16),.WL(WL231));
sram_cell_6t_5 inst_cell_231_17 (.BL(BL17),.BLN(BLN17),.WL(WL231));
sram_cell_6t_5 inst_cell_231_18 (.BL(BL18),.BLN(BLN18),.WL(WL231));
sram_cell_6t_5 inst_cell_231_19 (.BL(BL19),.BLN(BLN19),.WL(WL231));
sram_cell_6t_5 inst_cell_231_20 (.BL(BL20),.BLN(BLN20),.WL(WL231));
sram_cell_6t_5 inst_cell_231_21 (.BL(BL21),.BLN(BLN21),.WL(WL231));
sram_cell_6t_5 inst_cell_231_22 (.BL(BL22),.BLN(BLN22),.WL(WL231));
sram_cell_6t_5 inst_cell_231_23 (.BL(BL23),.BLN(BLN23),.WL(WL231));
sram_cell_6t_5 inst_cell_231_24 (.BL(BL24),.BLN(BLN24),.WL(WL231));
sram_cell_6t_5 inst_cell_231_25 (.BL(BL25),.BLN(BLN25),.WL(WL231));
sram_cell_6t_5 inst_cell_231_26 (.BL(BL26),.BLN(BLN26),.WL(WL231));
sram_cell_6t_5 inst_cell_231_27 (.BL(BL27),.BLN(BLN27),.WL(WL231));
sram_cell_6t_5 inst_cell_231_28 (.BL(BL28),.BLN(BLN28),.WL(WL231));
sram_cell_6t_5 inst_cell_231_29 (.BL(BL29),.BLN(BLN29),.WL(WL231));
sram_cell_6t_5 inst_cell_231_30 (.BL(BL30),.BLN(BLN30),.WL(WL231));
sram_cell_6t_5 inst_cell_231_31 (.BL(BL31),.BLN(BLN31),.WL(WL231));
sram_cell_6t_5 inst_cell_231_32 (.BL(BL32),.BLN(BLN32),.WL(WL231));
sram_cell_6t_5 inst_cell_231_33 (.BL(BL33),.BLN(BLN33),.WL(WL231));
sram_cell_6t_5 inst_cell_231_34 (.BL(BL34),.BLN(BLN34),.WL(WL231));
sram_cell_6t_5 inst_cell_231_35 (.BL(BL35),.BLN(BLN35),.WL(WL231));
sram_cell_6t_5 inst_cell_231_36 (.BL(BL36),.BLN(BLN36),.WL(WL231));
sram_cell_6t_5 inst_cell_231_37 (.BL(BL37),.BLN(BLN37),.WL(WL231));
sram_cell_6t_5 inst_cell_231_38 (.BL(BL38),.BLN(BLN38),.WL(WL231));
sram_cell_6t_5 inst_cell_231_39 (.BL(BL39),.BLN(BLN39),.WL(WL231));
sram_cell_6t_5 inst_cell_231_40 (.BL(BL40),.BLN(BLN40),.WL(WL231));
sram_cell_6t_5 inst_cell_231_41 (.BL(BL41),.BLN(BLN41),.WL(WL231));
sram_cell_6t_5 inst_cell_231_42 (.BL(BL42),.BLN(BLN42),.WL(WL231));
sram_cell_6t_5 inst_cell_231_43 (.BL(BL43),.BLN(BLN43),.WL(WL231));
sram_cell_6t_5 inst_cell_231_44 (.BL(BL44),.BLN(BLN44),.WL(WL231));
sram_cell_6t_5 inst_cell_231_45 (.BL(BL45),.BLN(BLN45),.WL(WL231));
sram_cell_6t_5 inst_cell_231_46 (.BL(BL46),.BLN(BLN46),.WL(WL231));
sram_cell_6t_5 inst_cell_231_47 (.BL(BL47),.BLN(BLN47),.WL(WL231));
sram_cell_6t_5 inst_cell_231_48 (.BL(BL48),.BLN(BLN48),.WL(WL231));
sram_cell_6t_5 inst_cell_231_49 (.BL(BL49),.BLN(BLN49),.WL(WL231));
sram_cell_6t_5 inst_cell_231_50 (.BL(BL50),.BLN(BLN50),.WL(WL231));
sram_cell_6t_5 inst_cell_231_51 (.BL(BL51),.BLN(BLN51),.WL(WL231));
sram_cell_6t_5 inst_cell_231_52 (.BL(BL52),.BLN(BLN52),.WL(WL231));
sram_cell_6t_5 inst_cell_231_53 (.BL(BL53),.BLN(BLN53),.WL(WL231));
sram_cell_6t_5 inst_cell_231_54 (.BL(BL54),.BLN(BLN54),.WL(WL231));
sram_cell_6t_5 inst_cell_231_55 (.BL(BL55),.BLN(BLN55),.WL(WL231));
sram_cell_6t_5 inst_cell_231_56 (.BL(BL56),.BLN(BLN56),.WL(WL231));
sram_cell_6t_5 inst_cell_231_57 (.BL(BL57),.BLN(BLN57),.WL(WL231));
sram_cell_6t_5 inst_cell_231_58 (.BL(BL58),.BLN(BLN58),.WL(WL231));
sram_cell_6t_5 inst_cell_231_59 (.BL(BL59),.BLN(BLN59),.WL(WL231));
sram_cell_6t_5 inst_cell_231_60 (.BL(BL60),.BLN(BLN60),.WL(WL231));
sram_cell_6t_5 inst_cell_231_61 (.BL(BL61),.BLN(BLN61),.WL(WL231));
sram_cell_6t_5 inst_cell_231_62 (.BL(BL62),.BLN(BLN62),.WL(WL231));
sram_cell_6t_5 inst_cell_231_63 (.BL(BL63),.BLN(BLN63),.WL(WL231));
sram_cell_6t_5 inst_cell_231_64 (.BL(BL64),.BLN(BLN64),.WL(WL231));
sram_cell_6t_5 inst_cell_231_65 (.BL(BL65),.BLN(BLN65),.WL(WL231));
sram_cell_6t_5 inst_cell_231_66 (.BL(BL66),.BLN(BLN66),.WL(WL231));
sram_cell_6t_5 inst_cell_231_67 (.BL(BL67),.BLN(BLN67),.WL(WL231));
sram_cell_6t_5 inst_cell_231_68 (.BL(BL68),.BLN(BLN68),.WL(WL231));
sram_cell_6t_5 inst_cell_231_69 (.BL(BL69),.BLN(BLN69),.WL(WL231));
sram_cell_6t_5 inst_cell_231_70 (.BL(BL70),.BLN(BLN70),.WL(WL231));
sram_cell_6t_5 inst_cell_231_71 (.BL(BL71),.BLN(BLN71),.WL(WL231));
sram_cell_6t_5 inst_cell_231_72 (.BL(BL72),.BLN(BLN72),.WL(WL231));
sram_cell_6t_5 inst_cell_231_73 (.BL(BL73),.BLN(BLN73),.WL(WL231));
sram_cell_6t_5 inst_cell_231_74 (.BL(BL74),.BLN(BLN74),.WL(WL231));
sram_cell_6t_5 inst_cell_231_75 (.BL(BL75),.BLN(BLN75),.WL(WL231));
sram_cell_6t_5 inst_cell_231_76 (.BL(BL76),.BLN(BLN76),.WL(WL231));
sram_cell_6t_5 inst_cell_231_77 (.BL(BL77),.BLN(BLN77),.WL(WL231));
sram_cell_6t_5 inst_cell_231_78 (.BL(BL78),.BLN(BLN78),.WL(WL231));
sram_cell_6t_5 inst_cell_231_79 (.BL(BL79),.BLN(BLN79),.WL(WL231));
sram_cell_6t_5 inst_cell_231_80 (.BL(BL80),.BLN(BLN80),.WL(WL231));
sram_cell_6t_5 inst_cell_231_81 (.BL(BL81),.BLN(BLN81),.WL(WL231));
sram_cell_6t_5 inst_cell_231_82 (.BL(BL82),.BLN(BLN82),.WL(WL231));
sram_cell_6t_5 inst_cell_231_83 (.BL(BL83),.BLN(BLN83),.WL(WL231));
sram_cell_6t_5 inst_cell_231_84 (.BL(BL84),.BLN(BLN84),.WL(WL231));
sram_cell_6t_5 inst_cell_231_85 (.BL(BL85),.BLN(BLN85),.WL(WL231));
sram_cell_6t_5 inst_cell_231_86 (.BL(BL86),.BLN(BLN86),.WL(WL231));
sram_cell_6t_5 inst_cell_231_87 (.BL(BL87),.BLN(BLN87),.WL(WL231));
sram_cell_6t_5 inst_cell_231_88 (.BL(BL88),.BLN(BLN88),.WL(WL231));
sram_cell_6t_5 inst_cell_231_89 (.BL(BL89),.BLN(BLN89),.WL(WL231));
sram_cell_6t_5 inst_cell_231_90 (.BL(BL90),.BLN(BLN90),.WL(WL231));
sram_cell_6t_5 inst_cell_231_91 (.BL(BL91),.BLN(BLN91),.WL(WL231));
sram_cell_6t_5 inst_cell_231_92 (.BL(BL92),.BLN(BLN92),.WL(WL231));
sram_cell_6t_5 inst_cell_231_93 (.BL(BL93),.BLN(BLN93),.WL(WL231));
sram_cell_6t_5 inst_cell_231_94 (.BL(BL94),.BLN(BLN94),.WL(WL231));
sram_cell_6t_5 inst_cell_231_95 (.BL(BL95),.BLN(BLN95),.WL(WL231));
sram_cell_6t_5 inst_cell_231_96 (.BL(BL96),.BLN(BLN96),.WL(WL231));
sram_cell_6t_5 inst_cell_231_97 (.BL(BL97),.BLN(BLN97),.WL(WL231));
sram_cell_6t_5 inst_cell_231_98 (.BL(BL98),.BLN(BLN98),.WL(WL231));
sram_cell_6t_5 inst_cell_231_99 (.BL(BL99),.BLN(BLN99),.WL(WL231));
sram_cell_6t_5 inst_cell_231_100 (.BL(BL100),.BLN(BLN100),.WL(WL231));
sram_cell_6t_5 inst_cell_231_101 (.BL(BL101),.BLN(BLN101),.WL(WL231));
sram_cell_6t_5 inst_cell_231_102 (.BL(BL102),.BLN(BLN102),.WL(WL231));
sram_cell_6t_5 inst_cell_231_103 (.BL(BL103),.BLN(BLN103),.WL(WL231));
sram_cell_6t_5 inst_cell_231_104 (.BL(BL104),.BLN(BLN104),.WL(WL231));
sram_cell_6t_5 inst_cell_231_105 (.BL(BL105),.BLN(BLN105),.WL(WL231));
sram_cell_6t_5 inst_cell_231_106 (.BL(BL106),.BLN(BLN106),.WL(WL231));
sram_cell_6t_5 inst_cell_231_107 (.BL(BL107),.BLN(BLN107),.WL(WL231));
sram_cell_6t_5 inst_cell_231_108 (.BL(BL108),.BLN(BLN108),.WL(WL231));
sram_cell_6t_5 inst_cell_231_109 (.BL(BL109),.BLN(BLN109),.WL(WL231));
sram_cell_6t_5 inst_cell_231_110 (.BL(BL110),.BLN(BLN110),.WL(WL231));
sram_cell_6t_5 inst_cell_231_111 (.BL(BL111),.BLN(BLN111),.WL(WL231));
sram_cell_6t_5 inst_cell_231_112 (.BL(BL112),.BLN(BLN112),.WL(WL231));
sram_cell_6t_5 inst_cell_231_113 (.BL(BL113),.BLN(BLN113),.WL(WL231));
sram_cell_6t_5 inst_cell_231_114 (.BL(BL114),.BLN(BLN114),.WL(WL231));
sram_cell_6t_5 inst_cell_231_115 (.BL(BL115),.BLN(BLN115),.WL(WL231));
sram_cell_6t_5 inst_cell_231_116 (.BL(BL116),.BLN(BLN116),.WL(WL231));
sram_cell_6t_5 inst_cell_231_117 (.BL(BL117),.BLN(BLN117),.WL(WL231));
sram_cell_6t_5 inst_cell_231_118 (.BL(BL118),.BLN(BLN118),.WL(WL231));
sram_cell_6t_5 inst_cell_231_119 (.BL(BL119),.BLN(BLN119),.WL(WL231));
sram_cell_6t_5 inst_cell_231_120 (.BL(BL120),.BLN(BLN120),.WL(WL231));
sram_cell_6t_5 inst_cell_231_121 (.BL(BL121),.BLN(BLN121),.WL(WL231));
sram_cell_6t_5 inst_cell_231_122 (.BL(BL122),.BLN(BLN122),.WL(WL231));
sram_cell_6t_5 inst_cell_231_123 (.BL(BL123),.BLN(BLN123),.WL(WL231));
sram_cell_6t_5 inst_cell_231_124 (.BL(BL124),.BLN(BLN124),.WL(WL231));
sram_cell_6t_5 inst_cell_231_125 (.BL(BL125),.BLN(BLN125),.WL(WL231));
sram_cell_6t_5 inst_cell_231_126 (.BL(BL126),.BLN(BLN126),.WL(WL231));
sram_cell_6t_5 inst_cell_231_127 (.BL(BL127),.BLN(BLN127),.WL(WL231));
sram_cell_6t_5 inst_cell_232_0 (.BL(BL0),.BLN(BLN0),.WL(WL232));
sram_cell_6t_5 inst_cell_232_1 (.BL(BL1),.BLN(BLN1),.WL(WL232));
sram_cell_6t_5 inst_cell_232_2 (.BL(BL2),.BLN(BLN2),.WL(WL232));
sram_cell_6t_5 inst_cell_232_3 (.BL(BL3),.BLN(BLN3),.WL(WL232));
sram_cell_6t_5 inst_cell_232_4 (.BL(BL4),.BLN(BLN4),.WL(WL232));
sram_cell_6t_5 inst_cell_232_5 (.BL(BL5),.BLN(BLN5),.WL(WL232));
sram_cell_6t_5 inst_cell_232_6 (.BL(BL6),.BLN(BLN6),.WL(WL232));
sram_cell_6t_5 inst_cell_232_7 (.BL(BL7),.BLN(BLN7),.WL(WL232));
sram_cell_6t_5 inst_cell_232_8 (.BL(BL8),.BLN(BLN8),.WL(WL232));
sram_cell_6t_5 inst_cell_232_9 (.BL(BL9),.BLN(BLN9),.WL(WL232));
sram_cell_6t_5 inst_cell_232_10 (.BL(BL10),.BLN(BLN10),.WL(WL232));
sram_cell_6t_5 inst_cell_232_11 (.BL(BL11),.BLN(BLN11),.WL(WL232));
sram_cell_6t_5 inst_cell_232_12 (.BL(BL12),.BLN(BLN12),.WL(WL232));
sram_cell_6t_5 inst_cell_232_13 (.BL(BL13),.BLN(BLN13),.WL(WL232));
sram_cell_6t_5 inst_cell_232_14 (.BL(BL14),.BLN(BLN14),.WL(WL232));
sram_cell_6t_5 inst_cell_232_15 (.BL(BL15),.BLN(BLN15),.WL(WL232));
sram_cell_6t_5 inst_cell_232_16 (.BL(BL16),.BLN(BLN16),.WL(WL232));
sram_cell_6t_5 inst_cell_232_17 (.BL(BL17),.BLN(BLN17),.WL(WL232));
sram_cell_6t_5 inst_cell_232_18 (.BL(BL18),.BLN(BLN18),.WL(WL232));
sram_cell_6t_5 inst_cell_232_19 (.BL(BL19),.BLN(BLN19),.WL(WL232));
sram_cell_6t_5 inst_cell_232_20 (.BL(BL20),.BLN(BLN20),.WL(WL232));
sram_cell_6t_5 inst_cell_232_21 (.BL(BL21),.BLN(BLN21),.WL(WL232));
sram_cell_6t_5 inst_cell_232_22 (.BL(BL22),.BLN(BLN22),.WL(WL232));
sram_cell_6t_5 inst_cell_232_23 (.BL(BL23),.BLN(BLN23),.WL(WL232));
sram_cell_6t_5 inst_cell_232_24 (.BL(BL24),.BLN(BLN24),.WL(WL232));
sram_cell_6t_5 inst_cell_232_25 (.BL(BL25),.BLN(BLN25),.WL(WL232));
sram_cell_6t_5 inst_cell_232_26 (.BL(BL26),.BLN(BLN26),.WL(WL232));
sram_cell_6t_5 inst_cell_232_27 (.BL(BL27),.BLN(BLN27),.WL(WL232));
sram_cell_6t_5 inst_cell_232_28 (.BL(BL28),.BLN(BLN28),.WL(WL232));
sram_cell_6t_5 inst_cell_232_29 (.BL(BL29),.BLN(BLN29),.WL(WL232));
sram_cell_6t_5 inst_cell_232_30 (.BL(BL30),.BLN(BLN30),.WL(WL232));
sram_cell_6t_5 inst_cell_232_31 (.BL(BL31),.BLN(BLN31),.WL(WL232));
sram_cell_6t_5 inst_cell_232_32 (.BL(BL32),.BLN(BLN32),.WL(WL232));
sram_cell_6t_5 inst_cell_232_33 (.BL(BL33),.BLN(BLN33),.WL(WL232));
sram_cell_6t_5 inst_cell_232_34 (.BL(BL34),.BLN(BLN34),.WL(WL232));
sram_cell_6t_5 inst_cell_232_35 (.BL(BL35),.BLN(BLN35),.WL(WL232));
sram_cell_6t_5 inst_cell_232_36 (.BL(BL36),.BLN(BLN36),.WL(WL232));
sram_cell_6t_5 inst_cell_232_37 (.BL(BL37),.BLN(BLN37),.WL(WL232));
sram_cell_6t_5 inst_cell_232_38 (.BL(BL38),.BLN(BLN38),.WL(WL232));
sram_cell_6t_5 inst_cell_232_39 (.BL(BL39),.BLN(BLN39),.WL(WL232));
sram_cell_6t_5 inst_cell_232_40 (.BL(BL40),.BLN(BLN40),.WL(WL232));
sram_cell_6t_5 inst_cell_232_41 (.BL(BL41),.BLN(BLN41),.WL(WL232));
sram_cell_6t_5 inst_cell_232_42 (.BL(BL42),.BLN(BLN42),.WL(WL232));
sram_cell_6t_5 inst_cell_232_43 (.BL(BL43),.BLN(BLN43),.WL(WL232));
sram_cell_6t_5 inst_cell_232_44 (.BL(BL44),.BLN(BLN44),.WL(WL232));
sram_cell_6t_5 inst_cell_232_45 (.BL(BL45),.BLN(BLN45),.WL(WL232));
sram_cell_6t_5 inst_cell_232_46 (.BL(BL46),.BLN(BLN46),.WL(WL232));
sram_cell_6t_5 inst_cell_232_47 (.BL(BL47),.BLN(BLN47),.WL(WL232));
sram_cell_6t_5 inst_cell_232_48 (.BL(BL48),.BLN(BLN48),.WL(WL232));
sram_cell_6t_5 inst_cell_232_49 (.BL(BL49),.BLN(BLN49),.WL(WL232));
sram_cell_6t_5 inst_cell_232_50 (.BL(BL50),.BLN(BLN50),.WL(WL232));
sram_cell_6t_5 inst_cell_232_51 (.BL(BL51),.BLN(BLN51),.WL(WL232));
sram_cell_6t_5 inst_cell_232_52 (.BL(BL52),.BLN(BLN52),.WL(WL232));
sram_cell_6t_5 inst_cell_232_53 (.BL(BL53),.BLN(BLN53),.WL(WL232));
sram_cell_6t_5 inst_cell_232_54 (.BL(BL54),.BLN(BLN54),.WL(WL232));
sram_cell_6t_5 inst_cell_232_55 (.BL(BL55),.BLN(BLN55),.WL(WL232));
sram_cell_6t_5 inst_cell_232_56 (.BL(BL56),.BLN(BLN56),.WL(WL232));
sram_cell_6t_5 inst_cell_232_57 (.BL(BL57),.BLN(BLN57),.WL(WL232));
sram_cell_6t_5 inst_cell_232_58 (.BL(BL58),.BLN(BLN58),.WL(WL232));
sram_cell_6t_5 inst_cell_232_59 (.BL(BL59),.BLN(BLN59),.WL(WL232));
sram_cell_6t_5 inst_cell_232_60 (.BL(BL60),.BLN(BLN60),.WL(WL232));
sram_cell_6t_5 inst_cell_232_61 (.BL(BL61),.BLN(BLN61),.WL(WL232));
sram_cell_6t_5 inst_cell_232_62 (.BL(BL62),.BLN(BLN62),.WL(WL232));
sram_cell_6t_5 inst_cell_232_63 (.BL(BL63),.BLN(BLN63),.WL(WL232));
sram_cell_6t_5 inst_cell_232_64 (.BL(BL64),.BLN(BLN64),.WL(WL232));
sram_cell_6t_5 inst_cell_232_65 (.BL(BL65),.BLN(BLN65),.WL(WL232));
sram_cell_6t_5 inst_cell_232_66 (.BL(BL66),.BLN(BLN66),.WL(WL232));
sram_cell_6t_5 inst_cell_232_67 (.BL(BL67),.BLN(BLN67),.WL(WL232));
sram_cell_6t_5 inst_cell_232_68 (.BL(BL68),.BLN(BLN68),.WL(WL232));
sram_cell_6t_5 inst_cell_232_69 (.BL(BL69),.BLN(BLN69),.WL(WL232));
sram_cell_6t_5 inst_cell_232_70 (.BL(BL70),.BLN(BLN70),.WL(WL232));
sram_cell_6t_5 inst_cell_232_71 (.BL(BL71),.BLN(BLN71),.WL(WL232));
sram_cell_6t_5 inst_cell_232_72 (.BL(BL72),.BLN(BLN72),.WL(WL232));
sram_cell_6t_5 inst_cell_232_73 (.BL(BL73),.BLN(BLN73),.WL(WL232));
sram_cell_6t_5 inst_cell_232_74 (.BL(BL74),.BLN(BLN74),.WL(WL232));
sram_cell_6t_5 inst_cell_232_75 (.BL(BL75),.BLN(BLN75),.WL(WL232));
sram_cell_6t_5 inst_cell_232_76 (.BL(BL76),.BLN(BLN76),.WL(WL232));
sram_cell_6t_5 inst_cell_232_77 (.BL(BL77),.BLN(BLN77),.WL(WL232));
sram_cell_6t_5 inst_cell_232_78 (.BL(BL78),.BLN(BLN78),.WL(WL232));
sram_cell_6t_5 inst_cell_232_79 (.BL(BL79),.BLN(BLN79),.WL(WL232));
sram_cell_6t_5 inst_cell_232_80 (.BL(BL80),.BLN(BLN80),.WL(WL232));
sram_cell_6t_5 inst_cell_232_81 (.BL(BL81),.BLN(BLN81),.WL(WL232));
sram_cell_6t_5 inst_cell_232_82 (.BL(BL82),.BLN(BLN82),.WL(WL232));
sram_cell_6t_5 inst_cell_232_83 (.BL(BL83),.BLN(BLN83),.WL(WL232));
sram_cell_6t_5 inst_cell_232_84 (.BL(BL84),.BLN(BLN84),.WL(WL232));
sram_cell_6t_5 inst_cell_232_85 (.BL(BL85),.BLN(BLN85),.WL(WL232));
sram_cell_6t_5 inst_cell_232_86 (.BL(BL86),.BLN(BLN86),.WL(WL232));
sram_cell_6t_5 inst_cell_232_87 (.BL(BL87),.BLN(BLN87),.WL(WL232));
sram_cell_6t_5 inst_cell_232_88 (.BL(BL88),.BLN(BLN88),.WL(WL232));
sram_cell_6t_5 inst_cell_232_89 (.BL(BL89),.BLN(BLN89),.WL(WL232));
sram_cell_6t_5 inst_cell_232_90 (.BL(BL90),.BLN(BLN90),.WL(WL232));
sram_cell_6t_5 inst_cell_232_91 (.BL(BL91),.BLN(BLN91),.WL(WL232));
sram_cell_6t_5 inst_cell_232_92 (.BL(BL92),.BLN(BLN92),.WL(WL232));
sram_cell_6t_5 inst_cell_232_93 (.BL(BL93),.BLN(BLN93),.WL(WL232));
sram_cell_6t_5 inst_cell_232_94 (.BL(BL94),.BLN(BLN94),.WL(WL232));
sram_cell_6t_5 inst_cell_232_95 (.BL(BL95),.BLN(BLN95),.WL(WL232));
sram_cell_6t_5 inst_cell_232_96 (.BL(BL96),.BLN(BLN96),.WL(WL232));
sram_cell_6t_5 inst_cell_232_97 (.BL(BL97),.BLN(BLN97),.WL(WL232));
sram_cell_6t_5 inst_cell_232_98 (.BL(BL98),.BLN(BLN98),.WL(WL232));
sram_cell_6t_5 inst_cell_232_99 (.BL(BL99),.BLN(BLN99),.WL(WL232));
sram_cell_6t_5 inst_cell_232_100 (.BL(BL100),.BLN(BLN100),.WL(WL232));
sram_cell_6t_5 inst_cell_232_101 (.BL(BL101),.BLN(BLN101),.WL(WL232));
sram_cell_6t_5 inst_cell_232_102 (.BL(BL102),.BLN(BLN102),.WL(WL232));
sram_cell_6t_5 inst_cell_232_103 (.BL(BL103),.BLN(BLN103),.WL(WL232));
sram_cell_6t_5 inst_cell_232_104 (.BL(BL104),.BLN(BLN104),.WL(WL232));
sram_cell_6t_5 inst_cell_232_105 (.BL(BL105),.BLN(BLN105),.WL(WL232));
sram_cell_6t_5 inst_cell_232_106 (.BL(BL106),.BLN(BLN106),.WL(WL232));
sram_cell_6t_5 inst_cell_232_107 (.BL(BL107),.BLN(BLN107),.WL(WL232));
sram_cell_6t_5 inst_cell_232_108 (.BL(BL108),.BLN(BLN108),.WL(WL232));
sram_cell_6t_5 inst_cell_232_109 (.BL(BL109),.BLN(BLN109),.WL(WL232));
sram_cell_6t_5 inst_cell_232_110 (.BL(BL110),.BLN(BLN110),.WL(WL232));
sram_cell_6t_5 inst_cell_232_111 (.BL(BL111),.BLN(BLN111),.WL(WL232));
sram_cell_6t_5 inst_cell_232_112 (.BL(BL112),.BLN(BLN112),.WL(WL232));
sram_cell_6t_5 inst_cell_232_113 (.BL(BL113),.BLN(BLN113),.WL(WL232));
sram_cell_6t_5 inst_cell_232_114 (.BL(BL114),.BLN(BLN114),.WL(WL232));
sram_cell_6t_5 inst_cell_232_115 (.BL(BL115),.BLN(BLN115),.WL(WL232));
sram_cell_6t_5 inst_cell_232_116 (.BL(BL116),.BLN(BLN116),.WL(WL232));
sram_cell_6t_5 inst_cell_232_117 (.BL(BL117),.BLN(BLN117),.WL(WL232));
sram_cell_6t_5 inst_cell_232_118 (.BL(BL118),.BLN(BLN118),.WL(WL232));
sram_cell_6t_5 inst_cell_232_119 (.BL(BL119),.BLN(BLN119),.WL(WL232));
sram_cell_6t_5 inst_cell_232_120 (.BL(BL120),.BLN(BLN120),.WL(WL232));
sram_cell_6t_5 inst_cell_232_121 (.BL(BL121),.BLN(BLN121),.WL(WL232));
sram_cell_6t_5 inst_cell_232_122 (.BL(BL122),.BLN(BLN122),.WL(WL232));
sram_cell_6t_5 inst_cell_232_123 (.BL(BL123),.BLN(BLN123),.WL(WL232));
sram_cell_6t_5 inst_cell_232_124 (.BL(BL124),.BLN(BLN124),.WL(WL232));
sram_cell_6t_5 inst_cell_232_125 (.BL(BL125),.BLN(BLN125),.WL(WL232));
sram_cell_6t_5 inst_cell_232_126 (.BL(BL126),.BLN(BLN126),.WL(WL232));
sram_cell_6t_5 inst_cell_232_127 (.BL(BL127),.BLN(BLN127),.WL(WL232));
sram_cell_6t_5 inst_cell_233_0 (.BL(BL0),.BLN(BLN0),.WL(WL233));
sram_cell_6t_5 inst_cell_233_1 (.BL(BL1),.BLN(BLN1),.WL(WL233));
sram_cell_6t_5 inst_cell_233_2 (.BL(BL2),.BLN(BLN2),.WL(WL233));
sram_cell_6t_5 inst_cell_233_3 (.BL(BL3),.BLN(BLN3),.WL(WL233));
sram_cell_6t_5 inst_cell_233_4 (.BL(BL4),.BLN(BLN4),.WL(WL233));
sram_cell_6t_5 inst_cell_233_5 (.BL(BL5),.BLN(BLN5),.WL(WL233));
sram_cell_6t_5 inst_cell_233_6 (.BL(BL6),.BLN(BLN6),.WL(WL233));
sram_cell_6t_5 inst_cell_233_7 (.BL(BL7),.BLN(BLN7),.WL(WL233));
sram_cell_6t_5 inst_cell_233_8 (.BL(BL8),.BLN(BLN8),.WL(WL233));
sram_cell_6t_5 inst_cell_233_9 (.BL(BL9),.BLN(BLN9),.WL(WL233));
sram_cell_6t_5 inst_cell_233_10 (.BL(BL10),.BLN(BLN10),.WL(WL233));
sram_cell_6t_5 inst_cell_233_11 (.BL(BL11),.BLN(BLN11),.WL(WL233));
sram_cell_6t_5 inst_cell_233_12 (.BL(BL12),.BLN(BLN12),.WL(WL233));
sram_cell_6t_5 inst_cell_233_13 (.BL(BL13),.BLN(BLN13),.WL(WL233));
sram_cell_6t_5 inst_cell_233_14 (.BL(BL14),.BLN(BLN14),.WL(WL233));
sram_cell_6t_5 inst_cell_233_15 (.BL(BL15),.BLN(BLN15),.WL(WL233));
sram_cell_6t_5 inst_cell_233_16 (.BL(BL16),.BLN(BLN16),.WL(WL233));
sram_cell_6t_5 inst_cell_233_17 (.BL(BL17),.BLN(BLN17),.WL(WL233));
sram_cell_6t_5 inst_cell_233_18 (.BL(BL18),.BLN(BLN18),.WL(WL233));
sram_cell_6t_5 inst_cell_233_19 (.BL(BL19),.BLN(BLN19),.WL(WL233));
sram_cell_6t_5 inst_cell_233_20 (.BL(BL20),.BLN(BLN20),.WL(WL233));
sram_cell_6t_5 inst_cell_233_21 (.BL(BL21),.BLN(BLN21),.WL(WL233));
sram_cell_6t_5 inst_cell_233_22 (.BL(BL22),.BLN(BLN22),.WL(WL233));
sram_cell_6t_5 inst_cell_233_23 (.BL(BL23),.BLN(BLN23),.WL(WL233));
sram_cell_6t_5 inst_cell_233_24 (.BL(BL24),.BLN(BLN24),.WL(WL233));
sram_cell_6t_5 inst_cell_233_25 (.BL(BL25),.BLN(BLN25),.WL(WL233));
sram_cell_6t_5 inst_cell_233_26 (.BL(BL26),.BLN(BLN26),.WL(WL233));
sram_cell_6t_5 inst_cell_233_27 (.BL(BL27),.BLN(BLN27),.WL(WL233));
sram_cell_6t_5 inst_cell_233_28 (.BL(BL28),.BLN(BLN28),.WL(WL233));
sram_cell_6t_5 inst_cell_233_29 (.BL(BL29),.BLN(BLN29),.WL(WL233));
sram_cell_6t_5 inst_cell_233_30 (.BL(BL30),.BLN(BLN30),.WL(WL233));
sram_cell_6t_5 inst_cell_233_31 (.BL(BL31),.BLN(BLN31),.WL(WL233));
sram_cell_6t_5 inst_cell_233_32 (.BL(BL32),.BLN(BLN32),.WL(WL233));
sram_cell_6t_5 inst_cell_233_33 (.BL(BL33),.BLN(BLN33),.WL(WL233));
sram_cell_6t_5 inst_cell_233_34 (.BL(BL34),.BLN(BLN34),.WL(WL233));
sram_cell_6t_5 inst_cell_233_35 (.BL(BL35),.BLN(BLN35),.WL(WL233));
sram_cell_6t_5 inst_cell_233_36 (.BL(BL36),.BLN(BLN36),.WL(WL233));
sram_cell_6t_5 inst_cell_233_37 (.BL(BL37),.BLN(BLN37),.WL(WL233));
sram_cell_6t_5 inst_cell_233_38 (.BL(BL38),.BLN(BLN38),.WL(WL233));
sram_cell_6t_5 inst_cell_233_39 (.BL(BL39),.BLN(BLN39),.WL(WL233));
sram_cell_6t_5 inst_cell_233_40 (.BL(BL40),.BLN(BLN40),.WL(WL233));
sram_cell_6t_5 inst_cell_233_41 (.BL(BL41),.BLN(BLN41),.WL(WL233));
sram_cell_6t_5 inst_cell_233_42 (.BL(BL42),.BLN(BLN42),.WL(WL233));
sram_cell_6t_5 inst_cell_233_43 (.BL(BL43),.BLN(BLN43),.WL(WL233));
sram_cell_6t_5 inst_cell_233_44 (.BL(BL44),.BLN(BLN44),.WL(WL233));
sram_cell_6t_5 inst_cell_233_45 (.BL(BL45),.BLN(BLN45),.WL(WL233));
sram_cell_6t_5 inst_cell_233_46 (.BL(BL46),.BLN(BLN46),.WL(WL233));
sram_cell_6t_5 inst_cell_233_47 (.BL(BL47),.BLN(BLN47),.WL(WL233));
sram_cell_6t_5 inst_cell_233_48 (.BL(BL48),.BLN(BLN48),.WL(WL233));
sram_cell_6t_5 inst_cell_233_49 (.BL(BL49),.BLN(BLN49),.WL(WL233));
sram_cell_6t_5 inst_cell_233_50 (.BL(BL50),.BLN(BLN50),.WL(WL233));
sram_cell_6t_5 inst_cell_233_51 (.BL(BL51),.BLN(BLN51),.WL(WL233));
sram_cell_6t_5 inst_cell_233_52 (.BL(BL52),.BLN(BLN52),.WL(WL233));
sram_cell_6t_5 inst_cell_233_53 (.BL(BL53),.BLN(BLN53),.WL(WL233));
sram_cell_6t_5 inst_cell_233_54 (.BL(BL54),.BLN(BLN54),.WL(WL233));
sram_cell_6t_5 inst_cell_233_55 (.BL(BL55),.BLN(BLN55),.WL(WL233));
sram_cell_6t_5 inst_cell_233_56 (.BL(BL56),.BLN(BLN56),.WL(WL233));
sram_cell_6t_5 inst_cell_233_57 (.BL(BL57),.BLN(BLN57),.WL(WL233));
sram_cell_6t_5 inst_cell_233_58 (.BL(BL58),.BLN(BLN58),.WL(WL233));
sram_cell_6t_5 inst_cell_233_59 (.BL(BL59),.BLN(BLN59),.WL(WL233));
sram_cell_6t_5 inst_cell_233_60 (.BL(BL60),.BLN(BLN60),.WL(WL233));
sram_cell_6t_5 inst_cell_233_61 (.BL(BL61),.BLN(BLN61),.WL(WL233));
sram_cell_6t_5 inst_cell_233_62 (.BL(BL62),.BLN(BLN62),.WL(WL233));
sram_cell_6t_5 inst_cell_233_63 (.BL(BL63),.BLN(BLN63),.WL(WL233));
sram_cell_6t_5 inst_cell_233_64 (.BL(BL64),.BLN(BLN64),.WL(WL233));
sram_cell_6t_5 inst_cell_233_65 (.BL(BL65),.BLN(BLN65),.WL(WL233));
sram_cell_6t_5 inst_cell_233_66 (.BL(BL66),.BLN(BLN66),.WL(WL233));
sram_cell_6t_5 inst_cell_233_67 (.BL(BL67),.BLN(BLN67),.WL(WL233));
sram_cell_6t_5 inst_cell_233_68 (.BL(BL68),.BLN(BLN68),.WL(WL233));
sram_cell_6t_5 inst_cell_233_69 (.BL(BL69),.BLN(BLN69),.WL(WL233));
sram_cell_6t_5 inst_cell_233_70 (.BL(BL70),.BLN(BLN70),.WL(WL233));
sram_cell_6t_5 inst_cell_233_71 (.BL(BL71),.BLN(BLN71),.WL(WL233));
sram_cell_6t_5 inst_cell_233_72 (.BL(BL72),.BLN(BLN72),.WL(WL233));
sram_cell_6t_5 inst_cell_233_73 (.BL(BL73),.BLN(BLN73),.WL(WL233));
sram_cell_6t_5 inst_cell_233_74 (.BL(BL74),.BLN(BLN74),.WL(WL233));
sram_cell_6t_5 inst_cell_233_75 (.BL(BL75),.BLN(BLN75),.WL(WL233));
sram_cell_6t_5 inst_cell_233_76 (.BL(BL76),.BLN(BLN76),.WL(WL233));
sram_cell_6t_5 inst_cell_233_77 (.BL(BL77),.BLN(BLN77),.WL(WL233));
sram_cell_6t_5 inst_cell_233_78 (.BL(BL78),.BLN(BLN78),.WL(WL233));
sram_cell_6t_5 inst_cell_233_79 (.BL(BL79),.BLN(BLN79),.WL(WL233));
sram_cell_6t_5 inst_cell_233_80 (.BL(BL80),.BLN(BLN80),.WL(WL233));
sram_cell_6t_5 inst_cell_233_81 (.BL(BL81),.BLN(BLN81),.WL(WL233));
sram_cell_6t_5 inst_cell_233_82 (.BL(BL82),.BLN(BLN82),.WL(WL233));
sram_cell_6t_5 inst_cell_233_83 (.BL(BL83),.BLN(BLN83),.WL(WL233));
sram_cell_6t_5 inst_cell_233_84 (.BL(BL84),.BLN(BLN84),.WL(WL233));
sram_cell_6t_5 inst_cell_233_85 (.BL(BL85),.BLN(BLN85),.WL(WL233));
sram_cell_6t_5 inst_cell_233_86 (.BL(BL86),.BLN(BLN86),.WL(WL233));
sram_cell_6t_5 inst_cell_233_87 (.BL(BL87),.BLN(BLN87),.WL(WL233));
sram_cell_6t_5 inst_cell_233_88 (.BL(BL88),.BLN(BLN88),.WL(WL233));
sram_cell_6t_5 inst_cell_233_89 (.BL(BL89),.BLN(BLN89),.WL(WL233));
sram_cell_6t_5 inst_cell_233_90 (.BL(BL90),.BLN(BLN90),.WL(WL233));
sram_cell_6t_5 inst_cell_233_91 (.BL(BL91),.BLN(BLN91),.WL(WL233));
sram_cell_6t_5 inst_cell_233_92 (.BL(BL92),.BLN(BLN92),.WL(WL233));
sram_cell_6t_5 inst_cell_233_93 (.BL(BL93),.BLN(BLN93),.WL(WL233));
sram_cell_6t_5 inst_cell_233_94 (.BL(BL94),.BLN(BLN94),.WL(WL233));
sram_cell_6t_5 inst_cell_233_95 (.BL(BL95),.BLN(BLN95),.WL(WL233));
sram_cell_6t_5 inst_cell_233_96 (.BL(BL96),.BLN(BLN96),.WL(WL233));
sram_cell_6t_5 inst_cell_233_97 (.BL(BL97),.BLN(BLN97),.WL(WL233));
sram_cell_6t_5 inst_cell_233_98 (.BL(BL98),.BLN(BLN98),.WL(WL233));
sram_cell_6t_5 inst_cell_233_99 (.BL(BL99),.BLN(BLN99),.WL(WL233));
sram_cell_6t_5 inst_cell_233_100 (.BL(BL100),.BLN(BLN100),.WL(WL233));
sram_cell_6t_5 inst_cell_233_101 (.BL(BL101),.BLN(BLN101),.WL(WL233));
sram_cell_6t_5 inst_cell_233_102 (.BL(BL102),.BLN(BLN102),.WL(WL233));
sram_cell_6t_5 inst_cell_233_103 (.BL(BL103),.BLN(BLN103),.WL(WL233));
sram_cell_6t_5 inst_cell_233_104 (.BL(BL104),.BLN(BLN104),.WL(WL233));
sram_cell_6t_5 inst_cell_233_105 (.BL(BL105),.BLN(BLN105),.WL(WL233));
sram_cell_6t_5 inst_cell_233_106 (.BL(BL106),.BLN(BLN106),.WL(WL233));
sram_cell_6t_5 inst_cell_233_107 (.BL(BL107),.BLN(BLN107),.WL(WL233));
sram_cell_6t_5 inst_cell_233_108 (.BL(BL108),.BLN(BLN108),.WL(WL233));
sram_cell_6t_5 inst_cell_233_109 (.BL(BL109),.BLN(BLN109),.WL(WL233));
sram_cell_6t_5 inst_cell_233_110 (.BL(BL110),.BLN(BLN110),.WL(WL233));
sram_cell_6t_5 inst_cell_233_111 (.BL(BL111),.BLN(BLN111),.WL(WL233));
sram_cell_6t_5 inst_cell_233_112 (.BL(BL112),.BLN(BLN112),.WL(WL233));
sram_cell_6t_5 inst_cell_233_113 (.BL(BL113),.BLN(BLN113),.WL(WL233));
sram_cell_6t_5 inst_cell_233_114 (.BL(BL114),.BLN(BLN114),.WL(WL233));
sram_cell_6t_5 inst_cell_233_115 (.BL(BL115),.BLN(BLN115),.WL(WL233));
sram_cell_6t_5 inst_cell_233_116 (.BL(BL116),.BLN(BLN116),.WL(WL233));
sram_cell_6t_5 inst_cell_233_117 (.BL(BL117),.BLN(BLN117),.WL(WL233));
sram_cell_6t_5 inst_cell_233_118 (.BL(BL118),.BLN(BLN118),.WL(WL233));
sram_cell_6t_5 inst_cell_233_119 (.BL(BL119),.BLN(BLN119),.WL(WL233));
sram_cell_6t_5 inst_cell_233_120 (.BL(BL120),.BLN(BLN120),.WL(WL233));
sram_cell_6t_5 inst_cell_233_121 (.BL(BL121),.BLN(BLN121),.WL(WL233));
sram_cell_6t_5 inst_cell_233_122 (.BL(BL122),.BLN(BLN122),.WL(WL233));
sram_cell_6t_5 inst_cell_233_123 (.BL(BL123),.BLN(BLN123),.WL(WL233));
sram_cell_6t_5 inst_cell_233_124 (.BL(BL124),.BLN(BLN124),.WL(WL233));
sram_cell_6t_5 inst_cell_233_125 (.BL(BL125),.BLN(BLN125),.WL(WL233));
sram_cell_6t_5 inst_cell_233_126 (.BL(BL126),.BLN(BLN126),.WL(WL233));
sram_cell_6t_5 inst_cell_233_127 (.BL(BL127),.BLN(BLN127),.WL(WL233));
sram_cell_6t_5 inst_cell_234_0 (.BL(BL0),.BLN(BLN0),.WL(WL234));
sram_cell_6t_5 inst_cell_234_1 (.BL(BL1),.BLN(BLN1),.WL(WL234));
sram_cell_6t_5 inst_cell_234_2 (.BL(BL2),.BLN(BLN2),.WL(WL234));
sram_cell_6t_5 inst_cell_234_3 (.BL(BL3),.BLN(BLN3),.WL(WL234));
sram_cell_6t_5 inst_cell_234_4 (.BL(BL4),.BLN(BLN4),.WL(WL234));
sram_cell_6t_5 inst_cell_234_5 (.BL(BL5),.BLN(BLN5),.WL(WL234));
sram_cell_6t_5 inst_cell_234_6 (.BL(BL6),.BLN(BLN6),.WL(WL234));
sram_cell_6t_5 inst_cell_234_7 (.BL(BL7),.BLN(BLN7),.WL(WL234));
sram_cell_6t_5 inst_cell_234_8 (.BL(BL8),.BLN(BLN8),.WL(WL234));
sram_cell_6t_5 inst_cell_234_9 (.BL(BL9),.BLN(BLN9),.WL(WL234));
sram_cell_6t_5 inst_cell_234_10 (.BL(BL10),.BLN(BLN10),.WL(WL234));
sram_cell_6t_5 inst_cell_234_11 (.BL(BL11),.BLN(BLN11),.WL(WL234));
sram_cell_6t_5 inst_cell_234_12 (.BL(BL12),.BLN(BLN12),.WL(WL234));
sram_cell_6t_5 inst_cell_234_13 (.BL(BL13),.BLN(BLN13),.WL(WL234));
sram_cell_6t_5 inst_cell_234_14 (.BL(BL14),.BLN(BLN14),.WL(WL234));
sram_cell_6t_5 inst_cell_234_15 (.BL(BL15),.BLN(BLN15),.WL(WL234));
sram_cell_6t_5 inst_cell_234_16 (.BL(BL16),.BLN(BLN16),.WL(WL234));
sram_cell_6t_5 inst_cell_234_17 (.BL(BL17),.BLN(BLN17),.WL(WL234));
sram_cell_6t_5 inst_cell_234_18 (.BL(BL18),.BLN(BLN18),.WL(WL234));
sram_cell_6t_5 inst_cell_234_19 (.BL(BL19),.BLN(BLN19),.WL(WL234));
sram_cell_6t_5 inst_cell_234_20 (.BL(BL20),.BLN(BLN20),.WL(WL234));
sram_cell_6t_5 inst_cell_234_21 (.BL(BL21),.BLN(BLN21),.WL(WL234));
sram_cell_6t_5 inst_cell_234_22 (.BL(BL22),.BLN(BLN22),.WL(WL234));
sram_cell_6t_5 inst_cell_234_23 (.BL(BL23),.BLN(BLN23),.WL(WL234));
sram_cell_6t_5 inst_cell_234_24 (.BL(BL24),.BLN(BLN24),.WL(WL234));
sram_cell_6t_5 inst_cell_234_25 (.BL(BL25),.BLN(BLN25),.WL(WL234));
sram_cell_6t_5 inst_cell_234_26 (.BL(BL26),.BLN(BLN26),.WL(WL234));
sram_cell_6t_5 inst_cell_234_27 (.BL(BL27),.BLN(BLN27),.WL(WL234));
sram_cell_6t_5 inst_cell_234_28 (.BL(BL28),.BLN(BLN28),.WL(WL234));
sram_cell_6t_5 inst_cell_234_29 (.BL(BL29),.BLN(BLN29),.WL(WL234));
sram_cell_6t_5 inst_cell_234_30 (.BL(BL30),.BLN(BLN30),.WL(WL234));
sram_cell_6t_5 inst_cell_234_31 (.BL(BL31),.BLN(BLN31),.WL(WL234));
sram_cell_6t_5 inst_cell_234_32 (.BL(BL32),.BLN(BLN32),.WL(WL234));
sram_cell_6t_5 inst_cell_234_33 (.BL(BL33),.BLN(BLN33),.WL(WL234));
sram_cell_6t_5 inst_cell_234_34 (.BL(BL34),.BLN(BLN34),.WL(WL234));
sram_cell_6t_5 inst_cell_234_35 (.BL(BL35),.BLN(BLN35),.WL(WL234));
sram_cell_6t_5 inst_cell_234_36 (.BL(BL36),.BLN(BLN36),.WL(WL234));
sram_cell_6t_5 inst_cell_234_37 (.BL(BL37),.BLN(BLN37),.WL(WL234));
sram_cell_6t_5 inst_cell_234_38 (.BL(BL38),.BLN(BLN38),.WL(WL234));
sram_cell_6t_5 inst_cell_234_39 (.BL(BL39),.BLN(BLN39),.WL(WL234));
sram_cell_6t_5 inst_cell_234_40 (.BL(BL40),.BLN(BLN40),.WL(WL234));
sram_cell_6t_5 inst_cell_234_41 (.BL(BL41),.BLN(BLN41),.WL(WL234));
sram_cell_6t_5 inst_cell_234_42 (.BL(BL42),.BLN(BLN42),.WL(WL234));
sram_cell_6t_5 inst_cell_234_43 (.BL(BL43),.BLN(BLN43),.WL(WL234));
sram_cell_6t_5 inst_cell_234_44 (.BL(BL44),.BLN(BLN44),.WL(WL234));
sram_cell_6t_5 inst_cell_234_45 (.BL(BL45),.BLN(BLN45),.WL(WL234));
sram_cell_6t_5 inst_cell_234_46 (.BL(BL46),.BLN(BLN46),.WL(WL234));
sram_cell_6t_5 inst_cell_234_47 (.BL(BL47),.BLN(BLN47),.WL(WL234));
sram_cell_6t_5 inst_cell_234_48 (.BL(BL48),.BLN(BLN48),.WL(WL234));
sram_cell_6t_5 inst_cell_234_49 (.BL(BL49),.BLN(BLN49),.WL(WL234));
sram_cell_6t_5 inst_cell_234_50 (.BL(BL50),.BLN(BLN50),.WL(WL234));
sram_cell_6t_5 inst_cell_234_51 (.BL(BL51),.BLN(BLN51),.WL(WL234));
sram_cell_6t_5 inst_cell_234_52 (.BL(BL52),.BLN(BLN52),.WL(WL234));
sram_cell_6t_5 inst_cell_234_53 (.BL(BL53),.BLN(BLN53),.WL(WL234));
sram_cell_6t_5 inst_cell_234_54 (.BL(BL54),.BLN(BLN54),.WL(WL234));
sram_cell_6t_5 inst_cell_234_55 (.BL(BL55),.BLN(BLN55),.WL(WL234));
sram_cell_6t_5 inst_cell_234_56 (.BL(BL56),.BLN(BLN56),.WL(WL234));
sram_cell_6t_5 inst_cell_234_57 (.BL(BL57),.BLN(BLN57),.WL(WL234));
sram_cell_6t_5 inst_cell_234_58 (.BL(BL58),.BLN(BLN58),.WL(WL234));
sram_cell_6t_5 inst_cell_234_59 (.BL(BL59),.BLN(BLN59),.WL(WL234));
sram_cell_6t_5 inst_cell_234_60 (.BL(BL60),.BLN(BLN60),.WL(WL234));
sram_cell_6t_5 inst_cell_234_61 (.BL(BL61),.BLN(BLN61),.WL(WL234));
sram_cell_6t_5 inst_cell_234_62 (.BL(BL62),.BLN(BLN62),.WL(WL234));
sram_cell_6t_5 inst_cell_234_63 (.BL(BL63),.BLN(BLN63),.WL(WL234));
sram_cell_6t_5 inst_cell_234_64 (.BL(BL64),.BLN(BLN64),.WL(WL234));
sram_cell_6t_5 inst_cell_234_65 (.BL(BL65),.BLN(BLN65),.WL(WL234));
sram_cell_6t_5 inst_cell_234_66 (.BL(BL66),.BLN(BLN66),.WL(WL234));
sram_cell_6t_5 inst_cell_234_67 (.BL(BL67),.BLN(BLN67),.WL(WL234));
sram_cell_6t_5 inst_cell_234_68 (.BL(BL68),.BLN(BLN68),.WL(WL234));
sram_cell_6t_5 inst_cell_234_69 (.BL(BL69),.BLN(BLN69),.WL(WL234));
sram_cell_6t_5 inst_cell_234_70 (.BL(BL70),.BLN(BLN70),.WL(WL234));
sram_cell_6t_5 inst_cell_234_71 (.BL(BL71),.BLN(BLN71),.WL(WL234));
sram_cell_6t_5 inst_cell_234_72 (.BL(BL72),.BLN(BLN72),.WL(WL234));
sram_cell_6t_5 inst_cell_234_73 (.BL(BL73),.BLN(BLN73),.WL(WL234));
sram_cell_6t_5 inst_cell_234_74 (.BL(BL74),.BLN(BLN74),.WL(WL234));
sram_cell_6t_5 inst_cell_234_75 (.BL(BL75),.BLN(BLN75),.WL(WL234));
sram_cell_6t_5 inst_cell_234_76 (.BL(BL76),.BLN(BLN76),.WL(WL234));
sram_cell_6t_5 inst_cell_234_77 (.BL(BL77),.BLN(BLN77),.WL(WL234));
sram_cell_6t_5 inst_cell_234_78 (.BL(BL78),.BLN(BLN78),.WL(WL234));
sram_cell_6t_5 inst_cell_234_79 (.BL(BL79),.BLN(BLN79),.WL(WL234));
sram_cell_6t_5 inst_cell_234_80 (.BL(BL80),.BLN(BLN80),.WL(WL234));
sram_cell_6t_5 inst_cell_234_81 (.BL(BL81),.BLN(BLN81),.WL(WL234));
sram_cell_6t_5 inst_cell_234_82 (.BL(BL82),.BLN(BLN82),.WL(WL234));
sram_cell_6t_5 inst_cell_234_83 (.BL(BL83),.BLN(BLN83),.WL(WL234));
sram_cell_6t_5 inst_cell_234_84 (.BL(BL84),.BLN(BLN84),.WL(WL234));
sram_cell_6t_5 inst_cell_234_85 (.BL(BL85),.BLN(BLN85),.WL(WL234));
sram_cell_6t_5 inst_cell_234_86 (.BL(BL86),.BLN(BLN86),.WL(WL234));
sram_cell_6t_5 inst_cell_234_87 (.BL(BL87),.BLN(BLN87),.WL(WL234));
sram_cell_6t_5 inst_cell_234_88 (.BL(BL88),.BLN(BLN88),.WL(WL234));
sram_cell_6t_5 inst_cell_234_89 (.BL(BL89),.BLN(BLN89),.WL(WL234));
sram_cell_6t_5 inst_cell_234_90 (.BL(BL90),.BLN(BLN90),.WL(WL234));
sram_cell_6t_5 inst_cell_234_91 (.BL(BL91),.BLN(BLN91),.WL(WL234));
sram_cell_6t_5 inst_cell_234_92 (.BL(BL92),.BLN(BLN92),.WL(WL234));
sram_cell_6t_5 inst_cell_234_93 (.BL(BL93),.BLN(BLN93),.WL(WL234));
sram_cell_6t_5 inst_cell_234_94 (.BL(BL94),.BLN(BLN94),.WL(WL234));
sram_cell_6t_5 inst_cell_234_95 (.BL(BL95),.BLN(BLN95),.WL(WL234));
sram_cell_6t_5 inst_cell_234_96 (.BL(BL96),.BLN(BLN96),.WL(WL234));
sram_cell_6t_5 inst_cell_234_97 (.BL(BL97),.BLN(BLN97),.WL(WL234));
sram_cell_6t_5 inst_cell_234_98 (.BL(BL98),.BLN(BLN98),.WL(WL234));
sram_cell_6t_5 inst_cell_234_99 (.BL(BL99),.BLN(BLN99),.WL(WL234));
sram_cell_6t_5 inst_cell_234_100 (.BL(BL100),.BLN(BLN100),.WL(WL234));
sram_cell_6t_5 inst_cell_234_101 (.BL(BL101),.BLN(BLN101),.WL(WL234));
sram_cell_6t_5 inst_cell_234_102 (.BL(BL102),.BLN(BLN102),.WL(WL234));
sram_cell_6t_5 inst_cell_234_103 (.BL(BL103),.BLN(BLN103),.WL(WL234));
sram_cell_6t_5 inst_cell_234_104 (.BL(BL104),.BLN(BLN104),.WL(WL234));
sram_cell_6t_5 inst_cell_234_105 (.BL(BL105),.BLN(BLN105),.WL(WL234));
sram_cell_6t_5 inst_cell_234_106 (.BL(BL106),.BLN(BLN106),.WL(WL234));
sram_cell_6t_5 inst_cell_234_107 (.BL(BL107),.BLN(BLN107),.WL(WL234));
sram_cell_6t_5 inst_cell_234_108 (.BL(BL108),.BLN(BLN108),.WL(WL234));
sram_cell_6t_5 inst_cell_234_109 (.BL(BL109),.BLN(BLN109),.WL(WL234));
sram_cell_6t_5 inst_cell_234_110 (.BL(BL110),.BLN(BLN110),.WL(WL234));
sram_cell_6t_5 inst_cell_234_111 (.BL(BL111),.BLN(BLN111),.WL(WL234));
sram_cell_6t_5 inst_cell_234_112 (.BL(BL112),.BLN(BLN112),.WL(WL234));
sram_cell_6t_5 inst_cell_234_113 (.BL(BL113),.BLN(BLN113),.WL(WL234));
sram_cell_6t_5 inst_cell_234_114 (.BL(BL114),.BLN(BLN114),.WL(WL234));
sram_cell_6t_5 inst_cell_234_115 (.BL(BL115),.BLN(BLN115),.WL(WL234));
sram_cell_6t_5 inst_cell_234_116 (.BL(BL116),.BLN(BLN116),.WL(WL234));
sram_cell_6t_5 inst_cell_234_117 (.BL(BL117),.BLN(BLN117),.WL(WL234));
sram_cell_6t_5 inst_cell_234_118 (.BL(BL118),.BLN(BLN118),.WL(WL234));
sram_cell_6t_5 inst_cell_234_119 (.BL(BL119),.BLN(BLN119),.WL(WL234));
sram_cell_6t_5 inst_cell_234_120 (.BL(BL120),.BLN(BLN120),.WL(WL234));
sram_cell_6t_5 inst_cell_234_121 (.BL(BL121),.BLN(BLN121),.WL(WL234));
sram_cell_6t_5 inst_cell_234_122 (.BL(BL122),.BLN(BLN122),.WL(WL234));
sram_cell_6t_5 inst_cell_234_123 (.BL(BL123),.BLN(BLN123),.WL(WL234));
sram_cell_6t_5 inst_cell_234_124 (.BL(BL124),.BLN(BLN124),.WL(WL234));
sram_cell_6t_5 inst_cell_234_125 (.BL(BL125),.BLN(BLN125),.WL(WL234));
sram_cell_6t_5 inst_cell_234_126 (.BL(BL126),.BLN(BLN126),.WL(WL234));
sram_cell_6t_5 inst_cell_234_127 (.BL(BL127),.BLN(BLN127),.WL(WL234));
sram_cell_6t_5 inst_cell_235_0 (.BL(BL0),.BLN(BLN0),.WL(WL235));
sram_cell_6t_5 inst_cell_235_1 (.BL(BL1),.BLN(BLN1),.WL(WL235));
sram_cell_6t_5 inst_cell_235_2 (.BL(BL2),.BLN(BLN2),.WL(WL235));
sram_cell_6t_5 inst_cell_235_3 (.BL(BL3),.BLN(BLN3),.WL(WL235));
sram_cell_6t_5 inst_cell_235_4 (.BL(BL4),.BLN(BLN4),.WL(WL235));
sram_cell_6t_5 inst_cell_235_5 (.BL(BL5),.BLN(BLN5),.WL(WL235));
sram_cell_6t_5 inst_cell_235_6 (.BL(BL6),.BLN(BLN6),.WL(WL235));
sram_cell_6t_5 inst_cell_235_7 (.BL(BL7),.BLN(BLN7),.WL(WL235));
sram_cell_6t_5 inst_cell_235_8 (.BL(BL8),.BLN(BLN8),.WL(WL235));
sram_cell_6t_5 inst_cell_235_9 (.BL(BL9),.BLN(BLN9),.WL(WL235));
sram_cell_6t_5 inst_cell_235_10 (.BL(BL10),.BLN(BLN10),.WL(WL235));
sram_cell_6t_5 inst_cell_235_11 (.BL(BL11),.BLN(BLN11),.WL(WL235));
sram_cell_6t_5 inst_cell_235_12 (.BL(BL12),.BLN(BLN12),.WL(WL235));
sram_cell_6t_5 inst_cell_235_13 (.BL(BL13),.BLN(BLN13),.WL(WL235));
sram_cell_6t_5 inst_cell_235_14 (.BL(BL14),.BLN(BLN14),.WL(WL235));
sram_cell_6t_5 inst_cell_235_15 (.BL(BL15),.BLN(BLN15),.WL(WL235));
sram_cell_6t_5 inst_cell_235_16 (.BL(BL16),.BLN(BLN16),.WL(WL235));
sram_cell_6t_5 inst_cell_235_17 (.BL(BL17),.BLN(BLN17),.WL(WL235));
sram_cell_6t_5 inst_cell_235_18 (.BL(BL18),.BLN(BLN18),.WL(WL235));
sram_cell_6t_5 inst_cell_235_19 (.BL(BL19),.BLN(BLN19),.WL(WL235));
sram_cell_6t_5 inst_cell_235_20 (.BL(BL20),.BLN(BLN20),.WL(WL235));
sram_cell_6t_5 inst_cell_235_21 (.BL(BL21),.BLN(BLN21),.WL(WL235));
sram_cell_6t_5 inst_cell_235_22 (.BL(BL22),.BLN(BLN22),.WL(WL235));
sram_cell_6t_5 inst_cell_235_23 (.BL(BL23),.BLN(BLN23),.WL(WL235));
sram_cell_6t_5 inst_cell_235_24 (.BL(BL24),.BLN(BLN24),.WL(WL235));
sram_cell_6t_5 inst_cell_235_25 (.BL(BL25),.BLN(BLN25),.WL(WL235));
sram_cell_6t_5 inst_cell_235_26 (.BL(BL26),.BLN(BLN26),.WL(WL235));
sram_cell_6t_5 inst_cell_235_27 (.BL(BL27),.BLN(BLN27),.WL(WL235));
sram_cell_6t_5 inst_cell_235_28 (.BL(BL28),.BLN(BLN28),.WL(WL235));
sram_cell_6t_5 inst_cell_235_29 (.BL(BL29),.BLN(BLN29),.WL(WL235));
sram_cell_6t_5 inst_cell_235_30 (.BL(BL30),.BLN(BLN30),.WL(WL235));
sram_cell_6t_5 inst_cell_235_31 (.BL(BL31),.BLN(BLN31),.WL(WL235));
sram_cell_6t_5 inst_cell_235_32 (.BL(BL32),.BLN(BLN32),.WL(WL235));
sram_cell_6t_5 inst_cell_235_33 (.BL(BL33),.BLN(BLN33),.WL(WL235));
sram_cell_6t_5 inst_cell_235_34 (.BL(BL34),.BLN(BLN34),.WL(WL235));
sram_cell_6t_5 inst_cell_235_35 (.BL(BL35),.BLN(BLN35),.WL(WL235));
sram_cell_6t_5 inst_cell_235_36 (.BL(BL36),.BLN(BLN36),.WL(WL235));
sram_cell_6t_5 inst_cell_235_37 (.BL(BL37),.BLN(BLN37),.WL(WL235));
sram_cell_6t_5 inst_cell_235_38 (.BL(BL38),.BLN(BLN38),.WL(WL235));
sram_cell_6t_5 inst_cell_235_39 (.BL(BL39),.BLN(BLN39),.WL(WL235));
sram_cell_6t_5 inst_cell_235_40 (.BL(BL40),.BLN(BLN40),.WL(WL235));
sram_cell_6t_5 inst_cell_235_41 (.BL(BL41),.BLN(BLN41),.WL(WL235));
sram_cell_6t_5 inst_cell_235_42 (.BL(BL42),.BLN(BLN42),.WL(WL235));
sram_cell_6t_5 inst_cell_235_43 (.BL(BL43),.BLN(BLN43),.WL(WL235));
sram_cell_6t_5 inst_cell_235_44 (.BL(BL44),.BLN(BLN44),.WL(WL235));
sram_cell_6t_5 inst_cell_235_45 (.BL(BL45),.BLN(BLN45),.WL(WL235));
sram_cell_6t_5 inst_cell_235_46 (.BL(BL46),.BLN(BLN46),.WL(WL235));
sram_cell_6t_5 inst_cell_235_47 (.BL(BL47),.BLN(BLN47),.WL(WL235));
sram_cell_6t_5 inst_cell_235_48 (.BL(BL48),.BLN(BLN48),.WL(WL235));
sram_cell_6t_5 inst_cell_235_49 (.BL(BL49),.BLN(BLN49),.WL(WL235));
sram_cell_6t_5 inst_cell_235_50 (.BL(BL50),.BLN(BLN50),.WL(WL235));
sram_cell_6t_5 inst_cell_235_51 (.BL(BL51),.BLN(BLN51),.WL(WL235));
sram_cell_6t_5 inst_cell_235_52 (.BL(BL52),.BLN(BLN52),.WL(WL235));
sram_cell_6t_5 inst_cell_235_53 (.BL(BL53),.BLN(BLN53),.WL(WL235));
sram_cell_6t_5 inst_cell_235_54 (.BL(BL54),.BLN(BLN54),.WL(WL235));
sram_cell_6t_5 inst_cell_235_55 (.BL(BL55),.BLN(BLN55),.WL(WL235));
sram_cell_6t_5 inst_cell_235_56 (.BL(BL56),.BLN(BLN56),.WL(WL235));
sram_cell_6t_5 inst_cell_235_57 (.BL(BL57),.BLN(BLN57),.WL(WL235));
sram_cell_6t_5 inst_cell_235_58 (.BL(BL58),.BLN(BLN58),.WL(WL235));
sram_cell_6t_5 inst_cell_235_59 (.BL(BL59),.BLN(BLN59),.WL(WL235));
sram_cell_6t_5 inst_cell_235_60 (.BL(BL60),.BLN(BLN60),.WL(WL235));
sram_cell_6t_5 inst_cell_235_61 (.BL(BL61),.BLN(BLN61),.WL(WL235));
sram_cell_6t_5 inst_cell_235_62 (.BL(BL62),.BLN(BLN62),.WL(WL235));
sram_cell_6t_5 inst_cell_235_63 (.BL(BL63),.BLN(BLN63),.WL(WL235));
sram_cell_6t_5 inst_cell_235_64 (.BL(BL64),.BLN(BLN64),.WL(WL235));
sram_cell_6t_5 inst_cell_235_65 (.BL(BL65),.BLN(BLN65),.WL(WL235));
sram_cell_6t_5 inst_cell_235_66 (.BL(BL66),.BLN(BLN66),.WL(WL235));
sram_cell_6t_5 inst_cell_235_67 (.BL(BL67),.BLN(BLN67),.WL(WL235));
sram_cell_6t_5 inst_cell_235_68 (.BL(BL68),.BLN(BLN68),.WL(WL235));
sram_cell_6t_5 inst_cell_235_69 (.BL(BL69),.BLN(BLN69),.WL(WL235));
sram_cell_6t_5 inst_cell_235_70 (.BL(BL70),.BLN(BLN70),.WL(WL235));
sram_cell_6t_5 inst_cell_235_71 (.BL(BL71),.BLN(BLN71),.WL(WL235));
sram_cell_6t_5 inst_cell_235_72 (.BL(BL72),.BLN(BLN72),.WL(WL235));
sram_cell_6t_5 inst_cell_235_73 (.BL(BL73),.BLN(BLN73),.WL(WL235));
sram_cell_6t_5 inst_cell_235_74 (.BL(BL74),.BLN(BLN74),.WL(WL235));
sram_cell_6t_5 inst_cell_235_75 (.BL(BL75),.BLN(BLN75),.WL(WL235));
sram_cell_6t_5 inst_cell_235_76 (.BL(BL76),.BLN(BLN76),.WL(WL235));
sram_cell_6t_5 inst_cell_235_77 (.BL(BL77),.BLN(BLN77),.WL(WL235));
sram_cell_6t_5 inst_cell_235_78 (.BL(BL78),.BLN(BLN78),.WL(WL235));
sram_cell_6t_5 inst_cell_235_79 (.BL(BL79),.BLN(BLN79),.WL(WL235));
sram_cell_6t_5 inst_cell_235_80 (.BL(BL80),.BLN(BLN80),.WL(WL235));
sram_cell_6t_5 inst_cell_235_81 (.BL(BL81),.BLN(BLN81),.WL(WL235));
sram_cell_6t_5 inst_cell_235_82 (.BL(BL82),.BLN(BLN82),.WL(WL235));
sram_cell_6t_5 inst_cell_235_83 (.BL(BL83),.BLN(BLN83),.WL(WL235));
sram_cell_6t_5 inst_cell_235_84 (.BL(BL84),.BLN(BLN84),.WL(WL235));
sram_cell_6t_5 inst_cell_235_85 (.BL(BL85),.BLN(BLN85),.WL(WL235));
sram_cell_6t_5 inst_cell_235_86 (.BL(BL86),.BLN(BLN86),.WL(WL235));
sram_cell_6t_5 inst_cell_235_87 (.BL(BL87),.BLN(BLN87),.WL(WL235));
sram_cell_6t_5 inst_cell_235_88 (.BL(BL88),.BLN(BLN88),.WL(WL235));
sram_cell_6t_5 inst_cell_235_89 (.BL(BL89),.BLN(BLN89),.WL(WL235));
sram_cell_6t_5 inst_cell_235_90 (.BL(BL90),.BLN(BLN90),.WL(WL235));
sram_cell_6t_5 inst_cell_235_91 (.BL(BL91),.BLN(BLN91),.WL(WL235));
sram_cell_6t_5 inst_cell_235_92 (.BL(BL92),.BLN(BLN92),.WL(WL235));
sram_cell_6t_5 inst_cell_235_93 (.BL(BL93),.BLN(BLN93),.WL(WL235));
sram_cell_6t_5 inst_cell_235_94 (.BL(BL94),.BLN(BLN94),.WL(WL235));
sram_cell_6t_5 inst_cell_235_95 (.BL(BL95),.BLN(BLN95),.WL(WL235));
sram_cell_6t_5 inst_cell_235_96 (.BL(BL96),.BLN(BLN96),.WL(WL235));
sram_cell_6t_5 inst_cell_235_97 (.BL(BL97),.BLN(BLN97),.WL(WL235));
sram_cell_6t_5 inst_cell_235_98 (.BL(BL98),.BLN(BLN98),.WL(WL235));
sram_cell_6t_5 inst_cell_235_99 (.BL(BL99),.BLN(BLN99),.WL(WL235));
sram_cell_6t_5 inst_cell_235_100 (.BL(BL100),.BLN(BLN100),.WL(WL235));
sram_cell_6t_5 inst_cell_235_101 (.BL(BL101),.BLN(BLN101),.WL(WL235));
sram_cell_6t_5 inst_cell_235_102 (.BL(BL102),.BLN(BLN102),.WL(WL235));
sram_cell_6t_5 inst_cell_235_103 (.BL(BL103),.BLN(BLN103),.WL(WL235));
sram_cell_6t_5 inst_cell_235_104 (.BL(BL104),.BLN(BLN104),.WL(WL235));
sram_cell_6t_5 inst_cell_235_105 (.BL(BL105),.BLN(BLN105),.WL(WL235));
sram_cell_6t_5 inst_cell_235_106 (.BL(BL106),.BLN(BLN106),.WL(WL235));
sram_cell_6t_5 inst_cell_235_107 (.BL(BL107),.BLN(BLN107),.WL(WL235));
sram_cell_6t_5 inst_cell_235_108 (.BL(BL108),.BLN(BLN108),.WL(WL235));
sram_cell_6t_5 inst_cell_235_109 (.BL(BL109),.BLN(BLN109),.WL(WL235));
sram_cell_6t_5 inst_cell_235_110 (.BL(BL110),.BLN(BLN110),.WL(WL235));
sram_cell_6t_5 inst_cell_235_111 (.BL(BL111),.BLN(BLN111),.WL(WL235));
sram_cell_6t_5 inst_cell_235_112 (.BL(BL112),.BLN(BLN112),.WL(WL235));
sram_cell_6t_5 inst_cell_235_113 (.BL(BL113),.BLN(BLN113),.WL(WL235));
sram_cell_6t_5 inst_cell_235_114 (.BL(BL114),.BLN(BLN114),.WL(WL235));
sram_cell_6t_5 inst_cell_235_115 (.BL(BL115),.BLN(BLN115),.WL(WL235));
sram_cell_6t_5 inst_cell_235_116 (.BL(BL116),.BLN(BLN116),.WL(WL235));
sram_cell_6t_5 inst_cell_235_117 (.BL(BL117),.BLN(BLN117),.WL(WL235));
sram_cell_6t_5 inst_cell_235_118 (.BL(BL118),.BLN(BLN118),.WL(WL235));
sram_cell_6t_5 inst_cell_235_119 (.BL(BL119),.BLN(BLN119),.WL(WL235));
sram_cell_6t_5 inst_cell_235_120 (.BL(BL120),.BLN(BLN120),.WL(WL235));
sram_cell_6t_5 inst_cell_235_121 (.BL(BL121),.BLN(BLN121),.WL(WL235));
sram_cell_6t_5 inst_cell_235_122 (.BL(BL122),.BLN(BLN122),.WL(WL235));
sram_cell_6t_5 inst_cell_235_123 (.BL(BL123),.BLN(BLN123),.WL(WL235));
sram_cell_6t_5 inst_cell_235_124 (.BL(BL124),.BLN(BLN124),.WL(WL235));
sram_cell_6t_5 inst_cell_235_125 (.BL(BL125),.BLN(BLN125),.WL(WL235));
sram_cell_6t_5 inst_cell_235_126 (.BL(BL126),.BLN(BLN126),.WL(WL235));
sram_cell_6t_5 inst_cell_235_127 (.BL(BL127),.BLN(BLN127),.WL(WL235));
sram_cell_6t_5 inst_cell_236_0 (.BL(BL0),.BLN(BLN0),.WL(WL236));
sram_cell_6t_5 inst_cell_236_1 (.BL(BL1),.BLN(BLN1),.WL(WL236));
sram_cell_6t_5 inst_cell_236_2 (.BL(BL2),.BLN(BLN2),.WL(WL236));
sram_cell_6t_5 inst_cell_236_3 (.BL(BL3),.BLN(BLN3),.WL(WL236));
sram_cell_6t_5 inst_cell_236_4 (.BL(BL4),.BLN(BLN4),.WL(WL236));
sram_cell_6t_5 inst_cell_236_5 (.BL(BL5),.BLN(BLN5),.WL(WL236));
sram_cell_6t_5 inst_cell_236_6 (.BL(BL6),.BLN(BLN6),.WL(WL236));
sram_cell_6t_5 inst_cell_236_7 (.BL(BL7),.BLN(BLN7),.WL(WL236));
sram_cell_6t_5 inst_cell_236_8 (.BL(BL8),.BLN(BLN8),.WL(WL236));
sram_cell_6t_5 inst_cell_236_9 (.BL(BL9),.BLN(BLN9),.WL(WL236));
sram_cell_6t_5 inst_cell_236_10 (.BL(BL10),.BLN(BLN10),.WL(WL236));
sram_cell_6t_5 inst_cell_236_11 (.BL(BL11),.BLN(BLN11),.WL(WL236));
sram_cell_6t_5 inst_cell_236_12 (.BL(BL12),.BLN(BLN12),.WL(WL236));
sram_cell_6t_5 inst_cell_236_13 (.BL(BL13),.BLN(BLN13),.WL(WL236));
sram_cell_6t_5 inst_cell_236_14 (.BL(BL14),.BLN(BLN14),.WL(WL236));
sram_cell_6t_5 inst_cell_236_15 (.BL(BL15),.BLN(BLN15),.WL(WL236));
sram_cell_6t_5 inst_cell_236_16 (.BL(BL16),.BLN(BLN16),.WL(WL236));
sram_cell_6t_5 inst_cell_236_17 (.BL(BL17),.BLN(BLN17),.WL(WL236));
sram_cell_6t_5 inst_cell_236_18 (.BL(BL18),.BLN(BLN18),.WL(WL236));
sram_cell_6t_5 inst_cell_236_19 (.BL(BL19),.BLN(BLN19),.WL(WL236));
sram_cell_6t_5 inst_cell_236_20 (.BL(BL20),.BLN(BLN20),.WL(WL236));
sram_cell_6t_5 inst_cell_236_21 (.BL(BL21),.BLN(BLN21),.WL(WL236));
sram_cell_6t_5 inst_cell_236_22 (.BL(BL22),.BLN(BLN22),.WL(WL236));
sram_cell_6t_5 inst_cell_236_23 (.BL(BL23),.BLN(BLN23),.WL(WL236));
sram_cell_6t_5 inst_cell_236_24 (.BL(BL24),.BLN(BLN24),.WL(WL236));
sram_cell_6t_5 inst_cell_236_25 (.BL(BL25),.BLN(BLN25),.WL(WL236));
sram_cell_6t_5 inst_cell_236_26 (.BL(BL26),.BLN(BLN26),.WL(WL236));
sram_cell_6t_5 inst_cell_236_27 (.BL(BL27),.BLN(BLN27),.WL(WL236));
sram_cell_6t_5 inst_cell_236_28 (.BL(BL28),.BLN(BLN28),.WL(WL236));
sram_cell_6t_5 inst_cell_236_29 (.BL(BL29),.BLN(BLN29),.WL(WL236));
sram_cell_6t_5 inst_cell_236_30 (.BL(BL30),.BLN(BLN30),.WL(WL236));
sram_cell_6t_5 inst_cell_236_31 (.BL(BL31),.BLN(BLN31),.WL(WL236));
sram_cell_6t_5 inst_cell_236_32 (.BL(BL32),.BLN(BLN32),.WL(WL236));
sram_cell_6t_5 inst_cell_236_33 (.BL(BL33),.BLN(BLN33),.WL(WL236));
sram_cell_6t_5 inst_cell_236_34 (.BL(BL34),.BLN(BLN34),.WL(WL236));
sram_cell_6t_5 inst_cell_236_35 (.BL(BL35),.BLN(BLN35),.WL(WL236));
sram_cell_6t_5 inst_cell_236_36 (.BL(BL36),.BLN(BLN36),.WL(WL236));
sram_cell_6t_5 inst_cell_236_37 (.BL(BL37),.BLN(BLN37),.WL(WL236));
sram_cell_6t_5 inst_cell_236_38 (.BL(BL38),.BLN(BLN38),.WL(WL236));
sram_cell_6t_5 inst_cell_236_39 (.BL(BL39),.BLN(BLN39),.WL(WL236));
sram_cell_6t_5 inst_cell_236_40 (.BL(BL40),.BLN(BLN40),.WL(WL236));
sram_cell_6t_5 inst_cell_236_41 (.BL(BL41),.BLN(BLN41),.WL(WL236));
sram_cell_6t_5 inst_cell_236_42 (.BL(BL42),.BLN(BLN42),.WL(WL236));
sram_cell_6t_5 inst_cell_236_43 (.BL(BL43),.BLN(BLN43),.WL(WL236));
sram_cell_6t_5 inst_cell_236_44 (.BL(BL44),.BLN(BLN44),.WL(WL236));
sram_cell_6t_5 inst_cell_236_45 (.BL(BL45),.BLN(BLN45),.WL(WL236));
sram_cell_6t_5 inst_cell_236_46 (.BL(BL46),.BLN(BLN46),.WL(WL236));
sram_cell_6t_5 inst_cell_236_47 (.BL(BL47),.BLN(BLN47),.WL(WL236));
sram_cell_6t_5 inst_cell_236_48 (.BL(BL48),.BLN(BLN48),.WL(WL236));
sram_cell_6t_5 inst_cell_236_49 (.BL(BL49),.BLN(BLN49),.WL(WL236));
sram_cell_6t_5 inst_cell_236_50 (.BL(BL50),.BLN(BLN50),.WL(WL236));
sram_cell_6t_5 inst_cell_236_51 (.BL(BL51),.BLN(BLN51),.WL(WL236));
sram_cell_6t_5 inst_cell_236_52 (.BL(BL52),.BLN(BLN52),.WL(WL236));
sram_cell_6t_5 inst_cell_236_53 (.BL(BL53),.BLN(BLN53),.WL(WL236));
sram_cell_6t_5 inst_cell_236_54 (.BL(BL54),.BLN(BLN54),.WL(WL236));
sram_cell_6t_5 inst_cell_236_55 (.BL(BL55),.BLN(BLN55),.WL(WL236));
sram_cell_6t_5 inst_cell_236_56 (.BL(BL56),.BLN(BLN56),.WL(WL236));
sram_cell_6t_5 inst_cell_236_57 (.BL(BL57),.BLN(BLN57),.WL(WL236));
sram_cell_6t_5 inst_cell_236_58 (.BL(BL58),.BLN(BLN58),.WL(WL236));
sram_cell_6t_5 inst_cell_236_59 (.BL(BL59),.BLN(BLN59),.WL(WL236));
sram_cell_6t_5 inst_cell_236_60 (.BL(BL60),.BLN(BLN60),.WL(WL236));
sram_cell_6t_5 inst_cell_236_61 (.BL(BL61),.BLN(BLN61),.WL(WL236));
sram_cell_6t_5 inst_cell_236_62 (.BL(BL62),.BLN(BLN62),.WL(WL236));
sram_cell_6t_5 inst_cell_236_63 (.BL(BL63),.BLN(BLN63),.WL(WL236));
sram_cell_6t_5 inst_cell_236_64 (.BL(BL64),.BLN(BLN64),.WL(WL236));
sram_cell_6t_5 inst_cell_236_65 (.BL(BL65),.BLN(BLN65),.WL(WL236));
sram_cell_6t_5 inst_cell_236_66 (.BL(BL66),.BLN(BLN66),.WL(WL236));
sram_cell_6t_5 inst_cell_236_67 (.BL(BL67),.BLN(BLN67),.WL(WL236));
sram_cell_6t_5 inst_cell_236_68 (.BL(BL68),.BLN(BLN68),.WL(WL236));
sram_cell_6t_5 inst_cell_236_69 (.BL(BL69),.BLN(BLN69),.WL(WL236));
sram_cell_6t_5 inst_cell_236_70 (.BL(BL70),.BLN(BLN70),.WL(WL236));
sram_cell_6t_5 inst_cell_236_71 (.BL(BL71),.BLN(BLN71),.WL(WL236));
sram_cell_6t_5 inst_cell_236_72 (.BL(BL72),.BLN(BLN72),.WL(WL236));
sram_cell_6t_5 inst_cell_236_73 (.BL(BL73),.BLN(BLN73),.WL(WL236));
sram_cell_6t_5 inst_cell_236_74 (.BL(BL74),.BLN(BLN74),.WL(WL236));
sram_cell_6t_5 inst_cell_236_75 (.BL(BL75),.BLN(BLN75),.WL(WL236));
sram_cell_6t_5 inst_cell_236_76 (.BL(BL76),.BLN(BLN76),.WL(WL236));
sram_cell_6t_5 inst_cell_236_77 (.BL(BL77),.BLN(BLN77),.WL(WL236));
sram_cell_6t_5 inst_cell_236_78 (.BL(BL78),.BLN(BLN78),.WL(WL236));
sram_cell_6t_5 inst_cell_236_79 (.BL(BL79),.BLN(BLN79),.WL(WL236));
sram_cell_6t_5 inst_cell_236_80 (.BL(BL80),.BLN(BLN80),.WL(WL236));
sram_cell_6t_5 inst_cell_236_81 (.BL(BL81),.BLN(BLN81),.WL(WL236));
sram_cell_6t_5 inst_cell_236_82 (.BL(BL82),.BLN(BLN82),.WL(WL236));
sram_cell_6t_5 inst_cell_236_83 (.BL(BL83),.BLN(BLN83),.WL(WL236));
sram_cell_6t_5 inst_cell_236_84 (.BL(BL84),.BLN(BLN84),.WL(WL236));
sram_cell_6t_5 inst_cell_236_85 (.BL(BL85),.BLN(BLN85),.WL(WL236));
sram_cell_6t_5 inst_cell_236_86 (.BL(BL86),.BLN(BLN86),.WL(WL236));
sram_cell_6t_5 inst_cell_236_87 (.BL(BL87),.BLN(BLN87),.WL(WL236));
sram_cell_6t_5 inst_cell_236_88 (.BL(BL88),.BLN(BLN88),.WL(WL236));
sram_cell_6t_5 inst_cell_236_89 (.BL(BL89),.BLN(BLN89),.WL(WL236));
sram_cell_6t_5 inst_cell_236_90 (.BL(BL90),.BLN(BLN90),.WL(WL236));
sram_cell_6t_5 inst_cell_236_91 (.BL(BL91),.BLN(BLN91),.WL(WL236));
sram_cell_6t_5 inst_cell_236_92 (.BL(BL92),.BLN(BLN92),.WL(WL236));
sram_cell_6t_5 inst_cell_236_93 (.BL(BL93),.BLN(BLN93),.WL(WL236));
sram_cell_6t_5 inst_cell_236_94 (.BL(BL94),.BLN(BLN94),.WL(WL236));
sram_cell_6t_5 inst_cell_236_95 (.BL(BL95),.BLN(BLN95),.WL(WL236));
sram_cell_6t_5 inst_cell_236_96 (.BL(BL96),.BLN(BLN96),.WL(WL236));
sram_cell_6t_5 inst_cell_236_97 (.BL(BL97),.BLN(BLN97),.WL(WL236));
sram_cell_6t_5 inst_cell_236_98 (.BL(BL98),.BLN(BLN98),.WL(WL236));
sram_cell_6t_5 inst_cell_236_99 (.BL(BL99),.BLN(BLN99),.WL(WL236));
sram_cell_6t_5 inst_cell_236_100 (.BL(BL100),.BLN(BLN100),.WL(WL236));
sram_cell_6t_5 inst_cell_236_101 (.BL(BL101),.BLN(BLN101),.WL(WL236));
sram_cell_6t_5 inst_cell_236_102 (.BL(BL102),.BLN(BLN102),.WL(WL236));
sram_cell_6t_5 inst_cell_236_103 (.BL(BL103),.BLN(BLN103),.WL(WL236));
sram_cell_6t_5 inst_cell_236_104 (.BL(BL104),.BLN(BLN104),.WL(WL236));
sram_cell_6t_5 inst_cell_236_105 (.BL(BL105),.BLN(BLN105),.WL(WL236));
sram_cell_6t_5 inst_cell_236_106 (.BL(BL106),.BLN(BLN106),.WL(WL236));
sram_cell_6t_5 inst_cell_236_107 (.BL(BL107),.BLN(BLN107),.WL(WL236));
sram_cell_6t_5 inst_cell_236_108 (.BL(BL108),.BLN(BLN108),.WL(WL236));
sram_cell_6t_5 inst_cell_236_109 (.BL(BL109),.BLN(BLN109),.WL(WL236));
sram_cell_6t_5 inst_cell_236_110 (.BL(BL110),.BLN(BLN110),.WL(WL236));
sram_cell_6t_5 inst_cell_236_111 (.BL(BL111),.BLN(BLN111),.WL(WL236));
sram_cell_6t_5 inst_cell_236_112 (.BL(BL112),.BLN(BLN112),.WL(WL236));
sram_cell_6t_5 inst_cell_236_113 (.BL(BL113),.BLN(BLN113),.WL(WL236));
sram_cell_6t_5 inst_cell_236_114 (.BL(BL114),.BLN(BLN114),.WL(WL236));
sram_cell_6t_5 inst_cell_236_115 (.BL(BL115),.BLN(BLN115),.WL(WL236));
sram_cell_6t_5 inst_cell_236_116 (.BL(BL116),.BLN(BLN116),.WL(WL236));
sram_cell_6t_5 inst_cell_236_117 (.BL(BL117),.BLN(BLN117),.WL(WL236));
sram_cell_6t_5 inst_cell_236_118 (.BL(BL118),.BLN(BLN118),.WL(WL236));
sram_cell_6t_5 inst_cell_236_119 (.BL(BL119),.BLN(BLN119),.WL(WL236));
sram_cell_6t_5 inst_cell_236_120 (.BL(BL120),.BLN(BLN120),.WL(WL236));
sram_cell_6t_5 inst_cell_236_121 (.BL(BL121),.BLN(BLN121),.WL(WL236));
sram_cell_6t_5 inst_cell_236_122 (.BL(BL122),.BLN(BLN122),.WL(WL236));
sram_cell_6t_5 inst_cell_236_123 (.BL(BL123),.BLN(BLN123),.WL(WL236));
sram_cell_6t_5 inst_cell_236_124 (.BL(BL124),.BLN(BLN124),.WL(WL236));
sram_cell_6t_5 inst_cell_236_125 (.BL(BL125),.BLN(BLN125),.WL(WL236));
sram_cell_6t_5 inst_cell_236_126 (.BL(BL126),.BLN(BLN126),.WL(WL236));
sram_cell_6t_5 inst_cell_236_127 (.BL(BL127),.BLN(BLN127),.WL(WL236));
sram_cell_6t_5 inst_cell_237_0 (.BL(BL0),.BLN(BLN0),.WL(WL237));
sram_cell_6t_5 inst_cell_237_1 (.BL(BL1),.BLN(BLN1),.WL(WL237));
sram_cell_6t_5 inst_cell_237_2 (.BL(BL2),.BLN(BLN2),.WL(WL237));
sram_cell_6t_5 inst_cell_237_3 (.BL(BL3),.BLN(BLN3),.WL(WL237));
sram_cell_6t_5 inst_cell_237_4 (.BL(BL4),.BLN(BLN4),.WL(WL237));
sram_cell_6t_5 inst_cell_237_5 (.BL(BL5),.BLN(BLN5),.WL(WL237));
sram_cell_6t_5 inst_cell_237_6 (.BL(BL6),.BLN(BLN6),.WL(WL237));
sram_cell_6t_5 inst_cell_237_7 (.BL(BL7),.BLN(BLN7),.WL(WL237));
sram_cell_6t_5 inst_cell_237_8 (.BL(BL8),.BLN(BLN8),.WL(WL237));
sram_cell_6t_5 inst_cell_237_9 (.BL(BL9),.BLN(BLN9),.WL(WL237));
sram_cell_6t_5 inst_cell_237_10 (.BL(BL10),.BLN(BLN10),.WL(WL237));
sram_cell_6t_5 inst_cell_237_11 (.BL(BL11),.BLN(BLN11),.WL(WL237));
sram_cell_6t_5 inst_cell_237_12 (.BL(BL12),.BLN(BLN12),.WL(WL237));
sram_cell_6t_5 inst_cell_237_13 (.BL(BL13),.BLN(BLN13),.WL(WL237));
sram_cell_6t_5 inst_cell_237_14 (.BL(BL14),.BLN(BLN14),.WL(WL237));
sram_cell_6t_5 inst_cell_237_15 (.BL(BL15),.BLN(BLN15),.WL(WL237));
sram_cell_6t_5 inst_cell_237_16 (.BL(BL16),.BLN(BLN16),.WL(WL237));
sram_cell_6t_5 inst_cell_237_17 (.BL(BL17),.BLN(BLN17),.WL(WL237));
sram_cell_6t_5 inst_cell_237_18 (.BL(BL18),.BLN(BLN18),.WL(WL237));
sram_cell_6t_5 inst_cell_237_19 (.BL(BL19),.BLN(BLN19),.WL(WL237));
sram_cell_6t_5 inst_cell_237_20 (.BL(BL20),.BLN(BLN20),.WL(WL237));
sram_cell_6t_5 inst_cell_237_21 (.BL(BL21),.BLN(BLN21),.WL(WL237));
sram_cell_6t_5 inst_cell_237_22 (.BL(BL22),.BLN(BLN22),.WL(WL237));
sram_cell_6t_5 inst_cell_237_23 (.BL(BL23),.BLN(BLN23),.WL(WL237));
sram_cell_6t_5 inst_cell_237_24 (.BL(BL24),.BLN(BLN24),.WL(WL237));
sram_cell_6t_5 inst_cell_237_25 (.BL(BL25),.BLN(BLN25),.WL(WL237));
sram_cell_6t_5 inst_cell_237_26 (.BL(BL26),.BLN(BLN26),.WL(WL237));
sram_cell_6t_5 inst_cell_237_27 (.BL(BL27),.BLN(BLN27),.WL(WL237));
sram_cell_6t_5 inst_cell_237_28 (.BL(BL28),.BLN(BLN28),.WL(WL237));
sram_cell_6t_5 inst_cell_237_29 (.BL(BL29),.BLN(BLN29),.WL(WL237));
sram_cell_6t_5 inst_cell_237_30 (.BL(BL30),.BLN(BLN30),.WL(WL237));
sram_cell_6t_5 inst_cell_237_31 (.BL(BL31),.BLN(BLN31),.WL(WL237));
sram_cell_6t_5 inst_cell_237_32 (.BL(BL32),.BLN(BLN32),.WL(WL237));
sram_cell_6t_5 inst_cell_237_33 (.BL(BL33),.BLN(BLN33),.WL(WL237));
sram_cell_6t_5 inst_cell_237_34 (.BL(BL34),.BLN(BLN34),.WL(WL237));
sram_cell_6t_5 inst_cell_237_35 (.BL(BL35),.BLN(BLN35),.WL(WL237));
sram_cell_6t_5 inst_cell_237_36 (.BL(BL36),.BLN(BLN36),.WL(WL237));
sram_cell_6t_5 inst_cell_237_37 (.BL(BL37),.BLN(BLN37),.WL(WL237));
sram_cell_6t_5 inst_cell_237_38 (.BL(BL38),.BLN(BLN38),.WL(WL237));
sram_cell_6t_5 inst_cell_237_39 (.BL(BL39),.BLN(BLN39),.WL(WL237));
sram_cell_6t_5 inst_cell_237_40 (.BL(BL40),.BLN(BLN40),.WL(WL237));
sram_cell_6t_5 inst_cell_237_41 (.BL(BL41),.BLN(BLN41),.WL(WL237));
sram_cell_6t_5 inst_cell_237_42 (.BL(BL42),.BLN(BLN42),.WL(WL237));
sram_cell_6t_5 inst_cell_237_43 (.BL(BL43),.BLN(BLN43),.WL(WL237));
sram_cell_6t_5 inst_cell_237_44 (.BL(BL44),.BLN(BLN44),.WL(WL237));
sram_cell_6t_5 inst_cell_237_45 (.BL(BL45),.BLN(BLN45),.WL(WL237));
sram_cell_6t_5 inst_cell_237_46 (.BL(BL46),.BLN(BLN46),.WL(WL237));
sram_cell_6t_5 inst_cell_237_47 (.BL(BL47),.BLN(BLN47),.WL(WL237));
sram_cell_6t_5 inst_cell_237_48 (.BL(BL48),.BLN(BLN48),.WL(WL237));
sram_cell_6t_5 inst_cell_237_49 (.BL(BL49),.BLN(BLN49),.WL(WL237));
sram_cell_6t_5 inst_cell_237_50 (.BL(BL50),.BLN(BLN50),.WL(WL237));
sram_cell_6t_5 inst_cell_237_51 (.BL(BL51),.BLN(BLN51),.WL(WL237));
sram_cell_6t_5 inst_cell_237_52 (.BL(BL52),.BLN(BLN52),.WL(WL237));
sram_cell_6t_5 inst_cell_237_53 (.BL(BL53),.BLN(BLN53),.WL(WL237));
sram_cell_6t_5 inst_cell_237_54 (.BL(BL54),.BLN(BLN54),.WL(WL237));
sram_cell_6t_5 inst_cell_237_55 (.BL(BL55),.BLN(BLN55),.WL(WL237));
sram_cell_6t_5 inst_cell_237_56 (.BL(BL56),.BLN(BLN56),.WL(WL237));
sram_cell_6t_5 inst_cell_237_57 (.BL(BL57),.BLN(BLN57),.WL(WL237));
sram_cell_6t_5 inst_cell_237_58 (.BL(BL58),.BLN(BLN58),.WL(WL237));
sram_cell_6t_5 inst_cell_237_59 (.BL(BL59),.BLN(BLN59),.WL(WL237));
sram_cell_6t_5 inst_cell_237_60 (.BL(BL60),.BLN(BLN60),.WL(WL237));
sram_cell_6t_5 inst_cell_237_61 (.BL(BL61),.BLN(BLN61),.WL(WL237));
sram_cell_6t_5 inst_cell_237_62 (.BL(BL62),.BLN(BLN62),.WL(WL237));
sram_cell_6t_5 inst_cell_237_63 (.BL(BL63),.BLN(BLN63),.WL(WL237));
sram_cell_6t_5 inst_cell_237_64 (.BL(BL64),.BLN(BLN64),.WL(WL237));
sram_cell_6t_5 inst_cell_237_65 (.BL(BL65),.BLN(BLN65),.WL(WL237));
sram_cell_6t_5 inst_cell_237_66 (.BL(BL66),.BLN(BLN66),.WL(WL237));
sram_cell_6t_5 inst_cell_237_67 (.BL(BL67),.BLN(BLN67),.WL(WL237));
sram_cell_6t_5 inst_cell_237_68 (.BL(BL68),.BLN(BLN68),.WL(WL237));
sram_cell_6t_5 inst_cell_237_69 (.BL(BL69),.BLN(BLN69),.WL(WL237));
sram_cell_6t_5 inst_cell_237_70 (.BL(BL70),.BLN(BLN70),.WL(WL237));
sram_cell_6t_5 inst_cell_237_71 (.BL(BL71),.BLN(BLN71),.WL(WL237));
sram_cell_6t_5 inst_cell_237_72 (.BL(BL72),.BLN(BLN72),.WL(WL237));
sram_cell_6t_5 inst_cell_237_73 (.BL(BL73),.BLN(BLN73),.WL(WL237));
sram_cell_6t_5 inst_cell_237_74 (.BL(BL74),.BLN(BLN74),.WL(WL237));
sram_cell_6t_5 inst_cell_237_75 (.BL(BL75),.BLN(BLN75),.WL(WL237));
sram_cell_6t_5 inst_cell_237_76 (.BL(BL76),.BLN(BLN76),.WL(WL237));
sram_cell_6t_5 inst_cell_237_77 (.BL(BL77),.BLN(BLN77),.WL(WL237));
sram_cell_6t_5 inst_cell_237_78 (.BL(BL78),.BLN(BLN78),.WL(WL237));
sram_cell_6t_5 inst_cell_237_79 (.BL(BL79),.BLN(BLN79),.WL(WL237));
sram_cell_6t_5 inst_cell_237_80 (.BL(BL80),.BLN(BLN80),.WL(WL237));
sram_cell_6t_5 inst_cell_237_81 (.BL(BL81),.BLN(BLN81),.WL(WL237));
sram_cell_6t_5 inst_cell_237_82 (.BL(BL82),.BLN(BLN82),.WL(WL237));
sram_cell_6t_5 inst_cell_237_83 (.BL(BL83),.BLN(BLN83),.WL(WL237));
sram_cell_6t_5 inst_cell_237_84 (.BL(BL84),.BLN(BLN84),.WL(WL237));
sram_cell_6t_5 inst_cell_237_85 (.BL(BL85),.BLN(BLN85),.WL(WL237));
sram_cell_6t_5 inst_cell_237_86 (.BL(BL86),.BLN(BLN86),.WL(WL237));
sram_cell_6t_5 inst_cell_237_87 (.BL(BL87),.BLN(BLN87),.WL(WL237));
sram_cell_6t_5 inst_cell_237_88 (.BL(BL88),.BLN(BLN88),.WL(WL237));
sram_cell_6t_5 inst_cell_237_89 (.BL(BL89),.BLN(BLN89),.WL(WL237));
sram_cell_6t_5 inst_cell_237_90 (.BL(BL90),.BLN(BLN90),.WL(WL237));
sram_cell_6t_5 inst_cell_237_91 (.BL(BL91),.BLN(BLN91),.WL(WL237));
sram_cell_6t_5 inst_cell_237_92 (.BL(BL92),.BLN(BLN92),.WL(WL237));
sram_cell_6t_5 inst_cell_237_93 (.BL(BL93),.BLN(BLN93),.WL(WL237));
sram_cell_6t_5 inst_cell_237_94 (.BL(BL94),.BLN(BLN94),.WL(WL237));
sram_cell_6t_5 inst_cell_237_95 (.BL(BL95),.BLN(BLN95),.WL(WL237));
sram_cell_6t_5 inst_cell_237_96 (.BL(BL96),.BLN(BLN96),.WL(WL237));
sram_cell_6t_5 inst_cell_237_97 (.BL(BL97),.BLN(BLN97),.WL(WL237));
sram_cell_6t_5 inst_cell_237_98 (.BL(BL98),.BLN(BLN98),.WL(WL237));
sram_cell_6t_5 inst_cell_237_99 (.BL(BL99),.BLN(BLN99),.WL(WL237));
sram_cell_6t_5 inst_cell_237_100 (.BL(BL100),.BLN(BLN100),.WL(WL237));
sram_cell_6t_5 inst_cell_237_101 (.BL(BL101),.BLN(BLN101),.WL(WL237));
sram_cell_6t_5 inst_cell_237_102 (.BL(BL102),.BLN(BLN102),.WL(WL237));
sram_cell_6t_5 inst_cell_237_103 (.BL(BL103),.BLN(BLN103),.WL(WL237));
sram_cell_6t_5 inst_cell_237_104 (.BL(BL104),.BLN(BLN104),.WL(WL237));
sram_cell_6t_5 inst_cell_237_105 (.BL(BL105),.BLN(BLN105),.WL(WL237));
sram_cell_6t_5 inst_cell_237_106 (.BL(BL106),.BLN(BLN106),.WL(WL237));
sram_cell_6t_5 inst_cell_237_107 (.BL(BL107),.BLN(BLN107),.WL(WL237));
sram_cell_6t_5 inst_cell_237_108 (.BL(BL108),.BLN(BLN108),.WL(WL237));
sram_cell_6t_5 inst_cell_237_109 (.BL(BL109),.BLN(BLN109),.WL(WL237));
sram_cell_6t_5 inst_cell_237_110 (.BL(BL110),.BLN(BLN110),.WL(WL237));
sram_cell_6t_5 inst_cell_237_111 (.BL(BL111),.BLN(BLN111),.WL(WL237));
sram_cell_6t_5 inst_cell_237_112 (.BL(BL112),.BLN(BLN112),.WL(WL237));
sram_cell_6t_5 inst_cell_237_113 (.BL(BL113),.BLN(BLN113),.WL(WL237));
sram_cell_6t_5 inst_cell_237_114 (.BL(BL114),.BLN(BLN114),.WL(WL237));
sram_cell_6t_5 inst_cell_237_115 (.BL(BL115),.BLN(BLN115),.WL(WL237));
sram_cell_6t_5 inst_cell_237_116 (.BL(BL116),.BLN(BLN116),.WL(WL237));
sram_cell_6t_5 inst_cell_237_117 (.BL(BL117),.BLN(BLN117),.WL(WL237));
sram_cell_6t_5 inst_cell_237_118 (.BL(BL118),.BLN(BLN118),.WL(WL237));
sram_cell_6t_5 inst_cell_237_119 (.BL(BL119),.BLN(BLN119),.WL(WL237));
sram_cell_6t_5 inst_cell_237_120 (.BL(BL120),.BLN(BLN120),.WL(WL237));
sram_cell_6t_5 inst_cell_237_121 (.BL(BL121),.BLN(BLN121),.WL(WL237));
sram_cell_6t_5 inst_cell_237_122 (.BL(BL122),.BLN(BLN122),.WL(WL237));
sram_cell_6t_5 inst_cell_237_123 (.BL(BL123),.BLN(BLN123),.WL(WL237));
sram_cell_6t_5 inst_cell_237_124 (.BL(BL124),.BLN(BLN124),.WL(WL237));
sram_cell_6t_5 inst_cell_237_125 (.BL(BL125),.BLN(BLN125),.WL(WL237));
sram_cell_6t_5 inst_cell_237_126 (.BL(BL126),.BLN(BLN126),.WL(WL237));
sram_cell_6t_5 inst_cell_237_127 (.BL(BL127),.BLN(BLN127),.WL(WL237));
sram_cell_6t_5 inst_cell_238_0 (.BL(BL0),.BLN(BLN0),.WL(WL238));
sram_cell_6t_5 inst_cell_238_1 (.BL(BL1),.BLN(BLN1),.WL(WL238));
sram_cell_6t_5 inst_cell_238_2 (.BL(BL2),.BLN(BLN2),.WL(WL238));
sram_cell_6t_5 inst_cell_238_3 (.BL(BL3),.BLN(BLN3),.WL(WL238));
sram_cell_6t_5 inst_cell_238_4 (.BL(BL4),.BLN(BLN4),.WL(WL238));
sram_cell_6t_5 inst_cell_238_5 (.BL(BL5),.BLN(BLN5),.WL(WL238));
sram_cell_6t_5 inst_cell_238_6 (.BL(BL6),.BLN(BLN6),.WL(WL238));
sram_cell_6t_5 inst_cell_238_7 (.BL(BL7),.BLN(BLN7),.WL(WL238));
sram_cell_6t_5 inst_cell_238_8 (.BL(BL8),.BLN(BLN8),.WL(WL238));
sram_cell_6t_5 inst_cell_238_9 (.BL(BL9),.BLN(BLN9),.WL(WL238));
sram_cell_6t_5 inst_cell_238_10 (.BL(BL10),.BLN(BLN10),.WL(WL238));
sram_cell_6t_5 inst_cell_238_11 (.BL(BL11),.BLN(BLN11),.WL(WL238));
sram_cell_6t_5 inst_cell_238_12 (.BL(BL12),.BLN(BLN12),.WL(WL238));
sram_cell_6t_5 inst_cell_238_13 (.BL(BL13),.BLN(BLN13),.WL(WL238));
sram_cell_6t_5 inst_cell_238_14 (.BL(BL14),.BLN(BLN14),.WL(WL238));
sram_cell_6t_5 inst_cell_238_15 (.BL(BL15),.BLN(BLN15),.WL(WL238));
sram_cell_6t_5 inst_cell_238_16 (.BL(BL16),.BLN(BLN16),.WL(WL238));
sram_cell_6t_5 inst_cell_238_17 (.BL(BL17),.BLN(BLN17),.WL(WL238));
sram_cell_6t_5 inst_cell_238_18 (.BL(BL18),.BLN(BLN18),.WL(WL238));
sram_cell_6t_5 inst_cell_238_19 (.BL(BL19),.BLN(BLN19),.WL(WL238));
sram_cell_6t_5 inst_cell_238_20 (.BL(BL20),.BLN(BLN20),.WL(WL238));
sram_cell_6t_5 inst_cell_238_21 (.BL(BL21),.BLN(BLN21),.WL(WL238));
sram_cell_6t_5 inst_cell_238_22 (.BL(BL22),.BLN(BLN22),.WL(WL238));
sram_cell_6t_5 inst_cell_238_23 (.BL(BL23),.BLN(BLN23),.WL(WL238));
sram_cell_6t_5 inst_cell_238_24 (.BL(BL24),.BLN(BLN24),.WL(WL238));
sram_cell_6t_5 inst_cell_238_25 (.BL(BL25),.BLN(BLN25),.WL(WL238));
sram_cell_6t_5 inst_cell_238_26 (.BL(BL26),.BLN(BLN26),.WL(WL238));
sram_cell_6t_5 inst_cell_238_27 (.BL(BL27),.BLN(BLN27),.WL(WL238));
sram_cell_6t_5 inst_cell_238_28 (.BL(BL28),.BLN(BLN28),.WL(WL238));
sram_cell_6t_5 inst_cell_238_29 (.BL(BL29),.BLN(BLN29),.WL(WL238));
sram_cell_6t_5 inst_cell_238_30 (.BL(BL30),.BLN(BLN30),.WL(WL238));
sram_cell_6t_5 inst_cell_238_31 (.BL(BL31),.BLN(BLN31),.WL(WL238));
sram_cell_6t_5 inst_cell_238_32 (.BL(BL32),.BLN(BLN32),.WL(WL238));
sram_cell_6t_5 inst_cell_238_33 (.BL(BL33),.BLN(BLN33),.WL(WL238));
sram_cell_6t_5 inst_cell_238_34 (.BL(BL34),.BLN(BLN34),.WL(WL238));
sram_cell_6t_5 inst_cell_238_35 (.BL(BL35),.BLN(BLN35),.WL(WL238));
sram_cell_6t_5 inst_cell_238_36 (.BL(BL36),.BLN(BLN36),.WL(WL238));
sram_cell_6t_5 inst_cell_238_37 (.BL(BL37),.BLN(BLN37),.WL(WL238));
sram_cell_6t_5 inst_cell_238_38 (.BL(BL38),.BLN(BLN38),.WL(WL238));
sram_cell_6t_5 inst_cell_238_39 (.BL(BL39),.BLN(BLN39),.WL(WL238));
sram_cell_6t_5 inst_cell_238_40 (.BL(BL40),.BLN(BLN40),.WL(WL238));
sram_cell_6t_5 inst_cell_238_41 (.BL(BL41),.BLN(BLN41),.WL(WL238));
sram_cell_6t_5 inst_cell_238_42 (.BL(BL42),.BLN(BLN42),.WL(WL238));
sram_cell_6t_5 inst_cell_238_43 (.BL(BL43),.BLN(BLN43),.WL(WL238));
sram_cell_6t_5 inst_cell_238_44 (.BL(BL44),.BLN(BLN44),.WL(WL238));
sram_cell_6t_5 inst_cell_238_45 (.BL(BL45),.BLN(BLN45),.WL(WL238));
sram_cell_6t_5 inst_cell_238_46 (.BL(BL46),.BLN(BLN46),.WL(WL238));
sram_cell_6t_5 inst_cell_238_47 (.BL(BL47),.BLN(BLN47),.WL(WL238));
sram_cell_6t_5 inst_cell_238_48 (.BL(BL48),.BLN(BLN48),.WL(WL238));
sram_cell_6t_5 inst_cell_238_49 (.BL(BL49),.BLN(BLN49),.WL(WL238));
sram_cell_6t_5 inst_cell_238_50 (.BL(BL50),.BLN(BLN50),.WL(WL238));
sram_cell_6t_5 inst_cell_238_51 (.BL(BL51),.BLN(BLN51),.WL(WL238));
sram_cell_6t_5 inst_cell_238_52 (.BL(BL52),.BLN(BLN52),.WL(WL238));
sram_cell_6t_5 inst_cell_238_53 (.BL(BL53),.BLN(BLN53),.WL(WL238));
sram_cell_6t_5 inst_cell_238_54 (.BL(BL54),.BLN(BLN54),.WL(WL238));
sram_cell_6t_5 inst_cell_238_55 (.BL(BL55),.BLN(BLN55),.WL(WL238));
sram_cell_6t_5 inst_cell_238_56 (.BL(BL56),.BLN(BLN56),.WL(WL238));
sram_cell_6t_5 inst_cell_238_57 (.BL(BL57),.BLN(BLN57),.WL(WL238));
sram_cell_6t_5 inst_cell_238_58 (.BL(BL58),.BLN(BLN58),.WL(WL238));
sram_cell_6t_5 inst_cell_238_59 (.BL(BL59),.BLN(BLN59),.WL(WL238));
sram_cell_6t_5 inst_cell_238_60 (.BL(BL60),.BLN(BLN60),.WL(WL238));
sram_cell_6t_5 inst_cell_238_61 (.BL(BL61),.BLN(BLN61),.WL(WL238));
sram_cell_6t_5 inst_cell_238_62 (.BL(BL62),.BLN(BLN62),.WL(WL238));
sram_cell_6t_5 inst_cell_238_63 (.BL(BL63),.BLN(BLN63),.WL(WL238));
sram_cell_6t_5 inst_cell_238_64 (.BL(BL64),.BLN(BLN64),.WL(WL238));
sram_cell_6t_5 inst_cell_238_65 (.BL(BL65),.BLN(BLN65),.WL(WL238));
sram_cell_6t_5 inst_cell_238_66 (.BL(BL66),.BLN(BLN66),.WL(WL238));
sram_cell_6t_5 inst_cell_238_67 (.BL(BL67),.BLN(BLN67),.WL(WL238));
sram_cell_6t_5 inst_cell_238_68 (.BL(BL68),.BLN(BLN68),.WL(WL238));
sram_cell_6t_5 inst_cell_238_69 (.BL(BL69),.BLN(BLN69),.WL(WL238));
sram_cell_6t_5 inst_cell_238_70 (.BL(BL70),.BLN(BLN70),.WL(WL238));
sram_cell_6t_5 inst_cell_238_71 (.BL(BL71),.BLN(BLN71),.WL(WL238));
sram_cell_6t_5 inst_cell_238_72 (.BL(BL72),.BLN(BLN72),.WL(WL238));
sram_cell_6t_5 inst_cell_238_73 (.BL(BL73),.BLN(BLN73),.WL(WL238));
sram_cell_6t_5 inst_cell_238_74 (.BL(BL74),.BLN(BLN74),.WL(WL238));
sram_cell_6t_5 inst_cell_238_75 (.BL(BL75),.BLN(BLN75),.WL(WL238));
sram_cell_6t_5 inst_cell_238_76 (.BL(BL76),.BLN(BLN76),.WL(WL238));
sram_cell_6t_5 inst_cell_238_77 (.BL(BL77),.BLN(BLN77),.WL(WL238));
sram_cell_6t_5 inst_cell_238_78 (.BL(BL78),.BLN(BLN78),.WL(WL238));
sram_cell_6t_5 inst_cell_238_79 (.BL(BL79),.BLN(BLN79),.WL(WL238));
sram_cell_6t_5 inst_cell_238_80 (.BL(BL80),.BLN(BLN80),.WL(WL238));
sram_cell_6t_5 inst_cell_238_81 (.BL(BL81),.BLN(BLN81),.WL(WL238));
sram_cell_6t_5 inst_cell_238_82 (.BL(BL82),.BLN(BLN82),.WL(WL238));
sram_cell_6t_5 inst_cell_238_83 (.BL(BL83),.BLN(BLN83),.WL(WL238));
sram_cell_6t_5 inst_cell_238_84 (.BL(BL84),.BLN(BLN84),.WL(WL238));
sram_cell_6t_5 inst_cell_238_85 (.BL(BL85),.BLN(BLN85),.WL(WL238));
sram_cell_6t_5 inst_cell_238_86 (.BL(BL86),.BLN(BLN86),.WL(WL238));
sram_cell_6t_5 inst_cell_238_87 (.BL(BL87),.BLN(BLN87),.WL(WL238));
sram_cell_6t_5 inst_cell_238_88 (.BL(BL88),.BLN(BLN88),.WL(WL238));
sram_cell_6t_5 inst_cell_238_89 (.BL(BL89),.BLN(BLN89),.WL(WL238));
sram_cell_6t_5 inst_cell_238_90 (.BL(BL90),.BLN(BLN90),.WL(WL238));
sram_cell_6t_5 inst_cell_238_91 (.BL(BL91),.BLN(BLN91),.WL(WL238));
sram_cell_6t_5 inst_cell_238_92 (.BL(BL92),.BLN(BLN92),.WL(WL238));
sram_cell_6t_5 inst_cell_238_93 (.BL(BL93),.BLN(BLN93),.WL(WL238));
sram_cell_6t_5 inst_cell_238_94 (.BL(BL94),.BLN(BLN94),.WL(WL238));
sram_cell_6t_5 inst_cell_238_95 (.BL(BL95),.BLN(BLN95),.WL(WL238));
sram_cell_6t_5 inst_cell_238_96 (.BL(BL96),.BLN(BLN96),.WL(WL238));
sram_cell_6t_5 inst_cell_238_97 (.BL(BL97),.BLN(BLN97),.WL(WL238));
sram_cell_6t_5 inst_cell_238_98 (.BL(BL98),.BLN(BLN98),.WL(WL238));
sram_cell_6t_5 inst_cell_238_99 (.BL(BL99),.BLN(BLN99),.WL(WL238));
sram_cell_6t_5 inst_cell_238_100 (.BL(BL100),.BLN(BLN100),.WL(WL238));
sram_cell_6t_5 inst_cell_238_101 (.BL(BL101),.BLN(BLN101),.WL(WL238));
sram_cell_6t_5 inst_cell_238_102 (.BL(BL102),.BLN(BLN102),.WL(WL238));
sram_cell_6t_5 inst_cell_238_103 (.BL(BL103),.BLN(BLN103),.WL(WL238));
sram_cell_6t_5 inst_cell_238_104 (.BL(BL104),.BLN(BLN104),.WL(WL238));
sram_cell_6t_5 inst_cell_238_105 (.BL(BL105),.BLN(BLN105),.WL(WL238));
sram_cell_6t_5 inst_cell_238_106 (.BL(BL106),.BLN(BLN106),.WL(WL238));
sram_cell_6t_5 inst_cell_238_107 (.BL(BL107),.BLN(BLN107),.WL(WL238));
sram_cell_6t_5 inst_cell_238_108 (.BL(BL108),.BLN(BLN108),.WL(WL238));
sram_cell_6t_5 inst_cell_238_109 (.BL(BL109),.BLN(BLN109),.WL(WL238));
sram_cell_6t_5 inst_cell_238_110 (.BL(BL110),.BLN(BLN110),.WL(WL238));
sram_cell_6t_5 inst_cell_238_111 (.BL(BL111),.BLN(BLN111),.WL(WL238));
sram_cell_6t_5 inst_cell_238_112 (.BL(BL112),.BLN(BLN112),.WL(WL238));
sram_cell_6t_5 inst_cell_238_113 (.BL(BL113),.BLN(BLN113),.WL(WL238));
sram_cell_6t_5 inst_cell_238_114 (.BL(BL114),.BLN(BLN114),.WL(WL238));
sram_cell_6t_5 inst_cell_238_115 (.BL(BL115),.BLN(BLN115),.WL(WL238));
sram_cell_6t_5 inst_cell_238_116 (.BL(BL116),.BLN(BLN116),.WL(WL238));
sram_cell_6t_5 inst_cell_238_117 (.BL(BL117),.BLN(BLN117),.WL(WL238));
sram_cell_6t_5 inst_cell_238_118 (.BL(BL118),.BLN(BLN118),.WL(WL238));
sram_cell_6t_5 inst_cell_238_119 (.BL(BL119),.BLN(BLN119),.WL(WL238));
sram_cell_6t_5 inst_cell_238_120 (.BL(BL120),.BLN(BLN120),.WL(WL238));
sram_cell_6t_5 inst_cell_238_121 (.BL(BL121),.BLN(BLN121),.WL(WL238));
sram_cell_6t_5 inst_cell_238_122 (.BL(BL122),.BLN(BLN122),.WL(WL238));
sram_cell_6t_5 inst_cell_238_123 (.BL(BL123),.BLN(BLN123),.WL(WL238));
sram_cell_6t_5 inst_cell_238_124 (.BL(BL124),.BLN(BLN124),.WL(WL238));
sram_cell_6t_5 inst_cell_238_125 (.BL(BL125),.BLN(BLN125),.WL(WL238));
sram_cell_6t_5 inst_cell_238_126 (.BL(BL126),.BLN(BLN126),.WL(WL238));
sram_cell_6t_5 inst_cell_238_127 (.BL(BL127),.BLN(BLN127),.WL(WL238));
sram_cell_6t_5 inst_cell_239_0 (.BL(BL0),.BLN(BLN0),.WL(WL239));
sram_cell_6t_5 inst_cell_239_1 (.BL(BL1),.BLN(BLN1),.WL(WL239));
sram_cell_6t_5 inst_cell_239_2 (.BL(BL2),.BLN(BLN2),.WL(WL239));
sram_cell_6t_5 inst_cell_239_3 (.BL(BL3),.BLN(BLN3),.WL(WL239));
sram_cell_6t_5 inst_cell_239_4 (.BL(BL4),.BLN(BLN4),.WL(WL239));
sram_cell_6t_5 inst_cell_239_5 (.BL(BL5),.BLN(BLN5),.WL(WL239));
sram_cell_6t_5 inst_cell_239_6 (.BL(BL6),.BLN(BLN6),.WL(WL239));
sram_cell_6t_5 inst_cell_239_7 (.BL(BL7),.BLN(BLN7),.WL(WL239));
sram_cell_6t_5 inst_cell_239_8 (.BL(BL8),.BLN(BLN8),.WL(WL239));
sram_cell_6t_5 inst_cell_239_9 (.BL(BL9),.BLN(BLN9),.WL(WL239));
sram_cell_6t_5 inst_cell_239_10 (.BL(BL10),.BLN(BLN10),.WL(WL239));
sram_cell_6t_5 inst_cell_239_11 (.BL(BL11),.BLN(BLN11),.WL(WL239));
sram_cell_6t_5 inst_cell_239_12 (.BL(BL12),.BLN(BLN12),.WL(WL239));
sram_cell_6t_5 inst_cell_239_13 (.BL(BL13),.BLN(BLN13),.WL(WL239));
sram_cell_6t_5 inst_cell_239_14 (.BL(BL14),.BLN(BLN14),.WL(WL239));
sram_cell_6t_5 inst_cell_239_15 (.BL(BL15),.BLN(BLN15),.WL(WL239));
sram_cell_6t_5 inst_cell_239_16 (.BL(BL16),.BLN(BLN16),.WL(WL239));
sram_cell_6t_5 inst_cell_239_17 (.BL(BL17),.BLN(BLN17),.WL(WL239));
sram_cell_6t_5 inst_cell_239_18 (.BL(BL18),.BLN(BLN18),.WL(WL239));
sram_cell_6t_5 inst_cell_239_19 (.BL(BL19),.BLN(BLN19),.WL(WL239));
sram_cell_6t_5 inst_cell_239_20 (.BL(BL20),.BLN(BLN20),.WL(WL239));
sram_cell_6t_5 inst_cell_239_21 (.BL(BL21),.BLN(BLN21),.WL(WL239));
sram_cell_6t_5 inst_cell_239_22 (.BL(BL22),.BLN(BLN22),.WL(WL239));
sram_cell_6t_5 inst_cell_239_23 (.BL(BL23),.BLN(BLN23),.WL(WL239));
sram_cell_6t_5 inst_cell_239_24 (.BL(BL24),.BLN(BLN24),.WL(WL239));
sram_cell_6t_5 inst_cell_239_25 (.BL(BL25),.BLN(BLN25),.WL(WL239));
sram_cell_6t_5 inst_cell_239_26 (.BL(BL26),.BLN(BLN26),.WL(WL239));
sram_cell_6t_5 inst_cell_239_27 (.BL(BL27),.BLN(BLN27),.WL(WL239));
sram_cell_6t_5 inst_cell_239_28 (.BL(BL28),.BLN(BLN28),.WL(WL239));
sram_cell_6t_5 inst_cell_239_29 (.BL(BL29),.BLN(BLN29),.WL(WL239));
sram_cell_6t_5 inst_cell_239_30 (.BL(BL30),.BLN(BLN30),.WL(WL239));
sram_cell_6t_5 inst_cell_239_31 (.BL(BL31),.BLN(BLN31),.WL(WL239));
sram_cell_6t_5 inst_cell_239_32 (.BL(BL32),.BLN(BLN32),.WL(WL239));
sram_cell_6t_5 inst_cell_239_33 (.BL(BL33),.BLN(BLN33),.WL(WL239));
sram_cell_6t_5 inst_cell_239_34 (.BL(BL34),.BLN(BLN34),.WL(WL239));
sram_cell_6t_5 inst_cell_239_35 (.BL(BL35),.BLN(BLN35),.WL(WL239));
sram_cell_6t_5 inst_cell_239_36 (.BL(BL36),.BLN(BLN36),.WL(WL239));
sram_cell_6t_5 inst_cell_239_37 (.BL(BL37),.BLN(BLN37),.WL(WL239));
sram_cell_6t_5 inst_cell_239_38 (.BL(BL38),.BLN(BLN38),.WL(WL239));
sram_cell_6t_5 inst_cell_239_39 (.BL(BL39),.BLN(BLN39),.WL(WL239));
sram_cell_6t_5 inst_cell_239_40 (.BL(BL40),.BLN(BLN40),.WL(WL239));
sram_cell_6t_5 inst_cell_239_41 (.BL(BL41),.BLN(BLN41),.WL(WL239));
sram_cell_6t_5 inst_cell_239_42 (.BL(BL42),.BLN(BLN42),.WL(WL239));
sram_cell_6t_5 inst_cell_239_43 (.BL(BL43),.BLN(BLN43),.WL(WL239));
sram_cell_6t_5 inst_cell_239_44 (.BL(BL44),.BLN(BLN44),.WL(WL239));
sram_cell_6t_5 inst_cell_239_45 (.BL(BL45),.BLN(BLN45),.WL(WL239));
sram_cell_6t_5 inst_cell_239_46 (.BL(BL46),.BLN(BLN46),.WL(WL239));
sram_cell_6t_5 inst_cell_239_47 (.BL(BL47),.BLN(BLN47),.WL(WL239));
sram_cell_6t_5 inst_cell_239_48 (.BL(BL48),.BLN(BLN48),.WL(WL239));
sram_cell_6t_5 inst_cell_239_49 (.BL(BL49),.BLN(BLN49),.WL(WL239));
sram_cell_6t_5 inst_cell_239_50 (.BL(BL50),.BLN(BLN50),.WL(WL239));
sram_cell_6t_5 inst_cell_239_51 (.BL(BL51),.BLN(BLN51),.WL(WL239));
sram_cell_6t_5 inst_cell_239_52 (.BL(BL52),.BLN(BLN52),.WL(WL239));
sram_cell_6t_5 inst_cell_239_53 (.BL(BL53),.BLN(BLN53),.WL(WL239));
sram_cell_6t_5 inst_cell_239_54 (.BL(BL54),.BLN(BLN54),.WL(WL239));
sram_cell_6t_5 inst_cell_239_55 (.BL(BL55),.BLN(BLN55),.WL(WL239));
sram_cell_6t_5 inst_cell_239_56 (.BL(BL56),.BLN(BLN56),.WL(WL239));
sram_cell_6t_5 inst_cell_239_57 (.BL(BL57),.BLN(BLN57),.WL(WL239));
sram_cell_6t_5 inst_cell_239_58 (.BL(BL58),.BLN(BLN58),.WL(WL239));
sram_cell_6t_5 inst_cell_239_59 (.BL(BL59),.BLN(BLN59),.WL(WL239));
sram_cell_6t_5 inst_cell_239_60 (.BL(BL60),.BLN(BLN60),.WL(WL239));
sram_cell_6t_5 inst_cell_239_61 (.BL(BL61),.BLN(BLN61),.WL(WL239));
sram_cell_6t_5 inst_cell_239_62 (.BL(BL62),.BLN(BLN62),.WL(WL239));
sram_cell_6t_5 inst_cell_239_63 (.BL(BL63),.BLN(BLN63),.WL(WL239));
sram_cell_6t_5 inst_cell_239_64 (.BL(BL64),.BLN(BLN64),.WL(WL239));
sram_cell_6t_5 inst_cell_239_65 (.BL(BL65),.BLN(BLN65),.WL(WL239));
sram_cell_6t_5 inst_cell_239_66 (.BL(BL66),.BLN(BLN66),.WL(WL239));
sram_cell_6t_5 inst_cell_239_67 (.BL(BL67),.BLN(BLN67),.WL(WL239));
sram_cell_6t_5 inst_cell_239_68 (.BL(BL68),.BLN(BLN68),.WL(WL239));
sram_cell_6t_5 inst_cell_239_69 (.BL(BL69),.BLN(BLN69),.WL(WL239));
sram_cell_6t_5 inst_cell_239_70 (.BL(BL70),.BLN(BLN70),.WL(WL239));
sram_cell_6t_5 inst_cell_239_71 (.BL(BL71),.BLN(BLN71),.WL(WL239));
sram_cell_6t_5 inst_cell_239_72 (.BL(BL72),.BLN(BLN72),.WL(WL239));
sram_cell_6t_5 inst_cell_239_73 (.BL(BL73),.BLN(BLN73),.WL(WL239));
sram_cell_6t_5 inst_cell_239_74 (.BL(BL74),.BLN(BLN74),.WL(WL239));
sram_cell_6t_5 inst_cell_239_75 (.BL(BL75),.BLN(BLN75),.WL(WL239));
sram_cell_6t_5 inst_cell_239_76 (.BL(BL76),.BLN(BLN76),.WL(WL239));
sram_cell_6t_5 inst_cell_239_77 (.BL(BL77),.BLN(BLN77),.WL(WL239));
sram_cell_6t_5 inst_cell_239_78 (.BL(BL78),.BLN(BLN78),.WL(WL239));
sram_cell_6t_5 inst_cell_239_79 (.BL(BL79),.BLN(BLN79),.WL(WL239));
sram_cell_6t_5 inst_cell_239_80 (.BL(BL80),.BLN(BLN80),.WL(WL239));
sram_cell_6t_5 inst_cell_239_81 (.BL(BL81),.BLN(BLN81),.WL(WL239));
sram_cell_6t_5 inst_cell_239_82 (.BL(BL82),.BLN(BLN82),.WL(WL239));
sram_cell_6t_5 inst_cell_239_83 (.BL(BL83),.BLN(BLN83),.WL(WL239));
sram_cell_6t_5 inst_cell_239_84 (.BL(BL84),.BLN(BLN84),.WL(WL239));
sram_cell_6t_5 inst_cell_239_85 (.BL(BL85),.BLN(BLN85),.WL(WL239));
sram_cell_6t_5 inst_cell_239_86 (.BL(BL86),.BLN(BLN86),.WL(WL239));
sram_cell_6t_5 inst_cell_239_87 (.BL(BL87),.BLN(BLN87),.WL(WL239));
sram_cell_6t_5 inst_cell_239_88 (.BL(BL88),.BLN(BLN88),.WL(WL239));
sram_cell_6t_5 inst_cell_239_89 (.BL(BL89),.BLN(BLN89),.WL(WL239));
sram_cell_6t_5 inst_cell_239_90 (.BL(BL90),.BLN(BLN90),.WL(WL239));
sram_cell_6t_5 inst_cell_239_91 (.BL(BL91),.BLN(BLN91),.WL(WL239));
sram_cell_6t_5 inst_cell_239_92 (.BL(BL92),.BLN(BLN92),.WL(WL239));
sram_cell_6t_5 inst_cell_239_93 (.BL(BL93),.BLN(BLN93),.WL(WL239));
sram_cell_6t_5 inst_cell_239_94 (.BL(BL94),.BLN(BLN94),.WL(WL239));
sram_cell_6t_5 inst_cell_239_95 (.BL(BL95),.BLN(BLN95),.WL(WL239));
sram_cell_6t_5 inst_cell_239_96 (.BL(BL96),.BLN(BLN96),.WL(WL239));
sram_cell_6t_5 inst_cell_239_97 (.BL(BL97),.BLN(BLN97),.WL(WL239));
sram_cell_6t_5 inst_cell_239_98 (.BL(BL98),.BLN(BLN98),.WL(WL239));
sram_cell_6t_5 inst_cell_239_99 (.BL(BL99),.BLN(BLN99),.WL(WL239));
sram_cell_6t_5 inst_cell_239_100 (.BL(BL100),.BLN(BLN100),.WL(WL239));
sram_cell_6t_5 inst_cell_239_101 (.BL(BL101),.BLN(BLN101),.WL(WL239));
sram_cell_6t_5 inst_cell_239_102 (.BL(BL102),.BLN(BLN102),.WL(WL239));
sram_cell_6t_5 inst_cell_239_103 (.BL(BL103),.BLN(BLN103),.WL(WL239));
sram_cell_6t_5 inst_cell_239_104 (.BL(BL104),.BLN(BLN104),.WL(WL239));
sram_cell_6t_5 inst_cell_239_105 (.BL(BL105),.BLN(BLN105),.WL(WL239));
sram_cell_6t_5 inst_cell_239_106 (.BL(BL106),.BLN(BLN106),.WL(WL239));
sram_cell_6t_5 inst_cell_239_107 (.BL(BL107),.BLN(BLN107),.WL(WL239));
sram_cell_6t_5 inst_cell_239_108 (.BL(BL108),.BLN(BLN108),.WL(WL239));
sram_cell_6t_5 inst_cell_239_109 (.BL(BL109),.BLN(BLN109),.WL(WL239));
sram_cell_6t_5 inst_cell_239_110 (.BL(BL110),.BLN(BLN110),.WL(WL239));
sram_cell_6t_5 inst_cell_239_111 (.BL(BL111),.BLN(BLN111),.WL(WL239));
sram_cell_6t_5 inst_cell_239_112 (.BL(BL112),.BLN(BLN112),.WL(WL239));
sram_cell_6t_5 inst_cell_239_113 (.BL(BL113),.BLN(BLN113),.WL(WL239));
sram_cell_6t_5 inst_cell_239_114 (.BL(BL114),.BLN(BLN114),.WL(WL239));
sram_cell_6t_5 inst_cell_239_115 (.BL(BL115),.BLN(BLN115),.WL(WL239));
sram_cell_6t_5 inst_cell_239_116 (.BL(BL116),.BLN(BLN116),.WL(WL239));
sram_cell_6t_5 inst_cell_239_117 (.BL(BL117),.BLN(BLN117),.WL(WL239));
sram_cell_6t_5 inst_cell_239_118 (.BL(BL118),.BLN(BLN118),.WL(WL239));
sram_cell_6t_5 inst_cell_239_119 (.BL(BL119),.BLN(BLN119),.WL(WL239));
sram_cell_6t_5 inst_cell_239_120 (.BL(BL120),.BLN(BLN120),.WL(WL239));
sram_cell_6t_5 inst_cell_239_121 (.BL(BL121),.BLN(BLN121),.WL(WL239));
sram_cell_6t_5 inst_cell_239_122 (.BL(BL122),.BLN(BLN122),.WL(WL239));
sram_cell_6t_5 inst_cell_239_123 (.BL(BL123),.BLN(BLN123),.WL(WL239));
sram_cell_6t_5 inst_cell_239_124 (.BL(BL124),.BLN(BLN124),.WL(WL239));
sram_cell_6t_5 inst_cell_239_125 (.BL(BL125),.BLN(BLN125),.WL(WL239));
sram_cell_6t_5 inst_cell_239_126 (.BL(BL126),.BLN(BLN126),.WL(WL239));
sram_cell_6t_5 inst_cell_239_127 (.BL(BL127),.BLN(BLN127),.WL(WL239));
sram_cell_6t_5 inst_cell_240_0 (.BL(BL0),.BLN(BLN0),.WL(WL240));
sram_cell_6t_5 inst_cell_240_1 (.BL(BL1),.BLN(BLN1),.WL(WL240));
sram_cell_6t_5 inst_cell_240_2 (.BL(BL2),.BLN(BLN2),.WL(WL240));
sram_cell_6t_5 inst_cell_240_3 (.BL(BL3),.BLN(BLN3),.WL(WL240));
sram_cell_6t_5 inst_cell_240_4 (.BL(BL4),.BLN(BLN4),.WL(WL240));
sram_cell_6t_5 inst_cell_240_5 (.BL(BL5),.BLN(BLN5),.WL(WL240));
sram_cell_6t_5 inst_cell_240_6 (.BL(BL6),.BLN(BLN6),.WL(WL240));
sram_cell_6t_5 inst_cell_240_7 (.BL(BL7),.BLN(BLN7),.WL(WL240));
sram_cell_6t_5 inst_cell_240_8 (.BL(BL8),.BLN(BLN8),.WL(WL240));
sram_cell_6t_5 inst_cell_240_9 (.BL(BL9),.BLN(BLN9),.WL(WL240));
sram_cell_6t_5 inst_cell_240_10 (.BL(BL10),.BLN(BLN10),.WL(WL240));
sram_cell_6t_5 inst_cell_240_11 (.BL(BL11),.BLN(BLN11),.WL(WL240));
sram_cell_6t_5 inst_cell_240_12 (.BL(BL12),.BLN(BLN12),.WL(WL240));
sram_cell_6t_5 inst_cell_240_13 (.BL(BL13),.BLN(BLN13),.WL(WL240));
sram_cell_6t_5 inst_cell_240_14 (.BL(BL14),.BLN(BLN14),.WL(WL240));
sram_cell_6t_5 inst_cell_240_15 (.BL(BL15),.BLN(BLN15),.WL(WL240));
sram_cell_6t_5 inst_cell_240_16 (.BL(BL16),.BLN(BLN16),.WL(WL240));
sram_cell_6t_5 inst_cell_240_17 (.BL(BL17),.BLN(BLN17),.WL(WL240));
sram_cell_6t_5 inst_cell_240_18 (.BL(BL18),.BLN(BLN18),.WL(WL240));
sram_cell_6t_5 inst_cell_240_19 (.BL(BL19),.BLN(BLN19),.WL(WL240));
sram_cell_6t_5 inst_cell_240_20 (.BL(BL20),.BLN(BLN20),.WL(WL240));
sram_cell_6t_5 inst_cell_240_21 (.BL(BL21),.BLN(BLN21),.WL(WL240));
sram_cell_6t_5 inst_cell_240_22 (.BL(BL22),.BLN(BLN22),.WL(WL240));
sram_cell_6t_5 inst_cell_240_23 (.BL(BL23),.BLN(BLN23),.WL(WL240));
sram_cell_6t_5 inst_cell_240_24 (.BL(BL24),.BLN(BLN24),.WL(WL240));
sram_cell_6t_5 inst_cell_240_25 (.BL(BL25),.BLN(BLN25),.WL(WL240));
sram_cell_6t_5 inst_cell_240_26 (.BL(BL26),.BLN(BLN26),.WL(WL240));
sram_cell_6t_5 inst_cell_240_27 (.BL(BL27),.BLN(BLN27),.WL(WL240));
sram_cell_6t_5 inst_cell_240_28 (.BL(BL28),.BLN(BLN28),.WL(WL240));
sram_cell_6t_5 inst_cell_240_29 (.BL(BL29),.BLN(BLN29),.WL(WL240));
sram_cell_6t_5 inst_cell_240_30 (.BL(BL30),.BLN(BLN30),.WL(WL240));
sram_cell_6t_5 inst_cell_240_31 (.BL(BL31),.BLN(BLN31),.WL(WL240));
sram_cell_6t_5 inst_cell_240_32 (.BL(BL32),.BLN(BLN32),.WL(WL240));
sram_cell_6t_5 inst_cell_240_33 (.BL(BL33),.BLN(BLN33),.WL(WL240));
sram_cell_6t_5 inst_cell_240_34 (.BL(BL34),.BLN(BLN34),.WL(WL240));
sram_cell_6t_5 inst_cell_240_35 (.BL(BL35),.BLN(BLN35),.WL(WL240));
sram_cell_6t_5 inst_cell_240_36 (.BL(BL36),.BLN(BLN36),.WL(WL240));
sram_cell_6t_5 inst_cell_240_37 (.BL(BL37),.BLN(BLN37),.WL(WL240));
sram_cell_6t_5 inst_cell_240_38 (.BL(BL38),.BLN(BLN38),.WL(WL240));
sram_cell_6t_5 inst_cell_240_39 (.BL(BL39),.BLN(BLN39),.WL(WL240));
sram_cell_6t_5 inst_cell_240_40 (.BL(BL40),.BLN(BLN40),.WL(WL240));
sram_cell_6t_5 inst_cell_240_41 (.BL(BL41),.BLN(BLN41),.WL(WL240));
sram_cell_6t_5 inst_cell_240_42 (.BL(BL42),.BLN(BLN42),.WL(WL240));
sram_cell_6t_5 inst_cell_240_43 (.BL(BL43),.BLN(BLN43),.WL(WL240));
sram_cell_6t_5 inst_cell_240_44 (.BL(BL44),.BLN(BLN44),.WL(WL240));
sram_cell_6t_5 inst_cell_240_45 (.BL(BL45),.BLN(BLN45),.WL(WL240));
sram_cell_6t_5 inst_cell_240_46 (.BL(BL46),.BLN(BLN46),.WL(WL240));
sram_cell_6t_5 inst_cell_240_47 (.BL(BL47),.BLN(BLN47),.WL(WL240));
sram_cell_6t_5 inst_cell_240_48 (.BL(BL48),.BLN(BLN48),.WL(WL240));
sram_cell_6t_5 inst_cell_240_49 (.BL(BL49),.BLN(BLN49),.WL(WL240));
sram_cell_6t_5 inst_cell_240_50 (.BL(BL50),.BLN(BLN50),.WL(WL240));
sram_cell_6t_5 inst_cell_240_51 (.BL(BL51),.BLN(BLN51),.WL(WL240));
sram_cell_6t_5 inst_cell_240_52 (.BL(BL52),.BLN(BLN52),.WL(WL240));
sram_cell_6t_5 inst_cell_240_53 (.BL(BL53),.BLN(BLN53),.WL(WL240));
sram_cell_6t_5 inst_cell_240_54 (.BL(BL54),.BLN(BLN54),.WL(WL240));
sram_cell_6t_5 inst_cell_240_55 (.BL(BL55),.BLN(BLN55),.WL(WL240));
sram_cell_6t_5 inst_cell_240_56 (.BL(BL56),.BLN(BLN56),.WL(WL240));
sram_cell_6t_5 inst_cell_240_57 (.BL(BL57),.BLN(BLN57),.WL(WL240));
sram_cell_6t_5 inst_cell_240_58 (.BL(BL58),.BLN(BLN58),.WL(WL240));
sram_cell_6t_5 inst_cell_240_59 (.BL(BL59),.BLN(BLN59),.WL(WL240));
sram_cell_6t_5 inst_cell_240_60 (.BL(BL60),.BLN(BLN60),.WL(WL240));
sram_cell_6t_5 inst_cell_240_61 (.BL(BL61),.BLN(BLN61),.WL(WL240));
sram_cell_6t_5 inst_cell_240_62 (.BL(BL62),.BLN(BLN62),.WL(WL240));
sram_cell_6t_5 inst_cell_240_63 (.BL(BL63),.BLN(BLN63),.WL(WL240));
sram_cell_6t_5 inst_cell_240_64 (.BL(BL64),.BLN(BLN64),.WL(WL240));
sram_cell_6t_5 inst_cell_240_65 (.BL(BL65),.BLN(BLN65),.WL(WL240));
sram_cell_6t_5 inst_cell_240_66 (.BL(BL66),.BLN(BLN66),.WL(WL240));
sram_cell_6t_5 inst_cell_240_67 (.BL(BL67),.BLN(BLN67),.WL(WL240));
sram_cell_6t_5 inst_cell_240_68 (.BL(BL68),.BLN(BLN68),.WL(WL240));
sram_cell_6t_5 inst_cell_240_69 (.BL(BL69),.BLN(BLN69),.WL(WL240));
sram_cell_6t_5 inst_cell_240_70 (.BL(BL70),.BLN(BLN70),.WL(WL240));
sram_cell_6t_5 inst_cell_240_71 (.BL(BL71),.BLN(BLN71),.WL(WL240));
sram_cell_6t_5 inst_cell_240_72 (.BL(BL72),.BLN(BLN72),.WL(WL240));
sram_cell_6t_5 inst_cell_240_73 (.BL(BL73),.BLN(BLN73),.WL(WL240));
sram_cell_6t_5 inst_cell_240_74 (.BL(BL74),.BLN(BLN74),.WL(WL240));
sram_cell_6t_5 inst_cell_240_75 (.BL(BL75),.BLN(BLN75),.WL(WL240));
sram_cell_6t_5 inst_cell_240_76 (.BL(BL76),.BLN(BLN76),.WL(WL240));
sram_cell_6t_5 inst_cell_240_77 (.BL(BL77),.BLN(BLN77),.WL(WL240));
sram_cell_6t_5 inst_cell_240_78 (.BL(BL78),.BLN(BLN78),.WL(WL240));
sram_cell_6t_5 inst_cell_240_79 (.BL(BL79),.BLN(BLN79),.WL(WL240));
sram_cell_6t_5 inst_cell_240_80 (.BL(BL80),.BLN(BLN80),.WL(WL240));
sram_cell_6t_5 inst_cell_240_81 (.BL(BL81),.BLN(BLN81),.WL(WL240));
sram_cell_6t_5 inst_cell_240_82 (.BL(BL82),.BLN(BLN82),.WL(WL240));
sram_cell_6t_5 inst_cell_240_83 (.BL(BL83),.BLN(BLN83),.WL(WL240));
sram_cell_6t_5 inst_cell_240_84 (.BL(BL84),.BLN(BLN84),.WL(WL240));
sram_cell_6t_5 inst_cell_240_85 (.BL(BL85),.BLN(BLN85),.WL(WL240));
sram_cell_6t_5 inst_cell_240_86 (.BL(BL86),.BLN(BLN86),.WL(WL240));
sram_cell_6t_5 inst_cell_240_87 (.BL(BL87),.BLN(BLN87),.WL(WL240));
sram_cell_6t_5 inst_cell_240_88 (.BL(BL88),.BLN(BLN88),.WL(WL240));
sram_cell_6t_5 inst_cell_240_89 (.BL(BL89),.BLN(BLN89),.WL(WL240));
sram_cell_6t_5 inst_cell_240_90 (.BL(BL90),.BLN(BLN90),.WL(WL240));
sram_cell_6t_5 inst_cell_240_91 (.BL(BL91),.BLN(BLN91),.WL(WL240));
sram_cell_6t_5 inst_cell_240_92 (.BL(BL92),.BLN(BLN92),.WL(WL240));
sram_cell_6t_5 inst_cell_240_93 (.BL(BL93),.BLN(BLN93),.WL(WL240));
sram_cell_6t_5 inst_cell_240_94 (.BL(BL94),.BLN(BLN94),.WL(WL240));
sram_cell_6t_5 inst_cell_240_95 (.BL(BL95),.BLN(BLN95),.WL(WL240));
sram_cell_6t_5 inst_cell_240_96 (.BL(BL96),.BLN(BLN96),.WL(WL240));
sram_cell_6t_5 inst_cell_240_97 (.BL(BL97),.BLN(BLN97),.WL(WL240));
sram_cell_6t_5 inst_cell_240_98 (.BL(BL98),.BLN(BLN98),.WL(WL240));
sram_cell_6t_5 inst_cell_240_99 (.BL(BL99),.BLN(BLN99),.WL(WL240));
sram_cell_6t_5 inst_cell_240_100 (.BL(BL100),.BLN(BLN100),.WL(WL240));
sram_cell_6t_5 inst_cell_240_101 (.BL(BL101),.BLN(BLN101),.WL(WL240));
sram_cell_6t_5 inst_cell_240_102 (.BL(BL102),.BLN(BLN102),.WL(WL240));
sram_cell_6t_5 inst_cell_240_103 (.BL(BL103),.BLN(BLN103),.WL(WL240));
sram_cell_6t_5 inst_cell_240_104 (.BL(BL104),.BLN(BLN104),.WL(WL240));
sram_cell_6t_5 inst_cell_240_105 (.BL(BL105),.BLN(BLN105),.WL(WL240));
sram_cell_6t_5 inst_cell_240_106 (.BL(BL106),.BLN(BLN106),.WL(WL240));
sram_cell_6t_5 inst_cell_240_107 (.BL(BL107),.BLN(BLN107),.WL(WL240));
sram_cell_6t_5 inst_cell_240_108 (.BL(BL108),.BLN(BLN108),.WL(WL240));
sram_cell_6t_5 inst_cell_240_109 (.BL(BL109),.BLN(BLN109),.WL(WL240));
sram_cell_6t_5 inst_cell_240_110 (.BL(BL110),.BLN(BLN110),.WL(WL240));
sram_cell_6t_5 inst_cell_240_111 (.BL(BL111),.BLN(BLN111),.WL(WL240));
sram_cell_6t_5 inst_cell_240_112 (.BL(BL112),.BLN(BLN112),.WL(WL240));
sram_cell_6t_5 inst_cell_240_113 (.BL(BL113),.BLN(BLN113),.WL(WL240));
sram_cell_6t_5 inst_cell_240_114 (.BL(BL114),.BLN(BLN114),.WL(WL240));
sram_cell_6t_5 inst_cell_240_115 (.BL(BL115),.BLN(BLN115),.WL(WL240));
sram_cell_6t_5 inst_cell_240_116 (.BL(BL116),.BLN(BLN116),.WL(WL240));
sram_cell_6t_5 inst_cell_240_117 (.BL(BL117),.BLN(BLN117),.WL(WL240));
sram_cell_6t_5 inst_cell_240_118 (.BL(BL118),.BLN(BLN118),.WL(WL240));
sram_cell_6t_5 inst_cell_240_119 (.BL(BL119),.BLN(BLN119),.WL(WL240));
sram_cell_6t_5 inst_cell_240_120 (.BL(BL120),.BLN(BLN120),.WL(WL240));
sram_cell_6t_5 inst_cell_240_121 (.BL(BL121),.BLN(BLN121),.WL(WL240));
sram_cell_6t_5 inst_cell_240_122 (.BL(BL122),.BLN(BLN122),.WL(WL240));
sram_cell_6t_5 inst_cell_240_123 (.BL(BL123),.BLN(BLN123),.WL(WL240));
sram_cell_6t_5 inst_cell_240_124 (.BL(BL124),.BLN(BLN124),.WL(WL240));
sram_cell_6t_5 inst_cell_240_125 (.BL(BL125),.BLN(BLN125),.WL(WL240));
sram_cell_6t_5 inst_cell_240_126 (.BL(BL126),.BLN(BLN126),.WL(WL240));
sram_cell_6t_5 inst_cell_240_127 (.BL(BL127),.BLN(BLN127),.WL(WL240));
sram_cell_6t_5 inst_cell_241_0 (.BL(BL0),.BLN(BLN0),.WL(WL241));
sram_cell_6t_5 inst_cell_241_1 (.BL(BL1),.BLN(BLN1),.WL(WL241));
sram_cell_6t_5 inst_cell_241_2 (.BL(BL2),.BLN(BLN2),.WL(WL241));
sram_cell_6t_5 inst_cell_241_3 (.BL(BL3),.BLN(BLN3),.WL(WL241));
sram_cell_6t_5 inst_cell_241_4 (.BL(BL4),.BLN(BLN4),.WL(WL241));
sram_cell_6t_5 inst_cell_241_5 (.BL(BL5),.BLN(BLN5),.WL(WL241));
sram_cell_6t_5 inst_cell_241_6 (.BL(BL6),.BLN(BLN6),.WL(WL241));
sram_cell_6t_5 inst_cell_241_7 (.BL(BL7),.BLN(BLN7),.WL(WL241));
sram_cell_6t_5 inst_cell_241_8 (.BL(BL8),.BLN(BLN8),.WL(WL241));
sram_cell_6t_5 inst_cell_241_9 (.BL(BL9),.BLN(BLN9),.WL(WL241));
sram_cell_6t_5 inst_cell_241_10 (.BL(BL10),.BLN(BLN10),.WL(WL241));
sram_cell_6t_5 inst_cell_241_11 (.BL(BL11),.BLN(BLN11),.WL(WL241));
sram_cell_6t_5 inst_cell_241_12 (.BL(BL12),.BLN(BLN12),.WL(WL241));
sram_cell_6t_5 inst_cell_241_13 (.BL(BL13),.BLN(BLN13),.WL(WL241));
sram_cell_6t_5 inst_cell_241_14 (.BL(BL14),.BLN(BLN14),.WL(WL241));
sram_cell_6t_5 inst_cell_241_15 (.BL(BL15),.BLN(BLN15),.WL(WL241));
sram_cell_6t_5 inst_cell_241_16 (.BL(BL16),.BLN(BLN16),.WL(WL241));
sram_cell_6t_5 inst_cell_241_17 (.BL(BL17),.BLN(BLN17),.WL(WL241));
sram_cell_6t_5 inst_cell_241_18 (.BL(BL18),.BLN(BLN18),.WL(WL241));
sram_cell_6t_5 inst_cell_241_19 (.BL(BL19),.BLN(BLN19),.WL(WL241));
sram_cell_6t_5 inst_cell_241_20 (.BL(BL20),.BLN(BLN20),.WL(WL241));
sram_cell_6t_5 inst_cell_241_21 (.BL(BL21),.BLN(BLN21),.WL(WL241));
sram_cell_6t_5 inst_cell_241_22 (.BL(BL22),.BLN(BLN22),.WL(WL241));
sram_cell_6t_5 inst_cell_241_23 (.BL(BL23),.BLN(BLN23),.WL(WL241));
sram_cell_6t_5 inst_cell_241_24 (.BL(BL24),.BLN(BLN24),.WL(WL241));
sram_cell_6t_5 inst_cell_241_25 (.BL(BL25),.BLN(BLN25),.WL(WL241));
sram_cell_6t_5 inst_cell_241_26 (.BL(BL26),.BLN(BLN26),.WL(WL241));
sram_cell_6t_5 inst_cell_241_27 (.BL(BL27),.BLN(BLN27),.WL(WL241));
sram_cell_6t_5 inst_cell_241_28 (.BL(BL28),.BLN(BLN28),.WL(WL241));
sram_cell_6t_5 inst_cell_241_29 (.BL(BL29),.BLN(BLN29),.WL(WL241));
sram_cell_6t_5 inst_cell_241_30 (.BL(BL30),.BLN(BLN30),.WL(WL241));
sram_cell_6t_5 inst_cell_241_31 (.BL(BL31),.BLN(BLN31),.WL(WL241));
sram_cell_6t_5 inst_cell_241_32 (.BL(BL32),.BLN(BLN32),.WL(WL241));
sram_cell_6t_5 inst_cell_241_33 (.BL(BL33),.BLN(BLN33),.WL(WL241));
sram_cell_6t_5 inst_cell_241_34 (.BL(BL34),.BLN(BLN34),.WL(WL241));
sram_cell_6t_5 inst_cell_241_35 (.BL(BL35),.BLN(BLN35),.WL(WL241));
sram_cell_6t_5 inst_cell_241_36 (.BL(BL36),.BLN(BLN36),.WL(WL241));
sram_cell_6t_5 inst_cell_241_37 (.BL(BL37),.BLN(BLN37),.WL(WL241));
sram_cell_6t_5 inst_cell_241_38 (.BL(BL38),.BLN(BLN38),.WL(WL241));
sram_cell_6t_5 inst_cell_241_39 (.BL(BL39),.BLN(BLN39),.WL(WL241));
sram_cell_6t_5 inst_cell_241_40 (.BL(BL40),.BLN(BLN40),.WL(WL241));
sram_cell_6t_5 inst_cell_241_41 (.BL(BL41),.BLN(BLN41),.WL(WL241));
sram_cell_6t_5 inst_cell_241_42 (.BL(BL42),.BLN(BLN42),.WL(WL241));
sram_cell_6t_5 inst_cell_241_43 (.BL(BL43),.BLN(BLN43),.WL(WL241));
sram_cell_6t_5 inst_cell_241_44 (.BL(BL44),.BLN(BLN44),.WL(WL241));
sram_cell_6t_5 inst_cell_241_45 (.BL(BL45),.BLN(BLN45),.WL(WL241));
sram_cell_6t_5 inst_cell_241_46 (.BL(BL46),.BLN(BLN46),.WL(WL241));
sram_cell_6t_5 inst_cell_241_47 (.BL(BL47),.BLN(BLN47),.WL(WL241));
sram_cell_6t_5 inst_cell_241_48 (.BL(BL48),.BLN(BLN48),.WL(WL241));
sram_cell_6t_5 inst_cell_241_49 (.BL(BL49),.BLN(BLN49),.WL(WL241));
sram_cell_6t_5 inst_cell_241_50 (.BL(BL50),.BLN(BLN50),.WL(WL241));
sram_cell_6t_5 inst_cell_241_51 (.BL(BL51),.BLN(BLN51),.WL(WL241));
sram_cell_6t_5 inst_cell_241_52 (.BL(BL52),.BLN(BLN52),.WL(WL241));
sram_cell_6t_5 inst_cell_241_53 (.BL(BL53),.BLN(BLN53),.WL(WL241));
sram_cell_6t_5 inst_cell_241_54 (.BL(BL54),.BLN(BLN54),.WL(WL241));
sram_cell_6t_5 inst_cell_241_55 (.BL(BL55),.BLN(BLN55),.WL(WL241));
sram_cell_6t_5 inst_cell_241_56 (.BL(BL56),.BLN(BLN56),.WL(WL241));
sram_cell_6t_5 inst_cell_241_57 (.BL(BL57),.BLN(BLN57),.WL(WL241));
sram_cell_6t_5 inst_cell_241_58 (.BL(BL58),.BLN(BLN58),.WL(WL241));
sram_cell_6t_5 inst_cell_241_59 (.BL(BL59),.BLN(BLN59),.WL(WL241));
sram_cell_6t_5 inst_cell_241_60 (.BL(BL60),.BLN(BLN60),.WL(WL241));
sram_cell_6t_5 inst_cell_241_61 (.BL(BL61),.BLN(BLN61),.WL(WL241));
sram_cell_6t_5 inst_cell_241_62 (.BL(BL62),.BLN(BLN62),.WL(WL241));
sram_cell_6t_5 inst_cell_241_63 (.BL(BL63),.BLN(BLN63),.WL(WL241));
sram_cell_6t_5 inst_cell_241_64 (.BL(BL64),.BLN(BLN64),.WL(WL241));
sram_cell_6t_5 inst_cell_241_65 (.BL(BL65),.BLN(BLN65),.WL(WL241));
sram_cell_6t_5 inst_cell_241_66 (.BL(BL66),.BLN(BLN66),.WL(WL241));
sram_cell_6t_5 inst_cell_241_67 (.BL(BL67),.BLN(BLN67),.WL(WL241));
sram_cell_6t_5 inst_cell_241_68 (.BL(BL68),.BLN(BLN68),.WL(WL241));
sram_cell_6t_5 inst_cell_241_69 (.BL(BL69),.BLN(BLN69),.WL(WL241));
sram_cell_6t_5 inst_cell_241_70 (.BL(BL70),.BLN(BLN70),.WL(WL241));
sram_cell_6t_5 inst_cell_241_71 (.BL(BL71),.BLN(BLN71),.WL(WL241));
sram_cell_6t_5 inst_cell_241_72 (.BL(BL72),.BLN(BLN72),.WL(WL241));
sram_cell_6t_5 inst_cell_241_73 (.BL(BL73),.BLN(BLN73),.WL(WL241));
sram_cell_6t_5 inst_cell_241_74 (.BL(BL74),.BLN(BLN74),.WL(WL241));
sram_cell_6t_5 inst_cell_241_75 (.BL(BL75),.BLN(BLN75),.WL(WL241));
sram_cell_6t_5 inst_cell_241_76 (.BL(BL76),.BLN(BLN76),.WL(WL241));
sram_cell_6t_5 inst_cell_241_77 (.BL(BL77),.BLN(BLN77),.WL(WL241));
sram_cell_6t_5 inst_cell_241_78 (.BL(BL78),.BLN(BLN78),.WL(WL241));
sram_cell_6t_5 inst_cell_241_79 (.BL(BL79),.BLN(BLN79),.WL(WL241));
sram_cell_6t_5 inst_cell_241_80 (.BL(BL80),.BLN(BLN80),.WL(WL241));
sram_cell_6t_5 inst_cell_241_81 (.BL(BL81),.BLN(BLN81),.WL(WL241));
sram_cell_6t_5 inst_cell_241_82 (.BL(BL82),.BLN(BLN82),.WL(WL241));
sram_cell_6t_5 inst_cell_241_83 (.BL(BL83),.BLN(BLN83),.WL(WL241));
sram_cell_6t_5 inst_cell_241_84 (.BL(BL84),.BLN(BLN84),.WL(WL241));
sram_cell_6t_5 inst_cell_241_85 (.BL(BL85),.BLN(BLN85),.WL(WL241));
sram_cell_6t_5 inst_cell_241_86 (.BL(BL86),.BLN(BLN86),.WL(WL241));
sram_cell_6t_5 inst_cell_241_87 (.BL(BL87),.BLN(BLN87),.WL(WL241));
sram_cell_6t_5 inst_cell_241_88 (.BL(BL88),.BLN(BLN88),.WL(WL241));
sram_cell_6t_5 inst_cell_241_89 (.BL(BL89),.BLN(BLN89),.WL(WL241));
sram_cell_6t_5 inst_cell_241_90 (.BL(BL90),.BLN(BLN90),.WL(WL241));
sram_cell_6t_5 inst_cell_241_91 (.BL(BL91),.BLN(BLN91),.WL(WL241));
sram_cell_6t_5 inst_cell_241_92 (.BL(BL92),.BLN(BLN92),.WL(WL241));
sram_cell_6t_5 inst_cell_241_93 (.BL(BL93),.BLN(BLN93),.WL(WL241));
sram_cell_6t_5 inst_cell_241_94 (.BL(BL94),.BLN(BLN94),.WL(WL241));
sram_cell_6t_5 inst_cell_241_95 (.BL(BL95),.BLN(BLN95),.WL(WL241));
sram_cell_6t_5 inst_cell_241_96 (.BL(BL96),.BLN(BLN96),.WL(WL241));
sram_cell_6t_5 inst_cell_241_97 (.BL(BL97),.BLN(BLN97),.WL(WL241));
sram_cell_6t_5 inst_cell_241_98 (.BL(BL98),.BLN(BLN98),.WL(WL241));
sram_cell_6t_5 inst_cell_241_99 (.BL(BL99),.BLN(BLN99),.WL(WL241));
sram_cell_6t_5 inst_cell_241_100 (.BL(BL100),.BLN(BLN100),.WL(WL241));
sram_cell_6t_5 inst_cell_241_101 (.BL(BL101),.BLN(BLN101),.WL(WL241));
sram_cell_6t_5 inst_cell_241_102 (.BL(BL102),.BLN(BLN102),.WL(WL241));
sram_cell_6t_5 inst_cell_241_103 (.BL(BL103),.BLN(BLN103),.WL(WL241));
sram_cell_6t_5 inst_cell_241_104 (.BL(BL104),.BLN(BLN104),.WL(WL241));
sram_cell_6t_5 inst_cell_241_105 (.BL(BL105),.BLN(BLN105),.WL(WL241));
sram_cell_6t_5 inst_cell_241_106 (.BL(BL106),.BLN(BLN106),.WL(WL241));
sram_cell_6t_5 inst_cell_241_107 (.BL(BL107),.BLN(BLN107),.WL(WL241));
sram_cell_6t_5 inst_cell_241_108 (.BL(BL108),.BLN(BLN108),.WL(WL241));
sram_cell_6t_5 inst_cell_241_109 (.BL(BL109),.BLN(BLN109),.WL(WL241));
sram_cell_6t_5 inst_cell_241_110 (.BL(BL110),.BLN(BLN110),.WL(WL241));
sram_cell_6t_5 inst_cell_241_111 (.BL(BL111),.BLN(BLN111),.WL(WL241));
sram_cell_6t_5 inst_cell_241_112 (.BL(BL112),.BLN(BLN112),.WL(WL241));
sram_cell_6t_5 inst_cell_241_113 (.BL(BL113),.BLN(BLN113),.WL(WL241));
sram_cell_6t_5 inst_cell_241_114 (.BL(BL114),.BLN(BLN114),.WL(WL241));
sram_cell_6t_5 inst_cell_241_115 (.BL(BL115),.BLN(BLN115),.WL(WL241));
sram_cell_6t_5 inst_cell_241_116 (.BL(BL116),.BLN(BLN116),.WL(WL241));
sram_cell_6t_5 inst_cell_241_117 (.BL(BL117),.BLN(BLN117),.WL(WL241));
sram_cell_6t_5 inst_cell_241_118 (.BL(BL118),.BLN(BLN118),.WL(WL241));
sram_cell_6t_5 inst_cell_241_119 (.BL(BL119),.BLN(BLN119),.WL(WL241));
sram_cell_6t_5 inst_cell_241_120 (.BL(BL120),.BLN(BLN120),.WL(WL241));
sram_cell_6t_5 inst_cell_241_121 (.BL(BL121),.BLN(BLN121),.WL(WL241));
sram_cell_6t_5 inst_cell_241_122 (.BL(BL122),.BLN(BLN122),.WL(WL241));
sram_cell_6t_5 inst_cell_241_123 (.BL(BL123),.BLN(BLN123),.WL(WL241));
sram_cell_6t_5 inst_cell_241_124 (.BL(BL124),.BLN(BLN124),.WL(WL241));
sram_cell_6t_5 inst_cell_241_125 (.BL(BL125),.BLN(BLN125),.WL(WL241));
sram_cell_6t_5 inst_cell_241_126 (.BL(BL126),.BLN(BLN126),.WL(WL241));
sram_cell_6t_5 inst_cell_241_127 (.BL(BL127),.BLN(BLN127),.WL(WL241));
sram_cell_6t_5 inst_cell_242_0 (.BL(BL0),.BLN(BLN0),.WL(WL242));
sram_cell_6t_5 inst_cell_242_1 (.BL(BL1),.BLN(BLN1),.WL(WL242));
sram_cell_6t_5 inst_cell_242_2 (.BL(BL2),.BLN(BLN2),.WL(WL242));
sram_cell_6t_5 inst_cell_242_3 (.BL(BL3),.BLN(BLN3),.WL(WL242));
sram_cell_6t_5 inst_cell_242_4 (.BL(BL4),.BLN(BLN4),.WL(WL242));
sram_cell_6t_5 inst_cell_242_5 (.BL(BL5),.BLN(BLN5),.WL(WL242));
sram_cell_6t_5 inst_cell_242_6 (.BL(BL6),.BLN(BLN6),.WL(WL242));
sram_cell_6t_5 inst_cell_242_7 (.BL(BL7),.BLN(BLN7),.WL(WL242));
sram_cell_6t_5 inst_cell_242_8 (.BL(BL8),.BLN(BLN8),.WL(WL242));
sram_cell_6t_5 inst_cell_242_9 (.BL(BL9),.BLN(BLN9),.WL(WL242));
sram_cell_6t_5 inst_cell_242_10 (.BL(BL10),.BLN(BLN10),.WL(WL242));
sram_cell_6t_5 inst_cell_242_11 (.BL(BL11),.BLN(BLN11),.WL(WL242));
sram_cell_6t_5 inst_cell_242_12 (.BL(BL12),.BLN(BLN12),.WL(WL242));
sram_cell_6t_5 inst_cell_242_13 (.BL(BL13),.BLN(BLN13),.WL(WL242));
sram_cell_6t_5 inst_cell_242_14 (.BL(BL14),.BLN(BLN14),.WL(WL242));
sram_cell_6t_5 inst_cell_242_15 (.BL(BL15),.BLN(BLN15),.WL(WL242));
sram_cell_6t_5 inst_cell_242_16 (.BL(BL16),.BLN(BLN16),.WL(WL242));
sram_cell_6t_5 inst_cell_242_17 (.BL(BL17),.BLN(BLN17),.WL(WL242));
sram_cell_6t_5 inst_cell_242_18 (.BL(BL18),.BLN(BLN18),.WL(WL242));
sram_cell_6t_5 inst_cell_242_19 (.BL(BL19),.BLN(BLN19),.WL(WL242));
sram_cell_6t_5 inst_cell_242_20 (.BL(BL20),.BLN(BLN20),.WL(WL242));
sram_cell_6t_5 inst_cell_242_21 (.BL(BL21),.BLN(BLN21),.WL(WL242));
sram_cell_6t_5 inst_cell_242_22 (.BL(BL22),.BLN(BLN22),.WL(WL242));
sram_cell_6t_5 inst_cell_242_23 (.BL(BL23),.BLN(BLN23),.WL(WL242));
sram_cell_6t_5 inst_cell_242_24 (.BL(BL24),.BLN(BLN24),.WL(WL242));
sram_cell_6t_5 inst_cell_242_25 (.BL(BL25),.BLN(BLN25),.WL(WL242));
sram_cell_6t_5 inst_cell_242_26 (.BL(BL26),.BLN(BLN26),.WL(WL242));
sram_cell_6t_5 inst_cell_242_27 (.BL(BL27),.BLN(BLN27),.WL(WL242));
sram_cell_6t_5 inst_cell_242_28 (.BL(BL28),.BLN(BLN28),.WL(WL242));
sram_cell_6t_5 inst_cell_242_29 (.BL(BL29),.BLN(BLN29),.WL(WL242));
sram_cell_6t_5 inst_cell_242_30 (.BL(BL30),.BLN(BLN30),.WL(WL242));
sram_cell_6t_5 inst_cell_242_31 (.BL(BL31),.BLN(BLN31),.WL(WL242));
sram_cell_6t_5 inst_cell_242_32 (.BL(BL32),.BLN(BLN32),.WL(WL242));
sram_cell_6t_5 inst_cell_242_33 (.BL(BL33),.BLN(BLN33),.WL(WL242));
sram_cell_6t_5 inst_cell_242_34 (.BL(BL34),.BLN(BLN34),.WL(WL242));
sram_cell_6t_5 inst_cell_242_35 (.BL(BL35),.BLN(BLN35),.WL(WL242));
sram_cell_6t_5 inst_cell_242_36 (.BL(BL36),.BLN(BLN36),.WL(WL242));
sram_cell_6t_5 inst_cell_242_37 (.BL(BL37),.BLN(BLN37),.WL(WL242));
sram_cell_6t_5 inst_cell_242_38 (.BL(BL38),.BLN(BLN38),.WL(WL242));
sram_cell_6t_5 inst_cell_242_39 (.BL(BL39),.BLN(BLN39),.WL(WL242));
sram_cell_6t_5 inst_cell_242_40 (.BL(BL40),.BLN(BLN40),.WL(WL242));
sram_cell_6t_5 inst_cell_242_41 (.BL(BL41),.BLN(BLN41),.WL(WL242));
sram_cell_6t_5 inst_cell_242_42 (.BL(BL42),.BLN(BLN42),.WL(WL242));
sram_cell_6t_5 inst_cell_242_43 (.BL(BL43),.BLN(BLN43),.WL(WL242));
sram_cell_6t_5 inst_cell_242_44 (.BL(BL44),.BLN(BLN44),.WL(WL242));
sram_cell_6t_5 inst_cell_242_45 (.BL(BL45),.BLN(BLN45),.WL(WL242));
sram_cell_6t_5 inst_cell_242_46 (.BL(BL46),.BLN(BLN46),.WL(WL242));
sram_cell_6t_5 inst_cell_242_47 (.BL(BL47),.BLN(BLN47),.WL(WL242));
sram_cell_6t_5 inst_cell_242_48 (.BL(BL48),.BLN(BLN48),.WL(WL242));
sram_cell_6t_5 inst_cell_242_49 (.BL(BL49),.BLN(BLN49),.WL(WL242));
sram_cell_6t_5 inst_cell_242_50 (.BL(BL50),.BLN(BLN50),.WL(WL242));
sram_cell_6t_5 inst_cell_242_51 (.BL(BL51),.BLN(BLN51),.WL(WL242));
sram_cell_6t_5 inst_cell_242_52 (.BL(BL52),.BLN(BLN52),.WL(WL242));
sram_cell_6t_5 inst_cell_242_53 (.BL(BL53),.BLN(BLN53),.WL(WL242));
sram_cell_6t_5 inst_cell_242_54 (.BL(BL54),.BLN(BLN54),.WL(WL242));
sram_cell_6t_5 inst_cell_242_55 (.BL(BL55),.BLN(BLN55),.WL(WL242));
sram_cell_6t_5 inst_cell_242_56 (.BL(BL56),.BLN(BLN56),.WL(WL242));
sram_cell_6t_5 inst_cell_242_57 (.BL(BL57),.BLN(BLN57),.WL(WL242));
sram_cell_6t_5 inst_cell_242_58 (.BL(BL58),.BLN(BLN58),.WL(WL242));
sram_cell_6t_5 inst_cell_242_59 (.BL(BL59),.BLN(BLN59),.WL(WL242));
sram_cell_6t_5 inst_cell_242_60 (.BL(BL60),.BLN(BLN60),.WL(WL242));
sram_cell_6t_5 inst_cell_242_61 (.BL(BL61),.BLN(BLN61),.WL(WL242));
sram_cell_6t_5 inst_cell_242_62 (.BL(BL62),.BLN(BLN62),.WL(WL242));
sram_cell_6t_5 inst_cell_242_63 (.BL(BL63),.BLN(BLN63),.WL(WL242));
sram_cell_6t_5 inst_cell_242_64 (.BL(BL64),.BLN(BLN64),.WL(WL242));
sram_cell_6t_5 inst_cell_242_65 (.BL(BL65),.BLN(BLN65),.WL(WL242));
sram_cell_6t_5 inst_cell_242_66 (.BL(BL66),.BLN(BLN66),.WL(WL242));
sram_cell_6t_5 inst_cell_242_67 (.BL(BL67),.BLN(BLN67),.WL(WL242));
sram_cell_6t_5 inst_cell_242_68 (.BL(BL68),.BLN(BLN68),.WL(WL242));
sram_cell_6t_5 inst_cell_242_69 (.BL(BL69),.BLN(BLN69),.WL(WL242));
sram_cell_6t_5 inst_cell_242_70 (.BL(BL70),.BLN(BLN70),.WL(WL242));
sram_cell_6t_5 inst_cell_242_71 (.BL(BL71),.BLN(BLN71),.WL(WL242));
sram_cell_6t_5 inst_cell_242_72 (.BL(BL72),.BLN(BLN72),.WL(WL242));
sram_cell_6t_5 inst_cell_242_73 (.BL(BL73),.BLN(BLN73),.WL(WL242));
sram_cell_6t_5 inst_cell_242_74 (.BL(BL74),.BLN(BLN74),.WL(WL242));
sram_cell_6t_5 inst_cell_242_75 (.BL(BL75),.BLN(BLN75),.WL(WL242));
sram_cell_6t_5 inst_cell_242_76 (.BL(BL76),.BLN(BLN76),.WL(WL242));
sram_cell_6t_5 inst_cell_242_77 (.BL(BL77),.BLN(BLN77),.WL(WL242));
sram_cell_6t_5 inst_cell_242_78 (.BL(BL78),.BLN(BLN78),.WL(WL242));
sram_cell_6t_5 inst_cell_242_79 (.BL(BL79),.BLN(BLN79),.WL(WL242));
sram_cell_6t_5 inst_cell_242_80 (.BL(BL80),.BLN(BLN80),.WL(WL242));
sram_cell_6t_5 inst_cell_242_81 (.BL(BL81),.BLN(BLN81),.WL(WL242));
sram_cell_6t_5 inst_cell_242_82 (.BL(BL82),.BLN(BLN82),.WL(WL242));
sram_cell_6t_5 inst_cell_242_83 (.BL(BL83),.BLN(BLN83),.WL(WL242));
sram_cell_6t_5 inst_cell_242_84 (.BL(BL84),.BLN(BLN84),.WL(WL242));
sram_cell_6t_5 inst_cell_242_85 (.BL(BL85),.BLN(BLN85),.WL(WL242));
sram_cell_6t_5 inst_cell_242_86 (.BL(BL86),.BLN(BLN86),.WL(WL242));
sram_cell_6t_5 inst_cell_242_87 (.BL(BL87),.BLN(BLN87),.WL(WL242));
sram_cell_6t_5 inst_cell_242_88 (.BL(BL88),.BLN(BLN88),.WL(WL242));
sram_cell_6t_5 inst_cell_242_89 (.BL(BL89),.BLN(BLN89),.WL(WL242));
sram_cell_6t_5 inst_cell_242_90 (.BL(BL90),.BLN(BLN90),.WL(WL242));
sram_cell_6t_5 inst_cell_242_91 (.BL(BL91),.BLN(BLN91),.WL(WL242));
sram_cell_6t_5 inst_cell_242_92 (.BL(BL92),.BLN(BLN92),.WL(WL242));
sram_cell_6t_5 inst_cell_242_93 (.BL(BL93),.BLN(BLN93),.WL(WL242));
sram_cell_6t_5 inst_cell_242_94 (.BL(BL94),.BLN(BLN94),.WL(WL242));
sram_cell_6t_5 inst_cell_242_95 (.BL(BL95),.BLN(BLN95),.WL(WL242));
sram_cell_6t_5 inst_cell_242_96 (.BL(BL96),.BLN(BLN96),.WL(WL242));
sram_cell_6t_5 inst_cell_242_97 (.BL(BL97),.BLN(BLN97),.WL(WL242));
sram_cell_6t_5 inst_cell_242_98 (.BL(BL98),.BLN(BLN98),.WL(WL242));
sram_cell_6t_5 inst_cell_242_99 (.BL(BL99),.BLN(BLN99),.WL(WL242));
sram_cell_6t_5 inst_cell_242_100 (.BL(BL100),.BLN(BLN100),.WL(WL242));
sram_cell_6t_5 inst_cell_242_101 (.BL(BL101),.BLN(BLN101),.WL(WL242));
sram_cell_6t_5 inst_cell_242_102 (.BL(BL102),.BLN(BLN102),.WL(WL242));
sram_cell_6t_5 inst_cell_242_103 (.BL(BL103),.BLN(BLN103),.WL(WL242));
sram_cell_6t_5 inst_cell_242_104 (.BL(BL104),.BLN(BLN104),.WL(WL242));
sram_cell_6t_5 inst_cell_242_105 (.BL(BL105),.BLN(BLN105),.WL(WL242));
sram_cell_6t_5 inst_cell_242_106 (.BL(BL106),.BLN(BLN106),.WL(WL242));
sram_cell_6t_5 inst_cell_242_107 (.BL(BL107),.BLN(BLN107),.WL(WL242));
sram_cell_6t_5 inst_cell_242_108 (.BL(BL108),.BLN(BLN108),.WL(WL242));
sram_cell_6t_5 inst_cell_242_109 (.BL(BL109),.BLN(BLN109),.WL(WL242));
sram_cell_6t_5 inst_cell_242_110 (.BL(BL110),.BLN(BLN110),.WL(WL242));
sram_cell_6t_5 inst_cell_242_111 (.BL(BL111),.BLN(BLN111),.WL(WL242));
sram_cell_6t_5 inst_cell_242_112 (.BL(BL112),.BLN(BLN112),.WL(WL242));
sram_cell_6t_5 inst_cell_242_113 (.BL(BL113),.BLN(BLN113),.WL(WL242));
sram_cell_6t_5 inst_cell_242_114 (.BL(BL114),.BLN(BLN114),.WL(WL242));
sram_cell_6t_5 inst_cell_242_115 (.BL(BL115),.BLN(BLN115),.WL(WL242));
sram_cell_6t_5 inst_cell_242_116 (.BL(BL116),.BLN(BLN116),.WL(WL242));
sram_cell_6t_5 inst_cell_242_117 (.BL(BL117),.BLN(BLN117),.WL(WL242));
sram_cell_6t_5 inst_cell_242_118 (.BL(BL118),.BLN(BLN118),.WL(WL242));
sram_cell_6t_5 inst_cell_242_119 (.BL(BL119),.BLN(BLN119),.WL(WL242));
sram_cell_6t_5 inst_cell_242_120 (.BL(BL120),.BLN(BLN120),.WL(WL242));
sram_cell_6t_5 inst_cell_242_121 (.BL(BL121),.BLN(BLN121),.WL(WL242));
sram_cell_6t_5 inst_cell_242_122 (.BL(BL122),.BLN(BLN122),.WL(WL242));
sram_cell_6t_5 inst_cell_242_123 (.BL(BL123),.BLN(BLN123),.WL(WL242));
sram_cell_6t_5 inst_cell_242_124 (.BL(BL124),.BLN(BLN124),.WL(WL242));
sram_cell_6t_5 inst_cell_242_125 (.BL(BL125),.BLN(BLN125),.WL(WL242));
sram_cell_6t_5 inst_cell_242_126 (.BL(BL126),.BLN(BLN126),.WL(WL242));
sram_cell_6t_5 inst_cell_242_127 (.BL(BL127),.BLN(BLN127),.WL(WL242));
sram_cell_6t_5 inst_cell_243_0 (.BL(BL0),.BLN(BLN0),.WL(WL243));
sram_cell_6t_5 inst_cell_243_1 (.BL(BL1),.BLN(BLN1),.WL(WL243));
sram_cell_6t_5 inst_cell_243_2 (.BL(BL2),.BLN(BLN2),.WL(WL243));
sram_cell_6t_5 inst_cell_243_3 (.BL(BL3),.BLN(BLN3),.WL(WL243));
sram_cell_6t_5 inst_cell_243_4 (.BL(BL4),.BLN(BLN4),.WL(WL243));
sram_cell_6t_5 inst_cell_243_5 (.BL(BL5),.BLN(BLN5),.WL(WL243));
sram_cell_6t_5 inst_cell_243_6 (.BL(BL6),.BLN(BLN6),.WL(WL243));
sram_cell_6t_5 inst_cell_243_7 (.BL(BL7),.BLN(BLN7),.WL(WL243));
sram_cell_6t_5 inst_cell_243_8 (.BL(BL8),.BLN(BLN8),.WL(WL243));
sram_cell_6t_5 inst_cell_243_9 (.BL(BL9),.BLN(BLN9),.WL(WL243));
sram_cell_6t_5 inst_cell_243_10 (.BL(BL10),.BLN(BLN10),.WL(WL243));
sram_cell_6t_5 inst_cell_243_11 (.BL(BL11),.BLN(BLN11),.WL(WL243));
sram_cell_6t_5 inst_cell_243_12 (.BL(BL12),.BLN(BLN12),.WL(WL243));
sram_cell_6t_5 inst_cell_243_13 (.BL(BL13),.BLN(BLN13),.WL(WL243));
sram_cell_6t_5 inst_cell_243_14 (.BL(BL14),.BLN(BLN14),.WL(WL243));
sram_cell_6t_5 inst_cell_243_15 (.BL(BL15),.BLN(BLN15),.WL(WL243));
sram_cell_6t_5 inst_cell_243_16 (.BL(BL16),.BLN(BLN16),.WL(WL243));
sram_cell_6t_5 inst_cell_243_17 (.BL(BL17),.BLN(BLN17),.WL(WL243));
sram_cell_6t_5 inst_cell_243_18 (.BL(BL18),.BLN(BLN18),.WL(WL243));
sram_cell_6t_5 inst_cell_243_19 (.BL(BL19),.BLN(BLN19),.WL(WL243));
sram_cell_6t_5 inst_cell_243_20 (.BL(BL20),.BLN(BLN20),.WL(WL243));
sram_cell_6t_5 inst_cell_243_21 (.BL(BL21),.BLN(BLN21),.WL(WL243));
sram_cell_6t_5 inst_cell_243_22 (.BL(BL22),.BLN(BLN22),.WL(WL243));
sram_cell_6t_5 inst_cell_243_23 (.BL(BL23),.BLN(BLN23),.WL(WL243));
sram_cell_6t_5 inst_cell_243_24 (.BL(BL24),.BLN(BLN24),.WL(WL243));
sram_cell_6t_5 inst_cell_243_25 (.BL(BL25),.BLN(BLN25),.WL(WL243));
sram_cell_6t_5 inst_cell_243_26 (.BL(BL26),.BLN(BLN26),.WL(WL243));
sram_cell_6t_5 inst_cell_243_27 (.BL(BL27),.BLN(BLN27),.WL(WL243));
sram_cell_6t_5 inst_cell_243_28 (.BL(BL28),.BLN(BLN28),.WL(WL243));
sram_cell_6t_5 inst_cell_243_29 (.BL(BL29),.BLN(BLN29),.WL(WL243));
sram_cell_6t_5 inst_cell_243_30 (.BL(BL30),.BLN(BLN30),.WL(WL243));
sram_cell_6t_5 inst_cell_243_31 (.BL(BL31),.BLN(BLN31),.WL(WL243));
sram_cell_6t_5 inst_cell_243_32 (.BL(BL32),.BLN(BLN32),.WL(WL243));
sram_cell_6t_5 inst_cell_243_33 (.BL(BL33),.BLN(BLN33),.WL(WL243));
sram_cell_6t_5 inst_cell_243_34 (.BL(BL34),.BLN(BLN34),.WL(WL243));
sram_cell_6t_5 inst_cell_243_35 (.BL(BL35),.BLN(BLN35),.WL(WL243));
sram_cell_6t_5 inst_cell_243_36 (.BL(BL36),.BLN(BLN36),.WL(WL243));
sram_cell_6t_5 inst_cell_243_37 (.BL(BL37),.BLN(BLN37),.WL(WL243));
sram_cell_6t_5 inst_cell_243_38 (.BL(BL38),.BLN(BLN38),.WL(WL243));
sram_cell_6t_5 inst_cell_243_39 (.BL(BL39),.BLN(BLN39),.WL(WL243));
sram_cell_6t_5 inst_cell_243_40 (.BL(BL40),.BLN(BLN40),.WL(WL243));
sram_cell_6t_5 inst_cell_243_41 (.BL(BL41),.BLN(BLN41),.WL(WL243));
sram_cell_6t_5 inst_cell_243_42 (.BL(BL42),.BLN(BLN42),.WL(WL243));
sram_cell_6t_5 inst_cell_243_43 (.BL(BL43),.BLN(BLN43),.WL(WL243));
sram_cell_6t_5 inst_cell_243_44 (.BL(BL44),.BLN(BLN44),.WL(WL243));
sram_cell_6t_5 inst_cell_243_45 (.BL(BL45),.BLN(BLN45),.WL(WL243));
sram_cell_6t_5 inst_cell_243_46 (.BL(BL46),.BLN(BLN46),.WL(WL243));
sram_cell_6t_5 inst_cell_243_47 (.BL(BL47),.BLN(BLN47),.WL(WL243));
sram_cell_6t_5 inst_cell_243_48 (.BL(BL48),.BLN(BLN48),.WL(WL243));
sram_cell_6t_5 inst_cell_243_49 (.BL(BL49),.BLN(BLN49),.WL(WL243));
sram_cell_6t_5 inst_cell_243_50 (.BL(BL50),.BLN(BLN50),.WL(WL243));
sram_cell_6t_5 inst_cell_243_51 (.BL(BL51),.BLN(BLN51),.WL(WL243));
sram_cell_6t_5 inst_cell_243_52 (.BL(BL52),.BLN(BLN52),.WL(WL243));
sram_cell_6t_5 inst_cell_243_53 (.BL(BL53),.BLN(BLN53),.WL(WL243));
sram_cell_6t_5 inst_cell_243_54 (.BL(BL54),.BLN(BLN54),.WL(WL243));
sram_cell_6t_5 inst_cell_243_55 (.BL(BL55),.BLN(BLN55),.WL(WL243));
sram_cell_6t_5 inst_cell_243_56 (.BL(BL56),.BLN(BLN56),.WL(WL243));
sram_cell_6t_5 inst_cell_243_57 (.BL(BL57),.BLN(BLN57),.WL(WL243));
sram_cell_6t_5 inst_cell_243_58 (.BL(BL58),.BLN(BLN58),.WL(WL243));
sram_cell_6t_5 inst_cell_243_59 (.BL(BL59),.BLN(BLN59),.WL(WL243));
sram_cell_6t_5 inst_cell_243_60 (.BL(BL60),.BLN(BLN60),.WL(WL243));
sram_cell_6t_5 inst_cell_243_61 (.BL(BL61),.BLN(BLN61),.WL(WL243));
sram_cell_6t_5 inst_cell_243_62 (.BL(BL62),.BLN(BLN62),.WL(WL243));
sram_cell_6t_5 inst_cell_243_63 (.BL(BL63),.BLN(BLN63),.WL(WL243));
sram_cell_6t_5 inst_cell_243_64 (.BL(BL64),.BLN(BLN64),.WL(WL243));
sram_cell_6t_5 inst_cell_243_65 (.BL(BL65),.BLN(BLN65),.WL(WL243));
sram_cell_6t_5 inst_cell_243_66 (.BL(BL66),.BLN(BLN66),.WL(WL243));
sram_cell_6t_5 inst_cell_243_67 (.BL(BL67),.BLN(BLN67),.WL(WL243));
sram_cell_6t_5 inst_cell_243_68 (.BL(BL68),.BLN(BLN68),.WL(WL243));
sram_cell_6t_5 inst_cell_243_69 (.BL(BL69),.BLN(BLN69),.WL(WL243));
sram_cell_6t_5 inst_cell_243_70 (.BL(BL70),.BLN(BLN70),.WL(WL243));
sram_cell_6t_5 inst_cell_243_71 (.BL(BL71),.BLN(BLN71),.WL(WL243));
sram_cell_6t_5 inst_cell_243_72 (.BL(BL72),.BLN(BLN72),.WL(WL243));
sram_cell_6t_5 inst_cell_243_73 (.BL(BL73),.BLN(BLN73),.WL(WL243));
sram_cell_6t_5 inst_cell_243_74 (.BL(BL74),.BLN(BLN74),.WL(WL243));
sram_cell_6t_5 inst_cell_243_75 (.BL(BL75),.BLN(BLN75),.WL(WL243));
sram_cell_6t_5 inst_cell_243_76 (.BL(BL76),.BLN(BLN76),.WL(WL243));
sram_cell_6t_5 inst_cell_243_77 (.BL(BL77),.BLN(BLN77),.WL(WL243));
sram_cell_6t_5 inst_cell_243_78 (.BL(BL78),.BLN(BLN78),.WL(WL243));
sram_cell_6t_5 inst_cell_243_79 (.BL(BL79),.BLN(BLN79),.WL(WL243));
sram_cell_6t_5 inst_cell_243_80 (.BL(BL80),.BLN(BLN80),.WL(WL243));
sram_cell_6t_5 inst_cell_243_81 (.BL(BL81),.BLN(BLN81),.WL(WL243));
sram_cell_6t_5 inst_cell_243_82 (.BL(BL82),.BLN(BLN82),.WL(WL243));
sram_cell_6t_5 inst_cell_243_83 (.BL(BL83),.BLN(BLN83),.WL(WL243));
sram_cell_6t_5 inst_cell_243_84 (.BL(BL84),.BLN(BLN84),.WL(WL243));
sram_cell_6t_5 inst_cell_243_85 (.BL(BL85),.BLN(BLN85),.WL(WL243));
sram_cell_6t_5 inst_cell_243_86 (.BL(BL86),.BLN(BLN86),.WL(WL243));
sram_cell_6t_5 inst_cell_243_87 (.BL(BL87),.BLN(BLN87),.WL(WL243));
sram_cell_6t_5 inst_cell_243_88 (.BL(BL88),.BLN(BLN88),.WL(WL243));
sram_cell_6t_5 inst_cell_243_89 (.BL(BL89),.BLN(BLN89),.WL(WL243));
sram_cell_6t_5 inst_cell_243_90 (.BL(BL90),.BLN(BLN90),.WL(WL243));
sram_cell_6t_5 inst_cell_243_91 (.BL(BL91),.BLN(BLN91),.WL(WL243));
sram_cell_6t_5 inst_cell_243_92 (.BL(BL92),.BLN(BLN92),.WL(WL243));
sram_cell_6t_5 inst_cell_243_93 (.BL(BL93),.BLN(BLN93),.WL(WL243));
sram_cell_6t_5 inst_cell_243_94 (.BL(BL94),.BLN(BLN94),.WL(WL243));
sram_cell_6t_5 inst_cell_243_95 (.BL(BL95),.BLN(BLN95),.WL(WL243));
sram_cell_6t_5 inst_cell_243_96 (.BL(BL96),.BLN(BLN96),.WL(WL243));
sram_cell_6t_5 inst_cell_243_97 (.BL(BL97),.BLN(BLN97),.WL(WL243));
sram_cell_6t_5 inst_cell_243_98 (.BL(BL98),.BLN(BLN98),.WL(WL243));
sram_cell_6t_5 inst_cell_243_99 (.BL(BL99),.BLN(BLN99),.WL(WL243));
sram_cell_6t_5 inst_cell_243_100 (.BL(BL100),.BLN(BLN100),.WL(WL243));
sram_cell_6t_5 inst_cell_243_101 (.BL(BL101),.BLN(BLN101),.WL(WL243));
sram_cell_6t_5 inst_cell_243_102 (.BL(BL102),.BLN(BLN102),.WL(WL243));
sram_cell_6t_5 inst_cell_243_103 (.BL(BL103),.BLN(BLN103),.WL(WL243));
sram_cell_6t_5 inst_cell_243_104 (.BL(BL104),.BLN(BLN104),.WL(WL243));
sram_cell_6t_5 inst_cell_243_105 (.BL(BL105),.BLN(BLN105),.WL(WL243));
sram_cell_6t_5 inst_cell_243_106 (.BL(BL106),.BLN(BLN106),.WL(WL243));
sram_cell_6t_5 inst_cell_243_107 (.BL(BL107),.BLN(BLN107),.WL(WL243));
sram_cell_6t_5 inst_cell_243_108 (.BL(BL108),.BLN(BLN108),.WL(WL243));
sram_cell_6t_5 inst_cell_243_109 (.BL(BL109),.BLN(BLN109),.WL(WL243));
sram_cell_6t_5 inst_cell_243_110 (.BL(BL110),.BLN(BLN110),.WL(WL243));
sram_cell_6t_5 inst_cell_243_111 (.BL(BL111),.BLN(BLN111),.WL(WL243));
sram_cell_6t_5 inst_cell_243_112 (.BL(BL112),.BLN(BLN112),.WL(WL243));
sram_cell_6t_5 inst_cell_243_113 (.BL(BL113),.BLN(BLN113),.WL(WL243));
sram_cell_6t_5 inst_cell_243_114 (.BL(BL114),.BLN(BLN114),.WL(WL243));
sram_cell_6t_5 inst_cell_243_115 (.BL(BL115),.BLN(BLN115),.WL(WL243));
sram_cell_6t_5 inst_cell_243_116 (.BL(BL116),.BLN(BLN116),.WL(WL243));
sram_cell_6t_5 inst_cell_243_117 (.BL(BL117),.BLN(BLN117),.WL(WL243));
sram_cell_6t_5 inst_cell_243_118 (.BL(BL118),.BLN(BLN118),.WL(WL243));
sram_cell_6t_5 inst_cell_243_119 (.BL(BL119),.BLN(BLN119),.WL(WL243));
sram_cell_6t_5 inst_cell_243_120 (.BL(BL120),.BLN(BLN120),.WL(WL243));
sram_cell_6t_5 inst_cell_243_121 (.BL(BL121),.BLN(BLN121),.WL(WL243));
sram_cell_6t_5 inst_cell_243_122 (.BL(BL122),.BLN(BLN122),.WL(WL243));
sram_cell_6t_5 inst_cell_243_123 (.BL(BL123),.BLN(BLN123),.WL(WL243));
sram_cell_6t_5 inst_cell_243_124 (.BL(BL124),.BLN(BLN124),.WL(WL243));
sram_cell_6t_5 inst_cell_243_125 (.BL(BL125),.BLN(BLN125),.WL(WL243));
sram_cell_6t_5 inst_cell_243_126 (.BL(BL126),.BLN(BLN126),.WL(WL243));
sram_cell_6t_5 inst_cell_243_127 (.BL(BL127),.BLN(BLN127),.WL(WL243));
sram_cell_6t_5 inst_cell_244_0 (.BL(BL0),.BLN(BLN0),.WL(WL244));
sram_cell_6t_5 inst_cell_244_1 (.BL(BL1),.BLN(BLN1),.WL(WL244));
sram_cell_6t_5 inst_cell_244_2 (.BL(BL2),.BLN(BLN2),.WL(WL244));
sram_cell_6t_5 inst_cell_244_3 (.BL(BL3),.BLN(BLN3),.WL(WL244));
sram_cell_6t_5 inst_cell_244_4 (.BL(BL4),.BLN(BLN4),.WL(WL244));
sram_cell_6t_5 inst_cell_244_5 (.BL(BL5),.BLN(BLN5),.WL(WL244));
sram_cell_6t_5 inst_cell_244_6 (.BL(BL6),.BLN(BLN6),.WL(WL244));
sram_cell_6t_5 inst_cell_244_7 (.BL(BL7),.BLN(BLN7),.WL(WL244));
sram_cell_6t_5 inst_cell_244_8 (.BL(BL8),.BLN(BLN8),.WL(WL244));
sram_cell_6t_5 inst_cell_244_9 (.BL(BL9),.BLN(BLN9),.WL(WL244));
sram_cell_6t_5 inst_cell_244_10 (.BL(BL10),.BLN(BLN10),.WL(WL244));
sram_cell_6t_5 inst_cell_244_11 (.BL(BL11),.BLN(BLN11),.WL(WL244));
sram_cell_6t_5 inst_cell_244_12 (.BL(BL12),.BLN(BLN12),.WL(WL244));
sram_cell_6t_5 inst_cell_244_13 (.BL(BL13),.BLN(BLN13),.WL(WL244));
sram_cell_6t_5 inst_cell_244_14 (.BL(BL14),.BLN(BLN14),.WL(WL244));
sram_cell_6t_5 inst_cell_244_15 (.BL(BL15),.BLN(BLN15),.WL(WL244));
sram_cell_6t_5 inst_cell_244_16 (.BL(BL16),.BLN(BLN16),.WL(WL244));
sram_cell_6t_5 inst_cell_244_17 (.BL(BL17),.BLN(BLN17),.WL(WL244));
sram_cell_6t_5 inst_cell_244_18 (.BL(BL18),.BLN(BLN18),.WL(WL244));
sram_cell_6t_5 inst_cell_244_19 (.BL(BL19),.BLN(BLN19),.WL(WL244));
sram_cell_6t_5 inst_cell_244_20 (.BL(BL20),.BLN(BLN20),.WL(WL244));
sram_cell_6t_5 inst_cell_244_21 (.BL(BL21),.BLN(BLN21),.WL(WL244));
sram_cell_6t_5 inst_cell_244_22 (.BL(BL22),.BLN(BLN22),.WL(WL244));
sram_cell_6t_5 inst_cell_244_23 (.BL(BL23),.BLN(BLN23),.WL(WL244));
sram_cell_6t_5 inst_cell_244_24 (.BL(BL24),.BLN(BLN24),.WL(WL244));
sram_cell_6t_5 inst_cell_244_25 (.BL(BL25),.BLN(BLN25),.WL(WL244));
sram_cell_6t_5 inst_cell_244_26 (.BL(BL26),.BLN(BLN26),.WL(WL244));
sram_cell_6t_5 inst_cell_244_27 (.BL(BL27),.BLN(BLN27),.WL(WL244));
sram_cell_6t_5 inst_cell_244_28 (.BL(BL28),.BLN(BLN28),.WL(WL244));
sram_cell_6t_5 inst_cell_244_29 (.BL(BL29),.BLN(BLN29),.WL(WL244));
sram_cell_6t_5 inst_cell_244_30 (.BL(BL30),.BLN(BLN30),.WL(WL244));
sram_cell_6t_5 inst_cell_244_31 (.BL(BL31),.BLN(BLN31),.WL(WL244));
sram_cell_6t_5 inst_cell_244_32 (.BL(BL32),.BLN(BLN32),.WL(WL244));
sram_cell_6t_5 inst_cell_244_33 (.BL(BL33),.BLN(BLN33),.WL(WL244));
sram_cell_6t_5 inst_cell_244_34 (.BL(BL34),.BLN(BLN34),.WL(WL244));
sram_cell_6t_5 inst_cell_244_35 (.BL(BL35),.BLN(BLN35),.WL(WL244));
sram_cell_6t_5 inst_cell_244_36 (.BL(BL36),.BLN(BLN36),.WL(WL244));
sram_cell_6t_5 inst_cell_244_37 (.BL(BL37),.BLN(BLN37),.WL(WL244));
sram_cell_6t_5 inst_cell_244_38 (.BL(BL38),.BLN(BLN38),.WL(WL244));
sram_cell_6t_5 inst_cell_244_39 (.BL(BL39),.BLN(BLN39),.WL(WL244));
sram_cell_6t_5 inst_cell_244_40 (.BL(BL40),.BLN(BLN40),.WL(WL244));
sram_cell_6t_5 inst_cell_244_41 (.BL(BL41),.BLN(BLN41),.WL(WL244));
sram_cell_6t_5 inst_cell_244_42 (.BL(BL42),.BLN(BLN42),.WL(WL244));
sram_cell_6t_5 inst_cell_244_43 (.BL(BL43),.BLN(BLN43),.WL(WL244));
sram_cell_6t_5 inst_cell_244_44 (.BL(BL44),.BLN(BLN44),.WL(WL244));
sram_cell_6t_5 inst_cell_244_45 (.BL(BL45),.BLN(BLN45),.WL(WL244));
sram_cell_6t_5 inst_cell_244_46 (.BL(BL46),.BLN(BLN46),.WL(WL244));
sram_cell_6t_5 inst_cell_244_47 (.BL(BL47),.BLN(BLN47),.WL(WL244));
sram_cell_6t_5 inst_cell_244_48 (.BL(BL48),.BLN(BLN48),.WL(WL244));
sram_cell_6t_5 inst_cell_244_49 (.BL(BL49),.BLN(BLN49),.WL(WL244));
sram_cell_6t_5 inst_cell_244_50 (.BL(BL50),.BLN(BLN50),.WL(WL244));
sram_cell_6t_5 inst_cell_244_51 (.BL(BL51),.BLN(BLN51),.WL(WL244));
sram_cell_6t_5 inst_cell_244_52 (.BL(BL52),.BLN(BLN52),.WL(WL244));
sram_cell_6t_5 inst_cell_244_53 (.BL(BL53),.BLN(BLN53),.WL(WL244));
sram_cell_6t_5 inst_cell_244_54 (.BL(BL54),.BLN(BLN54),.WL(WL244));
sram_cell_6t_5 inst_cell_244_55 (.BL(BL55),.BLN(BLN55),.WL(WL244));
sram_cell_6t_5 inst_cell_244_56 (.BL(BL56),.BLN(BLN56),.WL(WL244));
sram_cell_6t_5 inst_cell_244_57 (.BL(BL57),.BLN(BLN57),.WL(WL244));
sram_cell_6t_5 inst_cell_244_58 (.BL(BL58),.BLN(BLN58),.WL(WL244));
sram_cell_6t_5 inst_cell_244_59 (.BL(BL59),.BLN(BLN59),.WL(WL244));
sram_cell_6t_5 inst_cell_244_60 (.BL(BL60),.BLN(BLN60),.WL(WL244));
sram_cell_6t_5 inst_cell_244_61 (.BL(BL61),.BLN(BLN61),.WL(WL244));
sram_cell_6t_5 inst_cell_244_62 (.BL(BL62),.BLN(BLN62),.WL(WL244));
sram_cell_6t_5 inst_cell_244_63 (.BL(BL63),.BLN(BLN63),.WL(WL244));
sram_cell_6t_5 inst_cell_244_64 (.BL(BL64),.BLN(BLN64),.WL(WL244));
sram_cell_6t_5 inst_cell_244_65 (.BL(BL65),.BLN(BLN65),.WL(WL244));
sram_cell_6t_5 inst_cell_244_66 (.BL(BL66),.BLN(BLN66),.WL(WL244));
sram_cell_6t_5 inst_cell_244_67 (.BL(BL67),.BLN(BLN67),.WL(WL244));
sram_cell_6t_5 inst_cell_244_68 (.BL(BL68),.BLN(BLN68),.WL(WL244));
sram_cell_6t_5 inst_cell_244_69 (.BL(BL69),.BLN(BLN69),.WL(WL244));
sram_cell_6t_5 inst_cell_244_70 (.BL(BL70),.BLN(BLN70),.WL(WL244));
sram_cell_6t_5 inst_cell_244_71 (.BL(BL71),.BLN(BLN71),.WL(WL244));
sram_cell_6t_5 inst_cell_244_72 (.BL(BL72),.BLN(BLN72),.WL(WL244));
sram_cell_6t_5 inst_cell_244_73 (.BL(BL73),.BLN(BLN73),.WL(WL244));
sram_cell_6t_5 inst_cell_244_74 (.BL(BL74),.BLN(BLN74),.WL(WL244));
sram_cell_6t_5 inst_cell_244_75 (.BL(BL75),.BLN(BLN75),.WL(WL244));
sram_cell_6t_5 inst_cell_244_76 (.BL(BL76),.BLN(BLN76),.WL(WL244));
sram_cell_6t_5 inst_cell_244_77 (.BL(BL77),.BLN(BLN77),.WL(WL244));
sram_cell_6t_5 inst_cell_244_78 (.BL(BL78),.BLN(BLN78),.WL(WL244));
sram_cell_6t_5 inst_cell_244_79 (.BL(BL79),.BLN(BLN79),.WL(WL244));
sram_cell_6t_5 inst_cell_244_80 (.BL(BL80),.BLN(BLN80),.WL(WL244));
sram_cell_6t_5 inst_cell_244_81 (.BL(BL81),.BLN(BLN81),.WL(WL244));
sram_cell_6t_5 inst_cell_244_82 (.BL(BL82),.BLN(BLN82),.WL(WL244));
sram_cell_6t_5 inst_cell_244_83 (.BL(BL83),.BLN(BLN83),.WL(WL244));
sram_cell_6t_5 inst_cell_244_84 (.BL(BL84),.BLN(BLN84),.WL(WL244));
sram_cell_6t_5 inst_cell_244_85 (.BL(BL85),.BLN(BLN85),.WL(WL244));
sram_cell_6t_5 inst_cell_244_86 (.BL(BL86),.BLN(BLN86),.WL(WL244));
sram_cell_6t_5 inst_cell_244_87 (.BL(BL87),.BLN(BLN87),.WL(WL244));
sram_cell_6t_5 inst_cell_244_88 (.BL(BL88),.BLN(BLN88),.WL(WL244));
sram_cell_6t_5 inst_cell_244_89 (.BL(BL89),.BLN(BLN89),.WL(WL244));
sram_cell_6t_5 inst_cell_244_90 (.BL(BL90),.BLN(BLN90),.WL(WL244));
sram_cell_6t_5 inst_cell_244_91 (.BL(BL91),.BLN(BLN91),.WL(WL244));
sram_cell_6t_5 inst_cell_244_92 (.BL(BL92),.BLN(BLN92),.WL(WL244));
sram_cell_6t_5 inst_cell_244_93 (.BL(BL93),.BLN(BLN93),.WL(WL244));
sram_cell_6t_5 inst_cell_244_94 (.BL(BL94),.BLN(BLN94),.WL(WL244));
sram_cell_6t_5 inst_cell_244_95 (.BL(BL95),.BLN(BLN95),.WL(WL244));
sram_cell_6t_5 inst_cell_244_96 (.BL(BL96),.BLN(BLN96),.WL(WL244));
sram_cell_6t_5 inst_cell_244_97 (.BL(BL97),.BLN(BLN97),.WL(WL244));
sram_cell_6t_5 inst_cell_244_98 (.BL(BL98),.BLN(BLN98),.WL(WL244));
sram_cell_6t_5 inst_cell_244_99 (.BL(BL99),.BLN(BLN99),.WL(WL244));
sram_cell_6t_5 inst_cell_244_100 (.BL(BL100),.BLN(BLN100),.WL(WL244));
sram_cell_6t_5 inst_cell_244_101 (.BL(BL101),.BLN(BLN101),.WL(WL244));
sram_cell_6t_5 inst_cell_244_102 (.BL(BL102),.BLN(BLN102),.WL(WL244));
sram_cell_6t_5 inst_cell_244_103 (.BL(BL103),.BLN(BLN103),.WL(WL244));
sram_cell_6t_5 inst_cell_244_104 (.BL(BL104),.BLN(BLN104),.WL(WL244));
sram_cell_6t_5 inst_cell_244_105 (.BL(BL105),.BLN(BLN105),.WL(WL244));
sram_cell_6t_5 inst_cell_244_106 (.BL(BL106),.BLN(BLN106),.WL(WL244));
sram_cell_6t_5 inst_cell_244_107 (.BL(BL107),.BLN(BLN107),.WL(WL244));
sram_cell_6t_5 inst_cell_244_108 (.BL(BL108),.BLN(BLN108),.WL(WL244));
sram_cell_6t_5 inst_cell_244_109 (.BL(BL109),.BLN(BLN109),.WL(WL244));
sram_cell_6t_5 inst_cell_244_110 (.BL(BL110),.BLN(BLN110),.WL(WL244));
sram_cell_6t_5 inst_cell_244_111 (.BL(BL111),.BLN(BLN111),.WL(WL244));
sram_cell_6t_5 inst_cell_244_112 (.BL(BL112),.BLN(BLN112),.WL(WL244));
sram_cell_6t_5 inst_cell_244_113 (.BL(BL113),.BLN(BLN113),.WL(WL244));
sram_cell_6t_5 inst_cell_244_114 (.BL(BL114),.BLN(BLN114),.WL(WL244));
sram_cell_6t_5 inst_cell_244_115 (.BL(BL115),.BLN(BLN115),.WL(WL244));
sram_cell_6t_5 inst_cell_244_116 (.BL(BL116),.BLN(BLN116),.WL(WL244));
sram_cell_6t_5 inst_cell_244_117 (.BL(BL117),.BLN(BLN117),.WL(WL244));
sram_cell_6t_5 inst_cell_244_118 (.BL(BL118),.BLN(BLN118),.WL(WL244));
sram_cell_6t_5 inst_cell_244_119 (.BL(BL119),.BLN(BLN119),.WL(WL244));
sram_cell_6t_5 inst_cell_244_120 (.BL(BL120),.BLN(BLN120),.WL(WL244));
sram_cell_6t_5 inst_cell_244_121 (.BL(BL121),.BLN(BLN121),.WL(WL244));
sram_cell_6t_5 inst_cell_244_122 (.BL(BL122),.BLN(BLN122),.WL(WL244));
sram_cell_6t_5 inst_cell_244_123 (.BL(BL123),.BLN(BLN123),.WL(WL244));
sram_cell_6t_5 inst_cell_244_124 (.BL(BL124),.BLN(BLN124),.WL(WL244));
sram_cell_6t_5 inst_cell_244_125 (.BL(BL125),.BLN(BLN125),.WL(WL244));
sram_cell_6t_5 inst_cell_244_126 (.BL(BL126),.BLN(BLN126),.WL(WL244));
sram_cell_6t_5 inst_cell_244_127 (.BL(BL127),.BLN(BLN127),.WL(WL244));
sram_cell_6t_5 inst_cell_245_0 (.BL(BL0),.BLN(BLN0),.WL(WL245));
sram_cell_6t_5 inst_cell_245_1 (.BL(BL1),.BLN(BLN1),.WL(WL245));
sram_cell_6t_5 inst_cell_245_2 (.BL(BL2),.BLN(BLN2),.WL(WL245));
sram_cell_6t_5 inst_cell_245_3 (.BL(BL3),.BLN(BLN3),.WL(WL245));
sram_cell_6t_5 inst_cell_245_4 (.BL(BL4),.BLN(BLN4),.WL(WL245));
sram_cell_6t_5 inst_cell_245_5 (.BL(BL5),.BLN(BLN5),.WL(WL245));
sram_cell_6t_5 inst_cell_245_6 (.BL(BL6),.BLN(BLN6),.WL(WL245));
sram_cell_6t_5 inst_cell_245_7 (.BL(BL7),.BLN(BLN7),.WL(WL245));
sram_cell_6t_5 inst_cell_245_8 (.BL(BL8),.BLN(BLN8),.WL(WL245));
sram_cell_6t_5 inst_cell_245_9 (.BL(BL9),.BLN(BLN9),.WL(WL245));
sram_cell_6t_5 inst_cell_245_10 (.BL(BL10),.BLN(BLN10),.WL(WL245));
sram_cell_6t_5 inst_cell_245_11 (.BL(BL11),.BLN(BLN11),.WL(WL245));
sram_cell_6t_5 inst_cell_245_12 (.BL(BL12),.BLN(BLN12),.WL(WL245));
sram_cell_6t_5 inst_cell_245_13 (.BL(BL13),.BLN(BLN13),.WL(WL245));
sram_cell_6t_5 inst_cell_245_14 (.BL(BL14),.BLN(BLN14),.WL(WL245));
sram_cell_6t_5 inst_cell_245_15 (.BL(BL15),.BLN(BLN15),.WL(WL245));
sram_cell_6t_5 inst_cell_245_16 (.BL(BL16),.BLN(BLN16),.WL(WL245));
sram_cell_6t_5 inst_cell_245_17 (.BL(BL17),.BLN(BLN17),.WL(WL245));
sram_cell_6t_5 inst_cell_245_18 (.BL(BL18),.BLN(BLN18),.WL(WL245));
sram_cell_6t_5 inst_cell_245_19 (.BL(BL19),.BLN(BLN19),.WL(WL245));
sram_cell_6t_5 inst_cell_245_20 (.BL(BL20),.BLN(BLN20),.WL(WL245));
sram_cell_6t_5 inst_cell_245_21 (.BL(BL21),.BLN(BLN21),.WL(WL245));
sram_cell_6t_5 inst_cell_245_22 (.BL(BL22),.BLN(BLN22),.WL(WL245));
sram_cell_6t_5 inst_cell_245_23 (.BL(BL23),.BLN(BLN23),.WL(WL245));
sram_cell_6t_5 inst_cell_245_24 (.BL(BL24),.BLN(BLN24),.WL(WL245));
sram_cell_6t_5 inst_cell_245_25 (.BL(BL25),.BLN(BLN25),.WL(WL245));
sram_cell_6t_5 inst_cell_245_26 (.BL(BL26),.BLN(BLN26),.WL(WL245));
sram_cell_6t_5 inst_cell_245_27 (.BL(BL27),.BLN(BLN27),.WL(WL245));
sram_cell_6t_5 inst_cell_245_28 (.BL(BL28),.BLN(BLN28),.WL(WL245));
sram_cell_6t_5 inst_cell_245_29 (.BL(BL29),.BLN(BLN29),.WL(WL245));
sram_cell_6t_5 inst_cell_245_30 (.BL(BL30),.BLN(BLN30),.WL(WL245));
sram_cell_6t_5 inst_cell_245_31 (.BL(BL31),.BLN(BLN31),.WL(WL245));
sram_cell_6t_5 inst_cell_245_32 (.BL(BL32),.BLN(BLN32),.WL(WL245));
sram_cell_6t_5 inst_cell_245_33 (.BL(BL33),.BLN(BLN33),.WL(WL245));
sram_cell_6t_5 inst_cell_245_34 (.BL(BL34),.BLN(BLN34),.WL(WL245));
sram_cell_6t_5 inst_cell_245_35 (.BL(BL35),.BLN(BLN35),.WL(WL245));
sram_cell_6t_5 inst_cell_245_36 (.BL(BL36),.BLN(BLN36),.WL(WL245));
sram_cell_6t_5 inst_cell_245_37 (.BL(BL37),.BLN(BLN37),.WL(WL245));
sram_cell_6t_5 inst_cell_245_38 (.BL(BL38),.BLN(BLN38),.WL(WL245));
sram_cell_6t_5 inst_cell_245_39 (.BL(BL39),.BLN(BLN39),.WL(WL245));
sram_cell_6t_5 inst_cell_245_40 (.BL(BL40),.BLN(BLN40),.WL(WL245));
sram_cell_6t_5 inst_cell_245_41 (.BL(BL41),.BLN(BLN41),.WL(WL245));
sram_cell_6t_5 inst_cell_245_42 (.BL(BL42),.BLN(BLN42),.WL(WL245));
sram_cell_6t_5 inst_cell_245_43 (.BL(BL43),.BLN(BLN43),.WL(WL245));
sram_cell_6t_5 inst_cell_245_44 (.BL(BL44),.BLN(BLN44),.WL(WL245));
sram_cell_6t_5 inst_cell_245_45 (.BL(BL45),.BLN(BLN45),.WL(WL245));
sram_cell_6t_5 inst_cell_245_46 (.BL(BL46),.BLN(BLN46),.WL(WL245));
sram_cell_6t_5 inst_cell_245_47 (.BL(BL47),.BLN(BLN47),.WL(WL245));
sram_cell_6t_5 inst_cell_245_48 (.BL(BL48),.BLN(BLN48),.WL(WL245));
sram_cell_6t_5 inst_cell_245_49 (.BL(BL49),.BLN(BLN49),.WL(WL245));
sram_cell_6t_5 inst_cell_245_50 (.BL(BL50),.BLN(BLN50),.WL(WL245));
sram_cell_6t_5 inst_cell_245_51 (.BL(BL51),.BLN(BLN51),.WL(WL245));
sram_cell_6t_5 inst_cell_245_52 (.BL(BL52),.BLN(BLN52),.WL(WL245));
sram_cell_6t_5 inst_cell_245_53 (.BL(BL53),.BLN(BLN53),.WL(WL245));
sram_cell_6t_5 inst_cell_245_54 (.BL(BL54),.BLN(BLN54),.WL(WL245));
sram_cell_6t_5 inst_cell_245_55 (.BL(BL55),.BLN(BLN55),.WL(WL245));
sram_cell_6t_5 inst_cell_245_56 (.BL(BL56),.BLN(BLN56),.WL(WL245));
sram_cell_6t_5 inst_cell_245_57 (.BL(BL57),.BLN(BLN57),.WL(WL245));
sram_cell_6t_5 inst_cell_245_58 (.BL(BL58),.BLN(BLN58),.WL(WL245));
sram_cell_6t_5 inst_cell_245_59 (.BL(BL59),.BLN(BLN59),.WL(WL245));
sram_cell_6t_5 inst_cell_245_60 (.BL(BL60),.BLN(BLN60),.WL(WL245));
sram_cell_6t_5 inst_cell_245_61 (.BL(BL61),.BLN(BLN61),.WL(WL245));
sram_cell_6t_5 inst_cell_245_62 (.BL(BL62),.BLN(BLN62),.WL(WL245));
sram_cell_6t_5 inst_cell_245_63 (.BL(BL63),.BLN(BLN63),.WL(WL245));
sram_cell_6t_5 inst_cell_245_64 (.BL(BL64),.BLN(BLN64),.WL(WL245));
sram_cell_6t_5 inst_cell_245_65 (.BL(BL65),.BLN(BLN65),.WL(WL245));
sram_cell_6t_5 inst_cell_245_66 (.BL(BL66),.BLN(BLN66),.WL(WL245));
sram_cell_6t_5 inst_cell_245_67 (.BL(BL67),.BLN(BLN67),.WL(WL245));
sram_cell_6t_5 inst_cell_245_68 (.BL(BL68),.BLN(BLN68),.WL(WL245));
sram_cell_6t_5 inst_cell_245_69 (.BL(BL69),.BLN(BLN69),.WL(WL245));
sram_cell_6t_5 inst_cell_245_70 (.BL(BL70),.BLN(BLN70),.WL(WL245));
sram_cell_6t_5 inst_cell_245_71 (.BL(BL71),.BLN(BLN71),.WL(WL245));
sram_cell_6t_5 inst_cell_245_72 (.BL(BL72),.BLN(BLN72),.WL(WL245));
sram_cell_6t_5 inst_cell_245_73 (.BL(BL73),.BLN(BLN73),.WL(WL245));
sram_cell_6t_5 inst_cell_245_74 (.BL(BL74),.BLN(BLN74),.WL(WL245));
sram_cell_6t_5 inst_cell_245_75 (.BL(BL75),.BLN(BLN75),.WL(WL245));
sram_cell_6t_5 inst_cell_245_76 (.BL(BL76),.BLN(BLN76),.WL(WL245));
sram_cell_6t_5 inst_cell_245_77 (.BL(BL77),.BLN(BLN77),.WL(WL245));
sram_cell_6t_5 inst_cell_245_78 (.BL(BL78),.BLN(BLN78),.WL(WL245));
sram_cell_6t_5 inst_cell_245_79 (.BL(BL79),.BLN(BLN79),.WL(WL245));
sram_cell_6t_5 inst_cell_245_80 (.BL(BL80),.BLN(BLN80),.WL(WL245));
sram_cell_6t_5 inst_cell_245_81 (.BL(BL81),.BLN(BLN81),.WL(WL245));
sram_cell_6t_5 inst_cell_245_82 (.BL(BL82),.BLN(BLN82),.WL(WL245));
sram_cell_6t_5 inst_cell_245_83 (.BL(BL83),.BLN(BLN83),.WL(WL245));
sram_cell_6t_5 inst_cell_245_84 (.BL(BL84),.BLN(BLN84),.WL(WL245));
sram_cell_6t_5 inst_cell_245_85 (.BL(BL85),.BLN(BLN85),.WL(WL245));
sram_cell_6t_5 inst_cell_245_86 (.BL(BL86),.BLN(BLN86),.WL(WL245));
sram_cell_6t_5 inst_cell_245_87 (.BL(BL87),.BLN(BLN87),.WL(WL245));
sram_cell_6t_5 inst_cell_245_88 (.BL(BL88),.BLN(BLN88),.WL(WL245));
sram_cell_6t_5 inst_cell_245_89 (.BL(BL89),.BLN(BLN89),.WL(WL245));
sram_cell_6t_5 inst_cell_245_90 (.BL(BL90),.BLN(BLN90),.WL(WL245));
sram_cell_6t_5 inst_cell_245_91 (.BL(BL91),.BLN(BLN91),.WL(WL245));
sram_cell_6t_5 inst_cell_245_92 (.BL(BL92),.BLN(BLN92),.WL(WL245));
sram_cell_6t_5 inst_cell_245_93 (.BL(BL93),.BLN(BLN93),.WL(WL245));
sram_cell_6t_5 inst_cell_245_94 (.BL(BL94),.BLN(BLN94),.WL(WL245));
sram_cell_6t_5 inst_cell_245_95 (.BL(BL95),.BLN(BLN95),.WL(WL245));
sram_cell_6t_5 inst_cell_245_96 (.BL(BL96),.BLN(BLN96),.WL(WL245));
sram_cell_6t_5 inst_cell_245_97 (.BL(BL97),.BLN(BLN97),.WL(WL245));
sram_cell_6t_5 inst_cell_245_98 (.BL(BL98),.BLN(BLN98),.WL(WL245));
sram_cell_6t_5 inst_cell_245_99 (.BL(BL99),.BLN(BLN99),.WL(WL245));
sram_cell_6t_5 inst_cell_245_100 (.BL(BL100),.BLN(BLN100),.WL(WL245));
sram_cell_6t_5 inst_cell_245_101 (.BL(BL101),.BLN(BLN101),.WL(WL245));
sram_cell_6t_5 inst_cell_245_102 (.BL(BL102),.BLN(BLN102),.WL(WL245));
sram_cell_6t_5 inst_cell_245_103 (.BL(BL103),.BLN(BLN103),.WL(WL245));
sram_cell_6t_5 inst_cell_245_104 (.BL(BL104),.BLN(BLN104),.WL(WL245));
sram_cell_6t_5 inst_cell_245_105 (.BL(BL105),.BLN(BLN105),.WL(WL245));
sram_cell_6t_5 inst_cell_245_106 (.BL(BL106),.BLN(BLN106),.WL(WL245));
sram_cell_6t_5 inst_cell_245_107 (.BL(BL107),.BLN(BLN107),.WL(WL245));
sram_cell_6t_5 inst_cell_245_108 (.BL(BL108),.BLN(BLN108),.WL(WL245));
sram_cell_6t_5 inst_cell_245_109 (.BL(BL109),.BLN(BLN109),.WL(WL245));
sram_cell_6t_5 inst_cell_245_110 (.BL(BL110),.BLN(BLN110),.WL(WL245));
sram_cell_6t_5 inst_cell_245_111 (.BL(BL111),.BLN(BLN111),.WL(WL245));
sram_cell_6t_5 inst_cell_245_112 (.BL(BL112),.BLN(BLN112),.WL(WL245));
sram_cell_6t_5 inst_cell_245_113 (.BL(BL113),.BLN(BLN113),.WL(WL245));
sram_cell_6t_5 inst_cell_245_114 (.BL(BL114),.BLN(BLN114),.WL(WL245));
sram_cell_6t_5 inst_cell_245_115 (.BL(BL115),.BLN(BLN115),.WL(WL245));
sram_cell_6t_5 inst_cell_245_116 (.BL(BL116),.BLN(BLN116),.WL(WL245));
sram_cell_6t_5 inst_cell_245_117 (.BL(BL117),.BLN(BLN117),.WL(WL245));
sram_cell_6t_5 inst_cell_245_118 (.BL(BL118),.BLN(BLN118),.WL(WL245));
sram_cell_6t_5 inst_cell_245_119 (.BL(BL119),.BLN(BLN119),.WL(WL245));
sram_cell_6t_5 inst_cell_245_120 (.BL(BL120),.BLN(BLN120),.WL(WL245));
sram_cell_6t_5 inst_cell_245_121 (.BL(BL121),.BLN(BLN121),.WL(WL245));
sram_cell_6t_5 inst_cell_245_122 (.BL(BL122),.BLN(BLN122),.WL(WL245));
sram_cell_6t_5 inst_cell_245_123 (.BL(BL123),.BLN(BLN123),.WL(WL245));
sram_cell_6t_5 inst_cell_245_124 (.BL(BL124),.BLN(BLN124),.WL(WL245));
sram_cell_6t_5 inst_cell_245_125 (.BL(BL125),.BLN(BLN125),.WL(WL245));
sram_cell_6t_5 inst_cell_245_126 (.BL(BL126),.BLN(BLN126),.WL(WL245));
sram_cell_6t_5 inst_cell_245_127 (.BL(BL127),.BLN(BLN127),.WL(WL245));
sram_cell_6t_5 inst_cell_246_0 (.BL(BL0),.BLN(BLN0),.WL(WL246));
sram_cell_6t_5 inst_cell_246_1 (.BL(BL1),.BLN(BLN1),.WL(WL246));
sram_cell_6t_5 inst_cell_246_2 (.BL(BL2),.BLN(BLN2),.WL(WL246));
sram_cell_6t_5 inst_cell_246_3 (.BL(BL3),.BLN(BLN3),.WL(WL246));
sram_cell_6t_5 inst_cell_246_4 (.BL(BL4),.BLN(BLN4),.WL(WL246));
sram_cell_6t_5 inst_cell_246_5 (.BL(BL5),.BLN(BLN5),.WL(WL246));
sram_cell_6t_5 inst_cell_246_6 (.BL(BL6),.BLN(BLN6),.WL(WL246));
sram_cell_6t_5 inst_cell_246_7 (.BL(BL7),.BLN(BLN7),.WL(WL246));
sram_cell_6t_5 inst_cell_246_8 (.BL(BL8),.BLN(BLN8),.WL(WL246));
sram_cell_6t_5 inst_cell_246_9 (.BL(BL9),.BLN(BLN9),.WL(WL246));
sram_cell_6t_5 inst_cell_246_10 (.BL(BL10),.BLN(BLN10),.WL(WL246));
sram_cell_6t_5 inst_cell_246_11 (.BL(BL11),.BLN(BLN11),.WL(WL246));
sram_cell_6t_5 inst_cell_246_12 (.BL(BL12),.BLN(BLN12),.WL(WL246));
sram_cell_6t_5 inst_cell_246_13 (.BL(BL13),.BLN(BLN13),.WL(WL246));
sram_cell_6t_5 inst_cell_246_14 (.BL(BL14),.BLN(BLN14),.WL(WL246));
sram_cell_6t_5 inst_cell_246_15 (.BL(BL15),.BLN(BLN15),.WL(WL246));
sram_cell_6t_5 inst_cell_246_16 (.BL(BL16),.BLN(BLN16),.WL(WL246));
sram_cell_6t_5 inst_cell_246_17 (.BL(BL17),.BLN(BLN17),.WL(WL246));
sram_cell_6t_5 inst_cell_246_18 (.BL(BL18),.BLN(BLN18),.WL(WL246));
sram_cell_6t_5 inst_cell_246_19 (.BL(BL19),.BLN(BLN19),.WL(WL246));
sram_cell_6t_5 inst_cell_246_20 (.BL(BL20),.BLN(BLN20),.WL(WL246));
sram_cell_6t_5 inst_cell_246_21 (.BL(BL21),.BLN(BLN21),.WL(WL246));
sram_cell_6t_5 inst_cell_246_22 (.BL(BL22),.BLN(BLN22),.WL(WL246));
sram_cell_6t_5 inst_cell_246_23 (.BL(BL23),.BLN(BLN23),.WL(WL246));
sram_cell_6t_5 inst_cell_246_24 (.BL(BL24),.BLN(BLN24),.WL(WL246));
sram_cell_6t_5 inst_cell_246_25 (.BL(BL25),.BLN(BLN25),.WL(WL246));
sram_cell_6t_5 inst_cell_246_26 (.BL(BL26),.BLN(BLN26),.WL(WL246));
sram_cell_6t_5 inst_cell_246_27 (.BL(BL27),.BLN(BLN27),.WL(WL246));
sram_cell_6t_5 inst_cell_246_28 (.BL(BL28),.BLN(BLN28),.WL(WL246));
sram_cell_6t_5 inst_cell_246_29 (.BL(BL29),.BLN(BLN29),.WL(WL246));
sram_cell_6t_5 inst_cell_246_30 (.BL(BL30),.BLN(BLN30),.WL(WL246));
sram_cell_6t_5 inst_cell_246_31 (.BL(BL31),.BLN(BLN31),.WL(WL246));
sram_cell_6t_5 inst_cell_246_32 (.BL(BL32),.BLN(BLN32),.WL(WL246));
sram_cell_6t_5 inst_cell_246_33 (.BL(BL33),.BLN(BLN33),.WL(WL246));
sram_cell_6t_5 inst_cell_246_34 (.BL(BL34),.BLN(BLN34),.WL(WL246));
sram_cell_6t_5 inst_cell_246_35 (.BL(BL35),.BLN(BLN35),.WL(WL246));
sram_cell_6t_5 inst_cell_246_36 (.BL(BL36),.BLN(BLN36),.WL(WL246));
sram_cell_6t_5 inst_cell_246_37 (.BL(BL37),.BLN(BLN37),.WL(WL246));
sram_cell_6t_5 inst_cell_246_38 (.BL(BL38),.BLN(BLN38),.WL(WL246));
sram_cell_6t_5 inst_cell_246_39 (.BL(BL39),.BLN(BLN39),.WL(WL246));
sram_cell_6t_5 inst_cell_246_40 (.BL(BL40),.BLN(BLN40),.WL(WL246));
sram_cell_6t_5 inst_cell_246_41 (.BL(BL41),.BLN(BLN41),.WL(WL246));
sram_cell_6t_5 inst_cell_246_42 (.BL(BL42),.BLN(BLN42),.WL(WL246));
sram_cell_6t_5 inst_cell_246_43 (.BL(BL43),.BLN(BLN43),.WL(WL246));
sram_cell_6t_5 inst_cell_246_44 (.BL(BL44),.BLN(BLN44),.WL(WL246));
sram_cell_6t_5 inst_cell_246_45 (.BL(BL45),.BLN(BLN45),.WL(WL246));
sram_cell_6t_5 inst_cell_246_46 (.BL(BL46),.BLN(BLN46),.WL(WL246));
sram_cell_6t_5 inst_cell_246_47 (.BL(BL47),.BLN(BLN47),.WL(WL246));
sram_cell_6t_5 inst_cell_246_48 (.BL(BL48),.BLN(BLN48),.WL(WL246));
sram_cell_6t_5 inst_cell_246_49 (.BL(BL49),.BLN(BLN49),.WL(WL246));
sram_cell_6t_5 inst_cell_246_50 (.BL(BL50),.BLN(BLN50),.WL(WL246));
sram_cell_6t_5 inst_cell_246_51 (.BL(BL51),.BLN(BLN51),.WL(WL246));
sram_cell_6t_5 inst_cell_246_52 (.BL(BL52),.BLN(BLN52),.WL(WL246));
sram_cell_6t_5 inst_cell_246_53 (.BL(BL53),.BLN(BLN53),.WL(WL246));
sram_cell_6t_5 inst_cell_246_54 (.BL(BL54),.BLN(BLN54),.WL(WL246));
sram_cell_6t_5 inst_cell_246_55 (.BL(BL55),.BLN(BLN55),.WL(WL246));
sram_cell_6t_5 inst_cell_246_56 (.BL(BL56),.BLN(BLN56),.WL(WL246));
sram_cell_6t_5 inst_cell_246_57 (.BL(BL57),.BLN(BLN57),.WL(WL246));
sram_cell_6t_5 inst_cell_246_58 (.BL(BL58),.BLN(BLN58),.WL(WL246));
sram_cell_6t_5 inst_cell_246_59 (.BL(BL59),.BLN(BLN59),.WL(WL246));
sram_cell_6t_5 inst_cell_246_60 (.BL(BL60),.BLN(BLN60),.WL(WL246));
sram_cell_6t_5 inst_cell_246_61 (.BL(BL61),.BLN(BLN61),.WL(WL246));
sram_cell_6t_5 inst_cell_246_62 (.BL(BL62),.BLN(BLN62),.WL(WL246));
sram_cell_6t_5 inst_cell_246_63 (.BL(BL63),.BLN(BLN63),.WL(WL246));
sram_cell_6t_5 inst_cell_246_64 (.BL(BL64),.BLN(BLN64),.WL(WL246));
sram_cell_6t_5 inst_cell_246_65 (.BL(BL65),.BLN(BLN65),.WL(WL246));
sram_cell_6t_5 inst_cell_246_66 (.BL(BL66),.BLN(BLN66),.WL(WL246));
sram_cell_6t_5 inst_cell_246_67 (.BL(BL67),.BLN(BLN67),.WL(WL246));
sram_cell_6t_5 inst_cell_246_68 (.BL(BL68),.BLN(BLN68),.WL(WL246));
sram_cell_6t_5 inst_cell_246_69 (.BL(BL69),.BLN(BLN69),.WL(WL246));
sram_cell_6t_5 inst_cell_246_70 (.BL(BL70),.BLN(BLN70),.WL(WL246));
sram_cell_6t_5 inst_cell_246_71 (.BL(BL71),.BLN(BLN71),.WL(WL246));
sram_cell_6t_5 inst_cell_246_72 (.BL(BL72),.BLN(BLN72),.WL(WL246));
sram_cell_6t_5 inst_cell_246_73 (.BL(BL73),.BLN(BLN73),.WL(WL246));
sram_cell_6t_5 inst_cell_246_74 (.BL(BL74),.BLN(BLN74),.WL(WL246));
sram_cell_6t_5 inst_cell_246_75 (.BL(BL75),.BLN(BLN75),.WL(WL246));
sram_cell_6t_5 inst_cell_246_76 (.BL(BL76),.BLN(BLN76),.WL(WL246));
sram_cell_6t_5 inst_cell_246_77 (.BL(BL77),.BLN(BLN77),.WL(WL246));
sram_cell_6t_5 inst_cell_246_78 (.BL(BL78),.BLN(BLN78),.WL(WL246));
sram_cell_6t_5 inst_cell_246_79 (.BL(BL79),.BLN(BLN79),.WL(WL246));
sram_cell_6t_5 inst_cell_246_80 (.BL(BL80),.BLN(BLN80),.WL(WL246));
sram_cell_6t_5 inst_cell_246_81 (.BL(BL81),.BLN(BLN81),.WL(WL246));
sram_cell_6t_5 inst_cell_246_82 (.BL(BL82),.BLN(BLN82),.WL(WL246));
sram_cell_6t_5 inst_cell_246_83 (.BL(BL83),.BLN(BLN83),.WL(WL246));
sram_cell_6t_5 inst_cell_246_84 (.BL(BL84),.BLN(BLN84),.WL(WL246));
sram_cell_6t_5 inst_cell_246_85 (.BL(BL85),.BLN(BLN85),.WL(WL246));
sram_cell_6t_5 inst_cell_246_86 (.BL(BL86),.BLN(BLN86),.WL(WL246));
sram_cell_6t_5 inst_cell_246_87 (.BL(BL87),.BLN(BLN87),.WL(WL246));
sram_cell_6t_5 inst_cell_246_88 (.BL(BL88),.BLN(BLN88),.WL(WL246));
sram_cell_6t_5 inst_cell_246_89 (.BL(BL89),.BLN(BLN89),.WL(WL246));
sram_cell_6t_5 inst_cell_246_90 (.BL(BL90),.BLN(BLN90),.WL(WL246));
sram_cell_6t_5 inst_cell_246_91 (.BL(BL91),.BLN(BLN91),.WL(WL246));
sram_cell_6t_5 inst_cell_246_92 (.BL(BL92),.BLN(BLN92),.WL(WL246));
sram_cell_6t_5 inst_cell_246_93 (.BL(BL93),.BLN(BLN93),.WL(WL246));
sram_cell_6t_5 inst_cell_246_94 (.BL(BL94),.BLN(BLN94),.WL(WL246));
sram_cell_6t_5 inst_cell_246_95 (.BL(BL95),.BLN(BLN95),.WL(WL246));
sram_cell_6t_5 inst_cell_246_96 (.BL(BL96),.BLN(BLN96),.WL(WL246));
sram_cell_6t_5 inst_cell_246_97 (.BL(BL97),.BLN(BLN97),.WL(WL246));
sram_cell_6t_5 inst_cell_246_98 (.BL(BL98),.BLN(BLN98),.WL(WL246));
sram_cell_6t_5 inst_cell_246_99 (.BL(BL99),.BLN(BLN99),.WL(WL246));
sram_cell_6t_5 inst_cell_246_100 (.BL(BL100),.BLN(BLN100),.WL(WL246));
sram_cell_6t_5 inst_cell_246_101 (.BL(BL101),.BLN(BLN101),.WL(WL246));
sram_cell_6t_5 inst_cell_246_102 (.BL(BL102),.BLN(BLN102),.WL(WL246));
sram_cell_6t_5 inst_cell_246_103 (.BL(BL103),.BLN(BLN103),.WL(WL246));
sram_cell_6t_5 inst_cell_246_104 (.BL(BL104),.BLN(BLN104),.WL(WL246));
sram_cell_6t_5 inst_cell_246_105 (.BL(BL105),.BLN(BLN105),.WL(WL246));
sram_cell_6t_5 inst_cell_246_106 (.BL(BL106),.BLN(BLN106),.WL(WL246));
sram_cell_6t_5 inst_cell_246_107 (.BL(BL107),.BLN(BLN107),.WL(WL246));
sram_cell_6t_5 inst_cell_246_108 (.BL(BL108),.BLN(BLN108),.WL(WL246));
sram_cell_6t_5 inst_cell_246_109 (.BL(BL109),.BLN(BLN109),.WL(WL246));
sram_cell_6t_5 inst_cell_246_110 (.BL(BL110),.BLN(BLN110),.WL(WL246));
sram_cell_6t_5 inst_cell_246_111 (.BL(BL111),.BLN(BLN111),.WL(WL246));
sram_cell_6t_5 inst_cell_246_112 (.BL(BL112),.BLN(BLN112),.WL(WL246));
sram_cell_6t_5 inst_cell_246_113 (.BL(BL113),.BLN(BLN113),.WL(WL246));
sram_cell_6t_5 inst_cell_246_114 (.BL(BL114),.BLN(BLN114),.WL(WL246));
sram_cell_6t_5 inst_cell_246_115 (.BL(BL115),.BLN(BLN115),.WL(WL246));
sram_cell_6t_5 inst_cell_246_116 (.BL(BL116),.BLN(BLN116),.WL(WL246));
sram_cell_6t_5 inst_cell_246_117 (.BL(BL117),.BLN(BLN117),.WL(WL246));
sram_cell_6t_5 inst_cell_246_118 (.BL(BL118),.BLN(BLN118),.WL(WL246));
sram_cell_6t_5 inst_cell_246_119 (.BL(BL119),.BLN(BLN119),.WL(WL246));
sram_cell_6t_5 inst_cell_246_120 (.BL(BL120),.BLN(BLN120),.WL(WL246));
sram_cell_6t_5 inst_cell_246_121 (.BL(BL121),.BLN(BLN121),.WL(WL246));
sram_cell_6t_5 inst_cell_246_122 (.BL(BL122),.BLN(BLN122),.WL(WL246));
sram_cell_6t_5 inst_cell_246_123 (.BL(BL123),.BLN(BLN123),.WL(WL246));
sram_cell_6t_5 inst_cell_246_124 (.BL(BL124),.BLN(BLN124),.WL(WL246));
sram_cell_6t_5 inst_cell_246_125 (.BL(BL125),.BLN(BLN125),.WL(WL246));
sram_cell_6t_5 inst_cell_246_126 (.BL(BL126),.BLN(BLN126),.WL(WL246));
sram_cell_6t_5 inst_cell_246_127 (.BL(BL127),.BLN(BLN127),.WL(WL246));
sram_cell_6t_5 inst_cell_247_0 (.BL(BL0),.BLN(BLN0),.WL(WL247));
sram_cell_6t_5 inst_cell_247_1 (.BL(BL1),.BLN(BLN1),.WL(WL247));
sram_cell_6t_5 inst_cell_247_2 (.BL(BL2),.BLN(BLN2),.WL(WL247));
sram_cell_6t_5 inst_cell_247_3 (.BL(BL3),.BLN(BLN3),.WL(WL247));
sram_cell_6t_5 inst_cell_247_4 (.BL(BL4),.BLN(BLN4),.WL(WL247));
sram_cell_6t_5 inst_cell_247_5 (.BL(BL5),.BLN(BLN5),.WL(WL247));
sram_cell_6t_5 inst_cell_247_6 (.BL(BL6),.BLN(BLN6),.WL(WL247));
sram_cell_6t_5 inst_cell_247_7 (.BL(BL7),.BLN(BLN7),.WL(WL247));
sram_cell_6t_5 inst_cell_247_8 (.BL(BL8),.BLN(BLN8),.WL(WL247));
sram_cell_6t_5 inst_cell_247_9 (.BL(BL9),.BLN(BLN9),.WL(WL247));
sram_cell_6t_5 inst_cell_247_10 (.BL(BL10),.BLN(BLN10),.WL(WL247));
sram_cell_6t_5 inst_cell_247_11 (.BL(BL11),.BLN(BLN11),.WL(WL247));
sram_cell_6t_5 inst_cell_247_12 (.BL(BL12),.BLN(BLN12),.WL(WL247));
sram_cell_6t_5 inst_cell_247_13 (.BL(BL13),.BLN(BLN13),.WL(WL247));
sram_cell_6t_5 inst_cell_247_14 (.BL(BL14),.BLN(BLN14),.WL(WL247));
sram_cell_6t_5 inst_cell_247_15 (.BL(BL15),.BLN(BLN15),.WL(WL247));
sram_cell_6t_5 inst_cell_247_16 (.BL(BL16),.BLN(BLN16),.WL(WL247));
sram_cell_6t_5 inst_cell_247_17 (.BL(BL17),.BLN(BLN17),.WL(WL247));
sram_cell_6t_5 inst_cell_247_18 (.BL(BL18),.BLN(BLN18),.WL(WL247));
sram_cell_6t_5 inst_cell_247_19 (.BL(BL19),.BLN(BLN19),.WL(WL247));
sram_cell_6t_5 inst_cell_247_20 (.BL(BL20),.BLN(BLN20),.WL(WL247));
sram_cell_6t_5 inst_cell_247_21 (.BL(BL21),.BLN(BLN21),.WL(WL247));
sram_cell_6t_5 inst_cell_247_22 (.BL(BL22),.BLN(BLN22),.WL(WL247));
sram_cell_6t_5 inst_cell_247_23 (.BL(BL23),.BLN(BLN23),.WL(WL247));
sram_cell_6t_5 inst_cell_247_24 (.BL(BL24),.BLN(BLN24),.WL(WL247));
sram_cell_6t_5 inst_cell_247_25 (.BL(BL25),.BLN(BLN25),.WL(WL247));
sram_cell_6t_5 inst_cell_247_26 (.BL(BL26),.BLN(BLN26),.WL(WL247));
sram_cell_6t_5 inst_cell_247_27 (.BL(BL27),.BLN(BLN27),.WL(WL247));
sram_cell_6t_5 inst_cell_247_28 (.BL(BL28),.BLN(BLN28),.WL(WL247));
sram_cell_6t_5 inst_cell_247_29 (.BL(BL29),.BLN(BLN29),.WL(WL247));
sram_cell_6t_5 inst_cell_247_30 (.BL(BL30),.BLN(BLN30),.WL(WL247));
sram_cell_6t_5 inst_cell_247_31 (.BL(BL31),.BLN(BLN31),.WL(WL247));
sram_cell_6t_5 inst_cell_247_32 (.BL(BL32),.BLN(BLN32),.WL(WL247));
sram_cell_6t_5 inst_cell_247_33 (.BL(BL33),.BLN(BLN33),.WL(WL247));
sram_cell_6t_5 inst_cell_247_34 (.BL(BL34),.BLN(BLN34),.WL(WL247));
sram_cell_6t_5 inst_cell_247_35 (.BL(BL35),.BLN(BLN35),.WL(WL247));
sram_cell_6t_5 inst_cell_247_36 (.BL(BL36),.BLN(BLN36),.WL(WL247));
sram_cell_6t_5 inst_cell_247_37 (.BL(BL37),.BLN(BLN37),.WL(WL247));
sram_cell_6t_5 inst_cell_247_38 (.BL(BL38),.BLN(BLN38),.WL(WL247));
sram_cell_6t_5 inst_cell_247_39 (.BL(BL39),.BLN(BLN39),.WL(WL247));
sram_cell_6t_5 inst_cell_247_40 (.BL(BL40),.BLN(BLN40),.WL(WL247));
sram_cell_6t_5 inst_cell_247_41 (.BL(BL41),.BLN(BLN41),.WL(WL247));
sram_cell_6t_5 inst_cell_247_42 (.BL(BL42),.BLN(BLN42),.WL(WL247));
sram_cell_6t_5 inst_cell_247_43 (.BL(BL43),.BLN(BLN43),.WL(WL247));
sram_cell_6t_5 inst_cell_247_44 (.BL(BL44),.BLN(BLN44),.WL(WL247));
sram_cell_6t_5 inst_cell_247_45 (.BL(BL45),.BLN(BLN45),.WL(WL247));
sram_cell_6t_5 inst_cell_247_46 (.BL(BL46),.BLN(BLN46),.WL(WL247));
sram_cell_6t_5 inst_cell_247_47 (.BL(BL47),.BLN(BLN47),.WL(WL247));
sram_cell_6t_5 inst_cell_247_48 (.BL(BL48),.BLN(BLN48),.WL(WL247));
sram_cell_6t_5 inst_cell_247_49 (.BL(BL49),.BLN(BLN49),.WL(WL247));
sram_cell_6t_5 inst_cell_247_50 (.BL(BL50),.BLN(BLN50),.WL(WL247));
sram_cell_6t_5 inst_cell_247_51 (.BL(BL51),.BLN(BLN51),.WL(WL247));
sram_cell_6t_5 inst_cell_247_52 (.BL(BL52),.BLN(BLN52),.WL(WL247));
sram_cell_6t_5 inst_cell_247_53 (.BL(BL53),.BLN(BLN53),.WL(WL247));
sram_cell_6t_5 inst_cell_247_54 (.BL(BL54),.BLN(BLN54),.WL(WL247));
sram_cell_6t_5 inst_cell_247_55 (.BL(BL55),.BLN(BLN55),.WL(WL247));
sram_cell_6t_5 inst_cell_247_56 (.BL(BL56),.BLN(BLN56),.WL(WL247));
sram_cell_6t_5 inst_cell_247_57 (.BL(BL57),.BLN(BLN57),.WL(WL247));
sram_cell_6t_5 inst_cell_247_58 (.BL(BL58),.BLN(BLN58),.WL(WL247));
sram_cell_6t_5 inst_cell_247_59 (.BL(BL59),.BLN(BLN59),.WL(WL247));
sram_cell_6t_5 inst_cell_247_60 (.BL(BL60),.BLN(BLN60),.WL(WL247));
sram_cell_6t_5 inst_cell_247_61 (.BL(BL61),.BLN(BLN61),.WL(WL247));
sram_cell_6t_5 inst_cell_247_62 (.BL(BL62),.BLN(BLN62),.WL(WL247));
sram_cell_6t_5 inst_cell_247_63 (.BL(BL63),.BLN(BLN63),.WL(WL247));
sram_cell_6t_5 inst_cell_247_64 (.BL(BL64),.BLN(BLN64),.WL(WL247));
sram_cell_6t_5 inst_cell_247_65 (.BL(BL65),.BLN(BLN65),.WL(WL247));
sram_cell_6t_5 inst_cell_247_66 (.BL(BL66),.BLN(BLN66),.WL(WL247));
sram_cell_6t_5 inst_cell_247_67 (.BL(BL67),.BLN(BLN67),.WL(WL247));
sram_cell_6t_5 inst_cell_247_68 (.BL(BL68),.BLN(BLN68),.WL(WL247));
sram_cell_6t_5 inst_cell_247_69 (.BL(BL69),.BLN(BLN69),.WL(WL247));
sram_cell_6t_5 inst_cell_247_70 (.BL(BL70),.BLN(BLN70),.WL(WL247));
sram_cell_6t_5 inst_cell_247_71 (.BL(BL71),.BLN(BLN71),.WL(WL247));
sram_cell_6t_5 inst_cell_247_72 (.BL(BL72),.BLN(BLN72),.WL(WL247));
sram_cell_6t_5 inst_cell_247_73 (.BL(BL73),.BLN(BLN73),.WL(WL247));
sram_cell_6t_5 inst_cell_247_74 (.BL(BL74),.BLN(BLN74),.WL(WL247));
sram_cell_6t_5 inst_cell_247_75 (.BL(BL75),.BLN(BLN75),.WL(WL247));
sram_cell_6t_5 inst_cell_247_76 (.BL(BL76),.BLN(BLN76),.WL(WL247));
sram_cell_6t_5 inst_cell_247_77 (.BL(BL77),.BLN(BLN77),.WL(WL247));
sram_cell_6t_5 inst_cell_247_78 (.BL(BL78),.BLN(BLN78),.WL(WL247));
sram_cell_6t_5 inst_cell_247_79 (.BL(BL79),.BLN(BLN79),.WL(WL247));
sram_cell_6t_5 inst_cell_247_80 (.BL(BL80),.BLN(BLN80),.WL(WL247));
sram_cell_6t_5 inst_cell_247_81 (.BL(BL81),.BLN(BLN81),.WL(WL247));
sram_cell_6t_5 inst_cell_247_82 (.BL(BL82),.BLN(BLN82),.WL(WL247));
sram_cell_6t_5 inst_cell_247_83 (.BL(BL83),.BLN(BLN83),.WL(WL247));
sram_cell_6t_5 inst_cell_247_84 (.BL(BL84),.BLN(BLN84),.WL(WL247));
sram_cell_6t_5 inst_cell_247_85 (.BL(BL85),.BLN(BLN85),.WL(WL247));
sram_cell_6t_5 inst_cell_247_86 (.BL(BL86),.BLN(BLN86),.WL(WL247));
sram_cell_6t_5 inst_cell_247_87 (.BL(BL87),.BLN(BLN87),.WL(WL247));
sram_cell_6t_5 inst_cell_247_88 (.BL(BL88),.BLN(BLN88),.WL(WL247));
sram_cell_6t_5 inst_cell_247_89 (.BL(BL89),.BLN(BLN89),.WL(WL247));
sram_cell_6t_5 inst_cell_247_90 (.BL(BL90),.BLN(BLN90),.WL(WL247));
sram_cell_6t_5 inst_cell_247_91 (.BL(BL91),.BLN(BLN91),.WL(WL247));
sram_cell_6t_5 inst_cell_247_92 (.BL(BL92),.BLN(BLN92),.WL(WL247));
sram_cell_6t_5 inst_cell_247_93 (.BL(BL93),.BLN(BLN93),.WL(WL247));
sram_cell_6t_5 inst_cell_247_94 (.BL(BL94),.BLN(BLN94),.WL(WL247));
sram_cell_6t_5 inst_cell_247_95 (.BL(BL95),.BLN(BLN95),.WL(WL247));
sram_cell_6t_5 inst_cell_247_96 (.BL(BL96),.BLN(BLN96),.WL(WL247));
sram_cell_6t_5 inst_cell_247_97 (.BL(BL97),.BLN(BLN97),.WL(WL247));
sram_cell_6t_5 inst_cell_247_98 (.BL(BL98),.BLN(BLN98),.WL(WL247));
sram_cell_6t_5 inst_cell_247_99 (.BL(BL99),.BLN(BLN99),.WL(WL247));
sram_cell_6t_5 inst_cell_247_100 (.BL(BL100),.BLN(BLN100),.WL(WL247));
sram_cell_6t_5 inst_cell_247_101 (.BL(BL101),.BLN(BLN101),.WL(WL247));
sram_cell_6t_5 inst_cell_247_102 (.BL(BL102),.BLN(BLN102),.WL(WL247));
sram_cell_6t_5 inst_cell_247_103 (.BL(BL103),.BLN(BLN103),.WL(WL247));
sram_cell_6t_5 inst_cell_247_104 (.BL(BL104),.BLN(BLN104),.WL(WL247));
sram_cell_6t_5 inst_cell_247_105 (.BL(BL105),.BLN(BLN105),.WL(WL247));
sram_cell_6t_5 inst_cell_247_106 (.BL(BL106),.BLN(BLN106),.WL(WL247));
sram_cell_6t_5 inst_cell_247_107 (.BL(BL107),.BLN(BLN107),.WL(WL247));
sram_cell_6t_5 inst_cell_247_108 (.BL(BL108),.BLN(BLN108),.WL(WL247));
sram_cell_6t_5 inst_cell_247_109 (.BL(BL109),.BLN(BLN109),.WL(WL247));
sram_cell_6t_5 inst_cell_247_110 (.BL(BL110),.BLN(BLN110),.WL(WL247));
sram_cell_6t_5 inst_cell_247_111 (.BL(BL111),.BLN(BLN111),.WL(WL247));
sram_cell_6t_5 inst_cell_247_112 (.BL(BL112),.BLN(BLN112),.WL(WL247));
sram_cell_6t_5 inst_cell_247_113 (.BL(BL113),.BLN(BLN113),.WL(WL247));
sram_cell_6t_5 inst_cell_247_114 (.BL(BL114),.BLN(BLN114),.WL(WL247));
sram_cell_6t_5 inst_cell_247_115 (.BL(BL115),.BLN(BLN115),.WL(WL247));
sram_cell_6t_5 inst_cell_247_116 (.BL(BL116),.BLN(BLN116),.WL(WL247));
sram_cell_6t_5 inst_cell_247_117 (.BL(BL117),.BLN(BLN117),.WL(WL247));
sram_cell_6t_5 inst_cell_247_118 (.BL(BL118),.BLN(BLN118),.WL(WL247));
sram_cell_6t_5 inst_cell_247_119 (.BL(BL119),.BLN(BLN119),.WL(WL247));
sram_cell_6t_5 inst_cell_247_120 (.BL(BL120),.BLN(BLN120),.WL(WL247));
sram_cell_6t_5 inst_cell_247_121 (.BL(BL121),.BLN(BLN121),.WL(WL247));
sram_cell_6t_5 inst_cell_247_122 (.BL(BL122),.BLN(BLN122),.WL(WL247));
sram_cell_6t_5 inst_cell_247_123 (.BL(BL123),.BLN(BLN123),.WL(WL247));
sram_cell_6t_5 inst_cell_247_124 (.BL(BL124),.BLN(BLN124),.WL(WL247));
sram_cell_6t_5 inst_cell_247_125 (.BL(BL125),.BLN(BLN125),.WL(WL247));
sram_cell_6t_5 inst_cell_247_126 (.BL(BL126),.BLN(BLN126),.WL(WL247));
sram_cell_6t_5 inst_cell_247_127 (.BL(BL127),.BLN(BLN127),.WL(WL247));
sram_cell_6t_5 inst_cell_248_0 (.BL(BL0),.BLN(BLN0),.WL(WL248));
sram_cell_6t_5 inst_cell_248_1 (.BL(BL1),.BLN(BLN1),.WL(WL248));
sram_cell_6t_5 inst_cell_248_2 (.BL(BL2),.BLN(BLN2),.WL(WL248));
sram_cell_6t_5 inst_cell_248_3 (.BL(BL3),.BLN(BLN3),.WL(WL248));
sram_cell_6t_5 inst_cell_248_4 (.BL(BL4),.BLN(BLN4),.WL(WL248));
sram_cell_6t_5 inst_cell_248_5 (.BL(BL5),.BLN(BLN5),.WL(WL248));
sram_cell_6t_5 inst_cell_248_6 (.BL(BL6),.BLN(BLN6),.WL(WL248));
sram_cell_6t_5 inst_cell_248_7 (.BL(BL7),.BLN(BLN7),.WL(WL248));
sram_cell_6t_5 inst_cell_248_8 (.BL(BL8),.BLN(BLN8),.WL(WL248));
sram_cell_6t_5 inst_cell_248_9 (.BL(BL9),.BLN(BLN9),.WL(WL248));
sram_cell_6t_5 inst_cell_248_10 (.BL(BL10),.BLN(BLN10),.WL(WL248));
sram_cell_6t_5 inst_cell_248_11 (.BL(BL11),.BLN(BLN11),.WL(WL248));
sram_cell_6t_5 inst_cell_248_12 (.BL(BL12),.BLN(BLN12),.WL(WL248));
sram_cell_6t_5 inst_cell_248_13 (.BL(BL13),.BLN(BLN13),.WL(WL248));
sram_cell_6t_5 inst_cell_248_14 (.BL(BL14),.BLN(BLN14),.WL(WL248));
sram_cell_6t_5 inst_cell_248_15 (.BL(BL15),.BLN(BLN15),.WL(WL248));
sram_cell_6t_5 inst_cell_248_16 (.BL(BL16),.BLN(BLN16),.WL(WL248));
sram_cell_6t_5 inst_cell_248_17 (.BL(BL17),.BLN(BLN17),.WL(WL248));
sram_cell_6t_5 inst_cell_248_18 (.BL(BL18),.BLN(BLN18),.WL(WL248));
sram_cell_6t_5 inst_cell_248_19 (.BL(BL19),.BLN(BLN19),.WL(WL248));
sram_cell_6t_5 inst_cell_248_20 (.BL(BL20),.BLN(BLN20),.WL(WL248));
sram_cell_6t_5 inst_cell_248_21 (.BL(BL21),.BLN(BLN21),.WL(WL248));
sram_cell_6t_5 inst_cell_248_22 (.BL(BL22),.BLN(BLN22),.WL(WL248));
sram_cell_6t_5 inst_cell_248_23 (.BL(BL23),.BLN(BLN23),.WL(WL248));
sram_cell_6t_5 inst_cell_248_24 (.BL(BL24),.BLN(BLN24),.WL(WL248));
sram_cell_6t_5 inst_cell_248_25 (.BL(BL25),.BLN(BLN25),.WL(WL248));
sram_cell_6t_5 inst_cell_248_26 (.BL(BL26),.BLN(BLN26),.WL(WL248));
sram_cell_6t_5 inst_cell_248_27 (.BL(BL27),.BLN(BLN27),.WL(WL248));
sram_cell_6t_5 inst_cell_248_28 (.BL(BL28),.BLN(BLN28),.WL(WL248));
sram_cell_6t_5 inst_cell_248_29 (.BL(BL29),.BLN(BLN29),.WL(WL248));
sram_cell_6t_5 inst_cell_248_30 (.BL(BL30),.BLN(BLN30),.WL(WL248));
sram_cell_6t_5 inst_cell_248_31 (.BL(BL31),.BLN(BLN31),.WL(WL248));
sram_cell_6t_5 inst_cell_248_32 (.BL(BL32),.BLN(BLN32),.WL(WL248));
sram_cell_6t_5 inst_cell_248_33 (.BL(BL33),.BLN(BLN33),.WL(WL248));
sram_cell_6t_5 inst_cell_248_34 (.BL(BL34),.BLN(BLN34),.WL(WL248));
sram_cell_6t_5 inst_cell_248_35 (.BL(BL35),.BLN(BLN35),.WL(WL248));
sram_cell_6t_5 inst_cell_248_36 (.BL(BL36),.BLN(BLN36),.WL(WL248));
sram_cell_6t_5 inst_cell_248_37 (.BL(BL37),.BLN(BLN37),.WL(WL248));
sram_cell_6t_5 inst_cell_248_38 (.BL(BL38),.BLN(BLN38),.WL(WL248));
sram_cell_6t_5 inst_cell_248_39 (.BL(BL39),.BLN(BLN39),.WL(WL248));
sram_cell_6t_5 inst_cell_248_40 (.BL(BL40),.BLN(BLN40),.WL(WL248));
sram_cell_6t_5 inst_cell_248_41 (.BL(BL41),.BLN(BLN41),.WL(WL248));
sram_cell_6t_5 inst_cell_248_42 (.BL(BL42),.BLN(BLN42),.WL(WL248));
sram_cell_6t_5 inst_cell_248_43 (.BL(BL43),.BLN(BLN43),.WL(WL248));
sram_cell_6t_5 inst_cell_248_44 (.BL(BL44),.BLN(BLN44),.WL(WL248));
sram_cell_6t_5 inst_cell_248_45 (.BL(BL45),.BLN(BLN45),.WL(WL248));
sram_cell_6t_5 inst_cell_248_46 (.BL(BL46),.BLN(BLN46),.WL(WL248));
sram_cell_6t_5 inst_cell_248_47 (.BL(BL47),.BLN(BLN47),.WL(WL248));
sram_cell_6t_5 inst_cell_248_48 (.BL(BL48),.BLN(BLN48),.WL(WL248));
sram_cell_6t_5 inst_cell_248_49 (.BL(BL49),.BLN(BLN49),.WL(WL248));
sram_cell_6t_5 inst_cell_248_50 (.BL(BL50),.BLN(BLN50),.WL(WL248));
sram_cell_6t_5 inst_cell_248_51 (.BL(BL51),.BLN(BLN51),.WL(WL248));
sram_cell_6t_5 inst_cell_248_52 (.BL(BL52),.BLN(BLN52),.WL(WL248));
sram_cell_6t_5 inst_cell_248_53 (.BL(BL53),.BLN(BLN53),.WL(WL248));
sram_cell_6t_5 inst_cell_248_54 (.BL(BL54),.BLN(BLN54),.WL(WL248));
sram_cell_6t_5 inst_cell_248_55 (.BL(BL55),.BLN(BLN55),.WL(WL248));
sram_cell_6t_5 inst_cell_248_56 (.BL(BL56),.BLN(BLN56),.WL(WL248));
sram_cell_6t_5 inst_cell_248_57 (.BL(BL57),.BLN(BLN57),.WL(WL248));
sram_cell_6t_5 inst_cell_248_58 (.BL(BL58),.BLN(BLN58),.WL(WL248));
sram_cell_6t_5 inst_cell_248_59 (.BL(BL59),.BLN(BLN59),.WL(WL248));
sram_cell_6t_5 inst_cell_248_60 (.BL(BL60),.BLN(BLN60),.WL(WL248));
sram_cell_6t_5 inst_cell_248_61 (.BL(BL61),.BLN(BLN61),.WL(WL248));
sram_cell_6t_5 inst_cell_248_62 (.BL(BL62),.BLN(BLN62),.WL(WL248));
sram_cell_6t_5 inst_cell_248_63 (.BL(BL63),.BLN(BLN63),.WL(WL248));
sram_cell_6t_5 inst_cell_248_64 (.BL(BL64),.BLN(BLN64),.WL(WL248));
sram_cell_6t_5 inst_cell_248_65 (.BL(BL65),.BLN(BLN65),.WL(WL248));
sram_cell_6t_5 inst_cell_248_66 (.BL(BL66),.BLN(BLN66),.WL(WL248));
sram_cell_6t_5 inst_cell_248_67 (.BL(BL67),.BLN(BLN67),.WL(WL248));
sram_cell_6t_5 inst_cell_248_68 (.BL(BL68),.BLN(BLN68),.WL(WL248));
sram_cell_6t_5 inst_cell_248_69 (.BL(BL69),.BLN(BLN69),.WL(WL248));
sram_cell_6t_5 inst_cell_248_70 (.BL(BL70),.BLN(BLN70),.WL(WL248));
sram_cell_6t_5 inst_cell_248_71 (.BL(BL71),.BLN(BLN71),.WL(WL248));
sram_cell_6t_5 inst_cell_248_72 (.BL(BL72),.BLN(BLN72),.WL(WL248));
sram_cell_6t_5 inst_cell_248_73 (.BL(BL73),.BLN(BLN73),.WL(WL248));
sram_cell_6t_5 inst_cell_248_74 (.BL(BL74),.BLN(BLN74),.WL(WL248));
sram_cell_6t_5 inst_cell_248_75 (.BL(BL75),.BLN(BLN75),.WL(WL248));
sram_cell_6t_5 inst_cell_248_76 (.BL(BL76),.BLN(BLN76),.WL(WL248));
sram_cell_6t_5 inst_cell_248_77 (.BL(BL77),.BLN(BLN77),.WL(WL248));
sram_cell_6t_5 inst_cell_248_78 (.BL(BL78),.BLN(BLN78),.WL(WL248));
sram_cell_6t_5 inst_cell_248_79 (.BL(BL79),.BLN(BLN79),.WL(WL248));
sram_cell_6t_5 inst_cell_248_80 (.BL(BL80),.BLN(BLN80),.WL(WL248));
sram_cell_6t_5 inst_cell_248_81 (.BL(BL81),.BLN(BLN81),.WL(WL248));
sram_cell_6t_5 inst_cell_248_82 (.BL(BL82),.BLN(BLN82),.WL(WL248));
sram_cell_6t_5 inst_cell_248_83 (.BL(BL83),.BLN(BLN83),.WL(WL248));
sram_cell_6t_5 inst_cell_248_84 (.BL(BL84),.BLN(BLN84),.WL(WL248));
sram_cell_6t_5 inst_cell_248_85 (.BL(BL85),.BLN(BLN85),.WL(WL248));
sram_cell_6t_5 inst_cell_248_86 (.BL(BL86),.BLN(BLN86),.WL(WL248));
sram_cell_6t_5 inst_cell_248_87 (.BL(BL87),.BLN(BLN87),.WL(WL248));
sram_cell_6t_5 inst_cell_248_88 (.BL(BL88),.BLN(BLN88),.WL(WL248));
sram_cell_6t_5 inst_cell_248_89 (.BL(BL89),.BLN(BLN89),.WL(WL248));
sram_cell_6t_5 inst_cell_248_90 (.BL(BL90),.BLN(BLN90),.WL(WL248));
sram_cell_6t_5 inst_cell_248_91 (.BL(BL91),.BLN(BLN91),.WL(WL248));
sram_cell_6t_5 inst_cell_248_92 (.BL(BL92),.BLN(BLN92),.WL(WL248));
sram_cell_6t_5 inst_cell_248_93 (.BL(BL93),.BLN(BLN93),.WL(WL248));
sram_cell_6t_5 inst_cell_248_94 (.BL(BL94),.BLN(BLN94),.WL(WL248));
sram_cell_6t_5 inst_cell_248_95 (.BL(BL95),.BLN(BLN95),.WL(WL248));
sram_cell_6t_5 inst_cell_248_96 (.BL(BL96),.BLN(BLN96),.WL(WL248));
sram_cell_6t_5 inst_cell_248_97 (.BL(BL97),.BLN(BLN97),.WL(WL248));
sram_cell_6t_5 inst_cell_248_98 (.BL(BL98),.BLN(BLN98),.WL(WL248));
sram_cell_6t_5 inst_cell_248_99 (.BL(BL99),.BLN(BLN99),.WL(WL248));
sram_cell_6t_5 inst_cell_248_100 (.BL(BL100),.BLN(BLN100),.WL(WL248));
sram_cell_6t_5 inst_cell_248_101 (.BL(BL101),.BLN(BLN101),.WL(WL248));
sram_cell_6t_5 inst_cell_248_102 (.BL(BL102),.BLN(BLN102),.WL(WL248));
sram_cell_6t_5 inst_cell_248_103 (.BL(BL103),.BLN(BLN103),.WL(WL248));
sram_cell_6t_5 inst_cell_248_104 (.BL(BL104),.BLN(BLN104),.WL(WL248));
sram_cell_6t_5 inst_cell_248_105 (.BL(BL105),.BLN(BLN105),.WL(WL248));
sram_cell_6t_5 inst_cell_248_106 (.BL(BL106),.BLN(BLN106),.WL(WL248));
sram_cell_6t_5 inst_cell_248_107 (.BL(BL107),.BLN(BLN107),.WL(WL248));
sram_cell_6t_5 inst_cell_248_108 (.BL(BL108),.BLN(BLN108),.WL(WL248));
sram_cell_6t_5 inst_cell_248_109 (.BL(BL109),.BLN(BLN109),.WL(WL248));
sram_cell_6t_5 inst_cell_248_110 (.BL(BL110),.BLN(BLN110),.WL(WL248));
sram_cell_6t_5 inst_cell_248_111 (.BL(BL111),.BLN(BLN111),.WL(WL248));
sram_cell_6t_5 inst_cell_248_112 (.BL(BL112),.BLN(BLN112),.WL(WL248));
sram_cell_6t_5 inst_cell_248_113 (.BL(BL113),.BLN(BLN113),.WL(WL248));
sram_cell_6t_5 inst_cell_248_114 (.BL(BL114),.BLN(BLN114),.WL(WL248));
sram_cell_6t_5 inst_cell_248_115 (.BL(BL115),.BLN(BLN115),.WL(WL248));
sram_cell_6t_5 inst_cell_248_116 (.BL(BL116),.BLN(BLN116),.WL(WL248));
sram_cell_6t_5 inst_cell_248_117 (.BL(BL117),.BLN(BLN117),.WL(WL248));
sram_cell_6t_5 inst_cell_248_118 (.BL(BL118),.BLN(BLN118),.WL(WL248));
sram_cell_6t_5 inst_cell_248_119 (.BL(BL119),.BLN(BLN119),.WL(WL248));
sram_cell_6t_5 inst_cell_248_120 (.BL(BL120),.BLN(BLN120),.WL(WL248));
sram_cell_6t_5 inst_cell_248_121 (.BL(BL121),.BLN(BLN121),.WL(WL248));
sram_cell_6t_5 inst_cell_248_122 (.BL(BL122),.BLN(BLN122),.WL(WL248));
sram_cell_6t_5 inst_cell_248_123 (.BL(BL123),.BLN(BLN123),.WL(WL248));
sram_cell_6t_5 inst_cell_248_124 (.BL(BL124),.BLN(BLN124),.WL(WL248));
sram_cell_6t_5 inst_cell_248_125 (.BL(BL125),.BLN(BLN125),.WL(WL248));
sram_cell_6t_5 inst_cell_248_126 (.BL(BL126),.BLN(BLN126),.WL(WL248));
sram_cell_6t_5 inst_cell_248_127 (.BL(BL127),.BLN(BLN127),.WL(WL248));
sram_cell_6t_5 inst_cell_249_0 (.BL(BL0),.BLN(BLN0),.WL(WL249));
sram_cell_6t_5 inst_cell_249_1 (.BL(BL1),.BLN(BLN1),.WL(WL249));
sram_cell_6t_5 inst_cell_249_2 (.BL(BL2),.BLN(BLN2),.WL(WL249));
sram_cell_6t_5 inst_cell_249_3 (.BL(BL3),.BLN(BLN3),.WL(WL249));
sram_cell_6t_5 inst_cell_249_4 (.BL(BL4),.BLN(BLN4),.WL(WL249));
sram_cell_6t_5 inst_cell_249_5 (.BL(BL5),.BLN(BLN5),.WL(WL249));
sram_cell_6t_5 inst_cell_249_6 (.BL(BL6),.BLN(BLN6),.WL(WL249));
sram_cell_6t_5 inst_cell_249_7 (.BL(BL7),.BLN(BLN7),.WL(WL249));
sram_cell_6t_5 inst_cell_249_8 (.BL(BL8),.BLN(BLN8),.WL(WL249));
sram_cell_6t_5 inst_cell_249_9 (.BL(BL9),.BLN(BLN9),.WL(WL249));
sram_cell_6t_5 inst_cell_249_10 (.BL(BL10),.BLN(BLN10),.WL(WL249));
sram_cell_6t_5 inst_cell_249_11 (.BL(BL11),.BLN(BLN11),.WL(WL249));
sram_cell_6t_5 inst_cell_249_12 (.BL(BL12),.BLN(BLN12),.WL(WL249));
sram_cell_6t_5 inst_cell_249_13 (.BL(BL13),.BLN(BLN13),.WL(WL249));
sram_cell_6t_5 inst_cell_249_14 (.BL(BL14),.BLN(BLN14),.WL(WL249));
sram_cell_6t_5 inst_cell_249_15 (.BL(BL15),.BLN(BLN15),.WL(WL249));
sram_cell_6t_5 inst_cell_249_16 (.BL(BL16),.BLN(BLN16),.WL(WL249));
sram_cell_6t_5 inst_cell_249_17 (.BL(BL17),.BLN(BLN17),.WL(WL249));
sram_cell_6t_5 inst_cell_249_18 (.BL(BL18),.BLN(BLN18),.WL(WL249));
sram_cell_6t_5 inst_cell_249_19 (.BL(BL19),.BLN(BLN19),.WL(WL249));
sram_cell_6t_5 inst_cell_249_20 (.BL(BL20),.BLN(BLN20),.WL(WL249));
sram_cell_6t_5 inst_cell_249_21 (.BL(BL21),.BLN(BLN21),.WL(WL249));
sram_cell_6t_5 inst_cell_249_22 (.BL(BL22),.BLN(BLN22),.WL(WL249));
sram_cell_6t_5 inst_cell_249_23 (.BL(BL23),.BLN(BLN23),.WL(WL249));
sram_cell_6t_5 inst_cell_249_24 (.BL(BL24),.BLN(BLN24),.WL(WL249));
sram_cell_6t_5 inst_cell_249_25 (.BL(BL25),.BLN(BLN25),.WL(WL249));
sram_cell_6t_5 inst_cell_249_26 (.BL(BL26),.BLN(BLN26),.WL(WL249));
sram_cell_6t_5 inst_cell_249_27 (.BL(BL27),.BLN(BLN27),.WL(WL249));
sram_cell_6t_5 inst_cell_249_28 (.BL(BL28),.BLN(BLN28),.WL(WL249));
sram_cell_6t_5 inst_cell_249_29 (.BL(BL29),.BLN(BLN29),.WL(WL249));
sram_cell_6t_5 inst_cell_249_30 (.BL(BL30),.BLN(BLN30),.WL(WL249));
sram_cell_6t_5 inst_cell_249_31 (.BL(BL31),.BLN(BLN31),.WL(WL249));
sram_cell_6t_5 inst_cell_249_32 (.BL(BL32),.BLN(BLN32),.WL(WL249));
sram_cell_6t_5 inst_cell_249_33 (.BL(BL33),.BLN(BLN33),.WL(WL249));
sram_cell_6t_5 inst_cell_249_34 (.BL(BL34),.BLN(BLN34),.WL(WL249));
sram_cell_6t_5 inst_cell_249_35 (.BL(BL35),.BLN(BLN35),.WL(WL249));
sram_cell_6t_5 inst_cell_249_36 (.BL(BL36),.BLN(BLN36),.WL(WL249));
sram_cell_6t_5 inst_cell_249_37 (.BL(BL37),.BLN(BLN37),.WL(WL249));
sram_cell_6t_5 inst_cell_249_38 (.BL(BL38),.BLN(BLN38),.WL(WL249));
sram_cell_6t_5 inst_cell_249_39 (.BL(BL39),.BLN(BLN39),.WL(WL249));
sram_cell_6t_5 inst_cell_249_40 (.BL(BL40),.BLN(BLN40),.WL(WL249));
sram_cell_6t_5 inst_cell_249_41 (.BL(BL41),.BLN(BLN41),.WL(WL249));
sram_cell_6t_5 inst_cell_249_42 (.BL(BL42),.BLN(BLN42),.WL(WL249));
sram_cell_6t_5 inst_cell_249_43 (.BL(BL43),.BLN(BLN43),.WL(WL249));
sram_cell_6t_5 inst_cell_249_44 (.BL(BL44),.BLN(BLN44),.WL(WL249));
sram_cell_6t_5 inst_cell_249_45 (.BL(BL45),.BLN(BLN45),.WL(WL249));
sram_cell_6t_5 inst_cell_249_46 (.BL(BL46),.BLN(BLN46),.WL(WL249));
sram_cell_6t_5 inst_cell_249_47 (.BL(BL47),.BLN(BLN47),.WL(WL249));
sram_cell_6t_5 inst_cell_249_48 (.BL(BL48),.BLN(BLN48),.WL(WL249));
sram_cell_6t_5 inst_cell_249_49 (.BL(BL49),.BLN(BLN49),.WL(WL249));
sram_cell_6t_5 inst_cell_249_50 (.BL(BL50),.BLN(BLN50),.WL(WL249));
sram_cell_6t_5 inst_cell_249_51 (.BL(BL51),.BLN(BLN51),.WL(WL249));
sram_cell_6t_5 inst_cell_249_52 (.BL(BL52),.BLN(BLN52),.WL(WL249));
sram_cell_6t_5 inst_cell_249_53 (.BL(BL53),.BLN(BLN53),.WL(WL249));
sram_cell_6t_5 inst_cell_249_54 (.BL(BL54),.BLN(BLN54),.WL(WL249));
sram_cell_6t_5 inst_cell_249_55 (.BL(BL55),.BLN(BLN55),.WL(WL249));
sram_cell_6t_5 inst_cell_249_56 (.BL(BL56),.BLN(BLN56),.WL(WL249));
sram_cell_6t_5 inst_cell_249_57 (.BL(BL57),.BLN(BLN57),.WL(WL249));
sram_cell_6t_5 inst_cell_249_58 (.BL(BL58),.BLN(BLN58),.WL(WL249));
sram_cell_6t_5 inst_cell_249_59 (.BL(BL59),.BLN(BLN59),.WL(WL249));
sram_cell_6t_5 inst_cell_249_60 (.BL(BL60),.BLN(BLN60),.WL(WL249));
sram_cell_6t_5 inst_cell_249_61 (.BL(BL61),.BLN(BLN61),.WL(WL249));
sram_cell_6t_5 inst_cell_249_62 (.BL(BL62),.BLN(BLN62),.WL(WL249));
sram_cell_6t_5 inst_cell_249_63 (.BL(BL63),.BLN(BLN63),.WL(WL249));
sram_cell_6t_5 inst_cell_249_64 (.BL(BL64),.BLN(BLN64),.WL(WL249));
sram_cell_6t_5 inst_cell_249_65 (.BL(BL65),.BLN(BLN65),.WL(WL249));
sram_cell_6t_5 inst_cell_249_66 (.BL(BL66),.BLN(BLN66),.WL(WL249));
sram_cell_6t_5 inst_cell_249_67 (.BL(BL67),.BLN(BLN67),.WL(WL249));
sram_cell_6t_5 inst_cell_249_68 (.BL(BL68),.BLN(BLN68),.WL(WL249));
sram_cell_6t_5 inst_cell_249_69 (.BL(BL69),.BLN(BLN69),.WL(WL249));
sram_cell_6t_5 inst_cell_249_70 (.BL(BL70),.BLN(BLN70),.WL(WL249));
sram_cell_6t_5 inst_cell_249_71 (.BL(BL71),.BLN(BLN71),.WL(WL249));
sram_cell_6t_5 inst_cell_249_72 (.BL(BL72),.BLN(BLN72),.WL(WL249));
sram_cell_6t_5 inst_cell_249_73 (.BL(BL73),.BLN(BLN73),.WL(WL249));
sram_cell_6t_5 inst_cell_249_74 (.BL(BL74),.BLN(BLN74),.WL(WL249));
sram_cell_6t_5 inst_cell_249_75 (.BL(BL75),.BLN(BLN75),.WL(WL249));
sram_cell_6t_5 inst_cell_249_76 (.BL(BL76),.BLN(BLN76),.WL(WL249));
sram_cell_6t_5 inst_cell_249_77 (.BL(BL77),.BLN(BLN77),.WL(WL249));
sram_cell_6t_5 inst_cell_249_78 (.BL(BL78),.BLN(BLN78),.WL(WL249));
sram_cell_6t_5 inst_cell_249_79 (.BL(BL79),.BLN(BLN79),.WL(WL249));
sram_cell_6t_5 inst_cell_249_80 (.BL(BL80),.BLN(BLN80),.WL(WL249));
sram_cell_6t_5 inst_cell_249_81 (.BL(BL81),.BLN(BLN81),.WL(WL249));
sram_cell_6t_5 inst_cell_249_82 (.BL(BL82),.BLN(BLN82),.WL(WL249));
sram_cell_6t_5 inst_cell_249_83 (.BL(BL83),.BLN(BLN83),.WL(WL249));
sram_cell_6t_5 inst_cell_249_84 (.BL(BL84),.BLN(BLN84),.WL(WL249));
sram_cell_6t_5 inst_cell_249_85 (.BL(BL85),.BLN(BLN85),.WL(WL249));
sram_cell_6t_5 inst_cell_249_86 (.BL(BL86),.BLN(BLN86),.WL(WL249));
sram_cell_6t_5 inst_cell_249_87 (.BL(BL87),.BLN(BLN87),.WL(WL249));
sram_cell_6t_5 inst_cell_249_88 (.BL(BL88),.BLN(BLN88),.WL(WL249));
sram_cell_6t_5 inst_cell_249_89 (.BL(BL89),.BLN(BLN89),.WL(WL249));
sram_cell_6t_5 inst_cell_249_90 (.BL(BL90),.BLN(BLN90),.WL(WL249));
sram_cell_6t_5 inst_cell_249_91 (.BL(BL91),.BLN(BLN91),.WL(WL249));
sram_cell_6t_5 inst_cell_249_92 (.BL(BL92),.BLN(BLN92),.WL(WL249));
sram_cell_6t_5 inst_cell_249_93 (.BL(BL93),.BLN(BLN93),.WL(WL249));
sram_cell_6t_5 inst_cell_249_94 (.BL(BL94),.BLN(BLN94),.WL(WL249));
sram_cell_6t_5 inst_cell_249_95 (.BL(BL95),.BLN(BLN95),.WL(WL249));
sram_cell_6t_5 inst_cell_249_96 (.BL(BL96),.BLN(BLN96),.WL(WL249));
sram_cell_6t_5 inst_cell_249_97 (.BL(BL97),.BLN(BLN97),.WL(WL249));
sram_cell_6t_5 inst_cell_249_98 (.BL(BL98),.BLN(BLN98),.WL(WL249));
sram_cell_6t_5 inst_cell_249_99 (.BL(BL99),.BLN(BLN99),.WL(WL249));
sram_cell_6t_5 inst_cell_249_100 (.BL(BL100),.BLN(BLN100),.WL(WL249));
sram_cell_6t_5 inst_cell_249_101 (.BL(BL101),.BLN(BLN101),.WL(WL249));
sram_cell_6t_5 inst_cell_249_102 (.BL(BL102),.BLN(BLN102),.WL(WL249));
sram_cell_6t_5 inst_cell_249_103 (.BL(BL103),.BLN(BLN103),.WL(WL249));
sram_cell_6t_5 inst_cell_249_104 (.BL(BL104),.BLN(BLN104),.WL(WL249));
sram_cell_6t_5 inst_cell_249_105 (.BL(BL105),.BLN(BLN105),.WL(WL249));
sram_cell_6t_5 inst_cell_249_106 (.BL(BL106),.BLN(BLN106),.WL(WL249));
sram_cell_6t_5 inst_cell_249_107 (.BL(BL107),.BLN(BLN107),.WL(WL249));
sram_cell_6t_5 inst_cell_249_108 (.BL(BL108),.BLN(BLN108),.WL(WL249));
sram_cell_6t_5 inst_cell_249_109 (.BL(BL109),.BLN(BLN109),.WL(WL249));
sram_cell_6t_5 inst_cell_249_110 (.BL(BL110),.BLN(BLN110),.WL(WL249));
sram_cell_6t_5 inst_cell_249_111 (.BL(BL111),.BLN(BLN111),.WL(WL249));
sram_cell_6t_5 inst_cell_249_112 (.BL(BL112),.BLN(BLN112),.WL(WL249));
sram_cell_6t_5 inst_cell_249_113 (.BL(BL113),.BLN(BLN113),.WL(WL249));
sram_cell_6t_5 inst_cell_249_114 (.BL(BL114),.BLN(BLN114),.WL(WL249));
sram_cell_6t_5 inst_cell_249_115 (.BL(BL115),.BLN(BLN115),.WL(WL249));
sram_cell_6t_5 inst_cell_249_116 (.BL(BL116),.BLN(BLN116),.WL(WL249));
sram_cell_6t_5 inst_cell_249_117 (.BL(BL117),.BLN(BLN117),.WL(WL249));
sram_cell_6t_5 inst_cell_249_118 (.BL(BL118),.BLN(BLN118),.WL(WL249));
sram_cell_6t_5 inst_cell_249_119 (.BL(BL119),.BLN(BLN119),.WL(WL249));
sram_cell_6t_5 inst_cell_249_120 (.BL(BL120),.BLN(BLN120),.WL(WL249));
sram_cell_6t_5 inst_cell_249_121 (.BL(BL121),.BLN(BLN121),.WL(WL249));
sram_cell_6t_5 inst_cell_249_122 (.BL(BL122),.BLN(BLN122),.WL(WL249));
sram_cell_6t_5 inst_cell_249_123 (.BL(BL123),.BLN(BLN123),.WL(WL249));
sram_cell_6t_5 inst_cell_249_124 (.BL(BL124),.BLN(BLN124),.WL(WL249));
sram_cell_6t_5 inst_cell_249_125 (.BL(BL125),.BLN(BLN125),.WL(WL249));
sram_cell_6t_5 inst_cell_249_126 (.BL(BL126),.BLN(BLN126),.WL(WL249));
sram_cell_6t_5 inst_cell_249_127 (.BL(BL127),.BLN(BLN127),.WL(WL249));
sram_cell_6t_5 inst_cell_250_0 (.BL(BL0),.BLN(BLN0),.WL(WL250));
sram_cell_6t_5 inst_cell_250_1 (.BL(BL1),.BLN(BLN1),.WL(WL250));
sram_cell_6t_5 inst_cell_250_2 (.BL(BL2),.BLN(BLN2),.WL(WL250));
sram_cell_6t_5 inst_cell_250_3 (.BL(BL3),.BLN(BLN3),.WL(WL250));
sram_cell_6t_5 inst_cell_250_4 (.BL(BL4),.BLN(BLN4),.WL(WL250));
sram_cell_6t_5 inst_cell_250_5 (.BL(BL5),.BLN(BLN5),.WL(WL250));
sram_cell_6t_5 inst_cell_250_6 (.BL(BL6),.BLN(BLN6),.WL(WL250));
sram_cell_6t_5 inst_cell_250_7 (.BL(BL7),.BLN(BLN7),.WL(WL250));
sram_cell_6t_5 inst_cell_250_8 (.BL(BL8),.BLN(BLN8),.WL(WL250));
sram_cell_6t_5 inst_cell_250_9 (.BL(BL9),.BLN(BLN9),.WL(WL250));
sram_cell_6t_5 inst_cell_250_10 (.BL(BL10),.BLN(BLN10),.WL(WL250));
sram_cell_6t_5 inst_cell_250_11 (.BL(BL11),.BLN(BLN11),.WL(WL250));
sram_cell_6t_5 inst_cell_250_12 (.BL(BL12),.BLN(BLN12),.WL(WL250));
sram_cell_6t_5 inst_cell_250_13 (.BL(BL13),.BLN(BLN13),.WL(WL250));
sram_cell_6t_5 inst_cell_250_14 (.BL(BL14),.BLN(BLN14),.WL(WL250));
sram_cell_6t_5 inst_cell_250_15 (.BL(BL15),.BLN(BLN15),.WL(WL250));
sram_cell_6t_5 inst_cell_250_16 (.BL(BL16),.BLN(BLN16),.WL(WL250));
sram_cell_6t_5 inst_cell_250_17 (.BL(BL17),.BLN(BLN17),.WL(WL250));
sram_cell_6t_5 inst_cell_250_18 (.BL(BL18),.BLN(BLN18),.WL(WL250));
sram_cell_6t_5 inst_cell_250_19 (.BL(BL19),.BLN(BLN19),.WL(WL250));
sram_cell_6t_5 inst_cell_250_20 (.BL(BL20),.BLN(BLN20),.WL(WL250));
sram_cell_6t_5 inst_cell_250_21 (.BL(BL21),.BLN(BLN21),.WL(WL250));
sram_cell_6t_5 inst_cell_250_22 (.BL(BL22),.BLN(BLN22),.WL(WL250));
sram_cell_6t_5 inst_cell_250_23 (.BL(BL23),.BLN(BLN23),.WL(WL250));
sram_cell_6t_5 inst_cell_250_24 (.BL(BL24),.BLN(BLN24),.WL(WL250));
sram_cell_6t_5 inst_cell_250_25 (.BL(BL25),.BLN(BLN25),.WL(WL250));
sram_cell_6t_5 inst_cell_250_26 (.BL(BL26),.BLN(BLN26),.WL(WL250));
sram_cell_6t_5 inst_cell_250_27 (.BL(BL27),.BLN(BLN27),.WL(WL250));
sram_cell_6t_5 inst_cell_250_28 (.BL(BL28),.BLN(BLN28),.WL(WL250));
sram_cell_6t_5 inst_cell_250_29 (.BL(BL29),.BLN(BLN29),.WL(WL250));
sram_cell_6t_5 inst_cell_250_30 (.BL(BL30),.BLN(BLN30),.WL(WL250));
sram_cell_6t_5 inst_cell_250_31 (.BL(BL31),.BLN(BLN31),.WL(WL250));
sram_cell_6t_5 inst_cell_250_32 (.BL(BL32),.BLN(BLN32),.WL(WL250));
sram_cell_6t_5 inst_cell_250_33 (.BL(BL33),.BLN(BLN33),.WL(WL250));
sram_cell_6t_5 inst_cell_250_34 (.BL(BL34),.BLN(BLN34),.WL(WL250));
sram_cell_6t_5 inst_cell_250_35 (.BL(BL35),.BLN(BLN35),.WL(WL250));
sram_cell_6t_5 inst_cell_250_36 (.BL(BL36),.BLN(BLN36),.WL(WL250));
sram_cell_6t_5 inst_cell_250_37 (.BL(BL37),.BLN(BLN37),.WL(WL250));
sram_cell_6t_5 inst_cell_250_38 (.BL(BL38),.BLN(BLN38),.WL(WL250));
sram_cell_6t_5 inst_cell_250_39 (.BL(BL39),.BLN(BLN39),.WL(WL250));
sram_cell_6t_5 inst_cell_250_40 (.BL(BL40),.BLN(BLN40),.WL(WL250));
sram_cell_6t_5 inst_cell_250_41 (.BL(BL41),.BLN(BLN41),.WL(WL250));
sram_cell_6t_5 inst_cell_250_42 (.BL(BL42),.BLN(BLN42),.WL(WL250));
sram_cell_6t_5 inst_cell_250_43 (.BL(BL43),.BLN(BLN43),.WL(WL250));
sram_cell_6t_5 inst_cell_250_44 (.BL(BL44),.BLN(BLN44),.WL(WL250));
sram_cell_6t_5 inst_cell_250_45 (.BL(BL45),.BLN(BLN45),.WL(WL250));
sram_cell_6t_5 inst_cell_250_46 (.BL(BL46),.BLN(BLN46),.WL(WL250));
sram_cell_6t_5 inst_cell_250_47 (.BL(BL47),.BLN(BLN47),.WL(WL250));
sram_cell_6t_5 inst_cell_250_48 (.BL(BL48),.BLN(BLN48),.WL(WL250));
sram_cell_6t_5 inst_cell_250_49 (.BL(BL49),.BLN(BLN49),.WL(WL250));
sram_cell_6t_5 inst_cell_250_50 (.BL(BL50),.BLN(BLN50),.WL(WL250));
sram_cell_6t_5 inst_cell_250_51 (.BL(BL51),.BLN(BLN51),.WL(WL250));
sram_cell_6t_5 inst_cell_250_52 (.BL(BL52),.BLN(BLN52),.WL(WL250));
sram_cell_6t_5 inst_cell_250_53 (.BL(BL53),.BLN(BLN53),.WL(WL250));
sram_cell_6t_5 inst_cell_250_54 (.BL(BL54),.BLN(BLN54),.WL(WL250));
sram_cell_6t_5 inst_cell_250_55 (.BL(BL55),.BLN(BLN55),.WL(WL250));
sram_cell_6t_5 inst_cell_250_56 (.BL(BL56),.BLN(BLN56),.WL(WL250));
sram_cell_6t_5 inst_cell_250_57 (.BL(BL57),.BLN(BLN57),.WL(WL250));
sram_cell_6t_5 inst_cell_250_58 (.BL(BL58),.BLN(BLN58),.WL(WL250));
sram_cell_6t_5 inst_cell_250_59 (.BL(BL59),.BLN(BLN59),.WL(WL250));
sram_cell_6t_5 inst_cell_250_60 (.BL(BL60),.BLN(BLN60),.WL(WL250));
sram_cell_6t_5 inst_cell_250_61 (.BL(BL61),.BLN(BLN61),.WL(WL250));
sram_cell_6t_5 inst_cell_250_62 (.BL(BL62),.BLN(BLN62),.WL(WL250));
sram_cell_6t_5 inst_cell_250_63 (.BL(BL63),.BLN(BLN63),.WL(WL250));
sram_cell_6t_5 inst_cell_250_64 (.BL(BL64),.BLN(BLN64),.WL(WL250));
sram_cell_6t_5 inst_cell_250_65 (.BL(BL65),.BLN(BLN65),.WL(WL250));
sram_cell_6t_5 inst_cell_250_66 (.BL(BL66),.BLN(BLN66),.WL(WL250));
sram_cell_6t_5 inst_cell_250_67 (.BL(BL67),.BLN(BLN67),.WL(WL250));
sram_cell_6t_5 inst_cell_250_68 (.BL(BL68),.BLN(BLN68),.WL(WL250));
sram_cell_6t_5 inst_cell_250_69 (.BL(BL69),.BLN(BLN69),.WL(WL250));
sram_cell_6t_5 inst_cell_250_70 (.BL(BL70),.BLN(BLN70),.WL(WL250));
sram_cell_6t_5 inst_cell_250_71 (.BL(BL71),.BLN(BLN71),.WL(WL250));
sram_cell_6t_5 inst_cell_250_72 (.BL(BL72),.BLN(BLN72),.WL(WL250));
sram_cell_6t_5 inst_cell_250_73 (.BL(BL73),.BLN(BLN73),.WL(WL250));
sram_cell_6t_5 inst_cell_250_74 (.BL(BL74),.BLN(BLN74),.WL(WL250));
sram_cell_6t_5 inst_cell_250_75 (.BL(BL75),.BLN(BLN75),.WL(WL250));
sram_cell_6t_5 inst_cell_250_76 (.BL(BL76),.BLN(BLN76),.WL(WL250));
sram_cell_6t_5 inst_cell_250_77 (.BL(BL77),.BLN(BLN77),.WL(WL250));
sram_cell_6t_5 inst_cell_250_78 (.BL(BL78),.BLN(BLN78),.WL(WL250));
sram_cell_6t_5 inst_cell_250_79 (.BL(BL79),.BLN(BLN79),.WL(WL250));
sram_cell_6t_5 inst_cell_250_80 (.BL(BL80),.BLN(BLN80),.WL(WL250));
sram_cell_6t_5 inst_cell_250_81 (.BL(BL81),.BLN(BLN81),.WL(WL250));
sram_cell_6t_5 inst_cell_250_82 (.BL(BL82),.BLN(BLN82),.WL(WL250));
sram_cell_6t_5 inst_cell_250_83 (.BL(BL83),.BLN(BLN83),.WL(WL250));
sram_cell_6t_5 inst_cell_250_84 (.BL(BL84),.BLN(BLN84),.WL(WL250));
sram_cell_6t_5 inst_cell_250_85 (.BL(BL85),.BLN(BLN85),.WL(WL250));
sram_cell_6t_5 inst_cell_250_86 (.BL(BL86),.BLN(BLN86),.WL(WL250));
sram_cell_6t_5 inst_cell_250_87 (.BL(BL87),.BLN(BLN87),.WL(WL250));
sram_cell_6t_5 inst_cell_250_88 (.BL(BL88),.BLN(BLN88),.WL(WL250));
sram_cell_6t_5 inst_cell_250_89 (.BL(BL89),.BLN(BLN89),.WL(WL250));
sram_cell_6t_5 inst_cell_250_90 (.BL(BL90),.BLN(BLN90),.WL(WL250));
sram_cell_6t_5 inst_cell_250_91 (.BL(BL91),.BLN(BLN91),.WL(WL250));
sram_cell_6t_5 inst_cell_250_92 (.BL(BL92),.BLN(BLN92),.WL(WL250));
sram_cell_6t_5 inst_cell_250_93 (.BL(BL93),.BLN(BLN93),.WL(WL250));
sram_cell_6t_5 inst_cell_250_94 (.BL(BL94),.BLN(BLN94),.WL(WL250));
sram_cell_6t_5 inst_cell_250_95 (.BL(BL95),.BLN(BLN95),.WL(WL250));
sram_cell_6t_5 inst_cell_250_96 (.BL(BL96),.BLN(BLN96),.WL(WL250));
sram_cell_6t_5 inst_cell_250_97 (.BL(BL97),.BLN(BLN97),.WL(WL250));
sram_cell_6t_5 inst_cell_250_98 (.BL(BL98),.BLN(BLN98),.WL(WL250));
sram_cell_6t_5 inst_cell_250_99 (.BL(BL99),.BLN(BLN99),.WL(WL250));
sram_cell_6t_5 inst_cell_250_100 (.BL(BL100),.BLN(BLN100),.WL(WL250));
sram_cell_6t_5 inst_cell_250_101 (.BL(BL101),.BLN(BLN101),.WL(WL250));
sram_cell_6t_5 inst_cell_250_102 (.BL(BL102),.BLN(BLN102),.WL(WL250));
sram_cell_6t_5 inst_cell_250_103 (.BL(BL103),.BLN(BLN103),.WL(WL250));
sram_cell_6t_5 inst_cell_250_104 (.BL(BL104),.BLN(BLN104),.WL(WL250));
sram_cell_6t_5 inst_cell_250_105 (.BL(BL105),.BLN(BLN105),.WL(WL250));
sram_cell_6t_5 inst_cell_250_106 (.BL(BL106),.BLN(BLN106),.WL(WL250));
sram_cell_6t_5 inst_cell_250_107 (.BL(BL107),.BLN(BLN107),.WL(WL250));
sram_cell_6t_5 inst_cell_250_108 (.BL(BL108),.BLN(BLN108),.WL(WL250));
sram_cell_6t_5 inst_cell_250_109 (.BL(BL109),.BLN(BLN109),.WL(WL250));
sram_cell_6t_5 inst_cell_250_110 (.BL(BL110),.BLN(BLN110),.WL(WL250));
sram_cell_6t_5 inst_cell_250_111 (.BL(BL111),.BLN(BLN111),.WL(WL250));
sram_cell_6t_5 inst_cell_250_112 (.BL(BL112),.BLN(BLN112),.WL(WL250));
sram_cell_6t_5 inst_cell_250_113 (.BL(BL113),.BLN(BLN113),.WL(WL250));
sram_cell_6t_5 inst_cell_250_114 (.BL(BL114),.BLN(BLN114),.WL(WL250));
sram_cell_6t_5 inst_cell_250_115 (.BL(BL115),.BLN(BLN115),.WL(WL250));
sram_cell_6t_5 inst_cell_250_116 (.BL(BL116),.BLN(BLN116),.WL(WL250));
sram_cell_6t_5 inst_cell_250_117 (.BL(BL117),.BLN(BLN117),.WL(WL250));
sram_cell_6t_5 inst_cell_250_118 (.BL(BL118),.BLN(BLN118),.WL(WL250));
sram_cell_6t_5 inst_cell_250_119 (.BL(BL119),.BLN(BLN119),.WL(WL250));
sram_cell_6t_5 inst_cell_250_120 (.BL(BL120),.BLN(BLN120),.WL(WL250));
sram_cell_6t_5 inst_cell_250_121 (.BL(BL121),.BLN(BLN121),.WL(WL250));
sram_cell_6t_5 inst_cell_250_122 (.BL(BL122),.BLN(BLN122),.WL(WL250));
sram_cell_6t_5 inst_cell_250_123 (.BL(BL123),.BLN(BLN123),.WL(WL250));
sram_cell_6t_5 inst_cell_250_124 (.BL(BL124),.BLN(BLN124),.WL(WL250));
sram_cell_6t_5 inst_cell_250_125 (.BL(BL125),.BLN(BLN125),.WL(WL250));
sram_cell_6t_5 inst_cell_250_126 (.BL(BL126),.BLN(BLN126),.WL(WL250));
sram_cell_6t_5 inst_cell_250_127 (.BL(BL127),.BLN(BLN127),.WL(WL250));
sram_cell_6t_5 inst_cell_251_0 (.BL(BL0),.BLN(BLN0),.WL(WL251));
sram_cell_6t_5 inst_cell_251_1 (.BL(BL1),.BLN(BLN1),.WL(WL251));
sram_cell_6t_5 inst_cell_251_2 (.BL(BL2),.BLN(BLN2),.WL(WL251));
sram_cell_6t_5 inst_cell_251_3 (.BL(BL3),.BLN(BLN3),.WL(WL251));
sram_cell_6t_5 inst_cell_251_4 (.BL(BL4),.BLN(BLN4),.WL(WL251));
sram_cell_6t_5 inst_cell_251_5 (.BL(BL5),.BLN(BLN5),.WL(WL251));
sram_cell_6t_5 inst_cell_251_6 (.BL(BL6),.BLN(BLN6),.WL(WL251));
sram_cell_6t_5 inst_cell_251_7 (.BL(BL7),.BLN(BLN7),.WL(WL251));
sram_cell_6t_5 inst_cell_251_8 (.BL(BL8),.BLN(BLN8),.WL(WL251));
sram_cell_6t_5 inst_cell_251_9 (.BL(BL9),.BLN(BLN9),.WL(WL251));
sram_cell_6t_5 inst_cell_251_10 (.BL(BL10),.BLN(BLN10),.WL(WL251));
sram_cell_6t_5 inst_cell_251_11 (.BL(BL11),.BLN(BLN11),.WL(WL251));
sram_cell_6t_5 inst_cell_251_12 (.BL(BL12),.BLN(BLN12),.WL(WL251));
sram_cell_6t_5 inst_cell_251_13 (.BL(BL13),.BLN(BLN13),.WL(WL251));
sram_cell_6t_5 inst_cell_251_14 (.BL(BL14),.BLN(BLN14),.WL(WL251));
sram_cell_6t_5 inst_cell_251_15 (.BL(BL15),.BLN(BLN15),.WL(WL251));
sram_cell_6t_5 inst_cell_251_16 (.BL(BL16),.BLN(BLN16),.WL(WL251));
sram_cell_6t_5 inst_cell_251_17 (.BL(BL17),.BLN(BLN17),.WL(WL251));
sram_cell_6t_5 inst_cell_251_18 (.BL(BL18),.BLN(BLN18),.WL(WL251));
sram_cell_6t_5 inst_cell_251_19 (.BL(BL19),.BLN(BLN19),.WL(WL251));
sram_cell_6t_5 inst_cell_251_20 (.BL(BL20),.BLN(BLN20),.WL(WL251));
sram_cell_6t_5 inst_cell_251_21 (.BL(BL21),.BLN(BLN21),.WL(WL251));
sram_cell_6t_5 inst_cell_251_22 (.BL(BL22),.BLN(BLN22),.WL(WL251));
sram_cell_6t_5 inst_cell_251_23 (.BL(BL23),.BLN(BLN23),.WL(WL251));
sram_cell_6t_5 inst_cell_251_24 (.BL(BL24),.BLN(BLN24),.WL(WL251));
sram_cell_6t_5 inst_cell_251_25 (.BL(BL25),.BLN(BLN25),.WL(WL251));
sram_cell_6t_5 inst_cell_251_26 (.BL(BL26),.BLN(BLN26),.WL(WL251));
sram_cell_6t_5 inst_cell_251_27 (.BL(BL27),.BLN(BLN27),.WL(WL251));
sram_cell_6t_5 inst_cell_251_28 (.BL(BL28),.BLN(BLN28),.WL(WL251));
sram_cell_6t_5 inst_cell_251_29 (.BL(BL29),.BLN(BLN29),.WL(WL251));
sram_cell_6t_5 inst_cell_251_30 (.BL(BL30),.BLN(BLN30),.WL(WL251));
sram_cell_6t_5 inst_cell_251_31 (.BL(BL31),.BLN(BLN31),.WL(WL251));
sram_cell_6t_5 inst_cell_251_32 (.BL(BL32),.BLN(BLN32),.WL(WL251));
sram_cell_6t_5 inst_cell_251_33 (.BL(BL33),.BLN(BLN33),.WL(WL251));
sram_cell_6t_5 inst_cell_251_34 (.BL(BL34),.BLN(BLN34),.WL(WL251));
sram_cell_6t_5 inst_cell_251_35 (.BL(BL35),.BLN(BLN35),.WL(WL251));
sram_cell_6t_5 inst_cell_251_36 (.BL(BL36),.BLN(BLN36),.WL(WL251));
sram_cell_6t_5 inst_cell_251_37 (.BL(BL37),.BLN(BLN37),.WL(WL251));
sram_cell_6t_5 inst_cell_251_38 (.BL(BL38),.BLN(BLN38),.WL(WL251));
sram_cell_6t_5 inst_cell_251_39 (.BL(BL39),.BLN(BLN39),.WL(WL251));
sram_cell_6t_5 inst_cell_251_40 (.BL(BL40),.BLN(BLN40),.WL(WL251));
sram_cell_6t_5 inst_cell_251_41 (.BL(BL41),.BLN(BLN41),.WL(WL251));
sram_cell_6t_5 inst_cell_251_42 (.BL(BL42),.BLN(BLN42),.WL(WL251));
sram_cell_6t_5 inst_cell_251_43 (.BL(BL43),.BLN(BLN43),.WL(WL251));
sram_cell_6t_5 inst_cell_251_44 (.BL(BL44),.BLN(BLN44),.WL(WL251));
sram_cell_6t_5 inst_cell_251_45 (.BL(BL45),.BLN(BLN45),.WL(WL251));
sram_cell_6t_5 inst_cell_251_46 (.BL(BL46),.BLN(BLN46),.WL(WL251));
sram_cell_6t_5 inst_cell_251_47 (.BL(BL47),.BLN(BLN47),.WL(WL251));
sram_cell_6t_5 inst_cell_251_48 (.BL(BL48),.BLN(BLN48),.WL(WL251));
sram_cell_6t_5 inst_cell_251_49 (.BL(BL49),.BLN(BLN49),.WL(WL251));
sram_cell_6t_5 inst_cell_251_50 (.BL(BL50),.BLN(BLN50),.WL(WL251));
sram_cell_6t_5 inst_cell_251_51 (.BL(BL51),.BLN(BLN51),.WL(WL251));
sram_cell_6t_5 inst_cell_251_52 (.BL(BL52),.BLN(BLN52),.WL(WL251));
sram_cell_6t_5 inst_cell_251_53 (.BL(BL53),.BLN(BLN53),.WL(WL251));
sram_cell_6t_5 inst_cell_251_54 (.BL(BL54),.BLN(BLN54),.WL(WL251));
sram_cell_6t_5 inst_cell_251_55 (.BL(BL55),.BLN(BLN55),.WL(WL251));
sram_cell_6t_5 inst_cell_251_56 (.BL(BL56),.BLN(BLN56),.WL(WL251));
sram_cell_6t_5 inst_cell_251_57 (.BL(BL57),.BLN(BLN57),.WL(WL251));
sram_cell_6t_5 inst_cell_251_58 (.BL(BL58),.BLN(BLN58),.WL(WL251));
sram_cell_6t_5 inst_cell_251_59 (.BL(BL59),.BLN(BLN59),.WL(WL251));
sram_cell_6t_5 inst_cell_251_60 (.BL(BL60),.BLN(BLN60),.WL(WL251));
sram_cell_6t_5 inst_cell_251_61 (.BL(BL61),.BLN(BLN61),.WL(WL251));
sram_cell_6t_5 inst_cell_251_62 (.BL(BL62),.BLN(BLN62),.WL(WL251));
sram_cell_6t_5 inst_cell_251_63 (.BL(BL63),.BLN(BLN63),.WL(WL251));
sram_cell_6t_5 inst_cell_251_64 (.BL(BL64),.BLN(BLN64),.WL(WL251));
sram_cell_6t_5 inst_cell_251_65 (.BL(BL65),.BLN(BLN65),.WL(WL251));
sram_cell_6t_5 inst_cell_251_66 (.BL(BL66),.BLN(BLN66),.WL(WL251));
sram_cell_6t_5 inst_cell_251_67 (.BL(BL67),.BLN(BLN67),.WL(WL251));
sram_cell_6t_5 inst_cell_251_68 (.BL(BL68),.BLN(BLN68),.WL(WL251));
sram_cell_6t_5 inst_cell_251_69 (.BL(BL69),.BLN(BLN69),.WL(WL251));
sram_cell_6t_5 inst_cell_251_70 (.BL(BL70),.BLN(BLN70),.WL(WL251));
sram_cell_6t_5 inst_cell_251_71 (.BL(BL71),.BLN(BLN71),.WL(WL251));
sram_cell_6t_5 inst_cell_251_72 (.BL(BL72),.BLN(BLN72),.WL(WL251));
sram_cell_6t_5 inst_cell_251_73 (.BL(BL73),.BLN(BLN73),.WL(WL251));
sram_cell_6t_5 inst_cell_251_74 (.BL(BL74),.BLN(BLN74),.WL(WL251));
sram_cell_6t_5 inst_cell_251_75 (.BL(BL75),.BLN(BLN75),.WL(WL251));
sram_cell_6t_5 inst_cell_251_76 (.BL(BL76),.BLN(BLN76),.WL(WL251));
sram_cell_6t_5 inst_cell_251_77 (.BL(BL77),.BLN(BLN77),.WL(WL251));
sram_cell_6t_5 inst_cell_251_78 (.BL(BL78),.BLN(BLN78),.WL(WL251));
sram_cell_6t_5 inst_cell_251_79 (.BL(BL79),.BLN(BLN79),.WL(WL251));
sram_cell_6t_5 inst_cell_251_80 (.BL(BL80),.BLN(BLN80),.WL(WL251));
sram_cell_6t_5 inst_cell_251_81 (.BL(BL81),.BLN(BLN81),.WL(WL251));
sram_cell_6t_5 inst_cell_251_82 (.BL(BL82),.BLN(BLN82),.WL(WL251));
sram_cell_6t_5 inst_cell_251_83 (.BL(BL83),.BLN(BLN83),.WL(WL251));
sram_cell_6t_5 inst_cell_251_84 (.BL(BL84),.BLN(BLN84),.WL(WL251));
sram_cell_6t_5 inst_cell_251_85 (.BL(BL85),.BLN(BLN85),.WL(WL251));
sram_cell_6t_5 inst_cell_251_86 (.BL(BL86),.BLN(BLN86),.WL(WL251));
sram_cell_6t_5 inst_cell_251_87 (.BL(BL87),.BLN(BLN87),.WL(WL251));
sram_cell_6t_5 inst_cell_251_88 (.BL(BL88),.BLN(BLN88),.WL(WL251));
sram_cell_6t_5 inst_cell_251_89 (.BL(BL89),.BLN(BLN89),.WL(WL251));
sram_cell_6t_5 inst_cell_251_90 (.BL(BL90),.BLN(BLN90),.WL(WL251));
sram_cell_6t_5 inst_cell_251_91 (.BL(BL91),.BLN(BLN91),.WL(WL251));
sram_cell_6t_5 inst_cell_251_92 (.BL(BL92),.BLN(BLN92),.WL(WL251));
sram_cell_6t_5 inst_cell_251_93 (.BL(BL93),.BLN(BLN93),.WL(WL251));
sram_cell_6t_5 inst_cell_251_94 (.BL(BL94),.BLN(BLN94),.WL(WL251));
sram_cell_6t_5 inst_cell_251_95 (.BL(BL95),.BLN(BLN95),.WL(WL251));
sram_cell_6t_5 inst_cell_251_96 (.BL(BL96),.BLN(BLN96),.WL(WL251));
sram_cell_6t_5 inst_cell_251_97 (.BL(BL97),.BLN(BLN97),.WL(WL251));
sram_cell_6t_5 inst_cell_251_98 (.BL(BL98),.BLN(BLN98),.WL(WL251));
sram_cell_6t_5 inst_cell_251_99 (.BL(BL99),.BLN(BLN99),.WL(WL251));
sram_cell_6t_5 inst_cell_251_100 (.BL(BL100),.BLN(BLN100),.WL(WL251));
sram_cell_6t_5 inst_cell_251_101 (.BL(BL101),.BLN(BLN101),.WL(WL251));
sram_cell_6t_5 inst_cell_251_102 (.BL(BL102),.BLN(BLN102),.WL(WL251));
sram_cell_6t_5 inst_cell_251_103 (.BL(BL103),.BLN(BLN103),.WL(WL251));
sram_cell_6t_5 inst_cell_251_104 (.BL(BL104),.BLN(BLN104),.WL(WL251));
sram_cell_6t_5 inst_cell_251_105 (.BL(BL105),.BLN(BLN105),.WL(WL251));
sram_cell_6t_5 inst_cell_251_106 (.BL(BL106),.BLN(BLN106),.WL(WL251));
sram_cell_6t_5 inst_cell_251_107 (.BL(BL107),.BLN(BLN107),.WL(WL251));
sram_cell_6t_5 inst_cell_251_108 (.BL(BL108),.BLN(BLN108),.WL(WL251));
sram_cell_6t_5 inst_cell_251_109 (.BL(BL109),.BLN(BLN109),.WL(WL251));
sram_cell_6t_5 inst_cell_251_110 (.BL(BL110),.BLN(BLN110),.WL(WL251));
sram_cell_6t_5 inst_cell_251_111 (.BL(BL111),.BLN(BLN111),.WL(WL251));
sram_cell_6t_5 inst_cell_251_112 (.BL(BL112),.BLN(BLN112),.WL(WL251));
sram_cell_6t_5 inst_cell_251_113 (.BL(BL113),.BLN(BLN113),.WL(WL251));
sram_cell_6t_5 inst_cell_251_114 (.BL(BL114),.BLN(BLN114),.WL(WL251));
sram_cell_6t_5 inst_cell_251_115 (.BL(BL115),.BLN(BLN115),.WL(WL251));
sram_cell_6t_5 inst_cell_251_116 (.BL(BL116),.BLN(BLN116),.WL(WL251));
sram_cell_6t_5 inst_cell_251_117 (.BL(BL117),.BLN(BLN117),.WL(WL251));
sram_cell_6t_5 inst_cell_251_118 (.BL(BL118),.BLN(BLN118),.WL(WL251));
sram_cell_6t_5 inst_cell_251_119 (.BL(BL119),.BLN(BLN119),.WL(WL251));
sram_cell_6t_5 inst_cell_251_120 (.BL(BL120),.BLN(BLN120),.WL(WL251));
sram_cell_6t_5 inst_cell_251_121 (.BL(BL121),.BLN(BLN121),.WL(WL251));
sram_cell_6t_5 inst_cell_251_122 (.BL(BL122),.BLN(BLN122),.WL(WL251));
sram_cell_6t_5 inst_cell_251_123 (.BL(BL123),.BLN(BLN123),.WL(WL251));
sram_cell_6t_5 inst_cell_251_124 (.BL(BL124),.BLN(BLN124),.WL(WL251));
sram_cell_6t_5 inst_cell_251_125 (.BL(BL125),.BLN(BLN125),.WL(WL251));
sram_cell_6t_5 inst_cell_251_126 (.BL(BL126),.BLN(BLN126),.WL(WL251));
sram_cell_6t_5 inst_cell_251_127 (.BL(BL127),.BLN(BLN127),.WL(WL251));
sram_cell_6t_5 inst_cell_252_0 (.BL(BL0),.BLN(BLN0),.WL(WL252));
sram_cell_6t_5 inst_cell_252_1 (.BL(BL1),.BLN(BLN1),.WL(WL252));
sram_cell_6t_5 inst_cell_252_2 (.BL(BL2),.BLN(BLN2),.WL(WL252));
sram_cell_6t_5 inst_cell_252_3 (.BL(BL3),.BLN(BLN3),.WL(WL252));
sram_cell_6t_5 inst_cell_252_4 (.BL(BL4),.BLN(BLN4),.WL(WL252));
sram_cell_6t_5 inst_cell_252_5 (.BL(BL5),.BLN(BLN5),.WL(WL252));
sram_cell_6t_5 inst_cell_252_6 (.BL(BL6),.BLN(BLN6),.WL(WL252));
sram_cell_6t_5 inst_cell_252_7 (.BL(BL7),.BLN(BLN7),.WL(WL252));
sram_cell_6t_5 inst_cell_252_8 (.BL(BL8),.BLN(BLN8),.WL(WL252));
sram_cell_6t_5 inst_cell_252_9 (.BL(BL9),.BLN(BLN9),.WL(WL252));
sram_cell_6t_5 inst_cell_252_10 (.BL(BL10),.BLN(BLN10),.WL(WL252));
sram_cell_6t_5 inst_cell_252_11 (.BL(BL11),.BLN(BLN11),.WL(WL252));
sram_cell_6t_5 inst_cell_252_12 (.BL(BL12),.BLN(BLN12),.WL(WL252));
sram_cell_6t_5 inst_cell_252_13 (.BL(BL13),.BLN(BLN13),.WL(WL252));
sram_cell_6t_5 inst_cell_252_14 (.BL(BL14),.BLN(BLN14),.WL(WL252));
sram_cell_6t_5 inst_cell_252_15 (.BL(BL15),.BLN(BLN15),.WL(WL252));
sram_cell_6t_5 inst_cell_252_16 (.BL(BL16),.BLN(BLN16),.WL(WL252));
sram_cell_6t_5 inst_cell_252_17 (.BL(BL17),.BLN(BLN17),.WL(WL252));
sram_cell_6t_5 inst_cell_252_18 (.BL(BL18),.BLN(BLN18),.WL(WL252));
sram_cell_6t_5 inst_cell_252_19 (.BL(BL19),.BLN(BLN19),.WL(WL252));
sram_cell_6t_5 inst_cell_252_20 (.BL(BL20),.BLN(BLN20),.WL(WL252));
sram_cell_6t_5 inst_cell_252_21 (.BL(BL21),.BLN(BLN21),.WL(WL252));
sram_cell_6t_5 inst_cell_252_22 (.BL(BL22),.BLN(BLN22),.WL(WL252));
sram_cell_6t_5 inst_cell_252_23 (.BL(BL23),.BLN(BLN23),.WL(WL252));
sram_cell_6t_5 inst_cell_252_24 (.BL(BL24),.BLN(BLN24),.WL(WL252));
sram_cell_6t_5 inst_cell_252_25 (.BL(BL25),.BLN(BLN25),.WL(WL252));
sram_cell_6t_5 inst_cell_252_26 (.BL(BL26),.BLN(BLN26),.WL(WL252));
sram_cell_6t_5 inst_cell_252_27 (.BL(BL27),.BLN(BLN27),.WL(WL252));
sram_cell_6t_5 inst_cell_252_28 (.BL(BL28),.BLN(BLN28),.WL(WL252));
sram_cell_6t_5 inst_cell_252_29 (.BL(BL29),.BLN(BLN29),.WL(WL252));
sram_cell_6t_5 inst_cell_252_30 (.BL(BL30),.BLN(BLN30),.WL(WL252));
sram_cell_6t_5 inst_cell_252_31 (.BL(BL31),.BLN(BLN31),.WL(WL252));
sram_cell_6t_5 inst_cell_252_32 (.BL(BL32),.BLN(BLN32),.WL(WL252));
sram_cell_6t_5 inst_cell_252_33 (.BL(BL33),.BLN(BLN33),.WL(WL252));
sram_cell_6t_5 inst_cell_252_34 (.BL(BL34),.BLN(BLN34),.WL(WL252));
sram_cell_6t_5 inst_cell_252_35 (.BL(BL35),.BLN(BLN35),.WL(WL252));
sram_cell_6t_5 inst_cell_252_36 (.BL(BL36),.BLN(BLN36),.WL(WL252));
sram_cell_6t_5 inst_cell_252_37 (.BL(BL37),.BLN(BLN37),.WL(WL252));
sram_cell_6t_5 inst_cell_252_38 (.BL(BL38),.BLN(BLN38),.WL(WL252));
sram_cell_6t_5 inst_cell_252_39 (.BL(BL39),.BLN(BLN39),.WL(WL252));
sram_cell_6t_5 inst_cell_252_40 (.BL(BL40),.BLN(BLN40),.WL(WL252));
sram_cell_6t_5 inst_cell_252_41 (.BL(BL41),.BLN(BLN41),.WL(WL252));
sram_cell_6t_5 inst_cell_252_42 (.BL(BL42),.BLN(BLN42),.WL(WL252));
sram_cell_6t_5 inst_cell_252_43 (.BL(BL43),.BLN(BLN43),.WL(WL252));
sram_cell_6t_5 inst_cell_252_44 (.BL(BL44),.BLN(BLN44),.WL(WL252));
sram_cell_6t_5 inst_cell_252_45 (.BL(BL45),.BLN(BLN45),.WL(WL252));
sram_cell_6t_5 inst_cell_252_46 (.BL(BL46),.BLN(BLN46),.WL(WL252));
sram_cell_6t_5 inst_cell_252_47 (.BL(BL47),.BLN(BLN47),.WL(WL252));
sram_cell_6t_5 inst_cell_252_48 (.BL(BL48),.BLN(BLN48),.WL(WL252));
sram_cell_6t_5 inst_cell_252_49 (.BL(BL49),.BLN(BLN49),.WL(WL252));
sram_cell_6t_5 inst_cell_252_50 (.BL(BL50),.BLN(BLN50),.WL(WL252));
sram_cell_6t_5 inst_cell_252_51 (.BL(BL51),.BLN(BLN51),.WL(WL252));
sram_cell_6t_5 inst_cell_252_52 (.BL(BL52),.BLN(BLN52),.WL(WL252));
sram_cell_6t_5 inst_cell_252_53 (.BL(BL53),.BLN(BLN53),.WL(WL252));
sram_cell_6t_5 inst_cell_252_54 (.BL(BL54),.BLN(BLN54),.WL(WL252));
sram_cell_6t_5 inst_cell_252_55 (.BL(BL55),.BLN(BLN55),.WL(WL252));
sram_cell_6t_5 inst_cell_252_56 (.BL(BL56),.BLN(BLN56),.WL(WL252));
sram_cell_6t_5 inst_cell_252_57 (.BL(BL57),.BLN(BLN57),.WL(WL252));
sram_cell_6t_5 inst_cell_252_58 (.BL(BL58),.BLN(BLN58),.WL(WL252));
sram_cell_6t_5 inst_cell_252_59 (.BL(BL59),.BLN(BLN59),.WL(WL252));
sram_cell_6t_5 inst_cell_252_60 (.BL(BL60),.BLN(BLN60),.WL(WL252));
sram_cell_6t_5 inst_cell_252_61 (.BL(BL61),.BLN(BLN61),.WL(WL252));
sram_cell_6t_5 inst_cell_252_62 (.BL(BL62),.BLN(BLN62),.WL(WL252));
sram_cell_6t_5 inst_cell_252_63 (.BL(BL63),.BLN(BLN63),.WL(WL252));
sram_cell_6t_5 inst_cell_252_64 (.BL(BL64),.BLN(BLN64),.WL(WL252));
sram_cell_6t_5 inst_cell_252_65 (.BL(BL65),.BLN(BLN65),.WL(WL252));
sram_cell_6t_5 inst_cell_252_66 (.BL(BL66),.BLN(BLN66),.WL(WL252));
sram_cell_6t_5 inst_cell_252_67 (.BL(BL67),.BLN(BLN67),.WL(WL252));
sram_cell_6t_5 inst_cell_252_68 (.BL(BL68),.BLN(BLN68),.WL(WL252));
sram_cell_6t_5 inst_cell_252_69 (.BL(BL69),.BLN(BLN69),.WL(WL252));
sram_cell_6t_5 inst_cell_252_70 (.BL(BL70),.BLN(BLN70),.WL(WL252));
sram_cell_6t_5 inst_cell_252_71 (.BL(BL71),.BLN(BLN71),.WL(WL252));
sram_cell_6t_5 inst_cell_252_72 (.BL(BL72),.BLN(BLN72),.WL(WL252));
sram_cell_6t_5 inst_cell_252_73 (.BL(BL73),.BLN(BLN73),.WL(WL252));
sram_cell_6t_5 inst_cell_252_74 (.BL(BL74),.BLN(BLN74),.WL(WL252));
sram_cell_6t_5 inst_cell_252_75 (.BL(BL75),.BLN(BLN75),.WL(WL252));
sram_cell_6t_5 inst_cell_252_76 (.BL(BL76),.BLN(BLN76),.WL(WL252));
sram_cell_6t_5 inst_cell_252_77 (.BL(BL77),.BLN(BLN77),.WL(WL252));
sram_cell_6t_5 inst_cell_252_78 (.BL(BL78),.BLN(BLN78),.WL(WL252));
sram_cell_6t_5 inst_cell_252_79 (.BL(BL79),.BLN(BLN79),.WL(WL252));
sram_cell_6t_5 inst_cell_252_80 (.BL(BL80),.BLN(BLN80),.WL(WL252));
sram_cell_6t_5 inst_cell_252_81 (.BL(BL81),.BLN(BLN81),.WL(WL252));
sram_cell_6t_5 inst_cell_252_82 (.BL(BL82),.BLN(BLN82),.WL(WL252));
sram_cell_6t_5 inst_cell_252_83 (.BL(BL83),.BLN(BLN83),.WL(WL252));
sram_cell_6t_5 inst_cell_252_84 (.BL(BL84),.BLN(BLN84),.WL(WL252));
sram_cell_6t_5 inst_cell_252_85 (.BL(BL85),.BLN(BLN85),.WL(WL252));
sram_cell_6t_5 inst_cell_252_86 (.BL(BL86),.BLN(BLN86),.WL(WL252));
sram_cell_6t_5 inst_cell_252_87 (.BL(BL87),.BLN(BLN87),.WL(WL252));
sram_cell_6t_5 inst_cell_252_88 (.BL(BL88),.BLN(BLN88),.WL(WL252));
sram_cell_6t_5 inst_cell_252_89 (.BL(BL89),.BLN(BLN89),.WL(WL252));
sram_cell_6t_5 inst_cell_252_90 (.BL(BL90),.BLN(BLN90),.WL(WL252));
sram_cell_6t_5 inst_cell_252_91 (.BL(BL91),.BLN(BLN91),.WL(WL252));
sram_cell_6t_5 inst_cell_252_92 (.BL(BL92),.BLN(BLN92),.WL(WL252));
sram_cell_6t_5 inst_cell_252_93 (.BL(BL93),.BLN(BLN93),.WL(WL252));
sram_cell_6t_5 inst_cell_252_94 (.BL(BL94),.BLN(BLN94),.WL(WL252));
sram_cell_6t_5 inst_cell_252_95 (.BL(BL95),.BLN(BLN95),.WL(WL252));
sram_cell_6t_5 inst_cell_252_96 (.BL(BL96),.BLN(BLN96),.WL(WL252));
sram_cell_6t_5 inst_cell_252_97 (.BL(BL97),.BLN(BLN97),.WL(WL252));
sram_cell_6t_5 inst_cell_252_98 (.BL(BL98),.BLN(BLN98),.WL(WL252));
sram_cell_6t_5 inst_cell_252_99 (.BL(BL99),.BLN(BLN99),.WL(WL252));
sram_cell_6t_5 inst_cell_252_100 (.BL(BL100),.BLN(BLN100),.WL(WL252));
sram_cell_6t_5 inst_cell_252_101 (.BL(BL101),.BLN(BLN101),.WL(WL252));
sram_cell_6t_5 inst_cell_252_102 (.BL(BL102),.BLN(BLN102),.WL(WL252));
sram_cell_6t_5 inst_cell_252_103 (.BL(BL103),.BLN(BLN103),.WL(WL252));
sram_cell_6t_5 inst_cell_252_104 (.BL(BL104),.BLN(BLN104),.WL(WL252));
sram_cell_6t_5 inst_cell_252_105 (.BL(BL105),.BLN(BLN105),.WL(WL252));
sram_cell_6t_5 inst_cell_252_106 (.BL(BL106),.BLN(BLN106),.WL(WL252));
sram_cell_6t_5 inst_cell_252_107 (.BL(BL107),.BLN(BLN107),.WL(WL252));
sram_cell_6t_5 inst_cell_252_108 (.BL(BL108),.BLN(BLN108),.WL(WL252));
sram_cell_6t_5 inst_cell_252_109 (.BL(BL109),.BLN(BLN109),.WL(WL252));
sram_cell_6t_5 inst_cell_252_110 (.BL(BL110),.BLN(BLN110),.WL(WL252));
sram_cell_6t_5 inst_cell_252_111 (.BL(BL111),.BLN(BLN111),.WL(WL252));
sram_cell_6t_5 inst_cell_252_112 (.BL(BL112),.BLN(BLN112),.WL(WL252));
sram_cell_6t_5 inst_cell_252_113 (.BL(BL113),.BLN(BLN113),.WL(WL252));
sram_cell_6t_5 inst_cell_252_114 (.BL(BL114),.BLN(BLN114),.WL(WL252));
sram_cell_6t_5 inst_cell_252_115 (.BL(BL115),.BLN(BLN115),.WL(WL252));
sram_cell_6t_5 inst_cell_252_116 (.BL(BL116),.BLN(BLN116),.WL(WL252));
sram_cell_6t_5 inst_cell_252_117 (.BL(BL117),.BLN(BLN117),.WL(WL252));
sram_cell_6t_5 inst_cell_252_118 (.BL(BL118),.BLN(BLN118),.WL(WL252));
sram_cell_6t_5 inst_cell_252_119 (.BL(BL119),.BLN(BLN119),.WL(WL252));
sram_cell_6t_5 inst_cell_252_120 (.BL(BL120),.BLN(BLN120),.WL(WL252));
sram_cell_6t_5 inst_cell_252_121 (.BL(BL121),.BLN(BLN121),.WL(WL252));
sram_cell_6t_5 inst_cell_252_122 (.BL(BL122),.BLN(BLN122),.WL(WL252));
sram_cell_6t_5 inst_cell_252_123 (.BL(BL123),.BLN(BLN123),.WL(WL252));
sram_cell_6t_5 inst_cell_252_124 (.BL(BL124),.BLN(BLN124),.WL(WL252));
sram_cell_6t_5 inst_cell_252_125 (.BL(BL125),.BLN(BLN125),.WL(WL252));
sram_cell_6t_5 inst_cell_252_126 (.BL(BL126),.BLN(BLN126),.WL(WL252));
sram_cell_6t_5 inst_cell_252_127 (.BL(BL127),.BLN(BLN127),.WL(WL252));
sram_cell_6t_5 inst_cell_253_0 (.BL(BL0),.BLN(BLN0),.WL(WL253));
sram_cell_6t_5 inst_cell_253_1 (.BL(BL1),.BLN(BLN1),.WL(WL253));
sram_cell_6t_5 inst_cell_253_2 (.BL(BL2),.BLN(BLN2),.WL(WL253));
sram_cell_6t_5 inst_cell_253_3 (.BL(BL3),.BLN(BLN3),.WL(WL253));
sram_cell_6t_5 inst_cell_253_4 (.BL(BL4),.BLN(BLN4),.WL(WL253));
sram_cell_6t_5 inst_cell_253_5 (.BL(BL5),.BLN(BLN5),.WL(WL253));
sram_cell_6t_5 inst_cell_253_6 (.BL(BL6),.BLN(BLN6),.WL(WL253));
sram_cell_6t_5 inst_cell_253_7 (.BL(BL7),.BLN(BLN7),.WL(WL253));
sram_cell_6t_5 inst_cell_253_8 (.BL(BL8),.BLN(BLN8),.WL(WL253));
sram_cell_6t_5 inst_cell_253_9 (.BL(BL9),.BLN(BLN9),.WL(WL253));
sram_cell_6t_5 inst_cell_253_10 (.BL(BL10),.BLN(BLN10),.WL(WL253));
sram_cell_6t_5 inst_cell_253_11 (.BL(BL11),.BLN(BLN11),.WL(WL253));
sram_cell_6t_5 inst_cell_253_12 (.BL(BL12),.BLN(BLN12),.WL(WL253));
sram_cell_6t_5 inst_cell_253_13 (.BL(BL13),.BLN(BLN13),.WL(WL253));
sram_cell_6t_5 inst_cell_253_14 (.BL(BL14),.BLN(BLN14),.WL(WL253));
sram_cell_6t_5 inst_cell_253_15 (.BL(BL15),.BLN(BLN15),.WL(WL253));
sram_cell_6t_5 inst_cell_253_16 (.BL(BL16),.BLN(BLN16),.WL(WL253));
sram_cell_6t_5 inst_cell_253_17 (.BL(BL17),.BLN(BLN17),.WL(WL253));
sram_cell_6t_5 inst_cell_253_18 (.BL(BL18),.BLN(BLN18),.WL(WL253));
sram_cell_6t_5 inst_cell_253_19 (.BL(BL19),.BLN(BLN19),.WL(WL253));
sram_cell_6t_5 inst_cell_253_20 (.BL(BL20),.BLN(BLN20),.WL(WL253));
sram_cell_6t_5 inst_cell_253_21 (.BL(BL21),.BLN(BLN21),.WL(WL253));
sram_cell_6t_5 inst_cell_253_22 (.BL(BL22),.BLN(BLN22),.WL(WL253));
sram_cell_6t_5 inst_cell_253_23 (.BL(BL23),.BLN(BLN23),.WL(WL253));
sram_cell_6t_5 inst_cell_253_24 (.BL(BL24),.BLN(BLN24),.WL(WL253));
sram_cell_6t_5 inst_cell_253_25 (.BL(BL25),.BLN(BLN25),.WL(WL253));
sram_cell_6t_5 inst_cell_253_26 (.BL(BL26),.BLN(BLN26),.WL(WL253));
sram_cell_6t_5 inst_cell_253_27 (.BL(BL27),.BLN(BLN27),.WL(WL253));
sram_cell_6t_5 inst_cell_253_28 (.BL(BL28),.BLN(BLN28),.WL(WL253));
sram_cell_6t_5 inst_cell_253_29 (.BL(BL29),.BLN(BLN29),.WL(WL253));
sram_cell_6t_5 inst_cell_253_30 (.BL(BL30),.BLN(BLN30),.WL(WL253));
sram_cell_6t_5 inst_cell_253_31 (.BL(BL31),.BLN(BLN31),.WL(WL253));
sram_cell_6t_5 inst_cell_253_32 (.BL(BL32),.BLN(BLN32),.WL(WL253));
sram_cell_6t_5 inst_cell_253_33 (.BL(BL33),.BLN(BLN33),.WL(WL253));
sram_cell_6t_5 inst_cell_253_34 (.BL(BL34),.BLN(BLN34),.WL(WL253));
sram_cell_6t_5 inst_cell_253_35 (.BL(BL35),.BLN(BLN35),.WL(WL253));
sram_cell_6t_5 inst_cell_253_36 (.BL(BL36),.BLN(BLN36),.WL(WL253));
sram_cell_6t_5 inst_cell_253_37 (.BL(BL37),.BLN(BLN37),.WL(WL253));
sram_cell_6t_5 inst_cell_253_38 (.BL(BL38),.BLN(BLN38),.WL(WL253));
sram_cell_6t_5 inst_cell_253_39 (.BL(BL39),.BLN(BLN39),.WL(WL253));
sram_cell_6t_5 inst_cell_253_40 (.BL(BL40),.BLN(BLN40),.WL(WL253));
sram_cell_6t_5 inst_cell_253_41 (.BL(BL41),.BLN(BLN41),.WL(WL253));
sram_cell_6t_5 inst_cell_253_42 (.BL(BL42),.BLN(BLN42),.WL(WL253));
sram_cell_6t_5 inst_cell_253_43 (.BL(BL43),.BLN(BLN43),.WL(WL253));
sram_cell_6t_5 inst_cell_253_44 (.BL(BL44),.BLN(BLN44),.WL(WL253));
sram_cell_6t_5 inst_cell_253_45 (.BL(BL45),.BLN(BLN45),.WL(WL253));
sram_cell_6t_5 inst_cell_253_46 (.BL(BL46),.BLN(BLN46),.WL(WL253));
sram_cell_6t_5 inst_cell_253_47 (.BL(BL47),.BLN(BLN47),.WL(WL253));
sram_cell_6t_5 inst_cell_253_48 (.BL(BL48),.BLN(BLN48),.WL(WL253));
sram_cell_6t_5 inst_cell_253_49 (.BL(BL49),.BLN(BLN49),.WL(WL253));
sram_cell_6t_5 inst_cell_253_50 (.BL(BL50),.BLN(BLN50),.WL(WL253));
sram_cell_6t_5 inst_cell_253_51 (.BL(BL51),.BLN(BLN51),.WL(WL253));
sram_cell_6t_5 inst_cell_253_52 (.BL(BL52),.BLN(BLN52),.WL(WL253));
sram_cell_6t_5 inst_cell_253_53 (.BL(BL53),.BLN(BLN53),.WL(WL253));
sram_cell_6t_5 inst_cell_253_54 (.BL(BL54),.BLN(BLN54),.WL(WL253));
sram_cell_6t_5 inst_cell_253_55 (.BL(BL55),.BLN(BLN55),.WL(WL253));
sram_cell_6t_5 inst_cell_253_56 (.BL(BL56),.BLN(BLN56),.WL(WL253));
sram_cell_6t_5 inst_cell_253_57 (.BL(BL57),.BLN(BLN57),.WL(WL253));
sram_cell_6t_5 inst_cell_253_58 (.BL(BL58),.BLN(BLN58),.WL(WL253));
sram_cell_6t_5 inst_cell_253_59 (.BL(BL59),.BLN(BLN59),.WL(WL253));
sram_cell_6t_5 inst_cell_253_60 (.BL(BL60),.BLN(BLN60),.WL(WL253));
sram_cell_6t_5 inst_cell_253_61 (.BL(BL61),.BLN(BLN61),.WL(WL253));
sram_cell_6t_5 inst_cell_253_62 (.BL(BL62),.BLN(BLN62),.WL(WL253));
sram_cell_6t_5 inst_cell_253_63 (.BL(BL63),.BLN(BLN63),.WL(WL253));
sram_cell_6t_5 inst_cell_253_64 (.BL(BL64),.BLN(BLN64),.WL(WL253));
sram_cell_6t_5 inst_cell_253_65 (.BL(BL65),.BLN(BLN65),.WL(WL253));
sram_cell_6t_5 inst_cell_253_66 (.BL(BL66),.BLN(BLN66),.WL(WL253));
sram_cell_6t_5 inst_cell_253_67 (.BL(BL67),.BLN(BLN67),.WL(WL253));
sram_cell_6t_5 inst_cell_253_68 (.BL(BL68),.BLN(BLN68),.WL(WL253));
sram_cell_6t_5 inst_cell_253_69 (.BL(BL69),.BLN(BLN69),.WL(WL253));
sram_cell_6t_5 inst_cell_253_70 (.BL(BL70),.BLN(BLN70),.WL(WL253));
sram_cell_6t_5 inst_cell_253_71 (.BL(BL71),.BLN(BLN71),.WL(WL253));
sram_cell_6t_5 inst_cell_253_72 (.BL(BL72),.BLN(BLN72),.WL(WL253));
sram_cell_6t_5 inst_cell_253_73 (.BL(BL73),.BLN(BLN73),.WL(WL253));
sram_cell_6t_5 inst_cell_253_74 (.BL(BL74),.BLN(BLN74),.WL(WL253));
sram_cell_6t_5 inst_cell_253_75 (.BL(BL75),.BLN(BLN75),.WL(WL253));
sram_cell_6t_5 inst_cell_253_76 (.BL(BL76),.BLN(BLN76),.WL(WL253));
sram_cell_6t_5 inst_cell_253_77 (.BL(BL77),.BLN(BLN77),.WL(WL253));
sram_cell_6t_5 inst_cell_253_78 (.BL(BL78),.BLN(BLN78),.WL(WL253));
sram_cell_6t_5 inst_cell_253_79 (.BL(BL79),.BLN(BLN79),.WL(WL253));
sram_cell_6t_5 inst_cell_253_80 (.BL(BL80),.BLN(BLN80),.WL(WL253));
sram_cell_6t_5 inst_cell_253_81 (.BL(BL81),.BLN(BLN81),.WL(WL253));
sram_cell_6t_5 inst_cell_253_82 (.BL(BL82),.BLN(BLN82),.WL(WL253));
sram_cell_6t_5 inst_cell_253_83 (.BL(BL83),.BLN(BLN83),.WL(WL253));
sram_cell_6t_5 inst_cell_253_84 (.BL(BL84),.BLN(BLN84),.WL(WL253));
sram_cell_6t_5 inst_cell_253_85 (.BL(BL85),.BLN(BLN85),.WL(WL253));
sram_cell_6t_5 inst_cell_253_86 (.BL(BL86),.BLN(BLN86),.WL(WL253));
sram_cell_6t_5 inst_cell_253_87 (.BL(BL87),.BLN(BLN87),.WL(WL253));
sram_cell_6t_5 inst_cell_253_88 (.BL(BL88),.BLN(BLN88),.WL(WL253));
sram_cell_6t_5 inst_cell_253_89 (.BL(BL89),.BLN(BLN89),.WL(WL253));
sram_cell_6t_5 inst_cell_253_90 (.BL(BL90),.BLN(BLN90),.WL(WL253));
sram_cell_6t_5 inst_cell_253_91 (.BL(BL91),.BLN(BLN91),.WL(WL253));
sram_cell_6t_5 inst_cell_253_92 (.BL(BL92),.BLN(BLN92),.WL(WL253));
sram_cell_6t_5 inst_cell_253_93 (.BL(BL93),.BLN(BLN93),.WL(WL253));
sram_cell_6t_5 inst_cell_253_94 (.BL(BL94),.BLN(BLN94),.WL(WL253));
sram_cell_6t_5 inst_cell_253_95 (.BL(BL95),.BLN(BLN95),.WL(WL253));
sram_cell_6t_5 inst_cell_253_96 (.BL(BL96),.BLN(BLN96),.WL(WL253));
sram_cell_6t_5 inst_cell_253_97 (.BL(BL97),.BLN(BLN97),.WL(WL253));
sram_cell_6t_5 inst_cell_253_98 (.BL(BL98),.BLN(BLN98),.WL(WL253));
sram_cell_6t_5 inst_cell_253_99 (.BL(BL99),.BLN(BLN99),.WL(WL253));
sram_cell_6t_5 inst_cell_253_100 (.BL(BL100),.BLN(BLN100),.WL(WL253));
sram_cell_6t_5 inst_cell_253_101 (.BL(BL101),.BLN(BLN101),.WL(WL253));
sram_cell_6t_5 inst_cell_253_102 (.BL(BL102),.BLN(BLN102),.WL(WL253));
sram_cell_6t_5 inst_cell_253_103 (.BL(BL103),.BLN(BLN103),.WL(WL253));
sram_cell_6t_5 inst_cell_253_104 (.BL(BL104),.BLN(BLN104),.WL(WL253));
sram_cell_6t_5 inst_cell_253_105 (.BL(BL105),.BLN(BLN105),.WL(WL253));
sram_cell_6t_5 inst_cell_253_106 (.BL(BL106),.BLN(BLN106),.WL(WL253));
sram_cell_6t_5 inst_cell_253_107 (.BL(BL107),.BLN(BLN107),.WL(WL253));
sram_cell_6t_5 inst_cell_253_108 (.BL(BL108),.BLN(BLN108),.WL(WL253));
sram_cell_6t_5 inst_cell_253_109 (.BL(BL109),.BLN(BLN109),.WL(WL253));
sram_cell_6t_5 inst_cell_253_110 (.BL(BL110),.BLN(BLN110),.WL(WL253));
sram_cell_6t_5 inst_cell_253_111 (.BL(BL111),.BLN(BLN111),.WL(WL253));
sram_cell_6t_5 inst_cell_253_112 (.BL(BL112),.BLN(BLN112),.WL(WL253));
sram_cell_6t_5 inst_cell_253_113 (.BL(BL113),.BLN(BLN113),.WL(WL253));
sram_cell_6t_5 inst_cell_253_114 (.BL(BL114),.BLN(BLN114),.WL(WL253));
sram_cell_6t_5 inst_cell_253_115 (.BL(BL115),.BLN(BLN115),.WL(WL253));
sram_cell_6t_5 inst_cell_253_116 (.BL(BL116),.BLN(BLN116),.WL(WL253));
sram_cell_6t_5 inst_cell_253_117 (.BL(BL117),.BLN(BLN117),.WL(WL253));
sram_cell_6t_5 inst_cell_253_118 (.BL(BL118),.BLN(BLN118),.WL(WL253));
sram_cell_6t_5 inst_cell_253_119 (.BL(BL119),.BLN(BLN119),.WL(WL253));
sram_cell_6t_5 inst_cell_253_120 (.BL(BL120),.BLN(BLN120),.WL(WL253));
sram_cell_6t_5 inst_cell_253_121 (.BL(BL121),.BLN(BLN121),.WL(WL253));
sram_cell_6t_5 inst_cell_253_122 (.BL(BL122),.BLN(BLN122),.WL(WL253));
sram_cell_6t_5 inst_cell_253_123 (.BL(BL123),.BLN(BLN123),.WL(WL253));
sram_cell_6t_5 inst_cell_253_124 (.BL(BL124),.BLN(BLN124),.WL(WL253));
sram_cell_6t_5 inst_cell_253_125 (.BL(BL125),.BLN(BLN125),.WL(WL253));
sram_cell_6t_5 inst_cell_253_126 (.BL(BL126),.BLN(BLN126),.WL(WL253));
sram_cell_6t_5 inst_cell_253_127 (.BL(BL127),.BLN(BLN127),.WL(WL253));
sram_cell_6t_5 inst_cell_254_0 (.BL(BL0),.BLN(BLN0),.WL(WL254));
sram_cell_6t_5 inst_cell_254_1 (.BL(BL1),.BLN(BLN1),.WL(WL254));
sram_cell_6t_5 inst_cell_254_2 (.BL(BL2),.BLN(BLN2),.WL(WL254));
sram_cell_6t_5 inst_cell_254_3 (.BL(BL3),.BLN(BLN3),.WL(WL254));
sram_cell_6t_5 inst_cell_254_4 (.BL(BL4),.BLN(BLN4),.WL(WL254));
sram_cell_6t_5 inst_cell_254_5 (.BL(BL5),.BLN(BLN5),.WL(WL254));
sram_cell_6t_5 inst_cell_254_6 (.BL(BL6),.BLN(BLN6),.WL(WL254));
sram_cell_6t_5 inst_cell_254_7 (.BL(BL7),.BLN(BLN7),.WL(WL254));
sram_cell_6t_5 inst_cell_254_8 (.BL(BL8),.BLN(BLN8),.WL(WL254));
sram_cell_6t_5 inst_cell_254_9 (.BL(BL9),.BLN(BLN9),.WL(WL254));
sram_cell_6t_5 inst_cell_254_10 (.BL(BL10),.BLN(BLN10),.WL(WL254));
sram_cell_6t_5 inst_cell_254_11 (.BL(BL11),.BLN(BLN11),.WL(WL254));
sram_cell_6t_5 inst_cell_254_12 (.BL(BL12),.BLN(BLN12),.WL(WL254));
sram_cell_6t_5 inst_cell_254_13 (.BL(BL13),.BLN(BLN13),.WL(WL254));
sram_cell_6t_5 inst_cell_254_14 (.BL(BL14),.BLN(BLN14),.WL(WL254));
sram_cell_6t_5 inst_cell_254_15 (.BL(BL15),.BLN(BLN15),.WL(WL254));
sram_cell_6t_5 inst_cell_254_16 (.BL(BL16),.BLN(BLN16),.WL(WL254));
sram_cell_6t_5 inst_cell_254_17 (.BL(BL17),.BLN(BLN17),.WL(WL254));
sram_cell_6t_5 inst_cell_254_18 (.BL(BL18),.BLN(BLN18),.WL(WL254));
sram_cell_6t_5 inst_cell_254_19 (.BL(BL19),.BLN(BLN19),.WL(WL254));
sram_cell_6t_5 inst_cell_254_20 (.BL(BL20),.BLN(BLN20),.WL(WL254));
sram_cell_6t_5 inst_cell_254_21 (.BL(BL21),.BLN(BLN21),.WL(WL254));
sram_cell_6t_5 inst_cell_254_22 (.BL(BL22),.BLN(BLN22),.WL(WL254));
sram_cell_6t_5 inst_cell_254_23 (.BL(BL23),.BLN(BLN23),.WL(WL254));
sram_cell_6t_5 inst_cell_254_24 (.BL(BL24),.BLN(BLN24),.WL(WL254));
sram_cell_6t_5 inst_cell_254_25 (.BL(BL25),.BLN(BLN25),.WL(WL254));
sram_cell_6t_5 inst_cell_254_26 (.BL(BL26),.BLN(BLN26),.WL(WL254));
sram_cell_6t_5 inst_cell_254_27 (.BL(BL27),.BLN(BLN27),.WL(WL254));
sram_cell_6t_5 inst_cell_254_28 (.BL(BL28),.BLN(BLN28),.WL(WL254));
sram_cell_6t_5 inst_cell_254_29 (.BL(BL29),.BLN(BLN29),.WL(WL254));
sram_cell_6t_5 inst_cell_254_30 (.BL(BL30),.BLN(BLN30),.WL(WL254));
sram_cell_6t_5 inst_cell_254_31 (.BL(BL31),.BLN(BLN31),.WL(WL254));
sram_cell_6t_5 inst_cell_254_32 (.BL(BL32),.BLN(BLN32),.WL(WL254));
sram_cell_6t_5 inst_cell_254_33 (.BL(BL33),.BLN(BLN33),.WL(WL254));
sram_cell_6t_5 inst_cell_254_34 (.BL(BL34),.BLN(BLN34),.WL(WL254));
sram_cell_6t_5 inst_cell_254_35 (.BL(BL35),.BLN(BLN35),.WL(WL254));
sram_cell_6t_5 inst_cell_254_36 (.BL(BL36),.BLN(BLN36),.WL(WL254));
sram_cell_6t_5 inst_cell_254_37 (.BL(BL37),.BLN(BLN37),.WL(WL254));
sram_cell_6t_5 inst_cell_254_38 (.BL(BL38),.BLN(BLN38),.WL(WL254));
sram_cell_6t_5 inst_cell_254_39 (.BL(BL39),.BLN(BLN39),.WL(WL254));
sram_cell_6t_5 inst_cell_254_40 (.BL(BL40),.BLN(BLN40),.WL(WL254));
sram_cell_6t_5 inst_cell_254_41 (.BL(BL41),.BLN(BLN41),.WL(WL254));
sram_cell_6t_5 inst_cell_254_42 (.BL(BL42),.BLN(BLN42),.WL(WL254));
sram_cell_6t_5 inst_cell_254_43 (.BL(BL43),.BLN(BLN43),.WL(WL254));
sram_cell_6t_5 inst_cell_254_44 (.BL(BL44),.BLN(BLN44),.WL(WL254));
sram_cell_6t_5 inst_cell_254_45 (.BL(BL45),.BLN(BLN45),.WL(WL254));
sram_cell_6t_5 inst_cell_254_46 (.BL(BL46),.BLN(BLN46),.WL(WL254));
sram_cell_6t_5 inst_cell_254_47 (.BL(BL47),.BLN(BLN47),.WL(WL254));
sram_cell_6t_5 inst_cell_254_48 (.BL(BL48),.BLN(BLN48),.WL(WL254));
sram_cell_6t_5 inst_cell_254_49 (.BL(BL49),.BLN(BLN49),.WL(WL254));
sram_cell_6t_5 inst_cell_254_50 (.BL(BL50),.BLN(BLN50),.WL(WL254));
sram_cell_6t_5 inst_cell_254_51 (.BL(BL51),.BLN(BLN51),.WL(WL254));
sram_cell_6t_5 inst_cell_254_52 (.BL(BL52),.BLN(BLN52),.WL(WL254));
sram_cell_6t_5 inst_cell_254_53 (.BL(BL53),.BLN(BLN53),.WL(WL254));
sram_cell_6t_5 inst_cell_254_54 (.BL(BL54),.BLN(BLN54),.WL(WL254));
sram_cell_6t_5 inst_cell_254_55 (.BL(BL55),.BLN(BLN55),.WL(WL254));
sram_cell_6t_5 inst_cell_254_56 (.BL(BL56),.BLN(BLN56),.WL(WL254));
sram_cell_6t_5 inst_cell_254_57 (.BL(BL57),.BLN(BLN57),.WL(WL254));
sram_cell_6t_5 inst_cell_254_58 (.BL(BL58),.BLN(BLN58),.WL(WL254));
sram_cell_6t_5 inst_cell_254_59 (.BL(BL59),.BLN(BLN59),.WL(WL254));
sram_cell_6t_5 inst_cell_254_60 (.BL(BL60),.BLN(BLN60),.WL(WL254));
sram_cell_6t_5 inst_cell_254_61 (.BL(BL61),.BLN(BLN61),.WL(WL254));
sram_cell_6t_5 inst_cell_254_62 (.BL(BL62),.BLN(BLN62),.WL(WL254));
sram_cell_6t_5 inst_cell_254_63 (.BL(BL63),.BLN(BLN63),.WL(WL254));
sram_cell_6t_5 inst_cell_254_64 (.BL(BL64),.BLN(BLN64),.WL(WL254));
sram_cell_6t_5 inst_cell_254_65 (.BL(BL65),.BLN(BLN65),.WL(WL254));
sram_cell_6t_5 inst_cell_254_66 (.BL(BL66),.BLN(BLN66),.WL(WL254));
sram_cell_6t_5 inst_cell_254_67 (.BL(BL67),.BLN(BLN67),.WL(WL254));
sram_cell_6t_5 inst_cell_254_68 (.BL(BL68),.BLN(BLN68),.WL(WL254));
sram_cell_6t_5 inst_cell_254_69 (.BL(BL69),.BLN(BLN69),.WL(WL254));
sram_cell_6t_5 inst_cell_254_70 (.BL(BL70),.BLN(BLN70),.WL(WL254));
sram_cell_6t_5 inst_cell_254_71 (.BL(BL71),.BLN(BLN71),.WL(WL254));
sram_cell_6t_5 inst_cell_254_72 (.BL(BL72),.BLN(BLN72),.WL(WL254));
sram_cell_6t_5 inst_cell_254_73 (.BL(BL73),.BLN(BLN73),.WL(WL254));
sram_cell_6t_5 inst_cell_254_74 (.BL(BL74),.BLN(BLN74),.WL(WL254));
sram_cell_6t_5 inst_cell_254_75 (.BL(BL75),.BLN(BLN75),.WL(WL254));
sram_cell_6t_5 inst_cell_254_76 (.BL(BL76),.BLN(BLN76),.WL(WL254));
sram_cell_6t_5 inst_cell_254_77 (.BL(BL77),.BLN(BLN77),.WL(WL254));
sram_cell_6t_5 inst_cell_254_78 (.BL(BL78),.BLN(BLN78),.WL(WL254));
sram_cell_6t_5 inst_cell_254_79 (.BL(BL79),.BLN(BLN79),.WL(WL254));
sram_cell_6t_5 inst_cell_254_80 (.BL(BL80),.BLN(BLN80),.WL(WL254));
sram_cell_6t_5 inst_cell_254_81 (.BL(BL81),.BLN(BLN81),.WL(WL254));
sram_cell_6t_5 inst_cell_254_82 (.BL(BL82),.BLN(BLN82),.WL(WL254));
sram_cell_6t_5 inst_cell_254_83 (.BL(BL83),.BLN(BLN83),.WL(WL254));
sram_cell_6t_5 inst_cell_254_84 (.BL(BL84),.BLN(BLN84),.WL(WL254));
sram_cell_6t_5 inst_cell_254_85 (.BL(BL85),.BLN(BLN85),.WL(WL254));
sram_cell_6t_5 inst_cell_254_86 (.BL(BL86),.BLN(BLN86),.WL(WL254));
sram_cell_6t_5 inst_cell_254_87 (.BL(BL87),.BLN(BLN87),.WL(WL254));
sram_cell_6t_5 inst_cell_254_88 (.BL(BL88),.BLN(BLN88),.WL(WL254));
sram_cell_6t_5 inst_cell_254_89 (.BL(BL89),.BLN(BLN89),.WL(WL254));
sram_cell_6t_5 inst_cell_254_90 (.BL(BL90),.BLN(BLN90),.WL(WL254));
sram_cell_6t_5 inst_cell_254_91 (.BL(BL91),.BLN(BLN91),.WL(WL254));
sram_cell_6t_5 inst_cell_254_92 (.BL(BL92),.BLN(BLN92),.WL(WL254));
sram_cell_6t_5 inst_cell_254_93 (.BL(BL93),.BLN(BLN93),.WL(WL254));
sram_cell_6t_5 inst_cell_254_94 (.BL(BL94),.BLN(BLN94),.WL(WL254));
sram_cell_6t_5 inst_cell_254_95 (.BL(BL95),.BLN(BLN95),.WL(WL254));
sram_cell_6t_5 inst_cell_254_96 (.BL(BL96),.BLN(BLN96),.WL(WL254));
sram_cell_6t_5 inst_cell_254_97 (.BL(BL97),.BLN(BLN97),.WL(WL254));
sram_cell_6t_5 inst_cell_254_98 (.BL(BL98),.BLN(BLN98),.WL(WL254));
sram_cell_6t_5 inst_cell_254_99 (.BL(BL99),.BLN(BLN99),.WL(WL254));
sram_cell_6t_5 inst_cell_254_100 (.BL(BL100),.BLN(BLN100),.WL(WL254));
sram_cell_6t_5 inst_cell_254_101 (.BL(BL101),.BLN(BLN101),.WL(WL254));
sram_cell_6t_5 inst_cell_254_102 (.BL(BL102),.BLN(BLN102),.WL(WL254));
sram_cell_6t_5 inst_cell_254_103 (.BL(BL103),.BLN(BLN103),.WL(WL254));
sram_cell_6t_5 inst_cell_254_104 (.BL(BL104),.BLN(BLN104),.WL(WL254));
sram_cell_6t_5 inst_cell_254_105 (.BL(BL105),.BLN(BLN105),.WL(WL254));
sram_cell_6t_5 inst_cell_254_106 (.BL(BL106),.BLN(BLN106),.WL(WL254));
sram_cell_6t_5 inst_cell_254_107 (.BL(BL107),.BLN(BLN107),.WL(WL254));
sram_cell_6t_5 inst_cell_254_108 (.BL(BL108),.BLN(BLN108),.WL(WL254));
sram_cell_6t_5 inst_cell_254_109 (.BL(BL109),.BLN(BLN109),.WL(WL254));
sram_cell_6t_5 inst_cell_254_110 (.BL(BL110),.BLN(BLN110),.WL(WL254));
sram_cell_6t_5 inst_cell_254_111 (.BL(BL111),.BLN(BLN111),.WL(WL254));
sram_cell_6t_5 inst_cell_254_112 (.BL(BL112),.BLN(BLN112),.WL(WL254));
sram_cell_6t_5 inst_cell_254_113 (.BL(BL113),.BLN(BLN113),.WL(WL254));
sram_cell_6t_5 inst_cell_254_114 (.BL(BL114),.BLN(BLN114),.WL(WL254));
sram_cell_6t_5 inst_cell_254_115 (.BL(BL115),.BLN(BLN115),.WL(WL254));
sram_cell_6t_5 inst_cell_254_116 (.BL(BL116),.BLN(BLN116),.WL(WL254));
sram_cell_6t_5 inst_cell_254_117 (.BL(BL117),.BLN(BLN117),.WL(WL254));
sram_cell_6t_5 inst_cell_254_118 (.BL(BL118),.BLN(BLN118),.WL(WL254));
sram_cell_6t_5 inst_cell_254_119 (.BL(BL119),.BLN(BLN119),.WL(WL254));
sram_cell_6t_5 inst_cell_254_120 (.BL(BL120),.BLN(BLN120),.WL(WL254));
sram_cell_6t_5 inst_cell_254_121 (.BL(BL121),.BLN(BLN121),.WL(WL254));
sram_cell_6t_5 inst_cell_254_122 (.BL(BL122),.BLN(BLN122),.WL(WL254));
sram_cell_6t_5 inst_cell_254_123 (.BL(BL123),.BLN(BLN123),.WL(WL254));
sram_cell_6t_5 inst_cell_254_124 (.BL(BL124),.BLN(BLN124),.WL(WL254));
sram_cell_6t_5 inst_cell_254_125 (.BL(BL125),.BLN(BLN125),.WL(WL254));
sram_cell_6t_5 inst_cell_254_126 (.BL(BL126),.BLN(BLN126),.WL(WL254));
sram_cell_6t_5 inst_cell_254_127 (.BL(BL127),.BLN(BLN127),.WL(WL254));
sram_cell_6t_5 inst_cell_255_0 (.BL(BL0),.BLN(BLN0),.WL(WL255));
sram_cell_6t_5 inst_cell_255_1 (.BL(BL1),.BLN(BLN1),.WL(WL255));
sram_cell_6t_5 inst_cell_255_2 (.BL(BL2),.BLN(BLN2),.WL(WL255));
sram_cell_6t_5 inst_cell_255_3 (.BL(BL3),.BLN(BLN3),.WL(WL255));
sram_cell_6t_5 inst_cell_255_4 (.BL(BL4),.BLN(BLN4),.WL(WL255));
sram_cell_6t_5 inst_cell_255_5 (.BL(BL5),.BLN(BLN5),.WL(WL255));
sram_cell_6t_5 inst_cell_255_6 (.BL(BL6),.BLN(BLN6),.WL(WL255));
sram_cell_6t_5 inst_cell_255_7 (.BL(BL7),.BLN(BLN7),.WL(WL255));
sram_cell_6t_5 inst_cell_255_8 (.BL(BL8),.BLN(BLN8),.WL(WL255));
sram_cell_6t_5 inst_cell_255_9 (.BL(BL9),.BLN(BLN9),.WL(WL255));
sram_cell_6t_5 inst_cell_255_10 (.BL(BL10),.BLN(BLN10),.WL(WL255));
sram_cell_6t_5 inst_cell_255_11 (.BL(BL11),.BLN(BLN11),.WL(WL255));
sram_cell_6t_5 inst_cell_255_12 (.BL(BL12),.BLN(BLN12),.WL(WL255));
sram_cell_6t_5 inst_cell_255_13 (.BL(BL13),.BLN(BLN13),.WL(WL255));
sram_cell_6t_5 inst_cell_255_14 (.BL(BL14),.BLN(BLN14),.WL(WL255));
sram_cell_6t_5 inst_cell_255_15 (.BL(BL15),.BLN(BLN15),.WL(WL255));
sram_cell_6t_5 inst_cell_255_16 (.BL(BL16),.BLN(BLN16),.WL(WL255));
sram_cell_6t_5 inst_cell_255_17 (.BL(BL17),.BLN(BLN17),.WL(WL255));
sram_cell_6t_5 inst_cell_255_18 (.BL(BL18),.BLN(BLN18),.WL(WL255));
sram_cell_6t_5 inst_cell_255_19 (.BL(BL19),.BLN(BLN19),.WL(WL255));
sram_cell_6t_5 inst_cell_255_20 (.BL(BL20),.BLN(BLN20),.WL(WL255));
sram_cell_6t_5 inst_cell_255_21 (.BL(BL21),.BLN(BLN21),.WL(WL255));
sram_cell_6t_5 inst_cell_255_22 (.BL(BL22),.BLN(BLN22),.WL(WL255));
sram_cell_6t_5 inst_cell_255_23 (.BL(BL23),.BLN(BLN23),.WL(WL255));
sram_cell_6t_5 inst_cell_255_24 (.BL(BL24),.BLN(BLN24),.WL(WL255));
sram_cell_6t_5 inst_cell_255_25 (.BL(BL25),.BLN(BLN25),.WL(WL255));
sram_cell_6t_5 inst_cell_255_26 (.BL(BL26),.BLN(BLN26),.WL(WL255));
sram_cell_6t_5 inst_cell_255_27 (.BL(BL27),.BLN(BLN27),.WL(WL255));
sram_cell_6t_5 inst_cell_255_28 (.BL(BL28),.BLN(BLN28),.WL(WL255));
sram_cell_6t_5 inst_cell_255_29 (.BL(BL29),.BLN(BLN29),.WL(WL255));
sram_cell_6t_5 inst_cell_255_30 (.BL(BL30),.BLN(BLN30),.WL(WL255));
sram_cell_6t_5 inst_cell_255_31 (.BL(BL31),.BLN(BLN31),.WL(WL255));
sram_cell_6t_5 inst_cell_255_32 (.BL(BL32),.BLN(BLN32),.WL(WL255));
sram_cell_6t_5 inst_cell_255_33 (.BL(BL33),.BLN(BLN33),.WL(WL255));
sram_cell_6t_5 inst_cell_255_34 (.BL(BL34),.BLN(BLN34),.WL(WL255));
sram_cell_6t_5 inst_cell_255_35 (.BL(BL35),.BLN(BLN35),.WL(WL255));
sram_cell_6t_5 inst_cell_255_36 (.BL(BL36),.BLN(BLN36),.WL(WL255));
sram_cell_6t_5 inst_cell_255_37 (.BL(BL37),.BLN(BLN37),.WL(WL255));
sram_cell_6t_5 inst_cell_255_38 (.BL(BL38),.BLN(BLN38),.WL(WL255));
sram_cell_6t_5 inst_cell_255_39 (.BL(BL39),.BLN(BLN39),.WL(WL255));
sram_cell_6t_5 inst_cell_255_40 (.BL(BL40),.BLN(BLN40),.WL(WL255));
sram_cell_6t_5 inst_cell_255_41 (.BL(BL41),.BLN(BLN41),.WL(WL255));
sram_cell_6t_5 inst_cell_255_42 (.BL(BL42),.BLN(BLN42),.WL(WL255));
sram_cell_6t_5 inst_cell_255_43 (.BL(BL43),.BLN(BLN43),.WL(WL255));
sram_cell_6t_5 inst_cell_255_44 (.BL(BL44),.BLN(BLN44),.WL(WL255));
sram_cell_6t_5 inst_cell_255_45 (.BL(BL45),.BLN(BLN45),.WL(WL255));
sram_cell_6t_5 inst_cell_255_46 (.BL(BL46),.BLN(BLN46),.WL(WL255));
sram_cell_6t_5 inst_cell_255_47 (.BL(BL47),.BLN(BLN47),.WL(WL255));
sram_cell_6t_5 inst_cell_255_48 (.BL(BL48),.BLN(BLN48),.WL(WL255));
sram_cell_6t_5 inst_cell_255_49 (.BL(BL49),.BLN(BLN49),.WL(WL255));
sram_cell_6t_5 inst_cell_255_50 (.BL(BL50),.BLN(BLN50),.WL(WL255));
sram_cell_6t_5 inst_cell_255_51 (.BL(BL51),.BLN(BLN51),.WL(WL255));
sram_cell_6t_5 inst_cell_255_52 (.BL(BL52),.BLN(BLN52),.WL(WL255));
sram_cell_6t_5 inst_cell_255_53 (.BL(BL53),.BLN(BLN53),.WL(WL255));
sram_cell_6t_5 inst_cell_255_54 (.BL(BL54),.BLN(BLN54),.WL(WL255));
sram_cell_6t_5 inst_cell_255_55 (.BL(BL55),.BLN(BLN55),.WL(WL255));
sram_cell_6t_5 inst_cell_255_56 (.BL(BL56),.BLN(BLN56),.WL(WL255));
sram_cell_6t_5 inst_cell_255_57 (.BL(BL57),.BLN(BLN57),.WL(WL255));
sram_cell_6t_5 inst_cell_255_58 (.BL(BL58),.BLN(BLN58),.WL(WL255));
sram_cell_6t_5 inst_cell_255_59 (.BL(BL59),.BLN(BLN59),.WL(WL255));
sram_cell_6t_5 inst_cell_255_60 (.BL(BL60),.BLN(BLN60),.WL(WL255));
sram_cell_6t_5 inst_cell_255_61 (.BL(BL61),.BLN(BLN61),.WL(WL255));
sram_cell_6t_5 inst_cell_255_62 (.BL(BL62),.BLN(BLN62),.WL(WL255));
sram_cell_6t_5 inst_cell_255_63 (.BL(BL63),.BLN(BLN63),.WL(WL255));
sram_cell_6t_5 inst_cell_255_64 (.BL(BL64),.BLN(BLN64),.WL(WL255));
sram_cell_6t_5 inst_cell_255_65 (.BL(BL65),.BLN(BLN65),.WL(WL255));
sram_cell_6t_5 inst_cell_255_66 (.BL(BL66),.BLN(BLN66),.WL(WL255));
sram_cell_6t_5 inst_cell_255_67 (.BL(BL67),.BLN(BLN67),.WL(WL255));
sram_cell_6t_5 inst_cell_255_68 (.BL(BL68),.BLN(BLN68),.WL(WL255));
sram_cell_6t_5 inst_cell_255_69 (.BL(BL69),.BLN(BLN69),.WL(WL255));
sram_cell_6t_5 inst_cell_255_70 (.BL(BL70),.BLN(BLN70),.WL(WL255));
sram_cell_6t_5 inst_cell_255_71 (.BL(BL71),.BLN(BLN71),.WL(WL255));
sram_cell_6t_5 inst_cell_255_72 (.BL(BL72),.BLN(BLN72),.WL(WL255));
sram_cell_6t_5 inst_cell_255_73 (.BL(BL73),.BLN(BLN73),.WL(WL255));
sram_cell_6t_5 inst_cell_255_74 (.BL(BL74),.BLN(BLN74),.WL(WL255));
sram_cell_6t_5 inst_cell_255_75 (.BL(BL75),.BLN(BLN75),.WL(WL255));
sram_cell_6t_5 inst_cell_255_76 (.BL(BL76),.BLN(BLN76),.WL(WL255));
sram_cell_6t_5 inst_cell_255_77 (.BL(BL77),.BLN(BLN77),.WL(WL255));
sram_cell_6t_5 inst_cell_255_78 (.BL(BL78),.BLN(BLN78),.WL(WL255));
sram_cell_6t_5 inst_cell_255_79 (.BL(BL79),.BLN(BLN79),.WL(WL255));
sram_cell_6t_5 inst_cell_255_80 (.BL(BL80),.BLN(BLN80),.WL(WL255));
sram_cell_6t_5 inst_cell_255_81 (.BL(BL81),.BLN(BLN81),.WL(WL255));
sram_cell_6t_5 inst_cell_255_82 (.BL(BL82),.BLN(BLN82),.WL(WL255));
sram_cell_6t_5 inst_cell_255_83 (.BL(BL83),.BLN(BLN83),.WL(WL255));
sram_cell_6t_5 inst_cell_255_84 (.BL(BL84),.BLN(BLN84),.WL(WL255));
sram_cell_6t_5 inst_cell_255_85 (.BL(BL85),.BLN(BLN85),.WL(WL255));
sram_cell_6t_5 inst_cell_255_86 (.BL(BL86),.BLN(BLN86),.WL(WL255));
sram_cell_6t_5 inst_cell_255_87 (.BL(BL87),.BLN(BLN87),.WL(WL255));
sram_cell_6t_5 inst_cell_255_88 (.BL(BL88),.BLN(BLN88),.WL(WL255));
sram_cell_6t_5 inst_cell_255_89 (.BL(BL89),.BLN(BLN89),.WL(WL255));
sram_cell_6t_5 inst_cell_255_90 (.BL(BL90),.BLN(BLN90),.WL(WL255));
sram_cell_6t_5 inst_cell_255_91 (.BL(BL91),.BLN(BLN91),.WL(WL255));
sram_cell_6t_5 inst_cell_255_92 (.BL(BL92),.BLN(BLN92),.WL(WL255));
sram_cell_6t_5 inst_cell_255_93 (.BL(BL93),.BLN(BLN93),.WL(WL255));
sram_cell_6t_5 inst_cell_255_94 (.BL(BL94),.BLN(BLN94),.WL(WL255));
sram_cell_6t_5 inst_cell_255_95 (.BL(BL95),.BLN(BLN95),.WL(WL255));
sram_cell_6t_5 inst_cell_255_96 (.BL(BL96),.BLN(BLN96),.WL(WL255));
sram_cell_6t_5 inst_cell_255_97 (.BL(BL97),.BLN(BLN97),.WL(WL255));
sram_cell_6t_5 inst_cell_255_98 (.BL(BL98),.BLN(BLN98),.WL(WL255));
sram_cell_6t_5 inst_cell_255_99 (.BL(BL99),.BLN(BLN99),.WL(WL255));
sram_cell_6t_5 inst_cell_255_100 (.BL(BL100),.BLN(BLN100),.WL(WL255));
sram_cell_6t_5 inst_cell_255_101 (.BL(BL101),.BLN(BLN101),.WL(WL255));
sram_cell_6t_5 inst_cell_255_102 (.BL(BL102),.BLN(BLN102),.WL(WL255));
sram_cell_6t_5 inst_cell_255_103 (.BL(BL103),.BLN(BLN103),.WL(WL255));
sram_cell_6t_5 inst_cell_255_104 (.BL(BL104),.BLN(BLN104),.WL(WL255));
sram_cell_6t_5 inst_cell_255_105 (.BL(BL105),.BLN(BLN105),.WL(WL255));
sram_cell_6t_5 inst_cell_255_106 (.BL(BL106),.BLN(BLN106),.WL(WL255));
sram_cell_6t_5 inst_cell_255_107 (.BL(BL107),.BLN(BLN107),.WL(WL255));
sram_cell_6t_5 inst_cell_255_108 (.BL(BL108),.BLN(BLN108),.WL(WL255));
sram_cell_6t_5 inst_cell_255_109 (.BL(BL109),.BLN(BLN109),.WL(WL255));
sram_cell_6t_5 inst_cell_255_110 (.BL(BL110),.BLN(BLN110),.WL(WL255));
sram_cell_6t_5 inst_cell_255_111 (.BL(BL111),.BLN(BLN111),.WL(WL255));
sram_cell_6t_5 inst_cell_255_112 (.BL(BL112),.BLN(BLN112),.WL(WL255));
sram_cell_6t_5 inst_cell_255_113 (.BL(BL113),.BLN(BLN113),.WL(WL255));
sram_cell_6t_5 inst_cell_255_114 (.BL(BL114),.BLN(BLN114),.WL(WL255));
sram_cell_6t_5 inst_cell_255_115 (.BL(BL115),.BLN(BLN115),.WL(WL255));
sram_cell_6t_5 inst_cell_255_116 (.BL(BL116),.BLN(BLN116),.WL(WL255));
sram_cell_6t_5 inst_cell_255_117 (.BL(BL117),.BLN(BLN117),.WL(WL255));
sram_cell_6t_5 inst_cell_255_118 (.BL(BL118),.BLN(BLN118),.WL(WL255));
sram_cell_6t_5 inst_cell_255_119 (.BL(BL119),.BLN(BLN119),.WL(WL255));
sram_cell_6t_5 inst_cell_255_120 (.BL(BL120),.BLN(BLN120),.WL(WL255));
sram_cell_6t_5 inst_cell_255_121 (.BL(BL121),.BLN(BLN121),.WL(WL255));
sram_cell_6t_5 inst_cell_255_122 (.BL(BL122),.BLN(BLN122),.WL(WL255));
sram_cell_6t_5 inst_cell_255_123 (.BL(BL123),.BLN(BLN123),.WL(WL255));
sram_cell_6t_5 inst_cell_255_124 (.BL(BL124),.BLN(BLN124),.WL(WL255));
sram_cell_6t_5 inst_cell_255_125 (.BL(BL125),.BLN(BLN125),.WL(WL255));
sram_cell_6t_5 inst_cell_255_126 (.BL(BL126),.BLN(BLN126),.WL(WL255));
sram_cell_6t_5 inst_cell_255_127 (.BL(BL127),.BLN(BLN127),.WL(WL255));
columnMux inst_colMux0 (BL0,BLN0,BL1,BLN1,BL2,BLN2,BL3,BLN3,BL4,BLN4,BL5,BLN5,BL6,BLN6,BL7,BLN7,BL8,BLN8,BL9,BLN9,BL10,BLN10,BL11,BLN11,BL12,BLN12,BL13,BLN13,BL14,BLN14,BL15,BLN15,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL0,DLN0);
write_driver_compiler inst_writeDriver0 (.clk(clk_bar),.data(din0),.write_en(write_en),.BL(DL0),.BLN(DLN0));
sense_amp_clocked_compiler inst_senAmp0 (.bit(DL0),.bit_bar(DLN0),.sense_en(sense_en),.sense(dout0));
columnMux inst_colMux1 (BL16,BLN16,BL17,BLN17,BL18,BLN18,BL19,BLN19,BL20,BLN20,BL21,BLN21,BL22,BLN22,BL23,BLN23,BL24,BLN24,BL25,BLN25,BL26,BLN26,BL27,BLN27,BL28,BLN28,BL29,BLN29,BL30,BLN30,BL31,BLN31,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL1,DLN1);
write_driver_compiler inst_writeDriver1 (.clk(clk_bar),.data(din1),.write_en(write_en),.BL(DL1),.BLN(DLN1));
sense_amp_clocked_compiler inst_senAmp1 (.bit(DL1),.bit_bar(DLN1),.sense_en(sense_en),.sense(dout1));
columnMux inst_colMux2 (BL32,BLN32,BL33,BLN33,BL34,BLN34,BL35,BLN35,BL36,BLN36,BL37,BLN37,BL38,BLN38,BL39,BLN39,BL40,BLN40,BL41,BLN41,BL42,BLN42,BL43,BLN43,BL44,BLN44,BL45,BLN45,BL46,BLN46,BL47,BLN47,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL2,DLN2);
write_driver_compiler inst_writeDriver2 (.clk(clk_bar),.data(din2),.write_en(write_en),.BL(DL2),.BLN(DLN2));
sense_amp_clocked_compiler inst_senAmp2 (.bit(DL2),.bit_bar(DLN2),.sense_en(sense_en),.sense(dout2));
columnMux inst_colMux3 (BL48,BLN48,BL49,BLN49,BL50,BLN50,BL51,BLN51,BL52,BLN52,BL53,BLN53,BL54,BLN54,BL55,BLN55,BL56,BLN56,BL57,BLN57,BL58,BLN58,BL59,BLN59,BL60,BLN60,BL61,BLN61,BL62,BLN62,BL63,BLN63,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL3,DLN3);
write_driver_compiler inst_writeDriver3 (.clk(clk_bar),.data(din3),.write_en(write_en),.BL(DL3),.BLN(DLN3));
sense_amp_clocked_compiler inst_senAmp3 (.bit(DL3),.bit_bar(DLN3),.sense_en(sense_en),.sense(dout3));
columnMux inst_colMux4 (BL64,BLN64,BL65,BLN65,BL66,BLN66,BL67,BLN67,BL68,BLN68,BL69,BLN69,BL70,BLN70,BL71,BLN71,BL72,BLN72,BL73,BLN73,BL74,BLN74,BL75,BLN75,BL76,BLN76,BL77,BLN77,BL78,BLN78,BL79,BLN79,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL4,DLN4);
write_driver_compiler inst_writeDriver4 (.clk(clk_bar),.data(din4),.write_en(write_en),.BL(DL4),.BLN(DLN4));
sense_amp_clocked_compiler inst_senAmp4 (.bit(DL4),.bit_bar(DLN4),.sense_en(sense_en),.sense(dout4));
columnMux inst_colMux5 (BL80,BLN80,BL81,BLN81,BL82,BLN82,BL83,BLN83,BL84,BLN84,BL85,BLN85,BL86,BLN86,BL87,BLN87,BL88,BLN88,BL89,BLN89,BL90,BLN90,BL91,BLN91,BL92,BLN92,BL93,BLN93,BL94,BLN94,BL95,BLN95,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL5,DLN5);
write_driver_compiler inst_writeDriver5 (.clk(clk_bar),.data(din5),.write_en(write_en),.BL(DL5),.BLN(DLN5));
sense_amp_clocked_compiler inst_senAmp5 (.bit(DL5),.bit_bar(DLN5),.sense_en(sense_en),.sense(dout5));
columnMux inst_colMux6 (BL96,BLN96,BL97,BLN97,BL98,BLN98,BL99,BLN99,BL100,BLN100,BL101,BLN101,BL102,BLN102,BL103,BLN103,BL104,BLN104,BL105,BLN105,BL106,BLN106,BL107,BLN107,BL108,BLN108,BL109,BLN109,BL110,BLN110,BL111,BLN111,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL6,DLN6);
write_driver_compiler inst_writeDriver6 (.clk(clk_bar),.data(din6),.write_en(write_en),.BL(DL6),.BLN(DLN6));
sense_amp_clocked_compiler inst_senAmp6 (.bit(DL6),.bit_bar(DLN6),.sense_en(sense_en),.sense(dout6));
columnMux inst_colMux7 (BL112,BLN112,BL113,BLN113,BL114,BLN114,BL115,BLN115,BL116,BLN116,BL117,BLN117,BL118,BLN118,BL119,BLN119,BL120,BLN120,BL121,BLN121,BL122,BLN122,BL123,BLN123,BL124,BLN124,BL125,BLN125,BL126,BLN126,BL127,BLN127,SL0,SL1,SL2,SL3,SL4,SL5,SL6,SL7,SL8,SL9,SL10,SL11,SL12,SL13,SL14,SL15,DL7,DLN7);
write_driver_compiler inst_writeDriver7 (.clk(clk_bar),.data(din7),.write_en(write_en),.BL(DL7),.BLN(DLN7));
sense_amp_clocked_compiler inst_senAmp7 (.bit(DL7),.bit_bar(DLN7),.sense_en(sense_en),.sense(dout7));
precharge_compiler inst_precharge0 (.clk(clk_bar),.B(BL0),.B_bar(BLN0));
precharge_compiler inst_precharge1 (.clk(clk_bar),.B(BL1),.B_bar(BLN1));
precharge_compiler inst_precharge2 (.clk(clk_bar),.B(BL2),.B_bar(BLN2));
precharge_compiler inst_precharge3 (.clk(clk_bar),.B(BL3),.B_bar(BLN3));
precharge_compiler inst_precharge4 (.clk(clk_bar),.B(BL4),.B_bar(BLN4));
precharge_compiler inst_precharge5 (.clk(clk_bar),.B(BL5),.B_bar(BLN5));
precharge_compiler inst_precharge6 (.clk(clk_bar),.B(BL6),.B_bar(BLN6));
precharge_compiler inst_precharge7 (.clk(clk_bar),.B(BL7),.B_bar(BLN7));
precharge_compiler inst_precharge8 (.clk(clk_bar),.B(BL8),.B_bar(BLN8));
precharge_compiler inst_precharge9 (.clk(clk_bar),.B(BL9),.B_bar(BLN9));
precharge_compiler inst_precharge10 (.clk(clk_bar),.B(BL10),.B_bar(BLN10));
precharge_compiler inst_precharge11 (.clk(clk_bar),.B(BL11),.B_bar(BLN11));
precharge_compiler inst_precharge12 (.clk(clk_bar),.B(BL12),.B_bar(BLN12));
precharge_compiler inst_precharge13 (.clk(clk_bar),.B(BL13),.B_bar(BLN13));
precharge_compiler inst_precharge14 (.clk(clk_bar),.B(BL14),.B_bar(BLN14));
precharge_compiler inst_precharge15 (.clk(clk_bar),.B(BL15),.B_bar(BLN15));
precharge_compiler inst_precharge16 (.clk(clk_bar),.B(BL16),.B_bar(BLN16));
precharge_compiler inst_precharge17 (.clk(clk_bar),.B(BL17),.B_bar(BLN17));
precharge_compiler inst_precharge18 (.clk(clk_bar),.B(BL18),.B_bar(BLN18));
precharge_compiler inst_precharge19 (.clk(clk_bar),.B(BL19),.B_bar(BLN19));
precharge_compiler inst_precharge20 (.clk(clk_bar),.B(BL20),.B_bar(BLN20));
precharge_compiler inst_precharge21 (.clk(clk_bar),.B(BL21),.B_bar(BLN21));
precharge_compiler inst_precharge22 (.clk(clk_bar),.B(BL22),.B_bar(BLN22));
precharge_compiler inst_precharge23 (.clk(clk_bar),.B(BL23),.B_bar(BLN23));
precharge_compiler inst_precharge24 (.clk(clk_bar),.B(BL24),.B_bar(BLN24));
precharge_compiler inst_precharge25 (.clk(clk_bar),.B(BL25),.B_bar(BLN25));
precharge_compiler inst_precharge26 (.clk(clk_bar),.B(BL26),.B_bar(BLN26));
precharge_compiler inst_precharge27 (.clk(clk_bar),.B(BL27),.B_bar(BLN27));
precharge_compiler inst_precharge28 (.clk(clk_bar),.B(BL28),.B_bar(BLN28));
precharge_compiler inst_precharge29 (.clk(clk_bar),.B(BL29),.B_bar(BLN29));
precharge_compiler inst_precharge30 (.clk(clk_bar),.B(BL30),.B_bar(BLN30));
precharge_compiler inst_precharge31 (.clk(clk_bar),.B(BL31),.B_bar(BLN31));
precharge_compiler inst_precharge32 (.clk(clk_bar),.B(BL32),.B_bar(BLN32));
precharge_compiler inst_precharge33 (.clk(clk_bar),.B(BL33),.B_bar(BLN33));
precharge_compiler inst_precharge34 (.clk(clk_bar),.B(BL34),.B_bar(BLN34));
precharge_compiler inst_precharge35 (.clk(clk_bar),.B(BL35),.B_bar(BLN35));
precharge_compiler inst_precharge36 (.clk(clk_bar),.B(BL36),.B_bar(BLN36));
precharge_compiler inst_precharge37 (.clk(clk_bar),.B(BL37),.B_bar(BLN37));
precharge_compiler inst_precharge38 (.clk(clk_bar),.B(BL38),.B_bar(BLN38));
precharge_compiler inst_precharge39 (.clk(clk_bar),.B(BL39),.B_bar(BLN39));
precharge_compiler inst_precharge40 (.clk(clk_bar),.B(BL40),.B_bar(BLN40));
precharge_compiler inst_precharge41 (.clk(clk_bar),.B(BL41),.B_bar(BLN41));
precharge_compiler inst_precharge42 (.clk(clk_bar),.B(BL42),.B_bar(BLN42));
precharge_compiler inst_precharge43 (.clk(clk_bar),.B(BL43),.B_bar(BLN43));
precharge_compiler inst_precharge44 (.clk(clk_bar),.B(BL44),.B_bar(BLN44));
precharge_compiler inst_precharge45 (.clk(clk_bar),.B(BL45),.B_bar(BLN45));
precharge_compiler inst_precharge46 (.clk(clk_bar),.B(BL46),.B_bar(BLN46));
precharge_compiler inst_precharge47 (.clk(clk_bar),.B(BL47),.B_bar(BLN47));
precharge_compiler inst_precharge48 (.clk(clk_bar),.B(BL48),.B_bar(BLN48));
precharge_compiler inst_precharge49 (.clk(clk_bar),.B(BL49),.B_bar(BLN49));
precharge_compiler inst_precharge50 (.clk(clk_bar),.B(BL50),.B_bar(BLN50));
precharge_compiler inst_precharge51 (.clk(clk_bar),.B(BL51),.B_bar(BLN51));
precharge_compiler inst_precharge52 (.clk(clk_bar),.B(BL52),.B_bar(BLN52));
precharge_compiler inst_precharge53 (.clk(clk_bar),.B(BL53),.B_bar(BLN53));
precharge_compiler inst_precharge54 (.clk(clk_bar),.B(BL54),.B_bar(BLN54));
precharge_compiler inst_precharge55 (.clk(clk_bar),.B(BL55),.B_bar(BLN55));
precharge_compiler inst_precharge56 (.clk(clk_bar),.B(BL56),.B_bar(BLN56));
precharge_compiler inst_precharge57 (.clk(clk_bar),.B(BL57),.B_bar(BLN57));
precharge_compiler inst_precharge58 (.clk(clk_bar),.B(BL58),.B_bar(BLN58));
precharge_compiler inst_precharge59 (.clk(clk_bar),.B(BL59),.B_bar(BLN59));
precharge_compiler inst_precharge60 (.clk(clk_bar),.B(BL60),.B_bar(BLN60));
precharge_compiler inst_precharge61 (.clk(clk_bar),.B(BL61),.B_bar(BLN61));
precharge_compiler inst_precharge62 (.clk(clk_bar),.B(BL62),.B_bar(BLN62));
precharge_compiler inst_precharge63 (.clk(clk_bar),.B(BL63),.B_bar(BLN63));
precharge_compiler inst_precharge64 (.clk(clk_bar),.B(BL64),.B_bar(BLN64));
precharge_compiler inst_precharge65 (.clk(clk_bar),.B(BL65),.B_bar(BLN65));
precharge_compiler inst_precharge66 (.clk(clk_bar),.B(BL66),.B_bar(BLN66));
precharge_compiler inst_precharge67 (.clk(clk_bar),.B(BL67),.B_bar(BLN67));
precharge_compiler inst_precharge68 (.clk(clk_bar),.B(BL68),.B_bar(BLN68));
precharge_compiler inst_precharge69 (.clk(clk_bar),.B(BL69),.B_bar(BLN69));
precharge_compiler inst_precharge70 (.clk(clk_bar),.B(BL70),.B_bar(BLN70));
precharge_compiler inst_precharge71 (.clk(clk_bar),.B(BL71),.B_bar(BLN71));
precharge_compiler inst_precharge72 (.clk(clk_bar),.B(BL72),.B_bar(BLN72));
precharge_compiler inst_precharge73 (.clk(clk_bar),.B(BL73),.B_bar(BLN73));
precharge_compiler inst_precharge74 (.clk(clk_bar),.B(BL74),.B_bar(BLN74));
precharge_compiler inst_precharge75 (.clk(clk_bar),.B(BL75),.B_bar(BLN75));
precharge_compiler inst_precharge76 (.clk(clk_bar),.B(BL76),.B_bar(BLN76));
precharge_compiler inst_precharge77 (.clk(clk_bar),.B(BL77),.B_bar(BLN77));
precharge_compiler inst_precharge78 (.clk(clk_bar),.B(BL78),.B_bar(BLN78));
precharge_compiler inst_precharge79 (.clk(clk_bar),.B(BL79),.B_bar(BLN79));
precharge_compiler inst_precharge80 (.clk(clk_bar),.B(BL80),.B_bar(BLN80));
precharge_compiler inst_precharge81 (.clk(clk_bar),.B(BL81),.B_bar(BLN81));
precharge_compiler inst_precharge82 (.clk(clk_bar),.B(BL82),.B_bar(BLN82));
precharge_compiler inst_precharge83 (.clk(clk_bar),.B(BL83),.B_bar(BLN83));
precharge_compiler inst_precharge84 (.clk(clk_bar),.B(BL84),.B_bar(BLN84));
precharge_compiler inst_precharge85 (.clk(clk_bar),.B(BL85),.B_bar(BLN85));
precharge_compiler inst_precharge86 (.clk(clk_bar),.B(BL86),.B_bar(BLN86));
precharge_compiler inst_precharge87 (.clk(clk_bar),.B(BL87),.B_bar(BLN87));
precharge_compiler inst_precharge88 (.clk(clk_bar),.B(BL88),.B_bar(BLN88));
precharge_compiler inst_precharge89 (.clk(clk_bar),.B(BL89),.B_bar(BLN89));
precharge_compiler inst_precharge90 (.clk(clk_bar),.B(BL90),.B_bar(BLN90));
precharge_compiler inst_precharge91 (.clk(clk_bar),.B(BL91),.B_bar(BLN91));
precharge_compiler inst_precharge92 (.clk(clk_bar),.B(BL92),.B_bar(BLN92));
precharge_compiler inst_precharge93 (.clk(clk_bar),.B(BL93),.B_bar(BLN93));
precharge_compiler inst_precharge94 (.clk(clk_bar),.B(BL94),.B_bar(BLN94));
precharge_compiler inst_precharge95 (.clk(clk_bar),.B(BL95),.B_bar(BLN95));
precharge_compiler inst_precharge96 (.clk(clk_bar),.B(BL96),.B_bar(BLN96));
precharge_compiler inst_precharge97 (.clk(clk_bar),.B(BL97),.B_bar(BLN97));
precharge_compiler inst_precharge98 (.clk(clk_bar),.B(BL98),.B_bar(BLN98));
precharge_compiler inst_precharge99 (.clk(clk_bar),.B(BL99),.B_bar(BLN99));
precharge_compiler inst_precharge100 (.clk(clk_bar),.B(BL100),.B_bar(BLN100));
precharge_compiler inst_precharge101 (.clk(clk_bar),.B(BL101),.B_bar(BLN101));
precharge_compiler inst_precharge102 (.clk(clk_bar),.B(BL102),.B_bar(BLN102));
precharge_compiler inst_precharge103 (.clk(clk_bar),.B(BL103),.B_bar(BLN103));
precharge_compiler inst_precharge104 (.clk(clk_bar),.B(BL104),.B_bar(BLN104));
precharge_compiler inst_precharge105 (.clk(clk_bar),.B(BL105),.B_bar(BLN105));
precharge_compiler inst_precharge106 (.clk(clk_bar),.B(BL106),.B_bar(BLN106));
precharge_compiler inst_precharge107 (.clk(clk_bar),.B(BL107),.B_bar(BLN107));
precharge_compiler inst_precharge108 (.clk(clk_bar),.B(BL108),.B_bar(BLN108));
precharge_compiler inst_precharge109 (.clk(clk_bar),.B(BL109),.B_bar(BLN109));
precharge_compiler inst_precharge110 (.clk(clk_bar),.B(BL110),.B_bar(BLN110));
precharge_compiler inst_precharge111 (.clk(clk_bar),.B(BL111),.B_bar(BLN111));
precharge_compiler inst_precharge112 (.clk(clk_bar),.B(BL112),.B_bar(BLN112));
precharge_compiler inst_precharge113 (.clk(clk_bar),.B(BL113),.B_bar(BLN113));
precharge_compiler inst_precharge114 (.clk(clk_bar),.B(BL114),.B_bar(BLN114));
precharge_compiler inst_precharge115 (.clk(clk_bar),.B(BL115),.B_bar(BLN115));
precharge_compiler inst_precharge116 (.clk(clk_bar),.B(BL116),.B_bar(BLN116));
precharge_compiler inst_precharge117 (.clk(clk_bar),.B(BL117),.B_bar(BLN117));
precharge_compiler inst_precharge118 (.clk(clk_bar),.B(BL118),.B_bar(BLN118));
precharge_compiler inst_precharge119 (.clk(clk_bar),.B(BL119),.B_bar(BLN119));
precharge_compiler inst_precharge120 (.clk(clk_bar),.B(BL120),.B_bar(BLN120));
precharge_compiler inst_precharge121 (.clk(clk_bar),.B(BL121),.B_bar(BLN121));
precharge_compiler inst_precharge122 (.clk(clk_bar),.B(BL122),.B_bar(BLN122));
precharge_compiler inst_precharge123 (.clk(clk_bar),.B(BL123),.B_bar(BLN123));
precharge_compiler inst_precharge124 (.clk(clk_bar),.B(BL124),.B_bar(BLN124));
precharge_compiler inst_precharge125 (.clk(clk_bar),.B(BL125),.B_bar(BLN125));
precharge_compiler inst_precharge126 (.clk(clk_bar),.B(BL126),.B_bar(BLN126));
precharge_compiler inst_precharge127 (.clk(clk_bar),.B(BL127),.B_bar(BLN127));
endmodule
