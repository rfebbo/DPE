VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_1kb_64x128x32
  CLASS BLOCK ;
  ORIGIN 39.505 120.605 ;
  FOREIGN sram_1kb_64x128x32 -39.505 -120.605 ;
  SIZE 197.97 BY 130.5 ;
  SYMMETRY X Y R90 ;
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.235 -111.125 151.98 -111.035 ;
        RECT 151.8 -111.215 151.98 -111.035 ;
        RECT 147 -111.215 147.18 -111.035 ;
        RECT 142.2 -111.215 142.38 -111.035 ;
        RECT 137.4 -111.215 137.58 -111.035 ;
        RECT 132.6 -111.215 132.78 -111.035 ;
        RECT 127.8 -111.215 127.98 -111.035 ;
        RECT 123 -111.215 123.18 -111.035 ;
        RECT 118.2 -111.215 118.38 -111.035 ;
        RECT 113.4 -111.215 113.58 -111.035 ;
        RECT 108.6 -111.215 108.78 -111.035 ;
        RECT 103.8 -111.215 103.98 -111.035 ;
        RECT 99 -111.215 99.18 -111.035 ;
        RECT 94.2 -111.215 94.38 -111.035 ;
        RECT 89.4 -111.215 89.58 -111.035 ;
        RECT 84.6 -111.215 84.78 -111.035 ;
        RECT 79.8 -111.215 79.98 -111.035 ;
        RECT 75 -111.215 75.18 -111.035 ;
        RECT 70.2 -111.215 70.38 -111.035 ;
        RECT 65.4 -111.215 65.58 -111.035 ;
        RECT 60.6 -111.215 60.78 -111.035 ;
        RECT 55.8 -111.215 55.98 -111.035 ;
        RECT 51 -111.215 51.18 -111.035 ;
        RECT 46.2 -111.215 46.38 -111.035 ;
        RECT 41.4 -111.215 41.58 -111.035 ;
        RECT 36.6 -111.215 36.78 -111.035 ;
        RECT 31.8 -111.215 31.98 -111.035 ;
        RECT 27 -111.215 27.18 -111.035 ;
        RECT 22.2 -111.215 22.38 -111.035 ;
        RECT 17.4 -111.215 17.58 -111.035 ;
        RECT 12.6 -111.215 12.78 -111.035 ;
        RECT 7.8 -111.215 7.98 -111.035 ;
        RECT 3 -111.215 3.18 -111.035 ;
    END
  END write_en
  PIN din0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.29 -111.445 -0.06 -111.215 ;
      LAYER M3 ;
        RECT -0.29 -111.445 -0.06 -111.215 ;
      LAYER M1 ;
        RECT -0.29 -111.305 1.575 -111.215 ;
        RECT -0.29 -111.445 -0.06 -111.215 ;
    END
  END din0
  PIN din1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.51 -111.445 4.74 -111.215 ;
      LAYER M3 ;
        RECT 4.51 -111.445 4.74 -111.215 ;
      LAYER M1 ;
        RECT 4.51 -111.305 6.375 -111.215 ;
        RECT 4.51 -111.445 4.74 -111.215 ;
    END
  END din1
  PIN din2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.31 -111.445 9.54 -111.215 ;
      LAYER M3 ;
        RECT 9.31 -111.445 9.54 -111.215 ;
      LAYER M1 ;
        RECT 9.31 -111.305 11.175 -111.215 ;
        RECT 9.31 -111.445 9.54 -111.215 ;
    END
  END din2
  PIN din3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.11 -111.445 14.34 -111.215 ;
      LAYER M3 ;
        RECT 14.11 -111.445 14.34 -111.215 ;
      LAYER M1 ;
        RECT 14.11 -111.305 15.975 -111.215 ;
        RECT 14.11 -111.445 14.34 -111.215 ;
    END
  END din3
  PIN din4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.91 -111.445 19.14 -111.215 ;
      LAYER M3 ;
        RECT 18.91 -111.445 19.14 -111.215 ;
      LAYER M1 ;
        RECT 18.91 -111.305 20.775 -111.215 ;
        RECT 18.91 -111.445 19.14 -111.215 ;
    END
  END din4
  PIN din5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.71 -111.445 23.94 -111.215 ;
      LAYER M3 ;
        RECT 23.71 -111.445 23.94 -111.215 ;
      LAYER M1 ;
        RECT 23.71 -111.305 25.575 -111.215 ;
        RECT 23.71 -111.445 23.94 -111.215 ;
    END
  END din5
  PIN din6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.51 -111.445 28.74 -111.215 ;
      LAYER M3 ;
        RECT 28.51 -111.445 28.74 -111.215 ;
      LAYER M1 ;
        RECT 28.51 -111.305 30.375 -111.215 ;
        RECT 28.51 -111.445 28.74 -111.215 ;
    END
  END din6
  PIN din7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.31 -111.445 33.54 -111.215 ;
      LAYER M3 ;
        RECT 33.31 -111.445 33.54 -111.215 ;
      LAYER M1 ;
        RECT 33.31 -111.305 35.175 -111.215 ;
        RECT 33.31 -111.445 33.54 -111.215 ;
    END
  END din7
  PIN din8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.11 -111.445 38.34 -111.215 ;
      LAYER M3 ;
        RECT 38.11 -111.445 38.34 -111.215 ;
      LAYER M1 ;
        RECT 38.11 -111.305 39.975 -111.215 ;
        RECT 38.11 -111.445 38.34 -111.215 ;
    END
  END din8
  PIN din9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.91 -111.445 43.14 -111.215 ;
      LAYER M3 ;
        RECT 42.91 -111.445 43.14 -111.215 ;
      LAYER M1 ;
        RECT 42.91 -111.305 44.775 -111.215 ;
        RECT 42.91 -111.445 43.14 -111.215 ;
    END
  END din9
  PIN din10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.71 -111.445 47.94 -111.215 ;
      LAYER M3 ;
        RECT 47.71 -111.445 47.94 -111.215 ;
      LAYER M1 ;
        RECT 47.71 -111.305 49.575 -111.215 ;
        RECT 47.71 -111.445 47.94 -111.215 ;
    END
  END din10
  PIN din11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.51 -111.445 52.74 -111.215 ;
      LAYER M3 ;
        RECT 52.51 -111.445 52.74 -111.215 ;
      LAYER M1 ;
        RECT 52.51 -111.305 54.375 -111.215 ;
        RECT 52.51 -111.445 52.74 -111.215 ;
    END
  END din11
  PIN din12
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.31 -111.445 57.54 -111.215 ;
      LAYER M3 ;
        RECT 57.31 -111.445 57.54 -111.215 ;
      LAYER M1 ;
        RECT 57.31 -111.305 59.175 -111.215 ;
        RECT 57.31 -111.445 57.54 -111.215 ;
    END
  END din12
  PIN din13
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.11 -111.445 62.34 -111.215 ;
      LAYER M3 ;
        RECT 62.11 -111.445 62.34 -111.215 ;
      LAYER M1 ;
        RECT 62.11 -111.305 63.975 -111.215 ;
        RECT 62.11 -111.445 62.34 -111.215 ;
    END
  END din13
  PIN din14
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.91 -111.445 67.14 -111.215 ;
      LAYER M3 ;
        RECT 66.91 -111.445 67.14 -111.215 ;
      LAYER M1 ;
        RECT 66.91 -111.305 68.775 -111.215 ;
        RECT 66.91 -111.445 67.14 -111.215 ;
    END
  END din14
  PIN din15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.71 -111.445 71.94 -111.215 ;
      LAYER M3 ;
        RECT 71.71 -111.445 71.94 -111.215 ;
      LAYER M1 ;
        RECT 71.71 -111.305 73.575 -111.215 ;
        RECT 71.71 -111.445 71.94 -111.215 ;
    END
  END din15
  PIN din16
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.51 -111.445 76.74 -111.215 ;
      LAYER M3 ;
        RECT 76.51 -111.445 76.74 -111.215 ;
      LAYER M1 ;
        RECT 76.51 -111.305 78.375 -111.215 ;
        RECT 76.51 -111.445 76.74 -111.215 ;
    END
  END din16
  PIN din17
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.31 -111.445 81.54 -111.215 ;
      LAYER M3 ;
        RECT 81.31 -111.445 81.54 -111.215 ;
      LAYER M1 ;
        RECT 81.31 -111.305 83.175 -111.215 ;
        RECT 81.31 -111.445 81.54 -111.215 ;
    END
  END din17
  PIN din18
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.11 -111.445 86.34 -111.215 ;
      LAYER M3 ;
        RECT 86.11 -111.445 86.34 -111.215 ;
      LAYER M1 ;
        RECT 86.11 -111.305 87.975 -111.215 ;
        RECT 86.11 -111.445 86.34 -111.215 ;
    END
  END din18
  PIN din19
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.91 -111.445 91.14 -111.215 ;
      LAYER M3 ;
        RECT 90.91 -111.445 91.14 -111.215 ;
      LAYER M1 ;
        RECT 90.91 -111.305 92.775 -111.215 ;
        RECT 90.91 -111.445 91.14 -111.215 ;
    END
  END din19
  PIN din20
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.71 -111.445 95.94 -111.215 ;
      LAYER M3 ;
        RECT 95.71 -111.445 95.94 -111.215 ;
      LAYER M1 ;
        RECT 95.71 -111.305 97.575 -111.215 ;
        RECT 95.71 -111.445 95.94 -111.215 ;
    END
  END din20
  PIN din21
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.51 -111.445 100.74 -111.215 ;
      LAYER M3 ;
        RECT 100.51 -111.445 100.74 -111.215 ;
      LAYER M1 ;
        RECT 100.51 -111.305 102.375 -111.215 ;
        RECT 100.51 -111.445 100.74 -111.215 ;
    END
  END din21
  PIN din22
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.31 -111.445 105.54 -111.215 ;
      LAYER M3 ;
        RECT 105.31 -111.445 105.54 -111.215 ;
      LAYER M1 ;
        RECT 105.31 -111.305 107.175 -111.215 ;
        RECT 105.31 -111.445 105.54 -111.215 ;
    END
  END din22
  PIN din23
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.11 -111.445 110.34 -111.215 ;
      LAYER M3 ;
        RECT 110.11 -111.445 110.34 -111.215 ;
      LAYER M1 ;
        RECT 110.11 -111.305 111.975 -111.215 ;
        RECT 110.11 -111.445 110.34 -111.215 ;
    END
  END din23
  PIN din24
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.91 -111.445 115.14 -111.215 ;
      LAYER M3 ;
        RECT 114.91 -111.445 115.14 -111.215 ;
      LAYER M1 ;
        RECT 114.91 -111.305 116.775 -111.215 ;
        RECT 114.91 -111.445 115.14 -111.215 ;
    END
  END din24
  PIN din25
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.71 -111.445 119.94 -111.215 ;
      LAYER M3 ;
        RECT 119.71 -111.445 119.94 -111.215 ;
      LAYER M1 ;
        RECT 119.71 -111.305 121.575 -111.215 ;
        RECT 119.71 -111.445 119.94 -111.215 ;
    END
  END din25
  PIN din26
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.51 -111.445 124.74 -111.215 ;
      LAYER M3 ;
        RECT 124.51 -111.445 124.74 -111.215 ;
      LAYER M1 ;
        RECT 124.51 -111.305 126.375 -111.215 ;
        RECT 124.51 -111.445 124.74 -111.215 ;
    END
  END din26
  PIN din27
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.31 -111.445 129.54 -111.215 ;
      LAYER M3 ;
        RECT 129.31 -111.445 129.54 -111.215 ;
      LAYER M1 ;
        RECT 129.31 -111.305 131.175 -111.215 ;
        RECT 129.31 -111.445 129.54 -111.215 ;
    END
  END din27
  PIN din28
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.11 -111.445 134.34 -111.215 ;
      LAYER M3 ;
        RECT 134.11 -111.445 134.34 -111.215 ;
      LAYER M1 ;
        RECT 134.11 -111.305 135.975 -111.215 ;
        RECT 134.11 -111.445 134.34 -111.215 ;
    END
  END din28
  PIN din29
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.91 -111.445 139.14 -111.215 ;
      LAYER M3 ;
        RECT 138.91 -111.445 139.14 -111.215 ;
      LAYER M1 ;
        RECT 138.91 -111.305 140.775 -111.215 ;
        RECT 138.91 -111.445 139.14 -111.215 ;
    END
  END din29
  PIN din30
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.71 -111.445 143.94 -111.215 ;
      LAYER M3 ;
        RECT 143.71 -111.445 143.94 -111.215 ;
      LAYER M1 ;
        RECT 143.71 -111.305 145.575 -111.215 ;
        RECT 143.71 -111.445 143.94 -111.215 ;
    END
  END din30
  PIN din31
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.51 -111.445 148.74 -111.215 ;
      LAYER M3 ;
        RECT 148.51 -111.445 148.74 -111.215 ;
      LAYER M1 ;
        RECT 148.51 -111.305 150.375 -111.215 ;
        RECT 148.51 -111.445 148.74 -111.215 ;
    END
  END din31
  PIN sense_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.03 -114.105 149.685 -113.985 ;
    END
  END sense_en
  PIN dout0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9 -113.85 2 -113.1 ;
        RECT -0.03 -113.795 2 -113.675 ;
        RECT 1.53 -113.85 2 -113.675 ;
        RECT 0.355 -113.795 0.455 -113.09 ;
    END
  END dout0
  PIN dout1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.7 -113.85 6.8 -113.1 ;
        RECT 4.77 -113.795 6.8 -113.675 ;
        RECT 6.33 -113.85 6.8 -113.675 ;
        RECT 5.155 -113.795 5.255 -113.09 ;
    END
  END dout1
  PIN dout2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.5 -113.85 11.6 -113.1 ;
        RECT 9.57 -113.795 11.6 -113.675 ;
        RECT 11.13 -113.85 11.6 -113.675 ;
        RECT 9.955 -113.795 10.055 -113.09 ;
    END
  END dout2
  PIN dout3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.3 -113.85 16.4 -113.1 ;
        RECT 14.37 -113.795 16.4 -113.675 ;
        RECT 15.93 -113.85 16.4 -113.675 ;
        RECT 14.755 -113.795 14.855 -113.09 ;
    END
  END dout3
  PIN dout4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 21.1 -113.85 21.2 -113.1 ;
        RECT 19.17 -113.795 21.2 -113.675 ;
        RECT 20.73 -113.85 21.2 -113.675 ;
        RECT 19.555 -113.795 19.655 -113.09 ;
    END
  END dout4
  PIN dout5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 25.9 -113.85 26 -113.1 ;
        RECT 23.97 -113.795 26 -113.675 ;
        RECT 25.53 -113.85 26 -113.675 ;
        RECT 24.355 -113.795 24.455 -113.09 ;
    END
  END dout5
  PIN dout6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 30.7 -113.85 30.8 -113.1 ;
        RECT 28.77 -113.795 30.8 -113.675 ;
        RECT 30.33 -113.85 30.8 -113.675 ;
        RECT 29.155 -113.795 29.255 -113.09 ;
    END
  END dout6
  PIN dout7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 35.5 -113.85 35.6 -113.1 ;
        RECT 33.57 -113.795 35.6 -113.675 ;
        RECT 35.13 -113.85 35.6 -113.675 ;
        RECT 33.955 -113.795 34.055 -113.09 ;
    END
  END dout7
  PIN dout8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.3 -113.85 40.4 -113.1 ;
        RECT 38.37 -113.795 40.4 -113.675 ;
        RECT 39.93 -113.85 40.4 -113.675 ;
        RECT 38.755 -113.795 38.855 -113.09 ;
    END
  END dout8
  PIN dout9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 45.1 -113.85 45.2 -113.1 ;
        RECT 43.17 -113.795 45.2 -113.675 ;
        RECT 44.73 -113.85 45.2 -113.675 ;
        RECT 43.555 -113.795 43.655 -113.09 ;
    END
  END dout9
  PIN dout10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 49.9 -113.85 50 -113.1 ;
        RECT 47.97 -113.795 50 -113.675 ;
        RECT 49.53 -113.85 50 -113.675 ;
        RECT 48.355 -113.795 48.455 -113.09 ;
    END
  END dout10
  PIN dout11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 54.7 -113.85 54.8 -113.1 ;
        RECT 52.77 -113.795 54.8 -113.675 ;
        RECT 54.33 -113.85 54.8 -113.675 ;
        RECT 53.155 -113.795 53.255 -113.09 ;
    END
  END dout11
  PIN dout12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 59.5 -113.85 59.6 -113.1 ;
        RECT 57.57 -113.795 59.6 -113.675 ;
        RECT 59.13 -113.85 59.6 -113.675 ;
        RECT 57.955 -113.795 58.055 -113.09 ;
    END
  END dout12
  PIN dout13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 64.3 -113.85 64.4 -113.1 ;
        RECT 62.37 -113.795 64.4 -113.675 ;
        RECT 63.93 -113.85 64.4 -113.675 ;
        RECT 62.755 -113.795 62.855 -113.09 ;
    END
  END dout13
  PIN dout14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 69.1 -113.85 69.2 -113.1 ;
        RECT 67.17 -113.795 69.2 -113.675 ;
        RECT 68.73 -113.85 69.2 -113.675 ;
        RECT 67.555 -113.795 67.655 -113.09 ;
    END
  END dout14
  PIN dout15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 73.9 -113.85 74 -113.1 ;
        RECT 71.97 -113.795 74 -113.675 ;
        RECT 73.53 -113.85 74 -113.675 ;
        RECT 72.355 -113.795 72.455 -113.09 ;
    END
  END dout15
  PIN dout16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 78.7 -113.85 78.8 -113.1 ;
        RECT 76.77 -113.795 78.8 -113.675 ;
        RECT 78.33 -113.85 78.8 -113.675 ;
        RECT 77.155 -113.795 77.255 -113.09 ;
    END
  END dout16
  PIN dout17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 83.5 -113.85 83.6 -113.1 ;
        RECT 81.57 -113.795 83.6 -113.675 ;
        RECT 83.13 -113.85 83.6 -113.675 ;
        RECT 81.955 -113.795 82.055 -113.09 ;
    END
  END dout17
  PIN dout18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 88.3 -113.85 88.4 -113.1 ;
        RECT 86.37 -113.795 88.4 -113.675 ;
        RECT 87.93 -113.85 88.4 -113.675 ;
        RECT 86.755 -113.795 86.855 -113.09 ;
    END
  END dout18
  PIN dout19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 93.1 -113.85 93.2 -113.1 ;
        RECT 91.17 -113.795 93.2 -113.675 ;
        RECT 92.73 -113.85 93.2 -113.675 ;
        RECT 91.555 -113.795 91.655 -113.09 ;
    END
  END dout19
  PIN dout20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 97.9 -113.85 98 -113.1 ;
        RECT 95.97 -113.795 98 -113.675 ;
        RECT 97.53 -113.85 98 -113.675 ;
        RECT 96.355 -113.795 96.455 -113.09 ;
    END
  END dout20
  PIN dout21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 102.7 -113.85 102.8 -113.1 ;
        RECT 100.77 -113.795 102.8 -113.675 ;
        RECT 102.33 -113.85 102.8 -113.675 ;
        RECT 101.155 -113.795 101.255 -113.09 ;
    END
  END dout21
  PIN dout22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 107.5 -113.85 107.6 -113.1 ;
        RECT 105.57 -113.795 107.6 -113.675 ;
        RECT 107.13 -113.85 107.6 -113.675 ;
        RECT 105.955 -113.795 106.055 -113.09 ;
    END
  END dout22
  PIN dout23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 112.3 -113.85 112.4 -113.1 ;
        RECT 110.37 -113.795 112.4 -113.675 ;
        RECT 111.93 -113.85 112.4 -113.675 ;
        RECT 110.755 -113.795 110.855 -113.09 ;
    END
  END dout23
  PIN dout24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 117.1 -113.85 117.2 -113.1 ;
        RECT 115.17 -113.795 117.2 -113.675 ;
        RECT 116.73 -113.85 117.2 -113.675 ;
        RECT 115.555 -113.795 115.655 -113.09 ;
    END
  END dout24
  PIN dout25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 121.9 -113.85 122 -113.1 ;
        RECT 119.97 -113.795 122 -113.675 ;
        RECT 121.53 -113.85 122 -113.675 ;
        RECT 120.355 -113.795 120.455 -113.09 ;
    END
  END dout25
  PIN dout26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 126.7 -113.85 126.8 -113.1 ;
        RECT 124.77 -113.795 126.8 -113.675 ;
        RECT 126.33 -113.85 126.8 -113.675 ;
        RECT 125.155 -113.795 125.255 -113.09 ;
    END
  END dout26
  PIN dout27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 131.5 -113.85 131.6 -113.1 ;
        RECT 129.57 -113.795 131.6 -113.675 ;
        RECT 131.13 -113.85 131.6 -113.675 ;
        RECT 129.955 -113.795 130.055 -113.09 ;
    END
  END dout27
  PIN dout28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 136.3 -113.85 136.4 -113.1 ;
        RECT 134.37 -113.795 136.4 -113.675 ;
        RECT 135.93 -113.85 136.4 -113.675 ;
        RECT 134.755 -113.795 134.855 -113.09 ;
    END
  END dout28
  PIN dout29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 141.1 -113.85 141.2 -113.1 ;
        RECT 139.17 -113.795 141.2 -113.675 ;
        RECT 140.73 -113.85 141.2 -113.675 ;
        RECT 139.555 -113.795 139.655 -113.09 ;
    END
  END dout29
  PIN dout30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 145.9 -113.85 146 -113.1 ;
        RECT 143.97 -113.795 146 -113.675 ;
        RECT 145.53 -113.85 146 -113.675 ;
        RECT 144.355 -113.795 144.455 -113.09 ;
    END
  END dout30
  PIN dout31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 150.7 -113.85 150.8 -113.1 ;
        RECT 148.77 -113.795 150.8 -113.675 ;
        RECT 150.33 -113.85 150.8 -113.675 ;
        RECT 149.155 -113.795 149.255 -113.09 ;
    END
  END dout31
  PIN gnd!
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 155.747 7.175 158.465 9.895 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -39.325 -120.365 -36.607 -117.645 ;
    END
    PORT
      LAYER M1 ;
        RECT 155.747 -120.365 158.465 -117.645 ;
    END
  END vdd!
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -6.835 3.435 -5.845 3.535 ;
    END
  END clk
  PIN addr5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -35.545 -100.715 -35.365 0.645 ;
        RECT -35.545 -100.715 -35.445 3.005 ;
      LAYER M1 ;
        RECT -35.845 -98.715 -9.26 -98.615 ;
        RECT -35.845 -91.955 -9.26 -91.855 ;
        RECT -35.845 -85.795 -9.26 -85.695 ;
        RECT -35.845 -79.035 -9.26 -78.935 ;
        RECT -35.845 -72.875 -9.26 -72.775 ;
        RECT -35.845 -66.115 -9.26 -66.015 ;
        RECT -35.845 -59.955 -9.26 -59.855 ;
        RECT -35.845 -53.195 -9.26 -53.095 ;
        RECT -35.625 2.825 -35.24 3.005 ;
    END
  END addr5
  PIN addr4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -34.945 -100.715 -34.765 0.645 ;
        RECT -34.945 -100.715 -34.845 3.345 ;
      LAYER M1 ;
        RECT -35.845 -98.935 -9.52 -98.835 ;
        RECT -35.845 -91.735 -9.52 -91.635 ;
        RECT -35.845 -86.015 -9.52 -85.915 ;
        RECT -35.845 -78.815 -9.52 -78.715 ;
        RECT -35.845 -47.255 -9.52 -47.155 ;
        RECT -35.845 -40.055 -9.52 -39.955 ;
        RECT -35.845 -34.335 -9.52 -34.235 ;
        RECT -35.845 -27.135 -9.52 -27.035 ;
        RECT -35.625 3.165 -34.64 3.345 ;
    END
  END addr4
  PIN addr3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -34.345 -100.715 -34.165 0.645 ;
        RECT -34.345 -100.715 -34.245 3.685 ;
      LAYER M1 ;
        RECT -35.845 -99.155 -10.56 -99.055 ;
        RECT -35.845 -91.515 -10.56 -91.415 ;
        RECT -35.845 -73.315 -10.56 -73.215 ;
        RECT -35.845 -65.675 -10.56 -65.575 ;
        RECT -35.845 -47.475 -10.56 -47.375 ;
        RECT -35.845 -39.835 -10.56 -39.735 ;
        RECT -35.845 -21.635 -10.56 -21.535 ;
        RECT -35.845 -13.995 -10.56 -13.895 ;
        RECT -35.625 3.505 -34.04 3.685 ;
    END
  END addr3
  PIN addr2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -33.745 -100.715 -33.565 0.645 ;
        RECT -33.745 -100.715 -33.645 4.025 ;
      LAYER M1 ;
        RECT -35.845 -99.375 -10.82 -99.275 ;
        RECT -35.845 -86.455 -10.82 -86.355 ;
        RECT -35.845 -73.535 -10.82 -73.435 ;
        RECT -35.845 -60.615 -10.82 -60.515 ;
        RECT -35.845 -47.695 -10.82 -47.595 ;
        RECT -35.845 -34.775 -10.82 -34.675 ;
        RECT -35.845 -21.855 -10.82 -21.755 ;
        RECT -35.845 -8.935 -10.82 -8.835 ;
        RECT -35.625 3.845 -33.44 4.025 ;
    END
  END addr2
  PIN addr1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -33.145 -100.715 -32.965 0.645 ;
        RECT -33.145 -100.715 -33.045 4.365 ;
      LAYER M1 ;
        RECT -35.845 -99.595 -11.86 -99.495 ;
        RECT -35.845 -91.075 -11.86 -90.975 ;
        RECT -35.845 -86.675 -11.86 -86.575 ;
        RECT -35.845 -78.155 -11.86 -78.055 ;
        RECT -35.845 -73.755 -11.86 -73.655 ;
        RECT -35.845 -65.235 -11.86 -65.135 ;
        RECT -35.845 -60.835 -11.86 -60.735 ;
        RECT -35.845 -52.315 -11.86 -52.215 ;
        RECT -35.845 -47.915 -11.86 -47.815 ;
        RECT -35.845 -39.395 -11.86 -39.295 ;
        RECT -35.845 -34.995 -11.86 -34.895 ;
        RECT -35.845 -26.475 -11.86 -26.375 ;
        RECT -35.845 -22.075 -11.86 -21.975 ;
        RECT -35.845 -13.555 -11.86 -13.455 ;
        RECT -35.845 -9.155 -11.86 -9.055 ;
        RECT -35.845 -0.635 -11.86 -0.535 ;
        RECT -35.625 4.185 -32.84 4.365 ;
    END
  END addr1
  PIN addr0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -32.545 -100.715 -32.365 0.645 ;
        RECT -32.545 -100.715 -32.445 4.705 ;
      LAYER M1 ;
        RECT -35.845 -100.035 -12.12 -99.935 ;
        RECT -35.845 -90.635 -12.12 -90.535 ;
        RECT -35.845 -87.115 -12.12 -87.015 ;
        RECT -35.845 -77.715 -12.12 -77.615 ;
        RECT -35.845 -74.195 -12.12 -74.095 ;
        RECT -35.845 -64.795 -12.12 -64.695 ;
        RECT -35.845 -61.275 -12.12 -61.175 ;
        RECT -35.845 -51.875 -12.12 -51.775 ;
        RECT -35.845 -48.355 -12.12 -48.255 ;
        RECT -35.845 -38.955 -12.12 -38.855 ;
        RECT -35.845 -35.435 -12.12 -35.335 ;
        RECT -35.845 -26.035 -12.12 -25.935 ;
        RECT -35.845 -22.515 -12.12 -22.415 ;
        RECT -35.845 -13.115 -12.12 -13.015 ;
        RECT -35.845 -9.595 -12.12 -9.495 ;
        RECT -35.845 -0.195 -12.12 -0.095 ;
        RECT -35.625 4.525 -32.24 4.705 ;
    END
  END addr0
  PIN addr7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -12.345 -107.175 -12.165 -102.715 ;
        RECT -12.345 -109.975 -12.245 -102.715 ;
      LAYER M1 ;
        RECT -12.645 -103.995 -6.66 -103.895 ;
        RECT -12.425 -109.975 -12.04 -109.795 ;
    END
  END addr7
  PIN addr6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -11.745 -107.175 -11.565 -102.715 ;
        RECT -11.745 -109.635 -11.645 -102.715 ;
      LAYER M1 ;
        RECT -12.645 -103.555 -6.92 -103.455 ;
        RECT -12.425 -109.635 -11.44 -109.455 ;
    END
  END addr6
  OBS
    LAYER M1 SPACING 0.16 ;
      RECT 149.79 -115.455 149.89 -114.68 ;
      RECT 149.23 -115.455 149.33 -114.68 ;
      RECT 144.99 -115.455 145.09 -114.68 ;
      RECT 144.43 -115.455 144.53 -114.68 ;
      RECT 140.19 -115.455 140.29 -114.68 ;
      RECT 139.63 -115.455 139.73 -114.68 ;
      RECT 135.39 -115.455 135.49 -114.68 ;
      RECT 134.83 -115.455 134.93 -114.68 ;
      RECT 130.59 -115.455 130.69 -114.68 ;
      RECT 130.03 -115.455 130.13 -114.68 ;
      RECT 125.79 -115.455 125.89 -114.68 ;
      RECT 125.23 -115.455 125.33 -114.68 ;
      RECT 120.99 -115.455 121.09 -114.68 ;
      RECT 120.43 -115.455 120.53 -114.68 ;
      RECT 116.19 -115.455 116.29 -114.68 ;
      RECT 115.63 -115.455 115.73 -114.68 ;
      RECT 111.39 -115.455 111.49 -114.68 ;
      RECT 110.83 -115.455 110.93 -114.68 ;
      RECT 106.59 -115.455 106.69 -114.68 ;
      RECT 106.03 -115.455 106.13 -114.68 ;
      RECT 101.79 -115.455 101.89 -114.68 ;
      RECT 101.23 -115.455 101.33 -114.68 ;
      RECT 96.99 -115.455 97.09 -114.68 ;
      RECT 96.43 -115.455 96.53 -114.68 ;
      RECT 92.19 -115.455 92.29 -114.68 ;
      RECT 91.63 -115.455 91.73 -114.68 ;
      RECT 87.39 -115.455 87.49 -114.68 ;
      RECT 86.83 -115.455 86.93 -114.68 ;
      RECT 82.59 -115.455 82.69 -114.68 ;
      RECT 82.03 -115.455 82.13 -114.68 ;
      RECT 77.79 -115.455 77.89 -114.68 ;
      RECT 77.23 -115.455 77.33 -114.68 ;
      RECT 72.99 -115.455 73.09 -114.68 ;
      RECT 72.43 -115.455 72.53 -114.68 ;
      RECT 68.19 -115.455 68.29 -114.68 ;
      RECT 67.63 -115.455 67.73 -114.68 ;
      RECT 63.39 -115.455 63.49 -114.68 ;
      RECT 62.83 -115.455 62.93 -114.68 ;
      RECT 58.59 -115.455 58.69 -114.68 ;
      RECT 58.03 -115.455 58.13 -114.68 ;
      RECT 53.79 -115.455 53.89 -114.68 ;
      RECT 53.23 -115.455 53.33 -114.68 ;
      RECT 48.99 -115.455 49.09 -114.68 ;
      RECT 48.43 -115.455 48.53 -114.68 ;
      RECT 44.19 -115.455 44.29 -114.68 ;
      RECT 43.63 -115.455 43.73 -114.68 ;
      RECT 39.39 -115.455 39.49 -114.68 ;
      RECT 38.83 -115.455 38.93 -114.68 ;
      RECT 34.59 -115.455 34.69 -114.68 ;
      RECT 34.03 -115.455 34.13 -114.68 ;
      RECT 29.79 -115.455 29.89 -114.68 ;
      RECT 29.23 -115.455 29.33 -114.68 ;
      RECT 24.99 -115.455 25.09 -114.68 ;
      RECT 24.43 -115.455 24.53 -114.68 ;
      RECT 20.19 -115.455 20.29 -114.68 ;
      RECT 19.63 -115.455 19.73 -114.68 ;
      RECT 15.39 -115.455 15.49 -114.68 ;
      RECT 14.83 -115.455 14.93 -114.68 ;
      RECT 10.59 -115.455 10.69 -114.68 ;
      RECT 10.03 -115.455 10.13 -114.68 ;
      RECT 5.79 -115.455 5.89 -114.68 ;
      RECT 5.23 -115.455 5.33 -114.68 ;
      RECT 0.99 -115.455 1.09 -114.68 ;
      RECT 0.43 -115.455 0.53 -114.68 ;
      RECT 0.025 -115.455 158.465 -115.095 ;
      RECT 152.825 -110.195 152.925 -109.27 ;
      RECT 152.265 -110.195 152.365 -109.27 ;
      RECT 150.825 -110.195 150.925 -109.27 ;
      RECT 150.265 -110.195 150.365 -109.27 ;
      RECT 148.025 -110.195 148.125 -109.27 ;
      RECT 147.465 -110.195 147.565 -109.27 ;
      RECT 146.025 -110.195 146.125 -109.27 ;
      RECT 145.465 -110.195 145.565 -109.27 ;
      RECT 143.225 -110.195 143.325 -109.27 ;
      RECT 142.665 -110.195 142.765 -109.27 ;
      RECT 141.225 -110.195 141.325 -109.27 ;
      RECT 140.665 -110.195 140.765 -109.27 ;
      RECT 138.425 -110.195 138.525 -109.27 ;
      RECT 137.865 -110.195 137.965 -109.27 ;
      RECT 136.425 -110.195 136.525 -109.27 ;
      RECT 135.865 -110.195 135.965 -109.27 ;
      RECT 133.625 -110.195 133.725 -109.27 ;
      RECT 133.065 -110.195 133.165 -109.27 ;
      RECT 131.625 -110.195 131.725 -109.27 ;
      RECT 131.065 -110.195 131.165 -109.27 ;
      RECT 128.825 -110.195 128.925 -109.27 ;
      RECT 128.265 -110.195 128.365 -109.27 ;
      RECT 126.825 -110.195 126.925 -109.27 ;
      RECT 126.265 -110.195 126.365 -109.27 ;
      RECT 124.025 -110.195 124.125 -109.27 ;
      RECT 123.465 -110.195 123.565 -109.27 ;
      RECT 122.025 -110.195 122.125 -109.27 ;
      RECT 121.465 -110.195 121.565 -109.27 ;
      RECT 119.225 -110.195 119.325 -109.27 ;
      RECT 118.665 -110.195 118.765 -109.27 ;
      RECT 117.225 -110.195 117.325 -109.27 ;
      RECT 116.665 -110.195 116.765 -109.27 ;
      RECT 114.425 -110.195 114.525 -109.27 ;
      RECT 113.865 -110.195 113.965 -109.27 ;
      RECT 112.425 -110.195 112.525 -109.27 ;
      RECT 111.865 -110.195 111.965 -109.27 ;
      RECT 109.625 -110.195 109.725 -109.27 ;
      RECT 109.065 -110.195 109.165 -109.27 ;
      RECT 107.625 -110.195 107.725 -109.27 ;
      RECT 107.065 -110.195 107.165 -109.27 ;
      RECT 104.825 -110.195 104.925 -109.27 ;
      RECT 104.265 -110.195 104.365 -109.27 ;
      RECT 102.825 -110.195 102.925 -109.27 ;
      RECT 102.265 -110.195 102.365 -109.27 ;
      RECT 100.025 -110.195 100.125 -109.27 ;
      RECT 99.465 -110.195 99.565 -109.27 ;
      RECT 98.025 -110.195 98.125 -109.27 ;
      RECT 97.465 -110.195 97.565 -109.27 ;
      RECT 95.225 -110.195 95.325 -109.27 ;
      RECT 94.665 -110.195 94.765 -109.27 ;
      RECT 93.225 -110.195 93.325 -109.27 ;
      RECT 92.665 -110.195 92.765 -109.27 ;
      RECT 90.425 -110.195 90.525 -109.27 ;
      RECT 89.865 -110.195 89.965 -109.27 ;
      RECT 88.425 -110.195 88.525 -109.27 ;
      RECT 87.865 -110.195 87.965 -109.27 ;
      RECT 85.625 -110.195 85.725 -109.27 ;
      RECT 85.065 -110.195 85.165 -109.27 ;
      RECT 83.625 -110.195 83.725 -109.27 ;
      RECT 83.065 -110.195 83.165 -109.27 ;
      RECT 80.825 -110.195 80.925 -109.27 ;
      RECT 80.265 -110.195 80.365 -109.27 ;
      RECT 78.825 -110.195 78.925 -109.27 ;
      RECT 78.265 -110.195 78.365 -109.27 ;
      RECT 76.025 -110.195 76.125 -109.27 ;
      RECT 75.465 -110.195 75.565 -109.27 ;
      RECT 74.025 -110.195 74.125 -109.27 ;
      RECT 73.465 -110.195 73.565 -109.27 ;
      RECT 71.225 -110.195 71.325 -109.27 ;
      RECT 70.665 -110.195 70.765 -109.27 ;
      RECT 69.225 -110.195 69.325 -109.27 ;
      RECT 68.665 -110.195 68.765 -109.27 ;
      RECT 66.425 -110.195 66.525 -109.27 ;
      RECT 65.865 -110.195 65.965 -109.27 ;
      RECT 64.425 -110.195 64.525 -109.27 ;
      RECT 63.865 -110.195 63.965 -109.27 ;
      RECT 61.625 -110.195 61.725 -109.27 ;
      RECT 61.065 -110.195 61.165 -109.27 ;
      RECT 59.625 -110.195 59.725 -109.27 ;
      RECT 59.065 -110.195 59.165 -109.27 ;
      RECT 56.825 -110.195 56.925 -109.27 ;
      RECT 56.265 -110.195 56.365 -109.27 ;
      RECT 54.825 -110.195 54.925 -109.27 ;
      RECT 54.265 -110.195 54.365 -109.27 ;
      RECT 52.025 -110.195 52.125 -109.27 ;
      RECT 51.465 -110.195 51.565 -109.27 ;
      RECT 50.025 -110.195 50.125 -109.27 ;
      RECT 49.465 -110.195 49.565 -109.27 ;
      RECT 47.225 -110.195 47.325 -109.27 ;
      RECT 46.665 -110.195 46.765 -109.27 ;
      RECT 45.225 -110.195 45.325 -109.27 ;
      RECT 44.665 -110.195 44.765 -109.27 ;
      RECT 42.425 -110.195 42.525 -109.27 ;
      RECT 41.865 -110.195 41.965 -109.27 ;
      RECT 40.425 -110.195 40.525 -109.27 ;
      RECT 39.865 -110.195 39.965 -109.27 ;
      RECT 37.625 -110.195 37.725 -109.27 ;
      RECT 37.065 -110.195 37.165 -109.27 ;
      RECT 35.625 -110.195 35.725 -109.27 ;
      RECT 35.065 -110.195 35.165 -109.27 ;
      RECT 32.825 -110.195 32.925 -109.27 ;
      RECT 32.265 -110.195 32.365 -109.27 ;
      RECT 30.825 -110.195 30.925 -109.27 ;
      RECT 30.265 -110.195 30.365 -109.27 ;
      RECT 28.025 -110.195 28.125 -109.27 ;
      RECT 27.465 -110.195 27.565 -109.27 ;
      RECT 26.025 -110.195 26.125 -109.27 ;
      RECT 25.465 -110.195 25.565 -109.27 ;
      RECT 23.225 -110.195 23.325 -109.27 ;
      RECT 22.665 -110.195 22.765 -109.27 ;
      RECT 21.225 -110.195 21.325 -109.27 ;
      RECT 20.665 -110.195 20.765 -109.27 ;
      RECT 18.425 -110.195 18.525 -109.27 ;
      RECT 17.865 -110.195 17.965 -109.27 ;
      RECT 16.425 -110.195 16.525 -109.27 ;
      RECT 15.865 -110.195 15.965 -109.27 ;
      RECT 13.625 -110.195 13.725 -109.27 ;
      RECT 13.065 -110.195 13.165 -109.27 ;
      RECT 11.625 -110.195 11.725 -109.27 ;
      RECT 11.065 -110.195 11.165 -109.27 ;
      RECT 8.825 -110.195 8.925 -109.27 ;
      RECT 8.265 -110.195 8.365 -109.27 ;
      RECT 6.825 -110.195 6.925 -109.27 ;
      RECT 6.265 -110.195 6.365 -109.27 ;
      RECT 4.025 -110.195 4.125 -109.27 ;
      RECT 3.465 -110.195 3.565 -109.27 ;
      RECT 2.025 -110.195 2.125 -109.27 ;
      RECT 1.465 -110.195 1.565 -109.27 ;
      RECT -0.04 -110.195 158.465 -109.835 ;
      RECT 153.155 -110.765 153.255 -109.835 ;
      RECT 152.595 -110.765 152.695 -109.835 ;
      RECT 151.445 -110.75 151.545 -109.835 ;
      RECT 151.135 -110.765 151.235 -109.835 ;
      RECT 150.575 -110.765 150.675 -109.835 ;
      RECT 149.39 -110.765 149.565 -109.835 ;
      RECT 148.835 -110.73 148.935 -109.835 ;
      RECT 148.355 -110.765 148.455 -109.835 ;
      RECT 147.795 -110.765 147.895 -109.835 ;
      RECT 146.645 -110.75 146.745 -109.835 ;
      RECT 146.335 -110.765 146.435 -109.835 ;
      RECT 145.775 -110.765 145.875 -109.835 ;
      RECT 144.59 -110.765 144.765 -109.835 ;
      RECT 144.035 -110.73 144.135 -109.835 ;
      RECT 143.555 -110.765 143.655 -109.835 ;
      RECT 142.995 -110.765 143.095 -109.835 ;
      RECT 141.845 -110.75 141.945 -109.835 ;
      RECT 141.535 -110.765 141.635 -109.835 ;
      RECT 140.975 -110.765 141.075 -109.835 ;
      RECT 139.79 -110.765 139.965 -109.835 ;
      RECT 139.235 -110.73 139.335 -109.835 ;
      RECT 138.755 -110.765 138.855 -109.835 ;
      RECT 138.195 -110.765 138.295 -109.835 ;
      RECT 137.045 -110.75 137.145 -109.835 ;
      RECT 136.735 -110.765 136.835 -109.835 ;
      RECT 136.175 -110.765 136.275 -109.835 ;
      RECT 134.99 -110.765 135.165 -109.835 ;
      RECT 134.435 -110.73 134.535 -109.835 ;
      RECT 133.955 -110.765 134.055 -109.835 ;
      RECT 133.395 -110.765 133.495 -109.835 ;
      RECT 132.245 -110.75 132.345 -109.835 ;
      RECT 131.935 -110.765 132.035 -109.835 ;
      RECT 131.375 -110.765 131.475 -109.835 ;
      RECT 130.19 -110.765 130.365 -109.835 ;
      RECT 129.635 -110.73 129.735 -109.835 ;
      RECT 129.155 -110.765 129.255 -109.835 ;
      RECT 128.595 -110.765 128.695 -109.835 ;
      RECT 127.445 -110.75 127.545 -109.835 ;
      RECT 127.135 -110.765 127.235 -109.835 ;
      RECT 126.575 -110.765 126.675 -109.835 ;
      RECT 125.39 -110.765 125.565 -109.835 ;
      RECT 124.835 -110.73 124.935 -109.835 ;
      RECT 124.355 -110.765 124.455 -109.835 ;
      RECT 123.795 -110.765 123.895 -109.835 ;
      RECT 122.645 -110.75 122.745 -109.835 ;
      RECT 122.335 -110.765 122.435 -109.835 ;
      RECT 121.775 -110.765 121.875 -109.835 ;
      RECT 120.59 -110.765 120.765 -109.835 ;
      RECT 120.035 -110.73 120.135 -109.835 ;
      RECT 119.555 -110.765 119.655 -109.835 ;
      RECT 118.995 -110.765 119.095 -109.835 ;
      RECT 117.845 -110.75 117.945 -109.835 ;
      RECT 117.535 -110.765 117.635 -109.835 ;
      RECT 116.975 -110.765 117.075 -109.835 ;
      RECT 115.79 -110.765 115.965 -109.835 ;
      RECT 115.235 -110.73 115.335 -109.835 ;
      RECT 114.755 -110.765 114.855 -109.835 ;
      RECT 114.195 -110.765 114.295 -109.835 ;
      RECT 113.045 -110.75 113.145 -109.835 ;
      RECT 112.735 -110.765 112.835 -109.835 ;
      RECT 112.175 -110.765 112.275 -109.835 ;
      RECT 110.99 -110.765 111.165 -109.835 ;
      RECT 110.435 -110.73 110.535 -109.835 ;
      RECT 109.955 -110.765 110.055 -109.835 ;
      RECT 109.395 -110.765 109.495 -109.835 ;
      RECT 108.245 -110.75 108.345 -109.835 ;
      RECT 107.935 -110.765 108.035 -109.835 ;
      RECT 107.375 -110.765 107.475 -109.835 ;
      RECT 106.19 -110.765 106.365 -109.835 ;
      RECT 105.635 -110.73 105.735 -109.835 ;
      RECT 105.155 -110.765 105.255 -109.835 ;
      RECT 104.595 -110.765 104.695 -109.835 ;
      RECT 103.445 -110.75 103.545 -109.835 ;
      RECT 103.135 -110.765 103.235 -109.835 ;
      RECT 102.575 -110.765 102.675 -109.835 ;
      RECT 101.39 -110.765 101.565 -109.835 ;
      RECT 100.835 -110.73 100.935 -109.835 ;
      RECT 100.355 -110.765 100.455 -109.835 ;
      RECT 99.795 -110.765 99.895 -109.835 ;
      RECT 98.645 -110.75 98.745 -109.835 ;
      RECT 98.335 -110.765 98.435 -109.835 ;
      RECT 97.775 -110.765 97.875 -109.835 ;
      RECT 96.59 -110.765 96.765 -109.835 ;
      RECT 96.035 -110.73 96.135 -109.835 ;
      RECT 95.555 -110.765 95.655 -109.835 ;
      RECT 94.995 -110.765 95.095 -109.835 ;
      RECT 93.845 -110.75 93.945 -109.835 ;
      RECT 93.535 -110.765 93.635 -109.835 ;
      RECT 92.975 -110.765 93.075 -109.835 ;
      RECT 91.79 -110.765 91.965 -109.835 ;
      RECT 91.235 -110.73 91.335 -109.835 ;
      RECT 90.755 -110.765 90.855 -109.835 ;
      RECT 90.195 -110.765 90.295 -109.835 ;
      RECT 89.045 -110.75 89.145 -109.835 ;
      RECT 88.735 -110.765 88.835 -109.835 ;
      RECT 88.175 -110.765 88.275 -109.835 ;
      RECT 86.99 -110.765 87.165 -109.835 ;
      RECT 86.435 -110.73 86.535 -109.835 ;
      RECT 85.955 -110.765 86.055 -109.835 ;
      RECT 85.395 -110.765 85.495 -109.835 ;
      RECT 84.245 -110.75 84.345 -109.835 ;
      RECT 83.935 -110.765 84.035 -109.835 ;
      RECT 83.375 -110.765 83.475 -109.835 ;
      RECT 82.19 -110.765 82.365 -109.835 ;
      RECT 81.635 -110.73 81.735 -109.835 ;
      RECT 81.155 -110.765 81.255 -109.835 ;
      RECT 80.595 -110.765 80.695 -109.835 ;
      RECT 79.445 -110.75 79.545 -109.835 ;
      RECT 79.135 -110.765 79.235 -109.835 ;
      RECT 78.575 -110.765 78.675 -109.835 ;
      RECT 77.39 -110.765 77.565 -109.835 ;
      RECT 76.835 -110.73 76.935 -109.835 ;
      RECT 76.355 -110.765 76.455 -109.835 ;
      RECT 75.795 -110.765 75.895 -109.835 ;
      RECT 74.645 -110.75 74.745 -109.835 ;
      RECT 74.335 -110.765 74.435 -109.835 ;
      RECT 73.775 -110.765 73.875 -109.835 ;
      RECT 72.59 -110.765 72.765 -109.835 ;
      RECT 72.035 -110.73 72.135 -109.835 ;
      RECT 71.555 -110.765 71.655 -109.835 ;
      RECT 70.995 -110.765 71.095 -109.835 ;
      RECT 69.845 -110.75 69.945 -109.835 ;
      RECT 69.535 -110.765 69.635 -109.835 ;
      RECT 68.975 -110.765 69.075 -109.835 ;
      RECT 67.79 -110.765 67.965 -109.835 ;
      RECT 67.235 -110.73 67.335 -109.835 ;
      RECT 66.755 -110.765 66.855 -109.835 ;
      RECT 66.195 -110.765 66.295 -109.835 ;
      RECT 65.045 -110.75 65.145 -109.835 ;
      RECT 64.735 -110.765 64.835 -109.835 ;
      RECT 64.175 -110.765 64.275 -109.835 ;
      RECT 62.99 -110.765 63.165 -109.835 ;
      RECT 62.435 -110.73 62.535 -109.835 ;
      RECT 61.955 -110.765 62.055 -109.835 ;
      RECT 61.395 -110.765 61.495 -109.835 ;
      RECT 60.245 -110.75 60.345 -109.835 ;
      RECT 59.935 -110.765 60.035 -109.835 ;
      RECT 59.375 -110.765 59.475 -109.835 ;
      RECT 58.19 -110.765 58.365 -109.835 ;
      RECT 57.635 -110.73 57.735 -109.835 ;
      RECT 57.155 -110.765 57.255 -109.835 ;
      RECT 56.595 -110.765 56.695 -109.835 ;
      RECT 55.445 -110.75 55.545 -109.835 ;
      RECT 55.135 -110.765 55.235 -109.835 ;
      RECT 54.575 -110.765 54.675 -109.835 ;
      RECT 53.39 -110.765 53.565 -109.835 ;
      RECT 52.835 -110.73 52.935 -109.835 ;
      RECT 52.355 -110.765 52.455 -109.835 ;
      RECT 51.795 -110.765 51.895 -109.835 ;
      RECT 50.645 -110.75 50.745 -109.835 ;
      RECT 50.335 -110.765 50.435 -109.835 ;
      RECT 49.775 -110.765 49.875 -109.835 ;
      RECT 48.59 -110.765 48.765 -109.835 ;
      RECT 48.035 -110.73 48.135 -109.835 ;
      RECT 47.555 -110.765 47.655 -109.835 ;
      RECT 46.995 -110.765 47.095 -109.835 ;
      RECT 45.845 -110.75 45.945 -109.835 ;
      RECT 45.535 -110.765 45.635 -109.835 ;
      RECT 44.975 -110.765 45.075 -109.835 ;
      RECT 43.79 -110.765 43.965 -109.835 ;
      RECT 43.235 -110.73 43.335 -109.835 ;
      RECT 42.755 -110.765 42.855 -109.835 ;
      RECT 42.195 -110.765 42.295 -109.835 ;
      RECT 41.045 -110.75 41.145 -109.835 ;
      RECT 40.735 -110.765 40.835 -109.835 ;
      RECT 40.175 -110.765 40.275 -109.835 ;
      RECT 38.99 -110.765 39.165 -109.835 ;
      RECT 38.435 -110.73 38.535 -109.835 ;
      RECT 37.955 -110.765 38.055 -109.835 ;
      RECT 37.395 -110.765 37.495 -109.835 ;
      RECT 36.245 -110.75 36.345 -109.835 ;
      RECT 35.935 -110.765 36.035 -109.835 ;
      RECT 35.375 -110.765 35.475 -109.835 ;
      RECT 34.19 -110.765 34.365 -109.835 ;
      RECT 33.635 -110.73 33.735 -109.835 ;
      RECT 33.155 -110.765 33.255 -109.835 ;
      RECT 32.595 -110.765 32.695 -109.835 ;
      RECT 31.445 -110.75 31.545 -109.835 ;
      RECT 31.135 -110.765 31.235 -109.835 ;
      RECT 30.575 -110.765 30.675 -109.835 ;
      RECT 29.39 -110.765 29.565 -109.835 ;
      RECT 28.835 -110.73 28.935 -109.835 ;
      RECT 28.355 -110.765 28.455 -109.835 ;
      RECT 27.795 -110.765 27.895 -109.835 ;
      RECT 26.645 -110.75 26.745 -109.835 ;
      RECT 26.335 -110.765 26.435 -109.835 ;
      RECT 25.775 -110.765 25.875 -109.835 ;
      RECT 24.59 -110.765 24.765 -109.835 ;
      RECT 24.035 -110.73 24.135 -109.835 ;
      RECT 23.555 -110.765 23.655 -109.835 ;
      RECT 22.995 -110.765 23.095 -109.835 ;
      RECT 21.845 -110.75 21.945 -109.835 ;
      RECT 21.535 -110.765 21.635 -109.835 ;
      RECT 20.975 -110.765 21.075 -109.835 ;
      RECT 19.79 -110.765 19.965 -109.835 ;
      RECT 19.235 -110.73 19.335 -109.835 ;
      RECT 18.755 -110.765 18.855 -109.835 ;
      RECT 18.195 -110.765 18.295 -109.835 ;
      RECT 17.045 -110.75 17.145 -109.835 ;
      RECT 16.735 -110.765 16.835 -109.835 ;
      RECT 16.175 -110.765 16.275 -109.835 ;
      RECT 14.99 -110.765 15.165 -109.835 ;
      RECT 14.435 -110.73 14.535 -109.835 ;
      RECT 13.955 -110.765 14.055 -109.835 ;
      RECT 13.395 -110.765 13.495 -109.835 ;
      RECT 12.245 -110.75 12.345 -109.835 ;
      RECT 11.935 -110.765 12.035 -109.835 ;
      RECT 11.375 -110.765 11.475 -109.835 ;
      RECT 10.19 -110.765 10.365 -109.835 ;
      RECT 9.635 -110.73 9.735 -109.835 ;
      RECT 9.155 -110.765 9.255 -109.835 ;
      RECT 8.595 -110.765 8.695 -109.835 ;
      RECT 7.445 -110.75 7.545 -109.835 ;
      RECT 7.135 -110.765 7.235 -109.835 ;
      RECT 6.575 -110.765 6.675 -109.835 ;
      RECT 5.39 -110.765 5.565 -109.835 ;
      RECT 4.835 -110.73 4.935 -109.835 ;
      RECT 4.355 -110.765 4.455 -109.835 ;
      RECT 3.795 -110.765 3.895 -109.835 ;
      RECT 2.645 -110.75 2.745 -109.835 ;
      RECT 2.335 -110.765 2.435 -109.835 ;
      RECT 1.775 -110.765 1.875 -109.835 ;
      RECT 0.59 -110.765 0.765 -109.835 ;
      RECT 0.035 -110.73 0.135 -109.835 ;
      RECT 153.155 -112.825 153.255 -111.775 ;
      RECT 152.595 -112.825 152.695 -111.775 ;
      RECT 152.005 -112.825 152.105 -111.775 ;
      RECT 151.445 -112.825 151.545 -111.775 ;
      RECT 151.135 -112.825 151.235 -111.775 ;
      RECT 150.575 -112.825 150.675 -111.775 ;
      RECT 149.985 -112.825 150.085 -111.775 ;
      RECT 149.425 -112.825 149.525 -111.775 ;
      RECT 148.835 -112.825 148.935 -111.775 ;
      RECT 148.355 -112.825 148.455 -111.775 ;
      RECT 147.795 -112.825 147.895 -111.775 ;
      RECT 147.205 -112.825 147.305 -111.775 ;
      RECT 146.645 -112.825 146.745 -111.775 ;
      RECT 146.335 -112.825 146.435 -111.775 ;
      RECT 145.775 -112.825 145.875 -111.775 ;
      RECT 145.185 -112.825 145.285 -111.775 ;
      RECT 144.625 -112.825 144.725 -111.775 ;
      RECT 144.035 -112.825 144.135 -111.775 ;
      RECT 143.555 -112.825 143.655 -111.775 ;
      RECT 142.995 -112.825 143.095 -111.775 ;
      RECT 142.405 -112.825 142.505 -111.775 ;
      RECT 141.845 -112.825 141.945 -111.775 ;
      RECT 141.535 -112.825 141.635 -111.775 ;
      RECT 140.975 -112.825 141.075 -111.775 ;
      RECT 140.385 -112.825 140.485 -111.775 ;
      RECT 139.825 -112.825 139.925 -111.775 ;
      RECT 139.235 -112.825 139.335 -111.775 ;
      RECT 138.755 -112.825 138.855 -111.775 ;
      RECT 138.195 -112.825 138.295 -111.775 ;
      RECT 137.605 -112.825 137.705 -111.775 ;
      RECT 137.045 -112.825 137.145 -111.775 ;
      RECT 136.735 -112.825 136.835 -111.775 ;
      RECT 136.175 -112.825 136.275 -111.775 ;
      RECT 135.585 -112.825 135.685 -111.775 ;
      RECT 135.025 -112.825 135.125 -111.775 ;
      RECT 134.435 -112.825 134.535 -111.775 ;
      RECT 133.955 -112.825 134.055 -111.775 ;
      RECT 133.395 -112.825 133.495 -111.775 ;
      RECT 132.805 -112.825 132.905 -111.775 ;
      RECT 132.245 -112.825 132.345 -111.775 ;
      RECT 131.935 -112.825 132.035 -111.775 ;
      RECT 131.375 -112.825 131.475 -111.775 ;
      RECT 130.785 -112.825 130.885 -111.775 ;
      RECT 130.225 -112.825 130.325 -111.775 ;
      RECT 129.635 -112.825 129.735 -111.775 ;
      RECT 129.155 -112.825 129.255 -111.775 ;
      RECT 128.595 -112.825 128.695 -111.775 ;
      RECT 128.005 -112.825 128.105 -111.775 ;
      RECT 127.445 -112.825 127.545 -111.775 ;
      RECT 127.135 -112.825 127.235 -111.775 ;
      RECT 126.575 -112.825 126.675 -111.775 ;
      RECT 125.985 -112.825 126.085 -111.775 ;
      RECT 125.425 -112.825 125.525 -111.775 ;
      RECT 124.835 -112.825 124.935 -111.775 ;
      RECT 124.355 -112.825 124.455 -111.775 ;
      RECT 123.795 -112.825 123.895 -111.775 ;
      RECT 123.205 -112.825 123.305 -111.775 ;
      RECT 122.645 -112.825 122.745 -111.775 ;
      RECT 122.335 -112.825 122.435 -111.775 ;
      RECT 121.775 -112.825 121.875 -111.775 ;
      RECT 121.185 -112.825 121.285 -111.775 ;
      RECT 120.625 -112.825 120.725 -111.775 ;
      RECT 120.035 -112.825 120.135 -111.775 ;
      RECT 119.555 -112.825 119.655 -111.775 ;
      RECT 118.995 -112.825 119.095 -111.775 ;
      RECT 118.405 -112.825 118.505 -111.775 ;
      RECT 117.845 -112.825 117.945 -111.775 ;
      RECT 117.535 -112.825 117.635 -111.775 ;
      RECT 116.975 -112.825 117.075 -111.775 ;
      RECT 116.385 -112.825 116.485 -111.775 ;
      RECT 115.825 -112.825 115.925 -111.775 ;
      RECT 115.235 -112.825 115.335 -111.775 ;
      RECT 114.755 -112.825 114.855 -111.775 ;
      RECT 114.195 -112.825 114.295 -111.775 ;
      RECT 113.605 -112.825 113.705 -111.775 ;
      RECT 113.045 -112.825 113.145 -111.775 ;
      RECT 112.735 -112.825 112.835 -111.775 ;
      RECT 112.175 -112.825 112.275 -111.775 ;
      RECT 111.585 -112.825 111.685 -111.775 ;
      RECT 111.025 -112.825 111.125 -111.775 ;
      RECT 110.435 -112.825 110.535 -111.775 ;
      RECT 109.955 -112.825 110.055 -111.775 ;
      RECT 109.395 -112.825 109.495 -111.775 ;
      RECT 108.805 -112.825 108.905 -111.775 ;
      RECT 108.245 -112.825 108.345 -111.775 ;
      RECT 107.935 -112.825 108.035 -111.775 ;
      RECT 107.375 -112.825 107.475 -111.775 ;
      RECT 106.785 -112.825 106.885 -111.775 ;
      RECT 106.225 -112.825 106.325 -111.775 ;
      RECT 105.635 -112.825 105.735 -111.775 ;
      RECT 105.155 -112.825 105.255 -111.775 ;
      RECT 104.595 -112.825 104.695 -111.775 ;
      RECT 104.005 -112.825 104.105 -111.775 ;
      RECT 103.445 -112.825 103.545 -111.775 ;
      RECT 103.135 -112.825 103.235 -111.775 ;
      RECT 102.575 -112.825 102.675 -111.775 ;
      RECT 101.985 -112.825 102.085 -111.775 ;
      RECT 101.425 -112.825 101.525 -111.775 ;
      RECT 100.835 -112.825 100.935 -111.775 ;
      RECT 100.355 -112.825 100.455 -111.775 ;
      RECT 99.795 -112.825 99.895 -111.775 ;
      RECT 99.205 -112.825 99.305 -111.775 ;
      RECT 98.645 -112.825 98.745 -111.775 ;
      RECT 98.335 -112.825 98.435 -111.775 ;
      RECT 97.775 -112.825 97.875 -111.775 ;
      RECT 97.185 -112.825 97.285 -111.775 ;
      RECT 96.625 -112.825 96.725 -111.775 ;
      RECT 96.035 -112.825 96.135 -111.775 ;
      RECT 95.555 -112.825 95.655 -111.775 ;
      RECT 94.995 -112.825 95.095 -111.775 ;
      RECT 94.405 -112.825 94.505 -111.775 ;
      RECT 93.845 -112.825 93.945 -111.775 ;
      RECT 93.535 -112.825 93.635 -111.775 ;
      RECT 92.975 -112.825 93.075 -111.775 ;
      RECT 92.385 -112.825 92.485 -111.775 ;
      RECT 91.825 -112.825 91.925 -111.775 ;
      RECT 91.235 -112.825 91.335 -111.775 ;
      RECT 90.755 -112.825 90.855 -111.775 ;
      RECT 90.195 -112.825 90.295 -111.775 ;
      RECT 89.605 -112.825 89.705 -111.775 ;
      RECT 89.045 -112.825 89.145 -111.775 ;
      RECT 88.735 -112.825 88.835 -111.775 ;
      RECT 88.175 -112.825 88.275 -111.775 ;
      RECT 87.585 -112.825 87.685 -111.775 ;
      RECT 87.025 -112.825 87.125 -111.775 ;
      RECT 86.435 -112.825 86.535 -111.775 ;
      RECT 85.955 -112.825 86.055 -111.775 ;
      RECT 85.395 -112.825 85.495 -111.775 ;
      RECT 84.805 -112.825 84.905 -111.775 ;
      RECT 84.245 -112.825 84.345 -111.775 ;
      RECT 83.935 -112.825 84.035 -111.775 ;
      RECT 83.375 -112.825 83.475 -111.775 ;
      RECT 82.785 -112.825 82.885 -111.775 ;
      RECT 82.225 -112.825 82.325 -111.775 ;
      RECT 81.635 -112.825 81.735 -111.775 ;
      RECT 81.155 -112.825 81.255 -111.775 ;
      RECT 80.595 -112.825 80.695 -111.775 ;
      RECT 80.005 -112.825 80.105 -111.775 ;
      RECT 79.445 -112.825 79.545 -111.775 ;
      RECT 79.135 -112.825 79.235 -111.775 ;
      RECT 78.575 -112.825 78.675 -111.775 ;
      RECT 77.985 -112.825 78.085 -111.775 ;
      RECT 77.425 -112.825 77.525 -111.775 ;
      RECT 76.835 -112.825 76.935 -111.775 ;
      RECT 76.355 -112.825 76.455 -111.775 ;
      RECT 75.795 -112.825 75.895 -111.775 ;
      RECT 75.205 -112.825 75.305 -111.775 ;
      RECT 74.645 -112.825 74.745 -111.775 ;
      RECT 74.335 -112.825 74.435 -111.775 ;
      RECT 73.775 -112.825 73.875 -111.775 ;
      RECT 73.185 -112.825 73.285 -111.775 ;
      RECT 72.625 -112.825 72.725 -111.775 ;
      RECT 72.035 -112.825 72.135 -111.775 ;
      RECT 71.555 -112.825 71.655 -111.775 ;
      RECT 70.995 -112.825 71.095 -111.775 ;
      RECT 70.405 -112.825 70.505 -111.775 ;
      RECT 69.845 -112.825 69.945 -111.775 ;
      RECT 69.535 -112.825 69.635 -111.775 ;
      RECT 68.975 -112.825 69.075 -111.775 ;
      RECT 68.385 -112.825 68.485 -111.775 ;
      RECT 67.825 -112.825 67.925 -111.775 ;
      RECT 67.235 -112.825 67.335 -111.775 ;
      RECT 66.755 -112.825 66.855 -111.775 ;
      RECT 66.195 -112.825 66.295 -111.775 ;
      RECT 65.605 -112.825 65.705 -111.775 ;
      RECT 65.045 -112.825 65.145 -111.775 ;
      RECT 64.735 -112.825 64.835 -111.775 ;
      RECT 64.175 -112.825 64.275 -111.775 ;
      RECT 63.585 -112.825 63.685 -111.775 ;
      RECT 63.025 -112.825 63.125 -111.775 ;
      RECT 62.435 -112.825 62.535 -111.775 ;
      RECT 61.955 -112.825 62.055 -111.775 ;
      RECT 61.395 -112.825 61.495 -111.775 ;
      RECT 60.805 -112.825 60.905 -111.775 ;
      RECT 60.245 -112.825 60.345 -111.775 ;
      RECT 59.935 -112.825 60.035 -111.775 ;
      RECT 59.375 -112.825 59.475 -111.775 ;
      RECT 58.785 -112.825 58.885 -111.775 ;
      RECT 58.225 -112.825 58.325 -111.775 ;
      RECT 57.635 -112.825 57.735 -111.775 ;
      RECT 57.155 -112.825 57.255 -111.775 ;
      RECT 56.595 -112.825 56.695 -111.775 ;
      RECT 56.005 -112.825 56.105 -111.775 ;
      RECT 55.445 -112.825 55.545 -111.775 ;
      RECT 55.135 -112.825 55.235 -111.775 ;
      RECT 54.575 -112.825 54.675 -111.775 ;
      RECT 53.985 -112.825 54.085 -111.775 ;
      RECT 53.425 -112.825 53.525 -111.775 ;
      RECT 52.835 -112.825 52.935 -111.775 ;
      RECT 52.355 -112.825 52.455 -111.775 ;
      RECT 51.795 -112.825 51.895 -111.775 ;
      RECT 51.205 -112.825 51.305 -111.775 ;
      RECT 50.645 -112.825 50.745 -111.775 ;
      RECT 50.335 -112.825 50.435 -111.775 ;
      RECT 49.775 -112.825 49.875 -111.775 ;
      RECT 49.185 -112.825 49.285 -111.775 ;
      RECT 48.625 -112.825 48.725 -111.775 ;
      RECT 48.035 -112.825 48.135 -111.775 ;
      RECT 47.555 -112.825 47.655 -111.775 ;
      RECT 46.995 -112.825 47.095 -111.775 ;
      RECT 46.405 -112.825 46.505 -111.775 ;
      RECT 45.845 -112.825 45.945 -111.775 ;
      RECT 45.535 -112.825 45.635 -111.775 ;
      RECT 44.975 -112.825 45.075 -111.775 ;
      RECT 44.385 -112.825 44.485 -111.775 ;
      RECT 43.825 -112.825 43.925 -111.775 ;
      RECT 43.235 -112.825 43.335 -111.775 ;
      RECT 42.755 -112.825 42.855 -111.775 ;
      RECT 42.195 -112.825 42.295 -111.775 ;
      RECT 41.605 -112.825 41.705 -111.775 ;
      RECT 41.045 -112.825 41.145 -111.775 ;
      RECT 40.735 -112.825 40.835 -111.775 ;
      RECT 40.175 -112.825 40.275 -111.775 ;
      RECT 39.585 -112.825 39.685 -111.775 ;
      RECT 39.025 -112.825 39.125 -111.775 ;
      RECT 38.435 -112.825 38.535 -111.775 ;
      RECT 37.955 -112.825 38.055 -111.775 ;
      RECT 37.395 -112.825 37.495 -111.775 ;
      RECT 36.805 -112.825 36.905 -111.775 ;
      RECT 36.245 -112.825 36.345 -111.775 ;
      RECT 35.935 -112.825 36.035 -111.775 ;
      RECT 35.375 -112.825 35.475 -111.775 ;
      RECT 34.785 -112.825 34.885 -111.775 ;
      RECT 34.225 -112.825 34.325 -111.775 ;
      RECT 33.635 -112.825 33.735 -111.775 ;
      RECT 33.155 -112.825 33.255 -111.775 ;
      RECT 32.595 -112.825 32.695 -111.775 ;
      RECT 32.005 -112.825 32.105 -111.775 ;
      RECT 31.445 -112.825 31.545 -111.775 ;
      RECT 31.135 -112.825 31.235 -111.775 ;
      RECT 30.575 -112.825 30.675 -111.775 ;
      RECT 29.985 -112.825 30.085 -111.775 ;
      RECT 29.425 -112.825 29.525 -111.775 ;
      RECT 28.835 -112.825 28.935 -111.775 ;
      RECT 28.355 -112.825 28.455 -111.775 ;
      RECT 27.795 -112.825 27.895 -111.775 ;
      RECT 27.205 -112.825 27.305 -111.775 ;
      RECT 26.645 -112.825 26.745 -111.775 ;
      RECT 26.335 -112.825 26.435 -111.775 ;
      RECT 25.775 -112.825 25.875 -111.775 ;
      RECT 25.185 -112.825 25.285 -111.775 ;
      RECT 24.625 -112.825 24.725 -111.775 ;
      RECT 24.035 -112.825 24.135 -111.775 ;
      RECT 23.555 -112.825 23.655 -111.775 ;
      RECT 22.995 -112.825 23.095 -111.775 ;
      RECT 22.405 -112.825 22.505 -111.775 ;
      RECT 21.845 -112.825 21.945 -111.775 ;
      RECT 21.535 -112.825 21.635 -111.775 ;
      RECT 20.975 -112.825 21.075 -111.775 ;
      RECT 20.385 -112.825 20.485 -111.775 ;
      RECT 19.825 -112.825 19.925 -111.775 ;
      RECT 19.235 -112.825 19.335 -111.775 ;
      RECT 18.755 -112.825 18.855 -111.775 ;
      RECT 18.195 -112.825 18.295 -111.775 ;
      RECT 17.605 -112.825 17.705 -111.775 ;
      RECT 17.045 -112.825 17.145 -111.775 ;
      RECT 16.735 -112.825 16.835 -111.775 ;
      RECT 16.175 -112.825 16.275 -111.775 ;
      RECT 15.585 -112.825 15.685 -111.775 ;
      RECT 15.025 -112.825 15.125 -111.775 ;
      RECT 14.435 -112.825 14.535 -111.775 ;
      RECT 13.955 -112.825 14.055 -111.775 ;
      RECT 13.395 -112.825 13.495 -111.775 ;
      RECT 12.805 -112.825 12.905 -111.775 ;
      RECT 12.245 -112.825 12.345 -111.775 ;
      RECT 11.935 -112.825 12.035 -111.775 ;
      RECT 11.375 -112.825 11.475 -111.775 ;
      RECT 10.785 -112.825 10.885 -111.775 ;
      RECT 10.225 -112.825 10.325 -111.775 ;
      RECT 9.635 -112.825 9.735 -111.775 ;
      RECT 9.155 -112.825 9.255 -111.775 ;
      RECT 8.595 -112.825 8.695 -111.775 ;
      RECT 8.005 -112.825 8.105 -111.775 ;
      RECT 7.445 -112.825 7.545 -111.775 ;
      RECT 7.135 -112.825 7.235 -111.775 ;
      RECT 6.575 -112.825 6.675 -111.775 ;
      RECT 5.985 -112.825 6.085 -111.775 ;
      RECT 5.425 -112.825 5.525 -111.775 ;
      RECT 4.835 -112.825 4.935 -111.775 ;
      RECT 4.355 -112.825 4.455 -111.775 ;
      RECT 3.795 -112.825 3.895 -111.775 ;
      RECT 3.205 -112.825 3.305 -111.775 ;
      RECT 2.645 -112.825 2.745 -111.775 ;
      RECT 2.335 -112.825 2.435 -111.775 ;
      RECT 1.775 -112.825 1.875 -111.775 ;
      RECT 1.185 -112.825 1.285 -111.775 ;
      RECT 0.625 -112.825 0.725 -111.775 ;
      RECT 0.035 -112.825 0.135 -111.775 ;
      RECT -0.04 -112.825 156.465 -112.465 ;
      RECT 150.98 -113.275 151.08 -112.465 ;
      RECT 150.39 -113.275 150.49 -112.465 ;
      RECT 146.18 -113.275 146.28 -112.465 ;
      RECT 145.59 -113.275 145.69 -112.465 ;
      RECT 141.38 -113.275 141.48 -112.465 ;
      RECT 140.79 -113.275 140.89 -112.465 ;
      RECT 136.58 -113.275 136.68 -112.465 ;
      RECT 135.99 -113.275 136.09 -112.465 ;
      RECT 131.78 -113.275 131.88 -112.465 ;
      RECT 131.19 -113.275 131.29 -112.465 ;
      RECT 126.98 -113.275 127.08 -112.465 ;
      RECT 126.39 -113.275 126.49 -112.465 ;
      RECT 122.18 -113.275 122.28 -112.465 ;
      RECT 121.59 -113.275 121.69 -112.465 ;
      RECT 117.38 -113.275 117.48 -112.465 ;
      RECT 116.79 -113.275 116.89 -112.465 ;
      RECT 112.58 -113.275 112.68 -112.465 ;
      RECT 111.99 -113.275 112.09 -112.465 ;
      RECT 107.78 -113.275 107.88 -112.465 ;
      RECT 107.19 -113.275 107.29 -112.465 ;
      RECT 102.98 -113.275 103.08 -112.465 ;
      RECT 102.39 -113.275 102.49 -112.465 ;
      RECT 98.18 -113.275 98.28 -112.465 ;
      RECT 97.59 -113.275 97.69 -112.465 ;
      RECT 93.38 -113.275 93.48 -112.465 ;
      RECT 92.79 -113.275 92.89 -112.465 ;
      RECT 88.58 -113.275 88.68 -112.465 ;
      RECT 87.99 -113.275 88.09 -112.465 ;
      RECT 83.78 -113.275 83.88 -112.465 ;
      RECT 83.19 -113.275 83.29 -112.465 ;
      RECT 78.98 -113.275 79.08 -112.465 ;
      RECT 78.39 -113.275 78.49 -112.465 ;
      RECT 74.18 -113.275 74.28 -112.465 ;
      RECT 73.59 -113.275 73.69 -112.465 ;
      RECT 69.38 -113.275 69.48 -112.465 ;
      RECT 68.79 -113.275 68.89 -112.465 ;
      RECT 64.58 -113.275 64.68 -112.465 ;
      RECT 63.99 -113.275 64.09 -112.465 ;
      RECT 59.78 -113.275 59.88 -112.465 ;
      RECT 59.19 -113.275 59.29 -112.465 ;
      RECT 54.98 -113.275 55.08 -112.465 ;
      RECT 54.39 -113.275 54.49 -112.465 ;
      RECT 50.18 -113.275 50.28 -112.465 ;
      RECT 49.59 -113.275 49.69 -112.465 ;
      RECT 45.38 -113.275 45.48 -112.465 ;
      RECT 44.79 -113.275 44.89 -112.465 ;
      RECT 40.58 -113.275 40.68 -112.465 ;
      RECT 39.99 -113.275 40.09 -112.465 ;
      RECT 35.78 -113.275 35.88 -112.465 ;
      RECT 35.19 -113.275 35.29 -112.465 ;
      RECT 30.98 -113.275 31.08 -112.465 ;
      RECT 30.39 -113.275 30.49 -112.465 ;
      RECT 26.18 -113.275 26.28 -112.465 ;
      RECT 25.59 -113.275 25.69 -112.465 ;
      RECT 21.38 -113.275 21.48 -112.465 ;
      RECT 20.79 -113.275 20.89 -112.465 ;
      RECT 16.58 -113.275 16.68 -112.465 ;
      RECT 15.99 -113.275 16.09 -112.465 ;
      RECT 11.78 -113.275 11.88 -112.465 ;
      RECT 11.19 -113.275 11.29 -112.465 ;
      RECT 6.98 -113.275 7.08 -112.465 ;
      RECT 6.39 -113.275 6.49 -112.465 ;
      RECT 2.18 -113.275 2.28 -112.465 ;
      RECT 1.59 -113.275 1.69 -112.465 ;
      RECT 153.55 -101.805 153.65 -101.34 ;
      RECT 152.35 -101.805 152.45 -101.34 ;
      RECT 151.15 -101.805 151.25 -101.34 ;
      RECT 149.95 -101.805 150.05 -101.34 ;
      RECT 148.75 -101.805 148.85 -101.34 ;
      RECT 147.55 -101.805 147.65 -101.34 ;
      RECT 146.35 -101.805 146.45 -101.34 ;
      RECT 145.15 -101.805 145.25 -101.34 ;
      RECT 143.95 -101.805 144.05 -101.34 ;
      RECT 142.75 -101.805 142.85 -101.34 ;
      RECT 141.55 -101.805 141.65 -101.34 ;
      RECT 140.35 -101.805 140.45 -101.34 ;
      RECT 139.15 -101.805 139.25 -101.34 ;
      RECT 137.95 -101.805 138.05 -101.34 ;
      RECT 136.75 -101.805 136.85 -101.34 ;
      RECT 135.55 -101.805 135.65 -101.34 ;
      RECT 134.35 -101.805 134.45 -101.34 ;
      RECT 133.15 -101.805 133.25 -101.34 ;
      RECT 131.95 -101.805 132.05 -101.34 ;
      RECT 130.75 -101.805 130.85 -101.34 ;
      RECT 129.55 -101.805 129.65 -101.34 ;
      RECT 128.35 -101.805 128.45 -101.34 ;
      RECT 127.15 -101.805 127.25 -101.34 ;
      RECT 125.95 -101.805 126.05 -101.34 ;
      RECT 124.75 -101.805 124.85 -101.34 ;
      RECT 123.55 -101.805 123.65 -101.34 ;
      RECT 122.35 -101.805 122.45 -101.34 ;
      RECT 121.15 -101.805 121.25 -101.34 ;
      RECT 119.95 -101.805 120.05 -101.34 ;
      RECT 118.75 -101.805 118.85 -101.34 ;
      RECT 117.55 -101.805 117.65 -101.34 ;
      RECT 116.35 -101.805 116.45 -101.34 ;
      RECT 115.15 -101.805 115.25 -101.34 ;
      RECT 113.95 -101.805 114.05 -101.34 ;
      RECT 112.75 -101.805 112.85 -101.34 ;
      RECT 111.55 -101.805 111.65 -101.34 ;
      RECT 110.35 -101.805 110.45 -101.34 ;
      RECT 109.15 -101.805 109.25 -101.34 ;
      RECT 107.95 -101.805 108.05 -101.34 ;
      RECT 106.75 -101.805 106.85 -101.34 ;
      RECT 105.55 -101.805 105.65 -101.34 ;
      RECT 104.35 -101.805 104.45 -101.34 ;
      RECT 103.15 -101.805 103.25 -101.34 ;
      RECT 101.95 -101.805 102.05 -101.34 ;
      RECT 100.75 -101.805 100.85 -101.34 ;
      RECT 99.55 -101.805 99.65 -101.34 ;
      RECT 98.35 -101.805 98.45 -101.34 ;
      RECT 97.15 -101.805 97.25 -101.34 ;
      RECT 95.95 -101.805 96.05 -101.34 ;
      RECT 94.75 -101.805 94.85 -101.34 ;
      RECT 93.55 -101.805 93.65 -101.34 ;
      RECT 92.35 -101.805 92.45 -101.34 ;
      RECT 91.15 -101.805 91.25 -101.34 ;
      RECT 89.95 -101.805 90.05 -101.34 ;
      RECT 88.75 -101.805 88.85 -101.34 ;
      RECT 87.55 -101.805 87.65 -101.34 ;
      RECT 86.35 -101.805 86.45 -101.34 ;
      RECT 85.15 -101.805 85.25 -101.34 ;
      RECT 83.95 -101.805 84.05 -101.34 ;
      RECT 82.75 -101.805 82.85 -101.34 ;
      RECT 81.55 -101.805 81.65 -101.34 ;
      RECT 80.35 -101.805 80.45 -101.34 ;
      RECT 79.15 -101.805 79.25 -101.34 ;
      RECT 77.95 -101.805 78.05 -101.34 ;
      RECT 76.75 -101.805 76.85 -101.34 ;
      RECT 75.55 -101.805 75.65 -101.34 ;
      RECT 74.35 -101.805 74.45 -101.34 ;
      RECT 73.15 -101.805 73.25 -101.34 ;
      RECT 71.95 -101.805 72.05 -101.34 ;
      RECT 70.75 -101.805 70.85 -101.34 ;
      RECT 69.55 -101.805 69.65 -101.34 ;
      RECT 68.35 -101.805 68.45 -101.34 ;
      RECT 67.15 -101.805 67.25 -101.34 ;
      RECT 65.95 -101.805 66.05 -101.34 ;
      RECT 64.75 -101.805 64.85 -101.34 ;
      RECT 63.55 -101.805 63.65 -101.34 ;
      RECT 62.35 -101.805 62.45 -101.34 ;
      RECT 61.15 -101.805 61.25 -101.34 ;
      RECT 59.95 -101.805 60.05 -101.34 ;
      RECT 58.75 -101.805 58.85 -101.34 ;
      RECT 57.55 -101.805 57.65 -101.34 ;
      RECT 56.35 -101.805 56.45 -101.34 ;
      RECT 55.15 -101.805 55.25 -101.34 ;
      RECT 53.95 -101.805 54.05 -101.34 ;
      RECT 52.75 -101.805 52.85 -101.34 ;
      RECT 51.55 -101.805 51.65 -101.34 ;
      RECT 50.35 -101.805 50.45 -101.34 ;
      RECT 49.15 -101.805 49.25 -101.34 ;
      RECT 47.95 -101.805 48.05 -101.34 ;
      RECT 46.75 -101.805 46.85 -101.34 ;
      RECT 45.55 -101.805 45.65 -101.34 ;
      RECT 44.35 -101.805 44.45 -101.34 ;
      RECT 43.15 -101.805 43.25 -101.34 ;
      RECT 41.95 -101.805 42.05 -101.34 ;
      RECT 40.75 -101.805 40.85 -101.34 ;
      RECT 39.55 -101.805 39.65 -101.34 ;
      RECT 38.35 -101.805 38.45 -101.34 ;
      RECT 37.15 -101.805 37.25 -101.34 ;
      RECT 35.95 -101.805 36.05 -101.34 ;
      RECT 34.75 -101.805 34.85 -101.34 ;
      RECT 33.55 -101.805 33.65 -101.34 ;
      RECT 32.35 -101.805 32.45 -101.34 ;
      RECT 31.15 -101.805 31.25 -101.34 ;
      RECT 29.95 -101.805 30.05 -101.34 ;
      RECT 28.75 -101.805 28.85 -101.34 ;
      RECT 27.55 -101.805 27.65 -101.34 ;
      RECT 26.35 -101.805 26.45 -101.34 ;
      RECT 25.15 -101.805 25.25 -101.34 ;
      RECT 23.95 -101.805 24.05 -101.34 ;
      RECT 22.75 -101.805 22.85 -101.34 ;
      RECT 21.55 -101.805 21.65 -101.34 ;
      RECT 20.35 -101.805 20.45 -101.34 ;
      RECT 19.15 -101.805 19.25 -101.34 ;
      RECT 17.95 -101.805 18.05 -101.34 ;
      RECT 16.75 -101.805 16.85 -101.34 ;
      RECT 15.55 -101.805 15.65 -101.34 ;
      RECT 14.35 -101.805 14.45 -101.34 ;
      RECT 13.15 -101.805 13.25 -101.34 ;
      RECT 11.95 -101.805 12.05 -101.34 ;
      RECT 10.75 -101.805 10.85 -101.34 ;
      RECT 9.55 -101.805 9.65 -101.34 ;
      RECT 8.35 -101.805 8.45 -101.34 ;
      RECT 7.15 -101.805 7.25 -101.34 ;
      RECT 5.95 -101.805 6.05 -101.34 ;
      RECT 4.75 -101.805 4.85 -101.34 ;
      RECT 3.55 -101.805 3.65 -101.34 ;
      RECT 2.35 -101.805 2.45 -101.34 ;
      RECT 1.15 -101.805 1.25 -101.34 ;
      RECT -0.05 -101.805 0.05 -101.34 ;
      RECT -0.105 -101.805 156.465 -101.685 ;
      RECT 153.55 -98.92 153.65 -98.11 ;
      RECT 152.35 -98.92 152.45 -98.11 ;
      RECT 151.15 -98.92 151.25 -98.11 ;
      RECT 149.95 -98.92 150.05 -98.11 ;
      RECT 148.75 -98.92 148.85 -98.11 ;
      RECT 147.55 -98.92 147.65 -98.11 ;
      RECT 146.35 -98.92 146.45 -98.11 ;
      RECT 145.15 -98.92 145.25 -98.11 ;
      RECT 143.95 -98.92 144.05 -98.11 ;
      RECT 142.75 -98.92 142.85 -98.11 ;
      RECT 141.55 -98.92 141.65 -98.11 ;
      RECT 140.35 -98.92 140.45 -98.11 ;
      RECT 139.15 -98.92 139.25 -98.11 ;
      RECT 137.95 -98.92 138.05 -98.11 ;
      RECT 136.75 -98.92 136.85 -98.11 ;
      RECT 135.55 -98.92 135.65 -98.11 ;
      RECT 134.35 -98.92 134.45 -98.11 ;
      RECT 133.15 -98.92 133.25 -98.11 ;
      RECT 131.95 -98.92 132.05 -98.11 ;
      RECT 130.75 -98.92 130.85 -98.11 ;
      RECT 129.55 -98.92 129.65 -98.11 ;
      RECT 128.35 -98.92 128.45 -98.11 ;
      RECT 127.15 -98.92 127.25 -98.11 ;
      RECT 125.95 -98.92 126.05 -98.11 ;
      RECT 124.75 -98.92 124.85 -98.11 ;
      RECT 123.55 -98.92 123.65 -98.11 ;
      RECT 122.35 -98.92 122.45 -98.11 ;
      RECT 121.15 -98.92 121.25 -98.11 ;
      RECT 119.95 -98.92 120.05 -98.11 ;
      RECT 118.75 -98.92 118.85 -98.11 ;
      RECT 117.55 -98.92 117.65 -98.11 ;
      RECT 116.35 -98.92 116.45 -98.11 ;
      RECT 115.15 -98.92 115.25 -98.11 ;
      RECT 113.95 -98.92 114.05 -98.11 ;
      RECT 112.75 -98.92 112.85 -98.11 ;
      RECT 111.55 -98.92 111.65 -98.11 ;
      RECT 110.35 -98.92 110.45 -98.11 ;
      RECT 109.15 -98.92 109.25 -98.11 ;
      RECT 107.95 -98.92 108.05 -98.11 ;
      RECT 106.75 -98.92 106.85 -98.11 ;
      RECT 105.55 -98.92 105.65 -98.11 ;
      RECT 104.35 -98.92 104.45 -98.11 ;
      RECT 103.15 -98.92 103.25 -98.11 ;
      RECT 101.95 -98.92 102.05 -98.11 ;
      RECT 100.75 -98.92 100.85 -98.11 ;
      RECT 99.55 -98.92 99.65 -98.11 ;
      RECT 98.35 -98.92 98.45 -98.11 ;
      RECT 97.15 -98.92 97.25 -98.11 ;
      RECT 95.95 -98.92 96.05 -98.11 ;
      RECT 94.75 -98.92 94.85 -98.11 ;
      RECT 93.55 -98.92 93.65 -98.11 ;
      RECT 92.35 -98.92 92.45 -98.11 ;
      RECT 91.15 -98.92 91.25 -98.11 ;
      RECT 89.95 -98.92 90.05 -98.11 ;
      RECT 88.75 -98.92 88.85 -98.11 ;
      RECT 87.55 -98.92 87.65 -98.11 ;
      RECT 86.35 -98.92 86.45 -98.11 ;
      RECT 85.15 -98.92 85.25 -98.11 ;
      RECT 83.95 -98.92 84.05 -98.11 ;
      RECT 82.75 -98.92 82.85 -98.11 ;
      RECT 81.55 -98.92 81.65 -98.11 ;
      RECT 80.35 -98.92 80.45 -98.11 ;
      RECT 79.15 -98.92 79.25 -98.11 ;
      RECT 77.95 -98.92 78.05 -98.11 ;
      RECT 76.75 -98.92 76.85 -98.11 ;
      RECT 75.55 -98.92 75.65 -98.11 ;
      RECT 74.35 -98.92 74.45 -98.11 ;
      RECT 73.15 -98.92 73.25 -98.11 ;
      RECT 71.95 -98.92 72.05 -98.11 ;
      RECT 70.75 -98.92 70.85 -98.11 ;
      RECT 69.55 -98.92 69.65 -98.11 ;
      RECT 68.35 -98.92 68.45 -98.11 ;
      RECT 67.15 -98.92 67.25 -98.11 ;
      RECT 65.95 -98.92 66.05 -98.11 ;
      RECT 64.75 -98.92 64.85 -98.11 ;
      RECT 63.55 -98.92 63.65 -98.11 ;
      RECT 62.35 -98.92 62.45 -98.11 ;
      RECT 61.15 -98.92 61.25 -98.11 ;
      RECT 59.95 -98.92 60.05 -98.11 ;
      RECT 58.75 -98.92 58.85 -98.11 ;
      RECT 57.55 -98.92 57.65 -98.11 ;
      RECT 56.35 -98.92 56.45 -98.11 ;
      RECT 55.15 -98.92 55.25 -98.11 ;
      RECT 53.95 -98.92 54.05 -98.11 ;
      RECT 52.75 -98.92 52.85 -98.11 ;
      RECT 51.55 -98.92 51.65 -98.11 ;
      RECT 50.35 -98.92 50.45 -98.11 ;
      RECT 49.15 -98.92 49.25 -98.11 ;
      RECT 47.95 -98.92 48.05 -98.11 ;
      RECT 46.75 -98.92 46.85 -98.11 ;
      RECT 45.55 -98.92 45.65 -98.11 ;
      RECT 44.35 -98.92 44.45 -98.11 ;
      RECT 43.15 -98.92 43.25 -98.11 ;
      RECT 41.95 -98.92 42.05 -98.11 ;
      RECT 40.75 -98.92 40.85 -98.11 ;
      RECT 39.55 -98.92 39.65 -98.11 ;
      RECT 38.35 -98.92 38.45 -98.11 ;
      RECT 37.15 -98.92 37.25 -98.11 ;
      RECT 35.95 -98.92 36.05 -98.11 ;
      RECT 34.75 -98.92 34.85 -98.11 ;
      RECT 33.55 -98.92 33.65 -98.11 ;
      RECT 32.35 -98.92 32.45 -98.11 ;
      RECT 31.15 -98.92 31.25 -98.11 ;
      RECT 29.95 -98.92 30.05 -98.11 ;
      RECT 28.75 -98.92 28.85 -98.11 ;
      RECT 27.55 -98.92 27.65 -98.11 ;
      RECT 26.35 -98.92 26.45 -98.11 ;
      RECT 25.15 -98.92 25.25 -98.11 ;
      RECT 23.95 -98.92 24.05 -98.11 ;
      RECT 22.75 -98.92 22.85 -98.11 ;
      RECT 21.55 -98.92 21.65 -98.11 ;
      RECT 20.35 -98.92 20.45 -98.11 ;
      RECT 19.15 -98.92 19.25 -98.11 ;
      RECT 17.95 -98.92 18.05 -98.11 ;
      RECT 16.75 -98.92 16.85 -98.11 ;
      RECT 15.55 -98.92 15.65 -98.11 ;
      RECT 14.35 -98.92 14.45 -98.11 ;
      RECT 13.15 -98.92 13.25 -98.11 ;
      RECT 11.95 -98.92 12.05 -98.11 ;
      RECT 10.75 -98.92 10.85 -98.11 ;
      RECT 9.55 -98.92 9.65 -98.11 ;
      RECT 8.35 -98.92 8.45 -98.11 ;
      RECT 7.15 -98.92 7.25 -98.11 ;
      RECT 5.95 -98.92 6.05 -98.11 ;
      RECT 4.75 -98.92 4.85 -98.11 ;
      RECT 3.55 -98.92 3.65 -98.11 ;
      RECT 2.35 -98.92 2.45 -98.11 ;
      RECT 1.15 -98.92 1.25 -98.11 ;
      RECT -0.05 -98.92 0.05 -98.11 ;
      RECT -0.105 -98.575 156.465 -98.455 ;
      RECT 153.55 -95.69 153.65 -94.88 ;
      RECT 152.35 -95.69 152.45 -94.88 ;
      RECT 151.15 -95.69 151.25 -94.88 ;
      RECT 149.95 -95.69 150.05 -94.88 ;
      RECT 148.75 -95.69 148.85 -94.88 ;
      RECT 147.55 -95.69 147.65 -94.88 ;
      RECT 146.35 -95.69 146.45 -94.88 ;
      RECT 145.15 -95.69 145.25 -94.88 ;
      RECT 143.95 -95.69 144.05 -94.88 ;
      RECT 142.75 -95.69 142.85 -94.88 ;
      RECT 141.55 -95.69 141.65 -94.88 ;
      RECT 140.35 -95.69 140.45 -94.88 ;
      RECT 139.15 -95.69 139.25 -94.88 ;
      RECT 137.95 -95.69 138.05 -94.88 ;
      RECT 136.75 -95.69 136.85 -94.88 ;
      RECT 135.55 -95.69 135.65 -94.88 ;
      RECT 134.35 -95.69 134.45 -94.88 ;
      RECT 133.15 -95.69 133.25 -94.88 ;
      RECT 131.95 -95.69 132.05 -94.88 ;
      RECT 130.75 -95.69 130.85 -94.88 ;
      RECT 129.55 -95.69 129.65 -94.88 ;
      RECT 128.35 -95.69 128.45 -94.88 ;
      RECT 127.15 -95.69 127.25 -94.88 ;
      RECT 125.95 -95.69 126.05 -94.88 ;
      RECT 124.75 -95.69 124.85 -94.88 ;
      RECT 123.55 -95.69 123.65 -94.88 ;
      RECT 122.35 -95.69 122.45 -94.88 ;
      RECT 121.15 -95.69 121.25 -94.88 ;
      RECT 119.95 -95.69 120.05 -94.88 ;
      RECT 118.75 -95.69 118.85 -94.88 ;
      RECT 117.55 -95.69 117.65 -94.88 ;
      RECT 116.35 -95.69 116.45 -94.88 ;
      RECT 115.15 -95.69 115.25 -94.88 ;
      RECT 113.95 -95.69 114.05 -94.88 ;
      RECT 112.75 -95.69 112.85 -94.88 ;
      RECT 111.55 -95.69 111.65 -94.88 ;
      RECT 110.35 -95.69 110.45 -94.88 ;
      RECT 109.15 -95.69 109.25 -94.88 ;
      RECT 107.95 -95.69 108.05 -94.88 ;
      RECT 106.75 -95.69 106.85 -94.88 ;
      RECT 105.55 -95.69 105.65 -94.88 ;
      RECT 104.35 -95.69 104.45 -94.88 ;
      RECT 103.15 -95.69 103.25 -94.88 ;
      RECT 101.95 -95.69 102.05 -94.88 ;
      RECT 100.75 -95.69 100.85 -94.88 ;
      RECT 99.55 -95.69 99.65 -94.88 ;
      RECT 98.35 -95.69 98.45 -94.88 ;
      RECT 97.15 -95.69 97.25 -94.88 ;
      RECT 95.95 -95.69 96.05 -94.88 ;
      RECT 94.75 -95.69 94.85 -94.88 ;
      RECT 93.55 -95.69 93.65 -94.88 ;
      RECT 92.35 -95.69 92.45 -94.88 ;
      RECT 91.15 -95.69 91.25 -94.88 ;
      RECT 89.95 -95.69 90.05 -94.88 ;
      RECT 88.75 -95.69 88.85 -94.88 ;
      RECT 87.55 -95.69 87.65 -94.88 ;
      RECT 86.35 -95.69 86.45 -94.88 ;
      RECT 85.15 -95.69 85.25 -94.88 ;
      RECT 83.95 -95.69 84.05 -94.88 ;
      RECT 82.75 -95.69 82.85 -94.88 ;
      RECT 81.55 -95.69 81.65 -94.88 ;
      RECT 80.35 -95.69 80.45 -94.88 ;
      RECT 79.15 -95.69 79.25 -94.88 ;
      RECT 77.95 -95.69 78.05 -94.88 ;
      RECT 76.75 -95.69 76.85 -94.88 ;
      RECT 75.55 -95.69 75.65 -94.88 ;
      RECT 74.35 -95.69 74.45 -94.88 ;
      RECT 73.15 -95.69 73.25 -94.88 ;
      RECT 71.95 -95.69 72.05 -94.88 ;
      RECT 70.75 -95.69 70.85 -94.88 ;
      RECT 69.55 -95.69 69.65 -94.88 ;
      RECT 68.35 -95.69 68.45 -94.88 ;
      RECT 67.15 -95.69 67.25 -94.88 ;
      RECT 65.95 -95.69 66.05 -94.88 ;
      RECT 64.75 -95.69 64.85 -94.88 ;
      RECT 63.55 -95.69 63.65 -94.88 ;
      RECT 62.35 -95.69 62.45 -94.88 ;
      RECT 61.15 -95.69 61.25 -94.88 ;
      RECT 59.95 -95.69 60.05 -94.88 ;
      RECT 58.75 -95.69 58.85 -94.88 ;
      RECT 57.55 -95.69 57.65 -94.88 ;
      RECT 56.35 -95.69 56.45 -94.88 ;
      RECT 55.15 -95.69 55.25 -94.88 ;
      RECT 53.95 -95.69 54.05 -94.88 ;
      RECT 52.75 -95.69 52.85 -94.88 ;
      RECT 51.55 -95.69 51.65 -94.88 ;
      RECT 50.35 -95.69 50.45 -94.88 ;
      RECT 49.15 -95.69 49.25 -94.88 ;
      RECT 47.95 -95.69 48.05 -94.88 ;
      RECT 46.75 -95.69 46.85 -94.88 ;
      RECT 45.55 -95.69 45.65 -94.88 ;
      RECT 44.35 -95.69 44.45 -94.88 ;
      RECT 43.15 -95.69 43.25 -94.88 ;
      RECT 41.95 -95.69 42.05 -94.88 ;
      RECT 40.75 -95.69 40.85 -94.88 ;
      RECT 39.55 -95.69 39.65 -94.88 ;
      RECT 38.35 -95.69 38.45 -94.88 ;
      RECT 37.15 -95.69 37.25 -94.88 ;
      RECT 35.95 -95.69 36.05 -94.88 ;
      RECT 34.75 -95.69 34.85 -94.88 ;
      RECT 33.55 -95.69 33.65 -94.88 ;
      RECT 32.35 -95.69 32.45 -94.88 ;
      RECT 31.15 -95.69 31.25 -94.88 ;
      RECT 29.95 -95.69 30.05 -94.88 ;
      RECT 28.75 -95.69 28.85 -94.88 ;
      RECT 27.55 -95.69 27.65 -94.88 ;
      RECT 26.35 -95.69 26.45 -94.88 ;
      RECT 25.15 -95.69 25.25 -94.88 ;
      RECT 23.95 -95.69 24.05 -94.88 ;
      RECT 22.75 -95.69 22.85 -94.88 ;
      RECT 21.55 -95.69 21.65 -94.88 ;
      RECT 20.35 -95.69 20.45 -94.88 ;
      RECT 19.15 -95.69 19.25 -94.88 ;
      RECT 17.95 -95.69 18.05 -94.88 ;
      RECT 16.75 -95.69 16.85 -94.88 ;
      RECT 15.55 -95.69 15.65 -94.88 ;
      RECT 14.35 -95.69 14.45 -94.88 ;
      RECT 13.15 -95.69 13.25 -94.88 ;
      RECT 11.95 -95.69 12.05 -94.88 ;
      RECT 10.75 -95.69 10.85 -94.88 ;
      RECT 9.55 -95.69 9.65 -94.88 ;
      RECT 8.35 -95.69 8.45 -94.88 ;
      RECT 7.15 -95.69 7.25 -94.88 ;
      RECT 5.95 -95.69 6.05 -94.88 ;
      RECT 4.75 -95.69 4.85 -94.88 ;
      RECT 3.55 -95.69 3.65 -94.88 ;
      RECT 2.35 -95.69 2.45 -94.88 ;
      RECT 1.15 -95.69 1.25 -94.88 ;
      RECT -0.05 -95.69 0.05 -94.88 ;
      RECT -0.105 -95.345 156.465 -95.225 ;
      RECT 153.55 -92.46 153.65 -91.65 ;
      RECT 152.35 -92.46 152.45 -91.65 ;
      RECT 151.15 -92.46 151.25 -91.65 ;
      RECT 149.95 -92.46 150.05 -91.65 ;
      RECT 148.75 -92.46 148.85 -91.65 ;
      RECT 147.55 -92.46 147.65 -91.65 ;
      RECT 146.35 -92.46 146.45 -91.65 ;
      RECT 145.15 -92.46 145.25 -91.65 ;
      RECT 143.95 -92.46 144.05 -91.65 ;
      RECT 142.75 -92.46 142.85 -91.65 ;
      RECT 141.55 -92.46 141.65 -91.65 ;
      RECT 140.35 -92.46 140.45 -91.65 ;
      RECT 139.15 -92.46 139.25 -91.65 ;
      RECT 137.95 -92.46 138.05 -91.65 ;
      RECT 136.75 -92.46 136.85 -91.65 ;
      RECT 135.55 -92.46 135.65 -91.65 ;
      RECT 134.35 -92.46 134.45 -91.65 ;
      RECT 133.15 -92.46 133.25 -91.65 ;
      RECT 131.95 -92.46 132.05 -91.65 ;
      RECT 130.75 -92.46 130.85 -91.65 ;
      RECT 129.55 -92.46 129.65 -91.65 ;
      RECT 128.35 -92.46 128.45 -91.65 ;
      RECT 127.15 -92.46 127.25 -91.65 ;
      RECT 125.95 -92.46 126.05 -91.65 ;
      RECT 124.75 -92.46 124.85 -91.65 ;
      RECT 123.55 -92.46 123.65 -91.65 ;
      RECT 122.35 -92.46 122.45 -91.65 ;
      RECT 121.15 -92.46 121.25 -91.65 ;
      RECT 119.95 -92.46 120.05 -91.65 ;
      RECT 118.75 -92.46 118.85 -91.65 ;
      RECT 117.55 -92.46 117.65 -91.65 ;
      RECT 116.35 -92.46 116.45 -91.65 ;
      RECT 115.15 -92.46 115.25 -91.65 ;
      RECT 113.95 -92.46 114.05 -91.65 ;
      RECT 112.75 -92.46 112.85 -91.65 ;
      RECT 111.55 -92.46 111.65 -91.65 ;
      RECT 110.35 -92.46 110.45 -91.65 ;
      RECT 109.15 -92.46 109.25 -91.65 ;
      RECT 107.95 -92.46 108.05 -91.65 ;
      RECT 106.75 -92.46 106.85 -91.65 ;
      RECT 105.55 -92.46 105.65 -91.65 ;
      RECT 104.35 -92.46 104.45 -91.65 ;
      RECT 103.15 -92.46 103.25 -91.65 ;
      RECT 101.95 -92.46 102.05 -91.65 ;
      RECT 100.75 -92.46 100.85 -91.65 ;
      RECT 99.55 -92.46 99.65 -91.65 ;
      RECT 98.35 -92.46 98.45 -91.65 ;
      RECT 97.15 -92.46 97.25 -91.65 ;
      RECT 95.95 -92.46 96.05 -91.65 ;
      RECT 94.75 -92.46 94.85 -91.65 ;
      RECT 93.55 -92.46 93.65 -91.65 ;
      RECT 92.35 -92.46 92.45 -91.65 ;
      RECT 91.15 -92.46 91.25 -91.65 ;
      RECT 89.95 -92.46 90.05 -91.65 ;
      RECT 88.75 -92.46 88.85 -91.65 ;
      RECT 87.55 -92.46 87.65 -91.65 ;
      RECT 86.35 -92.46 86.45 -91.65 ;
      RECT 85.15 -92.46 85.25 -91.65 ;
      RECT 83.95 -92.46 84.05 -91.65 ;
      RECT 82.75 -92.46 82.85 -91.65 ;
      RECT 81.55 -92.46 81.65 -91.65 ;
      RECT 80.35 -92.46 80.45 -91.65 ;
      RECT 79.15 -92.46 79.25 -91.65 ;
      RECT 77.95 -92.46 78.05 -91.65 ;
      RECT 76.75 -92.46 76.85 -91.65 ;
      RECT 75.55 -92.46 75.65 -91.65 ;
      RECT 74.35 -92.46 74.45 -91.65 ;
      RECT 73.15 -92.46 73.25 -91.65 ;
      RECT 71.95 -92.46 72.05 -91.65 ;
      RECT 70.75 -92.46 70.85 -91.65 ;
      RECT 69.55 -92.46 69.65 -91.65 ;
      RECT 68.35 -92.46 68.45 -91.65 ;
      RECT 67.15 -92.46 67.25 -91.65 ;
      RECT 65.95 -92.46 66.05 -91.65 ;
      RECT 64.75 -92.46 64.85 -91.65 ;
      RECT 63.55 -92.46 63.65 -91.65 ;
      RECT 62.35 -92.46 62.45 -91.65 ;
      RECT 61.15 -92.46 61.25 -91.65 ;
      RECT 59.95 -92.46 60.05 -91.65 ;
      RECT 58.75 -92.46 58.85 -91.65 ;
      RECT 57.55 -92.46 57.65 -91.65 ;
      RECT 56.35 -92.46 56.45 -91.65 ;
      RECT 55.15 -92.46 55.25 -91.65 ;
      RECT 53.95 -92.46 54.05 -91.65 ;
      RECT 52.75 -92.46 52.85 -91.65 ;
      RECT 51.55 -92.46 51.65 -91.65 ;
      RECT 50.35 -92.46 50.45 -91.65 ;
      RECT 49.15 -92.46 49.25 -91.65 ;
      RECT 47.95 -92.46 48.05 -91.65 ;
      RECT 46.75 -92.46 46.85 -91.65 ;
      RECT 45.55 -92.46 45.65 -91.65 ;
      RECT 44.35 -92.46 44.45 -91.65 ;
      RECT 43.15 -92.46 43.25 -91.65 ;
      RECT 41.95 -92.46 42.05 -91.65 ;
      RECT 40.75 -92.46 40.85 -91.65 ;
      RECT 39.55 -92.46 39.65 -91.65 ;
      RECT 38.35 -92.46 38.45 -91.65 ;
      RECT 37.15 -92.46 37.25 -91.65 ;
      RECT 35.95 -92.46 36.05 -91.65 ;
      RECT 34.75 -92.46 34.85 -91.65 ;
      RECT 33.55 -92.46 33.65 -91.65 ;
      RECT 32.35 -92.46 32.45 -91.65 ;
      RECT 31.15 -92.46 31.25 -91.65 ;
      RECT 29.95 -92.46 30.05 -91.65 ;
      RECT 28.75 -92.46 28.85 -91.65 ;
      RECT 27.55 -92.46 27.65 -91.65 ;
      RECT 26.35 -92.46 26.45 -91.65 ;
      RECT 25.15 -92.46 25.25 -91.65 ;
      RECT 23.95 -92.46 24.05 -91.65 ;
      RECT 22.75 -92.46 22.85 -91.65 ;
      RECT 21.55 -92.46 21.65 -91.65 ;
      RECT 20.35 -92.46 20.45 -91.65 ;
      RECT 19.15 -92.46 19.25 -91.65 ;
      RECT 17.95 -92.46 18.05 -91.65 ;
      RECT 16.75 -92.46 16.85 -91.65 ;
      RECT 15.55 -92.46 15.65 -91.65 ;
      RECT 14.35 -92.46 14.45 -91.65 ;
      RECT 13.15 -92.46 13.25 -91.65 ;
      RECT 11.95 -92.46 12.05 -91.65 ;
      RECT 10.75 -92.46 10.85 -91.65 ;
      RECT 9.55 -92.46 9.65 -91.65 ;
      RECT 8.35 -92.46 8.45 -91.65 ;
      RECT 7.15 -92.46 7.25 -91.65 ;
      RECT 5.95 -92.46 6.05 -91.65 ;
      RECT 4.75 -92.46 4.85 -91.65 ;
      RECT 3.55 -92.46 3.65 -91.65 ;
      RECT 2.35 -92.46 2.45 -91.65 ;
      RECT 1.15 -92.46 1.25 -91.65 ;
      RECT -0.05 -92.46 0.05 -91.65 ;
      RECT -0.105 -92.115 156.465 -91.995 ;
      RECT 153.55 -89.23 153.65 -88.42 ;
      RECT 152.35 -89.23 152.45 -88.42 ;
      RECT 151.15 -89.23 151.25 -88.42 ;
      RECT 149.95 -89.23 150.05 -88.42 ;
      RECT 148.75 -89.23 148.85 -88.42 ;
      RECT 147.55 -89.23 147.65 -88.42 ;
      RECT 146.35 -89.23 146.45 -88.42 ;
      RECT 145.15 -89.23 145.25 -88.42 ;
      RECT 143.95 -89.23 144.05 -88.42 ;
      RECT 142.75 -89.23 142.85 -88.42 ;
      RECT 141.55 -89.23 141.65 -88.42 ;
      RECT 140.35 -89.23 140.45 -88.42 ;
      RECT 139.15 -89.23 139.25 -88.42 ;
      RECT 137.95 -89.23 138.05 -88.42 ;
      RECT 136.75 -89.23 136.85 -88.42 ;
      RECT 135.55 -89.23 135.65 -88.42 ;
      RECT 134.35 -89.23 134.45 -88.42 ;
      RECT 133.15 -89.23 133.25 -88.42 ;
      RECT 131.95 -89.23 132.05 -88.42 ;
      RECT 130.75 -89.23 130.85 -88.42 ;
      RECT 129.55 -89.23 129.65 -88.42 ;
      RECT 128.35 -89.23 128.45 -88.42 ;
      RECT 127.15 -89.23 127.25 -88.42 ;
      RECT 125.95 -89.23 126.05 -88.42 ;
      RECT 124.75 -89.23 124.85 -88.42 ;
      RECT 123.55 -89.23 123.65 -88.42 ;
      RECT 122.35 -89.23 122.45 -88.42 ;
      RECT 121.15 -89.23 121.25 -88.42 ;
      RECT 119.95 -89.23 120.05 -88.42 ;
      RECT 118.75 -89.23 118.85 -88.42 ;
      RECT 117.55 -89.23 117.65 -88.42 ;
      RECT 116.35 -89.23 116.45 -88.42 ;
      RECT 115.15 -89.23 115.25 -88.42 ;
      RECT 113.95 -89.23 114.05 -88.42 ;
      RECT 112.75 -89.23 112.85 -88.42 ;
      RECT 111.55 -89.23 111.65 -88.42 ;
      RECT 110.35 -89.23 110.45 -88.42 ;
      RECT 109.15 -89.23 109.25 -88.42 ;
      RECT 107.95 -89.23 108.05 -88.42 ;
      RECT 106.75 -89.23 106.85 -88.42 ;
      RECT 105.55 -89.23 105.65 -88.42 ;
      RECT 104.35 -89.23 104.45 -88.42 ;
      RECT 103.15 -89.23 103.25 -88.42 ;
      RECT 101.95 -89.23 102.05 -88.42 ;
      RECT 100.75 -89.23 100.85 -88.42 ;
      RECT 99.55 -89.23 99.65 -88.42 ;
      RECT 98.35 -89.23 98.45 -88.42 ;
      RECT 97.15 -89.23 97.25 -88.42 ;
      RECT 95.95 -89.23 96.05 -88.42 ;
      RECT 94.75 -89.23 94.85 -88.42 ;
      RECT 93.55 -89.23 93.65 -88.42 ;
      RECT 92.35 -89.23 92.45 -88.42 ;
      RECT 91.15 -89.23 91.25 -88.42 ;
      RECT 89.95 -89.23 90.05 -88.42 ;
      RECT 88.75 -89.23 88.85 -88.42 ;
      RECT 87.55 -89.23 87.65 -88.42 ;
      RECT 86.35 -89.23 86.45 -88.42 ;
      RECT 85.15 -89.23 85.25 -88.42 ;
      RECT 83.95 -89.23 84.05 -88.42 ;
      RECT 82.75 -89.23 82.85 -88.42 ;
      RECT 81.55 -89.23 81.65 -88.42 ;
      RECT 80.35 -89.23 80.45 -88.42 ;
      RECT 79.15 -89.23 79.25 -88.42 ;
      RECT 77.95 -89.23 78.05 -88.42 ;
      RECT 76.75 -89.23 76.85 -88.42 ;
      RECT 75.55 -89.23 75.65 -88.42 ;
      RECT 74.35 -89.23 74.45 -88.42 ;
      RECT 73.15 -89.23 73.25 -88.42 ;
      RECT 71.95 -89.23 72.05 -88.42 ;
      RECT 70.75 -89.23 70.85 -88.42 ;
      RECT 69.55 -89.23 69.65 -88.42 ;
      RECT 68.35 -89.23 68.45 -88.42 ;
      RECT 67.15 -89.23 67.25 -88.42 ;
      RECT 65.95 -89.23 66.05 -88.42 ;
      RECT 64.75 -89.23 64.85 -88.42 ;
      RECT 63.55 -89.23 63.65 -88.42 ;
      RECT 62.35 -89.23 62.45 -88.42 ;
      RECT 61.15 -89.23 61.25 -88.42 ;
      RECT 59.95 -89.23 60.05 -88.42 ;
      RECT 58.75 -89.23 58.85 -88.42 ;
      RECT 57.55 -89.23 57.65 -88.42 ;
      RECT 56.35 -89.23 56.45 -88.42 ;
      RECT 55.15 -89.23 55.25 -88.42 ;
      RECT 53.95 -89.23 54.05 -88.42 ;
      RECT 52.75 -89.23 52.85 -88.42 ;
      RECT 51.55 -89.23 51.65 -88.42 ;
      RECT 50.35 -89.23 50.45 -88.42 ;
      RECT 49.15 -89.23 49.25 -88.42 ;
      RECT 47.95 -89.23 48.05 -88.42 ;
      RECT 46.75 -89.23 46.85 -88.42 ;
      RECT 45.55 -89.23 45.65 -88.42 ;
      RECT 44.35 -89.23 44.45 -88.42 ;
      RECT 43.15 -89.23 43.25 -88.42 ;
      RECT 41.95 -89.23 42.05 -88.42 ;
      RECT 40.75 -89.23 40.85 -88.42 ;
      RECT 39.55 -89.23 39.65 -88.42 ;
      RECT 38.35 -89.23 38.45 -88.42 ;
      RECT 37.15 -89.23 37.25 -88.42 ;
      RECT 35.95 -89.23 36.05 -88.42 ;
      RECT 34.75 -89.23 34.85 -88.42 ;
      RECT 33.55 -89.23 33.65 -88.42 ;
      RECT 32.35 -89.23 32.45 -88.42 ;
      RECT 31.15 -89.23 31.25 -88.42 ;
      RECT 29.95 -89.23 30.05 -88.42 ;
      RECT 28.75 -89.23 28.85 -88.42 ;
      RECT 27.55 -89.23 27.65 -88.42 ;
      RECT 26.35 -89.23 26.45 -88.42 ;
      RECT 25.15 -89.23 25.25 -88.42 ;
      RECT 23.95 -89.23 24.05 -88.42 ;
      RECT 22.75 -89.23 22.85 -88.42 ;
      RECT 21.55 -89.23 21.65 -88.42 ;
      RECT 20.35 -89.23 20.45 -88.42 ;
      RECT 19.15 -89.23 19.25 -88.42 ;
      RECT 17.95 -89.23 18.05 -88.42 ;
      RECT 16.75 -89.23 16.85 -88.42 ;
      RECT 15.55 -89.23 15.65 -88.42 ;
      RECT 14.35 -89.23 14.45 -88.42 ;
      RECT 13.15 -89.23 13.25 -88.42 ;
      RECT 11.95 -89.23 12.05 -88.42 ;
      RECT 10.75 -89.23 10.85 -88.42 ;
      RECT 9.55 -89.23 9.65 -88.42 ;
      RECT 8.35 -89.23 8.45 -88.42 ;
      RECT 7.15 -89.23 7.25 -88.42 ;
      RECT 5.95 -89.23 6.05 -88.42 ;
      RECT 4.75 -89.23 4.85 -88.42 ;
      RECT 3.55 -89.23 3.65 -88.42 ;
      RECT 2.35 -89.23 2.45 -88.42 ;
      RECT 1.15 -89.23 1.25 -88.42 ;
      RECT -0.05 -89.23 0.05 -88.42 ;
      RECT -0.105 -88.885 156.465 -88.765 ;
      RECT 153.55 -86 153.65 -85.19 ;
      RECT 152.35 -86 152.45 -85.19 ;
      RECT 151.15 -86 151.25 -85.19 ;
      RECT 149.95 -86 150.05 -85.19 ;
      RECT 148.75 -86 148.85 -85.19 ;
      RECT 147.55 -86 147.65 -85.19 ;
      RECT 146.35 -86 146.45 -85.19 ;
      RECT 145.15 -86 145.25 -85.19 ;
      RECT 143.95 -86 144.05 -85.19 ;
      RECT 142.75 -86 142.85 -85.19 ;
      RECT 141.55 -86 141.65 -85.19 ;
      RECT 140.35 -86 140.45 -85.19 ;
      RECT 139.15 -86 139.25 -85.19 ;
      RECT 137.95 -86 138.05 -85.19 ;
      RECT 136.75 -86 136.85 -85.19 ;
      RECT 135.55 -86 135.65 -85.19 ;
      RECT 134.35 -86 134.45 -85.19 ;
      RECT 133.15 -86 133.25 -85.19 ;
      RECT 131.95 -86 132.05 -85.19 ;
      RECT 130.75 -86 130.85 -85.19 ;
      RECT 129.55 -86 129.65 -85.19 ;
      RECT 128.35 -86 128.45 -85.19 ;
      RECT 127.15 -86 127.25 -85.19 ;
      RECT 125.95 -86 126.05 -85.19 ;
      RECT 124.75 -86 124.85 -85.19 ;
      RECT 123.55 -86 123.65 -85.19 ;
      RECT 122.35 -86 122.45 -85.19 ;
      RECT 121.15 -86 121.25 -85.19 ;
      RECT 119.95 -86 120.05 -85.19 ;
      RECT 118.75 -86 118.85 -85.19 ;
      RECT 117.55 -86 117.65 -85.19 ;
      RECT 116.35 -86 116.45 -85.19 ;
      RECT 115.15 -86 115.25 -85.19 ;
      RECT 113.95 -86 114.05 -85.19 ;
      RECT 112.75 -86 112.85 -85.19 ;
      RECT 111.55 -86 111.65 -85.19 ;
      RECT 110.35 -86 110.45 -85.19 ;
      RECT 109.15 -86 109.25 -85.19 ;
      RECT 107.95 -86 108.05 -85.19 ;
      RECT 106.75 -86 106.85 -85.19 ;
      RECT 105.55 -86 105.65 -85.19 ;
      RECT 104.35 -86 104.45 -85.19 ;
      RECT 103.15 -86 103.25 -85.19 ;
      RECT 101.95 -86 102.05 -85.19 ;
      RECT 100.75 -86 100.85 -85.19 ;
      RECT 99.55 -86 99.65 -85.19 ;
      RECT 98.35 -86 98.45 -85.19 ;
      RECT 97.15 -86 97.25 -85.19 ;
      RECT 95.95 -86 96.05 -85.19 ;
      RECT 94.75 -86 94.85 -85.19 ;
      RECT 93.55 -86 93.65 -85.19 ;
      RECT 92.35 -86 92.45 -85.19 ;
      RECT 91.15 -86 91.25 -85.19 ;
      RECT 89.95 -86 90.05 -85.19 ;
      RECT 88.75 -86 88.85 -85.19 ;
      RECT 87.55 -86 87.65 -85.19 ;
      RECT 86.35 -86 86.45 -85.19 ;
      RECT 85.15 -86 85.25 -85.19 ;
      RECT 83.95 -86 84.05 -85.19 ;
      RECT 82.75 -86 82.85 -85.19 ;
      RECT 81.55 -86 81.65 -85.19 ;
      RECT 80.35 -86 80.45 -85.19 ;
      RECT 79.15 -86 79.25 -85.19 ;
      RECT 77.95 -86 78.05 -85.19 ;
      RECT 76.75 -86 76.85 -85.19 ;
      RECT 75.55 -86 75.65 -85.19 ;
      RECT 74.35 -86 74.45 -85.19 ;
      RECT 73.15 -86 73.25 -85.19 ;
      RECT 71.95 -86 72.05 -85.19 ;
      RECT 70.75 -86 70.85 -85.19 ;
      RECT 69.55 -86 69.65 -85.19 ;
      RECT 68.35 -86 68.45 -85.19 ;
      RECT 67.15 -86 67.25 -85.19 ;
      RECT 65.95 -86 66.05 -85.19 ;
      RECT 64.75 -86 64.85 -85.19 ;
      RECT 63.55 -86 63.65 -85.19 ;
      RECT 62.35 -86 62.45 -85.19 ;
      RECT 61.15 -86 61.25 -85.19 ;
      RECT 59.95 -86 60.05 -85.19 ;
      RECT 58.75 -86 58.85 -85.19 ;
      RECT 57.55 -86 57.65 -85.19 ;
      RECT 56.35 -86 56.45 -85.19 ;
      RECT 55.15 -86 55.25 -85.19 ;
      RECT 53.95 -86 54.05 -85.19 ;
      RECT 52.75 -86 52.85 -85.19 ;
      RECT 51.55 -86 51.65 -85.19 ;
      RECT 50.35 -86 50.45 -85.19 ;
      RECT 49.15 -86 49.25 -85.19 ;
      RECT 47.95 -86 48.05 -85.19 ;
      RECT 46.75 -86 46.85 -85.19 ;
      RECT 45.55 -86 45.65 -85.19 ;
      RECT 44.35 -86 44.45 -85.19 ;
      RECT 43.15 -86 43.25 -85.19 ;
      RECT 41.95 -86 42.05 -85.19 ;
      RECT 40.75 -86 40.85 -85.19 ;
      RECT 39.55 -86 39.65 -85.19 ;
      RECT 38.35 -86 38.45 -85.19 ;
      RECT 37.15 -86 37.25 -85.19 ;
      RECT 35.95 -86 36.05 -85.19 ;
      RECT 34.75 -86 34.85 -85.19 ;
      RECT 33.55 -86 33.65 -85.19 ;
      RECT 32.35 -86 32.45 -85.19 ;
      RECT 31.15 -86 31.25 -85.19 ;
      RECT 29.95 -86 30.05 -85.19 ;
      RECT 28.75 -86 28.85 -85.19 ;
      RECT 27.55 -86 27.65 -85.19 ;
      RECT 26.35 -86 26.45 -85.19 ;
      RECT 25.15 -86 25.25 -85.19 ;
      RECT 23.95 -86 24.05 -85.19 ;
      RECT 22.75 -86 22.85 -85.19 ;
      RECT 21.55 -86 21.65 -85.19 ;
      RECT 20.35 -86 20.45 -85.19 ;
      RECT 19.15 -86 19.25 -85.19 ;
      RECT 17.95 -86 18.05 -85.19 ;
      RECT 16.75 -86 16.85 -85.19 ;
      RECT 15.55 -86 15.65 -85.19 ;
      RECT 14.35 -86 14.45 -85.19 ;
      RECT 13.15 -86 13.25 -85.19 ;
      RECT 11.95 -86 12.05 -85.19 ;
      RECT 10.75 -86 10.85 -85.19 ;
      RECT 9.55 -86 9.65 -85.19 ;
      RECT 8.35 -86 8.45 -85.19 ;
      RECT 7.15 -86 7.25 -85.19 ;
      RECT 5.95 -86 6.05 -85.19 ;
      RECT 4.75 -86 4.85 -85.19 ;
      RECT 3.55 -86 3.65 -85.19 ;
      RECT 2.35 -86 2.45 -85.19 ;
      RECT 1.15 -86 1.25 -85.19 ;
      RECT -0.05 -86 0.05 -85.19 ;
      RECT -0.105 -85.655 156.465 -85.535 ;
      RECT 153.55 -82.77 153.65 -81.96 ;
      RECT 152.35 -82.77 152.45 -81.96 ;
      RECT 151.15 -82.77 151.25 -81.96 ;
      RECT 149.95 -82.77 150.05 -81.96 ;
      RECT 148.75 -82.77 148.85 -81.96 ;
      RECT 147.55 -82.77 147.65 -81.96 ;
      RECT 146.35 -82.77 146.45 -81.96 ;
      RECT 145.15 -82.77 145.25 -81.96 ;
      RECT 143.95 -82.77 144.05 -81.96 ;
      RECT 142.75 -82.77 142.85 -81.96 ;
      RECT 141.55 -82.77 141.65 -81.96 ;
      RECT 140.35 -82.77 140.45 -81.96 ;
      RECT 139.15 -82.77 139.25 -81.96 ;
      RECT 137.95 -82.77 138.05 -81.96 ;
      RECT 136.75 -82.77 136.85 -81.96 ;
      RECT 135.55 -82.77 135.65 -81.96 ;
      RECT 134.35 -82.77 134.45 -81.96 ;
      RECT 133.15 -82.77 133.25 -81.96 ;
      RECT 131.95 -82.77 132.05 -81.96 ;
      RECT 130.75 -82.77 130.85 -81.96 ;
      RECT 129.55 -82.77 129.65 -81.96 ;
      RECT 128.35 -82.77 128.45 -81.96 ;
      RECT 127.15 -82.77 127.25 -81.96 ;
      RECT 125.95 -82.77 126.05 -81.96 ;
      RECT 124.75 -82.77 124.85 -81.96 ;
      RECT 123.55 -82.77 123.65 -81.96 ;
      RECT 122.35 -82.77 122.45 -81.96 ;
      RECT 121.15 -82.77 121.25 -81.96 ;
      RECT 119.95 -82.77 120.05 -81.96 ;
      RECT 118.75 -82.77 118.85 -81.96 ;
      RECT 117.55 -82.77 117.65 -81.96 ;
      RECT 116.35 -82.77 116.45 -81.96 ;
      RECT 115.15 -82.77 115.25 -81.96 ;
      RECT 113.95 -82.77 114.05 -81.96 ;
      RECT 112.75 -82.77 112.85 -81.96 ;
      RECT 111.55 -82.77 111.65 -81.96 ;
      RECT 110.35 -82.77 110.45 -81.96 ;
      RECT 109.15 -82.77 109.25 -81.96 ;
      RECT 107.95 -82.77 108.05 -81.96 ;
      RECT 106.75 -82.77 106.85 -81.96 ;
      RECT 105.55 -82.77 105.65 -81.96 ;
      RECT 104.35 -82.77 104.45 -81.96 ;
      RECT 103.15 -82.77 103.25 -81.96 ;
      RECT 101.95 -82.77 102.05 -81.96 ;
      RECT 100.75 -82.77 100.85 -81.96 ;
      RECT 99.55 -82.77 99.65 -81.96 ;
      RECT 98.35 -82.77 98.45 -81.96 ;
      RECT 97.15 -82.77 97.25 -81.96 ;
      RECT 95.95 -82.77 96.05 -81.96 ;
      RECT 94.75 -82.77 94.85 -81.96 ;
      RECT 93.55 -82.77 93.65 -81.96 ;
      RECT 92.35 -82.77 92.45 -81.96 ;
      RECT 91.15 -82.77 91.25 -81.96 ;
      RECT 89.95 -82.77 90.05 -81.96 ;
      RECT 88.75 -82.77 88.85 -81.96 ;
      RECT 87.55 -82.77 87.65 -81.96 ;
      RECT 86.35 -82.77 86.45 -81.96 ;
      RECT 85.15 -82.77 85.25 -81.96 ;
      RECT 83.95 -82.77 84.05 -81.96 ;
      RECT 82.75 -82.77 82.85 -81.96 ;
      RECT 81.55 -82.77 81.65 -81.96 ;
      RECT 80.35 -82.77 80.45 -81.96 ;
      RECT 79.15 -82.77 79.25 -81.96 ;
      RECT 77.95 -82.77 78.05 -81.96 ;
      RECT 76.75 -82.77 76.85 -81.96 ;
      RECT 75.55 -82.77 75.65 -81.96 ;
      RECT 74.35 -82.77 74.45 -81.96 ;
      RECT 73.15 -82.77 73.25 -81.96 ;
      RECT 71.95 -82.77 72.05 -81.96 ;
      RECT 70.75 -82.77 70.85 -81.96 ;
      RECT 69.55 -82.77 69.65 -81.96 ;
      RECT 68.35 -82.77 68.45 -81.96 ;
      RECT 67.15 -82.77 67.25 -81.96 ;
      RECT 65.95 -82.77 66.05 -81.96 ;
      RECT 64.75 -82.77 64.85 -81.96 ;
      RECT 63.55 -82.77 63.65 -81.96 ;
      RECT 62.35 -82.77 62.45 -81.96 ;
      RECT 61.15 -82.77 61.25 -81.96 ;
      RECT 59.95 -82.77 60.05 -81.96 ;
      RECT 58.75 -82.77 58.85 -81.96 ;
      RECT 57.55 -82.77 57.65 -81.96 ;
      RECT 56.35 -82.77 56.45 -81.96 ;
      RECT 55.15 -82.77 55.25 -81.96 ;
      RECT 53.95 -82.77 54.05 -81.96 ;
      RECT 52.75 -82.77 52.85 -81.96 ;
      RECT 51.55 -82.77 51.65 -81.96 ;
      RECT 50.35 -82.77 50.45 -81.96 ;
      RECT 49.15 -82.77 49.25 -81.96 ;
      RECT 47.95 -82.77 48.05 -81.96 ;
      RECT 46.75 -82.77 46.85 -81.96 ;
      RECT 45.55 -82.77 45.65 -81.96 ;
      RECT 44.35 -82.77 44.45 -81.96 ;
      RECT 43.15 -82.77 43.25 -81.96 ;
      RECT 41.95 -82.77 42.05 -81.96 ;
      RECT 40.75 -82.77 40.85 -81.96 ;
      RECT 39.55 -82.77 39.65 -81.96 ;
      RECT 38.35 -82.77 38.45 -81.96 ;
      RECT 37.15 -82.77 37.25 -81.96 ;
      RECT 35.95 -82.77 36.05 -81.96 ;
      RECT 34.75 -82.77 34.85 -81.96 ;
      RECT 33.55 -82.77 33.65 -81.96 ;
      RECT 32.35 -82.77 32.45 -81.96 ;
      RECT 31.15 -82.77 31.25 -81.96 ;
      RECT 29.95 -82.77 30.05 -81.96 ;
      RECT 28.75 -82.77 28.85 -81.96 ;
      RECT 27.55 -82.77 27.65 -81.96 ;
      RECT 26.35 -82.77 26.45 -81.96 ;
      RECT 25.15 -82.77 25.25 -81.96 ;
      RECT 23.95 -82.77 24.05 -81.96 ;
      RECT 22.75 -82.77 22.85 -81.96 ;
      RECT 21.55 -82.77 21.65 -81.96 ;
      RECT 20.35 -82.77 20.45 -81.96 ;
      RECT 19.15 -82.77 19.25 -81.96 ;
      RECT 17.95 -82.77 18.05 -81.96 ;
      RECT 16.75 -82.77 16.85 -81.96 ;
      RECT 15.55 -82.77 15.65 -81.96 ;
      RECT 14.35 -82.77 14.45 -81.96 ;
      RECT 13.15 -82.77 13.25 -81.96 ;
      RECT 11.95 -82.77 12.05 -81.96 ;
      RECT 10.75 -82.77 10.85 -81.96 ;
      RECT 9.55 -82.77 9.65 -81.96 ;
      RECT 8.35 -82.77 8.45 -81.96 ;
      RECT 7.15 -82.77 7.25 -81.96 ;
      RECT 5.95 -82.77 6.05 -81.96 ;
      RECT 4.75 -82.77 4.85 -81.96 ;
      RECT 3.55 -82.77 3.65 -81.96 ;
      RECT 2.35 -82.77 2.45 -81.96 ;
      RECT 1.15 -82.77 1.25 -81.96 ;
      RECT -0.05 -82.77 0.05 -81.96 ;
      RECT -0.105 -82.425 156.465 -82.305 ;
      RECT 153.55 -79.54 153.65 -78.73 ;
      RECT 152.35 -79.54 152.45 -78.73 ;
      RECT 151.15 -79.54 151.25 -78.73 ;
      RECT 149.95 -79.54 150.05 -78.73 ;
      RECT 148.75 -79.54 148.85 -78.73 ;
      RECT 147.55 -79.54 147.65 -78.73 ;
      RECT 146.35 -79.54 146.45 -78.73 ;
      RECT 145.15 -79.54 145.25 -78.73 ;
      RECT 143.95 -79.54 144.05 -78.73 ;
      RECT 142.75 -79.54 142.85 -78.73 ;
      RECT 141.55 -79.54 141.65 -78.73 ;
      RECT 140.35 -79.54 140.45 -78.73 ;
      RECT 139.15 -79.54 139.25 -78.73 ;
      RECT 137.95 -79.54 138.05 -78.73 ;
      RECT 136.75 -79.54 136.85 -78.73 ;
      RECT 135.55 -79.54 135.65 -78.73 ;
      RECT 134.35 -79.54 134.45 -78.73 ;
      RECT 133.15 -79.54 133.25 -78.73 ;
      RECT 131.95 -79.54 132.05 -78.73 ;
      RECT 130.75 -79.54 130.85 -78.73 ;
      RECT 129.55 -79.54 129.65 -78.73 ;
      RECT 128.35 -79.54 128.45 -78.73 ;
      RECT 127.15 -79.54 127.25 -78.73 ;
      RECT 125.95 -79.54 126.05 -78.73 ;
      RECT 124.75 -79.54 124.85 -78.73 ;
      RECT 123.55 -79.54 123.65 -78.73 ;
      RECT 122.35 -79.54 122.45 -78.73 ;
      RECT 121.15 -79.54 121.25 -78.73 ;
      RECT 119.95 -79.54 120.05 -78.73 ;
      RECT 118.75 -79.54 118.85 -78.73 ;
      RECT 117.55 -79.54 117.65 -78.73 ;
      RECT 116.35 -79.54 116.45 -78.73 ;
      RECT 115.15 -79.54 115.25 -78.73 ;
      RECT 113.95 -79.54 114.05 -78.73 ;
      RECT 112.75 -79.54 112.85 -78.73 ;
      RECT 111.55 -79.54 111.65 -78.73 ;
      RECT 110.35 -79.54 110.45 -78.73 ;
      RECT 109.15 -79.54 109.25 -78.73 ;
      RECT 107.95 -79.54 108.05 -78.73 ;
      RECT 106.75 -79.54 106.85 -78.73 ;
      RECT 105.55 -79.54 105.65 -78.73 ;
      RECT 104.35 -79.54 104.45 -78.73 ;
      RECT 103.15 -79.54 103.25 -78.73 ;
      RECT 101.95 -79.54 102.05 -78.73 ;
      RECT 100.75 -79.54 100.85 -78.73 ;
      RECT 99.55 -79.54 99.65 -78.73 ;
      RECT 98.35 -79.54 98.45 -78.73 ;
      RECT 97.15 -79.54 97.25 -78.73 ;
      RECT 95.95 -79.54 96.05 -78.73 ;
      RECT 94.75 -79.54 94.85 -78.73 ;
      RECT 93.55 -79.54 93.65 -78.73 ;
      RECT 92.35 -79.54 92.45 -78.73 ;
      RECT 91.15 -79.54 91.25 -78.73 ;
      RECT 89.95 -79.54 90.05 -78.73 ;
      RECT 88.75 -79.54 88.85 -78.73 ;
      RECT 87.55 -79.54 87.65 -78.73 ;
      RECT 86.35 -79.54 86.45 -78.73 ;
      RECT 85.15 -79.54 85.25 -78.73 ;
      RECT 83.95 -79.54 84.05 -78.73 ;
      RECT 82.75 -79.54 82.85 -78.73 ;
      RECT 81.55 -79.54 81.65 -78.73 ;
      RECT 80.35 -79.54 80.45 -78.73 ;
      RECT 79.15 -79.54 79.25 -78.73 ;
      RECT 77.95 -79.54 78.05 -78.73 ;
      RECT 76.75 -79.54 76.85 -78.73 ;
      RECT 75.55 -79.54 75.65 -78.73 ;
      RECT 74.35 -79.54 74.45 -78.73 ;
      RECT 73.15 -79.54 73.25 -78.73 ;
      RECT 71.95 -79.54 72.05 -78.73 ;
      RECT 70.75 -79.54 70.85 -78.73 ;
      RECT 69.55 -79.54 69.65 -78.73 ;
      RECT 68.35 -79.54 68.45 -78.73 ;
      RECT 67.15 -79.54 67.25 -78.73 ;
      RECT 65.95 -79.54 66.05 -78.73 ;
      RECT 64.75 -79.54 64.85 -78.73 ;
      RECT 63.55 -79.54 63.65 -78.73 ;
      RECT 62.35 -79.54 62.45 -78.73 ;
      RECT 61.15 -79.54 61.25 -78.73 ;
      RECT 59.95 -79.54 60.05 -78.73 ;
      RECT 58.75 -79.54 58.85 -78.73 ;
      RECT 57.55 -79.54 57.65 -78.73 ;
      RECT 56.35 -79.54 56.45 -78.73 ;
      RECT 55.15 -79.54 55.25 -78.73 ;
      RECT 53.95 -79.54 54.05 -78.73 ;
      RECT 52.75 -79.54 52.85 -78.73 ;
      RECT 51.55 -79.54 51.65 -78.73 ;
      RECT 50.35 -79.54 50.45 -78.73 ;
      RECT 49.15 -79.54 49.25 -78.73 ;
      RECT 47.95 -79.54 48.05 -78.73 ;
      RECT 46.75 -79.54 46.85 -78.73 ;
      RECT 45.55 -79.54 45.65 -78.73 ;
      RECT 44.35 -79.54 44.45 -78.73 ;
      RECT 43.15 -79.54 43.25 -78.73 ;
      RECT 41.95 -79.54 42.05 -78.73 ;
      RECT 40.75 -79.54 40.85 -78.73 ;
      RECT 39.55 -79.54 39.65 -78.73 ;
      RECT 38.35 -79.54 38.45 -78.73 ;
      RECT 37.15 -79.54 37.25 -78.73 ;
      RECT 35.95 -79.54 36.05 -78.73 ;
      RECT 34.75 -79.54 34.85 -78.73 ;
      RECT 33.55 -79.54 33.65 -78.73 ;
      RECT 32.35 -79.54 32.45 -78.73 ;
      RECT 31.15 -79.54 31.25 -78.73 ;
      RECT 29.95 -79.54 30.05 -78.73 ;
      RECT 28.75 -79.54 28.85 -78.73 ;
      RECT 27.55 -79.54 27.65 -78.73 ;
      RECT 26.35 -79.54 26.45 -78.73 ;
      RECT 25.15 -79.54 25.25 -78.73 ;
      RECT 23.95 -79.54 24.05 -78.73 ;
      RECT 22.75 -79.54 22.85 -78.73 ;
      RECT 21.55 -79.54 21.65 -78.73 ;
      RECT 20.35 -79.54 20.45 -78.73 ;
      RECT 19.15 -79.54 19.25 -78.73 ;
      RECT 17.95 -79.54 18.05 -78.73 ;
      RECT 16.75 -79.54 16.85 -78.73 ;
      RECT 15.55 -79.54 15.65 -78.73 ;
      RECT 14.35 -79.54 14.45 -78.73 ;
      RECT 13.15 -79.54 13.25 -78.73 ;
      RECT 11.95 -79.54 12.05 -78.73 ;
      RECT 10.75 -79.54 10.85 -78.73 ;
      RECT 9.55 -79.54 9.65 -78.73 ;
      RECT 8.35 -79.54 8.45 -78.73 ;
      RECT 7.15 -79.54 7.25 -78.73 ;
      RECT 5.95 -79.54 6.05 -78.73 ;
      RECT 4.75 -79.54 4.85 -78.73 ;
      RECT 3.55 -79.54 3.65 -78.73 ;
      RECT 2.35 -79.54 2.45 -78.73 ;
      RECT 1.15 -79.54 1.25 -78.73 ;
      RECT -0.05 -79.54 0.05 -78.73 ;
      RECT -0.105 -79.195 156.465 -79.075 ;
      RECT 153.55 -76.31 153.65 -75.5 ;
      RECT 152.35 -76.31 152.45 -75.5 ;
      RECT 151.15 -76.31 151.25 -75.5 ;
      RECT 149.95 -76.31 150.05 -75.5 ;
      RECT 148.75 -76.31 148.85 -75.5 ;
      RECT 147.55 -76.31 147.65 -75.5 ;
      RECT 146.35 -76.31 146.45 -75.5 ;
      RECT 145.15 -76.31 145.25 -75.5 ;
      RECT 143.95 -76.31 144.05 -75.5 ;
      RECT 142.75 -76.31 142.85 -75.5 ;
      RECT 141.55 -76.31 141.65 -75.5 ;
      RECT 140.35 -76.31 140.45 -75.5 ;
      RECT 139.15 -76.31 139.25 -75.5 ;
      RECT 137.95 -76.31 138.05 -75.5 ;
      RECT 136.75 -76.31 136.85 -75.5 ;
      RECT 135.55 -76.31 135.65 -75.5 ;
      RECT 134.35 -76.31 134.45 -75.5 ;
      RECT 133.15 -76.31 133.25 -75.5 ;
      RECT 131.95 -76.31 132.05 -75.5 ;
      RECT 130.75 -76.31 130.85 -75.5 ;
      RECT 129.55 -76.31 129.65 -75.5 ;
      RECT 128.35 -76.31 128.45 -75.5 ;
      RECT 127.15 -76.31 127.25 -75.5 ;
      RECT 125.95 -76.31 126.05 -75.5 ;
      RECT 124.75 -76.31 124.85 -75.5 ;
      RECT 123.55 -76.31 123.65 -75.5 ;
      RECT 122.35 -76.31 122.45 -75.5 ;
      RECT 121.15 -76.31 121.25 -75.5 ;
      RECT 119.95 -76.31 120.05 -75.5 ;
      RECT 118.75 -76.31 118.85 -75.5 ;
      RECT 117.55 -76.31 117.65 -75.5 ;
      RECT 116.35 -76.31 116.45 -75.5 ;
      RECT 115.15 -76.31 115.25 -75.5 ;
      RECT 113.95 -76.31 114.05 -75.5 ;
      RECT 112.75 -76.31 112.85 -75.5 ;
      RECT 111.55 -76.31 111.65 -75.5 ;
      RECT 110.35 -76.31 110.45 -75.5 ;
      RECT 109.15 -76.31 109.25 -75.5 ;
      RECT 107.95 -76.31 108.05 -75.5 ;
      RECT 106.75 -76.31 106.85 -75.5 ;
      RECT 105.55 -76.31 105.65 -75.5 ;
      RECT 104.35 -76.31 104.45 -75.5 ;
      RECT 103.15 -76.31 103.25 -75.5 ;
      RECT 101.95 -76.31 102.05 -75.5 ;
      RECT 100.75 -76.31 100.85 -75.5 ;
      RECT 99.55 -76.31 99.65 -75.5 ;
      RECT 98.35 -76.31 98.45 -75.5 ;
      RECT 97.15 -76.31 97.25 -75.5 ;
      RECT 95.95 -76.31 96.05 -75.5 ;
      RECT 94.75 -76.31 94.85 -75.5 ;
      RECT 93.55 -76.31 93.65 -75.5 ;
      RECT 92.35 -76.31 92.45 -75.5 ;
      RECT 91.15 -76.31 91.25 -75.5 ;
      RECT 89.95 -76.31 90.05 -75.5 ;
      RECT 88.75 -76.31 88.85 -75.5 ;
      RECT 87.55 -76.31 87.65 -75.5 ;
      RECT 86.35 -76.31 86.45 -75.5 ;
      RECT 85.15 -76.31 85.25 -75.5 ;
      RECT 83.95 -76.31 84.05 -75.5 ;
      RECT 82.75 -76.31 82.85 -75.5 ;
      RECT 81.55 -76.31 81.65 -75.5 ;
      RECT 80.35 -76.31 80.45 -75.5 ;
      RECT 79.15 -76.31 79.25 -75.5 ;
      RECT 77.95 -76.31 78.05 -75.5 ;
      RECT 76.75 -76.31 76.85 -75.5 ;
      RECT 75.55 -76.31 75.65 -75.5 ;
      RECT 74.35 -76.31 74.45 -75.5 ;
      RECT 73.15 -76.31 73.25 -75.5 ;
      RECT 71.95 -76.31 72.05 -75.5 ;
      RECT 70.75 -76.31 70.85 -75.5 ;
      RECT 69.55 -76.31 69.65 -75.5 ;
      RECT 68.35 -76.31 68.45 -75.5 ;
      RECT 67.15 -76.31 67.25 -75.5 ;
      RECT 65.95 -76.31 66.05 -75.5 ;
      RECT 64.75 -76.31 64.85 -75.5 ;
      RECT 63.55 -76.31 63.65 -75.5 ;
      RECT 62.35 -76.31 62.45 -75.5 ;
      RECT 61.15 -76.31 61.25 -75.5 ;
      RECT 59.95 -76.31 60.05 -75.5 ;
      RECT 58.75 -76.31 58.85 -75.5 ;
      RECT 57.55 -76.31 57.65 -75.5 ;
      RECT 56.35 -76.31 56.45 -75.5 ;
      RECT 55.15 -76.31 55.25 -75.5 ;
      RECT 53.95 -76.31 54.05 -75.5 ;
      RECT 52.75 -76.31 52.85 -75.5 ;
      RECT 51.55 -76.31 51.65 -75.5 ;
      RECT 50.35 -76.31 50.45 -75.5 ;
      RECT 49.15 -76.31 49.25 -75.5 ;
      RECT 47.95 -76.31 48.05 -75.5 ;
      RECT 46.75 -76.31 46.85 -75.5 ;
      RECT 45.55 -76.31 45.65 -75.5 ;
      RECT 44.35 -76.31 44.45 -75.5 ;
      RECT 43.15 -76.31 43.25 -75.5 ;
      RECT 41.95 -76.31 42.05 -75.5 ;
      RECT 40.75 -76.31 40.85 -75.5 ;
      RECT 39.55 -76.31 39.65 -75.5 ;
      RECT 38.35 -76.31 38.45 -75.5 ;
      RECT 37.15 -76.31 37.25 -75.5 ;
      RECT 35.95 -76.31 36.05 -75.5 ;
      RECT 34.75 -76.31 34.85 -75.5 ;
      RECT 33.55 -76.31 33.65 -75.5 ;
      RECT 32.35 -76.31 32.45 -75.5 ;
      RECT 31.15 -76.31 31.25 -75.5 ;
      RECT 29.95 -76.31 30.05 -75.5 ;
      RECT 28.75 -76.31 28.85 -75.5 ;
      RECT 27.55 -76.31 27.65 -75.5 ;
      RECT 26.35 -76.31 26.45 -75.5 ;
      RECT 25.15 -76.31 25.25 -75.5 ;
      RECT 23.95 -76.31 24.05 -75.5 ;
      RECT 22.75 -76.31 22.85 -75.5 ;
      RECT 21.55 -76.31 21.65 -75.5 ;
      RECT 20.35 -76.31 20.45 -75.5 ;
      RECT 19.15 -76.31 19.25 -75.5 ;
      RECT 17.95 -76.31 18.05 -75.5 ;
      RECT 16.75 -76.31 16.85 -75.5 ;
      RECT 15.55 -76.31 15.65 -75.5 ;
      RECT 14.35 -76.31 14.45 -75.5 ;
      RECT 13.15 -76.31 13.25 -75.5 ;
      RECT 11.95 -76.31 12.05 -75.5 ;
      RECT 10.75 -76.31 10.85 -75.5 ;
      RECT 9.55 -76.31 9.65 -75.5 ;
      RECT 8.35 -76.31 8.45 -75.5 ;
      RECT 7.15 -76.31 7.25 -75.5 ;
      RECT 5.95 -76.31 6.05 -75.5 ;
      RECT 4.75 -76.31 4.85 -75.5 ;
      RECT 3.55 -76.31 3.65 -75.5 ;
      RECT 2.35 -76.31 2.45 -75.5 ;
      RECT 1.15 -76.31 1.25 -75.5 ;
      RECT -0.05 -76.31 0.05 -75.5 ;
      RECT -0.105 -75.965 156.465 -75.845 ;
      RECT 153.55 -73.08 153.65 -72.27 ;
      RECT 152.35 -73.08 152.45 -72.27 ;
      RECT 151.15 -73.08 151.25 -72.27 ;
      RECT 149.95 -73.08 150.05 -72.27 ;
      RECT 148.75 -73.08 148.85 -72.27 ;
      RECT 147.55 -73.08 147.65 -72.27 ;
      RECT 146.35 -73.08 146.45 -72.27 ;
      RECT 145.15 -73.08 145.25 -72.27 ;
      RECT 143.95 -73.08 144.05 -72.27 ;
      RECT 142.75 -73.08 142.85 -72.27 ;
      RECT 141.55 -73.08 141.65 -72.27 ;
      RECT 140.35 -73.08 140.45 -72.27 ;
      RECT 139.15 -73.08 139.25 -72.27 ;
      RECT 137.95 -73.08 138.05 -72.27 ;
      RECT 136.75 -73.08 136.85 -72.27 ;
      RECT 135.55 -73.08 135.65 -72.27 ;
      RECT 134.35 -73.08 134.45 -72.27 ;
      RECT 133.15 -73.08 133.25 -72.27 ;
      RECT 131.95 -73.08 132.05 -72.27 ;
      RECT 130.75 -73.08 130.85 -72.27 ;
      RECT 129.55 -73.08 129.65 -72.27 ;
      RECT 128.35 -73.08 128.45 -72.27 ;
      RECT 127.15 -73.08 127.25 -72.27 ;
      RECT 125.95 -73.08 126.05 -72.27 ;
      RECT 124.75 -73.08 124.85 -72.27 ;
      RECT 123.55 -73.08 123.65 -72.27 ;
      RECT 122.35 -73.08 122.45 -72.27 ;
      RECT 121.15 -73.08 121.25 -72.27 ;
      RECT 119.95 -73.08 120.05 -72.27 ;
      RECT 118.75 -73.08 118.85 -72.27 ;
      RECT 117.55 -73.08 117.65 -72.27 ;
      RECT 116.35 -73.08 116.45 -72.27 ;
      RECT 115.15 -73.08 115.25 -72.27 ;
      RECT 113.95 -73.08 114.05 -72.27 ;
      RECT 112.75 -73.08 112.85 -72.27 ;
      RECT 111.55 -73.08 111.65 -72.27 ;
      RECT 110.35 -73.08 110.45 -72.27 ;
      RECT 109.15 -73.08 109.25 -72.27 ;
      RECT 107.95 -73.08 108.05 -72.27 ;
      RECT 106.75 -73.08 106.85 -72.27 ;
      RECT 105.55 -73.08 105.65 -72.27 ;
      RECT 104.35 -73.08 104.45 -72.27 ;
      RECT 103.15 -73.08 103.25 -72.27 ;
      RECT 101.95 -73.08 102.05 -72.27 ;
      RECT 100.75 -73.08 100.85 -72.27 ;
      RECT 99.55 -73.08 99.65 -72.27 ;
      RECT 98.35 -73.08 98.45 -72.27 ;
      RECT 97.15 -73.08 97.25 -72.27 ;
      RECT 95.95 -73.08 96.05 -72.27 ;
      RECT 94.75 -73.08 94.85 -72.27 ;
      RECT 93.55 -73.08 93.65 -72.27 ;
      RECT 92.35 -73.08 92.45 -72.27 ;
      RECT 91.15 -73.08 91.25 -72.27 ;
      RECT 89.95 -73.08 90.05 -72.27 ;
      RECT 88.75 -73.08 88.85 -72.27 ;
      RECT 87.55 -73.08 87.65 -72.27 ;
      RECT 86.35 -73.08 86.45 -72.27 ;
      RECT 85.15 -73.08 85.25 -72.27 ;
      RECT 83.95 -73.08 84.05 -72.27 ;
      RECT 82.75 -73.08 82.85 -72.27 ;
      RECT 81.55 -73.08 81.65 -72.27 ;
      RECT 80.35 -73.08 80.45 -72.27 ;
      RECT 79.15 -73.08 79.25 -72.27 ;
      RECT 77.95 -73.08 78.05 -72.27 ;
      RECT 76.75 -73.08 76.85 -72.27 ;
      RECT 75.55 -73.08 75.65 -72.27 ;
      RECT 74.35 -73.08 74.45 -72.27 ;
      RECT 73.15 -73.08 73.25 -72.27 ;
      RECT 71.95 -73.08 72.05 -72.27 ;
      RECT 70.75 -73.08 70.85 -72.27 ;
      RECT 69.55 -73.08 69.65 -72.27 ;
      RECT 68.35 -73.08 68.45 -72.27 ;
      RECT 67.15 -73.08 67.25 -72.27 ;
      RECT 65.95 -73.08 66.05 -72.27 ;
      RECT 64.75 -73.08 64.85 -72.27 ;
      RECT 63.55 -73.08 63.65 -72.27 ;
      RECT 62.35 -73.08 62.45 -72.27 ;
      RECT 61.15 -73.08 61.25 -72.27 ;
      RECT 59.95 -73.08 60.05 -72.27 ;
      RECT 58.75 -73.08 58.85 -72.27 ;
      RECT 57.55 -73.08 57.65 -72.27 ;
      RECT 56.35 -73.08 56.45 -72.27 ;
      RECT 55.15 -73.08 55.25 -72.27 ;
      RECT 53.95 -73.08 54.05 -72.27 ;
      RECT 52.75 -73.08 52.85 -72.27 ;
      RECT 51.55 -73.08 51.65 -72.27 ;
      RECT 50.35 -73.08 50.45 -72.27 ;
      RECT 49.15 -73.08 49.25 -72.27 ;
      RECT 47.95 -73.08 48.05 -72.27 ;
      RECT 46.75 -73.08 46.85 -72.27 ;
      RECT 45.55 -73.08 45.65 -72.27 ;
      RECT 44.35 -73.08 44.45 -72.27 ;
      RECT 43.15 -73.08 43.25 -72.27 ;
      RECT 41.95 -73.08 42.05 -72.27 ;
      RECT 40.75 -73.08 40.85 -72.27 ;
      RECT 39.55 -73.08 39.65 -72.27 ;
      RECT 38.35 -73.08 38.45 -72.27 ;
      RECT 37.15 -73.08 37.25 -72.27 ;
      RECT 35.95 -73.08 36.05 -72.27 ;
      RECT 34.75 -73.08 34.85 -72.27 ;
      RECT 33.55 -73.08 33.65 -72.27 ;
      RECT 32.35 -73.08 32.45 -72.27 ;
      RECT 31.15 -73.08 31.25 -72.27 ;
      RECT 29.95 -73.08 30.05 -72.27 ;
      RECT 28.75 -73.08 28.85 -72.27 ;
      RECT 27.55 -73.08 27.65 -72.27 ;
      RECT 26.35 -73.08 26.45 -72.27 ;
      RECT 25.15 -73.08 25.25 -72.27 ;
      RECT 23.95 -73.08 24.05 -72.27 ;
      RECT 22.75 -73.08 22.85 -72.27 ;
      RECT 21.55 -73.08 21.65 -72.27 ;
      RECT 20.35 -73.08 20.45 -72.27 ;
      RECT 19.15 -73.08 19.25 -72.27 ;
      RECT 17.95 -73.08 18.05 -72.27 ;
      RECT 16.75 -73.08 16.85 -72.27 ;
      RECT 15.55 -73.08 15.65 -72.27 ;
      RECT 14.35 -73.08 14.45 -72.27 ;
      RECT 13.15 -73.08 13.25 -72.27 ;
      RECT 11.95 -73.08 12.05 -72.27 ;
      RECT 10.75 -73.08 10.85 -72.27 ;
      RECT 9.55 -73.08 9.65 -72.27 ;
      RECT 8.35 -73.08 8.45 -72.27 ;
      RECT 7.15 -73.08 7.25 -72.27 ;
      RECT 5.95 -73.08 6.05 -72.27 ;
      RECT 4.75 -73.08 4.85 -72.27 ;
      RECT 3.55 -73.08 3.65 -72.27 ;
      RECT 2.35 -73.08 2.45 -72.27 ;
      RECT 1.15 -73.08 1.25 -72.27 ;
      RECT -0.05 -73.08 0.05 -72.27 ;
      RECT -0.105 -72.735 156.465 -72.615 ;
      RECT 153.55 -69.85 153.65 -69.04 ;
      RECT 152.35 -69.85 152.45 -69.04 ;
      RECT 151.15 -69.85 151.25 -69.04 ;
      RECT 149.95 -69.85 150.05 -69.04 ;
      RECT 148.75 -69.85 148.85 -69.04 ;
      RECT 147.55 -69.85 147.65 -69.04 ;
      RECT 146.35 -69.85 146.45 -69.04 ;
      RECT 145.15 -69.85 145.25 -69.04 ;
      RECT 143.95 -69.85 144.05 -69.04 ;
      RECT 142.75 -69.85 142.85 -69.04 ;
      RECT 141.55 -69.85 141.65 -69.04 ;
      RECT 140.35 -69.85 140.45 -69.04 ;
      RECT 139.15 -69.85 139.25 -69.04 ;
      RECT 137.95 -69.85 138.05 -69.04 ;
      RECT 136.75 -69.85 136.85 -69.04 ;
      RECT 135.55 -69.85 135.65 -69.04 ;
      RECT 134.35 -69.85 134.45 -69.04 ;
      RECT 133.15 -69.85 133.25 -69.04 ;
      RECT 131.95 -69.85 132.05 -69.04 ;
      RECT 130.75 -69.85 130.85 -69.04 ;
      RECT 129.55 -69.85 129.65 -69.04 ;
      RECT 128.35 -69.85 128.45 -69.04 ;
      RECT 127.15 -69.85 127.25 -69.04 ;
      RECT 125.95 -69.85 126.05 -69.04 ;
      RECT 124.75 -69.85 124.85 -69.04 ;
      RECT 123.55 -69.85 123.65 -69.04 ;
      RECT 122.35 -69.85 122.45 -69.04 ;
      RECT 121.15 -69.85 121.25 -69.04 ;
      RECT 119.95 -69.85 120.05 -69.04 ;
      RECT 118.75 -69.85 118.85 -69.04 ;
      RECT 117.55 -69.85 117.65 -69.04 ;
      RECT 116.35 -69.85 116.45 -69.04 ;
      RECT 115.15 -69.85 115.25 -69.04 ;
      RECT 113.95 -69.85 114.05 -69.04 ;
      RECT 112.75 -69.85 112.85 -69.04 ;
      RECT 111.55 -69.85 111.65 -69.04 ;
      RECT 110.35 -69.85 110.45 -69.04 ;
      RECT 109.15 -69.85 109.25 -69.04 ;
      RECT 107.95 -69.85 108.05 -69.04 ;
      RECT 106.75 -69.85 106.85 -69.04 ;
      RECT 105.55 -69.85 105.65 -69.04 ;
      RECT 104.35 -69.85 104.45 -69.04 ;
      RECT 103.15 -69.85 103.25 -69.04 ;
      RECT 101.95 -69.85 102.05 -69.04 ;
      RECT 100.75 -69.85 100.85 -69.04 ;
      RECT 99.55 -69.85 99.65 -69.04 ;
      RECT 98.35 -69.85 98.45 -69.04 ;
      RECT 97.15 -69.85 97.25 -69.04 ;
      RECT 95.95 -69.85 96.05 -69.04 ;
      RECT 94.75 -69.85 94.85 -69.04 ;
      RECT 93.55 -69.85 93.65 -69.04 ;
      RECT 92.35 -69.85 92.45 -69.04 ;
      RECT 91.15 -69.85 91.25 -69.04 ;
      RECT 89.95 -69.85 90.05 -69.04 ;
      RECT 88.75 -69.85 88.85 -69.04 ;
      RECT 87.55 -69.85 87.65 -69.04 ;
      RECT 86.35 -69.85 86.45 -69.04 ;
      RECT 85.15 -69.85 85.25 -69.04 ;
      RECT 83.95 -69.85 84.05 -69.04 ;
      RECT 82.75 -69.85 82.85 -69.04 ;
      RECT 81.55 -69.85 81.65 -69.04 ;
      RECT 80.35 -69.85 80.45 -69.04 ;
      RECT 79.15 -69.85 79.25 -69.04 ;
      RECT 77.95 -69.85 78.05 -69.04 ;
      RECT 76.75 -69.85 76.85 -69.04 ;
      RECT 75.55 -69.85 75.65 -69.04 ;
      RECT 74.35 -69.85 74.45 -69.04 ;
      RECT 73.15 -69.85 73.25 -69.04 ;
      RECT 71.95 -69.85 72.05 -69.04 ;
      RECT 70.75 -69.85 70.85 -69.04 ;
      RECT 69.55 -69.85 69.65 -69.04 ;
      RECT 68.35 -69.85 68.45 -69.04 ;
      RECT 67.15 -69.85 67.25 -69.04 ;
      RECT 65.95 -69.85 66.05 -69.04 ;
      RECT 64.75 -69.85 64.85 -69.04 ;
      RECT 63.55 -69.85 63.65 -69.04 ;
      RECT 62.35 -69.85 62.45 -69.04 ;
      RECT 61.15 -69.85 61.25 -69.04 ;
      RECT 59.95 -69.85 60.05 -69.04 ;
      RECT 58.75 -69.85 58.85 -69.04 ;
      RECT 57.55 -69.85 57.65 -69.04 ;
      RECT 56.35 -69.85 56.45 -69.04 ;
      RECT 55.15 -69.85 55.25 -69.04 ;
      RECT 53.95 -69.85 54.05 -69.04 ;
      RECT 52.75 -69.85 52.85 -69.04 ;
      RECT 51.55 -69.85 51.65 -69.04 ;
      RECT 50.35 -69.85 50.45 -69.04 ;
      RECT 49.15 -69.85 49.25 -69.04 ;
      RECT 47.95 -69.85 48.05 -69.04 ;
      RECT 46.75 -69.85 46.85 -69.04 ;
      RECT 45.55 -69.85 45.65 -69.04 ;
      RECT 44.35 -69.85 44.45 -69.04 ;
      RECT 43.15 -69.85 43.25 -69.04 ;
      RECT 41.95 -69.85 42.05 -69.04 ;
      RECT 40.75 -69.85 40.85 -69.04 ;
      RECT 39.55 -69.85 39.65 -69.04 ;
      RECT 38.35 -69.85 38.45 -69.04 ;
      RECT 37.15 -69.85 37.25 -69.04 ;
      RECT 35.95 -69.85 36.05 -69.04 ;
      RECT 34.75 -69.85 34.85 -69.04 ;
      RECT 33.55 -69.85 33.65 -69.04 ;
      RECT 32.35 -69.85 32.45 -69.04 ;
      RECT 31.15 -69.85 31.25 -69.04 ;
      RECT 29.95 -69.85 30.05 -69.04 ;
      RECT 28.75 -69.85 28.85 -69.04 ;
      RECT 27.55 -69.85 27.65 -69.04 ;
      RECT 26.35 -69.85 26.45 -69.04 ;
      RECT 25.15 -69.85 25.25 -69.04 ;
      RECT 23.95 -69.85 24.05 -69.04 ;
      RECT 22.75 -69.85 22.85 -69.04 ;
      RECT 21.55 -69.85 21.65 -69.04 ;
      RECT 20.35 -69.85 20.45 -69.04 ;
      RECT 19.15 -69.85 19.25 -69.04 ;
      RECT 17.95 -69.85 18.05 -69.04 ;
      RECT 16.75 -69.85 16.85 -69.04 ;
      RECT 15.55 -69.85 15.65 -69.04 ;
      RECT 14.35 -69.85 14.45 -69.04 ;
      RECT 13.15 -69.85 13.25 -69.04 ;
      RECT 11.95 -69.85 12.05 -69.04 ;
      RECT 10.75 -69.85 10.85 -69.04 ;
      RECT 9.55 -69.85 9.65 -69.04 ;
      RECT 8.35 -69.85 8.45 -69.04 ;
      RECT 7.15 -69.85 7.25 -69.04 ;
      RECT 5.95 -69.85 6.05 -69.04 ;
      RECT 4.75 -69.85 4.85 -69.04 ;
      RECT 3.55 -69.85 3.65 -69.04 ;
      RECT 2.35 -69.85 2.45 -69.04 ;
      RECT 1.15 -69.85 1.25 -69.04 ;
      RECT -0.05 -69.85 0.05 -69.04 ;
      RECT -0.105 -69.505 156.465 -69.385 ;
      RECT 153.55 -66.62 153.65 -65.81 ;
      RECT 152.35 -66.62 152.45 -65.81 ;
      RECT 151.15 -66.62 151.25 -65.81 ;
      RECT 149.95 -66.62 150.05 -65.81 ;
      RECT 148.75 -66.62 148.85 -65.81 ;
      RECT 147.55 -66.62 147.65 -65.81 ;
      RECT 146.35 -66.62 146.45 -65.81 ;
      RECT 145.15 -66.62 145.25 -65.81 ;
      RECT 143.95 -66.62 144.05 -65.81 ;
      RECT 142.75 -66.62 142.85 -65.81 ;
      RECT 141.55 -66.62 141.65 -65.81 ;
      RECT 140.35 -66.62 140.45 -65.81 ;
      RECT 139.15 -66.62 139.25 -65.81 ;
      RECT 137.95 -66.62 138.05 -65.81 ;
      RECT 136.75 -66.62 136.85 -65.81 ;
      RECT 135.55 -66.62 135.65 -65.81 ;
      RECT 134.35 -66.62 134.45 -65.81 ;
      RECT 133.15 -66.62 133.25 -65.81 ;
      RECT 131.95 -66.62 132.05 -65.81 ;
      RECT 130.75 -66.62 130.85 -65.81 ;
      RECT 129.55 -66.62 129.65 -65.81 ;
      RECT 128.35 -66.62 128.45 -65.81 ;
      RECT 127.15 -66.62 127.25 -65.81 ;
      RECT 125.95 -66.62 126.05 -65.81 ;
      RECT 124.75 -66.62 124.85 -65.81 ;
      RECT 123.55 -66.62 123.65 -65.81 ;
      RECT 122.35 -66.62 122.45 -65.81 ;
      RECT 121.15 -66.62 121.25 -65.81 ;
      RECT 119.95 -66.62 120.05 -65.81 ;
      RECT 118.75 -66.62 118.85 -65.81 ;
      RECT 117.55 -66.62 117.65 -65.81 ;
      RECT 116.35 -66.62 116.45 -65.81 ;
      RECT 115.15 -66.62 115.25 -65.81 ;
      RECT 113.95 -66.62 114.05 -65.81 ;
      RECT 112.75 -66.62 112.85 -65.81 ;
      RECT 111.55 -66.62 111.65 -65.81 ;
      RECT 110.35 -66.62 110.45 -65.81 ;
      RECT 109.15 -66.62 109.25 -65.81 ;
      RECT 107.95 -66.62 108.05 -65.81 ;
      RECT 106.75 -66.62 106.85 -65.81 ;
      RECT 105.55 -66.62 105.65 -65.81 ;
      RECT 104.35 -66.62 104.45 -65.81 ;
      RECT 103.15 -66.62 103.25 -65.81 ;
      RECT 101.95 -66.62 102.05 -65.81 ;
      RECT 100.75 -66.62 100.85 -65.81 ;
      RECT 99.55 -66.62 99.65 -65.81 ;
      RECT 98.35 -66.62 98.45 -65.81 ;
      RECT 97.15 -66.62 97.25 -65.81 ;
      RECT 95.95 -66.62 96.05 -65.81 ;
      RECT 94.75 -66.62 94.85 -65.81 ;
      RECT 93.55 -66.62 93.65 -65.81 ;
      RECT 92.35 -66.62 92.45 -65.81 ;
      RECT 91.15 -66.62 91.25 -65.81 ;
      RECT 89.95 -66.62 90.05 -65.81 ;
      RECT 88.75 -66.62 88.85 -65.81 ;
      RECT 87.55 -66.62 87.65 -65.81 ;
      RECT 86.35 -66.62 86.45 -65.81 ;
      RECT 85.15 -66.62 85.25 -65.81 ;
      RECT 83.95 -66.62 84.05 -65.81 ;
      RECT 82.75 -66.62 82.85 -65.81 ;
      RECT 81.55 -66.62 81.65 -65.81 ;
      RECT 80.35 -66.62 80.45 -65.81 ;
      RECT 79.15 -66.62 79.25 -65.81 ;
      RECT 77.95 -66.62 78.05 -65.81 ;
      RECT 76.75 -66.62 76.85 -65.81 ;
      RECT 75.55 -66.62 75.65 -65.81 ;
      RECT 74.35 -66.62 74.45 -65.81 ;
      RECT 73.15 -66.62 73.25 -65.81 ;
      RECT 71.95 -66.62 72.05 -65.81 ;
      RECT 70.75 -66.62 70.85 -65.81 ;
      RECT 69.55 -66.62 69.65 -65.81 ;
      RECT 68.35 -66.62 68.45 -65.81 ;
      RECT 67.15 -66.62 67.25 -65.81 ;
      RECT 65.95 -66.62 66.05 -65.81 ;
      RECT 64.75 -66.62 64.85 -65.81 ;
      RECT 63.55 -66.62 63.65 -65.81 ;
      RECT 62.35 -66.62 62.45 -65.81 ;
      RECT 61.15 -66.62 61.25 -65.81 ;
      RECT 59.95 -66.62 60.05 -65.81 ;
      RECT 58.75 -66.62 58.85 -65.81 ;
      RECT 57.55 -66.62 57.65 -65.81 ;
      RECT 56.35 -66.62 56.45 -65.81 ;
      RECT 55.15 -66.62 55.25 -65.81 ;
      RECT 53.95 -66.62 54.05 -65.81 ;
      RECT 52.75 -66.62 52.85 -65.81 ;
      RECT 51.55 -66.62 51.65 -65.81 ;
      RECT 50.35 -66.62 50.45 -65.81 ;
      RECT 49.15 -66.62 49.25 -65.81 ;
      RECT 47.95 -66.62 48.05 -65.81 ;
      RECT 46.75 -66.62 46.85 -65.81 ;
      RECT 45.55 -66.62 45.65 -65.81 ;
      RECT 44.35 -66.62 44.45 -65.81 ;
      RECT 43.15 -66.62 43.25 -65.81 ;
      RECT 41.95 -66.62 42.05 -65.81 ;
      RECT 40.75 -66.62 40.85 -65.81 ;
      RECT 39.55 -66.62 39.65 -65.81 ;
      RECT 38.35 -66.62 38.45 -65.81 ;
      RECT 37.15 -66.62 37.25 -65.81 ;
      RECT 35.95 -66.62 36.05 -65.81 ;
      RECT 34.75 -66.62 34.85 -65.81 ;
      RECT 33.55 -66.62 33.65 -65.81 ;
      RECT 32.35 -66.62 32.45 -65.81 ;
      RECT 31.15 -66.62 31.25 -65.81 ;
      RECT 29.95 -66.62 30.05 -65.81 ;
      RECT 28.75 -66.62 28.85 -65.81 ;
      RECT 27.55 -66.62 27.65 -65.81 ;
      RECT 26.35 -66.62 26.45 -65.81 ;
      RECT 25.15 -66.62 25.25 -65.81 ;
      RECT 23.95 -66.62 24.05 -65.81 ;
      RECT 22.75 -66.62 22.85 -65.81 ;
      RECT 21.55 -66.62 21.65 -65.81 ;
      RECT 20.35 -66.62 20.45 -65.81 ;
      RECT 19.15 -66.62 19.25 -65.81 ;
      RECT 17.95 -66.62 18.05 -65.81 ;
      RECT 16.75 -66.62 16.85 -65.81 ;
      RECT 15.55 -66.62 15.65 -65.81 ;
      RECT 14.35 -66.62 14.45 -65.81 ;
      RECT 13.15 -66.62 13.25 -65.81 ;
      RECT 11.95 -66.62 12.05 -65.81 ;
      RECT 10.75 -66.62 10.85 -65.81 ;
      RECT 9.55 -66.62 9.65 -65.81 ;
      RECT 8.35 -66.62 8.45 -65.81 ;
      RECT 7.15 -66.62 7.25 -65.81 ;
      RECT 5.95 -66.62 6.05 -65.81 ;
      RECT 4.75 -66.62 4.85 -65.81 ;
      RECT 3.55 -66.62 3.65 -65.81 ;
      RECT 2.35 -66.62 2.45 -65.81 ;
      RECT 1.15 -66.62 1.25 -65.81 ;
      RECT -0.05 -66.62 0.05 -65.81 ;
      RECT -0.105 -66.275 156.465 -66.155 ;
      RECT 153.55 -63.39 153.65 -62.58 ;
      RECT 152.35 -63.39 152.45 -62.58 ;
      RECT 151.15 -63.39 151.25 -62.58 ;
      RECT 149.95 -63.39 150.05 -62.58 ;
      RECT 148.75 -63.39 148.85 -62.58 ;
      RECT 147.55 -63.39 147.65 -62.58 ;
      RECT 146.35 -63.39 146.45 -62.58 ;
      RECT 145.15 -63.39 145.25 -62.58 ;
      RECT 143.95 -63.39 144.05 -62.58 ;
      RECT 142.75 -63.39 142.85 -62.58 ;
      RECT 141.55 -63.39 141.65 -62.58 ;
      RECT 140.35 -63.39 140.45 -62.58 ;
      RECT 139.15 -63.39 139.25 -62.58 ;
      RECT 137.95 -63.39 138.05 -62.58 ;
      RECT 136.75 -63.39 136.85 -62.58 ;
      RECT 135.55 -63.39 135.65 -62.58 ;
      RECT 134.35 -63.39 134.45 -62.58 ;
      RECT 133.15 -63.39 133.25 -62.58 ;
      RECT 131.95 -63.39 132.05 -62.58 ;
      RECT 130.75 -63.39 130.85 -62.58 ;
      RECT 129.55 -63.39 129.65 -62.58 ;
      RECT 128.35 -63.39 128.45 -62.58 ;
      RECT 127.15 -63.39 127.25 -62.58 ;
      RECT 125.95 -63.39 126.05 -62.58 ;
      RECT 124.75 -63.39 124.85 -62.58 ;
      RECT 123.55 -63.39 123.65 -62.58 ;
      RECT 122.35 -63.39 122.45 -62.58 ;
      RECT 121.15 -63.39 121.25 -62.58 ;
      RECT 119.95 -63.39 120.05 -62.58 ;
      RECT 118.75 -63.39 118.85 -62.58 ;
      RECT 117.55 -63.39 117.65 -62.58 ;
      RECT 116.35 -63.39 116.45 -62.58 ;
      RECT 115.15 -63.39 115.25 -62.58 ;
      RECT 113.95 -63.39 114.05 -62.58 ;
      RECT 112.75 -63.39 112.85 -62.58 ;
      RECT 111.55 -63.39 111.65 -62.58 ;
      RECT 110.35 -63.39 110.45 -62.58 ;
      RECT 109.15 -63.39 109.25 -62.58 ;
      RECT 107.95 -63.39 108.05 -62.58 ;
      RECT 106.75 -63.39 106.85 -62.58 ;
      RECT 105.55 -63.39 105.65 -62.58 ;
      RECT 104.35 -63.39 104.45 -62.58 ;
      RECT 103.15 -63.39 103.25 -62.58 ;
      RECT 101.95 -63.39 102.05 -62.58 ;
      RECT 100.75 -63.39 100.85 -62.58 ;
      RECT 99.55 -63.39 99.65 -62.58 ;
      RECT 98.35 -63.39 98.45 -62.58 ;
      RECT 97.15 -63.39 97.25 -62.58 ;
      RECT 95.95 -63.39 96.05 -62.58 ;
      RECT 94.75 -63.39 94.85 -62.58 ;
      RECT 93.55 -63.39 93.65 -62.58 ;
      RECT 92.35 -63.39 92.45 -62.58 ;
      RECT 91.15 -63.39 91.25 -62.58 ;
      RECT 89.95 -63.39 90.05 -62.58 ;
      RECT 88.75 -63.39 88.85 -62.58 ;
      RECT 87.55 -63.39 87.65 -62.58 ;
      RECT 86.35 -63.39 86.45 -62.58 ;
      RECT 85.15 -63.39 85.25 -62.58 ;
      RECT 83.95 -63.39 84.05 -62.58 ;
      RECT 82.75 -63.39 82.85 -62.58 ;
      RECT 81.55 -63.39 81.65 -62.58 ;
      RECT 80.35 -63.39 80.45 -62.58 ;
      RECT 79.15 -63.39 79.25 -62.58 ;
      RECT 77.95 -63.39 78.05 -62.58 ;
      RECT 76.75 -63.39 76.85 -62.58 ;
      RECT 75.55 -63.39 75.65 -62.58 ;
      RECT 74.35 -63.39 74.45 -62.58 ;
      RECT 73.15 -63.39 73.25 -62.58 ;
      RECT 71.95 -63.39 72.05 -62.58 ;
      RECT 70.75 -63.39 70.85 -62.58 ;
      RECT 69.55 -63.39 69.65 -62.58 ;
      RECT 68.35 -63.39 68.45 -62.58 ;
      RECT 67.15 -63.39 67.25 -62.58 ;
      RECT 65.95 -63.39 66.05 -62.58 ;
      RECT 64.75 -63.39 64.85 -62.58 ;
      RECT 63.55 -63.39 63.65 -62.58 ;
      RECT 62.35 -63.39 62.45 -62.58 ;
      RECT 61.15 -63.39 61.25 -62.58 ;
      RECT 59.95 -63.39 60.05 -62.58 ;
      RECT 58.75 -63.39 58.85 -62.58 ;
      RECT 57.55 -63.39 57.65 -62.58 ;
      RECT 56.35 -63.39 56.45 -62.58 ;
      RECT 55.15 -63.39 55.25 -62.58 ;
      RECT 53.95 -63.39 54.05 -62.58 ;
      RECT 52.75 -63.39 52.85 -62.58 ;
      RECT 51.55 -63.39 51.65 -62.58 ;
      RECT 50.35 -63.39 50.45 -62.58 ;
      RECT 49.15 -63.39 49.25 -62.58 ;
      RECT 47.95 -63.39 48.05 -62.58 ;
      RECT 46.75 -63.39 46.85 -62.58 ;
      RECT 45.55 -63.39 45.65 -62.58 ;
      RECT 44.35 -63.39 44.45 -62.58 ;
      RECT 43.15 -63.39 43.25 -62.58 ;
      RECT 41.95 -63.39 42.05 -62.58 ;
      RECT 40.75 -63.39 40.85 -62.58 ;
      RECT 39.55 -63.39 39.65 -62.58 ;
      RECT 38.35 -63.39 38.45 -62.58 ;
      RECT 37.15 -63.39 37.25 -62.58 ;
      RECT 35.95 -63.39 36.05 -62.58 ;
      RECT 34.75 -63.39 34.85 -62.58 ;
      RECT 33.55 -63.39 33.65 -62.58 ;
      RECT 32.35 -63.39 32.45 -62.58 ;
      RECT 31.15 -63.39 31.25 -62.58 ;
      RECT 29.95 -63.39 30.05 -62.58 ;
      RECT 28.75 -63.39 28.85 -62.58 ;
      RECT 27.55 -63.39 27.65 -62.58 ;
      RECT 26.35 -63.39 26.45 -62.58 ;
      RECT 25.15 -63.39 25.25 -62.58 ;
      RECT 23.95 -63.39 24.05 -62.58 ;
      RECT 22.75 -63.39 22.85 -62.58 ;
      RECT 21.55 -63.39 21.65 -62.58 ;
      RECT 20.35 -63.39 20.45 -62.58 ;
      RECT 19.15 -63.39 19.25 -62.58 ;
      RECT 17.95 -63.39 18.05 -62.58 ;
      RECT 16.75 -63.39 16.85 -62.58 ;
      RECT 15.55 -63.39 15.65 -62.58 ;
      RECT 14.35 -63.39 14.45 -62.58 ;
      RECT 13.15 -63.39 13.25 -62.58 ;
      RECT 11.95 -63.39 12.05 -62.58 ;
      RECT 10.75 -63.39 10.85 -62.58 ;
      RECT 9.55 -63.39 9.65 -62.58 ;
      RECT 8.35 -63.39 8.45 -62.58 ;
      RECT 7.15 -63.39 7.25 -62.58 ;
      RECT 5.95 -63.39 6.05 -62.58 ;
      RECT 4.75 -63.39 4.85 -62.58 ;
      RECT 3.55 -63.39 3.65 -62.58 ;
      RECT 2.35 -63.39 2.45 -62.58 ;
      RECT 1.15 -63.39 1.25 -62.58 ;
      RECT -0.05 -63.39 0.05 -62.58 ;
      RECT -0.105 -63.045 156.465 -62.925 ;
      RECT 153.55 -60.16 153.65 -59.35 ;
      RECT 152.35 -60.16 152.45 -59.35 ;
      RECT 151.15 -60.16 151.25 -59.35 ;
      RECT 149.95 -60.16 150.05 -59.35 ;
      RECT 148.75 -60.16 148.85 -59.35 ;
      RECT 147.55 -60.16 147.65 -59.35 ;
      RECT 146.35 -60.16 146.45 -59.35 ;
      RECT 145.15 -60.16 145.25 -59.35 ;
      RECT 143.95 -60.16 144.05 -59.35 ;
      RECT 142.75 -60.16 142.85 -59.35 ;
      RECT 141.55 -60.16 141.65 -59.35 ;
      RECT 140.35 -60.16 140.45 -59.35 ;
      RECT 139.15 -60.16 139.25 -59.35 ;
      RECT 137.95 -60.16 138.05 -59.35 ;
      RECT 136.75 -60.16 136.85 -59.35 ;
      RECT 135.55 -60.16 135.65 -59.35 ;
      RECT 134.35 -60.16 134.45 -59.35 ;
      RECT 133.15 -60.16 133.25 -59.35 ;
      RECT 131.95 -60.16 132.05 -59.35 ;
      RECT 130.75 -60.16 130.85 -59.35 ;
      RECT 129.55 -60.16 129.65 -59.35 ;
      RECT 128.35 -60.16 128.45 -59.35 ;
      RECT 127.15 -60.16 127.25 -59.35 ;
      RECT 125.95 -60.16 126.05 -59.35 ;
      RECT 124.75 -60.16 124.85 -59.35 ;
      RECT 123.55 -60.16 123.65 -59.35 ;
      RECT 122.35 -60.16 122.45 -59.35 ;
      RECT 121.15 -60.16 121.25 -59.35 ;
      RECT 119.95 -60.16 120.05 -59.35 ;
      RECT 118.75 -60.16 118.85 -59.35 ;
      RECT 117.55 -60.16 117.65 -59.35 ;
      RECT 116.35 -60.16 116.45 -59.35 ;
      RECT 115.15 -60.16 115.25 -59.35 ;
      RECT 113.95 -60.16 114.05 -59.35 ;
      RECT 112.75 -60.16 112.85 -59.35 ;
      RECT 111.55 -60.16 111.65 -59.35 ;
      RECT 110.35 -60.16 110.45 -59.35 ;
      RECT 109.15 -60.16 109.25 -59.35 ;
      RECT 107.95 -60.16 108.05 -59.35 ;
      RECT 106.75 -60.16 106.85 -59.35 ;
      RECT 105.55 -60.16 105.65 -59.35 ;
      RECT 104.35 -60.16 104.45 -59.35 ;
      RECT 103.15 -60.16 103.25 -59.35 ;
      RECT 101.95 -60.16 102.05 -59.35 ;
      RECT 100.75 -60.16 100.85 -59.35 ;
      RECT 99.55 -60.16 99.65 -59.35 ;
      RECT 98.35 -60.16 98.45 -59.35 ;
      RECT 97.15 -60.16 97.25 -59.35 ;
      RECT 95.95 -60.16 96.05 -59.35 ;
      RECT 94.75 -60.16 94.85 -59.35 ;
      RECT 93.55 -60.16 93.65 -59.35 ;
      RECT 92.35 -60.16 92.45 -59.35 ;
      RECT 91.15 -60.16 91.25 -59.35 ;
      RECT 89.95 -60.16 90.05 -59.35 ;
      RECT 88.75 -60.16 88.85 -59.35 ;
      RECT 87.55 -60.16 87.65 -59.35 ;
      RECT 86.35 -60.16 86.45 -59.35 ;
      RECT 85.15 -60.16 85.25 -59.35 ;
      RECT 83.95 -60.16 84.05 -59.35 ;
      RECT 82.75 -60.16 82.85 -59.35 ;
      RECT 81.55 -60.16 81.65 -59.35 ;
      RECT 80.35 -60.16 80.45 -59.35 ;
      RECT 79.15 -60.16 79.25 -59.35 ;
      RECT 77.95 -60.16 78.05 -59.35 ;
      RECT 76.75 -60.16 76.85 -59.35 ;
      RECT 75.55 -60.16 75.65 -59.35 ;
      RECT 74.35 -60.16 74.45 -59.35 ;
      RECT 73.15 -60.16 73.25 -59.35 ;
      RECT 71.95 -60.16 72.05 -59.35 ;
      RECT 70.75 -60.16 70.85 -59.35 ;
      RECT 69.55 -60.16 69.65 -59.35 ;
      RECT 68.35 -60.16 68.45 -59.35 ;
      RECT 67.15 -60.16 67.25 -59.35 ;
      RECT 65.95 -60.16 66.05 -59.35 ;
      RECT 64.75 -60.16 64.85 -59.35 ;
      RECT 63.55 -60.16 63.65 -59.35 ;
      RECT 62.35 -60.16 62.45 -59.35 ;
      RECT 61.15 -60.16 61.25 -59.35 ;
      RECT 59.95 -60.16 60.05 -59.35 ;
      RECT 58.75 -60.16 58.85 -59.35 ;
      RECT 57.55 -60.16 57.65 -59.35 ;
      RECT 56.35 -60.16 56.45 -59.35 ;
      RECT 55.15 -60.16 55.25 -59.35 ;
      RECT 53.95 -60.16 54.05 -59.35 ;
      RECT 52.75 -60.16 52.85 -59.35 ;
      RECT 51.55 -60.16 51.65 -59.35 ;
      RECT 50.35 -60.16 50.45 -59.35 ;
      RECT 49.15 -60.16 49.25 -59.35 ;
      RECT 47.95 -60.16 48.05 -59.35 ;
      RECT 46.75 -60.16 46.85 -59.35 ;
      RECT 45.55 -60.16 45.65 -59.35 ;
      RECT 44.35 -60.16 44.45 -59.35 ;
      RECT 43.15 -60.16 43.25 -59.35 ;
      RECT 41.95 -60.16 42.05 -59.35 ;
      RECT 40.75 -60.16 40.85 -59.35 ;
      RECT 39.55 -60.16 39.65 -59.35 ;
      RECT 38.35 -60.16 38.45 -59.35 ;
      RECT 37.15 -60.16 37.25 -59.35 ;
      RECT 35.95 -60.16 36.05 -59.35 ;
      RECT 34.75 -60.16 34.85 -59.35 ;
      RECT 33.55 -60.16 33.65 -59.35 ;
      RECT 32.35 -60.16 32.45 -59.35 ;
      RECT 31.15 -60.16 31.25 -59.35 ;
      RECT 29.95 -60.16 30.05 -59.35 ;
      RECT 28.75 -60.16 28.85 -59.35 ;
      RECT 27.55 -60.16 27.65 -59.35 ;
      RECT 26.35 -60.16 26.45 -59.35 ;
      RECT 25.15 -60.16 25.25 -59.35 ;
      RECT 23.95 -60.16 24.05 -59.35 ;
      RECT 22.75 -60.16 22.85 -59.35 ;
      RECT 21.55 -60.16 21.65 -59.35 ;
      RECT 20.35 -60.16 20.45 -59.35 ;
      RECT 19.15 -60.16 19.25 -59.35 ;
      RECT 17.95 -60.16 18.05 -59.35 ;
      RECT 16.75 -60.16 16.85 -59.35 ;
      RECT 15.55 -60.16 15.65 -59.35 ;
      RECT 14.35 -60.16 14.45 -59.35 ;
      RECT 13.15 -60.16 13.25 -59.35 ;
      RECT 11.95 -60.16 12.05 -59.35 ;
      RECT 10.75 -60.16 10.85 -59.35 ;
      RECT 9.55 -60.16 9.65 -59.35 ;
      RECT 8.35 -60.16 8.45 -59.35 ;
      RECT 7.15 -60.16 7.25 -59.35 ;
      RECT 5.95 -60.16 6.05 -59.35 ;
      RECT 4.75 -60.16 4.85 -59.35 ;
      RECT 3.55 -60.16 3.65 -59.35 ;
      RECT 2.35 -60.16 2.45 -59.35 ;
      RECT 1.15 -60.16 1.25 -59.35 ;
      RECT -0.05 -60.16 0.05 -59.35 ;
      RECT -0.105 -59.815 156.465 -59.695 ;
      RECT 153.55 -56.93 153.65 -56.12 ;
      RECT 152.35 -56.93 152.45 -56.12 ;
      RECT 151.15 -56.93 151.25 -56.12 ;
      RECT 149.95 -56.93 150.05 -56.12 ;
      RECT 148.75 -56.93 148.85 -56.12 ;
      RECT 147.55 -56.93 147.65 -56.12 ;
      RECT 146.35 -56.93 146.45 -56.12 ;
      RECT 145.15 -56.93 145.25 -56.12 ;
      RECT 143.95 -56.93 144.05 -56.12 ;
      RECT 142.75 -56.93 142.85 -56.12 ;
      RECT 141.55 -56.93 141.65 -56.12 ;
      RECT 140.35 -56.93 140.45 -56.12 ;
      RECT 139.15 -56.93 139.25 -56.12 ;
      RECT 137.95 -56.93 138.05 -56.12 ;
      RECT 136.75 -56.93 136.85 -56.12 ;
      RECT 135.55 -56.93 135.65 -56.12 ;
      RECT 134.35 -56.93 134.45 -56.12 ;
      RECT 133.15 -56.93 133.25 -56.12 ;
      RECT 131.95 -56.93 132.05 -56.12 ;
      RECT 130.75 -56.93 130.85 -56.12 ;
      RECT 129.55 -56.93 129.65 -56.12 ;
      RECT 128.35 -56.93 128.45 -56.12 ;
      RECT 127.15 -56.93 127.25 -56.12 ;
      RECT 125.95 -56.93 126.05 -56.12 ;
      RECT 124.75 -56.93 124.85 -56.12 ;
      RECT 123.55 -56.93 123.65 -56.12 ;
      RECT 122.35 -56.93 122.45 -56.12 ;
      RECT 121.15 -56.93 121.25 -56.12 ;
      RECT 119.95 -56.93 120.05 -56.12 ;
      RECT 118.75 -56.93 118.85 -56.12 ;
      RECT 117.55 -56.93 117.65 -56.12 ;
      RECT 116.35 -56.93 116.45 -56.12 ;
      RECT 115.15 -56.93 115.25 -56.12 ;
      RECT 113.95 -56.93 114.05 -56.12 ;
      RECT 112.75 -56.93 112.85 -56.12 ;
      RECT 111.55 -56.93 111.65 -56.12 ;
      RECT 110.35 -56.93 110.45 -56.12 ;
      RECT 109.15 -56.93 109.25 -56.12 ;
      RECT 107.95 -56.93 108.05 -56.12 ;
      RECT 106.75 -56.93 106.85 -56.12 ;
      RECT 105.55 -56.93 105.65 -56.12 ;
      RECT 104.35 -56.93 104.45 -56.12 ;
      RECT 103.15 -56.93 103.25 -56.12 ;
      RECT 101.95 -56.93 102.05 -56.12 ;
      RECT 100.75 -56.93 100.85 -56.12 ;
      RECT 99.55 -56.93 99.65 -56.12 ;
      RECT 98.35 -56.93 98.45 -56.12 ;
      RECT 97.15 -56.93 97.25 -56.12 ;
      RECT 95.95 -56.93 96.05 -56.12 ;
      RECT 94.75 -56.93 94.85 -56.12 ;
      RECT 93.55 -56.93 93.65 -56.12 ;
      RECT 92.35 -56.93 92.45 -56.12 ;
      RECT 91.15 -56.93 91.25 -56.12 ;
      RECT 89.95 -56.93 90.05 -56.12 ;
      RECT 88.75 -56.93 88.85 -56.12 ;
      RECT 87.55 -56.93 87.65 -56.12 ;
      RECT 86.35 -56.93 86.45 -56.12 ;
      RECT 85.15 -56.93 85.25 -56.12 ;
      RECT 83.95 -56.93 84.05 -56.12 ;
      RECT 82.75 -56.93 82.85 -56.12 ;
      RECT 81.55 -56.93 81.65 -56.12 ;
      RECT 80.35 -56.93 80.45 -56.12 ;
      RECT 79.15 -56.93 79.25 -56.12 ;
      RECT 77.95 -56.93 78.05 -56.12 ;
      RECT 76.75 -56.93 76.85 -56.12 ;
      RECT 75.55 -56.93 75.65 -56.12 ;
      RECT 74.35 -56.93 74.45 -56.12 ;
      RECT 73.15 -56.93 73.25 -56.12 ;
      RECT 71.95 -56.93 72.05 -56.12 ;
      RECT 70.75 -56.93 70.85 -56.12 ;
      RECT 69.55 -56.93 69.65 -56.12 ;
      RECT 68.35 -56.93 68.45 -56.12 ;
      RECT 67.15 -56.93 67.25 -56.12 ;
      RECT 65.95 -56.93 66.05 -56.12 ;
      RECT 64.75 -56.93 64.85 -56.12 ;
      RECT 63.55 -56.93 63.65 -56.12 ;
      RECT 62.35 -56.93 62.45 -56.12 ;
      RECT 61.15 -56.93 61.25 -56.12 ;
      RECT 59.95 -56.93 60.05 -56.12 ;
      RECT 58.75 -56.93 58.85 -56.12 ;
      RECT 57.55 -56.93 57.65 -56.12 ;
      RECT 56.35 -56.93 56.45 -56.12 ;
      RECT 55.15 -56.93 55.25 -56.12 ;
      RECT 53.95 -56.93 54.05 -56.12 ;
      RECT 52.75 -56.93 52.85 -56.12 ;
      RECT 51.55 -56.93 51.65 -56.12 ;
      RECT 50.35 -56.93 50.45 -56.12 ;
      RECT 49.15 -56.93 49.25 -56.12 ;
      RECT 47.95 -56.93 48.05 -56.12 ;
      RECT 46.75 -56.93 46.85 -56.12 ;
      RECT 45.55 -56.93 45.65 -56.12 ;
      RECT 44.35 -56.93 44.45 -56.12 ;
      RECT 43.15 -56.93 43.25 -56.12 ;
      RECT 41.95 -56.93 42.05 -56.12 ;
      RECT 40.75 -56.93 40.85 -56.12 ;
      RECT 39.55 -56.93 39.65 -56.12 ;
      RECT 38.35 -56.93 38.45 -56.12 ;
      RECT 37.15 -56.93 37.25 -56.12 ;
      RECT 35.95 -56.93 36.05 -56.12 ;
      RECT 34.75 -56.93 34.85 -56.12 ;
      RECT 33.55 -56.93 33.65 -56.12 ;
      RECT 32.35 -56.93 32.45 -56.12 ;
      RECT 31.15 -56.93 31.25 -56.12 ;
      RECT 29.95 -56.93 30.05 -56.12 ;
      RECT 28.75 -56.93 28.85 -56.12 ;
      RECT 27.55 -56.93 27.65 -56.12 ;
      RECT 26.35 -56.93 26.45 -56.12 ;
      RECT 25.15 -56.93 25.25 -56.12 ;
      RECT 23.95 -56.93 24.05 -56.12 ;
      RECT 22.75 -56.93 22.85 -56.12 ;
      RECT 21.55 -56.93 21.65 -56.12 ;
      RECT 20.35 -56.93 20.45 -56.12 ;
      RECT 19.15 -56.93 19.25 -56.12 ;
      RECT 17.95 -56.93 18.05 -56.12 ;
      RECT 16.75 -56.93 16.85 -56.12 ;
      RECT 15.55 -56.93 15.65 -56.12 ;
      RECT 14.35 -56.93 14.45 -56.12 ;
      RECT 13.15 -56.93 13.25 -56.12 ;
      RECT 11.95 -56.93 12.05 -56.12 ;
      RECT 10.75 -56.93 10.85 -56.12 ;
      RECT 9.55 -56.93 9.65 -56.12 ;
      RECT 8.35 -56.93 8.45 -56.12 ;
      RECT 7.15 -56.93 7.25 -56.12 ;
      RECT 5.95 -56.93 6.05 -56.12 ;
      RECT 4.75 -56.93 4.85 -56.12 ;
      RECT 3.55 -56.93 3.65 -56.12 ;
      RECT 2.35 -56.93 2.45 -56.12 ;
      RECT 1.15 -56.93 1.25 -56.12 ;
      RECT -0.05 -56.93 0.05 -56.12 ;
      RECT -0.105 -56.585 156.465 -56.465 ;
      RECT 153.55 -53.7 153.65 -52.89 ;
      RECT 152.35 -53.7 152.45 -52.89 ;
      RECT 151.15 -53.7 151.25 -52.89 ;
      RECT 149.95 -53.7 150.05 -52.89 ;
      RECT 148.75 -53.7 148.85 -52.89 ;
      RECT 147.55 -53.7 147.65 -52.89 ;
      RECT 146.35 -53.7 146.45 -52.89 ;
      RECT 145.15 -53.7 145.25 -52.89 ;
      RECT 143.95 -53.7 144.05 -52.89 ;
      RECT 142.75 -53.7 142.85 -52.89 ;
      RECT 141.55 -53.7 141.65 -52.89 ;
      RECT 140.35 -53.7 140.45 -52.89 ;
      RECT 139.15 -53.7 139.25 -52.89 ;
      RECT 137.95 -53.7 138.05 -52.89 ;
      RECT 136.75 -53.7 136.85 -52.89 ;
      RECT 135.55 -53.7 135.65 -52.89 ;
      RECT 134.35 -53.7 134.45 -52.89 ;
      RECT 133.15 -53.7 133.25 -52.89 ;
      RECT 131.95 -53.7 132.05 -52.89 ;
      RECT 130.75 -53.7 130.85 -52.89 ;
      RECT 129.55 -53.7 129.65 -52.89 ;
      RECT 128.35 -53.7 128.45 -52.89 ;
      RECT 127.15 -53.7 127.25 -52.89 ;
      RECT 125.95 -53.7 126.05 -52.89 ;
      RECT 124.75 -53.7 124.85 -52.89 ;
      RECT 123.55 -53.7 123.65 -52.89 ;
      RECT 122.35 -53.7 122.45 -52.89 ;
      RECT 121.15 -53.7 121.25 -52.89 ;
      RECT 119.95 -53.7 120.05 -52.89 ;
      RECT 118.75 -53.7 118.85 -52.89 ;
      RECT 117.55 -53.7 117.65 -52.89 ;
      RECT 116.35 -53.7 116.45 -52.89 ;
      RECT 115.15 -53.7 115.25 -52.89 ;
      RECT 113.95 -53.7 114.05 -52.89 ;
      RECT 112.75 -53.7 112.85 -52.89 ;
      RECT 111.55 -53.7 111.65 -52.89 ;
      RECT 110.35 -53.7 110.45 -52.89 ;
      RECT 109.15 -53.7 109.25 -52.89 ;
      RECT 107.95 -53.7 108.05 -52.89 ;
      RECT 106.75 -53.7 106.85 -52.89 ;
      RECT 105.55 -53.7 105.65 -52.89 ;
      RECT 104.35 -53.7 104.45 -52.89 ;
      RECT 103.15 -53.7 103.25 -52.89 ;
      RECT 101.95 -53.7 102.05 -52.89 ;
      RECT 100.75 -53.7 100.85 -52.89 ;
      RECT 99.55 -53.7 99.65 -52.89 ;
      RECT 98.35 -53.7 98.45 -52.89 ;
      RECT 97.15 -53.7 97.25 -52.89 ;
      RECT 95.95 -53.7 96.05 -52.89 ;
      RECT 94.75 -53.7 94.85 -52.89 ;
      RECT 93.55 -53.7 93.65 -52.89 ;
      RECT 92.35 -53.7 92.45 -52.89 ;
      RECT 91.15 -53.7 91.25 -52.89 ;
      RECT 89.95 -53.7 90.05 -52.89 ;
      RECT 88.75 -53.7 88.85 -52.89 ;
      RECT 87.55 -53.7 87.65 -52.89 ;
      RECT 86.35 -53.7 86.45 -52.89 ;
      RECT 85.15 -53.7 85.25 -52.89 ;
      RECT 83.95 -53.7 84.05 -52.89 ;
      RECT 82.75 -53.7 82.85 -52.89 ;
      RECT 81.55 -53.7 81.65 -52.89 ;
      RECT 80.35 -53.7 80.45 -52.89 ;
      RECT 79.15 -53.7 79.25 -52.89 ;
      RECT 77.95 -53.7 78.05 -52.89 ;
      RECT 76.75 -53.7 76.85 -52.89 ;
      RECT 75.55 -53.7 75.65 -52.89 ;
      RECT 74.35 -53.7 74.45 -52.89 ;
      RECT 73.15 -53.7 73.25 -52.89 ;
      RECT 71.95 -53.7 72.05 -52.89 ;
      RECT 70.75 -53.7 70.85 -52.89 ;
      RECT 69.55 -53.7 69.65 -52.89 ;
      RECT 68.35 -53.7 68.45 -52.89 ;
      RECT 67.15 -53.7 67.25 -52.89 ;
      RECT 65.95 -53.7 66.05 -52.89 ;
      RECT 64.75 -53.7 64.85 -52.89 ;
      RECT 63.55 -53.7 63.65 -52.89 ;
      RECT 62.35 -53.7 62.45 -52.89 ;
      RECT 61.15 -53.7 61.25 -52.89 ;
      RECT 59.95 -53.7 60.05 -52.89 ;
      RECT 58.75 -53.7 58.85 -52.89 ;
      RECT 57.55 -53.7 57.65 -52.89 ;
      RECT 56.35 -53.7 56.45 -52.89 ;
      RECT 55.15 -53.7 55.25 -52.89 ;
      RECT 53.95 -53.7 54.05 -52.89 ;
      RECT 52.75 -53.7 52.85 -52.89 ;
      RECT 51.55 -53.7 51.65 -52.89 ;
      RECT 50.35 -53.7 50.45 -52.89 ;
      RECT 49.15 -53.7 49.25 -52.89 ;
      RECT 47.95 -53.7 48.05 -52.89 ;
      RECT 46.75 -53.7 46.85 -52.89 ;
      RECT 45.55 -53.7 45.65 -52.89 ;
      RECT 44.35 -53.7 44.45 -52.89 ;
      RECT 43.15 -53.7 43.25 -52.89 ;
      RECT 41.95 -53.7 42.05 -52.89 ;
      RECT 40.75 -53.7 40.85 -52.89 ;
      RECT 39.55 -53.7 39.65 -52.89 ;
      RECT 38.35 -53.7 38.45 -52.89 ;
      RECT 37.15 -53.7 37.25 -52.89 ;
      RECT 35.95 -53.7 36.05 -52.89 ;
      RECT 34.75 -53.7 34.85 -52.89 ;
      RECT 33.55 -53.7 33.65 -52.89 ;
      RECT 32.35 -53.7 32.45 -52.89 ;
      RECT 31.15 -53.7 31.25 -52.89 ;
      RECT 29.95 -53.7 30.05 -52.89 ;
      RECT 28.75 -53.7 28.85 -52.89 ;
      RECT 27.55 -53.7 27.65 -52.89 ;
      RECT 26.35 -53.7 26.45 -52.89 ;
      RECT 25.15 -53.7 25.25 -52.89 ;
      RECT 23.95 -53.7 24.05 -52.89 ;
      RECT 22.75 -53.7 22.85 -52.89 ;
      RECT 21.55 -53.7 21.65 -52.89 ;
      RECT 20.35 -53.7 20.45 -52.89 ;
      RECT 19.15 -53.7 19.25 -52.89 ;
      RECT 17.95 -53.7 18.05 -52.89 ;
      RECT 16.75 -53.7 16.85 -52.89 ;
      RECT 15.55 -53.7 15.65 -52.89 ;
      RECT 14.35 -53.7 14.45 -52.89 ;
      RECT 13.15 -53.7 13.25 -52.89 ;
      RECT 11.95 -53.7 12.05 -52.89 ;
      RECT 10.75 -53.7 10.85 -52.89 ;
      RECT 9.55 -53.7 9.65 -52.89 ;
      RECT 8.35 -53.7 8.45 -52.89 ;
      RECT 7.15 -53.7 7.25 -52.89 ;
      RECT 5.95 -53.7 6.05 -52.89 ;
      RECT 4.75 -53.7 4.85 -52.89 ;
      RECT 3.55 -53.7 3.65 -52.89 ;
      RECT 2.35 -53.7 2.45 -52.89 ;
      RECT 1.15 -53.7 1.25 -52.89 ;
      RECT -0.05 -53.7 0.05 -52.89 ;
      RECT -0.105 -53.355 156.465 -53.235 ;
      RECT 153.55 -50.47 153.65 -49.66 ;
      RECT 152.35 -50.47 152.45 -49.66 ;
      RECT 151.15 -50.47 151.25 -49.66 ;
      RECT 149.95 -50.47 150.05 -49.66 ;
      RECT 148.75 -50.47 148.85 -49.66 ;
      RECT 147.55 -50.47 147.65 -49.66 ;
      RECT 146.35 -50.47 146.45 -49.66 ;
      RECT 145.15 -50.47 145.25 -49.66 ;
      RECT 143.95 -50.47 144.05 -49.66 ;
      RECT 142.75 -50.47 142.85 -49.66 ;
      RECT 141.55 -50.47 141.65 -49.66 ;
      RECT 140.35 -50.47 140.45 -49.66 ;
      RECT 139.15 -50.47 139.25 -49.66 ;
      RECT 137.95 -50.47 138.05 -49.66 ;
      RECT 136.75 -50.47 136.85 -49.66 ;
      RECT 135.55 -50.47 135.65 -49.66 ;
      RECT 134.35 -50.47 134.45 -49.66 ;
      RECT 133.15 -50.47 133.25 -49.66 ;
      RECT 131.95 -50.47 132.05 -49.66 ;
      RECT 130.75 -50.47 130.85 -49.66 ;
      RECT 129.55 -50.47 129.65 -49.66 ;
      RECT 128.35 -50.47 128.45 -49.66 ;
      RECT 127.15 -50.47 127.25 -49.66 ;
      RECT 125.95 -50.47 126.05 -49.66 ;
      RECT 124.75 -50.47 124.85 -49.66 ;
      RECT 123.55 -50.47 123.65 -49.66 ;
      RECT 122.35 -50.47 122.45 -49.66 ;
      RECT 121.15 -50.47 121.25 -49.66 ;
      RECT 119.95 -50.47 120.05 -49.66 ;
      RECT 118.75 -50.47 118.85 -49.66 ;
      RECT 117.55 -50.47 117.65 -49.66 ;
      RECT 116.35 -50.47 116.45 -49.66 ;
      RECT 115.15 -50.47 115.25 -49.66 ;
      RECT 113.95 -50.47 114.05 -49.66 ;
      RECT 112.75 -50.47 112.85 -49.66 ;
      RECT 111.55 -50.47 111.65 -49.66 ;
      RECT 110.35 -50.47 110.45 -49.66 ;
      RECT 109.15 -50.47 109.25 -49.66 ;
      RECT 107.95 -50.47 108.05 -49.66 ;
      RECT 106.75 -50.47 106.85 -49.66 ;
      RECT 105.55 -50.47 105.65 -49.66 ;
      RECT 104.35 -50.47 104.45 -49.66 ;
      RECT 103.15 -50.47 103.25 -49.66 ;
      RECT 101.95 -50.47 102.05 -49.66 ;
      RECT 100.75 -50.47 100.85 -49.66 ;
      RECT 99.55 -50.47 99.65 -49.66 ;
      RECT 98.35 -50.47 98.45 -49.66 ;
      RECT 97.15 -50.47 97.25 -49.66 ;
      RECT 95.95 -50.47 96.05 -49.66 ;
      RECT 94.75 -50.47 94.85 -49.66 ;
      RECT 93.55 -50.47 93.65 -49.66 ;
      RECT 92.35 -50.47 92.45 -49.66 ;
      RECT 91.15 -50.47 91.25 -49.66 ;
      RECT 89.95 -50.47 90.05 -49.66 ;
      RECT 88.75 -50.47 88.85 -49.66 ;
      RECT 87.55 -50.47 87.65 -49.66 ;
      RECT 86.35 -50.47 86.45 -49.66 ;
      RECT 85.15 -50.47 85.25 -49.66 ;
      RECT 83.95 -50.47 84.05 -49.66 ;
      RECT 82.75 -50.47 82.85 -49.66 ;
      RECT 81.55 -50.47 81.65 -49.66 ;
      RECT 80.35 -50.47 80.45 -49.66 ;
      RECT 79.15 -50.47 79.25 -49.66 ;
      RECT 77.95 -50.47 78.05 -49.66 ;
      RECT 76.75 -50.47 76.85 -49.66 ;
      RECT 75.55 -50.47 75.65 -49.66 ;
      RECT 74.35 -50.47 74.45 -49.66 ;
      RECT 73.15 -50.47 73.25 -49.66 ;
      RECT 71.95 -50.47 72.05 -49.66 ;
      RECT 70.75 -50.47 70.85 -49.66 ;
      RECT 69.55 -50.47 69.65 -49.66 ;
      RECT 68.35 -50.47 68.45 -49.66 ;
      RECT 67.15 -50.47 67.25 -49.66 ;
      RECT 65.95 -50.47 66.05 -49.66 ;
      RECT 64.75 -50.47 64.85 -49.66 ;
      RECT 63.55 -50.47 63.65 -49.66 ;
      RECT 62.35 -50.47 62.45 -49.66 ;
      RECT 61.15 -50.47 61.25 -49.66 ;
      RECT 59.95 -50.47 60.05 -49.66 ;
      RECT 58.75 -50.47 58.85 -49.66 ;
      RECT 57.55 -50.47 57.65 -49.66 ;
      RECT 56.35 -50.47 56.45 -49.66 ;
      RECT 55.15 -50.47 55.25 -49.66 ;
      RECT 53.95 -50.47 54.05 -49.66 ;
      RECT 52.75 -50.47 52.85 -49.66 ;
      RECT 51.55 -50.47 51.65 -49.66 ;
      RECT 50.35 -50.47 50.45 -49.66 ;
      RECT 49.15 -50.47 49.25 -49.66 ;
      RECT 47.95 -50.47 48.05 -49.66 ;
      RECT 46.75 -50.47 46.85 -49.66 ;
      RECT 45.55 -50.47 45.65 -49.66 ;
      RECT 44.35 -50.47 44.45 -49.66 ;
      RECT 43.15 -50.47 43.25 -49.66 ;
      RECT 41.95 -50.47 42.05 -49.66 ;
      RECT 40.75 -50.47 40.85 -49.66 ;
      RECT 39.55 -50.47 39.65 -49.66 ;
      RECT 38.35 -50.47 38.45 -49.66 ;
      RECT 37.15 -50.47 37.25 -49.66 ;
      RECT 35.95 -50.47 36.05 -49.66 ;
      RECT 34.75 -50.47 34.85 -49.66 ;
      RECT 33.55 -50.47 33.65 -49.66 ;
      RECT 32.35 -50.47 32.45 -49.66 ;
      RECT 31.15 -50.47 31.25 -49.66 ;
      RECT 29.95 -50.47 30.05 -49.66 ;
      RECT 28.75 -50.47 28.85 -49.66 ;
      RECT 27.55 -50.47 27.65 -49.66 ;
      RECT 26.35 -50.47 26.45 -49.66 ;
      RECT 25.15 -50.47 25.25 -49.66 ;
      RECT 23.95 -50.47 24.05 -49.66 ;
      RECT 22.75 -50.47 22.85 -49.66 ;
      RECT 21.55 -50.47 21.65 -49.66 ;
      RECT 20.35 -50.47 20.45 -49.66 ;
      RECT 19.15 -50.47 19.25 -49.66 ;
      RECT 17.95 -50.47 18.05 -49.66 ;
      RECT 16.75 -50.47 16.85 -49.66 ;
      RECT 15.55 -50.47 15.65 -49.66 ;
      RECT 14.35 -50.47 14.45 -49.66 ;
      RECT 13.15 -50.47 13.25 -49.66 ;
      RECT 11.95 -50.47 12.05 -49.66 ;
      RECT 10.75 -50.47 10.85 -49.66 ;
      RECT 9.55 -50.47 9.65 -49.66 ;
      RECT 8.35 -50.47 8.45 -49.66 ;
      RECT 7.15 -50.47 7.25 -49.66 ;
      RECT 5.95 -50.47 6.05 -49.66 ;
      RECT 4.75 -50.47 4.85 -49.66 ;
      RECT 3.55 -50.47 3.65 -49.66 ;
      RECT 2.35 -50.47 2.45 -49.66 ;
      RECT 1.15 -50.47 1.25 -49.66 ;
      RECT -0.05 -50.47 0.05 -49.66 ;
      RECT -0.105 -50.125 156.465 -50.005 ;
      RECT 153.55 -47.24 153.65 -46.43 ;
      RECT 152.35 -47.24 152.45 -46.43 ;
      RECT 151.15 -47.24 151.25 -46.43 ;
      RECT 149.95 -47.24 150.05 -46.43 ;
      RECT 148.75 -47.24 148.85 -46.43 ;
      RECT 147.55 -47.24 147.65 -46.43 ;
      RECT 146.35 -47.24 146.45 -46.43 ;
      RECT 145.15 -47.24 145.25 -46.43 ;
      RECT 143.95 -47.24 144.05 -46.43 ;
      RECT 142.75 -47.24 142.85 -46.43 ;
      RECT 141.55 -47.24 141.65 -46.43 ;
      RECT 140.35 -47.24 140.45 -46.43 ;
      RECT 139.15 -47.24 139.25 -46.43 ;
      RECT 137.95 -47.24 138.05 -46.43 ;
      RECT 136.75 -47.24 136.85 -46.43 ;
      RECT 135.55 -47.24 135.65 -46.43 ;
      RECT 134.35 -47.24 134.45 -46.43 ;
      RECT 133.15 -47.24 133.25 -46.43 ;
      RECT 131.95 -47.24 132.05 -46.43 ;
      RECT 130.75 -47.24 130.85 -46.43 ;
      RECT 129.55 -47.24 129.65 -46.43 ;
      RECT 128.35 -47.24 128.45 -46.43 ;
      RECT 127.15 -47.24 127.25 -46.43 ;
      RECT 125.95 -47.24 126.05 -46.43 ;
      RECT 124.75 -47.24 124.85 -46.43 ;
      RECT 123.55 -47.24 123.65 -46.43 ;
      RECT 122.35 -47.24 122.45 -46.43 ;
      RECT 121.15 -47.24 121.25 -46.43 ;
      RECT 119.95 -47.24 120.05 -46.43 ;
      RECT 118.75 -47.24 118.85 -46.43 ;
      RECT 117.55 -47.24 117.65 -46.43 ;
      RECT 116.35 -47.24 116.45 -46.43 ;
      RECT 115.15 -47.24 115.25 -46.43 ;
      RECT 113.95 -47.24 114.05 -46.43 ;
      RECT 112.75 -47.24 112.85 -46.43 ;
      RECT 111.55 -47.24 111.65 -46.43 ;
      RECT 110.35 -47.24 110.45 -46.43 ;
      RECT 109.15 -47.24 109.25 -46.43 ;
      RECT 107.95 -47.24 108.05 -46.43 ;
      RECT 106.75 -47.24 106.85 -46.43 ;
      RECT 105.55 -47.24 105.65 -46.43 ;
      RECT 104.35 -47.24 104.45 -46.43 ;
      RECT 103.15 -47.24 103.25 -46.43 ;
      RECT 101.95 -47.24 102.05 -46.43 ;
      RECT 100.75 -47.24 100.85 -46.43 ;
      RECT 99.55 -47.24 99.65 -46.43 ;
      RECT 98.35 -47.24 98.45 -46.43 ;
      RECT 97.15 -47.24 97.25 -46.43 ;
      RECT 95.95 -47.24 96.05 -46.43 ;
      RECT 94.75 -47.24 94.85 -46.43 ;
      RECT 93.55 -47.24 93.65 -46.43 ;
      RECT 92.35 -47.24 92.45 -46.43 ;
      RECT 91.15 -47.24 91.25 -46.43 ;
      RECT 89.95 -47.24 90.05 -46.43 ;
      RECT 88.75 -47.24 88.85 -46.43 ;
      RECT 87.55 -47.24 87.65 -46.43 ;
      RECT 86.35 -47.24 86.45 -46.43 ;
      RECT 85.15 -47.24 85.25 -46.43 ;
      RECT 83.95 -47.24 84.05 -46.43 ;
      RECT 82.75 -47.24 82.85 -46.43 ;
      RECT 81.55 -47.24 81.65 -46.43 ;
      RECT 80.35 -47.24 80.45 -46.43 ;
      RECT 79.15 -47.24 79.25 -46.43 ;
      RECT 77.95 -47.24 78.05 -46.43 ;
      RECT 76.75 -47.24 76.85 -46.43 ;
      RECT 75.55 -47.24 75.65 -46.43 ;
      RECT 74.35 -47.24 74.45 -46.43 ;
      RECT 73.15 -47.24 73.25 -46.43 ;
      RECT 71.95 -47.24 72.05 -46.43 ;
      RECT 70.75 -47.24 70.85 -46.43 ;
      RECT 69.55 -47.24 69.65 -46.43 ;
      RECT 68.35 -47.24 68.45 -46.43 ;
      RECT 67.15 -47.24 67.25 -46.43 ;
      RECT 65.95 -47.24 66.05 -46.43 ;
      RECT 64.75 -47.24 64.85 -46.43 ;
      RECT 63.55 -47.24 63.65 -46.43 ;
      RECT 62.35 -47.24 62.45 -46.43 ;
      RECT 61.15 -47.24 61.25 -46.43 ;
      RECT 59.95 -47.24 60.05 -46.43 ;
      RECT 58.75 -47.24 58.85 -46.43 ;
      RECT 57.55 -47.24 57.65 -46.43 ;
      RECT 56.35 -47.24 56.45 -46.43 ;
      RECT 55.15 -47.24 55.25 -46.43 ;
      RECT 53.95 -47.24 54.05 -46.43 ;
      RECT 52.75 -47.24 52.85 -46.43 ;
      RECT 51.55 -47.24 51.65 -46.43 ;
      RECT 50.35 -47.24 50.45 -46.43 ;
      RECT 49.15 -47.24 49.25 -46.43 ;
      RECT 47.95 -47.24 48.05 -46.43 ;
      RECT 46.75 -47.24 46.85 -46.43 ;
      RECT 45.55 -47.24 45.65 -46.43 ;
      RECT 44.35 -47.24 44.45 -46.43 ;
      RECT 43.15 -47.24 43.25 -46.43 ;
      RECT 41.95 -47.24 42.05 -46.43 ;
      RECT 40.75 -47.24 40.85 -46.43 ;
      RECT 39.55 -47.24 39.65 -46.43 ;
      RECT 38.35 -47.24 38.45 -46.43 ;
      RECT 37.15 -47.24 37.25 -46.43 ;
      RECT 35.95 -47.24 36.05 -46.43 ;
      RECT 34.75 -47.24 34.85 -46.43 ;
      RECT 33.55 -47.24 33.65 -46.43 ;
      RECT 32.35 -47.24 32.45 -46.43 ;
      RECT 31.15 -47.24 31.25 -46.43 ;
      RECT 29.95 -47.24 30.05 -46.43 ;
      RECT 28.75 -47.24 28.85 -46.43 ;
      RECT 27.55 -47.24 27.65 -46.43 ;
      RECT 26.35 -47.24 26.45 -46.43 ;
      RECT 25.15 -47.24 25.25 -46.43 ;
      RECT 23.95 -47.24 24.05 -46.43 ;
      RECT 22.75 -47.24 22.85 -46.43 ;
      RECT 21.55 -47.24 21.65 -46.43 ;
      RECT 20.35 -47.24 20.45 -46.43 ;
      RECT 19.15 -47.24 19.25 -46.43 ;
      RECT 17.95 -47.24 18.05 -46.43 ;
      RECT 16.75 -47.24 16.85 -46.43 ;
      RECT 15.55 -47.24 15.65 -46.43 ;
      RECT 14.35 -47.24 14.45 -46.43 ;
      RECT 13.15 -47.24 13.25 -46.43 ;
      RECT 11.95 -47.24 12.05 -46.43 ;
      RECT 10.75 -47.24 10.85 -46.43 ;
      RECT 9.55 -47.24 9.65 -46.43 ;
      RECT 8.35 -47.24 8.45 -46.43 ;
      RECT 7.15 -47.24 7.25 -46.43 ;
      RECT 5.95 -47.24 6.05 -46.43 ;
      RECT 4.75 -47.24 4.85 -46.43 ;
      RECT 3.55 -47.24 3.65 -46.43 ;
      RECT 2.35 -47.24 2.45 -46.43 ;
      RECT 1.15 -47.24 1.25 -46.43 ;
      RECT -0.05 -47.24 0.05 -46.43 ;
      RECT -0.105 -46.895 156.465 -46.775 ;
      RECT 153.55 -44.01 153.65 -43.2 ;
      RECT 152.35 -44.01 152.45 -43.2 ;
      RECT 151.15 -44.01 151.25 -43.2 ;
      RECT 149.95 -44.01 150.05 -43.2 ;
      RECT 148.75 -44.01 148.85 -43.2 ;
      RECT 147.55 -44.01 147.65 -43.2 ;
      RECT 146.35 -44.01 146.45 -43.2 ;
      RECT 145.15 -44.01 145.25 -43.2 ;
      RECT 143.95 -44.01 144.05 -43.2 ;
      RECT 142.75 -44.01 142.85 -43.2 ;
      RECT 141.55 -44.01 141.65 -43.2 ;
      RECT 140.35 -44.01 140.45 -43.2 ;
      RECT 139.15 -44.01 139.25 -43.2 ;
      RECT 137.95 -44.01 138.05 -43.2 ;
      RECT 136.75 -44.01 136.85 -43.2 ;
      RECT 135.55 -44.01 135.65 -43.2 ;
      RECT 134.35 -44.01 134.45 -43.2 ;
      RECT 133.15 -44.01 133.25 -43.2 ;
      RECT 131.95 -44.01 132.05 -43.2 ;
      RECT 130.75 -44.01 130.85 -43.2 ;
      RECT 129.55 -44.01 129.65 -43.2 ;
      RECT 128.35 -44.01 128.45 -43.2 ;
      RECT 127.15 -44.01 127.25 -43.2 ;
      RECT 125.95 -44.01 126.05 -43.2 ;
      RECT 124.75 -44.01 124.85 -43.2 ;
      RECT 123.55 -44.01 123.65 -43.2 ;
      RECT 122.35 -44.01 122.45 -43.2 ;
      RECT 121.15 -44.01 121.25 -43.2 ;
      RECT 119.95 -44.01 120.05 -43.2 ;
      RECT 118.75 -44.01 118.85 -43.2 ;
      RECT 117.55 -44.01 117.65 -43.2 ;
      RECT 116.35 -44.01 116.45 -43.2 ;
      RECT 115.15 -44.01 115.25 -43.2 ;
      RECT 113.95 -44.01 114.05 -43.2 ;
      RECT 112.75 -44.01 112.85 -43.2 ;
      RECT 111.55 -44.01 111.65 -43.2 ;
      RECT 110.35 -44.01 110.45 -43.2 ;
      RECT 109.15 -44.01 109.25 -43.2 ;
      RECT 107.95 -44.01 108.05 -43.2 ;
      RECT 106.75 -44.01 106.85 -43.2 ;
      RECT 105.55 -44.01 105.65 -43.2 ;
      RECT 104.35 -44.01 104.45 -43.2 ;
      RECT 103.15 -44.01 103.25 -43.2 ;
      RECT 101.95 -44.01 102.05 -43.2 ;
      RECT 100.75 -44.01 100.85 -43.2 ;
      RECT 99.55 -44.01 99.65 -43.2 ;
      RECT 98.35 -44.01 98.45 -43.2 ;
      RECT 97.15 -44.01 97.25 -43.2 ;
      RECT 95.95 -44.01 96.05 -43.2 ;
      RECT 94.75 -44.01 94.85 -43.2 ;
      RECT 93.55 -44.01 93.65 -43.2 ;
      RECT 92.35 -44.01 92.45 -43.2 ;
      RECT 91.15 -44.01 91.25 -43.2 ;
      RECT 89.95 -44.01 90.05 -43.2 ;
      RECT 88.75 -44.01 88.85 -43.2 ;
      RECT 87.55 -44.01 87.65 -43.2 ;
      RECT 86.35 -44.01 86.45 -43.2 ;
      RECT 85.15 -44.01 85.25 -43.2 ;
      RECT 83.95 -44.01 84.05 -43.2 ;
      RECT 82.75 -44.01 82.85 -43.2 ;
      RECT 81.55 -44.01 81.65 -43.2 ;
      RECT 80.35 -44.01 80.45 -43.2 ;
      RECT 79.15 -44.01 79.25 -43.2 ;
      RECT 77.95 -44.01 78.05 -43.2 ;
      RECT 76.75 -44.01 76.85 -43.2 ;
      RECT 75.55 -44.01 75.65 -43.2 ;
      RECT 74.35 -44.01 74.45 -43.2 ;
      RECT 73.15 -44.01 73.25 -43.2 ;
      RECT 71.95 -44.01 72.05 -43.2 ;
      RECT 70.75 -44.01 70.85 -43.2 ;
      RECT 69.55 -44.01 69.65 -43.2 ;
      RECT 68.35 -44.01 68.45 -43.2 ;
      RECT 67.15 -44.01 67.25 -43.2 ;
      RECT 65.95 -44.01 66.05 -43.2 ;
      RECT 64.75 -44.01 64.85 -43.2 ;
      RECT 63.55 -44.01 63.65 -43.2 ;
      RECT 62.35 -44.01 62.45 -43.2 ;
      RECT 61.15 -44.01 61.25 -43.2 ;
      RECT 59.95 -44.01 60.05 -43.2 ;
      RECT 58.75 -44.01 58.85 -43.2 ;
      RECT 57.55 -44.01 57.65 -43.2 ;
      RECT 56.35 -44.01 56.45 -43.2 ;
      RECT 55.15 -44.01 55.25 -43.2 ;
      RECT 53.95 -44.01 54.05 -43.2 ;
      RECT 52.75 -44.01 52.85 -43.2 ;
      RECT 51.55 -44.01 51.65 -43.2 ;
      RECT 50.35 -44.01 50.45 -43.2 ;
      RECT 49.15 -44.01 49.25 -43.2 ;
      RECT 47.95 -44.01 48.05 -43.2 ;
      RECT 46.75 -44.01 46.85 -43.2 ;
      RECT 45.55 -44.01 45.65 -43.2 ;
      RECT 44.35 -44.01 44.45 -43.2 ;
      RECT 43.15 -44.01 43.25 -43.2 ;
      RECT 41.95 -44.01 42.05 -43.2 ;
      RECT 40.75 -44.01 40.85 -43.2 ;
      RECT 39.55 -44.01 39.65 -43.2 ;
      RECT 38.35 -44.01 38.45 -43.2 ;
      RECT 37.15 -44.01 37.25 -43.2 ;
      RECT 35.95 -44.01 36.05 -43.2 ;
      RECT 34.75 -44.01 34.85 -43.2 ;
      RECT 33.55 -44.01 33.65 -43.2 ;
      RECT 32.35 -44.01 32.45 -43.2 ;
      RECT 31.15 -44.01 31.25 -43.2 ;
      RECT 29.95 -44.01 30.05 -43.2 ;
      RECT 28.75 -44.01 28.85 -43.2 ;
      RECT 27.55 -44.01 27.65 -43.2 ;
      RECT 26.35 -44.01 26.45 -43.2 ;
      RECT 25.15 -44.01 25.25 -43.2 ;
      RECT 23.95 -44.01 24.05 -43.2 ;
      RECT 22.75 -44.01 22.85 -43.2 ;
      RECT 21.55 -44.01 21.65 -43.2 ;
      RECT 20.35 -44.01 20.45 -43.2 ;
      RECT 19.15 -44.01 19.25 -43.2 ;
      RECT 17.95 -44.01 18.05 -43.2 ;
      RECT 16.75 -44.01 16.85 -43.2 ;
      RECT 15.55 -44.01 15.65 -43.2 ;
      RECT 14.35 -44.01 14.45 -43.2 ;
      RECT 13.15 -44.01 13.25 -43.2 ;
      RECT 11.95 -44.01 12.05 -43.2 ;
      RECT 10.75 -44.01 10.85 -43.2 ;
      RECT 9.55 -44.01 9.65 -43.2 ;
      RECT 8.35 -44.01 8.45 -43.2 ;
      RECT 7.15 -44.01 7.25 -43.2 ;
      RECT 5.95 -44.01 6.05 -43.2 ;
      RECT 4.75 -44.01 4.85 -43.2 ;
      RECT 3.55 -44.01 3.65 -43.2 ;
      RECT 2.35 -44.01 2.45 -43.2 ;
      RECT 1.15 -44.01 1.25 -43.2 ;
      RECT -0.05 -44.01 0.05 -43.2 ;
      RECT -0.105 -43.665 156.465 -43.545 ;
      RECT 153.55 -40.78 153.65 -39.97 ;
      RECT 152.35 -40.78 152.45 -39.97 ;
      RECT 151.15 -40.78 151.25 -39.97 ;
      RECT 149.95 -40.78 150.05 -39.97 ;
      RECT 148.75 -40.78 148.85 -39.97 ;
      RECT 147.55 -40.78 147.65 -39.97 ;
      RECT 146.35 -40.78 146.45 -39.97 ;
      RECT 145.15 -40.78 145.25 -39.97 ;
      RECT 143.95 -40.78 144.05 -39.97 ;
      RECT 142.75 -40.78 142.85 -39.97 ;
      RECT 141.55 -40.78 141.65 -39.97 ;
      RECT 140.35 -40.78 140.45 -39.97 ;
      RECT 139.15 -40.78 139.25 -39.97 ;
      RECT 137.95 -40.78 138.05 -39.97 ;
      RECT 136.75 -40.78 136.85 -39.97 ;
      RECT 135.55 -40.78 135.65 -39.97 ;
      RECT 134.35 -40.78 134.45 -39.97 ;
      RECT 133.15 -40.78 133.25 -39.97 ;
      RECT 131.95 -40.78 132.05 -39.97 ;
      RECT 130.75 -40.78 130.85 -39.97 ;
      RECT 129.55 -40.78 129.65 -39.97 ;
      RECT 128.35 -40.78 128.45 -39.97 ;
      RECT 127.15 -40.78 127.25 -39.97 ;
      RECT 125.95 -40.78 126.05 -39.97 ;
      RECT 124.75 -40.78 124.85 -39.97 ;
      RECT 123.55 -40.78 123.65 -39.97 ;
      RECT 122.35 -40.78 122.45 -39.97 ;
      RECT 121.15 -40.78 121.25 -39.97 ;
      RECT 119.95 -40.78 120.05 -39.97 ;
      RECT 118.75 -40.78 118.85 -39.97 ;
      RECT 117.55 -40.78 117.65 -39.97 ;
      RECT 116.35 -40.78 116.45 -39.97 ;
      RECT 115.15 -40.78 115.25 -39.97 ;
      RECT 113.95 -40.78 114.05 -39.97 ;
      RECT 112.75 -40.78 112.85 -39.97 ;
      RECT 111.55 -40.78 111.65 -39.97 ;
      RECT 110.35 -40.78 110.45 -39.97 ;
      RECT 109.15 -40.78 109.25 -39.97 ;
      RECT 107.95 -40.78 108.05 -39.97 ;
      RECT 106.75 -40.78 106.85 -39.97 ;
      RECT 105.55 -40.78 105.65 -39.97 ;
      RECT 104.35 -40.78 104.45 -39.97 ;
      RECT 103.15 -40.78 103.25 -39.97 ;
      RECT 101.95 -40.78 102.05 -39.97 ;
      RECT 100.75 -40.78 100.85 -39.97 ;
      RECT 99.55 -40.78 99.65 -39.97 ;
      RECT 98.35 -40.78 98.45 -39.97 ;
      RECT 97.15 -40.78 97.25 -39.97 ;
      RECT 95.95 -40.78 96.05 -39.97 ;
      RECT 94.75 -40.78 94.85 -39.97 ;
      RECT 93.55 -40.78 93.65 -39.97 ;
      RECT 92.35 -40.78 92.45 -39.97 ;
      RECT 91.15 -40.78 91.25 -39.97 ;
      RECT 89.95 -40.78 90.05 -39.97 ;
      RECT 88.75 -40.78 88.85 -39.97 ;
      RECT 87.55 -40.78 87.65 -39.97 ;
      RECT 86.35 -40.78 86.45 -39.97 ;
      RECT 85.15 -40.78 85.25 -39.97 ;
      RECT 83.95 -40.78 84.05 -39.97 ;
      RECT 82.75 -40.78 82.85 -39.97 ;
      RECT 81.55 -40.78 81.65 -39.97 ;
      RECT 80.35 -40.78 80.45 -39.97 ;
      RECT 79.15 -40.78 79.25 -39.97 ;
      RECT 77.95 -40.78 78.05 -39.97 ;
      RECT 76.75 -40.78 76.85 -39.97 ;
      RECT 75.55 -40.78 75.65 -39.97 ;
      RECT 74.35 -40.78 74.45 -39.97 ;
      RECT 73.15 -40.78 73.25 -39.97 ;
      RECT 71.95 -40.78 72.05 -39.97 ;
      RECT 70.75 -40.78 70.85 -39.97 ;
      RECT 69.55 -40.78 69.65 -39.97 ;
      RECT 68.35 -40.78 68.45 -39.97 ;
      RECT 67.15 -40.78 67.25 -39.97 ;
      RECT 65.95 -40.78 66.05 -39.97 ;
      RECT 64.75 -40.78 64.85 -39.97 ;
      RECT 63.55 -40.78 63.65 -39.97 ;
      RECT 62.35 -40.78 62.45 -39.97 ;
      RECT 61.15 -40.78 61.25 -39.97 ;
      RECT 59.95 -40.78 60.05 -39.97 ;
      RECT 58.75 -40.78 58.85 -39.97 ;
      RECT 57.55 -40.78 57.65 -39.97 ;
      RECT 56.35 -40.78 56.45 -39.97 ;
      RECT 55.15 -40.78 55.25 -39.97 ;
      RECT 53.95 -40.78 54.05 -39.97 ;
      RECT 52.75 -40.78 52.85 -39.97 ;
      RECT 51.55 -40.78 51.65 -39.97 ;
      RECT 50.35 -40.78 50.45 -39.97 ;
      RECT 49.15 -40.78 49.25 -39.97 ;
      RECT 47.95 -40.78 48.05 -39.97 ;
      RECT 46.75 -40.78 46.85 -39.97 ;
      RECT 45.55 -40.78 45.65 -39.97 ;
      RECT 44.35 -40.78 44.45 -39.97 ;
      RECT 43.15 -40.78 43.25 -39.97 ;
      RECT 41.95 -40.78 42.05 -39.97 ;
      RECT 40.75 -40.78 40.85 -39.97 ;
      RECT 39.55 -40.78 39.65 -39.97 ;
      RECT 38.35 -40.78 38.45 -39.97 ;
      RECT 37.15 -40.78 37.25 -39.97 ;
      RECT 35.95 -40.78 36.05 -39.97 ;
      RECT 34.75 -40.78 34.85 -39.97 ;
      RECT 33.55 -40.78 33.65 -39.97 ;
      RECT 32.35 -40.78 32.45 -39.97 ;
      RECT 31.15 -40.78 31.25 -39.97 ;
      RECT 29.95 -40.78 30.05 -39.97 ;
      RECT 28.75 -40.78 28.85 -39.97 ;
      RECT 27.55 -40.78 27.65 -39.97 ;
      RECT 26.35 -40.78 26.45 -39.97 ;
      RECT 25.15 -40.78 25.25 -39.97 ;
      RECT 23.95 -40.78 24.05 -39.97 ;
      RECT 22.75 -40.78 22.85 -39.97 ;
      RECT 21.55 -40.78 21.65 -39.97 ;
      RECT 20.35 -40.78 20.45 -39.97 ;
      RECT 19.15 -40.78 19.25 -39.97 ;
      RECT 17.95 -40.78 18.05 -39.97 ;
      RECT 16.75 -40.78 16.85 -39.97 ;
      RECT 15.55 -40.78 15.65 -39.97 ;
      RECT 14.35 -40.78 14.45 -39.97 ;
      RECT 13.15 -40.78 13.25 -39.97 ;
      RECT 11.95 -40.78 12.05 -39.97 ;
      RECT 10.75 -40.78 10.85 -39.97 ;
      RECT 9.55 -40.78 9.65 -39.97 ;
      RECT 8.35 -40.78 8.45 -39.97 ;
      RECT 7.15 -40.78 7.25 -39.97 ;
      RECT 5.95 -40.78 6.05 -39.97 ;
      RECT 4.75 -40.78 4.85 -39.97 ;
      RECT 3.55 -40.78 3.65 -39.97 ;
      RECT 2.35 -40.78 2.45 -39.97 ;
      RECT 1.15 -40.78 1.25 -39.97 ;
      RECT -0.05 -40.78 0.05 -39.97 ;
      RECT -0.105 -40.435 156.465 -40.315 ;
      RECT 153.55 -37.55 153.65 -36.74 ;
      RECT 152.35 -37.55 152.45 -36.74 ;
      RECT 151.15 -37.55 151.25 -36.74 ;
      RECT 149.95 -37.55 150.05 -36.74 ;
      RECT 148.75 -37.55 148.85 -36.74 ;
      RECT 147.55 -37.55 147.65 -36.74 ;
      RECT 146.35 -37.55 146.45 -36.74 ;
      RECT 145.15 -37.55 145.25 -36.74 ;
      RECT 143.95 -37.55 144.05 -36.74 ;
      RECT 142.75 -37.55 142.85 -36.74 ;
      RECT 141.55 -37.55 141.65 -36.74 ;
      RECT 140.35 -37.55 140.45 -36.74 ;
      RECT 139.15 -37.55 139.25 -36.74 ;
      RECT 137.95 -37.55 138.05 -36.74 ;
      RECT 136.75 -37.55 136.85 -36.74 ;
      RECT 135.55 -37.55 135.65 -36.74 ;
      RECT 134.35 -37.55 134.45 -36.74 ;
      RECT 133.15 -37.55 133.25 -36.74 ;
      RECT 131.95 -37.55 132.05 -36.74 ;
      RECT 130.75 -37.55 130.85 -36.74 ;
      RECT 129.55 -37.55 129.65 -36.74 ;
      RECT 128.35 -37.55 128.45 -36.74 ;
      RECT 127.15 -37.55 127.25 -36.74 ;
      RECT 125.95 -37.55 126.05 -36.74 ;
      RECT 124.75 -37.55 124.85 -36.74 ;
      RECT 123.55 -37.55 123.65 -36.74 ;
      RECT 122.35 -37.55 122.45 -36.74 ;
      RECT 121.15 -37.55 121.25 -36.74 ;
      RECT 119.95 -37.55 120.05 -36.74 ;
      RECT 118.75 -37.55 118.85 -36.74 ;
      RECT 117.55 -37.55 117.65 -36.74 ;
      RECT 116.35 -37.55 116.45 -36.74 ;
      RECT 115.15 -37.55 115.25 -36.74 ;
      RECT 113.95 -37.55 114.05 -36.74 ;
      RECT 112.75 -37.55 112.85 -36.74 ;
      RECT 111.55 -37.55 111.65 -36.74 ;
      RECT 110.35 -37.55 110.45 -36.74 ;
      RECT 109.15 -37.55 109.25 -36.74 ;
      RECT 107.95 -37.55 108.05 -36.74 ;
      RECT 106.75 -37.55 106.85 -36.74 ;
      RECT 105.55 -37.55 105.65 -36.74 ;
      RECT 104.35 -37.55 104.45 -36.74 ;
      RECT 103.15 -37.55 103.25 -36.74 ;
      RECT 101.95 -37.55 102.05 -36.74 ;
      RECT 100.75 -37.55 100.85 -36.74 ;
      RECT 99.55 -37.55 99.65 -36.74 ;
      RECT 98.35 -37.55 98.45 -36.74 ;
      RECT 97.15 -37.55 97.25 -36.74 ;
      RECT 95.95 -37.55 96.05 -36.74 ;
      RECT 94.75 -37.55 94.85 -36.74 ;
      RECT 93.55 -37.55 93.65 -36.74 ;
      RECT 92.35 -37.55 92.45 -36.74 ;
      RECT 91.15 -37.55 91.25 -36.74 ;
      RECT 89.95 -37.55 90.05 -36.74 ;
      RECT 88.75 -37.55 88.85 -36.74 ;
      RECT 87.55 -37.55 87.65 -36.74 ;
      RECT 86.35 -37.55 86.45 -36.74 ;
      RECT 85.15 -37.55 85.25 -36.74 ;
      RECT 83.95 -37.55 84.05 -36.74 ;
      RECT 82.75 -37.55 82.85 -36.74 ;
      RECT 81.55 -37.55 81.65 -36.74 ;
      RECT 80.35 -37.55 80.45 -36.74 ;
      RECT 79.15 -37.55 79.25 -36.74 ;
      RECT 77.95 -37.55 78.05 -36.74 ;
      RECT 76.75 -37.55 76.85 -36.74 ;
      RECT 75.55 -37.55 75.65 -36.74 ;
      RECT 74.35 -37.55 74.45 -36.74 ;
      RECT 73.15 -37.55 73.25 -36.74 ;
      RECT 71.95 -37.55 72.05 -36.74 ;
      RECT 70.75 -37.55 70.85 -36.74 ;
      RECT 69.55 -37.55 69.65 -36.74 ;
      RECT 68.35 -37.55 68.45 -36.74 ;
      RECT 67.15 -37.55 67.25 -36.74 ;
      RECT 65.95 -37.55 66.05 -36.74 ;
      RECT 64.75 -37.55 64.85 -36.74 ;
      RECT 63.55 -37.55 63.65 -36.74 ;
      RECT 62.35 -37.55 62.45 -36.74 ;
      RECT 61.15 -37.55 61.25 -36.74 ;
      RECT 59.95 -37.55 60.05 -36.74 ;
      RECT 58.75 -37.55 58.85 -36.74 ;
      RECT 57.55 -37.55 57.65 -36.74 ;
      RECT 56.35 -37.55 56.45 -36.74 ;
      RECT 55.15 -37.55 55.25 -36.74 ;
      RECT 53.95 -37.55 54.05 -36.74 ;
      RECT 52.75 -37.55 52.85 -36.74 ;
      RECT 51.55 -37.55 51.65 -36.74 ;
      RECT 50.35 -37.55 50.45 -36.74 ;
      RECT 49.15 -37.55 49.25 -36.74 ;
      RECT 47.95 -37.55 48.05 -36.74 ;
      RECT 46.75 -37.55 46.85 -36.74 ;
      RECT 45.55 -37.55 45.65 -36.74 ;
      RECT 44.35 -37.55 44.45 -36.74 ;
      RECT 43.15 -37.55 43.25 -36.74 ;
      RECT 41.95 -37.55 42.05 -36.74 ;
      RECT 40.75 -37.55 40.85 -36.74 ;
      RECT 39.55 -37.55 39.65 -36.74 ;
      RECT 38.35 -37.55 38.45 -36.74 ;
      RECT 37.15 -37.55 37.25 -36.74 ;
      RECT 35.95 -37.55 36.05 -36.74 ;
      RECT 34.75 -37.55 34.85 -36.74 ;
      RECT 33.55 -37.55 33.65 -36.74 ;
      RECT 32.35 -37.55 32.45 -36.74 ;
      RECT 31.15 -37.55 31.25 -36.74 ;
      RECT 29.95 -37.55 30.05 -36.74 ;
      RECT 28.75 -37.55 28.85 -36.74 ;
      RECT 27.55 -37.55 27.65 -36.74 ;
      RECT 26.35 -37.55 26.45 -36.74 ;
      RECT 25.15 -37.55 25.25 -36.74 ;
      RECT 23.95 -37.55 24.05 -36.74 ;
      RECT 22.75 -37.55 22.85 -36.74 ;
      RECT 21.55 -37.55 21.65 -36.74 ;
      RECT 20.35 -37.55 20.45 -36.74 ;
      RECT 19.15 -37.55 19.25 -36.74 ;
      RECT 17.95 -37.55 18.05 -36.74 ;
      RECT 16.75 -37.55 16.85 -36.74 ;
      RECT 15.55 -37.55 15.65 -36.74 ;
      RECT 14.35 -37.55 14.45 -36.74 ;
      RECT 13.15 -37.55 13.25 -36.74 ;
      RECT 11.95 -37.55 12.05 -36.74 ;
      RECT 10.75 -37.55 10.85 -36.74 ;
      RECT 9.55 -37.55 9.65 -36.74 ;
      RECT 8.35 -37.55 8.45 -36.74 ;
      RECT 7.15 -37.55 7.25 -36.74 ;
      RECT 5.95 -37.55 6.05 -36.74 ;
      RECT 4.75 -37.55 4.85 -36.74 ;
      RECT 3.55 -37.55 3.65 -36.74 ;
      RECT 2.35 -37.55 2.45 -36.74 ;
      RECT 1.15 -37.55 1.25 -36.74 ;
      RECT -0.05 -37.55 0.05 -36.74 ;
      RECT -0.105 -37.205 156.465 -37.085 ;
      RECT 153.55 -34.32 153.65 -33.51 ;
      RECT 152.35 -34.32 152.45 -33.51 ;
      RECT 151.15 -34.32 151.25 -33.51 ;
      RECT 149.95 -34.32 150.05 -33.51 ;
      RECT 148.75 -34.32 148.85 -33.51 ;
      RECT 147.55 -34.32 147.65 -33.51 ;
      RECT 146.35 -34.32 146.45 -33.51 ;
      RECT 145.15 -34.32 145.25 -33.51 ;
      RECT 143.95 -34.32 144.05 -33.51 ;
      RECT 142.75 -34.32 142.85 -33.51 ;
      RECT 141.55 -34.32 141.65 -33.51 ;
      RECT 140.35 -34.32 140.45 -33.51 ;
      RECT 139.15 -34.32 139.25 -33.51 ;
      RECT 137.95 -34.32 138.05 -33.51 ;
      RECT 136.75 -34.32 136.85 -33.51 ;
      RECT 135.55 -34.32 135.65 -33.51 ;
      RECT 134.35 -34.32 134.45 -33.51 ;
      RECT 133.15 -34.32 133.25 -33.51 ;
      RECT 131.95 -34.32 132.05 -33.51 ;
      RECT 130.75 -34.32 130.85 -33.51 ;
      RECT 129.55 -34.32 129.65 -33.51 ;
      RECT 128.35 -34.32 128.45 -33.51 ;
      RECT 127.15 -34.32 127.25 -33.51 ;
      RECT 125.95 -34.32 126.05 -33.51 ;
      RECT 124.75 -34.32 124.85 -33.51 ;
      RECT 123.55 -34.32 123.65 -33.51 ;
      RECT 122.35 -34.32 122.45 -33.51 ;
      RECT 121.15 -34.32 121.25 -33.51 ;
      RECT 119.95 -34.32 120.05 -33.51 ;
      RECT 118.75 -34.32 118.85 -33.51 ;
      RECT 117.55 -34.32 117.65 -33.51 ;
      RECT 116.35 -34.32 116.45 -33.51 ;
      RECT 115.15 -34.32 115.25 -33.51 ;
      RECT 113.95 -34.32 114.05 -33.51 ;
      RECT 112.75 -34.32 112.85 -33.51 ;
      RECT 111.55 -34.32 111.65 -33.51 ;
      RECT 110.35 -34.32 110.45 -33.51 ;
      RECT 109.15 -34.32 109.25 -33.51 ;
      RECT 107.95 -34.32 108.05 -33.51 ;
      RECT 106.75 -34.32 106.85 -33.51 ;
      RECT 105.55 -34.32 105.65 -33.51 ;
      RECT 104.35 -34.32 104.45 -33.51 ;
      RECT 103.15 -34.32 103.25 -33.51 ;
      RECT 101.95 -34.32 102.05 -33.51 ;
      RECT 100.75 -34.32 100.85 -33.51 ;
      RECT 99.55 -34.32 99.65 -33.51 ;
      RECT 98.35 -34.32 98.45 -33.51 ;
      RECT 97.15 -34.32 97.25 -33.51 ;
      RECT 95.95 -34.32 96.05 -33.51 ;
      RECT 94.75 -34.32 94.85 -33.51 ;
      RECT 93.55 -34.32 93.65 -33.51 ;
      RECT 92.35 -34.32 92.45 -33.51 ;
      RECT 91.15 -34.32 91.25 -33.51 ;
      RECT 89.95 -34.32 90.05 -33.51 ;
      RECT 88.75 -34.32 88.85 -33.51 ;
      RECT 87.55 -34.32 87.65 -33.51 ;
      RECT 86.35 -34.32 86.45 -33.51 ;
      RECT 85.15 -34.32 85.25 -33.51 ;
      RECT 83.95 -34.32 84.05 -33.51 ;
      RECT 82.75 -34.32 82.85 -33.51 ;
      RECT 81.55 -34.32 81.65 -33.51 ;
      RECT 80.35 -34.32 80.45 -33.51 ;
      RECT 79.15 -34.32 79.25 -33.51 ;
      RECT 77.95 -34.32 78.05 -33.51 ;
      RECT 76.75 -34.32 76.85 -33.51 ;
      RECT 75.55 -34.32 75.65 -33.51 ;
      RECT 74.35 -34.32 74.45 -33.51 ;
      RECT 73.15 -34.32 73.25 -33.51 ;
      RECT 71.95 -34.32 72.05 -33.51 ;
      RECT 70.75 -34.32 70.85 -33.51 ;
      RECT 69.55 -34.32 69.65 -33.51 ;
      RECT 68.35 -34.32 68.45 -33.51 ;
      RECT 67.15 -34.32 67.25 -33.51 ;
      RECT 65.95 -34.32 66.05 -33.51 ;
      RECT 64.75 -34.32 64.85 -33.51 ;
      RECT 63.55 -34.32 63.65 -33.51 ;
      RECT 62.35 -34.32 62.45 -33.51 ;
      RECT 61.15 -34.32 61.25 -33.51 ;
      RECT 59.95 -34.32 60.05 -33.51 ;
      RECT 58.75 -34.32 58.85 -33.51 ;
      RECT 57.55 -34.32 57.65 -33.51 ;
      RECT 56.35 -34.32 56.45 -33.51 ;
      RECT 55.15 -34.32 55.25 -33.51 ;
      RECT 53.95 -34.32 54.05 -33.51 ;
      RECT 52.75 -34.32 52.85 -33.51 ;
      RECT 51.55 -34.32 51.65 -33.51 ;
      RECT 50.35 -34.32 50.45 -33.51 ;
      RECT 49.15 -34.32 49.25 -33.51 ;
      RECT 47.95 -34.32 48.05 -33.51 ;
      RECT 46.75 -34.32 46.85 -33.51 ;
      RECT 45.55 -34.32 45.65 -33.51 ;
      RECT 44.35 -34.32 44.45 -33.51 ;
      RECT 43.15 -34.32 43.25 -33.51 ;
      RECT 41.95 -34.32 42.05 -33.51 ;
      RECT 40.75 -34.32 40.85 -33.51 ;
      RECT 39.55 -34.32 39.65 -33.51 ;
      RECT 38.35 -34.32 38.45 -33.51 ;
      RECT 37.15 -34.32 37.25 -33.51 ;
      RECT 35.95 -34.32 36.05 -33.51 ;
      RECT 34.75 -34.32 34.85 -33.51 ;
      RECT 33.55 -34.32 33.65 -33.51 ;
      RECT 32.35 -34.32 32.45 -33.51 ;
      RECT 31.15 -34.32 31.25 -33.51 ;
      RECT 29.95 -34.32 30.05 -33.51 ;
      RECT 28.75 -34.32 28.85 -33.51 ;
      RECT 27.55 -34.32 27.65 -33.51 ;
      RECT 26.35 -34.32 26.45 -33.51 ;
      RECT 25.15 -34.32 25.25 -33.51 ;
      RECT 23.95 -34.32 24.05 -33.51 ;
      RECT 22.75 -34.32 22.85 -33.51 ;
      RECT 21.55 -34.32 21.65 -33.51 ;
      RECT 20.35 -34.32 20.45 -33.51 ;
      RECT 19.15 -34.32 19.25 -33.51 ;
      RECT 17.95 -34.32 18.05 -33.51 ;
      RECT 16.75 -34.32 16.85 -33.51 ;
      RECT 15.55 -34.32 15.65 -33.51 ;
      RECT 14.35 -34.32 14.45 -33.51 ;
      RECT 13.15 -34.32 13.25 -33.51 ;
      RECT 11.95 -34.32 12.05 -33.51 ;
      RECT 10.75 -34.32 10.85 -33.51 ;
      RECT 9.55 -34.32 9.65 -33.51 ;
      RECT 8.35 -34.32 8.45 -33.51 ;
      RECT 7.15 -34.32 7.25 -33.51 ;
      RECT 5.95 -34.32 6.05 -33.51 ;
      RECT 4.75 -34.32 4.85 -33.51 ;
      RECT 3.55 -34.32 3.65 -33.51 ;
      RECT 2.35 -34.32 2.45 -33.51 ;
      RECT 1.15 -34.32 1.25 -33.51 ;
      RECT -0.05 -34.32 0.05 -33.51 ;
      RECT -0.105 -33.975 156.465 -33.855 ;
      RECT 153.55 -31.09 153.65 -30.28 ;
      RECT 152.35 -31.09 152.45 -30.28 ;
      RECT 151.15 -31.09 151.25 -30.28 ;
      RECT 149.95 -31.09 150.05 -30.28 ;
      RECT 148.75 -31.09 148.85 -30.28 ;
      RECT 147.55 -31.09 147.65 -30.28 ;
      RECT 146.35 -31.09 146.45 -30.28 ;
      RECT 145.15 -31.09 145.25 -30.28 ;
      RECT 143.95 -31.09 144.05 -30.28 ;
      RECT 142.75 -31.09 142.85 -30.28 ;
      RECT 141.55 -31.09 141.65 -30.28 ;
      RECT 140.35 -31.09 140.45 -30.28 ;
      RECT 139.15 -31.09 139.25 -30.28 ;
      RECT 137.95 -31.09 138.05 -30.28 ;
      RECT 136.75 -31.09 136.85 -30.28 ;
      RECT 135.55 -31.09 135.65 -30.28 ;
      RECT 134.35 -31.09 134.45 -30.28 ;
      RECT 133.15 -31.09 133.25 -30.28 ;
      RECT 131.95 -31.09 132.05 -30.28 ;
      RECT 130.75 -31.09 130.85 -30.28 ;
      RECT 129.55 -31.09 129.65 -30.28 ;
      RECT 128.35 -31.09 128.45 -30.28 ;
      RECT 127.15 -31.09 127.25 -30.28 ;
      RECT 125.95 -31.09 126.05 -30.28 ;
      RECT 124.75 -31.09 124.85 -30.28 ;
      RECT 123.55 -31.09 123.65 -30.28 ;
      RECT 122.35 -31.09 122.45 -30.28 ;
      RECT 121.15 -31.09 121.25 -30.28 ;
      RECT 119.95 -31.09 120.05 -30.28 ;
      RECT 118.75 -31.09 118.85 -30.28 ;
      RECT 117.55 -31.09 117.65 -30.28 ;
      RECT 116.35 -31.09 116.45 -30.28 ;
      RECT 115.15 -31.09 115.25 -30.28 ;
      RECT 113.95 -31.09 114.05 -30.28 ;
      RECT 112.75 -31.09 112.85 -30.28 ;
      RECT 111.55 -31.09 111.65 -30.28 ;
      RECT 110.35 -31.09 110.45 -30.28 ;
      RECT 109.15 -31.09 109.25 -30.28 ;
      RECT 107.95 -31.09 108.05 -30.28 ;
      RECT 106.75 -31.09 106.85 -30.28 ;
      RECT 105.55 -31.09 105.65 -30.28 ;
      RECT 104.35 -31.09 104.45 -30.28 ;
      RECT 103.15 -31.09 103.25 -30.28 ;
      RECT 101.95 -31.09 102.05 -30.28 ;
      RECT 100.75 -31.09 100.85 -30.28 ;
      RECT 99.55 -31.09 99.65 -30.28 ;
      RECT 98.35 -31.09 98.45 -30.28 ;
      RECT 97.15 -31.09 97.25 -30.28 ;
      RECT 95.95 -31.09 96.05 -30.28 ;
      RECT 94.75 -31.09 94.85 -30.28 ;
      RECT 93.55 -31.09 93.65 -30.28 ;
      RECT 92.35 -31.09 92.45 -30.28 ;
      RECT 91.15 -31.09 91.25 -30.28 ;
      RECT 89.95 -31.09 90.05 -30.28 ;
      RECT 88.75 -31.09 88.85 -30.28 ;
      RECT 87.55 -31.09 87.65 -30.28 ;
      RECT 86.35 -31.09 86.45 -30.28 ;
      RECT 85.15 -31.09 85.25 -30.28 ;
      RECT 83.95 -31.09 84.05 -30.28 ;
      RECT 82.75 -31.09 82.85 -30.28 ;
      RECT 81.55 -31.09 81.65 -30.28 ;
      RECT 80.35 -31.09 80.45 -30.28 ;
      RECT 79.15 -31.09 79.25 -30.28 ;
      RECT 77.95 -31.09 78.05 -30.28 ;
      RECT 76.75 -31.09 76.85 -30.28 ;
      RECT 75.55 -31.09 75.65 -30.28 ;
      RECT 74.35 -31.09 74.45 -30.28 ;
      RECT 73.15 -31.09 73.25 -30.28 ;
      RECT 71.95 -31.09 72.05 -30.28 ;
      RECT 70.75 -31.09 70.85 -30.28 ;
      RECT 69.55 -31.09 69.65 -30.28 ;
      RECT 68.35 -31.09 68.45 -30.28 ;
      RECT 67.15 -31.09 67.25 -30.28 ;
      RECT 65.95 -31.09 66.05 -30.28 ;
      RECT 64.75 -31.09 64.85 -30.28 ;
      RECT 63.55 -31.09 63.65 -30.28 ;
      RECT 62.35 -31.09 62.45 -30.28 ;
      RECT 61.15 -31.09 61.25 -30.28 ;
      RECT 59.95 -31.09 60.05 -30.28 ;
      RECT 58.75 -31.09 58.85 -30.28 ;
      RECT 57.55 -31.09 57.65 -30.28 ;
      RECT 56.35 -31.09 56.45 -30.28 ;
      RECT 55.15 -31.09 55.25 -30.28 ;
      RECT 53.95 -31.09 54.05 -30.28 ;
      RECT 52.75 -31.09 52.85 -30.28 ;
      RECT 51.55 -31.09 51.65 -30.28 ;
      RECT 50.35 -31.09 50.45 -30.28 ;
      RECT 49.15 -31.09 49.25 -30.28 ;
      RECT 47.95 -31.09 48.05 -30.28 ;
      RECT 46.75 -31.09 46.85 -30.28 ;
      RECT 45.55 -31.09 45.65 -30.28 ;
      RECT 44.35 -31.09 44.45 -30.28 ;
      RECT 43.15 -31.09 43.25 -30.28 ;
      RECT 41.95 -31.09 42.05 -30.28 ;
      RECT 40.75 -31.09 40.85 -30.28 ;
      RECT 39.55 -31.09 39.65 -30.28 ;
      RECT 38.35 -31.09 38.45 -30.28 ;
      RECT 37.15 -31.09 37.25 -30.28 ;
      RECT 35.95 -31.09 36.05 -30.28 ;
      RECT 34.75 -31.09 34.85 -30.28 ;
      RECT 33.55 -31.09 33.65 -30.28 ;
      RECT 32.35 -31.09 32.45 -30.28 ;
      RECT 31.15 -31.09 31.25 -30.28 ;
      RECT 29.95 -31.09 30.05 -30.28 ;
      RECT 28.75 -31.09 28.85 -30.28 ;
      RECT 27.55 -31.09 27.65 -30.28 ;
      RECT 26.35 -31.09 26.45 -30.28 ;
      RECT 25.15 -31.09 25.25 -30.28 ;
      RECT 23.95 -31.09 24.05 -30.28 ;
      RECT 22.75 -31.09 22.85 -30.28 ;
      RECT 21.55 -31.09 21.65 -30.28 ;
      RECT 20.35 -31.09 20.45 -30.28 ;
      RECT 19.15 -31.09 19.25 -30.28 ;
      RECT 17.95 -31.09 18.05 -30.28 ;
      RECT 16.75 -31.09 16.85 -30.28 ;
      RECT 15.55 -31.09 15.65 -30.28 ;
      RECT 14.35 -31.09 14.45 -30.28 ;
      RECT 13.15 -31.09 13.25 -30.28 ;
      RECT 11.95 -31.09 12.05 -30.28 ;
      RECT 10.75 -31.09 10.85 -30.28 ;
      RECT 9.55 -31.09 9.65 -30.28 ;
      RECT 8.35 -31.09 8.45 -30.28 ;
      RECT 7.15 -31.09 7.25 -30.28 ;
      RECT 5.95 -31.09 6.05 -30.28 ;
      RECT 4.75 -31.09 4.85 -30.28 ;
      RECT 3.55 -31.09 3.65 -30.28 ;
      RECT 2.35 -31.09 2.45 -30.28 ;
      RECT 1.15 -31.09 1.25 -30.28 ;
      RECT -0.05 -31.09 0.05 -30.28 ;
      RECT -0.105 -30.745 156.465 -30.625 ;
      RECT 153.55 -27.86 153.65 -27.05 ;
      RECT 152.35 -27.86 152.45 -27.05 ;
      RECT 151.15 -27.86 151.25 -27.05 ;
      RECT 149.95 -27.86 150.05 -27.05 ;
      RECT 148.75 -27.86 148.85 -27.05 ;
      RECT 147.55 -27.86 147.65 -27.05 ;
      RECT 146.35 -27.86 146.45 -27.05 ;
      RECT 145.15 -27.86 145.25 -27.05 ;
      RECT 143.95 -27.86 144.05 -27.05 ;
      RECT 142.75 -27.86 142.85 -27.05 ;
      RECT 141.55 -27.86 141.65 -27.05 ;
      RECT 140.35 -27.86 140.45 -27.05 ;
      RECT 139.15 -27.86 139.25 -27.05 ;
      RECT 137.95 -27.86 138.05 -27.05 ;
      RECT 136.75 -27.86 136.85 -27.05 ;
      RECT 135.55 -27.86 135.65 -27.05 ;
      RECT 134.35 -27.86 134.45 -27.05 ;
      RECT 133.15 -27.86 133.25 -27.05 ;
      RECT 131.95 -27.86 132.05 -27.05 ;
      RECT 130.75 -27.86 130.85 -27.05 ;
      RECT 129.55 -27.86 129.65 -27.05 ;
      RECT 128.35 -27.86 128.45 -27.05 ;
      RECT 127.15 -27.86 127.25 -27.05 ;
      RECT 125.95 -27.86 126.05 -27.05 ;
      RECT 124.75 -27.86 124.85 -27.05 ;
      RECT 123.55 -27.86 123.65 -27.05 ;
      RECT 122.35 -27.86 122.45 -27.05 ;
      RECT 121.15 -27.86 121.25 -27.05 ;
      RECT 119.95 -27.86 120.05 -27.05 ;
      RECT 118.75 -27.86 118.85 -27.05 ;
      RECT 117.55 -27.86 117.65 -27.05 ;
      RECT 116.35 -27.86 116.45 -27.05 ;
      RECT 115.15 -27.86 115.25 -27.05 ;
      RECT 113.95 -27.86 114.05 -27.05 ;
      RECT 112.75 -27.86 112.85 -27.05 ;
      RECT 111.55 -27.86 111.65 -27.05 ;
      RECT 110.35 -27.86 110.45 -27.05 ;
      RECT 109.15 -27.86 109.25 -27.05 ;
      RECT 107.95 -27.86 108.05 -27.05 ;
      RECT 106.75 -27.86 106.85 -27.05 ;
      RECT 105.55 -27.86 105.65 -27.05 ;
      RECT 104.35 -27.86 104.45 -27.05 ;
      RECT 103.15 -27.86 103.25 -27.05 ;
      RECT 101.95 -27.86 102.05 -27.05 ;
      RECT 100.75 -27.86 100.85 -27.05 ;
      RECT 99.55 -27.86 99.65 -27.05 ;
      RECT 98.35 -27.86 98.45 -27.05 ;
      RECT 97.15 -27.86 97.25 -27.05 ;
      RECT 95.95 -27.86 96.05 -27.05 ;
      RECT 94.75 -27.86 94.85 -27.05 ;
      RECT 93.55 -27.86 93.65 -27.05 ;
      RECT 92.35 -27.86 92.45 -27.05 ;
      RECT 91.15 -27.86 91.25 -27.05 ;
      RECT 89.95 -27.86 90.05 -27.05 ;
      RECT 88.75 -27.86 88.85 -27.05 ;
      RECT 87.55 -27.86 87.65 -27.05 ;
      RECT 86.35 -27.86 86.45 -27.05 ;
      RECT 85.15 -27.86 85.25 -27.05 ;
      RECT 83.95 -27.86 84.05 -27.05 ;
      RECT 82.75 -27.86 82.85 -27.05 ;
      RECT 81.55 -27.86 81.65 -27.05 ;
      RECT 80.35 -27.86 80.45 -27.05 ;
      RECT 79.15 -27.86 79.25 -27.05 ;
      RECT 77.95 -27.86 78.05 -27.05 ;
      RECT 76.75 -27.86 76.85 -27.05 ;
      RECT 75.55 -27.86 75.65 -27.05 ;
      RECT 74.35 -27.86 74.45 -27.05 ;
      RECT 73.15 -27.86 73.25 -27.05 ;
      RECT 71.95 -27.86 72.05 -27.05 ;
      RECT 70.75 -27.86 70.85 -27.05 ;
      RECT 69.55 -27.86 69.65 -27.05 ;
      RECT 68.35 -27.86 68.45 -27.05 ;
      RECT 67.15 -27.86 67.25 -27.05 ;
      RECT 65.95 -27.86 66.05 -27.05 ;
      RECT 64.75 -27.86 64.85 -27.05 ;
      RECT 63.55 -27.86 63.65 -27.05 ;
      RECT 62.35 -27.86 62.45 -27.05 ;
      RECT 61.15 -27.86 61.25 -27.05 ;
      RECT 59.95 -27.86 60.05 -27.05 ;
      RECT 58.75 -27.86 58.85 -27.05 ;
      RECT 57.55 -27.86 57.65 -27.05 ;
      RECT 56.35 -27.86 56.45 -27.05 ;
      RECT 55.15 -27.86 55.25 -27.05 ;
      RECT 53.95 -27.86 54.05 -27.05 ;
      RECT 52.75 -27.86 52.85 -27.05 ;
      RECT 51.55 -27.86 51.65 -27.05 ;
      RECT 50.35 -27.86 50.45 -27.05 ;
      RECT 49.15 -27.86 49.25 -27.05 ;
      RECT 47.95 -27.86 48.05 -27.05 ;
      RECT 46.75 -27.86 46.85 -27.05 ;
      RECT 45.55 -27.86 45.65 -27.05 ;
      RECT 44.35 -27.86 44.45 -27.05 ;
      RECT 43.15 -27.86 43.25 -27.05 ;
      RECT 41.95 -27.86 42.05 -27.05 ;
      RECT 40.75 -27.86 40.85 -27.05 ;
      RECT 39.55 -27.86 39.65 -27.05 ;
      RECT 38.35 -27.86 38.45 -27.05 ;
      RECT 37.15 -27.86 37.25 -27.05 ;
      RECT 35.95 -27.86 36.05 -27.05 ;
      RECT 34.75 -27.86 34.85 -27.05 ;
      RECT 33.55 -27.86 33.65 -27.05 ;
      RECT 32.35 -27.86 32.45 -27.05 ;
      RECT 31.15 -27.86 31.25 -27.05 ;
      RECT 29.95 -27.86 30.05 -27.05 ;
      RECT 28.75 -27.86 28.85 -27.05 ;
      RECT 27.55 -27.86 27.65 -27.05 ;
      RECT 26.35 -27.86 26.45 -27.05 ;
      RECT 25.15 -27.86 25.25 -27.05 ;
      RECT 23.95 -27.86 24.05 -27.05 ;
      RECT 22.75 -27.86 22.85 -27.05 ;
      RECT 21.55 -27.86 21.65 -27.05 ;
      RECT 20.35 -27.86 20.45 -27.05 ;
      RECT 19.15 -27.86 19.25 -27.05 ;
      RECT 17.95 -27.86 18.05 -27.05 ;
      RECT 16.75 -27.86 16.85 -27.05 ;
      RECT 15.55 -27.86 15.65 -27.05 ;
      RECT 14.35 -27.86 14.45 -27.05 ;
      RECT 13.15 -27.86 13.25 -27.05 ;
      RECT 11.95 -27.86 12.05 -27.05 ;
      RECT 10.75 -27.86 10.85 -27.05 ;
      RECT 9.55 -27.86 9.65 -27.05 ;
      RECT 8.35 -27.86 8.45 -27.05 ;
      RECT 7.15 -27.86 7.25 -27.05 ;
      RECT 5.95 -27.86 6.05 -27.05 ;
      RECT 4.75 -27.86 4.85 -27.05 ;
      RECT 3.55 -27.86 3.65 -27.05 ;
      RECT 2.35 -27.86 2.45 -27.05 ;
      RECT 1.15 -27.86 1.25 -27.05 ;
      RECT -0.05 -27.86 0.05 -27.05 ;
      RECT -0.105 -27.515 156.465 -27.395 ;
      RECT 153.55 -24.63 153.65 -23.82 ;
      RECT 152.35 -24.63 152.45 -23.82 ;
      RECT 151.15 -24.63 151.25 -23.82 ;
      RECT 149.95 -24.63 150.05 -23.82 ;
      RECT 148.75 -24.63 148.85 -23.82 ;
      RECT 147.55 -24.63 147.65 -23.82 ;
      RECT 146.35 -24.63 146.45 -23.82 ;
      RECT 145.15 -24.63 145.25 -23.82 ;
      RECT 143.95 -24.63 144.05 -23.82 ;
      RECT 142.75 -24.63 142.85 -23.82 ;
      RECT 141.55 -24.63 141.65 -23.82 ;
      RECT 140.35 -24.63 140.45 -23.82 ;
      RECT 139.15 -24.63 139.25 -23.82 ;
      RECT 137.95 -24.63 138.05 -23.82 ;
      RECT 136.75 -24.63 136.85 -23.82 ;
      RECT 135.55 -24.63 135.65 -23.82 ;
      RECT 134.35 -24.63 134.45 -23.82 ;
      RECT 133.15 -24.63 133.25 -23.82 ;
      RECT 131.95 -24.63 132.05 -23.82 ;
      RECT 130.75 -24.63 130.85 -23.82 ;
      RECT 129.55 -24.63 129.65 -23.82 ;
      RECT 128.35 -24.63 128.45 -23.82 ;
      RECT 127.15 -24.63 127.25 -23.82 ;
      RECT 125.95 -24.63 126.05 -23.82 ;
      RECT 124.75 -24.63 124.85 -23.82 ;
      RECT 123.55 -24.63 123.65 -23.82 ;
      RECT 122.35 -24.63 122.45 -23.82 ;
      RECT 121.15 -24.63 121.25 -23.82 ;
      RECT 119.95 -24.63 120.05 -23.82 ;
      RECT 118.75 -24.63 118.85 -23.82 ;
      RECT 117.55 -24.63 117.65 -23.82 ;
      RECT 116.35 -24.63 116.45 -23.82 ;
      RECT 115.15 -24.63 115.25 -23.82 ;
      RECT 113.95 -24.63 114.05 -23.82 ;
      RECT 112.75 -24.63 112.85 -23.82 ;
      RECT 111.55 -24.63 111.65 -23.82 ;
      RECT 110.35 -24.63 110.45 -23.82 ;
      RECT 109.15 -24.63 109.25 -23.82 ;
      RECT 107.95 -24.63 108.05 -23.82 ;
      RECT 106.75 -24.63 106.85 -23.82 ;
      RECT 105.55 -24.63 105.65 -23.82 ;
      RECT 104.35 -24.63 104.45 -23.82 ;
      RECT 103.15 -24.63 103.25 -23.82 ;
      RECT 101.95 -24.63 102.05 -23.82 ;
      RECT 100.75 -24.63 100.85 -23.82 ;
      RECT 99.55 -24.63 99.65 -23.82 ;
      RECT 98.35 -24.63 98.45 -23.82 ;
      RECT 97.15 -24.63 97.25 -23.82 ;
      RECT 95.95 -24.63 96.05 -23.82 ;
      RECT 94.75 -24.63 94.85 -23.82 ;
      RECT 93.55 -24.63 93.65 -23.82 ;
      RECT 92.35 -24.63 92.45 -23.82 ;
      RECT 91.15 -24.63 91.25 -23.82 ;
      RECT 89.95 -24.63 90.05 -23.82 ;
      RECT 88.75 -24.63 88.85 -23.82 ;
      RECT 87.55 -24.63 87.65 -23.82 ;
      RECT 86.35 -24.63 86.45 -23.82 ;
      RECT 85.15 -24.63 85.25 -23.82 ;
      RECT 83.95 -24.63 84.05 -23.82 ;
      RECT 82.75 -24.63 82.85 -23.82 ;
      RECT 81.55 -24.63 81.65 -23.82 ;
      RECT 80.35 -24.63 80.45 -23.82 ;
      RECT 79.15 -24.63 79.25 -23.82 ;
      RECT 77.95 -24.63 78.05 -23.82 ;
      RECT 76.75 -24.63 76.85 -23.82 ;
      RECT 75.55 -24.63 75.65 -23.82 ;
      RECT 74.35 -24.63 74.45 -23.82 ;
      RECT 73.15 -24.63 73.25 -23.82 ;
      RECT 71.95 -24.63 72.05 -23.82 ;
      RECT 70.75 -24.63 70.85 -23.82 ;
      RECT 69.55 -24.63 69.65 -23.82 ;
      RECT 68.35 -24.63 68.45 -23.82 ;
      RECT 67.15 -24.63 67.25 -23.82 ;
      RECT 65.95 -24.63 66.05 -23.82 ;
      RECT 64.75 -24.63 64.85 -23.82 ;
      RECT 63.55 -24.63 63.65 -23.82 ;
      RECT 62.35 -24.63 62.45 -23.82 ;
      RECT 61.15 -24.63 61.25 -23.82 ;
      RECT 59.95 -24.63 60.05 -23.82 ;
      RECT 58.75 -24.63 58.85 -23.82 ;
      RECT 57.55 -24.63 57.65 -23.82 ;
      RECT 56.35 -24.63 56.45 -23.82 ;
      RECT 55.15 -24.63 55.25 -23.82 ;
      RECT 53.95 -24.63 54.05 -23.82 ;
      RECT 52.75 -24.63 52.85 -23.82 ;
      RECT 51.55 -24.63 51.65 -23.82 ;
      RECT 50.35 -24.63 50.45 -23.82 ;
      RECT 49.15 -24.63 49.25 -23.82 ;
      RECT 47.95 -24.63 48.05 -23.82 ;
      RECT 46.75 -24.63 46.85 -23.82 ;
      RECT 45.55 -24.63 45.65 -23.82 ;
      RECT 44.35 -24.63 44.45 -23.82 ;
      RECT 43.15 -24.63 43.25 -23.82 ;
      RECT 41.95 -24.63 42.05 -23.82 ;
      RECT 40.75 -24.63 40.85 -23.82 ;
      RECT 39.55 -24.63 39.65 -23.82 ;
      RECT 38.35 -24.63 38.45 -23.82 ;
      RECT 37.15 -24.63 37.25 -23.82 ;
      RECT 35.95 -24.63 36.05 -23.82 ;
      RECT 34.75 -24.63 34.85 -23.82 ;
      RECT 33.55 -24.63 33.65 -23.82 ;
      RECT 32.35 -24.63 32.45 -23.82 ;
      RECT 31.15 -24.63 31.25 -23.82 ;
      RECT 29.95 -24.63 30.05 -23.82 ;
      RECT 28.75 -24.63 28.85 -23.82 ;
      RECT 27.55 -24.63 27.65 -23.82 ;
      RECT 26.35 -24.63 26.45 -23.82 ;
      RECT 25.15 -24.63 25.25 -23.82 ;
      RECT 23.95 -24.63 24.05 -23.82 ;
      RECT 22.75 -24.63 22.85 -23.82 ;
      RECT 21.55 -24.63 21.65 -23.82 ;
      RECT 20.35 -24.63 20.45 -23.82 ;
      RECT 19.15 -24.63 19.25 -23.82 ;
      RECT 17.95 -24.63 18.05 -23.82 ;
      RECT 16.75 -24.63 16.85 -23.82 ;
      RECT 15.55 -24.63 15.65 -23.82 ;
      RECT 14.35 -24.63 14.45 -23.82 ;
      RECT 13.15 -24.63 13.25 -23.82 ;
      RECT 11.95 -24.63 12.05 -23.82 ;
      RECT 10.75 -24.63 10.85 -23.82 ;
      RECT 9.55 -24.63 9.65 -23.82 ;
      RECT 8.35 -24.63 8.45 -23.82 ;
      RECT 7.15 -24.63 7.25 -23.82 ;
      RECT 5.95 -24.63 6.05 -23.82 ;
      RECT 4.75 -24.63 4.85 -23.82 ;
      RECT 3.55 -24.63 3.65 -23.82 ;
      RECT 2.35 -24.63 2.45 -23.82 ;
      RECT 1.15 -24.63 1.25 -23.82 ;
      RECT -0.05 -24.63 0.05 -23.82 ;
      RECT -0.105 -24.285 156.465 -24.165 ;
      RECT 153.55 -21.4 153.65 -20.59 ;
      RECT 152.35 -21.4 152.45 -20.59 ;
      RECT 151.15 -21.4 151.25 -20.59 ;
      RECT 149.95 -21.4 150.05 -20.59 ;
      RECT 148.75 -21.4 148.85 -20.59 ;
      RECT 147.55 -21.4 147.65 -20.59 ;
      RECT 146.35 -21.4 146.45 -20.59 ;
      RECT 145.15 -21.4 145.25 -20.59 ;
      RECT 143.95 -21.4 144.05 -20.59 ;
      RECT 142.75 -21.4 142.85 -20.59 ;
      RECT 141.55 -21.4 141.65 -20.59 ;
      RECT 140.35 -21.4 140.45 -20.59 ;
      RECT 139.15 -21.4 139.25 -20.59 ;
      RECT 137.95 -21.4 138.05 -20.59 ;
      RECT 136.75 -21.4 136.85 -20.59 ;
      RECT 135.55 -21.4 135.65 -20.59 ;
      RECT 134.35 -21.4 134.45 -20.59 ;
      RECT 133.15 -21.4 133.25 -20.59 ;
      RECT 131.95 -21.4 132.05 -20.59 ;
      RECT 130.75 -21.4 130.85 -20.59 ;
      RECT 129.55 -21.4 129.65 -20.59 ;
      RECT 128.35 -21.4 128.45 -20.59 ;
      RECT 127.15 -21.4 127.25 -20.59 ;
      RECT 125.95 -21.4 126.05 -20.59 ;
      RECT 124.75 -21.4 124.85 -20.59 ;
      RECT 123.55 -21.4 123.65 -20.59 ;
      RECT 122.35 -21.4 122.45 -20.59 ;
      RECT 121.15 -21.4 121.25 -20.59 ;
      RECT 119.95 -21.4 120.05 -20.59 ;
      RECT 118.75 -21.4 118.85 -20.59 ;
      RECT 117.55 -21.4 117.65 -20.59 ;
      RECT 116.35 -21.4 116.45 -20.59 ;
      RECT 115.15 -21.4 115.25 -20.59 ;
      RECT 113.95 -21.4 114.05 -20.59 ;
      RECT 112.75 -21.4 112.85 -20.59 ;
      RECT 111.55 -21.4 111.65 -20.59 ;
      RECT 110.35 -21.4 110.45 -20.59 ;
      RECT 109.15 -21.4 109.25 -20.59 ;
      RECT 107.95 -21.4 108.05 -20.59 ;
      RECT 106.75 -21.4 106.85 -20.59 ;
      RECT 105.55 -21.4 105.65 -20.59 ;
      RECT 104.35 -21.4 104.45 -20.59 ;
      RECT 103.15 -21.4 103.25 -20.59 ;
      RECT 101.95 -21.4 102.05 -20.59 ;
      RECT 100.75 -21.4 100.85 -20.59 ;
      RECT 99.55 -21.4 99.65 -20.59 ;
      RECT 98.35 -21.4 98.45 -20.59 ;
      RECT 97.15 -21.4 97.25 -20.59 ;
      RECT 95.95 -21.4 96.05 -20.59 ;
      RECT 94.75 -21.4 94.85 -20.59 ;
      RECT 93.55 -21.4 93.65 -20.59 ;
      RECT 92.35 -21.4 92.45 -20.59 ;
      RECT 91.15 -21.4 91.25 -20.59 ;
      RECT 89.95 -21.4 90.05 -20.59 ;
      RECT 88.75 -21.4 88.85 -20.59 ;
      RECT 87.55 -21.4 87.65 -20.59 ;
      RECT 86.35 -21.4 86.45 -20.59 ;
      RECT 85.15 -21.4 85.25 -20.59 ;
      RECT 83.95 -21.4 84.05 -20.59 ;
      RECT 82.75 -21.4 82.85 -20.59 ;
      RECT 81.55 -21.4 81.65 -20.59 ;
      RECT 80.35 -21.4 80.45 -20.59 ;
      RECT 79.15 -21.4 79.25 -20.59 ;
      RECT 77.95 -21.4 78.05 -20.59 ;
      RECT 76.75 -21.4 76.85 -20.59 ;
      RECT 75.55 -21.4 75.65 -20.59 ;
      RECT 74.35 -21.4 74.45 -20.59 ;
      RECT 73.15 -21.4 73.25 -20.59 ;
      RECT 71.95 -21.4 72.05 -20.59 ;
      RECT 70.75 -21.4 70.85 -20.59 ;
      RECT 69.55 -21.4 69.65 -20.59 ;
      RECT 68.35 -21.4 68.45 -20.59 ;
      RECT 67.15 -21.4 67.25 -20.59 ;
      RECT 65.95 -21.4 66.05 -20.59 ;
      RECT 64.75 -21.4 64.85 -20.59 ;
      RECT 63.55 -21.4 63.65 -20.59 ;
      RECT 62.35 -21.4 62.45 -20.59 ;
      RECT 61.15 -21.4 61.25 -20.59 ;
      RECT 59.95 -21.4 60.05 -20.59 ;
      RECT 58.75 -21.4 58.85 -20.59 ;
      RECT 57.55 -21.4 57.65 -20.59 ;
      RECT 56.35 -21.4 56.45 -20.59 ;
      RECT 55.15 -21.4 55.25 -20.59 ;
      RECT 53.95 -21.4 54.05 -20.59 ;
      RECT 52.75 -21.4 52.85 -20.59 ;
      RECT 51.55 -21.4 51.65 -20.59 ;
      RECT 50.35 -21.4 50.45 -20.59 ;
      RECT 49.15 -21.4 49.25 -20.59 ;
      RECT 47.95 -21.4 48.05 -20.59 ;
      RECT 46.75 -21.4 46.85 -20.59 ;
      RECT 45.55 -21.4 45.65 -20.59 ;
      RECT 44.35 -21.4 44.45 -20.59 ;
      RECT 43.15 -21.4 43.25 -20.59 ;
      RECT 41.95 -21.4 42.05 -20.59 ;
      RECT 40.75 -21.4 40.85 -20.59 ;
      RECT 39.55 -21.4 39.65 -20.59 ;
      RECT 38.35 -21.4 38.45 -20.59 ;
      RECT 37.15 -21.4 37.25 -20.59 ;
      RECT 35.95 -21.4 36.05 -20.59 ;
      RECT 34.75 -21.4 34.85 -20.59 ;
      RECT 33.55 -21.4 33.65 -20.59 ;
      RECT 32.35 -21.4 32.45 -20.59 ;
      RECT 31.15 -21.4 31.25 -20.59 ;
      RECT 29.95 -21.4 30.05 -20.59 ;
      RECT 28.75 -21.4 28.85 -20.59 ;
      RECT 27.55 -21.4 27.65 -20.59 ;
      RECT 26.35 -21.4 26.45 -20.59 ;
      RECT 25.15 -21.4 25.25 -20.59 ;
      RECT 23.95 -21.4 24.05 -20.59 ;
      RECT 22.75 -21.4 22.85 -20.59 ;
      RECT 21.55 -21.4 21.65 -20.59 ;
      RECT 20.35 -21.4 20.45 -20.59 ;
      RECT 19.15 -21.4 19.25 -20.59 ;
      RECT 17.95 -21.4 18.05 -20.59 ;
      RECT 16.75 -21.4 16.85 -20.59 ;
      RECT 15.55 -21.4 15.65 -20.59 ;
      RECT 14.35 -21.4 14.45 -20.59 ;
      RECT 13.15 -21.4 13.25 -20.59 ;
      RECT 11.95 -21.4 12.05 -20.59 ;
      RECT 10.75 -21.4 10.85 -20.59 ;
      RECT 9.55 -21.4 9.65 -20.59 ;
      RECT 8.35 -21.4 8.45 -20.59 ;
      RECT 7.15 -21.4 7.25 -20.59 ;
      RECT 5.95 -21.4 6.05 -20.59 ;
      RECT 4.75 -21.4 4.85 -20.59 ;
      RECT 3.55 -21.4 3.65 -20.59 ;
      RECT 2.35 -21.4 2.45 -20.59 ;
      RECT 1.15 -21.4 1.25 -20.59 ;
      RECT -0.05 -21.4 0.05 -20.59 ;
      RECT -0.105 -21.055 156.465 -20.935 ;
      RECT 153.55 -18.17 153.65 -17.36 ;
      RECT 152.35 -18.17 152.45 -17.36 ;
      RECT 151.15 -18.17 151.25 -17.36 ;
      RECT 149.95 -18.17 150.05 -17.36 ;
      RECT 148.75 -18.17 148.85 -17.36 ;
      RECT 147.55 -18.17 147.65 -17.36 ;
      RECT 146.35 -18.17 146.45 -17.36 ;
      RECT 145.15 -18.17 145.25 -17.36 ;
      RECT 143.95 -18.17 144.05 -17.36 ;
      RECT 142.75 -18.17 142.85 -17.36 ;
      RECT 141.55 -18.17 141.65 -17.36 ;
      RECT 140.35 -18.17 140.45 -17.36 ;
      RECT 139.15 -18.17 139.25 -17.36 ;
      RECT 137.95 -18.17 138.05 -17.36 ;
      RECT 136.75 -18.17 136.85 -17.36 ;
      RECT 135.55 -18.17 135.65 -17.36 ;
      RECT 134.35 -18.17 134.45 -17.36 ;
      RECT 133.15 -18.17 133.25 -17.36 ;
      RECT 131.95 -18.17 132.05 -17.36 ;
      RECT 130.75 -18.17 130.85 -17.36 ;
      RECT 129.55 -18.17 129.65 -17.36 ;
      RECT 128.35 -18.17 128.45 -17.36 ;
      RECT 127.15 -18.17 127.25 -17.36 ;
      RECT 125.95 -18.17 126.05 -17.36 ;
      RECT 124.75 -18.17 124.85 -17.36 ;
      RECT 123.55 -18.17 123.65 -17.36 ;
      RECT 122.35 -18.17 122.45 -17.36 ;
      RECT 121.15 -18.17 121.25 -17.36 ;
      RECT 119.95 -18.17 120.05 -17.36 ;
      RECT 118.75 -18.17 118.85 -17.36 ;
      RECT 117.55 -18.17 117.65 -17.36 ;
      RECT 116.35 -18.17 116.45 -17.36 ;
      RECT 115.15 -18.17 115.25 -17.36 ;
      RECT 113.95 -18.17 114.05 -17.36 ;
      RECT 112.75 -18.17 112.85 -17.36 ;
      RECT 111.55 -18.17 111.65 -17.36 ;
      RECT 110.35 -18.17 110.45 -17.36 ;
      RECT 109.15 -18.17 109.25 -17.36 ;
      RECT 107.95 -18.17 108.05 -17.36 ;
      RECT 106.75 -18.17 106.85 -17.36 ;
      RECT 105.55 -18.17 105.65 -17.36 ;
      RECT 104.35 -18.17 104.45 -17.36 ;
      RECT 103.15 -18.17 103.25 -17.36 ;
      RECT 101.95 -18.17 102.05 -17.36 ;
      RECT 100.75 -18.17 100.85 -17.36 ;
      RECT 99.55 -18.17 99.65 -17.36 ;
      RECT 98.35 -18.17 98.45 -17.36 ;
      RECT 97.15 -18.17 97.25 -17.36 ;
      RECT 95.95 -18.17 96.05 -17.36 ;
      RECT 94.75 -18.17 94.85 -17.36 ;
      RECT 93.55 -18.17 93.65 -17.36 ;
      RECT 92.35 -18.17 92.45 -17.36 ;
      RECT 91.15 -18.17 91.25 -17.36 ;
      RECT 89.95 -18.17 90.05 -17.36 ;
      RECT 88.75 -18.17 88.85 -17.36 ;
      RECT 87.55 -18.17 87.65 -17.36 ;
      RECT 86.35 -18.17 86.45 -17.36 ;
      RECT 85.15 -18.17 85.25 -17.36 ;
      RECT 83.95 -18.17 84.05 -17.36 ;
      RECT 82.75 -18.17 82.85 -17.36 ;
      RECT 81.55 -18.17 81.65 -17.36 ;
      RECT 80.35 -18.17 80.45 -17.36 ;
      RECT 79.15 -18.17 79.25 -17.36 ;
      RECT 77.95 -18.17 78.05 -17.36 ;
      RECT 76.75 -18.17 76.85 -17.36 ;
      RECT 75.55 -18.17 75.65 -17.36 ;
      RECT 74.35 -18.17 74.45 -17.36 ;
      RECT 73.15 -18.17 73.25 -17.36 ;
      RECT 71.95 -18.17 72.05 -17.36 ;
      RECT 70.75 -18.17 70.85 -17.36 ;
      RECT 69.55 -18.17 69.65 -17.36 ;
      RECT 68.35 -18.17 68.45 -17.36 ;
      RECT 67.15 -18.17 67.25 -17.36 ;
      RECT 65.95 -18.17 66.05 -17.36 ;
      RECT 64.75 -18.17 64.85 -17.36 ;
      RECT 63.55 -18.17 63.65 -17.36 ;
      RECT 62.35 -18.17 62.45 -17.36 ;
      RECT 61.15 -18.17 61.25 -17.36 ;
      RECT 59.95 -18.17 60.05 -17.36 ;
      RECT 58.75 -18.17 58.85 -17.36 ;
      RECT 57.55 -18.17 57.65 -17.36 ;
      RECT 56.35 -18.17 56.45 -17.36 ;
      RECT 55.15 -18.17 55.25 -17.36 ;
      RECT 53.95 -18.17 54.05 -17.36 ;
      RECT 52.75 -18.17 52.85 -17.36 ;
      RECT 51.55 -18.17 51.65 -17.36 ;
      RECT 50.35 -18.17 50.45 -17.36 ;
      RECT 49.15 -18.17 49.25 -17.36 ;
      RECT 47.95 -18.17 48.05 -17.36 ;
      RECT 46.75 -18.17 46.85 -17.36 ;
      RECT 45.55 -18.17 45.65 -17.36 ;
      RECT 44.35 -18.17 44.45 -17.36 ;
      RECT 43.15 -18.17 43.25 -17.36 ;
      RECT 41.95 -18.17 42.05 -17.36 ;
      RECT 40.75 -18.17 40.85 -17.36 ;
      RECT 39.55 -18.17 39.65 -17.36 ;
      RECT 38.35 -18.17 38.45 -17.36 ;
      RECT 37.15 -18.17 37.25 -17.36 ;
      RECT 35.95 -18.17 36.05 -17.36 ;
      RECT 34.75 -18.17 34.85 -17.36 ;
      RECT 33.55 -18.17 33.65 -17.36 ;
      RECT 32.35 -18.17 32.45 -17.36 ;
      RECT 31.15 -18.17 31.25 -17.36 ;
      RECT 29.95 -18.17 30.05 -17.36 ;
      RECT 28.75 -18.17 28.85 -17.36 ;
      RECT 27.55 -18.17 27.65 -17.36 ;
      RECT 26.35 -18.17 26.45 -17.36 ;
      RECT 25.15 -18.17 25.25 -17.36 ;
      RECT 23.95 -18.17 24.05 -17.36 ;
      RECT 22.75 -18.17 22.85 -17.36 ;
      RECT 21.55 -18.17 21.65 -17.36 ;
      RECT 20.35 -18.17 20.45 -17.36 ;
      RECT 19.15 -18.17 19.25 -17.36 ;
      RECT 17.95 -18.17 18.05 -17.36 ;
      RECT 16.75 -18.17 16.85 -17.36 ;
      RECT 15.55 -18.17 15.65 -17.36 ;
      RECT 14.35 -18.17 14.45 -17.36 ;
      RECT 13.15 -18.17 13.25 -17.36 ;
      RECT 11.95 -18.17 12.05 -17.36 ;
      RECT 10.75 -18.17 10.85 -17.36 ;
      RECT 9.55 -18.17 9.65 -17.36 ;
      RECT 8.35 -18.17 8.45 -17.36 ;
      RECT 7.15 -18.17 7.25 -17.36 ;
      RECT 5.95 -18.17 6.05 -17.36 ;
      RECT 4.75 -18.17 4.85 -17.36 ;
      RECT 3.55 -18.17 3.65 -17.36 ;
      RECT 2.35 -18.17 2.45 -17.36 ;
      RECT 1.15 -18.17 1.25 -17.36 ;
      RECT -0.05 -18.17 0.05 -17.36 ;
      RECT -0.105 -17.825 156.465 -17.705 ;
      RECT 153.55 -14.94 153.65 -14.13 ;
      RECT 152.35 -14.94 152.45 -14.13 ;
      RECT 151.15 -14.94 151.25 -14.13 ;
      RECT 149.95 -14.94 150.05 -14.13 ;
      RECT 148.75 -14.94 148.85 -14.13 ;
      RECT 147.55 -14.94 147.65 -14.13 ;
      RECT 146.35 -14.94 146.45 -14.13 ;
      RECT 145.15 -14.94 145.25 -14.13 ;
      RECT 143.95 -14.94 144.05 -14.13 ;
      RECT 142.75 -14.94 142.85 -14.13 ;
      RECT 141.55 -14.94 141.65 -14.13 ;
      RECT 140.35 -14.94 140.45 -14.13 ;
      RECT 139.15 -14.94 139.25 -14.13 ;
      RECT 137.95 -14.94 138.05 -14.13 ;
      RECT 136.75 -14.94 136.85 -14.13 ;
      RECT 135.55 -14.94 135.65 -14.13 ;
      RECT 134.35 -14.94 134.45 -14.13 ;
      RECT 133.15 -14.94 133.25 -14.13 ;
      RECT 131.95 -14.94 132.05 -14.13 ;
      RECT 130.75 -14.94 130.85 -14.13 ;
      RECT 129.55 -14.94 129.65 -14.13 ;
      RECT 128.35 -14.94 128.45 -14.13 ;
      RECT 127.15 -14.94 127.25 -14.13 ;
      RECT 125.95 -14.94 126.05 -14.13 ;
      RECT 124.75 -14.94 124.85 -14.13 ;
      RECT 123.55 -14.94 123.65 -14.13 ;
      RECT 122.35 -14.94 122.45 -14.13 ;
      RECT 121.15 -14.94 121.25 -14.13 ;
      RECT 119.95 -14.94 120.05 -14.13 ;
      RECT 118.75 -14.94 118.85 -14.13 ;
      RECT 117.55 -14.94 117.65 -14.13 ;
      RECT 116.35 -14.94 116.45 -14.13 ;
      RECT 115.15 -14.94 115.25 -14.13 ;
      RECT 113.95 -14.94 114.05 -14.13 ;
      RECT 112.75 -14.94 112.85 -14.13 ;
      RECT 111.55 -14.94 111.65 -14.13 ;
      RECT 110.35 -14.94 110.45 -14.13 ;
      RECT 109.15 -14.94 109.25 -14.13 ;
      RECT 107.95 -14.94 108.05 -14.13 ;
      RECT 106.75 -14.94 106.85 -14.13 ;
      RECT 105.55 -14.94 105.65 -14.13 ;
      RECT 104.35 -14.94 104.45 -14.13 ;
      RECT 103.15 -14.94 103.25 -14.13 ;
      RECT 101.95 -14.94 102.05 -14.13 ;
      RECT 100.75 -14.94 100.85 -14.13 ;
      RECT 99.55 -14.94 99.65 -14.13 ;
      RECT 98.35 -14.94 98.45 -14.13 ;
      RECT 97.15 -14.94 97.25 -14.13 ;
      RECT 95.95 -14.94 96.05 -14.13 ;
      RECT 94.75 -14.94 94.85 -14.13 ;
      RECT 93.55 -14.94 93.65 -14.13 ;
      RECT 92.35 -14.94 92.45 -14.13 ;
      RECT 91.15 -14.94 91.25 -14.13 ;
      RECT 89.95 -14.94 90.05 -14.13 ;
      RECT 88.75 -14.94 88.85 -14.13 ;
      RECT 87.55 -14.94 87.65 -14.13 ;
      RECT 86.35 -14.94 86.45 -14.13 ;
      RECT 85.15 -14.94 85.25 -14.13 ;
      RECT 83.95 -14.94 84.05 -14.13 ;
      RECT 82.75 -14.94 82.85 -14.13 ;
      RECT 81.55 -14.94 81.65 -14.13 ;
      RECT 80.35 -14.94 80.45 -14.13 ;
      RECT 79.15 -14.94 79.25 -14.13 ;
      RECT 77.95 -14.94 78.05 -14.13 ;
      RECT 76.75 -14.94 76.85 -14.13 ;
      RECT 75.55 -14.94 75.65 -14.13 ;
      RECT 74.35 -14.94 74.45 -14.13 ;
      RECT 73.15 -14.94 73.25 -14.13 ;
      RECT 71.95 -14.94 72.05 -14.13 ;
      RECT 70.75 -14.94 70.85 -14.13 ;
      RECT 69.55 -14.94 69.65 -14.13 ;
      RECT 68.35 -14.94 68.45 -14.13 ;
      RECT 67.15 -14.94 67.25 -14.13 ;
      RECT 65.95 -14.94 66.05 -14.13 ;
      RECT 64.75 -14.94 64.85 -14.13 ;
      RECT 63.55 -14.94 63.65 -14.13 ;
      RECT 62.35 -14.94 62.45 -14.13 ;
      RECT 61.15 -14.94 61.25 -14.13 ;
      RECT 59.95 -14.94 60.05 -14.13 ;
      RECT 58.75 -14.94 58.85 -14.13 ;
      RECT 57.55 -14.94 57.65 -14.13 ;
      RECT 56.35 -14.94 56.45 -14.13 ;
      RECT 55.15 -14.94 55.25 -14.13 ;
      RECT 53.95 -14.94 54.05 -14.13 ;
      RECT 52.75 -14.94 52.85 -14.13 ;
      RECT 51.55 -14.94 51.65 -14.13 ;
      RECT 50.35 -14.94 50.45 -14.13 ;
      RECT 49.15 -14.94 49.25 -14.13 ;
      RECT 47.95 -14.94 48.05 -14.13 ;
      RECT 46.75 -14.94 46.85 -14.13 ;
      RECT 45.55 -14.94 45.65 -14.13 ;
      RECT 44.35 -14.94 44.45 -14.13 ;
      RECT 43.15 -14.94 43.25 -14.13 ;
      RECT 41.95 -14.94 42.05 -14.13 ;
      RECT 40.75 -14.94 40.85 -14.13 ;
      RECT 39.55 -14.94 39.65 -14.13 ;
      RECT 38.35 -14.94 38.45 -14.13 ;
      RECT 37.15 -14.94 37.25 -14.13 ;
      RECT 35.95 -14.94 36.05 -14.13 ;
      RECT 34.75 -14.94 34.85 -14.13 ;
      RECT 33.55 -14.94 33.65 -14.13 ;
      RECT 32.35 -14.94 32.45 -14.13 ;
      RECT 31.15 -14.94 31.25 -14.13 ;
      RECT 29.95 -14.94 30.05 -14.13 ;
      RECT 28.75 -14.94 28.85 -14.13 ;
      RECT 27.55 -14.94 27.65 -14.13 ;
      RECT 26.35 -14.94 26.45 -14.13 ;
      RECT 25.15 -14.94 25.25 -14.13 ;
      RECT 23.95 -14.94 24.05 -14.13 ;
      RECT 22.75 -14.94 22.85 -14.13 ;
      RECT 21.55 -14.94 21.65 -14.13 ;
      RECT 20.35 -14.94 20.45 -14.13 ;
      RECT 19.15 -14.94 19.25 -14.13 ;
      RECT 17.95 -14.94 18.05 -14.13 ;
      RECT 16.75 -14.94 16.85 -14.13 ;
      RECT 15.55 -14.94 15.65 -14.13 ;
      RECT 14.35 -14.94 14.45 -14.13 ;
      RECT 13.15 -14.94 13.25 -14.13 ;
      RECT 11.95 -14.94 12.05 -14.13 ;
      RECT 10.75 -14.94 10.85 -14.13 ;
      RECT 9.55 -14.94 9.65 -14.13 ;
      RECT 8.35 -14.94 8.45 -14.13 ;
      RECT 7.15 -14.94 7.25 -14.13 ;
      RECT 5.95 -14.94 6.05 -14.13 ;
      RECT 4.75 -14.94 4.85 -14.13 ;
      RECT 3.55 -14.94 3.65 -14.13 ;
      RECT 2.35 -14.94 2.45 -14.13 ;
      RECT 1.15 -14.94 1.25 -14.13 ;
      RECT -0.05 -14.94 0.05 -14.13 ;
      RECT -0.105 -14.595 156.465 -14.475 ;
      RECT 153.55 -11.71 153.65 -10.9 ;
      RECT 152.35 -11.71 152.45 -10.9 ;
      RECT 151.15 -11.71 151.25 -10.9 ;
      RECT 149.95 -11.71 150.05 -10.9 ;
      RECT 148.75 -11.71 148.85 -10.9 ;
      RECT 147.55 -11.71 147.65 -10.9 ;
      RECT 146.35 -11.71 146.45 -10.9 ;
      RECT 145.15 -11.71 145.25 -10.9 ;
      RECT 143.95 -11.71 144.05 -10.9 ;
      RECT 142.75 -11.71 142.85 -10.9 ;
      RECT 141.55 -11.71 141.65 -10.9 ;
      RECT 140.35 -11.71 140.45 -10.9 ;
      RECT 139.15 -11.71 139.25 -10.9 ;
      RECT 137.95 -11.71 138.05 -10.9 ;
      RECT 136.75 -11.71 136.85 -10.9 ;
      RECT 135.55 -11.71 135.65 -10.9 ;
      RECT 134.35 -11.71 134.45 -10.9 ;
      RECT 133.15 -11.71 133.25 -10.9 ;
      RECT 131.95 -11.71 132.05 -10.9 ;
      RECT 130.75 -11.71 130.85 -10.9 ;
      RECT 129.55 -11.71 129.65 -10.9 ;
      RECT 128.35 -11.71 128.45 -10.9 ;
      RECT 127.15 -11.71 127.25 -10.9 ;
      RECT 125.95 -11.71 126.05 -10.9 ;
      RECT 124.75 -11.71 124.85 -10.9 ;
      RECT 123.55 -11.71 123.65 -10.9 ;
      RECT 122.35 -11.71 122.45 -10.9 ;
      RECT 121.15 -11.71 121.25 -10.9 ;
      RECT 119.95 -11.71 120.05 -10.9 ;
      RECT 118.75 -11.71 118.85 -10.9 ;
      RECT 117.55 -11.71 117.65 -10.9 ;
      RECT 116.35 -11.71 116.45 -10.9 ;
      RECT 115.15 -11.71 115.25 -10.9 ;
      RECT 113.95 -11.71 114.05 -10.9 ;
      RECT 112.75 -11.71 112.85 -10.9 ;
      RECT 111.55 -11.71 111.65 -10.9 ;
      RECT 110.35 -11.71 110.45 -10.9 ;
      RECT 109.15 -11.71 109.25 -10.9 ;
      RECT 107.95 -11.71 108.05 -10.9 ;
      RECT 106.75 -11.71 106.85 -10.9 ;
      RECT 105.55 -11.71 105.65 -10.9 ;
      RECT 104.35 -11.71 104.45 -10.9 ;
      RECT 103.15 -11.71 103.25 -10.9 ;
      RECT 101.95 -11.71 102.05 -10.9 ;
      RECT 100.75 -11.71 100.85 -10.9 ;
      RECT 99.55 -11.71 99.65 -10.9 ;
      RECT 98.35 -11.71 98.45 -10.9 ;
      RECT 97.15 -11.71 97.25 -10.9 ;
      RECT 95.95 -11.71 96.05 -10.9 ;
      RECT 94.75 -11.71 94.85 -10.9 ;
      RECT 93.55 -11.71 93.65 -10.9 ;
      RECT 92.35 -11.71 92.45 -10.9 ;
      RECT 91.15 -11.71 91.25 -10.9 ;
      RECT 89.95 -11.71 90.05 -10.9 ;
      RECT 88.75 -11.71 88.85 -10.9 ;
      RECT 87.55 -11.71 87.65 -10.9 ;
      RECT 86.35 -11.71 86.45 -10.9 ;
      RECT 85.15 -11.71 85.25 -10.9 ;
      RECT 83.95 -11.71 84.05 -10.9 ;
      RECT 82.75 -11.71 82.85 -10.9 ;
      RECT 81.55 -11.71 81.65 -10.9 ;
      RECT 80.35 -11.71 80.45 -10.9 ;
      RECT 79.15 -11.71 79.25 -10.9 ;
      RECT 77.95 -11.71 78.05 -10.9 ;
      RECT 76.75 -11.71 76.85 -10.9 ;
      RECT 75.55 -11.71 75.65 -10.9 ;
      RECT 74.35 -11.71 74.45 -10.9 ;
      RECT 73.15 -11.71 73.25 -10.9 ;
      RECT 71.95 -11.71 72.05 -10.9 ;
      RECT 70.75 -11.71 70.85 -10.9 ;
      RECT 69.55 -11.71 69.65 -10.9 ;
      RECT 68.35 -11.71 68.45 -10.9 ;
      RECT 67.15 -11.71 67.25 -10.9 ;
      RECT 65.95 -11.71 66.05 -10.9 ;
      RECT 64.75 -11.71 64.85 -10.9 ;
      RECT 63.55 -11.71 63.65 -10.9 ;
      RECT 62.35 -11.71 62.45 -10.9 ;
      RECT 61.15 -11.71 61.25 -10.9 ;
      RECT 59.95 -11.71 60.05 -10.9 ;
      RECT 58.75 -11.71 58.85 -10.9 ;
      RECT 57.55 -11.71 57.65 -10.9 ;
      RECT 56.35 -11.71 56.45 -10.9 ;
      RECT 55.15 -11.71 55.25 -10.9 ;
      RECT 53.95 -11.71 54.05 -10.9 ;
      RECT 52.75 -11.71 52.85 -10.9 ;
      RECT 51.55 -11.71 51.65 -10.9 ;
      RECT 50.35 -11.71 50.45 -10.9 ;
      RECT 49.15 -11.71 49.25 -10.9 ;
      RECT 47.95 -11.71 48.05 -10.9 ;
      RECT 46.75 -11.71 46.85 -10.9 ;
      RECT 45.55 -11.71 45.65 -10.9 ;
      RECT 44.35 -11.71 44.45 -10.9 ;
      RECT 43.15 -11.71 43.25 -10.9 ;
      RECT 41.95 -11.71 42.05 -10.9 ;
      RECT 40.75 -11.71 40.85 -10.9 ;
      RECT 39.55 -11.71 39.65 -10.9 ;
      RECT 38.35 -11.71 38.45 -10.9 ;
      RECT 37.15 -11.71 37.25 -10.9 ;
      RECT 35.95 -11.71 36.05 -10.9 ;
      RECT 34.75 -11.71 34.85 -10.9 ;
      RECT 33.55 -11.71 33.65 -10.9 ;
      RECT 32.35 -11.71 32.45 -10.9 ;
      RECT 31.15 -11.71 31.25 -10.9 ;
      RECT 29.95 -11.71 30.05 -10.9 ;
      RECT 28.75 -11.71 28.85 -10.9 ;
      RECT 27.55 -11.71 27.65 -10.9 ;
      RECT 26.35 -11.71 26.45 -10.9 ;
      RECT 25.15 -11.71 25.25 -10.9 ;
      RECT 23.95 -11.71 24.05 -10.9 ;
      RECT 22.75 -11.71 22.85 -10.9 ;
      RECT 21.55 -11.71 21.65 -10.9 ;
      RECT 20.35 -11.71 20.45 -10.9 ;
      RECT 19.15 -11.71 19.25 -10.9 ;
      RECT 17.95 -11.71 18.05 -10.9 ;
      RECT 16.75 -11.71 16.85 -10.9 ;
      RECT 15.55 -11.71 15.65 -10.9 ;
      RECT 14.35 -11.71 14.45 -10.9 ;
      RECT 13.15 -11.71 13.25 -10.9 ;
      RECT 11.95 -11.71 12.05 -10.9 ;
      RECT 10.75 -11.71 10.85 -10.9 ;
      RECT 9.55 -11.71 9.65 -10.9 ;
      RECT 8.35 -11.71 8.45 -10.9 ;
      RECT 7.15 -11.71 7.25 -10.9 ;
      RECT 5.95 -11.71 6.05 -10.9 ;
      RECT 4.75 -11.71 4.85 -10.9 ;
      RECT 3.55 -11.71 3.65 -10.9 ;
      RECT 2.35 -11.71 2.45 -10.9 ;
      RECT 1.15 -11.71 1.25 -10.9 ;
      RECT -0.05 -11.71 0.05 -10.9 ;
      RECT -0.105 -11.365 156.465 -11.245 ;
      RECT 153.55 -8.48 153.65 -7.67 ;
      RECT 152.35 -8.48 152.45 -7.67 ;
      RECT 151.15 -8.48 151.25 -7.67 ;
      RECT 149.95 -8.48 150.05 -7.67 ;
      RECT 148.75 -8.48 148.85 -7.67 ;
      RECT 147.55 -8.48 147.65 -7.67 ;
      RECT 146.35 -8.48 146.45 -7.67 ;
      RECT 145.15 -8.48 145.25 -7.67 ;
      RECT 143.95 -8.48 144.05 -7.67 ;
      RECT 142.75 -8.48 142.85 -7.67 ;
      RECT 141.55 -8.48 141.65 -7.67 ;
      RECT 140.35 -8.48 140.45 -7.67 ;
      RECT 139.15 -8.48 139.25 -7.67 ;
      RECT 137.95 -8.48 138.05 -7.67 ;
      RECT 136.75 -8.48 136.85 -7.67 ;
      RECT 135.55 -8.48 135.65 -7.67 ;
      RECT 134.35 -8.48 134.45 -7.67 ;
      RECT 133.15 -8.48 133.25 -7.67 ;
      RECT 131.95 -8.48 132.05 -7.67 ;
      RECT 130.75 -8.48 130.85 -7.67 ;
      RECT 129.55 -8.48 129.65 -7.67 ;
      RECT 128.35 -8.48 128.45 -7.67 ;
      RECT 127.15 -8.48 127.25 -7.67 ;
      RECT 125.95 -8.48 126.05 -7.67 ;
      RECT 124.75 -8.48 124.85 -7.67 ;
      RECT 123.55 -8.48 123.65 -7.67 ;
      RECT 122.35 -8.48 122.45 -7.67 ;
      RECT 121.15 -8.48 121.25 -7.67 ;
      RECT 119.95 -8.48 120.05 -7.67 ;
      RECT 118.75 -8.48 118.85 -7.67 ;
      RECT 117.55 -8.48 117.65 -7.67 ;
      RECT 116.35 -8.48 116.45 -7.67 ;
      RECT 115.15 -8.48 115.25 -7.67 ;
      RECT 113.95 -8.48 114.05 -7.67 ;
      RECT 112.75 -8.48 112.85 -7.67 ;
      RECT 111.55 -8.48 111.65 -7.67 ;
      RECT 110.35 -8.48 110.45 -7.67 ;
      RECT 109.15 -8.48 109.25 -7.67 ;
      RECT 107.95 -8.48 108.05 -7.67 ;
      RECT 106.75 -8.48 106.85 -7.67 ;
      RECT 105.55 -8.48 105.65 -7.67 ;
      RECT 104.35 -8.48 104.45 -7.67 ;
      RECT 103.15 -8.48 103.25 -7.67 ;
      RECT 101.95 -8.48 102.05 -7.67 ;
      RECT 100.75 -8.48 100.85 -7.67 ;
      RECT 99.55 -8.48 99.65 -7.67 ;
      RECT 98.35 -8.48 98.45 -7.67 ;
      RECT 97.15 -8.48 97.25 -7.67 ;
      RECT 95.95 -8.48 96.05 -7.67 ;
      RECT 94.75 -8.48 94.85 -7.67 ;
      RECT 93.55 -8.48 93.65 -7.67 ;
      RECT 92.35 -8.48 92.45 -7.67 ;
      RECT 91.15 -8.48 91.25 -7.67 ;
      RECT 89.95 -8.48 90.05 -7.67 ;
      RECT 88.75 -8.48 88.85 -7.67 ;
      RECT 87.55 -8.48 87.65 -7.67 ;
      RECT 86.35 -8.48 86.45 -7.67 ;
      RECT 85.15 -8.48 85.25 -7.67 ;
      RECT 83.95 -8.48 84.05 -7.67 ;
      RECT 82.75 -8.48 82.85 -7.67 ;
      RECT 81.55 -8.48 81.65 -7.67 ;
      RECT 80.35 -8.48 80.45 -7.67 ;
      RECT 79.15 -8.48 79.25 -7.67 ;
      RECT 77.95 -8.48 78.05 -7.67 ;
      RECT 76.75 -8.48 76.85 -7.67 ;
      RECT 75.55 -8.48 75.65 -7.67 ;
      RECT 74.35 -8.48 74.45 -7.67 ;
      RECT 73.15 -8.48 73.25 -7.67 ;
      RECT 71.95 -8.48 72.05 -7.67 ;
      RECT 70.75 -8.48 70.85 -7.67 ;
      RECT 69.55 -8.48 69.65 -7.67 ;
      RECT 68.35 -8.48 68.45 -7.67 ;
      RECT 67.15 -8.48 67.25 -7.67 ;
      RECT 65.95 -8.48 66.05 -7.67 ;
      RECT 64.75 -8.48 64.85 -7.67 ;
      RECT 63.55 -8.48 63.65 -7.67 ;
      RECT 62.35 -8.48 62.45 -7.67 ;
      RECT 61.15 -8.48 61.25 -7.67 ;
      RECT 59.95 -8.48 60.05 -7.67 ;
      RECT 58.75 -8.48 58.85 -7.67 ;
      RECT 57.55 -8.48 57.65 -7.67 ;
      RECT 56.35 -8.48 56.45 -7.67 ;
      RECT 55.15 -8.48 55.25 -7.67 ;
      RECT 53.95 -8.48 54.05 -7.67 ;
      RECT 52.75 -8.48 52.85 -7.67 ;
      RECT 51.55 -8.48 51.65 -7.67 ;
      RECT 50.35 -8.48 50.45 -7.67 ;
      RECT 49.15 -8.48 49.25 -7.67 ;
      RECT 47.95 -8.48 48.05 -7.67 ;
      RECT 46.75 -8.48 46.85 -7.67 ;
      RECT 45.55 -8.48 45.65 -7.67 ;
      RECT 44.35 -8.48 44.45 -7.67 ;
      RECT 43.15 -8.48 43.25 -7.67 ;
      RECT 41.95 -8.48 42.05 -7.67 ;
      RECT 40.75 -8.48 40.85 -7.67 ;
      RECT 39.55 -8.48 39.65 -7.67 ;
      RECT 38.35 -8.48 38.45 -7.67 ;
      RECT 37.15 -8.48 37.25 -7.67 ;
      RECT 35.95 -8.48 36.05 -7.67 ;
      RECT 34.75 -8.48 34.85 -7.67 ;
      RECT 33.55 -8.48 33.65 -7.67 ;
      RECT 32.35 -8.48 32.45 -7.67 ;
      RECT 31.15 -8.48 31.25 -7.67 ;
      RECT 29.95 -8.48 30.05 -7.67 ;
      RECT 28.75 -8.48 28.85 -7.67 ;
      RECT 27.55 -8.48 27.65 -7.67 ;
      RECT 26.35 -8.48 26.45 -7.67 ;
      RECT 25.15 -8.48 25.25 -7.67 ;
      RECT 23.95 -8.48 24.05 -7.67 ;
      RECT 22.75 -8.48 22.85 -7.67 ;
      RECT 21.55 -8.48 21.65 -7.67 ;
      RECT 20.35 -8.48 20.45 -7.67 ;
      RECT 19.15 -8.48 19.25 -7.67 ;
      RECT 17.95 -8.48 18.05 -7.67 ;
      RECT 16.75 -8.48 16.85 -7.67 ;
      RECT 15.55 -8.48 15.65 -7.67 ;
      RECT 14.35 -8.48 14.45 -7.67 ;
      RECT 13.15 -8.48 13.25 -7.67 ;
      RECT 11.95 -8.48 12.05 -7.67 ;
      RECT 10.75 -8.48 10.85 -7.67 ;
      RECT 9.55 -8.48 9.65 -7.67 ;
      RECT 8.35 -8.48 8.45 -7.67 ;
      RECT 7.15 -8.48 7.25 -7.67 ;
      RECT 5.95 -8.48 6.05 -7.67 ;
      RECT 4.75 -8.48 4.85 -7.67 ;
      RECT 3.55 -8.48 3.65 -7.67 ;
      RECT 2.35 -8.48 2.45 -7.67 ;
      RECT 1.15 -8.48 1.25 -7.67 ;
      RECT -0.05 -8.48 0.05 -7.67 ;
      RECT -0.105 -8.135 156.465 -8.015 ;
      RECT 153.55 -5.25 153.65 -4.44 ;
      RECT 152.35 -5.25 152.45 -4.44 ;
      RECT 151.15 -5.25 151.25 -4.44 ;
      RECT 149.95 -5.25 150.05 -4.44 ;
      RECT 148.75 -5.25 148.85 -4.44 ;
      RECT 147.55 -5.25 147.65 -4.44 ;
      RECT 146.35 -5.25 146.45 -4.44 ;
      RECT 145.15 -5.25 145.25 -4.44 ;
      RECT 143.95 -5.25 144.05 -4.44 ;
      RECT 142.75 -5.25 142.85 -4.44 ;
      RECT 141.55 -5.25 141.65 -4.44 ;
      RECT 140.35 -5.25 140.45 -4.44 ;
      RECT 139.15 -5.25 139.25 -4.44 ;
      RECT 137.95 -5.25 138.05 -4.44 ;
      RECT 136.75 -5.25 136.85 -4.44 ;
      RECT 135.55 -5.25 135.65 -4.44 ;
      RECT 134.35 -5.25 134.45 -4.44 ;
      RECT 133.15 -5.25 133.25 -4.44 ;
      RECT 131.95 -5.25 132.05 -4.44 ;
      RECT 130.75 -5.25 130.85 -4.44 ;
      RECT 129.55 -5.25 129.65 -4.44 ;
      RECT 128.35 -5.25 128.45 -4.44 ;
      RECT 127.15 -5.25 127.25 -4.44 ;
      RECT 125.95 -5.25 126.05 -4.44 ;
      RECT 124.75 -5.25 124.85 -4.44 ;
      RECT 123.55 -5.25 123.65 -4.44 ;
      RECT 122.35 -5.25 122.45 -4.44 ;
      RECT 121.15 -5.25 121.25 -4.44 ;
      RECT 119.95 -5.25 120.05 -4.44 ;
      RECT 118.75 -5.25 118.85 -4.44 ;
      RECT 117.55 -5.25 117.65 -4.44 ;
      RECT 116.35 -5.25 116.45 -4.44 ;
      RECT 115.15 -5.25 115.25 -4.44 ;
      RECT 113.95 -5.25 114.05 -4.44 ;
      RECT 112.75 -5.25 112.85 -4.44 ;
      RECT 111.55 -5.25 111.65 -4.44 ;
      RECT 110.35 -5.25 110.45 -4.44 ;
      RECT 109.15 -5.25 109.25 -4.44 ;
      RECT 107.95 -5.25 108.05 -4.44 ;
      RECT 106.75 -5.25 106.85 -4.44 ;
      RECT 105.55 -5.25 105.65 -4.44 ;
      RECT 104.35 -5.25 104.45 -4.44 ;
      RECT 103.15 -5.25 103.25 -4.44 ;
      RECT 101.95 -5.25 102.05 -4.44 ;
      RECT 100.75 -5.25 100.85 -4.44 ;
      RECT 99.55 -5.25 99.65 -4.44 ;
      RECT 98.35 -5.25 98.45 -4.44 ;
      RECT 97.15 -5.25 97.25 -4.44 ;
      RECT 95.95 -5.25 96.05 -4.44 ;
      RECT 94.75 -5.25 94.85 -4.44 ;
      RECT 93.55 -5.25 93.65 -4.44 ;
      RECT 92.35 -5.25 92.45 -4.44 ;
      RECT 91.15 -5.25 91.25 -4.44 ;
      RECT 89.95 -5.25 90.05 -4.44 ;
      RECT 88.75 -5.25 88.85 -4.44 ;
      RECT 87.55 -5.25 87.65 -4.44 ;
      RECT 86.35 -5.25 86.45 -4.44 ;
      RECT 85.15 -5.25 85.25 -4.44 ;
      RECT 83.95 -5.25 84.05 -4.44 ;
      RECT 82.75 -5.25 82.85 -4.44 ;
      RECT 81.55 -5.25 81.65 -4.44 ;
      RECT 80.35 -5.25 80.45 -4.44 ;
      RECT 79.15 -5.25 79.25 -4.44 ;
      RECT 77.95 -5.25 78.05 -4.44 ;
      RECT 76.75 -5.25 76.85 -4.44 ;
      RECT 75.55 -5.25 75.65 -4.44 ;
      RECT 74.35 -5.25 74.45 -4.44 ;
      RECT 73.15 -5.25 73.25 -4.44 ;
      RECT 71.95 -5.25 72.05 -4.44 ;
      RECT 70.75 -5.25 70.85 -4.44 ;
      RECT 69.55 -5.25 69.65 -4.44 ;
      RECT 68.35 -5.25 68.45 -4.44 ;
      RECT 67.15 -5.25 67.25 -4.44 ;
      RECT 65.95 -5.25 66.05 -4.44 ;
      RECT 64.75 -5.25 64.85 -4.44 ;
      RECT 63.55 -5.25 63.65 -4.44 ;
      RECT 62.35 -5.25 62.45 -4.44 ;
      RECT 61.15 -5.25 61.25 -4.44 ;
      RECT 59.95 -5.25 60.05 -4.44 ;
      RECT 58.75 -5.25 58.85 -4.44 ;
      RECT 57.55 -5.25 57.65 -4.44 ;
      RECT 56.35 -5.25 56.45 -4.44 ;
      RECT 55.15 -5.25 55.25 -4.44 ;
      RECT 53.95 -5.25 54.05 -4.44 ;
      RECT 52.75 -5.25 52.85 -4.44 ;
      RECT 51.55 -5.25 51.65 -4.44 ;
      RECT 50.35 -5.25 50.45 -4.44 ;
      RECT 49.15 -5.25 49.25 -4.44 ;
      RECT 47.95 -5.25 48.05 -4.44 ;
      RECT 46.75 -5.25 46.85 -4.44 ;
      RECT 45.55 -5.25 45.65 -4.44 ;
      RECT 44.35 -5.25 44.45 -4.44 ;
      RECT 43.15 -5.25 43.25 -4.44 ;
      RECT 41.95 -5.25 42.05 -4.44 ;
      RECT 40.75 -5.25 40.85 -4.44 ;
      RECT 39.55 -5.25 39.65 -4.44 ;
      RECT 38.35 -5.25 38.45 -4.44 ;
      RECT 37.15 -5.25 37.25 -4.44 ;
      RECT 35.95 -5.25 36.05 -4.44 ;
      RECT 34.75 -5.25 34.85 -4.44 ;
      RECT 33.55 -5.25 33.65 -4.44 ;
      RECT 32.35 -5.25 32.45 -4.44 ;
      RECT 31.15 -5.25 31.25 -4.44 ;
      RECT 29.95 -5.25 30.05 -4.44 ;
      RECT 28.75 -5.25 28.85 -4.44 ;
      RECT 27.55 -5.25 27.65 -4.44 ;
      RECT 26.35 -5.25 26.45 -4.44 ;
      RECT 25.15 -5.25 25.25 -4.44 ;
      RECT 23.95 -5.25 24.05 -4.44 ;
      RECT 22.75 -5.25 22.85 -4.44 ;
      RECT 21.55 -5.25 21.65 -4.44 ;
      RECT 20.35 -5.25 20.45 -4.44 ;
      RECT 19.15 -5.25 19.25 -4.44 ;
      RECT 17.95 -5.25 18.05 -4.44 ;
      RECT 16.75 -5.25 16.85 -4.44 ;
      RECT 15.55 -5.25 15.65 -4.44 ;
      RECT 14.35 -5.25 14.45 -4.44 ;
      RECT 13.15 -5.25 13.25 -4.44 ;
      RECT 11.95 -5.25 12.05 -4.44 ;
      RECT 10.75 -5.25 10.85 -4.44 ;
      RECT 9.55 -5.25 9.65 -4.44 ;
      RECT 8.35 -5.25 8.45 -4.44 ;
      RECT 7.15 -5.25 7.25 -4.44 ;
      RECT 5.95 -5.25 6.05 -4.44 ;
      RECT 4.75 -5.25 4.85 -4.44 ;
      RECT 3.55 -5.25 3.65 -4.44 ;
      RECT 2.35 -5.25 2.45 -4.44 ;
      RECT 1.15 -5.25 1.25 -4.44 ;
      RECT -0.05 -5.25 0.05 -4.44 ;
      RECT -0.105 -4.905 156.465 -4.785 ;
      RECT 153.55 -2.02 153.65 -1.21 ;
      RECT 152.35 -2.02 152.45 -1.21 ;
      RECT 151.15 -2.02 151.25 -1.21 ;
      RECT 149.95 -2.02 150.05 -1.21 ;
      RECT 148.75 -2.02 148.85 -1.21 ;
      RECT 147.55 -2.02 147.65 -1.21 ;
      RECT 146.35 -2.02 146.45 -1.21 ;
      RECT 145.15 -2.02 145.25 -1.21 ;
      RECT 143.95 -2.02 144.05 -1.21 ;
      RECT 142.75 -2.02 142.85 -1.21 ;
      RECT 141.55 -2.02 141.65 -1.21 ;
      RECT 140.35 -2.02 140.45 -1.21 ;
      RECT 139.15 -2.02 139.25 -1.21 ;
      RECT 137.95 -2.02 138.05 -1.21 ;
      RECT 136.75 -2.02 136.85 -1.21 ;
      RECT 135.55 -2.02 135.65 -1.21 ;
      RECT 134.35 -2.02 134.45 -1.21 ;
      RECT 133.15 -2.02 133.25 -1.21 ;
      RECT 131.95 -2.02 132.05 -1.21 ;
      RECT 130.75 -2.02 130.85 -1.21 ;
      RECT 129.55 -2.02 129.65 -1.21 ;
      RECT 128.35 -2.02 128.45 -1.21 ;
      RECT 127.15 -2.02 127.25 -1.21 ;
      RECT 125.95 -2.02 126.05 -1.21 ;
      RECT 124.75 -2.02 124.85 -1.21 ;
      RECT 123.55 -2.02 123.65 -1.21 ;
      RECT 122.35 -2.02 122.45 -1.21 ;
      RECT 121.15 -2.02 121.25 -1.21 ;
      RECT 119.95 -2.02 120.05 -1.21 ;
      RECT 118.75 -2.02 118.85 -1.21 ;
      RECT 117.55 -2.02 117.65 -1.21 ;
      RECT 116.35 -2.02 116.45 -1.21 ;
      RECT 115.15 -2.02 115.25 -1.21 ;
      RECT 113.95 -2.02 114.05 -1.21 ;
      RECT 112.75 -2.02 112.85 -1.21 ;
      RECT 111.55 -2.02 111.65 -1.21 ;
      RECT 110.35 -2.02 110.45 -1.21 ;
      RECT 109.15 -2.02 109.25 -1.21 ;
      RECT 107.95 -2.02 108.05 -1.21 ;
      RECT 106.75 -2.02 106.85 -1.21 ;
      RECT 105.55 -2.02 105.65 -1.21 ;
      RECT 104.35 -2.02 104.45 -1.21 ;
      RECT 103.15 -2.02 103.25 -1.21 ;
      RECT 101.95 -2.02 102.05 -1.21 ;
      RECT 100.75 -2.02 100.85 -1.21 ;
      RECT 99.55 -2.02 99.65 -1.21 ;
      RECT 98.35 -2.02 98.45 -1.21 ;
      RECT 97.15 -2.02 97.25 -1.21 ;
      RECT 95.95 -2.02 96.05 -1.21 ;
      RECT 94.75 -2.02 94.85 -1.21 ;
      RECT 93.55 -2.02 93.65 -1.21 ;
      RECT 92.35 -2.02 92.45 -1.21 ;
      RECT 91.15 -2.02 91.25 -1.21 ;
      RECT 89.95 -2.02 90.05 -1.21 ;
      RECT 88.75 -2.02 88.85 -1.21 ;
      RECT 87.55 -2.02 87.65 -1.21 ;
      RECT 86.35 -2.02 86.45 -1.21 ;
      RECT 85.15 -2.02 85.25 -1.21 ;
      RECT 83.95 -2.02 84.05 -1.21 ;
      RECT 82.75 -2.02 82.85 -1.21 ;
      RECT 81.55 -2.02 81.65 -1.21 ;
      RECT 80.35 -2.02 80.45 -1.21 ;
      RECT 79.15 -2.02 79.25 -1.21 ;
      RECT 77.95 -2.02 78.05 -1.21 ;
      RECT 76.75 -2.02 76.85 -1.21 ;
      RECT 75.55 -2.02 75.65 -1.21 ;
      RECT 74.35 -2.02 74.45 -1.21 ;
      RECT 73.15 -2.02 73.25 -1.21 ;
      RECT 71.95 -2.02 72.05 -1.21 ;
      RECT 70.75 -2.02 70.85 -1.21 ;
      RECT 69.55 -2.02 69.65 -1.21 ;
      RECT 68.35 -2.02 68.45 -1.21 ;
      RECT 67.15 -2.02 67.25 -1.21 ;
      RECT 65.95 -2.02 66.05 -1.21 ;
      RECT 64.75 -2.02 64.85 -1.21 ;
      RECT 63.55 -2.02 63.65 -1.21 ;
      RECT 62.35 -2.02 62.45 -1.21 ;
      RECT 61.15 -2.02 61.25 -1.21 ;
      RECT 59.95 -2.02 60.05 -1.21 ;
      RECT 58.75 -2.02 58.85 -1.21 ;
      RECT 57.55 -2.02 57.65 -1.21 ;
      RECT 56.35 -2.02 56.45 -1.21 ;
      RECT 55.15 -2.02 55.25 -1.21 ;
      RECT 53.95 -2.02 54.05 -1.21 ;
      RECT 52.75 -2.02 52.85 -1.21 ;
      RECT 51.55 -2.02 51.65 -1.21 ;
      RECT 50.35 -2.02 50.45 -1.21 ;
      RECT 49.15 -2.02 49.25 -1.21 ;
      RECT 47.95 -2.02 48.05 -1.21 ;
      RECT 46.75 -2.02 46.85 -1.21 ;
      RECT 45.55 -2.02 45.65 -1.21 ;
      RECT 44.35 -2.02 44.45 -1.21 ;
      RECT 43.15 -2.02 43.25 -1.21 ;
      RECT 41.95 -2.02 42.05 -1.21 ;
      RECT 40.75 -2.02 40.85 -1.21 ;
      RECT 39.55 -2.02 39.65 -1.21 ;
      RECT 38.35 -2.02 38.45 -1.21 ;
      RECT 37.15 -2.02 37.25 -1.21 ;
      RECT 35.95 -2.02 36.05 -1.21 ;
      RECT 34.75 -2.02 34.85 -1.21 ;
      RECT 33.55 -2.02 33.65 -1.21 ;
      RECT 32.35 -2.02 32.45 -1.21 ;
      RECT 31.15 -2.02 31.25 -1.21 ;
      RECT 29.95 -2.02 30.05 -1.21 ;
      RECT 28.75 -2.02 28.85 -1.21 ;
      RECT 27.55 -2.02 27.65 -1.21 ;
      RECT 26.35 -2.02 26.45 -1.21 ;
      RECT 25.15 -2.02 25.25 -1.21 ;
      RECT 23.95 -2.02 24.05 -1.21 ;
      RECT 22.75 -2.02 22.85 -1.21 ;
      RECT 21.55 -2.02 21.65 -1.21 ;
      RECT 20.35 -2.02 20.45 -1.21 ;
      RECT 19.15 -2.02 19.25 -1.21 ;
      RECT 17.95 -2.02 18.05 -1.21 ;
      RECT 16.75 -2.02 16.85 -1.21 ;
      RECT 15.55 -2.02 15.65 -1.21 ;
      RECT 14.35 -2.02 14.45 -1.21 ;
      RECT 13.15 -2.02 13.25 -1.21 ;
      RECT 11.95 -2.02 12.05 -1.21 ;
      RECT 10.75 -2.02 10.85 -1.21 ;
      RECT 9.55 -2.02 9.65 -1.21 ;
      RECT 8.35 -2.02 8.45 -1.21 ;
      RECT 7.15 -2.02 7.25 -1.21 ;
      RECT 5.95 -2.02 6.05 -1.21 ;
      RECT 4.75 -2.02 4.85 -1.21 ;
      RECT 3.55 -2.02 3.65 -1.21 ;
      RECT 2.35 -2.02 2.45 -1.21 ;
      RECT 1.15 -2.02 1.25 -1.21 ;
      RECT -0.05 -2.02 0.05 -1.21 ;
      RECT -0.105 -1.675 156.465 -1.555 ;
      RECT -0.105 1.555 156.465 1.675 ;
      RECT 153.55 1.21 153.65 1.675 ;
      RECT 152.35 1.21 152.45 1.675 ;
      RECT 151.15 1.21 151.25 1.675 ;
      RECT 149.95 1.21 150.05 1.675 ;
      RECT 148.75 1.21 148.85 1.675 ;
      RECT 147.55 1.21 147.65 1.675 ;
      RECT 146.35 1.21 146.45 1.675 ;
      RECT 145.15 1.21 145.25 1.675 ;
      RECT 143.95 1.21 144.05 1.675 ;
      RECT 142.75 1.21 142.85 1.675 ;
      RECT 141.55 1.21 141.65 1.675 ;
      RECT 140.35 1.21 140.45 1.675 ;
      RECT 139.15 1.21 139.25 1.675 ;
      RECT 137.95 1.21 138.05 1.675 ;
      RECT 136.75 1.21 136.85 1.675 ;
      RECT 135.55 1.21 135.65 1.675 ;
      RECT 134.35 1.21 134.45 1.675 ;
      RECT 133.15 1.21 133.25 1.675 ;
      RECT 131.95 1.21 132.05 1.675 ;
      RECT 130.75 1.21 130.85 1.675 ;
      RECT 129.55 1.21 129.65 1.675 ;
      RECT 128.35 1.21 128.45 1.675 ;
      RECT 127.15 1.21 127.25 1.675 ;
      RECT 125.95 1.21 126.05 1.675 ;
      RECT 124.75 1.21 124.85 1.675 ;
      RECT 123.55 1.21 123.65 1.675 ;
      RECT 122.35 1.21 122.45 1.675 ;
      RECT 121.15 1.21 121.25 1.675 ;
      RECT 119.95 1.21 120.05 1.675 ;
      RECT 118.75 1.21 118.85 1.675 ;
      RECT 117.55 1.21 117.65 1.675 ;
      RECT 116.35 1.21 116.45 1.675 ;
      RECT 115.15 1.21 115.25 1.675 ;
      RECT 113.95 1.21 114.05 1.675 ;
      RECT 112.75 1.21 112.85 1.675 ;
      RECT 111.55 1.21 111.65 1.675 ;
      RECT 110.35 1.21 110.45 1.675 ;
      RECT 109.15 1.21 109.25 1.675 ;
      RECT 107.95 1.21 108.05 1.675 ;
      RECT 106.75 1.21 106.85 1.675 ;
      RECT 105.55 1.21 105.65 1.675 ;
      RECT 104.35 1.21 104.45 1.675 ;
      RECT 103.15 1.21 103.25 1.675 ;
      RECT 101.95 1.21 102.05 1.675 ;
      RECT 100.75 1.21 100.85 1.675 ;
      RECT 99.55 1.21 99.65 1.675 ;
      RECT 98.35 1.21 98.45 1.675 ;
      RECT 97.15 1.21 97.25 1.675 ;
      RECT 95.95 1.21 96.05 1.675 ;
      RECT 94.75 1.21 94.85 1.675 ;
      RECT 93.55 1.21 93.65 1.675 ;
      RECT 92.35 1.21 92.45 1.675 ;
      RECT 91.15 1.21 91.25 1.675 ;
      RECT 89.95 1.21 90.05 1.675 ;
      RECT 88.75 1.21 88.85 1.675 ;
      RECT 87.55 1.21 87.65 1.675 ;
      RECT 86.35 1.21 86.45 1.675 ;
      RECT 85.15 1.21 85.25 1.675 ;
      RECT 83.95 1.21 84.05 1.675 ;
      RECT 82.75 1.21 82.85 1.675 ;
      RECT 81.55 1.21 81.65 1.675 ;
      RECT 80.35 1.21 80.45 1.675 ;
      RECT 79.15 1.21 79.25 1.675 ;
      RECT 77.95 1.21 78.05 1.675 ;
      RECT 76.75 1.21 76.85 1.675 ;
      RECT 75.55 1.21 75.65 1.675 ;
      RECT 74.35 1.21 74.45 1.675 ;
      RECT 73.15 1.21 73.25 1.675 ;
      RECT 71.95 1.21 72.05 1.675 ;
      RECT 70.75 1.21 70.85 1.675 ;
      RECT 69.55 1.21 69.65 1.675 ;
      RECT 68.35 1.21 68.45 1.675 ;
      RECT 67.15 1.21 67.25 1.675 ;
      RECT 65.95 1.21 66.05 1.675 ;
      RECT 64.75 1.21 64.85 1.675 ;
      RECT 63.55 1.21 63.65 1.675 ;
      RECT 62.35 1.21 62.45 1.675 ;
      RECT 61.15 1.21 61.25 1.675 ;
      RECT 59.95 1.21 60.05 1.675 ;
      RECT 58.75 1.21 58.85 1.675 ;
      RECT 57.55 1.21 57.65 1.675 ;
      RECT 56.35 1.21 56.45 1.675 ;
      RECT 55.15 1.21 55.25 1.675 ;
      RECT 53.95 1.21 54.05 1.675 ;
      RECT 52.75 1.21 52.85 1.675 ;
      RECT 51.55 1.21 51.65 1.675 ;
      RECT 50.35 1.21 50.45 1.675 ;
      RECT 49.15 1.21 49.25 1.675 ;
      RECT 47.95 1.21 48.05 1.675 ;
      RECT 46.75 1.21 46.85 1.675 ;
      RECT 45.55 1.21 45.65 1.675 ;
      RECT 44.35 1.21 44.45 1.675 ;
      RECT 43.15 1.21 43.25 1.675 ;
      RECT 41.95 1.21 42.05 1.675 ;
      RECT 40.75 1.21 40.85 1.675 ;
      RECT 39.55 1.21 39.65 1.675 ;
      RECT 38.35 1.21 38.45 1.675 ;
      RECT 37.15 1.21 37.25 1.675 ;
      RECT 35.95 1.21 36.05 1.675 ;
      RECT 34.75 1.21 34.85 1.675 ;
      RECT 33.55 1.21 33.65 1.675 ;
      RECT 32.35 1.21 32.45 1.675 ;
      RECT 31.15 1.21 31.25 1.675 ;
      RECT 29.95 1.21 30.05 1.675 ;
      RECT 28.75 1.21 28.85 1.675 ;
      RECT 27.55 1.21 27.65 1.675 ;
      RECT 26.35 1.21 26.45 1.675 ;
      RECT 25.15 1.21 25.25 1.675 ;
      RECT 23.95 1.21 24.05 1.675 ;
      RECT 22.75 1.21 22.85 1.675 ;
      RECT 21.55 1.21 21.65 1.675 ;
      RECT 20.35 1.21 20.45 1.675 ;
      RECT 19.15 1.21 19.25 1.675 ;
      RECT 17.95 1.21 18.05 1.675 ;
      RECT 16.75 1.21 16.85 1.675 ;
      RECT 15.55 1.21 15.65 1.675 ;
      RECT 14.35 1.21 14.45 1.675 ;
      RECT 13.15 1.21 13.25 1.675 ;
      RECT 11.95 1.21 12.05 1.675 ;
      RECT 10.75 1.21 10.85 1.675 ;
      RECT 9.55 1.21 9.65 1.675 ;
      RECT 8.35 1.21 8.45 1.675 ;
      RECT 7.15 1.21 7.25 1.675 ;
      RECT 5.95 1.21 6.05 1.675 ;
      RECT 4.75 1.21 4.85 1.675 ;
      RECT 3.55 1.21 3.65 1.675 ;
      RECT 2.35 1.21 2.45 1.675 ;
      RECT 1.15 1.21 1.25 1.675 ;
      RECT -0.05 1.21 0.05 1.675 ;
      RECT -0.01 3.42 156.465 3.8 ;
      RECT 153.425 2.175 153.525 3.8 ;
      RECT 152.475 2.175 152.575 3.8 ;
      RECT 152.225 2.175 152.325 3.8 ;
      RECT 151.275 2.175 151.375 3.8 ;
      RECT 151.025 2.175 151.125 3.8 ;
      RECT 150.075 2.175 150.175 3.8 ;
      RECT 149.825 2.175 149.925 3.8 ;
      RECT 148.875 2.175 148.975 3.8 ;
      RECT 148.625 2.175 148.725 3.8 ;
      RECT 147.675 2.175 147.775 3.8 ;
      RECT 147.425 2.175 147.525 3.8 ;
      RECT 146.475 2.175 146.575 3.8 ;
      RECT 146.225 2.175 146.325 3.8 ;
      RECT 145.275 2.175 145.375 3.8 ;
      RECT 145.025 2.175 145.125 3.8 ;
      RECT 144.075 2.175 144.175 3.8 ;
      RECT 143.825 2.175 143.925 3.8 ;
      RECT 142.875 2.175 142.975 3.8 ;
      RECT 142.625 2.175 142.725 3.8 ;
      RECT 141.675 2.175 141.775 3.8 ;
      RECT 141.425 2.175 141.525 3.8 ;
      RECT 140.475 2.175 140.575 3.8 ;
      RECT 140.225 2.175 140.325 3.8 ;
      RECT 139.275 2.175 139.375 3.8 ;
      RECT 139.025 2.175 139.125 3.8 ;
      RECT 138.075 2.175 138.175 3.8 ;
      RECT 137.825 2.175 137.925 3.8 ;
      RECT 136.875 2.175 136.975 3.8 ;
      RECT 136.625 2.175 136.725 3.8 ;
      RECT 135.675 2.175 135.775 3.8 ;
      RECT 135.425 2.175 135.525 3.8 ;
      RECT 134.475 2.175 134.575 3.8 ;
      RECT 134.225 2.175 134.325 3.8 ;
      RECT 133.275 2.175 133.375 3.8 ;
      RECT 133.025 2.175 133.125 3.8 ;
      RECT 132.075 2.175 132.175 3.8 ;
      RECT 131.825 2.175 131.925 3.8 ;
      RECT 130.875 2.175 130.975 3.8 ;
      RECT 130.625 2.175 130.725 3.8 ;
      RECT 129.675 2.175 129.775 3.8 ;
      RECT 129.425 2.175 129.525 3.8 ;
      RECT 128.475 2.175 128.575 3.8 ;
      RECT 128.225 2.175 128.325 3.8 ;
      RECT 127.275 2.175 127.375 3.8 ;
      RECT 127.025 2.175 127.125 3.8 ;
      RECT 126.075 2.175 126.175 3.8 ;
      RECT 125.825 2.175 125.925 3.8 ;
      RECT 124.875 2.175 124.975 3.8 ;
      RECT 124.625 2.175 124.725 3.8 ;
      RECT 123.675 2.175 123.775 3.8 ;
      RECT 123.425 2.175 123.525 3.8 ;
      RECT 122.475 2.175 122.575 3.8 ;
      RECT 122.225 2.175 122.325 3.8 ;
      RECT 121.275 2.175 121.375 3.8 ;
      RECT 121.025 2.175 121.125 3.8 ;
      RECT 120.075 2.175 120.175 3.8 ;
      RECT 119.825 2.175 119.925 3.8 ;
      RECT 118.875 2.175 118.975 3.8 ;
      RECT 118.625 2.175 118.725 3.8 ;
      RECT 117.675 2.175 117.775 3.8 ;
      RECT 117.425 2.175 117.525 3.8 ;
      RECT 116.475 2.175 116.575 3.8 ;
      RECT 116.225 2.175 116.325 3.8 ;
      RECT 115.275 2.175 115.375 3.8 ;
      RECT 115.025 2.175 115.125 3.8 ;
      RECT 114.075 2.175 114.175 3.8 ;
      RECT 113.825 2.175 113.925 3.8 ;
      RECT 112.875 2.175 112.975 3.8 ;
      RECT 112.625 2.175 112.725 3.8 ;
      RECT 111.675 2.175 111.775 3.8 ;
      RECT 111.425 2.175 111.525 3.8 ;
      RECT 110.475 2.175 110.575 3.8 ;
      RECT 110.225 2.175 110.325 3.8 ;
      RECT 109.275 2.175 109.375 3.8 ;
      RECT 109.025 2.175 109.125 3.8 ;
      RECT 108.075 2.175 108.175 3.8 ;
      RECT 107.825 2.175 107.925 3.8 ;
      RECT 106.875 2.175 106.975 3.8 ;
      RECT 106.625 2.175 106.725 3.8 ;
      RECT 105.675 2.175 105.775 3.8 ;
      RECT 105.425 2.175 105.525 3.8 ;
      RECT 104.475 2.175 104.575 3.8 ;
      RECT 104.225 2.175 104.325 3.8 ;
      RECT 103.275 2.175 103.375 3.8 ;
      RECT 103.025 2.175 103.125 3.8 ;
      RECT 102.075 2.175 102.175 3.8 ;
      RECT 101.825 2.175 101.925 3.8 ;
      RECT 100.875 2.175 100.975 3.8 ;
      RECT 100.625 2.175 100.725 3.8 ;
      RECT 99.675 2.175 99.775 3.8 ;
      RECT 99.425 2.175 99.525 3.8 ;
      RECT 98.475 2.175 98.575 3.8 ;
      RECT 98.225 2.175 98.325 3.8 ;
      RECT 97.275 2.175 97.375 3.8 ;
      RECT 97.025 2.175 97.125 3.8 ;
      RECT 96.075 2.175 96.175 3.8 ;
      RECT 95.825 2.175 95.925 3.8 ;
      RECT 94.875 2.175 94.975 3.8 ;
      RECT 94.625 2.175 94.725 3.8 ;
      RECT 93.675 2.175 93.775 3.8 ;
      RECT 93.425 2.175 93.525 3.8 ;
      RECT 92.475 2.175 92.575 3.8 ;
      RECT 92.225 2.175 92.325 3.8 ;
      RECT 91.275 2.175 91.375 3.8 ;
      RECT 91.025 2.175 91.125 3.8 ;
      RECT 90.075 2.175 90.175 3.8 ;
      RECT 89.825 2.175 89.925 3.8 ;
      RECT 88.875 2.175 88.975 3.8 ;
      RECT 88.625 2.175 88.725 3.8 ;
      RECT 87.675 2.175 87.775 3.8 ;
      RECT 87.425 2.175 87.525 3.8 ;
      RECT 86.475 2.175 86.575 3.8 ;
      RECT 86.225 2.175 86.325 3.8 ;
      RECT 85.275 2.175 85.375 3.8 ;
      RECT 85.025 2.175 85.125 3.8 ;
      RECT 84.075 2.175 84.175 3.8 ;
      RECT 83.825 2.175 83.925 3.8 ;
      RECT 82.875 2.175 82.975 3.8 ;
      RECT 82.625 2.175 82.725 3.8 ;
      RECT 81.675 2.175 81.775 3.8 ;
      RECT 81.425 2.175 81.525 3.8 ;
      RECT 80.475 2.175 80.575 3.8 ;
      RECT 80.225 2.175 80.325 3.8 ;
      RECT 79.275 2.175 79.375 3.8 ;
      RECT 79.025 2.175 79.125 3.8 ;
      RECT 78.075 2.175 78.175 3.8 ;
      RECT 77.825 2.175 77.925 3.8 ;
      RECT 76.875 2.175 76.975 3.8 ;
      RECT 76.625 2.175 76.725 3.8 ;
      RECT 75.675 2.175 75.775 3.8 ;
      RECT 75.425 2.175 75.525 3.8 ;
      RECT 74.475 2.175 74.575 3.8 ;
      RECT 74.225 2.175 74.325 3.8 ;
      RECT 73.275 2.175 73.375 3.8 ;
      RECT 73.025 2.175 73.125 3.8 ;
      RECT 72.075 2.175 72.175 3.8 ;
      RECT 71.825 2.175 71.925 3.8 ;
      RECT 70.875 2.175 70.975 3.8 ;
      RECT 70.625 2.175 70.725 3.8 ;
      RECT 69.675 2.175 69.775 3.8 ;
      RECT 69.425 2.175 69.525 3.8 ;
      RECT 68.475 2.175 68.575 3.8 ;
      RECT 68.225 2.175 68.325 3.8 ;
      RECT 67.275 2.175 67.375 3.8 ;
      RECT 67.025 2.175 67.125 3.8 ;
      RECT 66.075 2.175 66.175 3.8 ;
      RECT 65.825 2.175 65.925 3.8 ;
      RECT 64.875 2.175 64.975 3.8 ;
      RECT 64.625 2.175 64.725 3.8 ;
      RECT 63.675 2.175 63.775 3.8 ;
      RECT 63.425 2.175 63.525 3.8 ;
      RECT 62.475 2.175 62.575 3.8 ;
      RECT 62.225 2.175 62.325 3.8 ;
      RECT 61.275 2.175 61.375 3.8 ;
      RECT 61.025 2.175 61.125 3.8 ;
      RECT 60.075 2.175 60.175 3.8 ;
      RECT 59.825 2.175 59.925 3.8 ;
      RECT 58.875 2.175 58.975 3.8 ;
      RECT 58.625 2.175 58.725 3.8 ;
      RECT 57.675 2.175 57.775 3.8 ;
      RECT 57.425 2.175 57.525 3.8 ;
      RECT 56.475 2.175 56.575 3.8 ;
      RECT 56.225 2.175 56.325 3.8 ;
      RECT 55.275 2.175 55.375 3.8 ;
      RECT 55.025 2.175 55.125 3.8 ;
      RECT 54.075 2.175 54.175 3.8 ;
      RECT 53.825 2.175 53.925 3.8 ;
      RECT 52.875 2.175 52.975 3.8 ;
      RECT 52.625 2.175 52.725 3.8 ;
      RECT 51.675 2.175 51.775 3.8 ;
      RECT 51.425 2.175 51.525 3.8 ;
      RECT 50.475 2.175 50.575 3.8 ;
      RECT 50.225 2.175 50.325 3.8 ;
      RECT 49.275 2.175 49.375 3.8 ;
      RECT 49.025 2.175 49.125 3.8 ;
      RECT 48.075 2.175 48.175 3.8 ;
      RECT 47.825 2.175 47.925 3.8 ;
      RECT 46.875 2.175 46.975 3.8 ;
      RECT 46.625 2.175 46.725 3.8 ;
      RECT 45.675 2.175 45.775 3.8 ;
      RECT 45.425 2.175 45.525 3.8 ;
      RECT 44.475 2.175 44.575 3.8 ;
      RECT 44.225 2.175 44.325 3.8 ;
      RECT 43.275 2.175 43.375 3.8 ;
      RECT 43.025 2.175 43.125 3.8 ;
      RECT 42.075 2.175 42.175 3.8 ;
      RECT 41.825 2.175 41.925 3.8 ;
      RECT 40.875 2.175 40.975 3.8 ;
      RECT 40.625 2.175 40.725 3.8 ;
      RECT 39.675 2.175 39.775 3.8 ;
      RECT 39.425 2.175 39.525 3.8 ;
      RECT 38.475 2.175 38.575 3.8 ;
      RECT 38.225 2.175 38.325 3.8 ;
      RECT 37.275 2.175 37.375 3.8 ;
      RECT 37.025 2.175 37.125 3.8 ;
      RECT 36.075 2.175 36.175 3.8 ;
      RECT 35.825 2.175 35.925 3.8 ;
      RECT 34.875 2.175 34.975 3.8 ;
      RECT 34.625 2.175 34.725 3.8 ;
      RECT 33.675 2.175 33.775 3.8 ;
      RECT 33.425 2.175 33.525 3.8 ;
      RECT 32.475 2.175 32.575 3.8 ;
      RECT 32.225 2.175 32.325 3.8 ;
      RECT 31.275 2.175 31.375 3.8 ;
      RECT 31.025 2.175 31.125 3.8 ;
      RECT 30.075 2.175 30.175 3.8 ;
      RECT 29.825 2.175 29.925 3.8 ;
      RECT 28.875 2.175 28.975 3.8 ;
      RECT 28.625 2.175 28.725 3.8 ;
      RECT 27.675 2.175 27.775 3.8 ;
      RECT 27.425 2.175 27.525 3.8 ;
      RECT 26.475 2.175 26.575 3.8 ;
      RECT 26.225 2.175 26.325 3.8 ;
      RECT 25.275 2.175 25.375 3.8 ;
      RECT 25.025 2.175 25.125 3.8 ;
      RECT 24.075 2.175 24.175 3.8 ;
      RECT 23.825 2.175 23.925 3.8 ;
      RECT 22.875 2.175 22.975 3.8 ;
      RECT 22.625 2.175 22.725 3.8 ;
      RECT 21.675 2.175 21.775 3.8 ;
      RECT 21.425 2.175 21.525 3.8 ;
      RECT 20.475 2.175 20.575 3.8 ;
      RECT 20.225 2.175 20.325 3.8 ;
      RECT 19.275 2.175 19.375 3.8 ;
      RECT 19.025 2.175 19.125 3.8 ;
      RECT 18.075 2.175 18.175 3.8 ;
      RECT 17.825 2.175 17.925 3.8 ;
      RECT 16.875 2.175 16.975 3.8 ;
      RECT 16.625 2.175 16.725 3.8 ;
      RECT 15.675 2.175 15.775 3.8 ;
      RECT 15.425 2.175 15.525 3.8 ;
      RECT 14.475 2.175 14.575 3.8 ;
      RECT 14.225 2.175 14.325 3.8 ;
      RECT 13.275 2.175 13.375 3.8 ;
      RECT 13.025 2.175 13.125 3.8 ;
      RECT 12.075 2.175 12.175 3.8 ;
      RECT 11.825 2.175 11.925 3.8 ;
      RECT 10.875 2.175 10.975 3.8 ;
      RECT 10.625 2.175 10.725 3.8 ;
      RECT 9.675 2.175 9.775 3.8 ;
      RECT 9.425 2.175 9.525 3.8 ;
      RECT 8.475 2.175 8.575 3.8 ;
      RECT 8.225 2.175 8.325 3.8 ;
      RECT 7.275 2.175 7.375 3.8 ;
      RECT 7.025 2.175 7.125 3.8 ;
      RECT 6.075 2.175 6.175 3.8 ;
      RECT 5.825 2.175 5.925 3.8 ;
      RECT 4.875 2.175 4.975 3.8 ;
      RECT 4.625 2.175 4.725 3.8 ;
      RECT 3.675 2.175 3.775 3.8 ;
      RECT 3.425 2.175 3.525 3.8 ;
      RECT 2.475 2.175 2.575 3.8 ;
      RECT 2.225 2.175 2.325 3.8 ;
      RECT 1.275 2.175 1.375 3.8 ;
      RECT 1.025 2.175 1.125 3.8 ;
      RECT 0.075 2.175 0.175 3.8 ;
      RECT -39.505 7.175 155.517 9.895 ;
      RECT -6.66 4.965 -5.425 9.895 ;
      RECT -6.065 4.385 -5.965 9.895 ;
      RECT -4.885 -100.48 -4.705 -100.3 ;
      RECT -4.885 -100.435 153.65 -100.345 ;
      RECT -3.585 -99.96 -3.405 -99.78 ;
      RECT -3.585 -99.915 153.65 -99.825 ;
      RECT -2.285 -97.25 -2.105 -97.07 ;
      RECT -2.285 -97.205 153.65 -97.115 ;
      RECT -0.985 -96.73 -0.805 -96.55 ;
      RECT -0.985 -96.685 153.65 -96.595 ;
      RECT -0.985 -94.02 -0.805 -93.84 ;
      RECT -0.985 -93.975 153.65 -93.885 ;
      RECT -2.285 -93.5 -2.105 -93.32 ;
      RECT -2.285 -93.455 153.65 -93.365 ;
      RECT -3.585 -90.79 -3.405 -90.61 ;
      RECT -3.585 -90.745 153.65 -90.655 ;
      RECT -4.885 -90.27 -4.705 -90.09 ;
      RECT -4.885 -90.225 153.65 -90.135 ;
      RECT -4.885 -87.56 -4.705 -87.38 ;
      RECT -4.885 -87.515 153.65 -87.425 ;
      RECT -3.585 -87.04 -3.405 -86.86 ;
      RECT -3.585 -86.995 153.65 -86.905 ;
      RECT -2.285 -84.33 -2.105 -84.15 ;
      RECT -2.285 -84.285 153.65 -84.195 ;
      RECT -0.985 -83.81 -0.805 -83.63 ;
      RECT -0.985 -83.765 153.65 -83.675 ;
      RECT -0.985 -81.1 -0.805 -80.92 ;
      RECT -0.985 -81.055 153.65 -80.965 ;
      RECT -2.285 -80.58 -2.105 -80.4 ;
      RECT -2.285 -80.535 153.65 -80.445 ;
      RECT -3.585 -77.87 -3.405 -77.69 ;
      RECT -3.585 -77.825 153.65 -77.735 ;
      RECT -4.885 -77.35 -4.705 -77.17 ;
      RECT -4.885 -77.305 153.65 -77.215 ;
      RECT -4.885 -74.64 -4.705 -74.46 ;
      RECT -4.885 -74.595 153.65 -74.505 ;
      RECT -3.585 -74.12 -3.405 -73.94 ;
      RECT -3.585 -74.075 153.65 -73.985 ;
      RECT -2.285 -71.41 -2.105 -71.23 ;
      RECT -2.285 -71.365 153.65 -71.275 ;
      RECT -0.985 -70.89 -0.805 -70.71 ;
      RECT -0.985 -70.845 153.65 -70.755 ;
      RECT -0.985 -68.18 -0.805 -68 ;
      RECT -0.985 -68.135 153.65 -68.045 ;
      RECT -2.285 -67.66 -2.105 -67.48 ;
      RECT -2.285 -67.615 153.65 -67.525 ;
      RECT -3.585 -64.95 -3.405 -64.77 ;
      RECT -3.585 -64.905 153.65 -64.815 ;
      RECT -4.885 -64.43 -4.705 -64.25 ;
      RECT -4.885 -64.385 153.65 -64.295 ;
      RECT -4.885 -61.72 -4.705 -61.54 ;
      RECT -4.885 -61.675 153.65 -61.585 ;
      RECT -3.585 -61.2 -3.405 -61.02 ;
      RECT -3.585 -61.155 153.65 -61.065 ;
      RECT -2.285 -58.49 -2.105 -58.31 ;
      RECT -2.285 -58.445 153.65 -58.355 ;
      RECT -0.985 -57.97 -0.805 -57.79 ;
      RECT -0.985 -57.925 153.65 -57.835 ;
      RECT -0.985 -55.26 -0.805 -55.08 ;
      RECT -0.985 -55.215 153.65 -55.125 ;
      RECT -2.285 -54.74 -2.105 -54.56 ;
      RECT -2.285 -54.695 153.65 -54.605 ;
      RECT -3.585 -52.03 -3.405 -51.85 ;
      RECT -3.585 -51.985 153.65 -51.895 ;
      RECT -4.885 -51.51 -4.705 -51.33 ;
      RECT -4.885 -51.465 153.65 -51.375 ;
      RECT -4.885 -48.8 -4.705 -48.62 ;
      RECT -4.885 -48.755 153.65 -48.665 ;
      RECT -3.585 -48.28 -3.405 -48.1 ;
      RECT -3.585 -48.235 153.65 -48.145 ;
      RECT -2.285 -45.57 -2.105 -45.39 ;
      RECT -2.285 -45.525 153.65 -45.435 ;
      RECT -0.985 -45.05 -0.805 -44.87 ;
      RECT -0.985 -45.005 153.65 -44.915 ;
      RECT -0.985 -42.34 -0.805 -42.16 ;
      RECT -0.985 -42.295 153.65 -42.205 ;
      RECT -2.285 -41.82 -2.105 -41.64 ;
      RECT -2.285 -41.775 153.65 -41.685 ;
      RECT -3.585 -39.11 -3.405 -38.93 ;
      RECT -3.585 -39.065 153.65 -38.975 ;
      RECT -4.885 -38.59 -4.705 -38.41 ;
      RECT -4.885 -38.545 153.65 -38.455 ;
      RECT -4.885 -35.88 -4.705 -35.7 ;
      RECT -4.885 -35.835 153.65 -35.745 ;
      RECT -3.585 -35.36 -3.405 -35.18 ;
      RECT -3.585 -35.315 153.65 -35.225 ;
      RECT -2.285 -32.65 -2.105 -32.47 ;
      RECT -2.285 -32.605 153.65 -32.515 ;
      RECT -0.985 -32.13 -0.805 -31.95 ;
      RECT -0.985 -32.085 153.65 -31.995 ;
      RECT -0.985 -29.42 -0.805 -29.24 ;
      RECT -0.985 -29.375 153.65 -29.285 ;
      RECT -2.285 -28.9 -2.105 -28.72 ;
      RECT -2.285 -28.855 153.65 -28.765 ;
      RECT -3.585 -26.19 -3.405 -26.01 ;
      RECT -3.585 -26.145 153.65 -26.055 ;
      RECT -4.885 -25.67 -4.705 -25.49 ;
      RECT -4.885 -25.625 153.65 -25.535 ;
      RECT -4.885 -22.96 -4.705 -22.78 ;
      RECT -4.885 -22.915 153.65 -22.825 ;
      RECT -3.585 -22.44 -3.405 -22.26 ;
      RECT -3.585 -22.395 153.65 -22.305 ;
      RECT -2.285 -19.73 -2.105 -19.55 ;
      RECT -2.285 -19.685 153.65 -19.595 ;
      RECT -0.985 -19.21 -0.805 -19.03 ;
      RECT -0.985 -19.165 153.65 -19.075 ;
      RECT -0.985 -16.5 -0.805 -16.32 ;
      RECT -0.985 -16.455 153.65 -16.365 ;
      RECT -2.285 -15.98 -2.105 -15.8 ;
      RECT -2.285 -15.935 153.65 -15.845 ;
      RECT -3.585 -13.27 -3.405 -13.09 ;
      RECT -3.585 -13.225 153.65 -13.135 ;
      RECT -4.885 -12.75 -4.705 -12.57 ;
      RECT -4.885 -12.705 153.65 -12.615 ;
      RECT -4.885 -10.04 -4.705 -9.86 ;
      RECT -4.885 -9.995 153.65 -9.905 ;
      RECT -3.585 -9.52 -3.405 -9.34 ;
      RECT -3.585 -9.475 153.65 -9.385 ;
      RECT -2.285 -6.81 -2.105 -6.63 ;
      RECT -2.285 -6.765 153.65 -6.675 ;
      RECT -0.985 -6.29 -0.805 -6.11 ;
      RECT -0.985 -6.245 153.65 -6.155 ;
      RECT -0.985 -3.58 -0.805 -3.4 ;
      RECT -0.985 -3.535 153.65 -3.445 ;
      RECT -2.285 -3.06 -2.105 -2.88 ;
      RECT -2.285 -3.015 153.65 -2.925 ;
      RECT -3.585 -0.35 -3.405 -0.17 ;
      RECT -3.585 -0.305 153.65 -0.215 ;
      RECT -4.885 0.17 -4.705 0.35 ;
      RECT -4.885 0.215 153.65 0.305 ;
      RECT 149.785 -108.935 153.565 -108.815 ;
      RECT 151.105 -109.475 151.205 -108.815 ;
      RECT 150.545 -109.475 150.645 -108.815 ;
      RECT 149.985 -109.475 150.085 -108.815 ;
      RECT -4.885 -103.19 -4.705 -103.01 ;
      RECT -4.885 -103.145 153.43 -103.055 ;
      RECT 153.155 -101.538 153.245 -100.53 ;
      RECT 153.105 -100.935 153.245 -100.765 ;
      RECT 153.155 -99.73 153.245 -98.722 ;
      RECT 153.105 -99.495 153.245 -99.325 ;
      RECT 153.155 -98.308 153.245 -97.3 ;
      RECT 153.105 -97.705 153.245 -97.535 ;
      RECT 153.155 -96.5 153.245 -95.492 ;
      RECT 153.105 -96.265 153.245 -96.095 ;
      RECT 153.155 -95.078 153.245 -94.07 ;
      RECT 153.105 -94.475 153.245 -94.305 ;
      RECT 153.155 -93.27 153.245 -92.262 ;
      RECT 153.105 -93.035 153.245 -92.865 ;
      RECT 153.155 -91.848 153.245 -90.84 ;
      RECT 153.105 -91.245 153.245 -91.075 ;
      RECT 153.155 -90.04 153.245 -89.032 ;
      RECT 153.105 -89.805 153.245 -89.635 ;
      RECT 153.155 -88.618 153.245 -87.61 ;
      RECT 153.105 -88.015 153.245 -87.845 ;
      RECT 153.155 -86.81 153.245 -85.802 ;
      RECT 153.105 -86.575 153.245 -86.405 ;
      RECT 153.155 -85.388 153.245 -84.38 ;
      RECT 153.105 -84.785 153.245 -84.615 ;
      RECT 153.155 -83.58 153.245 -82.572 ;
      RECT 153.105 -83.345 153.245 -83.175 ;
      RECT 153.155 -82.158 153.245 -81.15 ;
      RECT 153.105 -81.555 153.245 -81.385 ;
      RECT 153.155 -80.35 153.245 -79.342 ;
      RECT 153.105 -80.115 153.245 -79.945 ;
      RECT 153.155 -78.928 153.245 -77.92 ;
      RECT 153.105 -78.325 153.245 -78.155 ;
      RECT 153.155 -77.12 153.245 -76.112 ;
      RECT 153.105 -76.885 153.245 -76.715 ;
      RECT 153.155 -75.698 153.245 -74.69 ;
      RECT 153.105 -75.095 153.245 -74.925 ;
      RECT 153.155 -73.89 153.245 -72.882 ;
      RECT 153.105 -73.655 153.245 -73.485 ;
      RECT 153.155 -72.468 153.245 -71.46 ;
      RECT 153.105 -71.865 153.245 -71.695 ;
      RECT 153.155 -70.66 153.245 -69.652 ;
      RECT 153.105 -70.425 153.245 -70.255 ;
      RECT 153.155 -69.238 153.245 -68.23 ;
      RECT 153.105 -68.635 153.245 -68.465 ;
      RECT 153.155 -67.43 153.245 -66.422 ;
      RECT 153.105 -67.195 153.245 -67.025 ;
      RECT 153.155 -66.008 153.245 -65 ;
      RECT 153.105 -65.405 153.245 -65.235 ;
      RECT 153.155 -64.2 153.245 -63.192 ;
      RECT 153.105 -63.965 153.245 -63.795 ;
      RECT 153.155 -62.778 153.245 -61.77 ;
      RECT 153.105 -62.175 153.245 -62.005 ;
      RECT 153.155 -60.97 153.245 -59.962 ;
      RECT 153.105 -60.735 153.245 -60.565 ;
      RECT 153.155 -59.548 153.245 -58.54 ;
      RECT 153.105 -58.945 153.245 -58.775 ;
      RECT 153.155 -57.74 153.245 -56.732 ;
      RECT 153.105 -57.505 153.245 -57.335 ;
      RECT 153.155 -56.318 153.245 -55.31 ;
      RECT 153.105 -55.715 153.245 -55.545 ;
      RECT 153.155 -54.51 153.245 -53.502 ;
      RECT 153.105 -54.275 153.245 -54.105 ;
      RECT 153.155 -53.088 153.245 -52.08 ;
      RECT 153.105 -52.485 153.245 -52.315 ;
      RECT 153.155 -51.28 153.245 -50.272 ;
      RECT 153.105 -51.045 153.245 -50.875 ;
      RECT 153.155 -49.858 153.245 -48.85 ;
      RECT 153.105 -49.255 153.245 -49.085 ;
      RECT 153.155 -48.05 153.245 -47.042 ;
      RECT 153.105 -47.815 153.245 -47.645 ;
      RECT 153.155 -46.628 153.245 -45.62 ;
      RECT 153.105 -46.025 153.245 -45.855 ;
      RECT 153.155 -44.82 153.245 -43.812 ;
      RECT 153.105 -44.585 153.245 -44.415 ;
      RECT 153.155 -43.398 153.245 -42.39 ;
      RECT 153.105 -42.795 153.245 -42.625 ;
      RECT 153.155 -41.59 153.245 -40.582 ;
      RECT 153.105 -41.355 153.245 -41.185 ;
      RECT 153.155 -40.168 153.245 -39.16 ;
      RECT 153.105 -39.565 153.245 -39.395 ;
      RECT 153.155 -38.36 153.245 -37.352 ;
      RECT 153.105 -38.125 153.245 -37.955 ;
      RECT 153.155 -36.938 153.245 -35.93 ;
      RECT 153.105 -36.335 153.245 -36.165 ;
      RECT 153.155 -35.13 153.245 -34.122 ;
      RECT 153.105 -34.895 153.245 -34.725 ;
      RECT 153.155 -33.708 153.245 -32.7 ;
      RECT 153.105 -33.105 153.245 -32.935 ;
      RECT 153.155 -31.9 153.245 -30.892 ;
      RECT 153.105 -31.665 153.245 -31.495 ;
      RECT 153.155 -30.478 153.245 -29.47 ;
      RECT 153.105 -29.875 153.245 -29.705 ;
      RECT 153.155 -28.67 153.245 -27.662 ;
      RECT 153.105 -28.435 153.245 -28.265 ;
      RECT 153.155 -27.248 153.245 -26.24 ;
      RECT 153.105 -26.645 153.245 -26.475 ;
      RECT 153.155 -25.44 153.245 -24.432 ;
      RECT 153.105 -25.205 153.245 -25.035 ;
      RECT 153.155 -24.018 153.245 -23.01 ;
      RECT 153.105 -23.415 153.245 -23.245 ;
      RECT 153.155 -22.21 153.245 -21.202 ;
      RECT 153.105 -21.975 153.245 -21.805 ;
      RECT 153.155 -20.788 153.245 -19.78 ;
      RECT 153.105 -20.185 153.245 -20.015 ;
      RECT 153.155 -18.98 153.245 -17.972 ;
      RECT 153.105 -18.745 153.245 -18.575 ;
      RECT 153.155 -17.558 153.245 -16.55 ;
      RECT 153.105 -16.955 153.245 -16.785 ;
      RECT 153.155 -15.75 153.245 -14.742 ;
      RECT 153.105 -15.515 153.245 -15.345 ;
      RECT 153.155 -14.328 153.245 -13.32 ;
      RECT 153.105 -13.725 153.245 -13.555 ;
      RECT 153.155 -12.52 153.245 -11.512 ;
      RECT 153.105 -12.285 153.245 -12.115 ;
      RECT 153.155 -11.098 153.245 -10.09 ;
      RECT 153.105 -10.495 153.245 -10.325 ;
      RECT 153.155 -9.29 153.245 -8.282 ;
      RECT 153.105 -9.055 153.245 -8.885 ;
      RECT 153.155 -7.868 153.245 -6.86 ;
      RECT 153.105 -7.265 153.245 -7.095 ;
      RECT 153.155 -6.06 153.245 -5.052 ;
      RECT 153.105 -5.825 153.245 -5.655 ;
      RECT 153.155 -4.638 153.245 -3.63 ;
      RECT 153.105 -4.035 153.245 -3.865 ;
      RECT 153.155 -2.83 153.245 -1.822 ;
      RECT 153.105 -2.595 153.245 -2.425 ;
      RECT 153.155 -1.408 153.245 -0.4 ;
      RECT 153.105 -0.805 153.245 -0.635 ;
      RECT 153.155 0.4 153.245 1.408 ;
      RECT 153.105 0.635 153.245 0.805 ;
      RECT 151.725 -111.685 153.205 -111.585 ;
      RECT 151.725 -112.195 151.825 -111.585 ;
      RECT 151.945 -109.15 153.205 -109.05 ;
      RECT 153.105 -109.475 153.205 -109.05 ;
      RECT 152.545 -109.475 152.645 -109.05 ;
      RECT 151.985 -109.475 152.085 -109.05 ;
      RECT 152.755 -101.538 152.845 -100.531 ;
      RECT 152.755 -101.225 152.895 -101.055 ;
      RECT 152.755 -99.729 152.845 -98.722 ;
      RECT 152.755 -99.205 152.895 -99.035 ;
      RECT 152.755 -98.308 152.845 -97.301 ;
      RECT 152.755 -97.995 152.895 -97.825 ;
      RECT 152.755 -96.499 152.845 -95.492 ;
      RECT 152.755 -95.975 152.895 -95.805 ;
      RECT 152.755 -95.078 152.845 -94.071 ;
      RECT 152.755 -94.765 152.895 -94.595 ;
      RECT 152.755 -93.269 152.845 -92.262 ;
      RECT 152.755 -92.745 152.895 -92.575 ;
      RECT 152.755 -91.848 152.845 -90.841 ;
      RECT 152.755 -91.535 152.895 -91.365 ;
      RECT 152.755 -90.039 152.845 -89.032 ;
      RECT 152.755 -89.515 152.895 -89.345 ;
      RECT 152.755 -88.618 152.845 -87.611 ;
      RECT 152.755 -88.305 152.895 -88.135 ;
      RECT 152.755 -86.809 152.845 -85.802 ;
      RECT 152.755 -86.285 152.895 -86.115 ;
      RECT 152.755 -85.388 152.845 -84.381 ;
      RECT 152.755 -85.075 152.895 -84.905 ;
      RECT 152.755 -83.579 152.845 -82.572 ;
      RECT 152.755 -83.055 152.895 -82.885 ;
      RECT 152.755 -82.158 152.845 -81.151 ;
      RECT 152.755 -81.845 152.895 -81.675 ;
      RECT 152.755 -80.349 152.845 -79.342 ;
      RECT 152.755 -79.825 152.895 -79.655 ;
      RECT 152.755 -78.928 152.845 -77.921 ;
      RECT 152.755 -78.615 152.895 -78.445 ;
      RECT 152.755 -77.119 152.845 -76.112 ;
      RECT 152.755 -76.595 152.895 -76.425 ;
      RECT 152.755 -75.698 152.845 -74.691 ;
      RECT 152.755 -75.385 152.895 -75.215 ;
      RECT 152.755 -73.889 152.845 -72.882 ;
      RECT 152.755 -73.365 152.895 -73.195 ;
      RECT 152.755 -72.468 152.845 -71.461 ;
      RECT 152.755 -72.155 152.895 -71.985 ;
      RECT 152.755 -70.659 152.845 -69.652 ;
      RECT 152.755 -70.135 152.895 -69.965 ;
      RECT 152.755 -69.238 152.845 -68.231 ;
      RECT 152.755 -68.925 152.895 -68.755 ;
      RECT 152.755 -67.429 152.845 -66.422 ;
      RECT 152.755 -66.905 152.895 -66.735 ;
      RECT 152.755 -66.008 152.845 -65.001 ;
      RECT 152.755 -65.695 152.895 -65.525 ;
      RECT 152.755 -64.199 152.845 -63.192 ;
      RECT 152.755 -63.675 152.895 -63.505 ;
      RECT 152.755 -62.778 152.845 -61.771 ;
      RECT 152.755 -62.465 152.895 -62.295 ;
      RECT 152.755 -60.969 152.845 -59.962 ;
      RECT 152.755 -60.445 152.895 -60.275 ;
      RECT 152.755 -59.548 152.845 -58.541 ;
      RECT 152.755 -59.235 152.895 -59.065 ;
      RECT 152.755 -57.739 152.845 -56.732 ;
      RECT 152.755 -57.215 152.895 -57.045 ;
      RECT 152.755 -56.318 152.845 -55.311 ;
      RECT 152.755 -56.005 152.895 -55.835 ;
      RECT 152.755 -54.509 152.845 -53.502 ;
      RECT 152.755 -53.985 152.895 -53.815 ;
      RECT 152.755 -53.088 152.845 -52.081 ;
      RECT 152.755 -52.775 152.895 -52.605 ;
      RECT 152.755 -51.279 152.845 -50.272 ;
      RECT 152.755 -50.755 152.895 -50.585 ;
      RECT 152.755 -49.858 152.845 -48.851 ;
      RECT 152.755 -49.545 152.895 -49.375 ;
      RECT 152.755 -48.049 152.845 -47.042 ;
      RECT 152.755 -47.525 152.895 -47.355 ;
      RECT 152.755 -46.628 152.845 -45.621 ;
      RECT 152.755 -46.315 152.895 -46.145 ;
      RECT 152.755 -44.819 152.845 -43.812 ;
      RECT 152.755 -44.295 152.895 -44.125 ;
      RECT 152.755 -43.398 152.845 -42.391 ;
      RECT 152.755 -43.085 152.895 -42.915 ;
      RECT 152.755 -41.589 152.845 -40.582 ;
      RECT 152.755 -41.065 152.895 -40.895 ;
      RECT 152.755 -40.168 152.845 -39.161 ;
      RECT 152.755 -39.855 152.895 -39.685 ;
      RECT 152.755 -38.359 152.845 -37.352 ;
      RECT 152.755 -37.835 152.895 -37.665 ;
      RECT 152.755 -36.938 152.845 -35.931 ;
      RECT 152.755 -36.625 152.895 -36.455 ;
      RECT 152.755 -35.129 152.845 -34.122 ;
      RECT 152.755 -34.605 152.895 -34.435 ;
      RECT 152.755 -33.708 152.845 -32.701 ;
      RECT 152.755 -33.395 152.895 -33.225 ;
      RECT 152.755 -31.899 152.845 -30.892 ;
      RECT 152.755 -31.375 152.895 -31.205 ;
      RECT 152.755 -30.478 152.845 -29.471 ;
      RECT 152.755 -30.165 152.895 -29.995 ;
      RECT 152.755 -28.669 152.845 -27.662 ;
      RECT 152.755 -28.145 152.895 -27.975 ;
      RECT 152.755 -27.248 152.845 -26.241 ;
      RECT 152.755 -26.935 152.895 -26.765 ;
      RECT 152.755 -25.439 152.845 -24.432 ;
      RECT 152.755 -24.915 152.895 -24.745 ;
      RECT 152.755 -24.018 152.845 -23.011 ;
      RECT 152.755 -23.705 152.895 -23.535 ;
      RECT 152.755 -22.209 152.845 -21.202 ;
      RECT 152.755 -21.685 152.895 -21.515 ;
      RECT 152.755 -20.788 152.845 -19.781 ;
      RECT 152.755 -20.475 152.895 -20.305 ;
      RECT 152.755 -18.979 152.845 -17.972 ;
      RECT 152.755 -18.455 152.895 -18.285 ;
      RECT 152.755 -17.558 152.845 -16.551 ;
      RECT 152.755 -17.245 152.895 -17.075 ;
      RECT 152.755 -15.749 152.845 -14.742 ;
      RECT 152.755 -15.225 152.895 -15.055 ;
      RECT 152.755 -14.328 152.845 -13.321 ;
      RECT 152.755 -14.015 152.895 -13.845 ;
      RECT 152.755 -12.519 152.845 -11.512 ;
      RECT 152.755 -11.995 152.895 -11.825 ;
      RECT 152.755 -11.098 152.845 -10.091 ;
      RECT 152.755 -10.785 152.895 -10.615 ;
      RECT 152.755 -9.289 152.845 -8.282 ;
      RECT 152.755 -8.765 152.895 -8.595 ;
      RECT 152.755 -7.868 152.845 -6.861 ;
      RECT 152.755 -7.555 152.895 -7.385 ;
      RECT 152.755 -6.059 152.845 -5.052 ;
      RECT 152.755 -5.535 152.895 -5.365 ;
      RECT 152.755 -4.638 152.845 -3.631 ;
      RECT 152.755 -4.325 152.895 -4.155 ;
      RECT 152.755 -2.829 152.845 -1.822 ;
      RECT 152.755 -2.305 152.895 -2.135 ;
      RECT 152.755 -1.408 152.845 -0.401 ;
      RECT 152.755 -1.095 152.895 -0.925 ;
      RECT 152.755 0.401 152.845 1.408 ;
      RECT 152.755 0.925 152.895 1.095 ;
      RECT 152.085 -111.495 152.255 -111.385 ;
      RECT 148.935 -111.495 152.255 -111.395 ;
      RECT -3.585 -103.71 -3.405 -103.53 ;
      RECT -3.585 -103.665 152.23 -103.575 ;
      RECT 151.955 -101.538 152.045 -100.53 ;
      RECT 151.905 -100.935 152.045 -100.765 ;
      RECT 151.955 -99.73 152.045 -98.722 ;
      RECT 151.905 -99.495 152.045 -99.325 ;
      RECT 151.955 -98.308 152.045 -97.3 ;
      RECT 151.905 -97.705 152.045 -97.535 ;
      RECT 151.955 -96.5 152.045 -95.492 ;
      RECT 151.905 -96.265 152.045 -96.095 ;
      RECT 151.955 -95.078 152.045 -94.07 ;
      RECT 151.905 -94.475 152.045 -94.305 ;
      RECT 151.955 -93.27 152.045 -92.262 ;
      RECT 151.905 -93.035 152.045 -92.865 ;
      RECT 151.955 -91.848 152.045 -90.84 ;
      RECT 151.905 -91.245 152.045 -91.075 ;
      RECT 151.955 -90.04 152.045 -89.032 ;
      RECT 151.905 -89.805 152.045 -89.635 ;
      RECT 151.955 -88.618 152.045 -87.61 ;
      RECT 151.905 -88.015 152.045 -87.845 ;
      RECT 151.955 -86.81 152.045 -85.802 ;
      RECT 151.905 -86.575 152.045 -86.405 ;
      RECT 151.955 -85.388 152.045 -84.38 ;
      RECT 151.905 -84.785 152.045 -84.615 ;
      RECT 151.955 -83.58 152.045 -82.572 ;
      RECT 151.905 -83.345 152.045 -83.175 ;
      RECT 151.955 -82.158 152.045 -81.15 ;
      RECT 151.905 -81.555 152.045 -81.385 ;
      RECT 151.955 -80.35 152.045 -79.342 ;
      RECT 151.905 -80.115 152.045 -79.945 ;
      RECT 151.955 -78.928 152.045 -77.92 ;
      RECT 151.905 -78.325 152.045 -78.155 ;
      RECT 151.955 -77.12 152.045 -76.112 ;
      RECT 151.905 -76.885 152.045 -76.715 ;
      RECT 151.955 -75.698 152.045 -74.69 ;
      RECT 151.905 -75.095 152.045 -74.925 ;
      RECT 151.955 -73.89 152.045 -72.882 ;
      RECT 151.905 -73.655 152.045 -73.485 ;
      RECT 151.955 -72.468 152.045 -71.46 ;
      RECT 151.905 -71.865 152.045 -71.695 ;
      RECT 151.955 -70.66 152.045 -69.652 ;
      RECT 151.905 -70.425 152.045 -70.255 ;
      RECT 151.955 -69.238 152.045 -68.23 ;
      RECT 151.905 -68.635 152.045 -68.465 ;
      RECT 151.955 -67.43 152.045 -66.422 ;
      RECT 151.905 -67.195 152.045 -67.025 ;
      RECT 151.955 -66.008 152.045 -65 ;
      RECT 151.905 -65.405 152.045 -65.235 ;
      RECT 151.955 -64.2 152.045 -63.192 ;
      RECT 151.905 -63.965 152.045 -63.795 ;
      RECT 151.955 -62.778 152.045 -61.77 ;
      RECT 151.905 -62.175 152.045 -62.005 ;
      RECT 151.955 -60.97 152.045 -59.962 ;
      RECT 151.905 -60.735 152.045 -60.565 ;
      RECT 151.955 -59.548 152.045 -58.54 ;
      RECT 151.905 -58.945 152.045 -58.775 ;
      RECT 151.955 -57.74 152.045 -56.732 ;
      RECT 151.905 -57.505 152.045 -57.335 ;
      RECT 151.955 -56.318 152.045 -55.31 ;
      RECT 151.905 -55.715 152.045 -55.545 ;
      RECT 151.955 -54.51 152.045 -53.502 ;
      RECT 151.905 -54.275 152.045 -54.105 ;
      RECT 151.955 -53.088 152.045 -52.08 ;
      RECT 151.905 -52.485 152.045 -52.315 ;
      RECT 151.955 -51.28 152.045 -50.272 ;
      RECT 151.905 -51.045 152.045 -50.875 ;
      RECT 151.955 -49.858 152.045 -48.85 ;
      RECT 151.905 -49.255 152.045 -49.085 ;
      RECT 151.955 -48.05 152.045 -47.042 ;
      RECT 151.905 -47.815 152.045 -47.645 ;
      RECT 151.955 -46.628 152.045 -45.62 ;
      RECT 151.905 -46.025 152.045 -45.855 ;
      RECT 151.955 -44.82 152.045 -43.812 ;
      RECT 151.905 -44.585 152.045 -44.415 ;
      RECT 151.955 -43.398 152.045 -42.39 ;
      RECT 151.905 -42.795 152.045 -42.625 ;
      RECT 151.955 -41.59 152.045 -40.582 ;
      RECT 151.905 -41.355 152.045 -41.185 ;
      RECT 151.955 -40.168 152.045 -39.16 ;
      RECT 151.905 -39.565 152.045 -39.395 ;
      RECT 151.955 -38.36 152.045 -37.352 ;
      RECT 151.905 -38.125 152.045 -37.955 ;
      RECT 151.955 -36.938 152.045 -35.93 ;
      RECT 151.905 -36.335 152.045 -36.165 ;
      RECT 151.955 -35.13 152.045 -34.122 ;
      RECT 151.905 -34.895 152.045 -34.725 ;
      RECT 151.955 -33.708 152.045 -32.7 ;
      RECT 151.905 -33.105 152.045 -32.935 ;
      RECT 151.955 -31.9 152.045 -30.892 ;
      RECT 151.905 -31.665 152.045 -31.495 ;
      RECT 151.955 -30.478 152.045 -29.47 ;
      RECT 151.905 -29.875 152.045 -29.705 ;
      RECT 151.955 -28.67 152.045 -27.662 ;
      RECT 151.905 -28.435 152.045 -28.265 ;
      RECT 151.955 -27.248 152.045 -26.24 ;
      RECT 151.905 -26.645 152.045 -26.475 ;
      RECT 151.955 -25.44 152.045 -24.432 ;
      RECT 151.905 -25.205 152.045 -25.035 ;
      RECT 151.955 -24.018 152.045 -23.01 ;
      RECT 151.905 -23.415 152.045 -23.245 ;
      RECT 151.955 -22.21 152.045 -21.202 ;
      RECT 151.905 -21.975 152.045 -21.805 ;
      RECT 151.955 -20.788 152.045 -19.78 ;
      RECT 151.905 -20.185 152.045 -20.015 ;
      RECT 151.955 -18.98 152.045 -17.972 ;
      RECT 151.905 -18.745 152.045 -18.575 ;
      RECT 151.955 -17.558 152.045 -16.55 ;
      RECT 151.905 -16.955 152.045 -16.785 ;
      RECT 151.955 -15.75 152.045 -14.742 ;
      RECT 151.905 -15.515 152.045 -15.345 ;
      RECT 151.955 -14.328 152.045 -13.32 ;
      RECT 151.905 -13.725 152.045 -13.555 ;
      RECT 151.955 -12.52 152.045 -11.512 ;
      RECT 151.905 -12.285 152.045 -12.115 ;
      RECT 151.955 -11.098 152.045 -10.09 ;
      RECT 151.905 -10.495 152.045 -10.325 ;
      RECT 151.955 -9.29 152.045 -8.282 ;
      RECT 151.905 -9.055 152.045 -8.885 ;
      RECT 151.955 -7.868 152.045 -6.86 ;
      RECT 151.905 -7.265 152.045 -7.095 ;
      RECT 151.955 -6.06 152.045 -5.052 ;
      RECT 151.905 -5.825 152.045 -5.655 ;
      RECT 151.955 -4.638 152.045 -3.63 ;
      RECT 151.905 -4.035 152.045 -3.865 ;
      RECT 151.955 -2.83 152.045 -1.822 ;
      RECT 151.905 -2.595 152.045 -2.425 ;
      RECT 151.955 -1.408 152.045 -0.4 ;
      RECT 151.905 -0.805 152.045 -0.635 ;
      RECT 151.955 0.4 152.045 1.408 ;
      RECT 151.905 0.635 152.045 0.805 ;
      RECT 151.555 -101.538 151.645 -100.531 ;
      RECT 151.555 -101.225 151.695 -101.055 ;
      RECT 151.555 -99.729 151.645 -98.722 ;
      RECT 151.555 -99.205 151.695 -99.035 ;
      RECT 151.555 -98.308 151.645 -97.301 ;
      RECT 151.555 -97.995 151.695 -97.825 ;
      RECT 151.555 -96.499 151.645 -95.492 ;
      RECT 151.555 -95.975 151.695 -95.805 ;
      RECT 151.555 -95.078 151.645 -94.071 ;
      RECT 151.555 -94.765 151.695 -94.595 ;
      RECT 151.555 -93.269 151.645 -92.262 ;
      RECT 151.555 -92.745 151.695 -92.575 ;
      RECT 151.555 -91.848 151.645 -90.841 ;
      RECT 151.555 -91.535 151.695 -91.365 ;
      RECT 151.555 -90.039 151.645 -89.032 ;
      RECT 151.555 -89.515 151.695 -89.345 ;
      RECT 151.555 -88.618 151.645 -87.611 ;
      RECT 151.555 -88.305 151.695 -88.135 ;
      RECT 151.555 -86.809 151.645 -85.802 ;
      RECT 151.555 -86.285 151.695 -86.115 ;
      RECT 151.555 -85.388 151.645 -84.381 ;
      RECT 151.555 -85.075 151.695 -84.905 ;
      RECT 151.555 -83.579 151.645 -82.572 ;
      RECT 151.555 -83.055 151.695 -82.885 ;
      RECT 151.555 -82.158 151.645 -81.151 ;
      RECT 151.555 -81.845 151.695 -81.675 ;
      RECT 151.555 -80.349 151.645 -79.342 ;
      RECT 151.555 -79.825 151.695 -79.655 ;
      RECT 151.555 -78.928 151.645 -77.921 ;
      RECT 151.555 -78.615 151.695 -78.445 ;
      RECT 151.555 -77.119 151.645 -76.112 ;
      RECT 151.555 -76.595 151.695 -76.425 ;
      RECT 151.555 -75.698 151.645 -74.691 ;
      RECT 151.555 -75.385 151.695 -75.215 ;
      RECT 151.555 -73.889 151.645 -72.882 ;
      RECT 151.555 -73.365 151.695 -73.195 ;
      RECT 151.555 -72.468 151.645 -71.461 ;
      RECT 151.555 -72.155 151.695 -71.985 ;
      RECT 151.555 -70.659 151.645 -69.652 ;
      RECT 151.555 -70.135 151.695 -69.965 ;
      RECT 151.555 -69.238 151.645 -68.231 ;
      RECT 151.555 -68.925 151.695 -68.755 ;
      RECT 151.555 -67.429 151.645 -66.422 ;
      RECT 151.555 -66.905 151.695 -66.735 ;
      RECT 151.555 -66.008 151.645 -65.001 ;
      RECT 151.555 -65.695 151.695 -65.525 ;
      RECT 151.555 -64.199 151.645 -63.192 ;
      RECT 151.555 -63.675 151.695 -63.505 ;
      RECT 151.555 -62.778 151.645 -61.771 ;
      RECT 151.555 -62.465 151.695 -62.295 ;
      RECT 151.555 -60.969 151.645 -59.962 ;
      RECT 151.555 -60.445 151.695 -60.275 ;
      RECT 151.555 -59.548 151.645 -58.541 ;
      RECT 151.555 -59.235 151.695 -59.065 ;
      RECT 151.555 -57.739 151.645 -56.732 ;
      RECT 151.555 -57.215 151.695 -57.045 ;
      RECT 151.555 -56.318 151.645 -55.311 ;
      RECT 151.555 -56.005 151.695 -55.835 ;
      RECT 151.555 -54.509 151.645 -53.502 ;
      RECT 151.555 -53.985 151.695 -53.815 ;
      RECT 151.555 -53.088 151.645 -52.081 ;
      RECT 151.555 -52.775 151.695 -52.605 ;
      RECT 151.555 -51.279 151.645 -50.272 ;
      RECT 151.555 -50.755 151.695 -50.585 ;
      RECT 151.555 -49.858 151.645 -48.851 ;
      RECT 151.555 -49.545 151.695 -49.375 ;
      RECT 151.555 -48.049 151.645 -47.042 ;
      RECT 151.555 -47.525 151.695 -47.355 ;
      RECT 151.555 -46.628 151.645 -45.621 ;
      RECT 151.555 -46.315 151.695 -46.145 ;
      RECT 151.555 -44.819 151.645 -43.812 ;
      RECT 151.555 -44.295 151.695 -44.125 ;
      RECT 151.555 -43.398 151.645 -42.391 ;
      RECT 151.555 -43.085 151.695 -42.915 ;
      RECT 151.555 -41.589 151.645 -40.582 ;
      RECT 151.555 -41.065 151.695 -40.895 ;
      RECT 151.555 -40.168 151.645 -39.161 ;
      RECT 151.555 -39.855 151.695 -39.685 ;
      RECT 151.555 -38.359 151.645 -37.352 ;
      RECT 151.555 -37.835 151.695 -37.665 ;
      RECT 151.555 -36.938 151.645 -35.931 ;
      RECT 151.555 -36.625 151.695 -36.455 ;
      RECT 151.555 -35.129 151.645 -34.122 ;
      RECT 151.555 -34.605 151.695 -34.435 ;
      RECT 151.555 -33.708 151.645 -32.701 ;
      RECT 151.555 -33.395 151.695 -33.225 ;
      RECT 151.555 -31.899 151.645 -30.892 ;
      RECT 151.555 -31.375 151.695 -31.205 ;
      RECT 151.555 -30.478 151.645 -29.471 ;
      RECT 151.555 -30.165 151.695 -29.995 ;
      RECT 151.555 -28.669 151.645 -27.662 ;
      RECT 151.555 -28.145 151.695 -27.975 ;
      RECT 151.555 -27.248 151.645 -26.241 ;
      RECT 151.555 -26.935 151.695 -26.765 ;
      RECT 151.555 -25.439 151.645 -24.432 ;
      RECT 151.555 -24.915 151.695 -24.745 ;
      RECT 151.555 -24.018 151.645 -23.011 ;
      RECT 151.555 -23.705 151.695 -23.535 ;
      RECT 151.555 -22.209 151.645 -21.202 ;
      RECT 151.555 -21.685 151.695 -21.515 ;
      RECT 151.555 -20.788 151.645 -19.781 ;
      RECT 151.555 -20.475 151.695 -20.305 ;
      RECT 151.555 -18.979 151.645 -17.972 ;
      RECT 151.555 -18.455 151.695 -18.285 ;
      RECT 151.555 -17.558 151.645 -16.551 ;
      RECT 151.555 -17.245 151.695 -17.075 ;
      RECT 151.555 -15.749 151.645 -14.742 ;
      RECT 151.555 -15.225 151.695 -15.055 ;
      RECT 151.555 -14.328 151.645 -13.321 ;
      RECT 151.555 -14.015 151.695 -13.845 ;
      RECT 151.555 -12.519 151.645 -11.512 ;
      RECT 151.555 -11.995 151.695 -11.825 ;
      RECT 151.555 -11.098 151.645 -10.091 ;
      RECT 151.555 -10.785 151.695 -10.615 ;
      RECT 151.555 -9.289 151.645 -8.282 ;
      RECT 151.555 -8.765 151.695 -8.595 ;
      RECT 151.555 -7.868 151.645 -6.861 ;
      RECT 151.555 -7.555 151.695 -7.385 ;
      RECT 151.555 -6.059 151.645 -5.052 ;
      RECT 151.555 -5.535 151.695 -5.365 ;
      RECT 151.555 -4.638 151.645 -3.631 ;
      RECT 151.555 -4.325 151.695 -4.155 ;
      RECT 151.555 -2.829 151.645 -1.822 ;
      RECT 151.555 -2.305 151.695 -2.135 ;
      RECT 151.555 -1.408 151.645 -0.401 ;
      RECT 151.555 -1.095 151.695 -0.925 ;
      RECT 151.555 0.401 151.645 1.408 ;
      RECT 151.555 0.925 151.695 1.095 ;
      RECT -5.145 -110.99 -4.965 -110.81 ;
      RECT -5.145 -110.945 151.665 -110.855 ;
      RECT 149.705 -111.685 151.185 -111.585 ;
      RECT 149.705 -112.055 149.805 -111.585 ;
      RECT 149.51 -114.395 151.085 -114.275 ;
      RECT 150.985 -114.895 151.085 -114.275 ;
      RECT 150.39 -114.895 150.49 -114.275 ;
      RECT 149.51 -114.85 149.61 -114.275 ;
      RECT -2.285 -106.42 -2.105 -106.24 ;
      RECT -2.285 -106.375 151.03 -106.285 ;
      RECT 150.755 -101.538 150.845 -100.53 ;
      RECT 150.705 -100.935 150.845 -100.765 ;
      RECT 150.755 -99.73 150.845 -98.722 ;
      RECT 150.705 -99.495 150.845 -99.325 ;
      RECT 150.755 -98.308 150.845 -97.3 ;
      RECT 150.705 -97.705 150.845 -97.535 ;
      RECT 150.755 -96.5 150.845 -95.492 ;
      RECT 150.705 -96.265 150.845 -96.095 ;
      RECT 150.755 -95.078 150.845 -94.07 ;
      RECT 150.705 -94.475 150.845 -94.305 ;
      RECT 150.755 -93.27 150.845 -92.262 ;
      RECT 150.705 -93.035 150.845 -92.865 ;
      RECT 150.755 -91.848 150.845 -90.84 ;
      RECT 150.705 -91.245 150.845 -91.075 ;
      RECT 150.755 -90.04 150.845 -89.032 ;
      RECT 150.705 -89.805 150.845 -89.635 ;
      RECT 150.755 -88.618 150.845 -87.61 ;
      RECT 150.705 -88.015 150.845 -87.845 ;
      RECT 150.755 -86.81 150.845 -85.802 ;
      RECT 150.705 -86.575 150.845 -86.405 ;
      RECT 150.755 -85.388 150.845 -84.38 ;
      RECT 150.705 -84.785 150.845 -84.615 ;
      RECT 150.755 -83.58 150.845 -82.572 ;
      RECT 150.705 -83.345 150.845 -83.175 ;
      RECT 150.755 -82.158 150.845 -81.15 ;
      RECT 150.705 -81.555 150.845 -81.385 ;
      RECT 150.755 -80.35 150.845 -79.342 ;
      RECT 150.705 -80.115 150.845 -79.945 ;
      RECT 150.755 -78.928 150.845 -77.92 ;
      RECT 150.705 -78.325 150.845 -78.155 ;
      RECT 150.755 -77.12 150.845 -76.112 ;
      RECT 150.705 -76.885 150.845 -76.715 ;
      RECT 150.755 -75.698 150.845 -74.69 ;
      RECT 150.705 -75.095 150.845 -74.925 ;
      RECT 150.755 -73.89 150.845 -72.882 ;
      RECT 150.705 -73.655 150.845 -73.485 ;
      RECT 150.755 -72.468 150.845 -71.46 ;
      RECT 150.705 -71.865 150.845 -71.695 ;
      RECT 150.755 -70.66 150.845 -69.652 ;
      RECT 150.705 -70.425 150.845 -70.255 ;
      RECT 150.755 -69.238 150.845 -68.23 ;
      RECT 150.705 -68.635 150.845 -68.465 ;
      RECT 150.755 -67.43 150.845 -66.422 ;
      RECT 150.705 -67.195 150.845 -67.025 ;
      RECT 150.755 -66.008 150.845 -65 ;
      RECT 150.705 -65.405 150.845 -65.235 ;
      RECT 150.755 -64.2 150.845 -63.192 ;
      RECT 150.705 -63.965 150.845 -63.795 ;
      RECT 150.755 -62.778 150.845 -61.77 ;
      RECT 150.705 -62.175 150.845 -62.005 ;
      RECT 150.755 -60.97 150.845 -59.962 ;
      RECT 150.705 -60.735 150.845 -60.565 ;
      RECT 150.755 -59.548 150.845 -58.54 ;
      RECT 150.705 -58.945 150.845 -58.775 ;
      RECT 150.755 -57.74 150.845 -56.732 ;
      RECT 150.705 -57.505 150.845 -57.335 ;
      RECT 150.755 -56.318 150.845 -55.31 ;
      RECT 150.705 -55.715 150.845 -55.545 ;
      RECT 150.755 -54.51 150.845 -53.502 ;
      RECT 150.705 -54.275 150.845 -54.105 ;
      RECT 150.755 -53.088 150.845 -52.08 ;
      RECT 150.705 -52.485 150.845 -52.315 ;
      RECT 150.755 -51.28 150.845 -50.272 ;
      RECT 150.705 -51.045 150.845 -50.875 ;
      RECT 150.755 -49.858 150.845 -48.85 ;
      RECT 150.705 -49.255 150.845 -49.085 ;
      RECT 150.755 -48.05 150.845 -47.042 ;
      RECT 150.705 -47.815 150.845 -47.645 ;
      RECT 150.755 -46.628 150.845 -45.62 ;
      RECT 150.705 -46.025 150.845 -45.855 ;
      RECT 150.755 -44.82 150.845 -43.812 ;
      RECT 150.705 -44.585 150.845 -44.415 ;
      RECT 150.755 -43.398 150.845 -42.39 ;
      RECT 150.705 -42.795 150.845 -42.625 ;
      RECT 150.755 -41.59 150.845 -40.582 ;
      RECT 150.705 -41.355 150.845 -41.185 ;
      RECT 150.755 -40.168 150.845 -39.16 ;
      RECT 150.705 -39.565 150.845 -39.395 ;
      RECT 150.755 -38.36 150.845 -37.352 ;
      RECT 150.705 -38.125 150.845 -37.955 ;
      RECT 150.755 -36.938 150.845 -35.93 ;
      RECT 150.705 -36.335 150.845 -36.165 ;
      RECT 150.755 -35.13 150.845 -34.122 ;
      RECT 150.705 -34.895 150.845 -34.725 ;
      RECT 150.755 -33.708 150.845 -32.7 ;
      RECT 150.705 -33.105 150.845 -32.935 ;
      RECT 150.755 -31.9 150.845 -30.892 ;
      RECT 150.705 -31.665 150.845 -31.495 ;
      RECT 150.755 -30.478 150.845 -29.47 ;
      RECT 150.705 -29.875 150.845 -29.705 ;
      RECT 150.755 -28.67 150.845 -27.662 ;
      RECT 150.705 -28.435 150.845 -28.265 ;
      RECT 150.755 -27.248 150.845 -26.24 ;
      RECT 150.705 -26.645 150.845 -26.475 ;
      RECT 150.755 -25.44 150.845 -24.432 ;
      RECT 150.705 -25.205 150.845 -25.035 ;
      RECT 150.755 -24.018 150.845 -23.01 ;
      RECT 150.705 -23.415 150.845 -23.245 ;
      RECT 150.755 -22.21 150.845 -21.202 ;
      RECT 150.705 -21.975 150.845 -21.805 ;
      RECT 150.755 -20.788 150.845 -19.78 ;
      RECT 150.705 -20.185 150.845 -20.015 ;
      RECT 150.755 -18.98 150.845 -17.972 ;
      RECT 150.705 -18.745 150.845 -18.575 ;
      RECT 150.755 -17.558 150.845 -16.55 ;
      RECT 150.705 -16.955 150.845 -16.785 ;
      RECT 150.755 -15.75 150.845 -14.742 ;
      RECT 150.705 -15.515 150.845 -15.345 ;
      RECT 150.755 -14.328 150.845 -13.32 ;
      RECT 150.705 -13.725 150.845 -13.555 ;
      RECT 150.755 -12.52 150.845 -11.512 ;
      RECT 150.705 -12.285 150.845 -12.115 ;
      RECT 150.755 -11.098 150.845 -10.09 ;
      RECT 150.705 -10.495 150.845 -10.325 ;
      RECT 150.755 -9.29 150.845 -8.282 ;
      RECT 150.705 -9.055 150.845 -8.885 ;
      RECT 150.755 -7.868 150.845 -6.86 ;
      RECT 150.705 -7.265 150.845 -7.095 ;
      RECT 150.755 -6.06 150.845 -5.052 ;
      RECT 150.705 -5.825 150.845 -5.655 ;
      RECT 150.755 -4.638 150.845 -3.63 ;
      RECT 150.705 -4.035 150.845 -3.865 ;
      RECT 150.755 -2.83 150.845 -1.822 ;
      RECT 150.705 -2.595 150.845 -2.425 ;
      RECT 150.755 -1.408 150.845 -0.4 ;
      RECT 150.705 -0.805 150.845 -0.635 ;
      RECT 150.755 0.4 150.845 1.408 ;
      RECT 150.705 0.635 150.845 0.805 ;
      RECT 150.63 -114.685 150.805 -114.515 ;
      RECT 150.705 -114.895 150.805 -114.515 ;
      RECT 149.745 -113.555 149.845 -113.09 ;
      RECT 150.11 -113.555 150.21 -113.1 ;
      RECT 149.745 -113.555 150.59 -113.385 ;
      RECT 150.355 -101.538 150.445 -100.531 ;
      RECT 150.355 -101.225 150.495 -101.055 ;
      RECT 150.355 -99.729 150.445 -98.722 ;
      RECT 150.355 -99.205 150.495 -99.035 ;
      RECT 150.355 -98.308 150.445 -97.301 ;
      RECT 150.355 -97.995 150.495 -97.825 ;
      RECT 150.355 -96.499 150.445 -95.492 ;
      RECT 150.355 -95.975 150.495 -95.805 ;
      RECT 150.355 -95.078 150.445 -94.071 ;
      RECT 150.355 -94.765 150.495 -94.595 ;
      RECT 150.355 -93.269 150.445 -92.262 ;
      RECT 150.355 -92.745 150.495 -92.575 ;
      RECT 150.355 -91.848 150.445 -90.841 ;
      RECT 150.355 -91.535 150.495 -91.365 ;
      RECT 150.355 -90.039 150.445 -89.032 ;
      RECT 150.355 -89.515 150.495 -89.345 ;
      RECT 150.355 -88.618 150.445 -87.611 ;
      RECT 150.355 -88.305 150.495 -88.135 ;
      RECT 150.355 -86.809 150.445 -85.802 ;
      RECT 150.355 -86.285 150.495 -86.115 ;
      RECT 150.355 -85.388 150.445 -84.381 ;
      RECT 150.355 -85.075 150.495 -84.905 ;
      RECT 150.355 -83.579 150.445 -82.572 ;
      RECT 150.355 -83.055 150.495 -82.885 ;
      RECT 150.355 -82.158 150.445 -81.151 ;
      RECT 150.355 -81.845 150.495 -81.675 ;
      RECT 150.355 -80.349 150.445 -79.342 ;
      RECT 150.355 -79.825 150.495 -79.655 ;
      RECT 150.355 -78.928 150.445 -77.921 ;
      RECT 150.355 -78.615 150.495 -78.445 ;
      RECT 150.355 -77.119 150.445 -76.112 ;
      RECT 150.355 -76.595 150.495 -76.425 ;
      RECT 150.355 -75.698 150.445 -74.691 ;
      RECT 150.355 -75.385 150.495 -75.215 ;
      RECT 150.355 -73.889 150.445 -72.882 ;
      RECT 150.355 -73.365 150.495 -73.195 ;
      RECT 150.355 -72.468 150.445 -71.461 ;
      RECT 150.355 -72.155 150.495 -71.985 ;
      RECT 150.355 -70.659 150.445 -69.652 ;
      RECT 150.355 -70.135 150.495 -69.965 ;
      RECT 150.355 -69.238 150.445 -68.231 ;
      RECT 150.355 -68.925 150.495 -68.755 ;
      RECT 150.355 -67.429 150.445 -66.422 ;
      RECT 150.355 -66.905 150.495 -66.735 ;
      RECT 150.355 -66.008 150.445 -65.001 ;
      RECT 150.355 -65.695 150.495 -65.525 ;
      RECT 150.355 -64.199 150.445 -63.192 ;
      RECT 150.355 -63.675 150.495 -63.505 ;
      RECT 150.355 -62.778 150.445 -61.771 ;
      RECT 150.355 -62.465 150.495 -62.295 ;
      RECT 150.355 -60.969 150.445 -59.962 ;
      RECT 150.355 -60.445 150.495 -60.275 ;
      RECT 150.355 -59.548 150.445 -58.541 ;
      RECT 150.355 -59.235 150.495 -59.065 ;
      RECT 150.355 -57.739 150.445 -56.732 ;
      RECT 150.355 -57.215 150.495 -57.045 ;
      RECT 150.355 -56.318 150.445 -55.311 ;
      RECT 150.355 -56.005 150.495 -55.835 ;
      RECT 150.355 -54.509 150.445 -53.502 ;
      RECT 150.355 -53.985 150.495 -53.815 ;
      RECT 150.355 -53.088 150.445 -52.081 ;
      RECT 150.355 -52.775 150.495 -52.605 ;
      RECT 150.355 -51.279 150.445 -50.272 ;
      RECT 150.355 -50.755 150.495 -50.585 ;
      RECT 150.355 -49.858 150.445 -48.851 ;
      RECT 150.355 -49.545 150.495 -49.375 ;
      RECT 150.355 -48.049 150.445 -47.042 ;
      RECT 150.355 -47.525 150.495 -47.355 ;
      RECT 150.355 -46.628 150.445 -45.621 ;
      RECT 150.355 -46.315 150.495 -46.145 ;
      RECT 150.355 -44.819 150.445 -43.812 ;
      RECT 150.355 -44.295 150.495 -44.125 ;
      RECT 150.355 -43.398 150.445 -42.391 ;
      RECT 150.355 -43.085 150.495 -42.915 ;
      RECT 150.355 -41.589 150.445 -40.582 ;
      RECT 150.355 -41.065 150.495 -40.895 ;
      RECT 150.355 -40.168 150.445 -39.161 ;
      RECT 150.355 -39.855 150.495 -39.685 ;
      RECT 150.355 -38.359 150.445 -37.352 ;
      RECT 150.355 -37.835 150.495 -37.665 ;
      RECT 150.355 -36.938 150.445 -35.931 ;
      RECT 150.355 -36.625 150.495 -36.455 ;
      RECT 150.355 -35.129 150.445 -34.122 ;
      RECT 150.355 -34.605 150.495 -34.435 ;
      RECT 150.355 -33.708 150.445 -32.701 ;
      RECT 150.355 -33.395 150.495 -33.225 ;
      RECT 150.355 -31.899 150.445 -30.892 ;
      RECT 150.355 -31.375 150.495 -31.205 ;
      RECT 150.355 -30.478 150.445 -29.471 ;
      RECT 150.355 -30.165 150.495 -29.995 ;
      RECT 150.355 -28.669 150.445 -27.662 ;
      RECT 150.355 -28.145 150.495 -27.975 ;
      RECT 150.355 -27.248 150.445 -26.241 ;
      RECT 150.355 -26.935 150.495 -26.765 ;
      RECT 150.355 -25.439 150.445 -24.432 ;
      RECT 150.355 -24.915 150.495 -24.745 ;
      RECT 150.355 -24.018 150.445 -23.011 ;
      RECT 150.355 -23.705 150.495 -23.535 ;
      RECT 150.355 -22.209 150.445 -21.202 ;
      RECT 150.355 -21.685 150.495 -21.515 ;
      RECT 150.355 -20.788 150.445 -19.781 ;
      RECT 150.355 -20.475 150.495 -20.305 ;
      RECT 150.355 -18.979 150.445 -17.972 ;
      RECT 150.355 -18.455 150.495 -18.285 ;
      RECT 150.355 -17.558 150.445 -16.551 ;
      RECT 150.355 -17.245 150.495 -17.075 ;
      RECT 150.355 -15.749 150.445 -14.742 ;
      RECT 150.355 -15.225 150.495 -15.055 ;
      RECT 150.355 -14.328 150.445 -13.321 ;
      RECT 150.355 -14.015 150.495 -13.845 ;
      RECT 150.355 -12.519 150.445 -11.512 ;
      RECT 150.355 -11.995 150.495 -11.825 ;
      RECT 150.355 -11.098 150.445 -10.091 ;
      RECT 150.355 -10.785 150.495 -10.615 ;
      RECT 150.355 -9.289 150.445 -8.282 ;
      RECT 150.355 -8.765 150.495 -8.595 ;
      RECT 150.355 -7.868 150.445 -6.861 ;
      RECT 150.355 -7.555 150.495 -7.385 ;
      RECT 150.355 -6.059 150.445 -5.052 ;
      RECT 150.355 -5.535 150.495 -5.365 ;
      RECT 150.355 -4.638 150.445 -3.631 ;
      RECT 150.355 -4.325 150.495 -4.155 ;
      RECT 150.355 -2.829 150.445 -1.822 ;
      RECT 150.355 -2.305 150.495 -2.135 ;
      RECT 150.355 -1.408 150.445 -0.401 ;
      RECT 150.355 -1.095 150.495 -0.925 ;
      RECT 150.355 0.401 150.445 1.408 ;
      RECT 150.355 0.925 150.495 1.095 ;
      RECT 150.04 -114.685 150.21 -114.515 ;
      RECT 150.11 -114.895 150.21 -114.515 ;
      RECT -0.985 -106.94 -0.805 -106.76 ;
      RECT -1.925 -106.895 149.83 -106.805 ;
      RECT 149.555 -101.538 149.645 -100.53 ;
      RECT 149.505 -100.935 149.645 -100.765 ;
      RECT 149.555 -99.73 149.645 -98.722 ;
      RECT 149.505 -99.495 149.645 -99.325 ;
      RECT 149.555 -98.308 149.645 -97.3 ;
      RECT 149.505 -97.705 149.645 -97.535 ;
      RECT 149.555 -96.5 149.645 -95.492 ;
      RECT 149.505 -96.265 149.645 -96.095 ;
      RECT 149.555 -95.078 149.645 -94.07 ;
      RECT 149.505 -94.475 149.645 -94.305 ;
      RECT 149.555 -93.27 149.645 -92.262 ;
      RECT 149.505 -93.035 149.645 -92.865 ;
      RECT 149.555 -91.848 149.645 -90.84 ;
      RECT 149.505 -91.245 149.645 -91.075 ;
      RECT 149.555 -90.04 149.645 -89.032 ;
      RECT 149.505 -89.805 149.645 -89.635 ;
      RECT 149.555 -88.618 149.645 -87.61 ;
      RECT 149.505 -88.015 149.645 -87.845 ;
      RECT 149.555 -86.81 149.645 -85.802 ;
      RECT 149.505 -86.575 149.645 -86.405 ;
      RECT 149.555 -85.388 149.645 -84.38 ;
      RECT 149.505 -84.785 149.645 -84.615 ;
      RECT 149.555 -83.58 149.645 -82.572 ;
      RECT 149.505 -83.345 149.645 -83.175 ;
      RECT 149.555 -82.158 149.645 -81.15 ;
      RECT 149.505 -81.555 149.645 -81.385 ;
      RECT 149.555 -80.35 149.645 -79.342 ;
      RECT 149.505 -80.115 149.645 -79.945 ;
      RECT 149.555 -78.928 149.645 -77.92 ;
      RECT 149.505 -78.325 149.645 -78.155 ;
      RECT 149.555 -77.12 149.645 -76.112 ;
      RECT 149.505 -76.885 149.645 -76.715 ;
      RECT 149.555 -75.698 149.645 -74.69 ;
      RECT 149.505 -75.095 149.645 -74.925 ;
      RECT 149.555 -73.89 149.645 -72.882 ;
      RECT 149.505 -73.655 149.645 -73.485 ;
      RECT 149.555 -72.468 149.645 -71.46 ;
      RECT 149.505 -71.865 149.645 -71.695 ;
      RECT 149.555 -70.66 149.645 -69.652 ;
      RECT 149.505 -70.425 149.645 -70.255 ;
      RECT 149.555 -69.238 149.645 -68.23 ;
      RECT 149.505 -68.635 149.645 -68.465 ;
      RECT 149.555 -67.43 149.645 -66.422 ;
      RECT 149.505 -67.195 149.645 -67.025 ;
      RECT 149.555 -66.008 149.645 -65 ;
      RECT 149.505 -65.405 149.645 -65.235 ;
      RECT 149.555 -64.2 149.645 -63.192 ;
      RECT 149.505 -63.965 149.645 -63.795 ;
      RECT 149.555 -62.778 149.645 -61.77 ;
      RECT 149.505 -62.175 149.645 -62.005 ;
      RECT 149.555 -60.97 149.645 -59.962 ;
      RECT 149.505 -60.735 149.645 -60.565 ;
      RECT 149.555 -59.548 149.645 -58.54 ;
      RECT 149.505 -58.945 149.645 -58.775 ;
      RECT 149.555 -57.74 149.645 -56.732 ;
      RECT 149.505 -57.505 149.645 -57.335 ;
      RECT 149.555 -56.318 149.645 -55.31 ;
      RECT 149.505 -55.715 149.645 -55.545 ;
      RECT 149.555 -54.51 149.645 -53.502 ;
      RECT 149.505 -54.275 149.645 -54.105 ;
      RECT 149.555 -53.088 149.645 -52.08 ;
      RECT 149.505 -52.485 149.645 -52.315 ;
      RECT 149.555 -51.28 149.645 -50.272 ;
      RECT 149.505 -51.045 149.645 -50.875 ;
      RECT 149.555 -49.858 149.645 -48.85 ;
      RECT 149.505 -49.255 149.645 -49.085 ;
      RECT 149.555 -48.05 149.645 -47.042 ;
      RECT 149.505 -47.815 149.645 -47.645 ;
      RECT 149.555 -46.628 149.645 -45.62 ;
      RECT 149.505 -46.025 149.645 -45.855 ;
      RECT 149.555 -44.82 149.645 -43.812 ;
      RECT 149.505 -44.585 149.645 -44.415 ;
      RECT 149.555 -43.398 149.645 -42.39 ;
      RECT 149.505 -42.795 149.645 -42.625 ;
      RECT 149.555 -41.59 149.645 -40.582 ;
      RECT 149.505 -41.355 149.645 -41.185 ;
      RECT 149.555 -40.168 149.645 -39.16 ;
      RECT 149.505 -39.565 149.645 -39.395 ;
      RECT 149.555 -38.36 149.645 -37.352 ;
      RECT 149.505 -38.125 149.645 -37.955 ;
      RECT 149.555 -36.938 149.645 -35.93 ;
      RECT 149.505 -36.335 149.645 -36.165 ;
      RECT 149.555 -35.13 149.645 -34.122 ;
      RECT 149.505 -34.895 149.645 -34.725 ;
      RECT 149.555 -33.708 149.645 -32.7 ;
      RECT 149.505 -33.105 149.645 -32.935 ;
      RECT 149.555 -31.9 149.645 -30.892 ;
      RECT 149.505 -31.665 149.645 -31.495 ;
      RECT 149.555 -30.478 149.645 -29.47 ;
      RECT 149.505 -29.875 149.645 -29.705 ;
      RECT 149.555 -28.67 149.645 -27.662 ;
      RECT 149.505 -28.435 149.645 -28.265 ;
      RECT 149.555 -27.248 149.645 -26.24 ;
      RECT 149.505 -26.645 149.645 -26.475 ;
      RECT 149.555 -25.44 149.645 -24.432 ;
      RECT 149.505 -25.205 149.645 -25.035 ;
      RECT 149.555 -24.018 149.645 -23.01 ;
      RECT 149.505 -23.415 149.645 -23.245 ;
      RECT 149.555 -22.21 149.645 -21.202 ;
      RECT 149.505 -21.975 149.645 -21.805 ;
      RECT 149.555 -20.788 149.645 -19.78 ;
      RECT 149.505 -20.185 149.645 -20.015 ;
      RECT 149.555 -18.98 149.645 -17.972 ;
      RECT 149.505 -18.745 149.645 -18.575 ;
      RECT 149.555 -17.558 149.645 -16.55 ;
      RECT 149.505 -16.955 149.645 -16.785 ;
      RECT 149.555 -15.75 149.645 -14.742 ;
      RECT 149.505 -15.515 149.645 -15.345 ;
      RECT 149.555 -14.328 149.645 -13.32 ;
      RECT 149.505 -13.725 149.645 -13.555 ;
      RECT 149.555 -12.52 149.645 -11.512 ;
      RECT 149.505 -12.285 149.645 -12.115 ;
      RECT 149.555 -11.098 149.645 -10.09 ;
      RECT 149.505 -10.495 149.645 -10.325 ;
      RECT 149.555 -9.29 149.645 -8.282 ;
      RECT 149.505 -9.055 149.645 -8.885 ;
      RECT 149.555 -7.868 149.645 -6.86 ;
      RECT 149.505 -7.265 149.645 -7.095 ;
      RECT 149.555 -6.06 149.645 -5.052 ;
      RECT 149.505 -5.825 149.645 -5.655 ;
      RECT 149.555 -4.638 149.645 -3.63 ;
      RECT 149.505 -4.035 149.645 -3.865 ;
      RECT 149.555 -2.83 149.645 -1.822 ;
      RECT 149.505 -2.595 149.645 -2.425 ;
      RECT 149.555 -1.408 149.645 -0.4 ;
      RECT 149.505 -0.805 149.645 -0.635 ;
      RECT 149.555 0.4 149.645 1.408 ;
      RECT 149.505 0.635 149.645 0.805 ;
      RECT 149.155 -101.538 149.245 -100.531 ;
      RECT 149.155 -101.225 149.295 -101.055 ;
      RECT 149.155 -99.729 149.245 -98.722 ;
      RECT 149.155 -99.205 149.295 -99.035 ;
      RECT 149.155 -98.308 149.245 -97.301 ;
      RECT 149.155 -97.995 149.295 -97.825 ;
      RECT 149.155 -96.499 149.245 -95.492 ;
      RECT 149.155 -95.975 149.295 -95.805 ;
      RECT 149.155 -95.078 149.245 -94.071 ;
      RECT 149.155 -94.765 149.295 -94.595 ;
      RECT 149.155 -93.269 149.245 -92.262 ;
      RECT 149.155 -92.745 149.295 -92.575 ;
      RECT 149.155 -91.848 149.245 -90.841 ;
      RECT 149.155 -91.535 149.295 -91.365 ;
      RECT 149.155 -90.039 149.245 -89.032 ;
      RECT 149.155 -89.515 149.295 -89.345 ;
      RECT 149.155 -88.618 149.245 -87.611 ;
      RECT 149.155 -88.305 149.295 -88.135 ;
      RECT 149.155 -86.809 149.245 -85.802 ;
      RECT 149.155 -86.285 149.295 -86.115 ;
      RECT 149.155 -85.388 149.245 -84.381 ;
      RECT 149.155 -85.075 149.295 -84.905 ;
      RECT 149.155 -83.579 149.245 -82.572 ;
      RECT 149.155 -83.055 149.295 -82.885 ;
      RECT 149.155 -82.158 149.245 -81.151 ;
      RECT 149.155 -81.845 149.295 -81.675 ;
      RECT 149.155 -80.349 149.245 -79.342 ;
      RECT 149.155 -79.825 149.295 -79.655 ;
      RECT 149.155 -78.928 149.245 -77.921 ;
      RECT 149.155 -78.615 149.295 -78.445 ;
      RECT 149.155 -77.119 149.245 -76.112 ;
      RECT 149.155 -76.595 149.295 -76.425 ;
      RECT 149.155 -75.698 149.245 -74.691 ;
      RECT 149.155 -75.385 149.295 -75.215 ;
      RECT 149.155 -73.889 149.245 -72.882 ;
      RECT 149.155 -73.365 149.295 -73.195 ;
      RECT 149.155 -72.468 149.245 -71.461 ;
      RECT 149.155 -72.155 149.295 -71.985 ;
      RECT 149.155 -70.659 149.245 -69.652 ;
      RECT 149.155 -70.135 149.295 -69.965 ;
      RECT 149.155 -69.238 149.245 -68.231 ;
      RECT 149.155 -68.925 149.295 -68.755 ;
      RECT 149.155 -67.429 149.245 -66.422 ;
      RECT 149.155 -66.905 149.295 -66.735 ;
      RECT 149.155 -66.008 149.245 -65.001 ;
      RECT 149.155 -65.695 149.295 -65.525 ;
      RECT 149.155 -64.199 149.245 -63.192 ;
      RECT 149.155 -63.675 149.295 -63.505 ;
      RECT 149.155 -62.778 149.245 -61.771 ;
      RECT 149.155 -62.465 149.295 -62.295 ;
      RECT 149.155 -60.969 149.245 -59.962 ;
      RECT 149.155 -60.445 149.295 -60.275 ;
      RECT 149.155 -59.548 149.245 -58.541 ;
      RECT 149.155 -59.235 149.295 -59.065 ;
      RECT 149.155 -57.739 149.245 -56.732 ;
      RECT 149.155 -57.215 149.295 -57.045 ;
      RECT 149.155 -56.318 149.245 -55.311 ;
      RECT 149.155 -56.005 149.295 -55.835 ;
      RECT 149.155 -54.509 149.245 -53.502 ;
      RECT 149.155 -53.985 149.295 -53.815 ;
      RECT 149.155 -53.088 149.245 -52.081 ;
      RECT 149.155 -52.775 149.295 -52.605 ;
      RECT 149.155 -51.279 149.245 -50.272 ;
      RECT 149.155 -50.755 149.295 -50.585 ;
      RECT 149.155 -49.858 149.245 -48.851 ;
      RECT 149.155 -49.545 149.295 -49.375 ;
      RECT 149.155 -48.049 149.245 -47.042 ;
      RECT 149.155 -47.525 149.295 -47.355 ;
      RECT 149.155 -46.628 149.245 -45.621 ;
      RECT 149.155 -46.315 149.295 -46.145 ;
      RECT 149.155 -44.819 149.245 -43.812 ;
      RECT 149.155 -44.295 149.295 -44.125 ;
      RECT 149.155 -43.398 149.245 -42.391 ;
      RECT 149.155 -43.085 149.295 -42.915 ;
      RECT 149.155 -41.589 149.245 -40.582 ;
      RECT 149.155 -41.065 149.295 -40.895 ;
      RECT 149.155 -40.168 149.245 -39.161 ;
      RECT 149.155 -39.855 149.295 -39.685 ;
      RECT 149.155 -38.359 149.245 -37.352 ;
      RECT 149.155 -37.835 149.295 -37.665 ;
      RECT 149.155 -36.938 149.245 -35.931 ;
      RECT 149.155 -36.625 149.295 -36.455 ;
      RECT 149.155 -35.129 149.245 -34.122 ;
      RECT 149.155 -34.605 149.295 -34.435 ;
      RECT 149.155 -33.708 149.245 -32.701 ;
      RECT 149.155 -33.395 149.295 -33.225 ;
      RECT 149.155 -31.899 149.245 -30.892 ;
      RECT 149.155 -31.375 149.295 -31.205 ;
      RECT 149.155 -30.478 149.245 -29.471 ;
      RECT 149.155 -30.165 149.295 -29.995 ;
      RECT 149.155 -28.669 149.245 -27.662 ;
      RECT 149.155 -28.145 149.295 -27.975 ;
      RECT 149.155 -27.248 149.245 -26.241 ;
      RECT 149.155 -26.935 149.295 -26.765 ;
      RECT 149.155 -25.439 149.245 -24.432 ;
      RECT 149.155 -24.915 149.295 -24.745 ;
      RECT 149.155 -24.018 149.245 -23.011 ;
      RECT 149.155 -23.705 149.295 -23.535 ;
      RECT 149.155 -22.209 149.245 -21.202 ;
      RECT 149.155 -21.685 149.295 -21.515 ;
      RECT 149.155 -20.788 149.245 -19.781 ;
      RECT 149.155 -20.475 149.295 -20.305 ;
      RECT 149.155 -18.979 149.245 -17.972 ;
      RECT 149.155 -18.455 149.295 -18.285 ;
      RECT 149.155 -17.558 149.245 -16.551 ;
      RECT 149.155 -17.245 149.295 -17.075 ;
      RECT 149.155 -15.749 149.245 -14.742 ;
      RECT 149.155 -15.225 149.295 -15.055 ;
      RECT 149.155 -14.328 149.245 -13.321 ;
      RECT 149.155 -14.015 149.295 -13.845 ;
      RECT 149.155 -12.519 149.245 -11.512 ;
      RECT 149.155 -11.995 149.295 -11.825 ;
      RECT 149.155 -11.098 149.245 -10.091 ;
      RECT 149.155 -10.785 149.295 -10.615 ;
      RECT 149.155 -9.289 149.245 -8.282 ;
      RECT 149.155 -8.765 149.295 -8.595 ;
      RECT 149.155 -7.868 149.245 -6.861 ;
      RECT 149.155 -7.555 149.295 -7.385 ;
      RECT 149.155 -6.059 149.245 -5.052 ;
      RECT 149.155 -5.535 149.295 -5.365 ;
      RECT 149.155 -4.638 149.245 -3.631 ;
      RECT 149.155 -4.325 149.295 -4.155 ;
      RECT 149.155 -2.829 149.245 -1.822 ;
      RECT 149.155 -2.305 149.295 -2.135 ;
      RECT 149.155 -1.408 149.245 -0.401 ;
      RECT 149.155 -1.095 149.295 -0.925 ;
      RECT 149.155 0.401 149.245 1.408 ;
      RECT 149.155 0.925 149.295 1.095 ;
      RECT 144.985 -108.935 148.765 -108.815 ;
      RECT 146.305 -109.475 146.405 -108.815 ;
      RECT 145.745 -109.475 145.845 -108.815 ;
      RECT 145.185 -109.475 145.285 -108.815 ;
      RECT 148.355 -101.538 148.445 -100.53 ;
      RECT 148.305 -100.935 148.445 -100.765 ;
      RECT 148.355 -99.73 148.445 -98.722 ;
      RECT 148.305 -99.495 148.445 -99.325 ;
      RECT 148.355 -98.308 148.445 -97.3 ;
      RECT 148.305 -97.705 148.445 -97.535 ;
      RECT 148.355 -96.5 148.445 -95.492 ;
      RECT 148.305 -96.265 148.445 -96.095 ;
      RECT 148.355 -95.078 148.445 -94.07 ;
      RECT 148.305 -94.475 148.445 -94.305 ;
      RECT 148.355 -93.27 148.445 -92.262 ;
      RECT 148.305 -93.035 148.445 -92.865 ;
      RECT 148.355 -91.848 148.445 -90.84 ;
      RECT 148.305 -91.245 148.445 -91.075 ;
      RECT 148.355 -90.04 148.445 -89.032 ;
      RECT 148.305 -89.805 148.445 -89.635 ;
      RECT 148.355 -88.618 148.445 -87.61 ;
      RECT 148.305 -88.015 148.445 -87.845 ;
      RECT 148.355 -86.81 148.445 -85.802 ;
      RECT 148.305 -86.575 148.445 -86.405 ;
      RECT 148.355 -85.388 148.445 -84.38 ;
      RECT 148.305 -84.785 148.445 -84.615 ;
      RECT 148.355 -83.58 148.445 -82.572 ;
      RECT 148.305 -83.345 148.445 -83.175 ;
      RECT 148.355 -82.158 148.445 -81.15 ;
      RECT 148.305 -81.555 148.445 -81.385 ;
      RECT 148.355 -80.35 148.445 -79.342 ;
      RECT 148.305 -80.115 148.445 -79.945 ;
      RECT 148.355 -78.928 148.445 -77.92 ;
      RECT 148.305 -78.325 148.445 -78.155 ;
      RECT 148.355 -77.12 148.445 -76.112 ;
      RECT 148.305 -76.885 148.445 -76.715 ;
      RECT 148.355 -75.698 148.445 -74.69 ;
      RECT 148.305 -75.095 148.445 -74.925 ;
      RECT 148.355 -73.89 148.445 -72.882 ;
      RECT 148.305 -73.655 148.445 -73.485 ;
      RECT 148.355 -72.468 148.445 -71.46 ;
      RECT 148.305 -71.865 148.445 -71.695 ;
      RECT 148.355 -70.66 148.445 -69.652 ;
      RECT 148.305 -70.425 148.445 -70.255 ;
      RECT 148.355 -69.238 148.445 -68.23 ;
      RECT 148.305 -68.635 148.445 -68.465 ;
      RECT 148.355 -67.43 148.445 -66.422 ;
      RECT 148.305 -67.195 148.445 -67.025 ;
      RECT 148.355 -66.008 148.445 -65 ;
      RECT 148.305 -65.405 148.445 -65.235 ;
      RECT 148.355 -64.2 148.445 -63.192 ;
      RECT 148.305 -63.965 148.445 -63.795 ;
      RECT 148.355 -62.778 148.445 -61.77 ;
      RECT 148.305 -62.175 148.445 -62.005 ;
      RECT 148.355 -60.97 148.445 -59.962 ;
      RECT 148.305 -60.735 148.445 -60.565 ;
      RECT 148.355 -59.548 148.445 -58.54 ;
      RECT 148.305 -58.945 148.445 -58.775 ;
      RECT 148.355 -57.74 148.445 -56.732 ;
      RECT 148.305 -57.505 148.445 -57.335 ;
      RECT 148.355 -56.318 148.445 -55.31 ;
      RECT 148.305 -55.715 148.445 -55.545 ;
      RECT 148.355 -54.51 148.445 -53.502 ;
      RECT 148.305 -54.275 148.445 -54.105 ;
      RECT 148.355 -53.088 148.445 -52.08 ;
      RECT 148.305 -52.485 148.445 -52.315 ;
      RECT 148.355 -51.28 148.445 -50.272 ;
      RECT 148.305 -51.045 148.445 -50.875 ;
      RECT 148.355 -49.858 148.445 -48.85 ;
      RECT 148.305 -49.255 148.445 -49.085 ;
      RECT 148.355 -48.05 148.445 -47.042 ;
      RECT 148.305 -47.815 148.445 -47.645 ;
      RECT 148.355 -46.628 148.445 -45.62 ;
      RECT 148.305 -46.025 148.445 -45.855 ;
      RECT 148.355 -44.82 148.445 -43.812 ;
      RECT 148.305 -44.585 148.445 -44.415 ;
      RECT 148.355 -43.398 148.445 -42.39 ;
      RECT 148.305 -42.795 148.445 -42.625 ;
      RECT 148.355 -41.59 148.445 -40.582 ;
      RECT 148.305 -41.355 148.445 -41.185 ;
      RECT 148.355 -40.168 148.445 -39.16 ;
      RECT 148.305 -39.565 148.445 -39.395 ;
      RECT 148.355 -38.36 148.445 -37.352 ;
      RECT 148.305 -38.125 148.445 -37.955 ;
      RECT 148.355 -36.938 148.445 -35.93 ;
      RECT 148.305 -36.335 148.445 -36.165 ;
      RECT 148.355 -35.13 148.445 -34.122 ;
      RECT 148.305 -34.895 148.445 -34.725 ;
      RECT 148.355 -33.708 148.445 -32.7 ;
      RECT 148.305 -33.105 148.445 -32.935 ;
      RECT 148.355 -31.9 148.445 -30.892 ;
      RECT 148.305 -31.665 148.445 -31.495 ;
      RECT 148.355 -30.478 148.445 -29.47 ;
      RECT 148.305 -29.875 148.445 -29.705 ;
      RECT 148.355 -28.67 148.445 -27.662 ;
      RECT 148.305 -28.435 148.445 -28.265 ;
      RECT 148.355 -27.248 148.445 -26.24 ;
      RECT 148.305 -26.645 148.445 -26.475 ;
      RECT 148.355 -25.44 148.445 -24.432 ;
      RECT 148.305 -25.205 148.445 -25.035 ;
      RECT 148.355 -24.018 148.445 -23.01 ;
      RECT 148.305 -23.415 148.445 -23.245 ;
      RECT 148.355 -22.21 148.445 -21.202 ;
      RECT 148.305 -21.975 148.445 -21.805 ;
      RECT 148.355 -20.788 148.445 -19.78 ;
      RECT 148.305 -20.185 148.445 -20.015 ;
      RECT 148.355 -18.98 148.445 -17.972 ;
      RECT 148.305 -18.745 148.445 -18.575 ;
      RECT 148.355 -17.558 148.445 -16.55 ;
      RECT 148.305 -16.955 148.445 -16.785 ;
      RECT 148.355 -15.75 148.445 -14.742 ;
      RECT 148.305 -15.515 148.445 -15.345 ;
      RECT 148.355 -14.328 148.445 -13.32 ;
      RECT 148.305 -13.725 148.445 -13.555 ;
      RECT 148.355 -12.52 148.445 -11.512 ;
      RECT 148.305 -12.285 148.445 -12.115 ;
      RECT 148.355 -11.098 148.445 -10.09 ;
      RECT 148.305 -10.495 148.445 -10.325 ;
      RECT 148.355 -9.29 148.445 -8.282 ;
      RECT 148.305 -9.055 148.445 -8.885 ;
      RECT 148.355 -7.868 148.445 -6.86 ;
      RECT 148.305 -7.265 148.445 -7.095 ;
      RECT 148.355 -6.06 148.445 -5.052 ;
      RECT 148.305 -5.825 148.445 -5.655 ;
      RECT 148.355 -4.638 148.445 -3.63 ;
      RECT 148.305 -4.035 148.445 -3.865 ;
      RECT 148.355 -2.83 148.445 -1.822 ;
      RECT 148.305 -2.595 148.445 -2.425 ;
      RECT 148.355 -1.408 148.445 -0.4 ;
      RECT 148.305 -0.805 148.445 -0.635 ;
      RECT 148.355 0.4 148.445 1.408 ;
      RECT 148.305 0.635 148.445 0.805 ;
      RECT 146.925 -111.685 148.405 -111.585 ;
      RECT 146.925 -112.195 147.025 -111.585 ;
      RECT 147.145 -109.15 148.405 -109.05 ;
      RECT 148.305 -109.475 148.405 -109.05 ;
      RECT 147.745 -109.475 147.845 -109.05 ;
      RECT 147.185 -109.475 147.285 -109.05 ;
      RECT 147.955 -101.538 148.045 -100.531 ;
      RECT 147.955 -101.225 148.095 -101.055 ;
      RECT 147.955 -99.729 148.045 -98.722 ;
      RECT 147.955 -99.205 148.095 -99.035 ;
      RECT 147.955 -98.308 148.045 -97.301 ;
      RECT 147.955 -97.995 148.095 -97.825 ;
      RECT 147.955 -96.499 148.045 -95.492 ;
      RECT 147.955 -95.975 148.095 -95.805 ;
      RECT 147.955 -95.078 148.045 -94.071 ;
      RECT 147.955 -94.765 148.095 -94.595 ;
      RECT 147.955 -93.269 148.045 -92.262 ;
      RECT 147.955 -92.745 148.095 -92.575 ;
      RECT 147.955 -91.848 148.045 -90.841 ;
      RECT 147.955 -91.535 148.095 -91.365 ;
      RECT 147.955 -90.039 148.045 -89.032 ;
      RECT 147.955 -89.515 148.095 -89.345 ;
      RECT 147.955 -88.618 148.045 -87.611 ;
      RECT 147.955 -88.305 148.095 -88.135 ;
      RECT 147.955 -86.809 148.045 -85.802 ;
      RECT 147.955 -86.285 148.095 -86.115 ;
      RECT 147.955 -85.388 148.045 -84.381 ;
      RECT 147.955 -85.075 148.095 -84.905 ;
      RECT 147.955 -83.579 148.045 -82.572 ;
      RECT 147.955 -83.055 148.095 -82.885 ;
      RECT 147.955 -82.158 148.045 -81.151 ;
      RECT 147.955 -81.845 148.095 -81.675 ;
      RECT 147.955 -80.349 148.045 -79.342 ;
      RECT 147.955 -79.825 148.095 -79.655 ;
      RECT 147.955 -78.928 148.045 -77.921 ;
      RECT 147.955 -78.615 148.095 -78.445 ;
      RECT 147.955 -77.119 148.045 -76.112 ;
      RECT 147.955 -76.595 148.095 -76.425 ;
      RECT 147.955 -75.698 148.045 -74.691 ;
      RECT 147.955 -75.385 148.095 -75.215 ;
      RECT 147.955 -73.889 148.045 -72.882 ;
      RECT 147.955 -73.365 148.095 -73.195 ;
      RECT 147.955 -72.468 148.045 -71.461 ;
      RECT 147.955 -72.155 148.095 -71.985 ;
      RECT 147.955 -70.659 148.045 -69.652 ;
      RECT 147.955 -70.135 148.095 -69.965 ;
      RECT 147.955 -69.238 148.045 -68.231 ;
      RECT 147.955 -68.925 148.095 -68.755 ;
      RECT 147.955 -67.429 148.045 -66.422 ;
      RECT 147.955 -66.905 148.095 -66.735 ;
      RECT 147.955 -66.008 148.045 -65.001 ;
      RECT 147.955 -65.695 148.095 -65.525 ;
      RECT 147.955 -64.199 148.045 -63.192 ;
      RECT 147.955 -63.675 148.095 -63.505 ;
      RECT 147.955 -62.778 148.045 -61.771 ;
      RECT 147.955 -62.465 148.095 -62.295 ;
      RECT 147.955 -60.969 148.045 -59.962 ;
      RECT 147.955 -60.445 148.095 -60.275 ;
      RECT 147.955 -59.548 148.045 -58.541 ;
      RECT 147.955 -59.235 148.095 -59.065 ;
      RECT 147.955 -57.739 148.045 -56.732 ;
      RECT 147.955 -57.215 148.095 -57.045 ;
      RECT 147.955 -56.318 148.045 -55.311 ;
      RECT 147.955 -56.005 148.095 -55.835 ;
      RECT 147.955 -54.509 148.045 -53.502 ;
      RECT 147.955 -53.985 148.095 -53.815 ;
      RECT 147.955 -53.088 148.045 -52.081 ;
      RECT 147.955 -52.775 148.095 -52.605 ;
      RECT 147.955 -51.279 148.045 -50.272 ;
      RECT 147.955 -50.755 148.095 -50.585 ;
      RECT 147.955 -49.858 148.045 -48.851 ;
      RECT 147.955 -49.545 148.095 -49.375 ;
      RECT 147.955 -48.049 148.045 -47.042 ;
      RECT 147.955 -47.525 148.095 -47.355 ;
      RECT 147.955 -46.628 148.045 -45.621 ;
      RECT 147.955 -46.315 148.095 -46.145 ;
      RECT 147.955 -44.819 148.045 -43.812 ;
      RECT 147.955 -44.295 148.095 -44.125 ;
      RECT 147.955 -43.398 148.045 -42.391 ;
      RECT 147.955 -43.085 148.095 -42.915 ;
      RECT 147.955 -41.589 148.045 -40.582 ;
      RECT 147.955 -41.065 148.095 -40.895 ;
      RECT 147.955 -40.168 148.045 -39.161 ;
      RECT 147.955 -39.855 148.095 -39.685 ;
      RECT 147.955 -38.359 148.045 -37.352 ;
      RECT 147.955 -37.835 148.095 -37.665 ;
      RECT 147.955 -36.938 148.045 -35.931 ;
      RECT 147.955 -36.625 148.095 -36.455 ;
      RECT 147.955 -35.129 148.045 -34.122 ;
      RECT 147.955 -34.605 148.095 -34.435 ;
      RECT 147.955 -33.708 148.045 -32.701 ;
      RECT 147.955 -33.395 148.095 -33.225 ;
      RECT 147.955 -31.899 148.045 -30.892 ;
      RECT 147.955 -31.375 148.095 -31.205 ;
      RECT 147.955 -30.478 148.045 -29.471 ;
      RECT 147.955 -30.165 148.095 -29.995 ;
      RECT 147.955 -28.669 148.045 -27.662 ;
      RECT 147.955 -28.145 148.095 -27.975 ;
      RECT 147.955 -27.248 148.045 -26.241 ;
      RECT 147.955 -26.935 148.095 -26.765 ;
      RECT 147.955 -25.439 148.045 -24.432 ;
      RECT 147.955 -24.915 148.095 -24.745 ;
      RECT 147.955 -24.018 148.045 -23.011 ;
      RECT 147.955 -23.705 148.095 -23.535 ;
      RECT 147.955 -22.209 148.045 -21.202 ;
      RECT 147.955 -21.685 148.095 -21.515 ;
      RECT 147.955 -20.788 148.045 -19.781 ;
      RECT 147.955 -20.475 148.095 -20.305 ;
      RECT 147.955 -18.979 148.045 -17.972 ;
      RECT 147.955 -18.455 148.095 -18.285 ;
      RECT 147.955 -17.558 148.045 -16.551 ;
      RECT 147.955 -17.245 148.095 -17.075 ;
      RECT 147.955 -15.749 148.045 -14.742 ;
      RECT 147.955 -15.225 148.095 -15.055 ;
      RECT 147.955 -14.328 148.045 -13.321 ;
      RECT 147.955 -14.015 148.095 -13.845 ;
      RECT 147.955 -12.519 148.045 -11.512 ;
      RECT 147.955 -11.995 148.095 -11.825 ;
      RECT 147.955 -11.098 148.045 -10.091 ;
      RECT 147.955 -10.785 148.095 -10.615 ;
      RECT 147.955 -9.289 148.045 -8.282 ;
      RECT 147.955 -8.765 148.095 -8.595 ;
      RECT 147.955 -7.868 148.045 -6.861 ;
      RECT 147.955 -7.555 148.095 -7.385 ;
      RECT 147.955 -6.059 148.045 -5.052 ;
      RECT 147.955 -5.535 148.095 -5.365 ;
      RECT 147.955 -4.638 148.045 -3.631 ;
      RECT 147.955 -4.325 148.095 -4.155 ;
      RECT 147.955 -2.829 148.045 -1.822 ;
      RECT 147.955 -2.305 148.095 -2.135 ;
      RECT 147.955 -1.408 148.045 -0.401 ;
      RECT 147.955 -1.095 148.095 -0.925 ;
      RECT 147.955 0.401 148.045 1.408 ;
      RECT 147.955 0.925 148.095 1.095 ;
      RECT 147.285 -111.495 147.455 -111.385 ;
      RECT 144.135 -111.495 147.455 -111.395 ;
      RECT 147.155 -101.538 147.245 -100.53 ;
      RECT 147.105 -100.935 147.245 -100.765 ;
      RECT 147.155 -99.73 147.245 -98.722 ;
      RECT 147.105 -99.495 147.245 -99.325 ;
      RECT 147.155 -98.308 147.245 -97.3 ;
      RECT 147.105 -97.705 147.245 -97.535 ;
      RECT 147.155 -96.5 147.245 -95.492 ;
      RECT 147.105 -96.265 147.245 -96.095 ;
      RECT 147.155 -95.078 147.245 -94.07 ;
      RECT 147.105 -94.475 147.245 -94.305 ;
      RECT 147.155 -93.27 147.245 -92.262 ;
      RECT 147.105 -93.035 147.245 -92.865 ;
      RECT 147.155 -91.848 147.245 -90.84 ;
      RECT 147.105 -91.245 147.245 -91.075 ;
      RECT 147.155 -90.04 147.245 -89.032 ;
      RECT 147.105 -89.805 147.245 -89.635 ;
      RECT 147.155 -88.618 147.245 -87.61 ;
      RECT 147.105 -88.015 147.245 -87.845 ;
      RECT 147.155 -86.81 147.245 -85.802 ;
      RECT 147.105 -86.575 147.245 -86.405 ;
      RECT 147.155 -85.388 147.245 -84.38 ;
      RECT 147.105 -84.785 147.245 -84.615 ;
      RECT 147.155 -83.58 147.245 -82.572 ;
      RECT 147.105 -83.345 147.245 -83.175 ;
      RECT 147.155 -82.158 147.245 -81.15 ;
      RECT 147.105 -81.555 147.245 -81.385 ;
      RECT 147.155 -80.35 147.245 -79.342 ;
      RECT 147.105 -80.115 147.245 -79.945 ;
      RECT 147.155 -78.928 147.245 -77.92 ;
      RECT 147.105 -78.325 147.245 -78.155 ;
      RECT 147.155 -77.12 147.245 -76.112 ;
      RECT 147.105 -76.885 147.245 -76.715 ;
      RECT 147.155 -75.698 147.245 -74.69 ;
      RECT 147.105 -75.095 147.245 -74.925 ;
      RECT 147.155 -73.89 147.245 -72.882 ;
      RECT 147.105 -73.655 147.245 -73.485 ;
      RECT 147.155 -72.468 147.245 -71.46 ;
      RECT 147.105 -71.865 147.245 -71.695 ;
      RECT 147.155 -70.66 147.245 -69.652 ;
      RECT 147.105 -70.425 147.245 -70.255 ;
      RECT 147.155 -69.238 147.245 -68.23 ;
      RECT 147.105 -68.635 147.245 -68.465 ;
      RECT 147.155 -67.43 147.245 -66.422 ;
      RECT 147.105 -67.195 147.245 -67.025 ;
      RECT 147.155 -66.008 147.245 -65 ;
      RECT 147.105 -65.405 147.245 -65.235 ;
      RECT 147.155 -64.2 147.245 -63.192 ;
      RECT 147.105 -63.965 147.245 -63.795 ;
      RECT 147.155 -62.778 147.245 -61.77 ;
      RECT 147.105 -62.175 147.245 -62.005 ;
      RECT 147.155 -60.97 147.245 -59.962 ;
      RECT 147.105 -60.735 147.245 -60.565 ;
      RECT 147.155 -59.548 147.245 -58.54 ;
      RECT 147.105 -58.945 147.245 -58.775 ;
      RECT 147.155 -57.74 147.245 -56.732 ;
      RECT 147.105 -57.505 147.245 -57.335 ;
      RECT 147.155 -56.318 147.245 -55.31 ;
      RECT 147.105 -55.715 147.245 -55.545 ;
      RECT 147.155 -54.51 147.245 -53.502 ;
      RECT 147.105 -54.275 147.245 -54.105 ;
      RECT 147.155 -53.088 147.245 -52.08 ;
      RECT 147.105 -52.485 147.245 -52.315 ;
      RECT 147.155 -51.28 147.245 -50.272 ;
      RECT 147.105 -51.045 147.245 -50.875 ;
      RECT 147.155 -49.858 147.245 -48.85 ;
      RECT 147.105 -49.255 147.245 -49.085 ;
      RECT 147.155 -48.05 147.245 -47.042 ;
      RECT 147.105 -47.815 147.245 -47.645 ;
      RECT 147.155 -46.628 147.245 -45.62 ;
      RECT 147.105 -46.025 147.245 -45.855 ;
      RECT 147.155 -44.82 147.245 -43.812 ;
      RECT 147.105 -44.585 147.245 -44.415 ;
      RECT 147.155 -43.398 147.245 -42.39 ;
      RECT 147.105 -42.795 147.245 -42.625 ;
      RECT 147.155 -41.59 147.245 -40.582 ;
      RECT 147.105 -41.355 147.245 -41.185 ;
      RECT 147.155 -40.168 147.245 -39.16 ;
      RECT 147.105 -39.565 147.245 -39.395 ;
      RECT 147.155 -38.36 147.245 -37.352 ;
      RECT 147.105 -38.125 147.245 -37.955 ;
      RECT 147.155 -36.938 147.245 -35.93 ;
      RECT 147.105 -36.335 147.245 -36.165 ;
      RECT 147.155 -35.13 147.245 -34.122 ;
      RECT 147.105 -34.895 147.245 -34.725 ;
      RECT 147.155 -33.708 147.245 -32.7 ;
      RECT 147.105 -33.105 147.245 -32.935 ;
      RECT 147.155 -31.9 147.245 -30.892 ;
      RECT 147.105 -31.665 147.245 -31.495 ;
      RECT 147.155 -30.478 147.245 -29.47 ;
      RECT 147.105 -29.875 147.245 -29.705 ;
      RECT 147.155 -28.67 147.245 -27.662 ;
      RECT 147.105 -28.435 147.245 -28.265 ;
      RECT 147.155 -27.248 147.245 -26.24 ;
      RECT 147.105 -26.645 147.245 -26.475 ;
      RECT 147.155 -25.44 147.245 -24.432 ;
      RECT 147.105 -25.205 147.245 -25.035 ;
      RECT 147.155 -24.018 147.245 -23.01 ;
      RECT 147.105 -23.415 147.245 -23.245 ;
      RECT 147.155 -22.21 147.245 -21.202 ;
      RECT 147.105 -21.975 147.245 -21.805 ;
      RECT 147.155 -20.788 147.245 -19.78 ;
      RECT 147.105 -20.185 147.245 -20.015 ;
      RECT 147.155 -18.98 147.245 -17.972 ;
      RECT 147.105 -18.745 147.245 -18.575 ;
      RECT 147.155 -17.558 147.245 -16.55 ;
      RECT 147.105 -16.955 147.245 -16.785 ;
      RECT 147.155 -15.75 147.245 -14.742 ;
      RECT 147.105 -15.515 147.245 -15.345 ;
      RECT 147.155 -14.328 147.245 -13.32 ;
      RECT 147.105 -13.725 147.245 -13.555 ;
      RECT 147.155 -12.52 147.245 -11.512 ;
      RECT 147.105 -12.285 147.245 -12.115 ;
      RECT 147.155 -11.098 147.245 -10.09 ;
      RECT 147.105 -10.495 147.245 -10.325 ;
      RECT 147.155 -9.29 147.245 -8.282 ;
      RECT 147.105 -9.055 147.245 -8.885 ;
      RECT 147.155 -7.868 147.245 -6.86 ;
      RECT 147.105 -7.265 147.245 -7.095 ;
      RECT 147.155 -6.06 147.245 -5.052 ;
      RECT 147.105 -5.825 147.245 -5.655 ;
      RECT 147.155 -4.638 147.245 -3.63 ;
      RECT 147.105 -4.035 147.245 -3.865 ;
      RECT 147.155 -2.83 147.245 -1.822 ;
      RECT 147.105 -2.595 147.245 -2.425 ;
      RECT 147.155 -1.408 147.245 -0.4 ;
      RECT 147.105 -0.805 147.245 -0.635 ;
      RECT 147.155 0.4 147.245 1.408 ;
      RECT 147.105 0.635 147.245 0.805 ;
      RECT 146.755 -101.538 146.845 -100.531 ;
      RECT 146.755 -101.225 146.895 -101.055 ;
      RECT 146.755 -99.729 146.845 -98.722 ;
      RECT 146.755 -99.205 146.895 -99.035 ;
      RECT 146.755 -98.308 146.845 -97.301 ;
      RECT 146.755 -97.995 146.895 -97.825 ;
      RECT 146.755 -96.499 146.845 -95.492 ;
      RECT 146.755 -95.975 146.895 -95.805 ;
      RECT 146.755 -95.078 146.845 -94.071 ;
      RECT 146.755 -94.765 146.895 -94.595 ;
      RECT 146.755 -93.269 146.845 -92.262 ;
      RECT 146.755 -92.745 146.895 -92.575 ;
      RECT 146.755 -91.848 146.845 -90.841 ;
      RECT 146.755 -91.535 146.895 -91.365 ;
      RECT 146.755 -90.039 146.845 -89.032 ;
      RECT 146.755 -89.515 146.895 -89.345 ;
      RECT 146.755 -88.618 146.845 -87.611 ;
      RECT 146.755 -88.305 146.895 -88.135 ;
      RECT 146.755 -86.809 146.845 -85.802 ;
      RECT 146.755 -86.285 146.895 -86.115 ;
      RECT 146.755 -85.388 146.845 -84.381 ;
      RECT 146.755 -85.075 146.895 -84.905 ;
      RECT 146.755 -83.579 146.845 -82.572 ;
      RECT 146.755 -83.055 146.895 -82.885 ;
      RECT 146.755 -82.158 146.845 -81.151 ;
      RECT 146.755 -81.845 146.895 -81.675 ;
      RECT 146.755 -80.349 146.845 -79.342 ;
      RECT 146.755 -79.825 146.895 -79.655 ;
      RECT 146.755 -78.928 146.845 -77.921 ;
      RECT 146.755 -78.615 146.895 -78.445 ;
      RECT 146.755 -77.119 146.845 -76.112 ;
      RECT 146.755 -76.595 146.895 -76.425 ;
      RECT 146.755 -75.698 146.845 -74.691 ;
      RECT 146.755 -75.385 146.895 -75.215 ;
      RECT 146.755 -73.889 146.845 -72.882 ;
      RECT 146.755 -73.365 146.895 -73.195 ;
      RECT 146.755 -72.468 146.845 -71.461 ;
      RECT 146.755 -72.155 146.895 -71.985 ;
      RECT 146.755 -70.659 146.845 -69.652 ;
      RECT 146.755 -70.135 146.895 -69.965 ;
      RECT 146.755 -69.238 146.845 -68.231 ;
      RECT 146.755 -68.925 146.895 -68.755 ;
      RECT 146.755 -67.429 146.845 -66.422 ;
      RECT 146.755 -66.905 146.895 -66.735 ;
      RECT 146.755 -66.008 146.845 -65.001 ;
      RECT 146.755 -65.695 146.895 -65.525 ;
      RECT 146.755 -64.199 146.845 -63.192 ;
      RECT 146.755 -63.675 146.895 -63.505 ;
      RECT 146.755 -62.778 146.845 -61.771 ;
      RECT 146.755 -62.465 146.895 -62.295 ;
      RECT 146.755 -60.969 146.845 -59.962 ;
      RECT 146.755 -60.445 146.895 -60.275 ;
      RECT 146.755 -59.548 146.845 -58.541 ;
      RECT 146.755 -59.235 146.895 -59.065 ;
      RECT 146.755 -57.739 146.845 -56.732 ;
      RECT 146.755 -57.215 146.895 -57.045 ;
      RECT 146.755 -56.318 146.845 -55.311 ;
      RECT 146.755 -56.005 146.895 -55.835 ;
      RECT 146.755 -54.509 146.845 -53.502 ;
      RECT 146.755 -53.985 146.895 -53.815 ;
      RECT 146.755 -53.088 146.845 -52.081 ;
      RECT 146.755 -52.775 146.895 -52.605 ;
      RECT 146.755 -51.279 146.845 -50.272 ;
      RECT 146.755 -50.755 146.895 -50.585 ;
      RECT 146.755 -49.858 146.845 -48.851 ;
      RECT 146.755 -49.545 146.895 -49.375 ;
      RECT 146.755 -48.049 146.845 -47.042 ;
      RECT 146.755 -47.525 146.895 -47.355 ;
      RECT 146.755 -46.628 146.845 -45.621 ;
      RECT 146.755 -46.315 146.895 -46.145 ;
      RECT 146.755 -44.819 146.845 -43.812 ;
      RECT 146.755 -44.295 146.895 -44.125 ;
      RECT 146.755 -43.398 146.845 -42.391 ;
      RECT 146.755 -43.085 146.895 -42.915 ;
      RECT 146.755 -41.589 146.845 -40.582 ;
      RECT 146.755 -41.065 146.895 -40.895 ;
      RECT 146.755 -40.168 146.845 -39.161 ;
      RECT 146.755 -39.855 146.895 -39.685 ;
      RECT 146.755 -38.359 146.845 -37.352 ;
      RECT 146.755 -37.835 146.895 -37.665 ;
      RECT 146.755 -36.938 146.845 -35.931 ;
      RECT 146.755 -36.625 146.895 -36.455 ;
      RECT 146.755 -35.129 146.845 -34.122 ;
      RECT 146.755 -34.605 146.895 -34.435 ;
      RECT 146.755 -33.708 146.845 -32.701 ;
      RECT 146.755 -33.395 146.895 -33.225 ;
      RECT 146.755 -31.899 146.845 -30.892 ;
      RECT 146.755 -31.375 146.895 -31.205 ;
      RECT 146.755 -30.478 146.845 -29.471 ;
      RECT 146.755 -30.165 146.895 -29.995 ;
      RECT 146.755 -28.669 146.845 -27.662 ;
      RECT 146.755 -28.145 146.895 -27.975 ;
      RECT 146.755 -27.248 146.845 -26.241 ;
      RECT 146.755 -26.935 146.895 -26.765 ;
      RECT 146.755 -25.439 146.845 -24.432 ;
      RECT 146.755 -24.915 146.895 -24.745 ;
      RECT 146.755 -24.018 146.845 -23.011 ;
      RECT 146.755 -23.705 146.895 -23.535 ;
      RECT 146.755 -22.209 146.845 -21.202 ;
      RECT 146.755 -21.685 146.895 -21.515 ;
      RECT 146.755 -20.788 146.845 -19.781 ;
      RECT 146.755 -20.475 146.895 -20.305 ;
      RECT 146.755 -18.979 146.845 -17.972 ;
      RECT 146.755 -18.455 146.895 -18.285 ;
      RECT 146.755 -17.558 146.845 -16.551 ;
      RECT 146.755 -17.245 146.895 -17.075 ;
      RECT 146.755 -15.749 146.845 -14.742 ;
      RECT 146.755 -15.225 146.895 -15.055 ;
      RECT 146.755 -14.328 146.845 -13.321 ;
      RECT 146.755 -14.015 146.895 -13.845 ;
      RECT 146.755 -12.519 146.845 -11.512 ;
      RECT 146.755 -11.995 146.895 -11.825 ;
      RECT 146.755 -11.098 146.845 -10.091 ;
      RECT 146.755 -10.785 146.895 -10.615 ;
      RECT 146.755 -9.289 146.845 -8.282 ;
      RECT 146.755 -8.765 146.895 -8.595 ;
      RECT 146.755 -7.868 146.845 -6.861 ;
      RECT 146.755 -7.555 146.895 -7.385 ;
      RECT 146.755 -6.059 146.845 -5.052 ;
      RECT 146.755 -5.535 146.895 -5.365 ;
      RECT 146.755 -4.638 146.845 -3.631 ;
      RECT 146.755 -4.325 146.895 -4.155 ;
      RECT 146.755 -2.829 146.845 -1.822 ;
      RECT 146.755 -2.305 146.895 -2.135 ;
      RECT 146.755 -1.408 146.845 -0.401 ;
      RECT 146.755 -1.095 146.895 -0.925 ;
      RECT 146.755 0.401 146.845 1.408 ;
      RECT 146.755 0.925 146.895 1.095 ;
      RECT 144.905 -111.685 146.385 -111.585 ;
      RECT 144.905 -112.055 145.005 -111.585 ;
      RECT 144.71 -114.395 146.285 -114.275 ;
      RECT 146.185 -114.895 146.285 -114.275 ;
      RECT 145.59 -114.895 145.69 -114.275 ;
      RECT 144.71 -114.85 144.81 -114.275 ;
      RECT 145.955 -101.538 146.045 -100.53 ;
      RECT 145.905 -100.935 146.045 -100.765 ;
      RECT 145.955 -99.73 146.045 -98.722 ;
      RECT 145.905 -99.495 146.045 -99.325 ;
      RECT 145.955 -98.308 146.045 -97.3 ;
      RECT 145.905 -97.705 146.045 -97.535 ;
      RECT 145.955 -96.5 146.045 -95.492 ;
      RECT 145.905 -96.265 146.045 -96.095 ;
      RECT 145.955 -95.078 146.045 -94.07 ;
      RECT 145.905 -94.475 146.045 -94.305 ;
      RECT 145.955 -93.27 146.045 -92.262 ;
      RECT 145.905 -93.035 146.045 -92.865 ;
      RECT 145.955 -91.848 146.045 -90.84 ;
      RECT 145.905 -91.245 146.045 -91.075 ;
      RECT 145.955 -90.04 146.045 -89.032 ;
      RECT 145.905 -89.805 146.045 -89.635 ;
      RECT 145.955 -88.618 146.045 -87.61 ;
      RECT 145.905 -88.015 146.045 -87.845 ;
      RECT 145.955 -86.81 146.045 -85.802 ;
      RECT 145.905 -86.575 146.045 -86.405 ;
      RECT 145.955 -85.388 146.045 -84.38 ;
      RECT 145.905 -84.785 146.045 -84.615 ;
      RECT 145.955 -83.58 146.045 -82.572 ;
      RECT 145.905 -83.345 146.045 -83.175 ;
      RECT 145.955 -82.158 146.045 -81.15 ;
      RECT 145.905 -81.555 146.045 -81.385 ;
      RECT 145.955 -80.35 146.045 -79.342 ;
      RECT 145.905 -80.115 146.045 -79.945 ;
      RECT 145.955 -78.928 146.045 -77.92 ;
      RECT 145.905 -78.325 146.045 -78.155 ;
      RECT 145.955 -77.12 146.045 -76.112 ;
      RECT 145.905 -76.885 146.045 -76.715 ;
      RECT 145.955 -75.698 146.045 -74.69 ;
      RECT 145.905 -75.095 146.045 -74.925 ;
      RECT 145.955 -73.89 146.045 -72.882 ;
      RECT 145.905 -73.655 146.045 -73.485 ;
      RECT 145.955 -72.468 146.045 -71.46 ;
      RECT 145.905 -71.865 146.045 -71.695 ;
      RECT 145.955 -70.66 146.045 -69.652 ;
      RECT 145.905 -70.425 146.045 -70.255 ;
      RECT 145.955 -69.238 146.045 -68.23 ;
      RECT 145.905 -68.635 146.045 -68.465 ;
      RECT 145.955 -67.43 146.045 -66.422 ;
      RECT 145.905 -67.195 146.045 -67.025 ;
      RECT 145.955 -66.008 146.045 -65 ;
      RECT 145.905 -65.405 146.045 -65.235 ;
      RECT 145.955 -64.2 146.045 -63.192 ;
      RECT 145.905 -63.965 146.045 -63.795 ;
      RECT 145.955 -62.778 146.045 -61.77 ;
      RECT 145.905 -62.175 146.045 -62.005 ;
      RECT 145.955 -60.97 146.045 -59.962 ;
      RECT 145.905 -60.735 146.045 -60.565 ;
      RECT 145.955 -59.548 146.045 -58.54 ;
      RECT 145.905 -58.945 146.045 -58.775 ;
      RECT 145.955 -57.74 146.045 -56.732 ;
      RECT 145.905 -57.505 146.045 -57.335 ;
      RECT 145.955 -56.318 146.045 -55.31 ;
      RECT 145.905 -55.715 146.045 -55.545 ;
      RECT 145.955 -54.51 146.045 -53.502 ;
      RECT 145.905 -54.275 146.045 -54.105 ;
      RECT 145.955 -53.088 146.045 -52.08 ;
      RECT 145.905 -52.485 146.045 -52.315 ;
      RECT 145.955 -51.28 146.045 -50.272 ;
      RECT 145.905 -51.045 146.045 -50.875 ;
      RECT 145.955 -49.858 146.045 -48.85 ;
      RECT 145.905 -49.255 146.045 -49.085 ;
      RECT 145.955 -48.05 146.045 -47.042 ;
      RECT 145.905 -47.815 146.045 -47.645 ;
      RECT 145.955 -46.628 146.045 -45.62 ;
      RECT 145.905 -46.025 146.045 -45.855 ;
      RECT 145.955 -44.82 146.045 -43.812 ;
      RECT 145.905 -44.585 146.045 -44.415 ;
      RECT 145.955 -43.398 146.045 -42.39 ;
      RECT 145.905 -42.795 146.045 -42.625 ;
      RECT 145.955 -41.59 146.045 -40.582 ;
      RECT 145.905 -41.355 146.045 -41.185 ;
      RECT 145.955 -40.168 146.045 -39.16 ;
      RECT 145.905 -39.565 146.045 -39.395 ;
      RECT 145.955 -38.36 146.045 -37.352 ;
      RECT 145.905 -38.125 146.045 -37.955 ;
      RECT 145.955 -36.938 146.045 -35.93 ;
      RECT 145.905 -36.335 146.045 -36.165 ;
      RECT 145.955 -35.13 146.045 -34.122 ;
      RECT 145.905 -34.895 146.045 -34.725 ;
      RECT 145.955 -33.708 146.045 -32.7 ;
      RECT 145.905 -33.105 146.045 -32.935 ;
      RECT 145.955 -31.9 146.045 -30.892 ;
      RECT 145.905 -31.665 146.045 -31.495 ;
      RECT 145.955 -30.478 146.045 -29.47 ;
      RECT 145.905 -29.875 146.045 -29.705 ;
      RECT 145.955 -28.67 146.045 -27.662 ;
      RECT 145.905 -28.435 146.045 -28.265 ;
      RECT 145.955 -27.248 146.045 -26.24 ;
      RECT 145.905 -26.645 146.045 -26.475 ;
      RECT 145.955 -25.44 146.045 -24.432 ;
      RECT 145.905 -25.205 146.045 -25.035 ;
      RECT 145.955 -24.018 146.045 -23.01 ;
      RECT 145.905 -23.415 146.045 -23.245 ;
      RECT 145.955 -22.21 146.045 -21.202 ;
      RECT 145.905 -21.975 146.045 -21.805 ;
      RECT 145.955 -20.788 146.045 -19.78 ;
      RECT 145.905 -20.185 146.045 -20.015 ;
      RECT 145.955 -18.98 146.045 -17.972 ;
      RECT 145.905 -18.745 146.045 -18.575 ;
      RECT 145.955 -17.558 146.045 -16.55 ;
      RECT 145.905 -16.955 146.045 -16.785 ;
      RECT 145.955 -15.75 146.045 -14.742 ;
      RECT 145.905 -15.515 146.045 -15.345 ;
      RECT 145.955 -14.328 146.045 -13.32 ;
      RECT 145.905 -13.725 146.045 -13.555 ;
      RECT 145.955 -12.52 146.045 -11.512 ;
      RECT 145.905 -12.285 146.045 -12.115 ;
      RECT 145.955 -11.098 146.045 -10.09 ;
      RECT 145.905 -10.495 146.045 -10.325 ;
      RECT 145.955 -9.29 146.045 -8.282 ;
      RECT 145.905 -9.055 146.045 -8.885 ;
      RECT 145.955 -7.868 146.045 -6.86 ;
      RECT 145.905 -7.265 146.045 -7.095 ;
      RECT 145.955 -6.06 146.045 -5.052 ;
      RECT 145.905 -5.825 146.045 -5.655 ;
      RECT 145.955 -4.638 146.045 -3.63 ;
      RECT 145.905 -4.035 146.045 -3.865 ;
      RECT 145.955 -2.83 146.045 -1.822 ;
      RECT 145.905 -2.595 146.045 -2.425 ;
      RECT 145.955 -1.408 146.045 -0.4 ;
      RECT 145.905 -0.805 146.045 -0.635 ;
      RECT 145.955 0.4 146.045 1.408 ;
      RECT 145.905 0.635 146.045 0.805 ;
      RECT 145.83 -114.685 146.005 -114.515 ;
      RECT 145.905 -114.895 146.005 -114.515 ;
      RECT 144.945 -113.555 145.045 -113.09 ;
      RECT 145.31 -113.555 145.41 -113.1 ;
      RECT 144.945 -113.555 145.79 -113.385 ;
      RECT 145.555 -101.538 145.645 -100.531 ;
      RECT 145.555 -101.225 145.695 -101.055 ;
      RECT 145.555 -99.729 145.645 -98.722 ;
      RECT 145.555 -99.205 145.695 -99.035 ;
      RECT 145.555 -98.308 145.645 -97.301 ;
      RECT 145.555 -97.995 145.695 -97.825 ;
      RECT 145.555 -96.499 145.645 -95.492 ;
      RECT 145.555 -95.975 145.695 -95.805 ;
      RECT 145.555 -95.078 145.645 -94.071 ;
      RECT 145.555 -94.765 145.695 -94.595 ;
      RECT 145.555 -93.269 145.645 -92.262 ;
      RECT 145.555 -92.745 145.695 -92.575 ;
      RECT 145.555 -91.848 145.645 -90.841 ;
      RECT 145.555 -91.535 145.695 -91.365 ;
      RECT 145.555 -90.039 145.645 -89.032 ;
      RECT 145.555 -89.515 145.695 -89.345 ;
      RECT 145.555 -88.618 145.645 -87.611 ;
      RECT 145.555 -88.305 145.695 -88.135 ;
      RECT 145.555 -86.809 145.645 -85.802 ;
      RECT 145.555 -86.285 145.695 -86.115 ;
      RECT 145.555 -85.388 145.645 -84.381 ;
      RECT 145.555 -85.075 145.695 -84.905 ;
      RECT 145.555 -83.579 145.645 -82.572 ;
      RECT 145.555 -83.055 145.695 -82.885 ;
      RECT 145.555 -82.158 145.645 -81.151 ;
      RECT 145.555 -81.845 145.695 -81.675 ;
      RECT 145.555 -80.349 145.645 -79.342 ;
      RECT 145.555 -79.825 145.695 -79.655 ;
      RECT 145.555 -78.928 145.645 -77.921 ;
      RECT 145.555 -78.615 145.695 -78.445 ;
      RECT 145.555 -77.119 145.645 -76.112 ;
      RECT 145.555 -76.595 145.695 -76.425 ;
      RECT 145.555 -75.698 145.645 -74.691 ;
      RECT 145.555 -75.385 145.695 -75.215 ;
      RECT 145.555 -73.889 145.645 -72.882 ;
      RECT 145.555 -73.365 145.695 -73.195 ;
      RECT 145.555 -72.468 145.645 -71.461 ;
      RECT 145.555 -72.155 145.695 -71.985 ;
      RECT 145.555 -70.659 145.645 -69.652 ;
      RECT 145.555 -70.135 145.695 -69.965 ;
      RECT 145.555 -69.238 145.645 -68.231 ;
      RECT 145.555 -68.925 145.695 -68.755 ;
      RECT 145.555 -67.429 145.645 -66.422 ;
      RECT 145.555 -66.905 145.695 -66.735 ;
      RECT 145.555 -66.008 145.645 -65.001 ;
      RECT 145.555 -65.695 145.695 -65.525 ;
      RECT 145.555 -64.199 145.645 -63.192 ;
      RECT 145.555 -63.675 145.695 -63.505 ;
      RECT 145.555 -62.778 145.645 -61.771 ;
      RECT 145.555 -62.465 145.695 -62.295 ;
      RECT 145.555 -60.969 145.645 -59.962 ;
      RECT 145.555 -60.445 145.695 -60.275 ;
      RECT 145.555 -59.548 145.645 -58.541 ;
      RECT 145.555 -59.235 145.695 -59.065 ;
      RECT 145.555 -57.739 145.645 -56.732 ;
      RECT 145.555 -57.215 145.695 -57.045 ;
      RECT 145.555 -56.318 145.645 -55.311 ;
      RECT 145.555 -56.005 145.695 -55.835 ;
      RECT 145.555 -54.509 145.645 -53.502 ;
      RECT 145.555 -53.985 145.695 -53.815 ;
      RECT 145.555 -53.088 145.645 -52.081 ;
      RECT 145.555 -52.775 145.695 -52.605 ;
      RECT 145.555 -51.279 145.645 -50.272 ;
      RECT 145.555 -50.755 145.695 -50.585 ;
      RECT 145.555 -49.858 145.645 -48.851 ;
      RECT 145.555 -49.545 145.695 -49.375 ;
      RECT 145.555 -48.049 145.645 -47.042 ;
      RECT 145.555 -47.525 145.695 -47.355 ;
      RECT 145.555 -46.628 145.645 -45.621 ;
      RECT 145.555 -46.315 145.695 -46.145 ;
      RECT 145.555 -44.819 145.645 -43.812 ;
      RECT 145.555 -44.295 145.695 -44.125 ;
      RECT 145.555 -43.398 145.645 -42.391 ;
      RECT 145.555 -43.085 145.695 -42.915 ;
      RECT 145.555 -41.589 145.645 -40.582 ;
      RECT 145.555 -41.065 145.695 -40.895 ;
      RECT 145.555 -40.168 145.645 -39.161 ;
      RECT 145.555 -39.855 145.695 -39.685 ;
      RECT 145.555 -38.359 145.645 -37.352 ;
      RECT 145.555 -37.835 145.695 -37.665 ;
      RECT 145.555 -36.938 145.645 -35.931 ;
      RECT 145.555 -36.625 145.695 -36.455 ;
      RECT 145.555 -35.129 145.645 -34.122 ;
      RECT 145.555 -34.605 145.695 -34.435 ;
      RECT 145.555 -33.708 145.645 -32.701 ;
      RECT 145.555 -33.395 145.695 -33.225 ;
      RECT 145.555 -31.899 145.645 -30.892 ;
      RECT 145.555 -31.375 145.695 -31.205 ;
      RECT 145.555 -30.478 145.645 -29.471 ;
      RECT 145.555 -30.165 145.695 -29.995 ;
      RECT 145.555 -28.669 145.645 -27.662 ;
      RECT 145.555 -28.145 145.695 -27.975 ;
      RECT 145.555 -27.248 145.645 -26.241 ;
      RECT 145.555 -26.935 145.695 -26.765 ;
      RECT 145.555 -25.439 145.645 -24.432 ;
      RECT 145.555 -24.915 145.695 -24.745 ;
      RECT 145.555 -24.018 145.645 -23.011 ;
      RECT 145.555 -23.705 145.695 -23.535 ;
      RECT 145.555 -22.209 145.645 -21.202 ;
      RECT 145.555 -21.685 145.695 -21.515 ;
      RECT 145.555 -20.788 145.645 -19.781 ;
      RECT 145.555 -20.475 145.695 -20.305 ;
      RECT 145.555 -18.979 145.645 -17.972 ;
      RECT 145.555 -18.455 145.695 -18.285 ;
      RECT 145.555 -17.558 145.645 -16.551 ;
      RECT 145.555 -17.245 145.695 -17.075 ;
      RECT 145.555 -15.749 145.645 -14.742 ;
      RECT 145.555 -15.225 145.695 -15.055 ;
      RECT 145.555 -14.328 145.645 -13.321 ;
      RECT 145.555 -14.015 145.695 -13.845 ;
      RECT 145.555 -12.519 145.645 -11.512 ;
      RECT 145.555 -11.995 145.695 -11.825 ;
      RECT 145.555 -11.098 145.645 -10.091 ;
      RECT 145.555 -10.785 145.695 -10.615 ;
      RECT 145.555 -9.289 145.645 -8.282 ;
      RECT 145.555 -8.765 145.695 -8.595 ;
      RECT 145.555 -7.868 145.645 -6.861 ;
      RECT 145.555 -7.555 145.695 -7.385 ;
      RECT 145.555 -6.059 145.645 -5.052 ;
      RECT 145.555 -5.535 145.695 -5.365 ;
      RECT 145.555 -4.638 145.645 -3.631 ;
      RECT 145.555 -4.325 145.695 -4.155 ;
      RECT 145.555 -2.829 145.645 -1.822 ;
      RECT 145.555 -2.305 145.695 -2.135 ;
      RECT 145.555 -1.408 145.645 -0.401 ;
      RECT 145.555 -1.095 145.695 -0.925 ;
      RECT 145.555 0.401 145.645 1.408 ;
      RECT 145.555 0.925 145.695 1.095 ;
      RECT 145.24 -114.685 145.41 -114.515 ;
      RECT 145.31 -114.895 145.41 -114.515 ;
      RECT 144.755 -101.538 144.845 -100.53 ;
      RECT 144.705 -100.935 144.845 -100.765 ;
      RECT 144.755 -99.73 144.845 -98.722 ;
      RECT 144.705 -99.495 144.845 -99.325 ;
      RECT 144.755 -98.308 144.845 -97.3 ;
      RECT 144.705 -97.705 144.845 -97.535 ;
      RECT 144.755 -96.5 144.845 -95.492 ;
      RECT 144.705 -96.265 144.845 -96.095 ;
      RECT 144.755 -95.078 144.845 -94.07 ;
      RECT 144.705 -94.475 144.845 -94.305 ;
      RECT 144.755 -93.27 144.845 -92.262 ;
      RECT 144.705 -93.035 144.845 -92.865 ;
      RECT 144.755 -91.848 144.845 -90.84 ;
      RECT 144.705 -91.245 144.845 -91.075 ;
      RECT 144.755 -90.04 144.845 -89.032 ;
      RECT 144.705 -89.805 144.845 -89.635 ;
      RECT 144.755 -88.618 144.845 -87.61 ;
      RECT 144.705 -88.015 144.845 -87.845 ;
      RECT 144.755 -86.81 144.845 -85.802 ;
      RECT 144.705 -86.575 144.845 -86.405 ;
      RECT 144.755 -85.388 144.845 -84.38 ;
      RECT 144.705 -84.785 144.845 -84.615 ;
      RECT 144.755 -83.58 144.845 -82.572 ;
      RECT 144.705 -83.345 144.845 -83.175 ;
      RECT 144.755 -82.158 144.845 -81.15 ;
      RECT 144.705 -81.555 144.845 -81.385 ;
      RECT 144.755 -80.35 144.845 -79.342 ;
      RECT 144.705 -80.115 144.845 -79.945 ;
      RECT 144.755 -78.928 144.845 -77.92 ;
      RECT 144.705 -78.325 144.845 -78.155 ;
      RECT 144.755 -77.12 144.845 -76.112 ;
      RECT 144.705 -76.885 144.845 -76.715 ;
      RECT 144.755 -75.698 144.845 -74.69 ;
      RECT 144.705 -75.095 144.845 -74.925 ;
      RECT 144.755 -73.89 144.845 -72.882 ;
      RECT 144.705 -73.655 144.845 -73.485 ;
      RECT 144.755 -72.468 144.845 -71.46 ;
      RECT 144.705 -71.865 144.845 -71.695 ;
      RECT 144.755 -70.66 144.845 -69.652 ;
      RECT 144.705 -70.425 144.845 -70.255 ;
      RECT 144.755 -69.238 144.845 -68.23 ;
      RECT 144.705 -68.635 144.845 -68.465 ;
      RECT 144.755 -67.43 144.845 -66.422 ;
      RECT 144.705 -67.195 144.845 -67.025 ;
      RECT 144.755 -66.008 144.845 -65 ;
      RECT 144.705 -65.405 144.845 -65.235 ;
      RECT 144.755 -64.2 144.845 -63.192 ;
      RECT 144.705 -63.965 144.845 -63.795 ;
      RECT 144.755 -62.778 144.845 -61.77 ;
      RECT 144.705 -62.175 144.845 -62.005 ;
      RECT 144.755 -60.97 144.845 -59.962 ;
      RECT 144.705 -60.735 144.845 -60.565 ;
      RECT 144.755 -59.548 144.845 -58.54 ;
      RECT 144.705 -58.945 144.845 -58.775 ;
      RECT 144.755 -57.74 144.845 -56.732 ;
      RECT 144.705 -57.505 144.845 -57.335 ;
      RECT 144.755 -56.318 144.845 -55.31 ;
      RECT 144.705 -55.715 144.845 -55.545 ;
      RECT 144.755 -54.51 144.845 -53.502 ;
      RECT 144.705 -54.275 144.845 -54.105 ;
      RECT 144.755 -53.088 144.845 -52.08 ;
      RECT 144.705 -52.485 144.845 -52.315 ;
      RECT 144.755 -51.28 144.845 -50.272 ;
      RECT 144.705 -51.045 144.845 -50.875 ;
      RECT 144.755 -49.858 144.845 -48.85 ;
      RECT 144.705 -49.255 144.845 -49.085 ;
      RECT 144.755 -48.05 144.845 -47.042 ;
      RECT 144.705 -47.815 144.845 -47.645 ;
      RECT 144.755 -46.628 144.845 -45.62 ;
      RECT 144.705 -46.025 144.845 -45.855 ;
      RECT 144.755 -44.82 144.845 -43.812 ;
      RECT 144.705 -44.585 144.845 -44.415 ;
      RECT 144.755 -43.398 144.845 -42.39 ;
      RECT 144.705 -42.795 144.845 -42.625 ;
      RECT 144.755 -41.59 144.845 -40.582 ;
      RECT 144.705 -41.355 144.845 -41.185 ;
      RECT 144.755 -40.168 144.845 -39.16 ;
      RECT 144.705 -39.565 144.845 -39.395 ;
      RECT 144.755 -38.36 144.845 -37.352 ;
      RECT 144.705 -38.125 144.845 -37.955 ;
      RECT 144.755 -36.938 144.845 -35.93 ;
      RECT 144.705 -36.335 144.845 -36.165 ;
      RECT 144.755 -35.13 144.845 -34.122 ;
      RECT 144.705 -34.895 144.845 -34.725 ;
      RECT 144.755 -33.708 144.845 -32.7 ;
      RECT 144.705 -33.105 144.845 -32.935 ;
      RECT 144.755 -31.9 144.845 -30.892 ;
      RECT 144.705 -31.665 144.845 -31.495 ;
      RECT 144.755 -30.478 144.845 -29.47 ;
      RECT 144.705 -29.875 144.845 -29.705 ;
      RECT 144.755 -28.67 144.845 -27.662 ;
      RECT 144.705 -28.435 144.845 -28.265 ;
      RECT 144.755 -27.248 144.845 -26.24 ;
      RECT 144.705 -26.645 144.845 -26.475 ;
      RECT 144.755 -25.44 144.845 -24.432 ;
      RECT 144.705 -25.205 144.845 -25.035 ;
      RECT 144.755 -24.018 144.845 -23.01 ;
      RECT 144.705 -23.415 144.845 -23.245 ;
      RECT 144.755 -22.21 144.845 -21.202 ;
      RECT 144.705 -21.975 144.845 -21.805 ;
      RECT 144.755 -20.788 144.845 -19.78 ;
      RECT 144.705 -20.185 144.845 -20.015 ;
      RECT 144.755 -18.98 144.845 -17.972 ;
      RECT 144.705 -18.745 144.845 -18.575 ;
      RECT 144.755 -17.558 144.845 -16.55 ;
      RECT 144.705 -16.955 144.845 -16.785 ;
      RECT 144.755 -15.75 144.845 -14.742 ;
      RECT 144.705 -15.515 144.845 -15.345 ;
      RECT 144.755 -14.328 144.845 -13.32 ;
      RECT 144.705 -13.725 144.845 -13.555 ;
      RECT 144.755 -12.52 144.845 -11.512 ;
      RECT 144.705 -12.285 144.845 -12.115 ;
      RECT 144.755 -11.098 144.845 -10.09 ;
      RECT 144.705 -10.495 144.845 -10.325 ;
      RECT 144.755 -9.29 144.845 -8.282 ;
      RECT 144.705 -9.055 144.845 -8.885 ;
      RECT 144.755 -7.868 144.845 -6.86 ;
      RECT 144.705 -7.265 144.845 -7.095 ;
      RECT 144.755 -6.06 144.845 -5.052 ;
      RECT 144.705 -5.825 144.845 -5.655 ;
      RECT 144.755 -4.638 144.845 -3.63 ;
      RECT 144.705 -4.035 144.845 -3.865 ;
      RECT 144.755 -2.83 144.845 -1.822 ;
      RECT 144.705 -2.595 144.845 -2.425 ;
      RECT 144.755 -1.408 144.845 -0.4 ;
      RECT 144.705 -0.805 144.845 -0.635 ;
      RECT 144.755 0.4 144.845 1.408 ;
      RECT 144.705 0.635 144.845 0.805 ;
      RECT 144.355 -101.538 144.445 -100.531 ;
      RECT 144.355 -101.225 144.495 -101.055 ;
      RECT 144.355 -99.729 144.445 -98.722 ;
      RECT 144.355 -99.205 144.495 -99.035 ;
      RECT 144.355 -98.308 144.445 -97.301 ;
      RECT 144.355 -97.995 144.495 -97.825 ;
      RECT 144.355 -96.499 144.445 -95.492 ;
      RECT 144.355 -95.975 144.495 -95.805 ;
      RECT 144.355 -95.078 144.445 -94.071 ;
      RECT 144.355 -94.765 144.495 -94.595 ;
      RECT 144.355 -93.269 144.445 -92.262 ;
      RECT 144.355 -92.745 144.495 -92.575 ;
      RECT 144.355 -91.848 144.445 -90.841 ;
      RECT 144.355 -91.535 144.495 -91.365 ;
      RECT 144.355 -90.039 144.445 -89.032 ;
      RECT 144.355 -89.515 144.495 -89.345 ;
      RECT 144.355 -88.618 144.445 -87.611 ;
      RECT 144.355 -88.305 144.495 -88.135 ;
      RECT 144.355 -86.809 144.445 -85.802 ;
      RECT 144.355 -86.285 144.495 -86.115 ;
      RECT 144.355 -85.388 144.445 -84.381 ;
      RECT 144.355 -85.075 144.495 -84.905 ;
      RECT 144.355 -83.579 144.445 -82.572 ;
      RECT 144.355 -83.055 144.495 -82.885 ;
      RECT 144.355 -82.158 144.445 -81.151 ;
      RECT 144.355 -81.845 144.495 -81.675 ;
      RECT 144.355 -80.349 144.445 -79.342 ;
      RECT 144.355 -79.825 144.495 -79.655 ;
      RECT 144.355 -78.928 144.445 -77.921 ;
      RECT 144.355 -78.615 144.495 -78.445 ;
      RECT 144.355 -77.119 144.445 -76.112 ;
      RECT 144.355 -76.595 144.495 -76.425 ;
      RECT 144.355 -75.698 144.445 -74.691 ;
      RECT 144.355 -75.385 144.495 -75.215 ;
      RECT 144.355 -73.889 144.445 -72.882 ;
      RECT 144.355 -73.365 144.495 -73.195 ;
      RECT 144.355 -72.468 144.445 -71.461 ;
      RECT 144.355 -72.155 144.495 -71.985 ;
      RECT 144.355 -70.659 144.445 -69.652 ;
      RECT 144.355 -70.135 144.495 -69.965 ;
      RECT 144.355 -69.238 144.445 -68.231 ;
      RECT 144.355 -68.925 144.495 -68.755 ;
      RECT 144.355 -67.429 144.445 -66.422 ;
      RECT 144.355 -66.905 144.495 -66.735 ;
      RECT 144.355 -66.008 144.445 -65.001 ;
      RECT 144.355 -65.695 144.495 -65.525 ;
      RECT 144.355 -64.199 144.445 -63.192 ;
      RECT 144.355 -63.675 144.495 -63.505 ;
      RECT 144.355 -62.778 144.445 -61.771 ;
      RECT 144.355 -62.465 144.495 -62.295 ;
      RECT 144.355 -60.969 144.445 -59.962 ;
      RECT 144.355 -60.445 144.495 -60.275 ;
      RECT 144.355 -59.548 144.445 -58.541 ;
      RECT 144.355 -59.235 144.495 -59.065 ;
      RECT 144.355 -57.739 144.445 -56.732 ;
      RECT 144.355 -57.215 144.495 -57.045 ;
      RECT 144.355 -56.318 144.445 -55.311 ;
      RECT 144.355 -56.005 144.495 -55.835 ;
      RECT 144.355 -54.509 144.445 -53.502 ;
      RECT 144.355 -53.985 144.495 -53.815 ;
      RECT 144.355 -53.088 144.445 -52.081 ;
      RECT 144.355 -52.775 144.495 -52.605 ;
      RECT 144.355 -51.279 144.445 -50.272 ;
      RECT 144.355 -50.755 144.495 -50.585 ;
      RECT 144.355 -49.858 144.445 -48.851 ;
      RECT 144.355 -49.545 144.495 -49.375 ;
      RECT 144.355 -48.049 144.445 -47.042 ;
      RECT 144.355 -47.525 144.495 -47.355 ;
      RECT 144.355 -46.628 144.445 -45.621 ;
      RECT 144.355 -46.315 144.495 -46.145 ;
      RECT 144.355 -44.819 144.445 -43.812 ;
      RECT 144.355 -44.295 144.495 -44.125 ;
      RECT 144.355 -43.398 144.445 -42.391 ;
      RECT 144.355 -43.085 144.495 -42.915 ;
      RECT 144.355 -41.589 144.445 -40.582 ;
      RECT 144.355 -41.065 144.495 -40.895 ;
      RECT 144.355 -40.168 144.445 -39.161 ;
      RECT 144.355 -39.855 144.495 -39.685 ;
      RECT 144.355 -38.359 144.445 -37.352 ;
      RECT 144.355 -37.835 144.495 -37.665 ;
      RECT 144.355 -36.938 144.445 -35.931 ;
      RECT 144.355 -36.625 144.495 -36.455 ;
      RECT 144.355 -35.129 144.445 -34.122 ;
      RECT 144.355 -34.605 144.495 -34.435 ;
      RECT 144.355 -33.708 144.445 -32.701 ;
      RECT 144.355 -33.395 144.495 -33.225 ;
      RECT 144.355 -31.899 144.445 -30.892 ;
      RECT 144.355 -31.375 144.495 -31.205 ;
      RECT 144.355 -30.478 144.445 -29.471 ;
      RECT 144.355 -30.165 144.495 -29.995 ;
      RECT 144.355 -28.669 144.445 -27.662 ;
      RECT 144.355 -28.145 144.495 -27.975 ;
      RECT 144.355 -27.248 144.445 -26.241 ;
      RECT 144.355 -26.935 144.495 -26.765 ;
      RECT 144.355 -25.439 144.445 -24.432 ;
      RECT 144.355 -24.915 144.495 -24.745 ;
      RECT 144.355 -24.018 144.445 -23.011 ;
      RECT 144.355 -23.705 144.495 -23.535 ;
      RECT 144.355 -22.209 144.445 -21.202 ;
      RECT 144.355 -21.685 144.495 -21.515 ;
      RECT 144.355 -20.788 144.445 -19.781 ;
      RECT 144.355 -20.475 144.495 -20.305 ;
      RECT 144.355 -18.979 144.445 -17.972 ;
      RECT 144.355 -18.455 144.495 -18.285 ;
      RECT 144.355 -17.558 144.445 -16.551 ;
      RECT 144.355 -17.245 144.495 -17.075 ;
      RECT 144.355 -15.749 144.445 -14.742 ;
      RECT 144.355 -15.225 144.495 -15.055 ;
      RECT 144.355 -14.328 144.445 -13.321 ;
      RECT 144.355 -14.015 144.495 -13.845 ;
      RECT 144.355 -12.519 144.445 -11.512 ;
      RECT 144.355 -11.995 144.495 -11.825 ;
      RECT 144.355 -11.098 144.445 -10.091 ;
      RECT 144.355 -10.785 144.495 -10.615 ;
      RECT 144.355 -9.289 144.445 -8.282 ;
      RECT 144.355 -8.765 144.495 -8.595 ;
      RECT 144.355 -7.868 144.445 -6.861 ;
      RECT 144.355 -7.555 144.495 -7.385 ;
      RECT 144.355 -6.059 144.445 -5.052 ;
      RECT 144.355 -5.535 144.495 -5.365 ;
      RECT 144.355 -4.638 144.445 -3.631 ;
      RECT 144.355 -4.325 144.495 -4.155 ;
      RECT 144.355 -2.829 144.445 -1.822 ;
      RECT 144.355 -2.305 144.495 -2.135 ;
      RECT 144.355 -1.408 144.445 -0.401 ;
      RECT 144.355 -1.095 144.495 -0.925 ;
      RECT 144.355 0.401 144.445 1.408 ;
      RECT 144.355 0.925 144.495 1.095 ;
      RECT 140.185 -108.935 143.965 -108.815 ;
      RECT 141.505 -109.475 141.605 -108.815 ;
      RECT 140.945 -109.475 141.045 -108.815 ;
      RECT 140.385 -109.475 140.485 -108.815 ;
      RECT 143.555 -101.538 143.645 -100.53 ;
      RECT 143.505 -100.935 143.645 -100.765 ;
      RECT 143.555 -99.73 143.645 -98.722 ;
      RECT 143.505 -99.495 143.645 -99.325 ;
      RECT 143.555 -98.308 143.645 -97.3 ;
      RECT 143.505 -97.705 143.645 -97.535 ;
      RECT 143.555 -96.5 143.645 -95.492 ;
      RECT 143.505 -96.265 143.645 -96.095 ;
      RECT 143.555 -95.078 143.645 -94.07 ;
      RECT 143.505 -94.475 143.645 -94.305 ;
      RECT 143.555 -93.27 143.645 -92.262 ;
      RECT 143.505 -93.035 143.645 -92.865 ;
      RECT 143.555 -91.848 143.645 -90.84 ;
      RECT 143.505 -91.245 143.645 -91.075 ;
      RECT 143.555 -90.04 143.645 -89.032 ;
      RECT 143.505 -89.805 143.645 -89.635 ;
      RECT 143.555 -88.618 143.645 -87.61 ;
      RECT 143.505 -88.015 143.645 -87.845 ;
      RECT 143.555 -86.81 143.645 -85.802 ;
      RECT 143.505 -86.575 143.645 -86.405 ;
      RECT 143.555 -85.388 143.645 -84.38 ;
      RECT 143.505 -84.785 143.645 -84.615 ;
      RECT 143.555 -83.58 143.645 -82.572 ;
      RECT 143.505 -83.345 143.645 -83.175 ;
      RECT 143.555 -82.158 143.645 -81.15 ;
      RECT 143.505 -81.555 143.645 -81.385 ;
      RECT 143.555 -80.35 143.645 -79.342 ;
      RECT 143.505 -80.115 143.645 -79.945 ;
      RECT 143.555 -78.928 143.645 -77.92 ;
      RECT 143.505 -78.325 143.645 -78.155 ;
      RECT 143.555 -77.12 143.645 -76.112 ;
      RECT 143.505 -76.885 143.645 -76.715 ;
      RECT 143.555 -75.698 143.645 -74.69 ;
      RECT 143.505 -75.095 143.645 -74.925 ;
      RECT 143.555 -73.89 143.645 -72.882 ;
      RECT 143.505 -73.655 143.645 -73.485 ;
      RECT 143.555 -72.468 143.645 -71.46 ;
      RECT 143.505 -71.865 143.645 -71.695 ;
      RECT 143.555 -70.66 143.645 -69.652 ;
      RECT 143.505 -70.425 143.645 -70.255 ;
      RECT 143.555 -69.238 143.645 -68.23 ;
      RECT 143.505 -68.635 143.645 -68.465 ;
      RECT 143.555 -67.43 143.645 -66.422 ;
      RECT 143.505 -67.195 143.645 -67.025 ;
      RECT 143.555 -66.008 143.645 -65 ;
      RECT 143.505 -65.405 143.645 -65.235 ;
      RECT 143.555 -64.2 143.645 -63.192 ;
      RECT 143.505 -63.965 143.645 -63.795 ;
      RECT 143.555 -62.778 143.645 -61.77 ;
      RECT 143.505 -62.175 143.645 -62.005 ;
      RECT 143.555 -60.97 143.645 -59.962 ;
      RECT 143.505 -60.735 143.645 -60.565 ;
      RECT 143.555 -59.548 143.645 -58.54 ;
      RECT 143.505 -58.945 143.645 -58.775 ;
      RECT 143.555 -57.74 143.645 -56.732 ;
      RECT 143.505 -57.505 143.645 -57.335 ;
      RECT 143.555 -56.318 143.645 -55.31 ;
      RECT 143.505 -55.715 143.645 -55.545 ;
      RECT 143.555 -54.51 143.645 -53.502 ;
      RECT 143.505 -54.275 143.645 -54.105 ;
      RECT 143.555 -53.088 143.645 -52.08 ;
      RECT 143.505 -52.485 143.645 -52.315 ;
      RECT 143.555 -51.28 143.645 -50.272 ;
      RECT 143.505 -51.045 143.645 -50.875 ;
      RECT 143.555 -49.858 143.645 -48.85 ;
      RECT 143.505 -49.255 143.645 -49.085 ;
      RECT 143.555 -48.05 143.645 -47.042 ;
      RECT 143.505 -47.815 143.645 -47.645 ;
      RECT 143.555 -46.628 143.645 -45.62 ;
      RECT 143.505 -46.025 143.645 -45.855 ;
      RECT 143.555 -44.82 143.645 -43.812 ;
      RECT 143.505 -44.585 143.645 -44.415 ;
      RECT 143.555 -43.398 143.645 -42.39 ;
      RECT 143.505 -42.795 143.645 -42.625 ;
      RECT 143.555 -41.59 143.645 -40.582 ;
      RECT 143.505 -41.355 143.645 -41.185 ;
      RECT 143.555 -40.168 143.645 -39.16 ;
      RECT 143.505 -39.565 143.645 -39.395 ;
      RECT 143.555 -38.36 143.645 -37.352 ;
      RECT 143.505 -38.125 143.645 -37.955 ;
      RECT 143.555 -36.938 143.645 -35.93 ;
      RECT 143.505 -36.335 143.645 -36.165 ;
      RECT 143.555 -35.13 143.645 -34.122 ;
      RECT 143.505 -34.895 143.645 -34.725 ;
      RECT 143.555 -33.708 143.645 -32.7 ;
      RECT 143.505 -33.105 143.645 -32.935 ;
      RECT 143.555 -31.9 143.645 -30.892 ;
      RECT 143.505 -31.665 143.645 -31.495 ;
      RECT 143.555 -30.478 143.645 -29.47 ;
      RECT 143.505 -29.875 143.645 -29.705 ;
      RECT 143.555 -28.67 143.645 -27.662 ;
      RECT 143.505 -28.435 143.645 -28.265 ;
      RECT 143.555 -27.248 143.645 -26.24 ;
      RECT 143.505 -26.645 143.645 -26.475 ;
      RECT 143.555 -25.44 143.645 -24.432 ;
      RECT 143.505 -25.205 143.645 -25.035 ;
      RECT 143.555 -24.018 143.645 -23.01 ;
      RECT 143.505 -23.415 143.645 -23.245 ;
      RECT 143.555 -22.21 143.645 -21.202 ;
      RECT 143.505 -21.975 143.645 -21.805 ;
      RECT 143.555 -20.788 143.645 -19.78 ;
      RECT 143.505 -20.185 143.645 -20.015 ;
      RECT 143.555 -18.98 143.645 -17.972 ;
      RECT 143.505 -18.745 143.645 -18.575 ;
      RECT 143.555 -17.558 143.645 -16.55 ;
      RECT 143.505 -16.955 143.645 -16.785 ;
      RECT 143.555 -15.75 143.645 -14.742 ;
      RECT 143.505 -15.515 143.645 -15.345 ;
      RECT 143.555 -14.328 143.645 -13.32 ;
      RECT 143.505 -13.725 143.645 -13.555 ;
      RECT 143.555 -12.52 143.645 -11.512 ;
      RECT 143.505 -12.285 143.645 -12.115 ;
      RECT 143.555 -11.098 143.645 -10.09 ;
      RECT 143.505 -10.495 143.645 -10.325 ;
      RECT 143.555 -9.29 143.645 -8.282 ;
      RECT 143.505 -9.055 143.645 -8.885 ;
      RECT 143.555 -7.868 143.645 -6.86 ;
      RECT 143.505 -7.265 143.645 -7.095 ;
      RECT 143.555 -6.06 143.645 -5.052 ;
      RECT 143.505 -5.825 143.645 -5.655 ;
      RECT 143.555 -4.638 143.645 -3.63 ;
      RECT 143.505 -4.035 143.645 -3.865 ;
      RECT 143.555 -2.83 143.645 -1.822 ;
      RECT 143.505 -2.595 143.645 -2.425 ;
      RECT 143.555 -1.408 143.645 -0.4 ;
      RECT 143.505 -0.805 143.645 -0.635 ;
      RECT 143.555 0.4 143.645 1.408 ;
      RECT 143.505 0.635 143.645 0.805 ;
      RECT 142.125 -111.685 143.605 -111.585 ;
      RECT 142.125 -112.195 142.225 -111.585 ;
      RECT 142.345 -109.15 143.605 -109.05 ;
      RECT 143.505 -109.475 143.605 -109.05 ;
      RECT 142.945 -109.475 143.045 -109.05 ;
      RECT 142.385 -109.475 142.485 -109.05 ;
      RECT 143.155 -101.538 143.245 -100.531 ;
      RECT 143.155 -101.225 143.295 -101.055 ;
      RECT 143.155 -99.729 143.245 -98.722 ;
      RECT 143.155 -99.205 143.295 -99.035 ;
      RECT 143.155 -98.308 143.245 -97.301 ;
      RECT 143.155 -97.995 143.295 -97.825 ;
      RECT 143.155 -96.499 143.245 -95.492 ;
      RECT 143.155 -95.975 143.295 -95.805 ;
      RECT 143.155 -95.078 143.245 -94.071 ;
      RECT 143.155 -94.765 143.295 -94.595 ;
      RECT 143.155 -93.269 143.245 -92.262 ;
      RECT 143.155 -92.745 143.295 -92.575 ;
      RECT 143.155 -91.848 143.245 -90.841 ;
      RECT 143.155 -91.535 143.295 -91.365 ;
      RECT 143.155 -90.039 143.245 -89.032 ;
      RECT 143.155 -89.515 143.295 -89.345 ;
      RECT 143.155 -88.618 143.245 -87.611 ;
      RECT 143.155 -88.305 143.295 -88.135 ;
      RECT 143.155 -86.809 143.245 -85.802 ;
      RECT 143.155 -86.285 143.295 -86.115 ;
      RECT 143.155 -85.388 143.245 -84.381 ;
      RECT 143.155 -85.075 143.295 -84.905 ;
      RECT 143.155 -83.579 143.245 -82.572 ;
      RECT 143.155 -83.055 143.295 -82.885 ;
      RECT 143.155 -82.158 143.245 -81.151 ;
      RECT 143.155 -81.845 143.295 -81.675 ;
      RECT 143.155 -80.349 143.245 -79.342 ;
      RECT 143.155 -79.825 143.295 -79.655 ;
      RECT 143.155 -78.928 143.245 -77.921 ;
      RECT 143.155 -78.615 143.295 -78.445 ;
      RECT 143.155 -77.119 143.245 -76.112 ;
      RECT 143.155 -76.595 143.295 -76.425 ;
      RECT 143.155 -75.698 143.245 -74.691 ;
      RECT 143.155 -75.385 143.295 -75.215 ;
      RECT 143.155 -73.889 143.245 -72.882 ;
      RECT 143.155 -73.365 143.295 -73.195 ;
      RECT 143.155 -72.468 143.245 -71.461 ;
      RECT 143.155 -72.155 143.295 -71.985 ;
      RECT 143.155 -70.659 143.245 -69.652 ;
      RECT 143.155 -70.135 143.295 -69.965 ;
      RECT 143.155 -69.238 143.245 -68.231 ;
      RECT 143.155 -68.925 143.295 -68.755 ;
      RECT 143.155 -67.429 143.245 -66.422 ;
      RECT 143.155 -66.905 143.295 -66.735 ;
      RECT 143.155 -66.008 143.245 -65.001 ;
      RECT 143.155 -65.695 143.295 -65.525 ;
      RECT 143.155 -64.199 143.245 -63.192 ;
      RECT 143.155 -63.675 143.295 -63.505 ;
      RECT 143.155 -62.778 143.245 -61.771 ;
      RECT 143.155 -62.465 143.295 -62.295 ;
      RECT 143.155 -60.969 143.245 -59.962 ;
      RECT 143.155 -60.445 143.295 -60.275 ;
      RECT 143.155 -59.548 143.245 -58.541 ;
      RECT 143.155 -59.235 143.295 -59.065 ;
      RECT 143.155 -57.739 143.245 -56.732 ;
      RECT 143.155 -57.215 143.295 -57.045 ;
      RECT 143.155 -56.318 143.245 -55.311 ;
      RECT 143.155 -56.005 143.295 -55.835 ;
      RECT 143.155 -54.509 143.245 -53.502 ;
      RECT 143.155 -53.985 143.295 -53.815 ;
      RECT 143.155 -53.088 143.245 -52.081 ;
      RECT 143.155 -52.775 143.295 -52.605 ;
      RECT 143.155 -51.279 143.245 -50.272 ;
      RECT 143.155 -50.755 143.295 -50.585 ;
      RECT 143.155 -49.858 143.245 -48.851 ;
      RECT 143.155 -49.545 143.295 -49.375 ;
      RECT 143.155 -48.049 143.245 -47.042 ;
      RECT 143.155 -47.525 143.295 -47.355 ;
      RECT 143.155 -46.628 143.245 -45.621 ;
      RECT 143.155 -46.315 143.295 -46.145 ;
      RECT 143.155 -44.819 143.245 -43.812 ;
      RECT 143.155 -44.295 143.295 -44.125 ;
      RECT 143.155 -43.398 143.245 -42.391 ;
      RECT 143.155 -43.085 143.295 -42.915 ;
      RECT 143.155 -41.589 143.245 -40.582 ;
      RECT 143.155 -41.065 143.295 -40.895 ;
      RECT 143.155 -40.168 143.245 -39.161 ;
      RECT 143.155 -39.855 143.295 -39.685 ;
      RECT 143.155 -38.359 143.245 -37.352 ;
      RECT 143.155 -37.835 143.295 -37.665 ;
      RECT 143.155 -36.938 143.245 -35.931 ;
      RECT 143.155 -36.625 143.295 -36.455 ;
      RECT 143.155 -35.129 143.245 -34.122 ;
      RECT 143.155 -34.605 143.295 -34.435 ;
      RECT 143.155 -33.708 143.245 -32.701 ;
      RECT 143.155 -33.395 143.295 -33.225 ;
      RECT 143.155 -31.899 143.245 -30.892 ;
      RECT 143.155 -31.375 143.295 -31.205 ;
      RECT 143.155 -30.478 143.245 -29.471 ;
      RECT 143.155 -30.165 143.295 -29.995 ;
      RECT 143.155 -28.669 143.245 -27.662 ;
      RECT 143.155 -28.145 143.295 -27.975 ;
      RECT 143.155 -27.248 143.245 -26.241 ;
      RECT 143.155 -26.935 143.295 -26.765 ;
      RECT 143.155 -25.439 143.245 -24.432 ;
      RECT 143.155 -24.915 143.295 -24.745 ;
      RECT 143.155 -24.018 143.245 -23.011 ;
      RECT 143.155 -23.705 143.295 -23.535 ;
      RECT 143.155 -22.209 143.245 -21.202 ;
      RECT 143.155 -21.685 143.295 -21.515 ;
      RECT 143.155 -20.788 143.245 -19.781 ;
      RECT 143.155 -20.475 143.295 -20.305 ;
      RECT 143.155 -18.979 143.245 -17.972 ;
      RECT 143.155 -18.455 143.295 -18.285 ;
      RECT 143.155 -17.558 143.245 -16.551 ;
      RECT 143.155 -17.245 143.295 -17.075 ;
      RECT 143.155 -15.749 143.245 -14.742 ;
      RECT 143.155 -15.225 143.295 -15.055 ;
      RECT 143.155 -14.328 143.245 -13.321 ;
      RECT 143.155 -14.015 143.295 -13.845 ;
      RECT 143.155 -12.519 143.245 -11.512 ;
      RECT 143.155 -11.995 143.295 -11.825 ;
      RECT 143.155 -11.098 143.245 -10.091 ;
      RECT 143.155 -10.785 143.295 -10.615 ;
      RECT 143.155 -9.289 143.245 -8.282 ;
      RECT 143.155 -8.765 143.295 -8.595 ;
      RECT 143.155 -7.868 143.245 -6.861 ;
      RECT 143.155 -7.555 143.295 -7.385 ;
      RECT 143.155 -6.059 143.245 -5.052 ;
      RECT 143.155 -5.535 143.295 -5.365 ;
      RECT 143.155 -4.638 143.245 -3.631 ;
      RECT 143.155 -4.325 143.295 -4.155 ;
      RECT 143.155 -2.829 143.245 -1.822 ;
      RECT 143.155 -2.305 143.295 -2.135 ;
      RECT 143.155 -1.408 143.245 -0.401 ;
      RECT 143.155 -1.095 143.295 -0.925 ;
      RECT 143.155 0.401 143.245 1.408 ;
      RECT 143.155 0.925 143.295 1.095 ;
      RECT 142.485 -111.495 142.655 -111.385 ;
      RECT 139.335 -111.495 142.655 -111.395 ;
      RECT 142.355 -101.538 142.445 -100.53 ;
      RECT 142.305 -100.935 142.445 -100.765 ;
      RECT 142.355 -99.73 142.445 -98.722 ;
      RECT 142.305 -99.495 142.445 -99.325 ;
      RECT 142.355 -98.308 142.445 -97.3 ;
      RECT 142.305 -97.705 142.445 -97.535 ;
      RECT 142.355 -96.5 142.445 -95.492 ;
      RECT 142.305 -96.265 142.445 -96.095 ;
      RECT 142.355 -95.078 142.445 -94.07 ;
      RECT 142.305 -94.475 142.445 -94.305 ;
      RECT 142.355 -93.27 142.445 -92.262 ;
      RECT 142.305 -93.035 142.445 -92.865 ;
      RECT 142.355 -91.848 142.445 -90.84 ;
      RECT 142.305 -91.245 142.445 -91.075 ;
      RECT 142.355 -90.04 142.445 -89.032 ;
      RECT 142.305 -89.805 142.445 -89.635 ;
      RECT 142.355 -88.618 142.445 -87.61 ;
      RECT 142.305 -88.015 142.445 -87.845 ;
      RECT 142.355 -86.81 142.445 -85.802 ;
      RECT 142.305 -86.575 142.445 -86.405 ;
      RECT 142.355 -85.388 142.445 -84.38 ;
      RECT 142.305 -84.785 142.445 -84.615 ;
      RECT 142.355 -83.58 142.445 -82.572 ;
      RECT 142.305 -83.345 142.445 -83.175 ;
      RECT 142.355 -82.158 142.445 -81.15 ;
      RECT 142.305 -81.555 142.445 -81.385 ;
      RECT 142.355 -80.35 142.445 -79.342 ;
      RECT 142.305 -80.115 142.445 -79.945 ;
      RECT 142.355 -78.928 142.445 -77.92 ;
      RECT 142.305 -78.325 142.445 -78.155 ;
      RECT 142.355 -77.12 142.445 -76.112 ;
      RECT 142.305 -76.885 142.445 -76.715 ;
      RECT 142.355 -75.698 142.445 -74.69 ;
      RECT 142.305 -75.095 142.445 -74.925 ;
      RECT 142.355 -73.89 142.445 -72.882 ;
      RECT 142.305 -73.655 142.445 -73.485 ;
      RECT 142.355 -72.468 142.445 -71.46 ;
      RECT 142.305 -71.865 142.445 -71.695 ;
      RECT 142.355 -70.66 142.445 -69.652 ;
      RECT 142.305 -70.425 142.445 -70.255 ;
      RECT 142.355 -69.238 142.445 -68.23 ;
      RECT 142.305 -68.635 142.445 -68.465 ;
      RECT 142.355 -67.43 142.445 -66.422 ;
      RECT 142.305 -67.195 142.445 -67.025 ;
      RECT 142.355 -66.008 142.445 -65 ;
      RECT 142.305 -65.405 142.445 -65.235 ;
      RECT 142.355 -64.2 142.445 -63.192 ;
      RECT 142.305 -63.965 142.445 -63.795 ;
      RECT 142.355 -62.778 142.445 -61.77 ;
      RECT 142.305 -62.175 142.445 -62.005 ;
      RECT 142.355 -60.97 142.445 -59.962 ;
      RECT 142.305 -60.735 142.445 -60.565 ;
      RECT 142.355 -59.548 142.445 -58.54 ;
      RECT 142.305 -58.945 142.445 -58.775 ;
      RECT 142.355 -57.74 142.445 -56.732 ;
      RECT 142.305 -57.505 142.445 -57.335 ;
      RECT 142.355 -56.318 142.445 -55.31 ;
      RECT 142.305 -55.715 142.445 -55.545 ;
      RECT 142.355 -54.51 142.445 -53.502 ;
      RECT 142.305 -54.275 142.445 -54.105 ;
      RECT 142.355 -53.088 142.445 -52.08 ;
      RECT 142.305 -52.485 142.445 -52.315 ;
      RECT 142.355 -51.28 142.445 -50.272 ;
      RECT 142.305 -51.045 142.445 -50.875 ;
      RECT 142.355 -49.858 142.445 -48.85 ;
      RECT 142.305 -49.255 142.445 -49.085 ;
      RECT 142.355 -48.05 142.445 -47.042 ;
      RECT 142.305 -47.815 142.445 -47.645 ;
      RECT 142.355 -46.628 142.445 -45.62 ;
      RECT 142.305 -46.025 142.445 -45.855 ;
      RECT 142.355 -44.82 142.445 -43.812 ;
      RECT 142.305 -44.585 142.445 -44.415 ;
      RECT 142.355 -43.398 142.445 -42.39 ;
      RECT 142.305 -42.795 142.445 -42.625 ;
      RECT 142.355 -41.59 142.445 -40.582 ;
      RECT 142.305 -41.355 142.445 -41.185 ;
      RECT 142.355 -40.168 142.445 -39.16 ;
      RECT 142.305 -39.565 142.445 -39.395 ;
      RECT 142.355 -38.36 142.445 -37.352 ;
      RECT 142.305 -38.125 142.445 -37.955 ;
      RECT 142.355 -36.938 142.445 -35.93 ;
      RECT 142.305 -36.335 142.445 -36.165 ;
      RECT 142.355 -35.13 142.445 -34.122 ;
      RECT 142.305 -34.895 142.445 -34.725 ;
      RECT 142.355 -33.708 142.445 -32.7 ;
      RECT 142.305 -33.105 142.445 -32.935 ;
      RECT 142.355 -31.9 142.445 -30.892 ;
      RECT 142.305 -31.665 142.445 -31.495 ;
      RECT 142.355 -30.478 142.445 -29.47 ;
      RECT 142.305 -29.875 142.445 -29.705 ;
      RECT 142.355 -28.67 142.445 -27.662 ;
      RECT 142.305 -28.435 142.445 -28.265 ;
      RECT 142.355 -27.248 142.445 -26.24 ;
      RECT 142.305 -26.645 142.445 -26.475 ;
      RECT 142.355 -25.44 142.445 -24.432 ;
      RECT 142.305 -25.205 142.445 -25.035 ;
      RECT 142.355 -24.018 142.445 -23.01 ;
      RECT 142.305 -23.415 142.445 -23.245 ;
      RECT 142.355 -22.21 142.445 -21.202 ;
      RECT 142.305 -21.975 142.445 -21.805 ;
      RECT 142.355 -20.788 142.445 -19.78 ;
      RECT 142.305 -20.185 142.445 -20.015 ;
      RECT 142.355 -18.98 142.445 -17.972 ;
      RECT 142.305 -18.745 142.445 -18.575 ;
      RECT 142.355 -17.558 142.445 -16.55 ;
      RECT 142.305 -16.955 142.445 -16.785 ;
      RECT 142.355 -15.75 142.445 -14.742 ;
      RECT 142.305 -15.515 142.445 -15.345 ;
      RECT 142.355 -14.328 142.445 -13.32 ;
      RECT 142.305 -13.725 142.445 -13.555 ;
      RECT 142.355 -12.52 142.445 -11.512 ;
      RECT 142.305 -12.285 142.445 -12.115 ;
      RECT 142.355 -11.098 142.445 -10.09 ;
      RECT 142.305 -10.495 142.445 -10.325 ;
      RECT 142.355 -9.29 142.445 -8.282 ;
      RECT 142.305 -9.055 142.445 -8.885 ;
      RECT 142.355 -7.868 142.445 -6.86 ;
      RECT 142.305 -7.265 142.445 -7.095 ;
      RECT 142.355 -6.06 142.445 -5.052 ;
      RECT 142.305 -5.825 142.445 -5.655 ;
      RECT 142.355 -4.638 142.445 -3.63 ;
      RECT 142.305 -4.035 142.445 -3.865 ;
      RECT 142.355 -2.83 142.445 -1.822 ;
      RECT 142.305 -2.595 142.445 -2.425 ;
      RECT 142.355 -1.408 142.445 -0.4 ;
      RECT 142.305 -0.805 142.445 -0.635 ;
      RECT 142.355 0.4 142.445 1.408 ;
      RECT 142.305 0.635 142.445 0.805 ;
      RECT 141.955 -101.538 142.045 -100.531 ;
      RECT 141.955 -101.225 142.095 -101.055 ;
      RECT 141.955 -99.729 142.045 -98.722 ;
      RECT 141.955 -99.205 142.095 -99.035 ;
      RECT 141.955 -98.308 142.045 -97.301 ;
      RECT 141.955 -97.995 142.095 -97.825 ;
      RECT 141.955 -96.499 142.045 -95.492 ;
      RECT 141.955 -95.975 142.095 -95.805 ;
      RECT 141.955 -95.078 142.045 -94.071 ;
      RECT 141.955 -94.765 142.095 -94.595 ;
      RECT 141.955 -93.269 142.045 -92.262 ;
      RECT 141.955 -92.745 142.095 -92.575 ;
      RECT 141.955 -91.848 142.045 -90.841 ;
      RECT 141.955 -91.535 142.095 -91.365 ;
      RECT 141.955 -90.039 142.045 -89.032 ;
      RECT 141.955 -89.515 142.095 -89.345 ;
      RECT 141.955 -88.618 142.045 -87.611 ;
      RECT 141.955 -88.305 142.095 -88.135 ;
      RECT 141.955 -86.809 142.045 -85.802 ;
      RECT 141.955 -86.285 142.095 -86.115 ;
      RECT 141.955 -85.388 142.045 -84.381 ;
      RECT 141.955 -85.075 142.095 -84.905 ;
      RECT 141.955 -83.579 142.045 -82.572 ;
      RECT 141.955 -83.055 142.095 -82.885 ;
      RECT 141.955 -82.158 142.045 -81.151 ;
      RECT 141.955 -81.845 142.095 -81.675 ;
      RECT 141.955 -80.349 142.045 -79.342 ;
      RECT 141.955 -79.825 142.095 -79.655 ;
      RECT 141.955 -78.928 142.045 -77.921 ;
      RECT 141.955 -78.615 142.095 -78.445 ;
      RECT 141.955 -77.119 142.045 -76.112 ;
      RECT 141.955 -76.595 142.095 -76.425 ;
      RECT 141.955 -75.698 142.045 -74.691 ;
      RECT 141.955 -75.385 142.095 -75.215 ;
      RECT 141.955 -73.889 142.045 -72.882 ;
      RECT 141.955 -73.365 142.095 -73.195 ;
      RECT 141.955 -72.468 142.045 -71.461 ;
      RECT 141.955 -72.155 142.095 -71.985 ;
      RECT 141.955 -70.659 142.045 -69.652 ;
      RECT 141.955 -70.135 142.095 -69.965 ;
      RECT 141.955 -69.238 142.045 -68.231 ;
      RECT 141.955 -68.925 142.095 -68.755 ;
      RECT 141.955 -67.429 142.045 -66.422 ;
      RECT 141.955 -66.905 142.095 -66.735 ;
      RECT 141.955 -66.008 142.045 -65.001 ;
      RECT 141.955 -65.695 142.095 -65.525 ;
      RECT 141.955 -64.199 142.045 -63.192 ;
      RECT 141.955 -63.675 142.095 -63.505 ;
      RECT 141.955 -62.778 142.045 -61.771 ;
      RECT 141.955 -62.465 142.095 -62.295 ;
      RECT 141.955 -60.969 142.045 -59.962 ;
      RECT 141.955 -60.445 142.095 -60.275 ;
      RECT 141.955 -59.548 142.045 -58.541 ;
      RECT 141.955 -59.235 142.095 -59.065 ;
      RECT 141.955 -57.739 142.045 -56.732 ;
      RECT 141.955 -57.215 142.095 -57.045 ;
      RECT 141.955 -56.318 142.045 -55.311 ;
      RECT 141.955 -56.005 142.095 -55.835 ;
      RECT 141.955 -54.509 142.045 -53.502 ;
      RECT 141.955 -53.985 142.095 -53.815 ;
      RECT 141.955 -53.088 142.045 -52.081 ;
      RECT 141.955 -52.775 142.095 -52.605 ;
      RECT 141.955 -51.279 142.045 -50.272 ;
      RECT 141.955 -50.755 142.095 -50.585 ;
      RECT 141.955 -49.858 142.045 -48.851 ;
      RECT 141.955 -49.545 142.095 -49.375 ;
      RECT 141.955 -48.049 142.045 -47.042 ;
      RECT 141.955 -47.525 142.095 -47.355 ;
      RECT 141.955 -46.628 142.045 -45.621 ;
      RECT 141.955 -46.315 142.095 -46.145 ;
      RECT 141.955 -44.819 142.045 -43.812 ;
      RECT 141.955 -44.295 142.095 -44.125 ;
      RECT 141.955 -43.398 142.045 -42.391 ;
      RECT 141.955 -43.085 142.095 -42.915 ;
      RECT 141.955 -41.589 142.045 -40.582 ;
      RECT 141.955 -41.065 142.095 -40.895 ;
      RECT 141.955 -40.168 142.045 -39.161 ;
      RECT 141.955 -39.855 142.095 -39.685 ;
      RECT 141.955 -38.359 142.045 -37.352 ;
      RECT 141.955 -37.835 142.095 -37.665 ;
      RECT 141.955 -36.938 142.045 -35.931 ;
      RECT 141.955 -36.625 142.095 -36.455 ;
      RECT 141.955 -35.129 142.045 -34.122 ;
      RECT 141.955 -34.605 142.095 -34.435 ;
      RECT 141.955 -33.708 142.045 -32.701 ;
      RECT 141.955 -33.395 142.095 -33.225 ;
      RECT 141.955 -31.899 142.045 -30.892 ;
      RECT 141.955 -31.375 142.095 -31.205 ;
      RECT 141.955 -30.478 142.045 -29.471 ;
      RECT 141.955 -30.165 142.095 -29.995 ;
      RECT 141.955 -28.669 142.045 -27.662 ;
      RECT 141.955 -28.145 142.095 -27.975 ;
      RECT 141.955 -27.248 142.045 -26.241 ;
      RECT 141.955 -26.935 142.095 -26.765 ;
      RECT 141.955 -25.439 142.045 -24.432 ;
      RECT 141.955 -24.915 142.095 -24.745 ;
      RECT 141.955 -24.018 142.045 -23.011 ;
      RECT 141.955 -23.705 142.095 -23.535 ;
      RECT 141.955 -22.209 142.045 -21.202 ;
      RECT 141.955 -21.685 142.095 -21.515 ;
      RECT 141.955 -20.788 142.045 -19.781 ;
      RECT 141.955 -20.475 142.095 -20.305 ;
      RECT 141.955 -18.979 142.045 -17.972 ;
      RECT 141.955 -18.455 142.095 -18.285 ;
      RECT 141.955 -17.558 142.045 -16.551 ;
      RECT 141.955 -17.245 142.095 -17.075 ;
      RECT 141.955 -15.749 142.045 -14.742 ;
      RECT 141.955 -15.225 142.095 -15.055 ;
      RECT 141.955 -14.328 142.045 -13.321 ;
      RECT 141.955 -14.015 142.095 -13.845 ;
      RECT 141.955 -12.519 142.045 -11.512 ;
      RECT 141.955 -11.995 142.095 -11.825 ;
      RECT 141.955 -11.098 142.045 -10.091 ;
      RECT 141.955 -10.785 142.095 -10.615 ;
      RECT 141.955 -9.289 142.045 -8.282 ;
      RECT 141.955 -8.765 142.095 -8.595 ;
      RECT 141.955 -7.868 142.045 -6.861 ;
      RECT 141.955 -7.555 142.095 -7.385 ;
      RECT 141.955 -6.059 142.045 -5.052 ;
      RECT 141.955 -5.535 142.095 -5.365 ;
      RECT 141.955 -4.638 142.045 -3.631 ;
      RECT 141.955 -4.325 142.095 -4.155 ;
      RECT 141.955 -2.829 142.045 -1.822 ;
      RECT 141.955 -2.305 142.095 -2.135 ;
      RECT 141.955 -1.408 142.045 -0.401 ;
      RECT 141.955 -1.095 142.095 -0.925 ;
      RECT 141.955 0.401 142.045 1.408 ;
      RECT 141.955 0.925 142.095 1.095 ;
      RECT 140.105 -111.685 141.585 -111.585 ;
      RECT 140.105 -112.055 140.205 -111.585 ;
      RECT 139.91 -114.395 141.485 -114.275 ;
      RECT 141.385 -114.895 141.485 -114.275 ;
      RECT 140.79 -114.895 140.89 -114.275 ;
      RECT 139.91 -114.85 140.01 -114.275 ;
      RECT 141.155 -101.538 141.245 -100.53 ;
      RECT 141.105 -100.935 141.245 -100.765 ;
      RECT 141.155 -99.73 141.245 -98.722 ;
      RECT 141.105 -99.495 141.245 -99.325 ;
      RECT 141.155 -98.308 141.245 -97.3 ;
      RECT 141.105 -97.705 141.245 -97.535 ;
      RECT 141.155 -96.5 141.245 -95.492 ;
      RECT 141.105 -96.265 141.245 -96.095 ;
      RECT 141.155 -95.078 141.245 -94.07 ;
      RECT 141.105 -94.475 141.245 -94.305 ;
      RECT 141.155 -93.27 141.245 -92.262 ;
      RECT 141.105 -93.035 141.245 -92.865 ;
      RECT 141.155 -91.848 141.245 -90.84 ;
      RECT 141.105 -91.245 141.245 -91.075 ;
      RECT 141.155 -90.04 141.245 -89.032 ;
      RECT 141.105 -89.805 141.245 -89.635 ;
      RECT 141.155 -88.618 141.245 -87.61 ;
      RECT 141.105 -88.015 141.245 -87.845 ;
      RECT 141.155 -86.81 141.245 -85.802 ;
      RECT 141.105 -86.575 141.245 -86.405 ;
      RECT 141.155 -85.388 141.245 -84.38 ;
      RECT 141.105 -84.785 141.245 -84.615 ;
      RECT 141.155 -83.58 141.245 -82.572 ;
      RECT 141.105 -83.345 141.245 -83.175 ;
      RECT 141.155 -82.158 141.245 -81.15 ;
      RECT 141.105 -81.555 141.245 -81.385 ;
      RECT 141.155 -80.35 141.245 -79.342 ;
      RECT 141.105 -80.115 141.245 -79.945 ;
      RECT 141.155 -78.928 141.245 -77.92 ;
      RECT 141.105 -78.325 141.245 -78.155 ;
      RECT 141.155 -77.12 141.245 -76.112 ;
      RECT 141.105 -76.885 141.245 -76.715 ;
      RECT 141.155 -75.698 141.245 -74.69 ;
      RECT 141.105 -75.095 141.245 -74.925 ;
      RECT 141.155 -73.89 141.245 -72.882 ;
      RECT 141.105 -73.655 141.245 -73.485 ;
      RECT 141.155 -72.468 141.245 -71.46 ;
      RECT 141.105 -71.865 141.245 -71.695 ;
      RECT 141.155 -70.66 141.245 -69.652 ;
      RECT 141.105 -70.425 141.245 -70.255 ;
      RECT 141.155 -69.238 141.245 -68.23 ;
      RECT 141.105 -68.635 141.245 -68.465 ;
      RECT 141.155 -67.43 141.245 -66.422 ;
      RECT 141.105 -67.195 141.245 -67.025 ;
      RECT 141.155 -66.008 141.245 -65 ;
      RECT 141.105 -65.405 141.245 -65.235 ;
      RECT 141.155 -64.2 141.245 -63.192 ;
      RECT 141.105 -63.965 141.245 -63.795 ;
      RECT 141.155 -62.778 141.245 -61.77 ;
      RECT 141.105 -62.175 141.245 -62.005 ;
      RECT 141.155 -60.97 141.245 -59.962 ;
      RECT 141.105 -60.735 141.245 -60.565 ;
      RECT 141.155 -59.548 141.245 -58.54 ;
      RECT 141.105 -58.945 141.245 -58.775 ;
      RECT 141.155 -57.74 141.245 -56.732 ;
      RECT 141.105 -57.505 141.245 -57.335 ;
      RECT 141.155 -56.318 141.245 -55.31 ;
      RECT 141.105 -55.715 141.245 -55.545 ;
      RECT 141.155 -54.51 141.245 -53.502 ;
      RECT 141.105 -54.275 141.245 -54.105 ;
      RECT 141.155 -53.088 141.245 -52.08 ;
      RECT 141.105 -52.485 141.245 -52.315 ;
      RECT 141.155 -51.28 141.245 -50.272 ;
      RECT 141.105 -51.045 141.245 -50.875 ;
      RECT 141.155 -49.858 141.245 -48.85 ;
      RECT 141.105 -49.255 141.245 -49.085 ;
      RECT 141.155 -48.05 141.245 -47.042 ;
      RECT 141.105 -47.815 141.245 -47.645 ;
      RECT 141.155 -46.628 141.245 -45.62 ;
      RECT 141.105 -46.025 141.245 -45.855 ;
      RECT 141.155 -44.82 141.245 -43.812 ;
      RECT 141.105 -44.585 141.245 -44.415 ;
      RECT 141.155 -43.398 141.245 -42.39 ;
      RECT 141.105 -42.795 141.245 -42.625 ;
      RECT 141.155 -41.59 141.245 -40.582 ;
      RECT 141.105 -41.355 141.245 -41.185 ;
      RECT 141.155 -40.168 141.245 -39.16 ;
      RECT 141.105 -39.565 141.245 -39.395 ;
      RECT 141.155 -38.36 141.245 -37.352 ;
      RECT 141.105 -38.125 141.245 -37.955 ;
      RECT 141.155 -36.938 141.245 -35.93 ;
      RECT 141.105 -36.335 141.245 -36.165 ;
      RECT 141.155 -35.13 141.245 -34.122 ;
      RECT 141.105 -34.895 141.245 -34.725 ;
      RECT 141.155 -33.708 141.245 -32.7 ;
      RECT 141.105 -33.105 141.245 -32.935 ;
      RECT 141.155 -31.9 141.245 -30.892 ;
      RECT 141.105 -31.665 141.245 -31.495 ;
      RECT 141.155 -30.478 141.245 -29.47 ;
      RECT 141.105 -29.875 141.245 -29.705 ;
      RECT 141.155 -28.67 141.245 -27.662 ;
      RECT 141.105 -28.435 141.245 -28.265 ;
      RECT 141.155 -27.248 141.245 -26.24 ;
      RECT 141.105 -26.645 141.245 -26.475 ;
      RECT 141.155 -25.44 141.245 -24.432 ;
      RECT 141.105 -25.205 141.245 -25.035 ;
      RECT 141.155 -24.018 141.245 -23.01 ;
      RECT 141.105 -23.415 141.245 -23.245 ;
      RECT 141.155 -22.21 141.245 -21.202 ;
      RECT 141.105 -21.975 141.245 -21.805 ;
      RECT 141.155 -20.788 141.245 -19.78 ;
      RECT 141.105 -20.185 141.245 -20.015 ;
      RECT 141.155 -18.98 141.245 -17.972 ;
      RECT 141.105 -18.745 141.245 -18.575 ;
      RECT 141.155 -17.558 141.245 -16.55 ;
      RECT 141.105 -16.955 141.245 -16.785 ;
      RECT 141.155 -15.75 141.245 -14.742 ;
      RECT 141.105 -15.515 141.245 -15.345 ;
      RECT 141.155 -14.328 141.245 -13.32 ;
      RECT 141.105 -13.725 141.245 -13.555 ;
      RECT 141.155 -12.52 141.245 -11.512 ;
      RECT 141.105 -12.285 141.245 -12.115 ;
      RECT 141.155 -11.098 141.245 -10.09 ;
      RECT 141.105 -10.495 141.245 -10.325 ;
      RECT 141.155 -9.29 141.245 -8.282 ;
      RECT 141.105 -9.055 141.245 -8.885 ;
      RECT 141.155 -7.868 141.245 -6.86 ;
      RECT 141.105 -7.265 141.245 -7.095 ;
      RECT 141.155 -6.06 141.245 -5.052 ;
      RECT 141.105 -5.825 141.245 -5.655 ;
      RECT 141.155 -4.638 141.245 -3.63 ;
      RECT 141.105 -4.035 141.245 -3.865 ;
      RECT 141.155 -2.83 141.245 -1.822 ;
      RECT 141.105 -2.595 141.245 -2.425 ;
      RECT 141.155 -1.408 141.245 -0.4 ;
      RECT 141.105 -0.805 141.245 -0.635 ;
      RECT 141.155 0.4 141.245 1.408 ;
      RECT 141.105 0.635 141.245 0.805 ;
      RECT 141.03 -114.685 141.205 -114.515 ;
      RECT 141.105 -114.895 141.205 -114.515 ;
      RECT 140.145 -113.555 140.245 -113.09 ;
      RECT 140.51 -113.555 140.61 -113.1 ;
      RECT 140.145 -113.555 140.99 -113.385 ;
      RECT 140.755 -101.538 140.845 -100.531 ;
      RECT 140.755 -101.225 140.895 -101.055 ;
      RECT 140.755 -99.729 140.845 -98.722 ;
      RECT 140.755 -99.205 140.895 -99.035 ;
      RECT 140.755 -98.308 140.845 -97.301 ;
      RECT 140.755 -97.995 140.895 -97.825 ;
      RECT 140.755 -96.499 140.845 -95.492 ;
      RECT 140.755 -95.975 140.895 -95.805 ;
      RECT 140.755 -95.078 140.845 -94.071 ;
      RECT 140.755 -94.765 140.895 -94.595 ;
      RECT 140.755 -93.269 140.845 -92.262 ;
      RECT 140.755 -92.745 140.895 -92.575 ;
      RECT 140.755 -91.848 140.845 -90.841 ;
      RECT 140.755 -91.535 140.895 -91.365 ;
      RECT 140.755 -90.039 140.845 -89.032 ;
      RECT 140.755 -89.515 140.895 -89.345 ;
      RECT 140.755 -88.618 140.845 -87.611 ;
      RECT 140.755 -88.305 140.895 -88.135 ;
      RECT 140.755 -86.809 140.845 -85.802 ;
      RECT 140.755 -86.285 140.895 -86.115 ;
      RECT 140.755 -85.388 140.845 -84.381 ;
      RECT 140.755 -85.075 140.895 -84.905 ;
      RECT 140.755 -83.579 140.845 -82.572 ;
      RECT 140.755 -83.055 140.895 -82.885 ;
      RECT 140.755 -82.158 140.845 -81.151 ;
      RECT 140.755 -81.845 140.895 -81.675 ;
      RECT 140.755 -80.349 140.845 -79.342 ;
      RECT 140.755 -79.825 140.895 -79.655 ;
      RECT 140.755 -78.928 140.845 -77.921 ;
      RECT 140.755 -78.615 140.895 -78.445 ;
      RECT 140.755 -77.119 140.845 -76.112 ;
      RECT 140.755 -76.595 140.895 -76.425 ;
      RECT 140.755 -75.698 140.845 -74.691 ;
      RECT 140.755 -75.385 140.895 -75.215 ;
      RECT 140.755 -73.889 140.845 -72.882 ;
      RECT 140.755 -73.365 140.895 -73.195 ;
      RECT 140.755 -72.468 140.845 -71.461 ;
      RECT 140.755 -72.155 140.895 -71.985 ;
      RECT 140.755 -70.659 140.845 -69.652 ;
      RECT 140.755 -70.135 140.895 -69.965 ;
      RECT 140.755 -69.238 140.845 -68.231 ;
      RECT 140.755 -68.925 140.895 -68.755 ;
      RECT 140.755 -67.429 140.845 -66.422 ;
      RECT 140.755 -66.905 140.895 -66.735 ;
      RECT 140.755 -66.008 140.845 -65.001 ;
      RECT 140.755 -65.695 140.895 -65.525 ;
      RECT 140.755 -64.199 140.845 -63.192 ;
      RECT 140.755 -63.675 140.895 -63.505 ;
      RECT 140.755 -62.778 140.845 -61.771 ;
      RECT 140.755 -62.465 140.895 -62.295 ;
      RECT 140.755 -60.969 140.845 -59.962 ;
      RECT 140.755 -60.445 140.895 -60.275 ;
      RECT 140.755 -59.548 140.845 -58.541 ;
      RECT 140.755 -59.235 140.895 -59.065 ;
      RECT 140.755 -57.739 140.845 -56.732 ;
      RECT 140.755 -57.215 140.895 -57.045 ;
      RECT 140.755 -56.318 140.845 -55.311 ;
      RECT 140.755 -56.005 140.895 -55.835 ;
      RECT 140.755 -54.509 140.845 -53.502 ;
      RECT 140.755 -53.985 140.895 -53.815 ;
      RECT 140.755 -53.088 140.845 -52.081 ;
      RECT 140.755 -52.775 140.895 -52.605 ;
      RECT 140.755 -51.279 140.845 -50.272 ;
      RECT 140.755 -50.755 140.895 -50.585 ;
      RECT 140.755 -49.858 140.845 -48.851 ;
      RECT 140.755 -49.545 140.895 -49.375 ;
      RECT 140.755 -48.049 140.845 -47.042 ;
      RECT 140.755 -47.525 140.895 -47.355 ;
      RECT 140.755 -46.628 140.845 -45.621 ;
      RECT 140.755 -46.315 140.895 -46.145 ;
      RECT 140.755 -44.819 140.845 -43.812 ;
      RECT 140.755 -44.295 140.895 -44.125 ;
      RECT 140.755 -43.398 140.845 -42.391 ;
      RECT 140.755 -43.085 140.895 -42.915 ;
      RECT 140.755 -41.589 140.845 -40.582 ;
      RECT 140.755 -41.065 140.895 -40.895 ;
      RECT 140.755 -40.168 140.845 -39.161 ;
      RECT 140.755 -39.855 140.895 -39.685 ;
      RECT 140.755 -38.359 140.845 -37.352 ;
      RECT 140.755 -37.835 140.895 -37.665 ;
      RECT 140.755 -36.938 140.845 -35.931 ;
      RECT 140.755 -36.625 140.895 -36.455 ;
      RECT 140.755 -35.129 140.845 -34.122 ;
      RECT 140.755 -34.605 140.895 -34.435 ;
      RECT 140.755 -33.708 140.845 -32.701 ;
      RECT 140.755 -33.395 140.895 -33.225 ;
      RECT 140.755 -31.899 140.845 -30.892 ;
      RECT 140.755 -31.375 140.895 -31.205 ;
      RECT 140.755 -30.478 140.845 -29.471 ;
      RECT 140.755 -30.165 140.895 -29.995 ;
      RECT 140.755 -28.669 140.845 -27.662 ;
      RECT 140.755 -28.145 140.895 -27.975 ;
      RECT 140.755 -27.248 140.845 -26.241 ;
      RECT 140.755 -26.935 140.895 -26.765 ;
      RECT 140.755 -25.439 140.845 -24.432 ;
      RECT 140.755 -24.915 140.895 -24.745 ;
      RECT 140.755 -24.018 140.845 -23.011 ;
      RECT 140.755 -23.705 140.895 -23.535 ;
      RECT 140.755 -22.209 140.845 -21.202 ;
      RECT 140.755 -21.685 140.895 -21.515 ;
      RECT 140.755 -20.788 140.845 -19.781 ;
      RECT 140.755 -20.475 140.895 -20.305 ;
      RECT 140.755 -18.979 140.845 -17.972 ;
      RECT 140.755 -18.455 140.895 -18.285 ;
      RECT 140.755 -17.558 140.845 -16.551 ;
      RECT 140.755 -17.245 140.895 -17.075 ;
      RECT 140.755 -15.749 140.845 -14.742 ;
      RECT 140.755 -15.225 140.895 -15.055 ;
      RECT 140.755 -14.328 140.845 -13.321 ;
      RECT 140.755 -14.015 140.895 -13.845 ;
      RECT 140.755 -12.519 140.845 -11.512 ;
      RECT 140.755 -11.995 140.895 -11.825 ;
      RECT 140.755 -11.098 140.845 -10.091 ;
      RECT 140.755 -10.785 140.895 -10.615 ;
      RECT 140.755 -9.289 140.845 -8.282 ;
      RECT 140.755 -8.765 140.895 -8.595 ;
      RECT 140.755 -7.868 140.845 -6.861 ;
      RECT 140.755 -7.555 140.895 -7.385 ;
      RECT 140.755 -6.059 140.845 -5.052 ;
      RECT 140.755 -5.535 140.895 -5.365 ;
      RECT 140.755 -4.638 140.845 -3.631 ;
      RECT 140.755 -4.325 140.895 -4.155 ;
      RECT 140.755 -2.829 140.845 -1.822 ;
      RECT 140.755 -2.305 140.895 -2.135 ;
      RECT 140.755 -1.408 140.845 -0.401 ;
      RECT 140.755 -1.095 140.895 -0.925 ;
      RECT 140.755 0.401 140.845 1.408 ;
      RECT 140.755 0.925 140.895 1.095 ;
      RECT 140.44 -114.685 140.61 -114.515 ;
      RECT 140.51 -114.895 140.61 -114.515 ;
      RECT 139.955 -101.538 140.045 -100.53 ;
      RECT 139.905 -100.935 140.045 -100.765 ;
      RECT 139.955 -99.73 140.045 -98.722 ;
      RECT 139.905 -99.495 140.045 -99.325 ;
      RECT 139.955 -98.308 140.045 -97.3 ;
      RECT 139.905 -97.705 140.045 -97.535 ;
      RECT 139.955 -96.5 140.045 -95.492 ;
      RECT 139.905 -96.265 140.045 -96.095 ;
      RECT 139.955 -95.078 140.045 -94.07 ;
      RECT 139.905 -94.475 140.045 -94.305 ;
      RECT 139.955 -93.27 140.045 -92.262 ;
      RECT 139.905 -93.035 140.045 -92.865 ;
      RECT 139.955 -91.848 140.045 -90.84 ;
      RECT 139.905 -91.245 140.045 -91.075 ;
      RECT 139.955 -90.04 140.045 -89.032 ;
      RECT 139.905 -89.805 140.045 -89.635 ;
      RECT 139.955 -88.618 140.045 -87.61 ;
      RECT 139.905 -88.015 140.045 -87.845 ;
      RECT 139.955 -86.81 140.045 -85.802 ;
      RECT 139.905 -86.575 140.045 -86.405 ;
      RECT 139.955 -85.388 140.045 -84.38 ;
      RECT 139.905 -84.785 140.045 -84.615 ;
      RECT 139.955 -83.58 140.045 -82.572 ;
      RECT 139.905 -83.345 140.045 -83.175 ;
      RECT 139.955 -82.158 140.045 -81.15 ;
      RECT 139.905 -81.555 140.045 -81.385 ;
      RECT 139.955 -80.35 140.045 -79.342 ;
      RECT 139.905 -80.115 140.045 -79.945 ;
      RECT 139.955 -78.928 140.045 -77.92 ;
      RECT 139.905 -78.325 140.045 -78.155 ;
      RECT 139.955 -77.12 140.045 -76.112 ;
      RECT 139.905 -76.885 140.045 -76.715 ;
      RECT 139.955 -75.698 140.045 -74.69 ;
      RECT 139.905 -75.095 140.045 -74.925 ;
      RECT 139.955 -73.89 140.045 -72.882 ;
      RECT 139.905 -73.655 140.045 -73.485 ;
      RECT 139.955 -72.468 140.045 -71.46 ;
      RECT 139.905 -71.865 140.045 -71.695 ;
      RECT 139.955 -70.66 140.045 -69.652 ;
      RECT 139.905 -70.425 140.045 -70.255 ;
      RECT 139.955 -69.238 140.045 -68.23 ;
      RECT 139.905 -68.635 140.045 -68.465 ;
      RECT 139.955 -67.43 140.045 -66.422 ;
      RECT 139.905 -67.195 140.045 -67.025 ;
      RECT 139.955 -66.008 140.045 -65 ;
      RECT 139.905 -65.405 140.045 -65.235 ;
      RECT 139.955 -64.2 140.045 -63.192 ;
      RECT 139.905 -63.965 140.045 -63.795 ;
      RECT 139.955 -62.778 140.045 -61.77 ;
      RECT 139.905 -62.175 140.045 -62.005 ;
      RECT 139.955 -60.97 140.045 -59.962 ;
      RECT 139.905 -60.735 140.045 -60.565 ;
      RECT 139.955 -59.548 140.045 -58.54 ;
      RECT 139.905 -58.945 140.045 -58.775 ;
      RECT 139.955 -57.74 140.045 -56.732 ;
      RECT 139.905 -57.505 140.045 -57.335 ;
      RECT 139.955 -56.318 140.045 -55.31 ;
      RECT 139.905 -55.715 140.045 -55.545 ;
      RECT 139.955 -54.51 140.045 -53.502 ;
      RECT 139.905 -54.275 140.045 -54.105 ;
      RECT 139.955 -53.088 140.045 -52.08 ;
      RECT 139.905 -52.485 140.045 -52.315 ;
      RECT 139.955 -51.28 140.045 -50.272 ;
      RECT 139.905 -51.045 140.045 -50.875 ;
      RECT 139.955 -49.858 140.045 -48.85 ;
      RECT 139.905 -49.255 140.045 -49.085 ;
      RECT 139.955 -48.05 140.045 -47.042 ;
      RECT 139.905 -47.815 140.045 -47.645 ;
      RECT 139.955 -46.628 140.045 -45.62 ;
      RECT 139.905 -46.025 140.045 -45.855 ;
      RECT 139.955 -44.82 140.045 -43.812 ;
      RECT 139.905 -44.585 140.045 -44.415 ;
      RECT 139.955 -43.398 140.045 -42.39 ;
      RECT 139.905 -42.795 140.045 -42.625 ;
      RECT 139.955 -41.59 140.045 -40.582 ;
      RECT 139.905 -41.355 140.045 -41.185 ;
      RECT 139.955 -40.168 140.045 -39.16 ;
      RECT 139.905 -39.565 140.045 -39.395 ;
      RECT 139.955 -38.36 140.045 -37.352 ;
      RECT 139.905 -38.125 140.045 -37.955 ;
      RECT 139.955 -36.938 140.045 -35.93 ;
      RECT 139.905 -36.335 140.045 -36.165 ;
      RECT 139.955 -35.13 140.045 -34.122 ;
      RECT 139.905 -34.895 140.045 -34.725 ;
      RECT 139.955 -33.708 140.045 -32.7 ;
      RECT 139.905 -33.105 140.045 -32.935 ;
      RECT 139.955 -31.9 140.045 -30.892 ;
      RECT 139.905 -31.665 140.045 -31.495 ;
      RECT 139.955 -30.478 140.045 -29.47 ;
      RECT 139.905 -29.875 140.045 -29.705 ;
      RECT 139.955 -28.67 140.045 -27.662 ;
      RECT 139.905 -28.435 140.045 -28.265 ;
      RECT 139.955 -27.248 140.045 -26.24 ;
      RECT 139.905 -26.645 140.045 -26.475 ;
      RECT 139.955 -25.44 140.045 -24.432 ;
      RECT 139.905 -25.205 140.045 -25.035 ;
      RECT 139.955 -24.018 140.045 -23.01 ;
      RECT 139.905 -23.415 140.045 -23.245 ;
      RECT 139.955 -22.21 140.045 -21.202 ;
      RECT 139.905 -21.975 140.045 -21.805 ;
      RECT 139.955 -20.788 140.045 -19.78 ;
      RECT 139.905 -20.185 140.045 -20.015 ;
      RECT 139.955 -18.98 140.045 -17.972 ;
      RECT 139.905 -18.745 140.045 -18.575 ;
      RECT 139.955 -17.558 140.045 -16.55 ;
      RECT 139.905 -16.955 140.045 -16.785 ;
      RECT 139.955 -15.75 140.045 -14.742 ;
      RECT 139.905 -15.515 140.045 -15.345 ;
      RECT 139.955 -14.328 140.045 -13.32 ;
      RECT 139.905 -13.725 140.045 -13.555 ;
      RECT 139.955 -12.52 140.045 -11.512 ;
      RECT 139.905 -12.285 140.045 -12.115 ;
      RECT 139.955 -11.098 140.045 -10.09 ;
      RECT 139.905 -10.495 140.045 -10.325 ;
      RECT 139.955 -9.29 140.045 -8.282 ;
      RECT 139.905 -9.055 140.045 -8.885 ;
      RECT 139.955 -7.868 140.045 -6.86 ;
      RECT 139.905 -7.265 140.045 -7.095 ;
      RECT 139.955 -6.06 140.045 -5.052 ;
      RECT 139.905 -5.825 140.045 -5.655 ;
      RECT 139.955 -4.638 140.045 -3.63 ;
      RECT 139.905 -4.035 140.045 -3.865 ;
      RECT 139.955 -2.83 140.045 -1.822 ;
      RECT 139.905 -2.595 140.045 -2.425 ;
      RECT 139.955 -1.408 140.045 -0.4 ;
      RECT 139.905 -0.805 140.045 -0.635 ;
      RECT 139.955 0.4 140.045 1.408 ;
      RECT 139.905 0.635 140.045 0.805 ;
      RECT 139.555 -101.538 139.645 -100.531 ;
      RECT 139.555 -101.225 139.695 -101.055 ;
      RECT 139.555 -99.729 139.645 -98.722 ;
      RECT 139.555 -99.205 139.695 -99.035 ;
      RECT 139.555 -98.308 139.645 -97.301 ;
      RECT 139.555 -97.995 139.695 -97.825 ;
      RECT 139.555 -96.499 139.645 -95.492 ;
      RECT 139.555 -95.975 139.695 -95.805 ;
      RECT 139.555 -95.078 139.645 -94.071 ;
      RECT 139.555 -94.765 139.695 -94.595 ;
      RECT 139.555 -93.269 139.645 -92.262 ;
      RECT 139.555 -92.745 139.695 -92.575 ;
      RECT 139.555 -91.848 139.645 -90.841 ;
      RECT 139.555 -91.535 139.695 -91.365 ;
      RECT 139.555 -90.039 139.645 -89.032 ;
      RECT 139.555 -89.515 139.695 -89.345 ;
      RECT 139.555 -88.618 139.645 -87.611 ;
      RECT 139.555 -88.305 139.695 -88.135 ;
      RECT 139.555 -86.809 139.645 -85.802 ;
      RECT 139.555 -86.285 139.695 -86.115 ;
      RECT 139.555 -85.388 139.645 -84.381 ;
      RECT 139.555 -85.075 139.695 -84.905 ;
      RECT 139.555 -83.579 139.645 -82.572 ;
      RECT 139.555 -83.055 139.695 -82.885 ;
      RECT 139.555 -82.158 139.645 -81.151 ;
      RECT 139.555 -81.845 139.695 -81.675 ;
      RECT 139.555 -80.349 139.645 -79.342 ;
      RECT 139.555 -79.825 139.695 -79.655 ;
      RECT 139.555 -78.928 139.645 -77.921 ;
      RECT 139.555 -78.615 139.695 -78.445 ;
      RECT 139.555 -77.119 139.645 -76.112 ;
      RECT 139.555 -76.595 139.695 -76.425 ;
      RECT 139.555 -75.698 139.645 -74.691 ;
      RECT 139.555 -75.385 139.695 -75.215 ;
      RECT 139.555 -73.889 139.645 -72.882 ;
      RECT 139.555 -73.365 139.695 -73.195 ;
      RECT 139.555 -72.468 139.645 -71.461 ;
      RECT 139.555 -72.155 139.695 -71.985 ;
      RECT 139.555 -70.659 139.645 -69.652 ;
      RECT 139.555 -70.135 139.695 -69.965 ;
      RECT 139.555 -69.238 139.645 -68.231 ;
      RECT 139.555 -68.925 139.695 -68.755 ;
      RECT 139.555 -67.429 139.645 -66.422 ;
      RECT 139.555 -66.905 139.695 -66.735 ;
      RECT 139.555 -66.008 139.645 -65.001 ;
      RECT 139.555 -65.695 139.695 -65.525 ;
      RECT 139.555 -64.199 139.645 -63.192 ;
      RECT 139.555 -63.675 139.695 -63.505 ;
      RECT 139.555 -62.778 139.645 -61.771 ;
      RECT 139.555 -62.465 139.695 -62.295 ;
      RECT 139.555 -60.969 139.645 -59.962 ;
      RECT 139.555 -60.445 139.695 -60.275 ;
      RECT 139.555 -59.548 139.645 -58.541 ;
      RECT 139.555 -59.235 139.695 -59.065 ;
      RECT 139.555 -57.739 139.645 -56.732 ;
      RECT 139.555 -57.215 139.695 -57.045 ;
      RECT 139.555 -56.318 139.645 -55.311 ;
      RECT 139.555 -56.005 139.695 -55.835 ;
      RECT 139.555 -54.509 139.645 -53.502 ;
      RECT 139.555 -53.985 139.695 -53.815 ;
      RECT 139.555 -53.088 139.645 -52.081 ;
      RECT 139.555 -52.775 139.695 -52.605 ;
      RECT 139.555 -51.279 139.645 -50.272 ;
      RECT 139.555 -50.755 139.695 -50.585 ;
      RECT 139.555 -49.858 139.645 -48.851 ;
      RECT 139.555 -49.545 139.695 -49.375 ;
      RECT 139.555 -48.049 139.645 -47.042 ;
      RECT 139.555 -47.525 139.695 -47.355 ;
      RECT 139.555 -46.628 139.645 -45.621 ;
      RECT 139.555 -46.315 139.695 -46.145 ;
      RECT 139.555 -44.819 139.645 -43.812 ;
      RECT 139.555 -44.295 139.695 -44.125 ;
      RECT 139.555 -43.398 139.645 -42.391 ;
      RECT 139.555 -43.085 139.695 -42.915 ;
      RECT 139.555 -41.589 139.645 -40.582 ;
      RECT 139.555 -41.065 139.695 -40.895 ;
      RECT 139.555 -40.168 139.645 -39.161 ;
      RECT 139.555 -39.855 139.695 -39.685 ;
      RECT 139.555 -38.359 139.645 -37.352 ;
      RECT 139.555 -37.835 139.695 -37.665 ;
      RECT 139.555 -36.938 139.645 -35.931 ;
      RECT 139.555 -36.625 139.695 -36.455 ;
      RECT 139.555 -35.129 139.645 -34.122 ;
      RECT 139.555 -34.605 139.695 -34.435 ;
      RECT 139.555 -33.708 139.645 -32.701 ;
      RECT 139.555 -33.395 139.695 -33.225 ;
      RECT 139.555 -31.899 139.645 -30.892 ;
      RECT 139.555 -31.375 139.695 -31.205 ;
      RECT 139.555 -30.478 139.645 -29.471 ;
      RECT 139.555 -30.165 139.695 -29.995 ;
      RECT 139.555 -28.669 139.645 -27.662 ;
      RECT 139.555 -28.145 139.695 -27.975 ;
      RECT 139.555 -27.248 139.645 -26.241 ;
      RECT 139.555 -26.935 139.695 -26.765 ;
      RECT 139.555 -25.439 139.645 -24.432 ;
      RECT 139.555 -24.915 139.695 -24.745 ;
      RECT 139.555 -24.018 139.645 -23.011 ;
      RECT 139.555 -23.705 139.695 -23.535 ;
      RECT 139.555 -22.209 139.645 -21.202 ;
      RECT 139.555 -21.685 139.695 -21.515 ;
      RECT 139.555 -20.788 139.645 -19.781 ;
      RECT 139.555 -20.475 139.695 -20.305 ;
      RECT 139.555 -18.979 139.645 -17.972 ;
      RECT 139.555 -18.455 139.695 -18.285 ;
      RECT 139.555 -17.558 139.645 -16.551 ;
      RECT 139.555 -17.245 139.695 -17.075 ;
      RECT 139.555 -15.749 139.645 -14.742 ;
      RECT 139.555 -15.225 139.695 -15.055 ;
      RECT 139.555 -14.328 139.645 -13.321 ;
      RECT 139.555 -14.015 139.695 -13.845 ;
      RECT 139.555 -12.519 139.645 -11.512 ;
      RECT 139.555 -11.995 139.695 -11.825 ;
      RECT 139.555 -11.098 139.645 -10.091 ;
      RECT 139.555 -10.785 139.695 -10.615 ;
      RECT 139.555 -9.289 139.645 -8.282 ;
      RECT 139.555 -8.765 139.695 -8.595 ;
      RECT 139.555 -7.868 139.645 -6.861 ;
      RECT 139.555 -7.555 139.695 -7.385 ;
      RECT 139.555 -6.059 139.645 -5.052 ;
      RECT 139.555 -5.535 139.695 -5.365 ;
      RECT 139.555 -4.638 139.645 -3.631 ;
      RECT 139.555 -4.325 139.695 -4.155 ;
      RECT 139.555 -2.829 139.645 -1.822 ;
      RECT 139.555 -2.305 139.695 -2.135 ;
      RECT 139.555 -1.408 139.645 -0.401 ;
      RECT 139.555 -1.095 139.695 -0.925 ;
      RECT 139.555 0.401 139.645 1.408 ;
      RECT 139.555 0.925 139.695 1.095 ;
      RECT 135.385 -108.935 139.165 -108.815 ;
      RECT 136.705 -109.475 136.805 -108.815 ;
      RECT 136.145 -109.475 136.245 -108.815 ;
      RECT 135.585 -109.475 135.685 -108.815 ;
      RECT 138.755 -101.538 138.845 -100.53 ;
      RECT 138.705 -100.935 138.845 -100.765 ;
      RECT 138.755 -99.73 138.845 -98.722 ;
      RECT 138.705 -99.495 138.845 -99.325 ;
      RECT 138.755 -98.308 138.845 -97.3 ;
      RECT 138.705 -97.705 138.845 -97.535 ;
      RECT 138.755 -96.5 138.845 -95.492 ;
      RECT 138.705 -96.265 138.845 -96.095 ;
      RECT 138.755 -95.078 138.845 -94.07 ;
      RECT 138.705 -94.475 138.845 -94.305 ;
      RECT 138.755 -93.27 138.845 -92.262 ;
      RECT 138.705 -93.035 138.845 -92.865 ;
      RECT 138.755 -91.848 138.845 -90.84 ;
      RECT 138.705 -91.245 138.845 -91.075 ;
      RECT 138.755 -90.04 138.845 -89.032 ;
      RECT 138.705 -89.805 138.845 -89.635 ;
      RECT 138.755 -88.618 138.845 -87.61 ;
      RECT 138.705 -88.015 138.845 -87.845 ;
      RECT 138.755 -86.81 138.845 -85.802 ;
      RECT 138.705 -86.575 138.845 -86.405 ;
      RECT 138.755 -85.388 138.845 -84.38 ;
      RECT 138.705 -84.785 138.845 -84.615 ;
      RECT 138.755 -83.58 138.845 -82.572 ;
      RECT 138.705 -83.345 138.845 -83.175 ;
      RECT 138.755 -82.158 138.845 -81.15 ;
      RECT 138.705 -81.555 138.845 -81.385 ;
      RECT 138.755 -80.35 138.845 -79.342 ;
      RECT 138.705 -80.115 138.845 -79.945 ;
      RECT 138.755 -78.928 138.845 -77.92 ;
      RECT 138.705 -78.325 138.845 -78.155 ;
      RECT 138.755 -77.12 138.845 -76.112 ;
      RECT 138.705 -76.885 138.845 -76.715 ;
      RECT 138.755 -75.698 138.845 -74.69 ;
      RECT 138.705 -75.095 138.845 -74.925 ;
      RECT 138.755 -73.89 138.845 -72.882 ;
      RECT 138.705 -73.655 138.845 -73.485 ;
      RECT 138.755 -72.468 138.845 -71.46 ;
      RECT 138.705 -71.865 138.845 -71.695 ;
      RECT 138.755 -70.66 138.845 -69.652 ;
      RECT 138.705 -70.425 138.845 -70.255 ;
      RECT 138.755 -69.238 138.845 -68.23 ;
      RECT 138.705 -68.635 138.845 -68.465 ;
      RECT 138.755 -67.43 138.845 -66.422 ;
      RECT 138.705 -67.195 138.845 -67.025 ;
      RECT 138.755 -66.008 138.845 -65 ;
      RECT 138.705 -65.405 138.845 -65.235 ;
      RECT 138.755 -64.2 138.845 -63.192 ;
      RECT 138.705 -63.965 138.845 -63.795 ;
      RECT 138.755 -62.778 138.845 -61.77 ;
      RECT 138.705 -62.175 138.845 -62.005 ;
      RECT 138.755 -60.97 138.845 -59.962 ;
      RECT 138.705 -60.735 138.845 -60.565 ;
      RECT 138.755 -59.548 138.845 -58.54 ;
      RECT 138.705 -58.945 138.845 -58.775 ;
      RECT 138.755 -57.74 138.845 -56.732 ;
      RECT 138.705 -57.505 138.845 -57.335 ;
      RECT 138.755 -56.318 138.845 -55.31 ;
      RECT 138.705 -55.715 138.845 -55.545 ;
      RECT 138.755 -54.51 138.845 -53.502 ;
      RECT 138.705 -54.275 138.845 -54.105 ;
      RECT 138.755 -53.088 138.845 -52.08 ;
      RECT 138.705 -52.485 138.845 -52.315 ;
      RECT 138.755 -51.28 138.845 -50.272 ;
      RECT 138.705 -51.045 138.845 -50.875 ;
      RECT 138.755 -49.858 138.845 -48.85 ;
      RECT 138.705 -49.255 138.845 -49.085 ;
      RECT 138.755 -48.05 138.845 -47.042 ;
      RECT 138.705 -47.815 138.845 -47.645 ;
      RECT 138.755 -46.628 138.845 -45.62 ;
      RECT 138.705 -46.025 138.845 -45.855 ;
      RECT 138.755 -44.82 138.845 -43.812 ;
      RECT 138.705 -44.585 138.845 -44.415 ;
      RECT 138.755 -43.398 138.845 -42.39 ;
      RECT 138.705 -42.795 138.845 -42.625 ;
      RECT 138.755 -41.59 138.845 -40.582 ;
      RECT 138.705 -41.355 138.845 -41.185 ;
      RECT 138.755 -40.168 138.845 -39.16 ;
      RECT 138.705 -39.565 138.845 -39.395 ;
      RECT 138.755 -38.36 138.845 -37.352 ;
      RECT 138.705 -38.125 138.845 -37.955 ;
      RECT 138.755 -36.938 138.845 -35.93 ;
      RECT 138.705 -36.335 138.845 -36.165 ;
      RECT 138.755 -35.13 138.845 -34.122 ;
      RECT 138.705 -34.895 138.845 -34.725 ;
      RECT 138.755 -33.708 138.845 -32.7 ;
      RECT 138.705 -33.105 138.845 -32.935 ;
      RECT 138.755 -31.9 138.845 -30.892 ;
      RECT 138.705 -31.665 138.845 -31.495 ;
      RECT 138.755 -30.478 138.845 -29.47 ;
      RECT 138.705 -29.875 138.845 -29.705 ;
      RECT 138.755 -28.67 138.845 -27.662 ;
      RECT 138.705 -28.435 138.845 -28.265 ;
      RECT 138.755 -27.248 138.845 -26.24 ;
      RECT 138.705 -26.645 138.845 -26.475 ;
      RECT 138.755 -25.44 138.845 -24.432 ;
      RECT 138.705 -25.205 138.845 -25.035 ;
      RECT 138.755 -24.018 138.845 -23.01 ;
      RECT 138.705 -23.415 138.845 -23.245 ;
      RECT 138.755 -22.21 138.845 -21.202 ;
      RECT 138.705 -21.975 138.845 -21.805 ;
      RECT 138.755 -20.788 138.845 -19.78 ;
      RECT 138.705 -20.185 138.845 -20.015 ;
      RECT 138.755 -18.98 138.845 -17.972 ;
      RECT 138.705 -18.745 138.845 -18.575 ;
      RECT 138.755 -17.558 138.845 -16.55 ;
      RECT 138.705 -16.955 138.845 -16.785 ;
      RECT 138.755 -15.75 138.845 -14.742 ;
      RECT 138.705 -15.515 138.845 -15.345 ;
      RECT 138.755 -14.328 138.845 -13.32 ;
      RECT 138.705 -13.725 138.845 -13.555 ;
      RECT 138.755 -12.52 138.845 -11.512 ;
      RECT 138.705 -12.285 138.845 -12.115 ;
      RECT 138.755 -11.098 138.845 -10.09 ;
      RECT 138.705 -10.495 138.845 -10.325 ;
      RECT 138.755 -9.29 138.845 -8.282 ;
      RECT 138.705 -9.055 138.845 -8.885 ;
      RECT 138.755 -7.868 138.845 -6.86 ;
      RECT 138.705 -7.265 138.845 -7.095 ;
      RECT 138.755 -6.06 138.845 -5.052 ;
      RECT 138.705 -5.825 138.845 -5.655 ;
      RECT 138.755 -4.638 138.845 -3.63 ;
      RECT 138.705 -4.035 138.845 -3.865 ;
      RECT 138.755 -2.83 138.845 -1.822 ;
      RECT 138.705 -2.595 138.845 -2.425 ;
      RECT 138.755 -1.408 138.845 -0.4 ;
      RECT 138.705 -0.805 138.845 -0.635 ;
      RECT 138.755 0.4 138.845 1.408 ;
      RECT 138.705 0.635 138.845 0.805 ;
      RECT 137.325 -111.685 138.805 -111.585 ;
      RECT 137.325 -112.195 137.425 -111.585 ;
      RECT 137.545 -109.15 138.805 -109.05 ;
      RECT 138.705 -109.475 138.805 -109.05 ;
      RECT 138.145 -109.475 138.245 -109.05 ;
      RECT 137.585 -109.475 137.685 -109.05 ;
      RECT 138.355 -101.538 138.445 -100.531 ;
      RECT 138.355 -101.225 138.495 -101.055 ;
      RECT 138.355 -99.729 138.445 -98.722 ;
      RECT 138.355 -99.205 138.495 -99.035 ;
      RECT 138.355 -98.308 138.445 -97.301 ;
      RECT 138.355 -97.995 138.495 -97.825 ;
      RECT 138.355 -96.499 138.445 -95.492 ;
      RECT 138.355 -95.975 138.495 -95.805 ;
      RECT 138.355 -95.078 138.445 -94.071 ;
      RECT 138.355 -94.765 138.495 -94.595 ;
      RECT 138.355 -93.269 138.445 -92.262 ;
      RECT 138.355 -92.745 138.495 -92.575 ;
      RECT 138.355 -91.848 138.445 -90.841 ;
      RECT 138.355 -91.535 138.495 -91.365 ;
      RECT 138.355 -90.039 138.445 -89.032 ;
      RECT 138.355 -89.515 138.495 -89.345 ;
      RECT 138.355 -88.618 138.445 -87.611 ;
      RECT 138.355 -88.305 138.495 -88.135 ;
      RECT 138.355 -86.809 138.445 -85.802 ;
      RECT 138.355 -86.285 138.495 -86.115 ;
      RECT 138.355 -85.388 138.445 -84.381 ;
      RECT 138.355 -85.075 138.495 -84.905 ;
      RECT 138.355 -83.579 138.445 -82.572 ;
      RECT 138.355 -83.055 138.495 -82.885 ;
      RECT 138.355 -82.158 138.445 -81.151 ;
      RECT 138.355 -81.845 138.495 -81.675 ;
      RECT 138.355 -80.349 138.445 -79.342 ;
      RECT 138.355 -79.825 138.495 -79.655 ;
      RECT 138.355 -78.928 138.445 -77.921 ;
      RECT 138.355 -78.615 138.495 -78.445 ;
      RECT 138.355 -77.119 138.445 -76.112 ;
      RECT 138.355 -76.595 138.495 -76.425 ;
      RECT 138.355 -75.698 138.445 -74.691 ;
      RECT 138.355 -75.385 138.495 -75.215 ;
      RECT 138.355 -73.889 138.445 -72.882 ;
      RECT 138.355 -73.365 138.495 -73.195 ;
      RECT 138.355 -72.468 138.445 -71.461 ;
      RECT 138.355 -72.155 138.495 -71.985 ;
      RECT 138.355 -70.659 138.445 -69.652 ;
      RECT 138.355 -70.135 138.495 -69.965 ;
      RECT 138.355 -69.238 138.445 -68.231 ;
      RECT 138.355 -68.925 138.495 -68.755 ;
      RECT 138.355 -67.429 138.445 -66.422 ;
      RECT 138.355 -66.905 138.495 -66.735 ;
      RECT 138.355 -66.008 138.445 -65.001 ;
      RECT 138.355 -65.695 138.495 -65.525 ;
      RECT 138.355 -64.199 138.445 -63.192 ;
      RECT 138.355 -63.675 138.495 -63.505 ;
      RECT 138.355 -62.778 138.445 -61.771 ;
      RECT 138.355 -62.465 138.495 -62.295 ;
      RECT 138.355 -60.969 138.445 -59.962 ;
      RECT 138.355 -60.445 138.495 -60.275 ;
      RECT 138.355 -59.548 138.445 -58.541 ;
      RECT 138.355 -59.235 138.495 -59.065 ;
      RECT 138.355 -57.739 138.445 -56.732 ;
      RECT 138.355 -57.215 138.495 -57.045 ;
      RECT 138.355 -56.318 138.445 -55.311 ;
      RECT 138.355 -56.005 138.495 -55.835 ;
      RECT 138.355 -54.509 138.445 -53.502 ;
      RECT 138.355 -53.985 138.495 -53.815 ;
      RECT 138.355 -53.088 138.445 -52.081 ;
      RECT 138.355 -52.775 138.495 -52.605 ;
      RECT 138.355 -51.279 138.445 -50.272 ;
      RECT 138.355 -50.755 138.495 -50.585 ;
      RECT 138.355 -49.858 138.445 -48.851 ;
      RECT 138.355 -49.545 138.495 -49.375 ;
      RECT 138.355 -48.049 138.445 -47.042 ;
      RECT 138.355 -47.525 138.495 -47.355 ;
      RECT 138.355 -46.628 138.445 -45.621 ;
      RECT 138.355 -46.315 138.495 -46.145 ;
      RECT 138.355 -44.819 138.445 -43.812 ;
      RECT 138.355 -44.295 138.495 -44.125 ;
      RECT 138.355 -43.398 138.445 -42.391 ;
      RECT 138.355 -43.085 138.495 -42.915 ;
      RECT 138.355 -41.589 138.445 -40.582 ;
      RECT 138.355 -41.065 138.495 -40.895 ;
      RECT 138.355 -40.168 138.445 -39.161 ;
      RECT 138.355 -39.855 138.495 -39.685 ;
      RECT 138.355 -38.359 138.445 -37.352 ;
      RECT 138.355 -37.835 138.495 -37.665 ;
      RECT 138.355 -36.938 138.445 -35.931 ;
      RECT 138.355 -36.625 138.495 -36.455 ;
      RECT 138.355 -35.129 138.445 -34.122 ;
      RECT 138.355 -34.605 138.495 -34.435 ;
      RECT 138.355 -33.708 138.445 -32.701 ;
      RECT 138.355 -33.395 138.495 -33.225 ;
      RECT 138.355 -31.899 138.445 -30.892 ;
      RECT 138.355 -31.375 138.495 -31.205 ;
      RECT 138.355 -30.478 138.445 -29.471 ;
      RECT 138.355 -30.165 138.495 -29.995 ;
      RECT 138.355 -28.669 138.445 -27.662 ;
      RECT 138.355 -28.145 138.495 -27.975 ;
      RECT 138.355 -27.248 138.445 -26.241 ;
      RECT 138.355 -26.935 138.495 -26.765 ;
      RECT 138.355 -25.439 138.445 -24.432 ;
      RECT 138.355 -24.915 138.495 -24.745 ;
      RECT 138.355 -24.018 138.445 -23.011 ;
      RECT 138.355 -23.705 138.495 -23.535 ;
      RECT 138.355 -22.209 138.445 -21.202 ;
      RECT 138.355 -21.685 138.495 -21.515 ;
      RECT 138.355 -20.788 138.445 -19.781 ;
      RECT 138.355 -20.475 138.495 -20.305 ;
      RECT 138.355 -18.979 138.445 -17.972 ;
      RECT 138.355 -18.455 138.495 -18.285 ;
      RECT 138.355 -17.558 138.445 -16.551 ;
      RECT 138.355 -17.245 138.495 -17.075 ;
      RECT 138.355 -15.749 138.445 -14.742 ;
      RECT 138.355 -15.225 138.495 -15.055 ;
      RECT 138.355 -14.328 138.445 -13.321 ;
      RECT 138.355 -14.015 138.495 -13.845 ;
      RECT 138.355 -12.519 138.445 -11.512 ;
      RECT 138.355 -11.995 138.495 -11.825 ;
      RECT 138.355 -11.098 138.445 -10.091 ;
      RECT 138.355 -10.785 138.495 -10.615 ;
      RECT 138.355 -9.289 138.445 -8.282 ;
      RECT 138.355 -8.765 138.495 -8.595 ;
      RECT 138.355 -7.868 138.445 -6.861 ;
      RECT 138.355 -7.555 138.495 -7.385 ;
      RECT 138.355 -6.059 138.445 -5.052 ;
      RECT 138.355 -5.535 138.495 -5.365 ;
      RECT 138.355 -4.638 138.445 -3.631 ;
      RECT 138.355 -4.325 138.495 -4.155 ;
      RECT 138.355 -2.829 138.445 -1.822 ;
      RECT 138.355 -2.305 138.495 -2.135 ;
      RECT 138.355 -1.408 138.445 -0.401 ;
      RECT 138.355 -1.095 138.495 -0.925 ;
      RECT 138.355 0.401 138.445 1.408 ;
      RECT 138.355 0.925 138.495 1.095 ;
      RECT 137.685 -111.495 137.855 -111.385 ;
      RECT 134.535 -111.495 137.855 -111.395 ;
      RECT 137.555 -101.538 137.645 -100.53 ;
      RECT 137.505 -100.935 137.645 -100.765 ;
      RECT 137.555 -99.73 137.645 -98.722 ;
      RECT 137.505 -99.495 137.645 -99.325 ;
      RECT 137.555 -98.308 137.645 -97.3 ;
      RECT 137.505 -97.705 137.645 -97.535 ;
      RECT 137.555 -96.5 137.645 -95.492 ;
      RECT 137.505 -96.265 137.645 -96.095 ;
      RECT 137.555 -95.078 137.645 -94.07 ;
      RECT 137.505 -94.475 137.645 -94.305 ;
      RECT 137.555 -93.27 137.645 -92.262 ;
      RECT 137.505 -93.035 137.645 -92.865 ;
      RECT 137.555 -91.848 137.645 -90.84 ;
      RECT 137.505 -91.245 137.645 -91.075 ;
      RECT 137.555 -90.04 137.645 -89.032 ;
      RECT 137.505 -89.805 137.645 -89.635 ;
      RECT 137.555 -88.618 137.645 -87.61 ;
      RECT 137.505 -88.015 137.645 -87.845 ;
      RECT 137.555 -86.81 137.645 -85.802 ;
      RECT 137.505 -86.575 137.645 -86.405 ;
      RECT 137.555 -85.388 137.645 -84.38 ;
      RECT 137.505 -84.785 137.645 -84.615 ;
      RECT 137.555 -83.58 137.645 -82.572 ;
      RECT 137.505 -83.345 137.645 -83.175 ;
      RECT 137.555 -82.158 137.645 -81.15 ;
      RECT 137.505 -81.555 137.645 -81.385 ;
      RECT 137.555 -80.35 137.645 -79.342 ;
      RECT 137.505 -80.115 137.645 -79.945 ;
      RECT 137.555 -78.928 137.645 -77.92 ;
      RECT 137.505 -78.325 137.645 -78.155 ;
      RECT 137.555 -77.12 137.645 -76.112 ;
      RECT 137.505 -76.885 137.645 -76.715 ;
      RECT 137.555 -75.698 137.645 -74.69 ;
      RECT 137.505 -75.095 137.645 -74.925 ;
      RECT 137.555 -73.89 137.645 -72.882 ;
      RECT 137.505 -73.655 137.645 -73.485 ;
      RECT 137.555 -72.468 137.645 -71.46 ;
      RECT 137.505 -71.865 137.645 -71.695 ;
      RECT 137.555 -70.66 137.645 -69.652 ;
      RECT 137.505 -70.425 137.645 -70.255 ;
      RECT 137.555 -69.238 137.645 -68.23 ;
      RECT 137.505 -68.635 137.645 -68.465 ;
      RECT 137.555 -67.43 137.645 -66.422 ;
      RECT 137.505 -67.195 137.645 -67.025 ;
      RECT 137.555 -66.008 137.645 -65 ;
      RECT 137.505 -65.405 137.645 -65.235 ;
      RECT 137.555 -64.2 137.645 -63.192 ;
      RECT 137.505 -63.965 137.645 -63.795 ;
      RECT 137.555 -62.778 137.645 -61.77 ;
      RECT 137.505 -62.175 137.645 -62.005 ;
      RECT 137.555 -60.97 137.645 -59.962 ;
      RECT 137.505 -60.735 137.645 -60.565 ;
      RECT 137.555 -59.548 137.645 -58.54 ;
      RECT 137.505 -58.945 137.645 -58.775 ;
      RECT 137.555 -57.74 137.645 -56.732 ;
      RECT 137.505 -57.505 137.645 -57.335 ;
      RECT 137.555 -56.318 137.645 -55.31 ;
      RECT 137.505 -55.715 137.645 -55.545 ;
      RECT 137.555 -54.51 137.645 -53.502 ;
      RECT 137.505 -54.275 137.645 -54.105 ;
      RECT 137.555 -53.088 137.645 -52.08 ;
      RECT 137.505 -52.485 137.645 -52.315 ;
      RECT 137.555 -51.28 137.645 -50.272 ;
      RECT 137.505 -51.045 137.645 -50.875 ;
      RECT 137.555 -49.858 137.645 -48.85 ;
      RECT 137.505 -49.255 137.645 -49.085 ;
      RECT 137.555 -48.05 137.645 -47.042 ;
      RECT 137.505 -47.815 137.645 -47.645 ;
      RECT 137.555 -46.628 137.645 -45.62 ;
      RECT 137.505 -46.025 137.645 -45.855 ;
      RECT 137.555 -44.82 137.645 -43.812 ;
      RECT 137.505 -44.585 137.645 -44.415 ;
      RECT 137.555 -43.398 137.645 -42.39 ;
      RECT 137.505 -42.795 137.645 -42.625 ;
      RECT 137.555 -41.59 137.645 -40.582 ;
      RECT 137.505 -41.355 137.645 -41.185 ;
      RECT 137.555 -40.168 137.645 -39.16 ;
      RECT 137.505 -39.565 137.645 -39.395 ;
      RECT 137.555 -38.36 137.645 -37.352 ;
      RECT 137.505 -38.125 137.645 -37.955 ;
      RECT 137.555 -36.938 137.645 -35.93 ;
      RECT 137.505 -36.335 137.645 -36.165 ;
      RECT 137.555 -35.13 137.645 -34.122 ;
      RECT 137.505 -34.895 137.645 -34.725 ;
      RECT 137.555 -33.708 137.645 -32.7 ;
      RECT 137.505 -33.105 137.645 -32.935 ;
      RECT 137.555 -31.9 137.645 -30.892 ;
      RECT 137.505 -31.665 137.645 -31.495 ;
      RECT 137.555 -30.478 137.645 -29.47 ;
      RECT 137.505 -29.875 137.645 -29.705 ;
      RECT 137.555 -28.67 137.645 -27.662 ;
      RECT 137.505 -28.435 137.645 -28.265 ;
      RECT 137.555 -27.248 137.645 -26.24 ;
      RECT 137.505 -26.645 137.645 -26.475 ;
      RECT 137.555 -25.44 137.645 -24.432 ;
      RECT 137.505 -25.205 137.645 -25.035 ;
      RECT 137.555 -24.018 137.645 -23.01 ;
      RECT 137.505 -23.415 137.645 -23.245 ;
      RECT 137.555 -22.21 137.645 -21.202 ;
      RECT 137.505 -21.975 137.645 -21.805 ;
      RECT 137.555 -20.788 137.645 -19.78 ;
      RECT 137.505 -20.185 137.645 -20.015 ;
      RECT 137.555 -18.98 137.645 -17.972 ;
      RECT 137.505 -18.745 137.645 -18.575 ;
      RECT 137.555 -17.558 137.645 -16.55 ;
      RECT 137.505 -16.955 137.645 -16.785 ;
      RECT 137.555 -15.75 137.645 -14.742 ;
      RECT 137.505 -15.515 137.645 -15.345 ;
      RECT 137.555 -14.328 137.645 -13.32 ;
      RECT 137.505 -13.725 137.645 -13.555 ;
      RECT 137.555 -12.52 137.645 -11.512 ;
      RECT 137.505 -12.285 137.645 -12.115 ;
      RECT 137.555 -11.098 137.645 -10.09 ;
      RECT 137.505 -10.495 137.645 -10.325 ;
      RECT 137.555 -9.29 137.645 -8.282 ;
      RECT 137.505 -9.055 137.645 -8.885 ;
      RECT 137.555 -7.868 137.645 -6.86 ;
      RECT 137.505 -7.265 137.645 -7.095 ;
      RECT 137.555 -6.06 137.645 -5.052 ;
      RECT 137.505 -5.825 137.645 -5.655 ;
      RECT 137.555 -4.638 137.645 -3.63 ;
      RECT 137.505 -4.035 137.645 -3.865 ;
      RECT 137.555 -2.83 137.645 -1.822 ;
      RECT 137.505 -2.595 137.645 -2.425 ;
      RECT 137.555 -1.408 137.645 -0.4 ;
      RECT 137.505 -0.805 137.645 -0.635 ;
      RECT 137.555 0.4 137.645 1.408 ;
      RECT 137.505 0.635 137.645 0.805 ;
      RECT 137.155 -101.538 137.245 -100.531 ;
      RECT 137.155 -101.225 137.295 -101.055 ;
      RECT 137.155 -99.729 137.245 -98.722 ;
      RECT 137.155 -99.205 137.295 -99.035 ;
      RECT 137.155 -98.308 137.245 -97.301 ;
      RECT 137.155 -97.995 137.295 -97.825 ;
      RECT 137.155 -96.499 137.245 -95.492 ;
      RECT 137.155 -95.975 137.295 -95.805 ;
      RECT 137.155 -95.078 137.245 -94.071 ;
      RECT 137.155 -94.765 137.295 -94.595 ;
      RECT 137.155 -93.269 137.245 -92.262 ;
      RECT 137.155 -92.745 137.295 -92.575 ;
      RECT 137.155 -91.848 137.245 -90.841 ;
      RECT 137.155 -91.535 137.295 -91.365 ;
      RECT 137.155 -90.039 137.245 -89.032 ;
      RECT 137.155 -89.515 137.295 -89.345 ;
      RECT 137.155 -88.618 137.245 -87.611 ;
      RECT 137.155 -88.305 137.295 -88.135 ;
      RECT 137.155 -86.809 137.245 -85.802 ;
      RECT 137.155 -86.285 137.295 -86.115 ;
      RECT 137.155 -85.388 137.245 -84.381 ;
      RECT 137.155 -85.075 137.295 -84.905 ;
      RECT 137.155 -83.579 137.245 -82.572 ;
      RECT 137.155 -83.055 137.295 -82.885 ;
      RECT 137.155 -82.158 137.245 -81.151 ;
      RECT 137.155 -81.845 137.295 -81.675 ;
      RECT 137.155 -80.349 137.245 -79.342 ;
      RECT 137.155 -79.825 137.295 -79.655 ;
      RECT 137.155 -78.928 137.245 -77.921 ;
      RECT 137.155 -78.615 137.295 -78.445 ;
      RECT 137.155 -77.119 137.245 -76.112 ;
      RECT 137.155 -76.595 137.295 -76.425 ;
      RECT 137.155 -75.698 137.245 -74.691 ;
      RECT 137.155 -75.385 137.295 -75.215 ;
      RECT 137.155 -73.889 137.245 -72.882 ;
      RECT 137.155 -73.365 137.295 -73.195 ;
      RECT 137.155 -72.468 137.245 -71.461 ;
      RECT 137.155 -72.155 137.295 -71.985 ;
      RECT 137.155 -70.659 137.245 -69.652 ;
      RECT 137.155 -70.135 137.295 -69.965 ;
      RECT 137.155 -69.238 137.245 -68.231 ;
      RECT 137.155 -68.925 137.295 -68.755 ;
      RECT 137.155 -67.429 137.245 -66.422 ;
      RECT 137.155 -66.905 137.295 -66.735 ;
      RECT 137.155 -66.008 137.245 -65.001 ;
      RECT 137.155 -65.695 137.295 -65.525 ;
      RECT 137.155 -64.199 137.245 -63.192 ;
      RECT 137.155 -63.675 137.295 -63.505 ;
      RECT 137.155 -62.778 137.245 -61.771 ;
      RECT 137.155 -62.465 137.295 -62.295 ;
      RECT 137.155 -60.969 137.245 -59.962 ;
      RECT 137.155 -60.445 137.295 -60.275 ;
      RECT 137.155 -59.548 137.245 -58.541 ;
      RECT 137.155 -59.235 137.295 -59.065 ;
      RECT 137.155 -57.739 137.245 -56.732 ;
      RECT 137.155 -57.215 137.295 -57.045 ;
      RECT 137.155 -56.318 137.245 -55.311 ;
      RECT 137.155 -56.005 137.295 -55.835 ;
      RECT 137.155 -54.509 137.245 -53.502 ;
      RECT 137.155 -53.985 137.295 -53.815 ;
      RECT 137.155 -53.088 137.245 -52.081 ;
      RECT 137.155 -52.775 137.295 -52.605 ;
      RECT 137.155 -51.279 137.245 -50.272 ;
      RECT 137.155 -50.755 137.295 -50.585 ;
      RECT 137.155 -49.858 137.245 -48.851 ;
      RECT 137.155 -49.545 137.295 -49.375 ;
      RECT 137.155 -48.049 137.245 -47.042 ;
      RECT 137.155 -47.525 137.295 -47.355 ;
      RECT 137.155 -46.628 137.245 -45.621 ;
      RECT 137.155 -46.315 137.295 -46.145 ;
      RECT 137.155 -44.819 137.245 -43.812 ;
      RECT 137.155 -44.295 137.295 -44.125 ;
      RECT 137.155 -43.398 137.245 -42.391 ;
      RECT 137.155 -43.085 137.295 -42.915 ;
      RECT 137.155 -41.589 137.245 -40.582 ;
      RECT 137.155 -41.065 137.295 -40.895 ;
      RECT 137.155 -40.168 137.245 -39.161 ;
      RECT 137.155 -39.855 137.295 -39.685 ;
      RECT 137.155 -38.359 137.245 -37.352 ;
      RECT 137.155 -37.835 137.295 -37.665 ;
      RECT 137.155 -36.938 137.245 -35.931 ;
      RECT 137.155 -36.625 137.295 -36.455 ;
      RECT 137.155 -35.129 137.245 -34.122 ;
      RECT 137.155 -34.605 137.295 -34.435 ;
      RECT 137.155 -33.708 137.245 -32.701 ;
      RECT 137.155 -33.395 137.295 -33.225 ;
      RECT 137.155 -31.899 137.245 -30.892 ;
      RECT 137.155 -31.375 137.295 -31.205 ;
      RECT 137.155 -30.478 137.245 -29.471 ;
      RECT 137.155 -30.165 137.295 -29.995 ;
      RECT 137.155 -28.669 137.245 -27.662 ;
      RECT 137.155 -28.145 137.295 -27.975 ;
      RECT 137.155 -27.248 137.245 -26.241 ;
      RECT 137.155 -26.935 137.295 -26.765 ;
      RECT 137.155 -25.439 137.245 -24.432 ;
      RECT 137.155 -24.915 137.295 -24.745 ;
      RECT 137.155 -24.018 137.245 -23.011 ;
      RECT 137.155 -23.705 137.295 -23.535 ;
      RECT 137.155 -22.209 137.245 -21.202 ;
      RECT 137.155 -21.685 137.295 -21.515 ;
      RECT 137.155 -20.788 137.245 -19.781 ;
      RECT 137.155 -20.475 137.295 -20.305 ;
      RECT 137.155 -18.979 137.245 -17.972 ;
      RECT 137.155 -18.455 137.295 -18.285 ;
      RECT 137.155 -17.558 137.245 -16.551 ;
      RECT 137.155 -17.245 137.295 -17.075 ;
      RECT 137.155 -15.749 137.245 -14.742 ;
      RECT 137.155 -15.225 137.295 -15.055 ;
      RECT 137.155 -14.328 137.245 -13.321 ;
      RECT 137.155 -14.015 137.295 -13.845 ;
      RECT 137.155 -12.519 137.245 -11.512 ;
      RECT 137.155 -11.995 137.295 -11.825 ;
      RECT 137.155 -11.098 137.245 -10.091 ;
      RECT 137.155 -10.785 137.295 -10.615 ;
      RECT 137.155 -9.289 137.245 -8.282 ;
      RECT 137.155 -8.765 137.295 -8.595 ;
      RECT 137.155 -7.868 137.245 -6.861 ;
      RECT 137.155 -7.555 137.295 -7.385 ;
      RECT 137.155 -6.059 137.245 -5.052 ;
      RECT 137.155 -5.535 137.295 -5.365 ;
      RECT 137.155 -4.638 137.245 -3.631 ;
      RECT 137.155 -4.325 137.295 -4.155 ;
      RECT 137.155 -2.829 137.245 -1.822 ;
      RECT 137.155 -2.305 137.295 -2.135 ;
      RECT 137.155 -1.408 137.245 -0.401 ;
      RECT 137.155 -1.095 137.295 -0.925 ;
      RECT 137.155 0.401 137.245 1.408 ;
      RECT 137.155 0.925 137.295 1.095 ;
      RECT 135.305 -111.685 136.785 -111.585 ;
      RECT 135.305 -112.055 135.405 -111.585 ;
      RECT 135.11 -114.395 136.685 -114.275 ;
      RECT 136.585 -114.895 136.685 -114.275 ;
      RECT 135.99 -114.895 136.09 -114.275 ;
      RECT 135.11 -114.85 135.21 -114.275 ;
      RECT 136.355 -101.538 136.445 -100.53 ;
      RECT 136.305 -100.935 136.445 -100.765 ;
      RECT 136.355 -99.73 136.445 -98.722 ;
      RECT 136.305 -99.495 136.445 -99.325 ;
      RECT 136.355 -98.308 136.445 -97.3 ;
      RECT 136.305 -97.705 136.445 -97.535 ;
      RECT 136.355 -96.5 136.445 -95.492 ;
      RECT 136.305 -96.265 136.445 -96.095 ;
      RECT 136.355 -95.078 136.445 -94.07 ;
      RECT 136.305 -94.475 136.445 -94.305 ;
      RECT 136.355 -93.27 136.445 -92.262 ;
      RECT 136.305 -93.035 136.445 -92.865 ;
      RECT 136.355 -91.848 136.445 -90.84 ;
      RECT 136.305 -91.245 136.445 -91.075 ;
      RECT 136.355 -90.04 136.445 -89.032 ;
      RECT 136.305 -89.805 136.445 -89.635 ;
      RECT 136.355 -88.618 136.445 -87.61 ;
      RECT 136.305 -88.015 136.445 -87.845 ;
      RECT 136.355 -86.81 136.445 -85.802 ;
      RECT 136.305 -86.575 136.445 -86.405 ;
      RECT 136.355 -85.388 136.445 -84.38 ;
      RECT 136.305 -84.785 136.445 -84.615 ;
      RECT 136.355 -83.58 136.445 -82.572 ;
      RECT 136.305 -83.345 136.445 -83.175 ;
      RECT 136.355 -82.158 136.445 -81.15 ;
      RECT 136.305 -81.555 136.445 -81.385 ;
      RECT 136.355 -80.35 136.445 -79.342 ;
      RECT 136.305 -80.115 136.445 -79.945 ;
      RECT 136.355 -78.928 136.445 -77.92 ;
      RECT 136.305 -78.325 136.445 -78.155 ;
      RECT 136.355 -77.12 136.445 -76.112 ;
      RECT 136.305 -76.885 136.445 -76.715 ;
      RECT 136.355 -75.698 136.445 -74.69 ;
      RECT 136.305 -75.095 136.445 -74.925 ;
      RECT 136.355 -73.89 136.445 -72.882 ;
      RECT 136.305 -73.655 136.445 -73.485 ;
      RECT 136.355 -72.468 136.445 -71.46 ;
      RECT 136.305 -71.865 136.445 -71.695 ;
      RECT 136.355 -70.66 136.445 -69.652 ;
      RECT 136.305 -70.425 136.445 -70.255 ;
      RECT 136.355 -69.238 136.445 -68.23 ;
      RECT 136.305 -68.635 136.445 -68.465 ;
      RECT 136.355 -67.43 136.445 -66.422 ;
      RECT 136.305 -67.195 136.445 -67.025 ;
      RECT 136.355 -66.008 136.445 -65 ;
      RECT 136.305 -65.405 136.445 -65.235 ;
      RECT 136.355 -64.2 136.445 -63.192 ;
      RECT 136.305 -63.965 136.445 -63.795 ;
      RECT 136.355 -62.778 136.445 -61.77 ;
      RECT 136.305 -62.175 136.445 -62.005 ;
      RECT 136.355 -60.97 136.445 -59.962 ;
      RECT 136.305 -60.735 136.445 -60.565 ;
      RECT 136.355 -59.548 136.445 -58.54 ;
      RECT 136.305 -58.945 136.445 -58.775 ;
      RECT 136.355 -57.74 136.445 -56.732 ;
      RECT 136.305 -57.505 136.445 -57.335 ;
      RECT 136.355 -56.318 136.445 -55.31 ;
      RECT 136.305 -55.715 136.445 -55.545 ;
      RECT 136.355 -54.51 136.445 -53.502 ;
      RECT 136.305 -54.275 136.445 -54.105 ;
      RECT 136.355 -53.088 136.445 -52.08 ;
      RECT 136.305 -52.485 136.445 -52.315 ;
      RECT 136.355 -51.28 136.445 -50.272 ;
      RECT 136.305 -51.045 136.445 -50.875 ;
      RECT 136.355 -49.858 136.445 -48.85 ;
      RECT 136.305 -49.255 136.445 -49.085 ;
      RECT 136.355 -48.05 136.445 -47.042 ;
      RECT 136.305 -47.815 136.445 -47.645 ;
      RECT 136.355 -46.628 136.445 -45.62 ;
      RECT 136.305 -46.025 136.445 -45.855 ;
      RECT 136.355 -44.82 136.445 -43.812 ;
      RECT 136.305 -44.585 136.445 -44.415 ;
      RECT 136.355 -43.398 136.445 -42.39 ;
      RECT 136.305 -42.795 136.445 -42.625 ;
      RECT 136.355 -41.59 136.445 -40.582 ;
      RECT 136.305 -41.355 136.445 -41.185 ;
      RECT 136.355 -40.168 136.445 -39.16 ;
      RECT 136.305 -39.565 136.445 -39.395 ;
      RECT 136.355 -38.36 136.445 -37.352 ;
      RECT 136.305 -38.125 136.445 -37.955 ;
      RECT 136.355 -36.938 136.445 -35.93 ;
      RECT 136.305 -36.335 136.445 -36.165 ;
      RECT 136.355 -35.13 136.445 -34.122 ;
      RECT 136.305 -34.895 136.445 -34.725 ;
      RECT 136.355 -33.708 136.445 -32.7 ;
      RECT 136.305 -33.105 136.445 -32.935 ;
      RECT 136.355 -31.9 136.445 -30.892 ;
      RECT 136.305 -31.665 136.445 -31.495 ;
      RECT 136.355 -30.478 136.445 -29.47 ;
      RECT 136.305 -29.875 136.445 -29.705 ;
      RECT 136.355 -28.67 136.445 -27.662 ;
      RECT 136.305 -28.435 136.445 -28.265 ;
      RECT 136.355 -27.248 136.445 -26.24 ;
      RECT 136.305 -26.645 136.445 -26.475 ;
      RECT 136.355 -25.44 136.445 -24.432 ;
      RECT 136.305 -25.205 136.445 -25.035 ;
      RECT 136.355 -24.018 136.445 -23.01 ;
      RECT 136.305 -23.415 136.445 -23.245 ;
      RECT 136.355 -22.21 136.445 -21.202 ;
      RECT 136.305 -21.975 136.445 -21.805 ;
      RECT 136.355 -20.788 136.445 -19.78 ;
      RECT 136.305 -20.185 136.445 -20.015 ;
      RECT 136.355 -18.98 136.445 -17.972 ;
      RECT 136.305 -18.745 136.445 -18.575 ;
      RECT 136.355 -17.558 136.445 -16.55 ;
      RECT 136.305 -16.955 136.445 -16.785 ;
      RECT 136.355 -15.75 136.445 -14.742 ;
      RECT 136.305 -15.515 136.445 -15.345 ;
      RECT 136.355 -14.328 136.445 -13.32 ;
      RECT 136.305 -13.725 136.445 -13.555 ;
      RECT 136.355 -12.52 136.445 -11.512 ;
      RECT 136.305 -12.285 136.445 -12.115 ;
      RECT 136.355 -11.098 136.445 -10.09 ;
      RECT 136.305 -10.495 136.445 -10.325 ;
      RECT 136.355 -9.29 136.445 -8.282 ;
      RECT 136.305 -9.055 136.445 -8.885 ;
      RECT 136.355 -7.868 136.445 -6.86 ;
      RECT 136.305 -7.265 136.445 -7.095 ;
      RECT 136.355 -6.06 136.445 -5.052 ;
      RECT 136.305 -5.825 136.445 -5.655 ;
      RECT 136.355 -4.638 136.445 -3.63 ;
      RECT 136.305 -4.035 136.445 -3.865 ;
      RECT 136.355 -2.83 136.445 -1.822 ;
      RECT 136.305 -2.595 136.445 -2.425 ;
      RECT 136.355 -1.408 136.445 -0.4 ;
      RECT 136.305 -0.805 136.445 -0.635 ;
      RECT 136.355 0.4 136.445 1.408 ;
      RECT 136.305 0.635 136.445 0.805 ;
      RECT 136.23 -114.685 136.405 -114.515 ;
      RECT 136.305 -114.895 136.405 -114.515 ;
      RECT 135.345 -113.555 135.445 -113.09 ;
      RECT 135.71 -113.555 135.81 -113.1 ;
      RECT 135.345 -113.555 136.19 -113.385 ;
      RECT 135.955 -101.538 136.045 -100.531 ;
      RECT 135.955 -101.225 136.095 -101.055 ;
      RECT 135.955 -99.729 136.045 -98.722 ;
      RECT 135.955 -99.205 136.095 -99.035 ;
      RECT 135.955 -98.308 136.045 -97.301 ;
      RECT 135.955 -97.995 136.095 -97.825 ;
      RECT 135.955 -96.499 136.045 -95.492 ;
      RECT 135.955 -95.975 136.095 -95.805 ;
      RECT 135.955 -95.078 136.045 -94.071 ;
      RECT 135.955 -94.765 136.095 -94.595 ;
      RECT 135.955 -93.269 136.045 -92.262 ;
      RECT 135.955 -92.745 136.095 -92.575 ;
      RECT 135.955 -91.848 136.045 -90.841 ;
      RECT 135.955 -91.535 136.095 -91.365 ;
      RECT 135.955 -90.039 136.045 -89.032 ;
      RECT 135.955 -89.515 136.095 -89.345 ;
      RECT 135.955 -88.618 136.045 -87.611 ;
      RECT 135.955 -88.305 136.095 -88.135 ;
      RECT 135.955 -86.809 136.045 -85.802 ;
      RECT 135.955 -86.285 136.095 -86.115 ;
      RECT 135.955 -85.388 136.045 -84.381 ;
      RECT 135.955 -85.075 136.095 -84.905 ;
      RECT 135.955 -83.579 136.045 -82.572 ;
      RECT 135.955 -83.055 136.095 -82.885 ;
      RECT 135.955 -82.158 136.045 -81.151 ;
      RECT 135.955 -81.845 136.095 -81.675 ;
      RECT 135.955 -80.349 136.045 -79.342 ;
      RECT 135.955 -79.825 136.095 -79.655 ;
      RECT 135.955 -78.928 136.045 -77.921 ;
      RECT 135.955 -78.615 136.095 -78.445 ;
      RECT 135.955 -77.119 136.045 -76.112 ;
      RECT 135.955 -76.595 136.095 -76.425 ;
      RECT 135.955 -75.698 136.045 -74.691 ;
      RECT 135.955 -75.385 136.095 -75.215 ;
      RECT 135.955 -73.889 136.045 -72.882 ;
      RECT 135.955 -73.365 136.095 -73.195 ;
      RECT 135.955 -72.468 136.045 -71.461 ;
      RECT 135.955 -72.155 136.095 -71.985 ;
      RECT 135.955 -70.659 136.045 -69.652 ;
      RECT 135.955 -70.135 136.095 -69.965 ;
      RECT 135.955 -69.238 136.045 -68.231 ;
      RECT 135.955 -68.925 136.095 -68.755 ;
      RECT 135.955 -67.429 136.045 -66.422 ;
      RECT 135.955 -66.905 136.095 -66.735 ;
      RECT 135.955 -66.008 136.045 -65.001 ;
      RECT 135.955 -65.695 136.095 -65.525 ;
      RECT 135.955 -64.199 136.045 -63.192 ;
      RECT 135.955 -63.675 136.095 -63.505 ;
      RECT 135.955 -62.778 136.045 -61.771 ;
      RECT 135.955 -62.465 136.095 -62.295 ;
      RECT 135.955 -60.969 136.045 -59.962 ;
      RECT 135.955 -60.445 136.095 -60.275 ;
      RECT 135.955 -59.548 136.045 -58.541 ;
      RECT 135.955 -59.235 136.095 -59.065 ;
      RECT 135.955 -57.739 136.045 -56.732 ;
      RECT 135.955 -57.215 136.095 -57.045 ;
      RECT 135.955 -56.318 136.045 -55.311 ;
      RECT 135.955 -56.005 136.095 -55.835 ;
      RECT 135.955 -54.509 136.045 -53.502 ;
      RECT 135.955 -53.985 136.095 -53.815 ;
      RECT 135.955 -53.088 136.045 -52.081 ;
      RECT 135.955 -52.775 136.095 -52.605 ;
      RECT 135.955 -51.279 136.045 -50.272 ;
      RECT 135.955 -50.755 136.095 -50.585 ;
      RECT 135.955 -49.858 136.045 -48.851 ;
      RECT 135.955 -49.545 136.095 -49.375 ;
      RECT 135.955 -48.049 136.045 -47.042 ;
      RECT 135.955 -47.525 136.095 -47.355 ;
      RECT 135.955 -46.628 136.045 -45.621 ;
      RECT 135.955 -46.315 136.095 -46.145 ;
      RECT 135.955 -44.819 136.045 -43.812 ;
      RECT 135.955 -44.295 136.095 -44.125 ;
      RECT 135.955 -43.398 136.045 -42.391 ;
      RECT 135.955 -43.085 136.095 -42.915 ;
      RECT 135.955 -41.589 136.045 -40.582 ;
      RECT 135.955 -41.065 136.095 -40.895 ;
      RECT 135.955 -40.168 136.045 -39.161 ;
      RECT 135.955 -39.855 136.095 -39.685 ;
      RECT 135.955 -38.359 136.045 -37.352 ;
      RECT 135.955 -37.835 136.095 -37.665 ;
      RECT 135.955 -36.938 136.045 -35.931 ;
      RECT 135.955 -36.625 136.095 -36.455 ;
      RECT 135.955 -35.129 136.045 -34.122 ;
      RECT 135.955 -34.605 136.095 -34.435 ;
      RECT 135.955 -33.708 136.045 -32.701 ;
      RECT 135.955 -33.395 136.095 -33.225 ;
      RECT 135.955 -31.899 136.045 -30.892 ;
      RECT 135.955 -31.375 136.095 -31.205 ;
      RECT 135.955 -30.478 136.045 -29.471 ;
      RECT 135.955 -30.165 136.095 -29.995 ;
      RECT 135.955 -28.669 136.045 -27.662 ;
      RECT 135.955 -28.145 136.095 -27.975 ;
      RECT 135.955 -27.248 136.045 -26.241 ;
      RECT 135.955 -26.935 136.095 -26.765 ;
      RECT 135.955 -25.439 136.045 -24.432 ;
      RECT 135.955 -24.915 136.095 -24.745 ;
      RECT 135.955 -24.018 136.045 -23.011 ;
      RECT 135.955 -23.705 136.095 -23.535 ;
      RECT 135.955 -22.209 136.045 -21.202 ;
      RECT 135.955 -21.685 136.095 -21.515 ;
      RECT 135.955 -20.788 136.045 -19.781 ;
      RECT 135.955 -20.475 136.095 -20.305 ;
      RECT 135.955 -18.979 136.045 -17.972 ;
      RECT 135.955 -18.455 136.095 -18.285 ;
      RECT 135.955 -17.558 136.045 -16.551 ;
      RECT 135.955 -17.245 136.095 -17.075 ;
      RECT 135.955 -15.749 136.045 -14.742 ;
      RECT 135.955 -15.225 136.095 -15.055 ;
      RECT 135.955 -14.328 136.045 -13.321 ;
      RECT 135.955 -14.015 136.095 -13.845 ;
      RECT 135.955 -12.519 136.045 -11.512 ;
      RECT 135.955 -11.995 136.095 -11.825 ;
      RECT 135.955 -11.098 136.045 -10.091 ;
      RECT 135.955 -10.785 136.095 -10.615 ;
      RECT 135.955 -9.289 136.045 -8.282 ;
      RECT 135.955 -8.765 136.095 -8.595 ;
      RECT 135.955 -7.868 136.045 -6.861 ;
      RECT 135.955 -7.555 136.095 -7.385 ;
      RECT 135.955 -6.059 136.045 -5.052 ;
      RECT 135.955 -5.535 136.095 -5.365 ;
      RECT 135.955 -4.638 136.045 -3.631 ;
      RECT 135.955 -4.325 136.095 -4.155 ;
      RECT 135.955 -2.829 136.045 -1.822 ;
      RECT 135.955 -2.305 136.095 -2.135 ;
      RECT 135.955 -1.408 136.045 -0.401 ;
      RECT 135.955 -1.095 136.095 -0.925 ;
      RECT 135.955 0.401 136.045 1.408 ;
      RECT 135.955 0.925 136.095 1.095 ;
      RECT 135.64 -114.685 135.81 -114.515 ;
      RECT 135.71 -114.895 135.81 -114.515 ;
      RECT 135.155 -101.538 135.245 -100.53 ;
      RECT 135.105 -100.935 135.245 -100.765 ;
      RECT 135.155 -99.73 135.245 -98.722 ;
      RECT 135.105 -99.495 135.245 -99.325 ;
      RECT 135.155 -98.308 135.245 -97.3 ;
      RECT 135.105 -97.705 135.245 -97.535 ;
      RECT 135.155 -96.5 135.245 -95.492 ;
      RECT 135.105 -96.265 135.245 -96.095 ;
      RECT 135.155 -95.078 135.245 -94.07 ;
      RECT 135.105 -94.475 135.245 -94.305 ;
      RECT 135.155 -93.27 135.245 -92.262 ;
      RECT 135.105 -93.035 135.245 -92.865 ;
      RECT 135.155 -91.848 135.245 -90.84 ;
      RECT 135.105 -91.245 135.245 -91.075 ;
      RECT 135.155 -90.04 135.245 -89.032 ;
      RECT 135.105 -89.805 135.245 -89.635 ;
      RECT 135.155 -88.618 135.245 -87.61 ;
      RECT 135.105 -88.015 135.245 -87.845 ;
      RECT 135.155 -86.81 135.245 -85.802 ;
      RECT 135.105 -86.575 135.245 -86.405 ;
      RECT 135.155 -85.388 135.245 -84.38 ;
      RECT 135.105 -84.785 135.245 -84.615 ;
      RECT 135.155 -83.58 135.245 -82.572 ;
      RECT 135.105 -83.345 135.245 -83.175 ;
      RECT 135.155 -82.158 135.245 -81.15 ;
      RECT 135.105 -81.555 135.245 -81.385 ;
      RECT 135.155 -80.35 135.245 -79.342 ;
      RECT 135.105 -80.115 135.245 -79.945 ;
      RECT 135.155 -78.928 135.245 -77.92 ;
      RECT 135.105 -78.325 135.245 -78.155 ;
      RECT 135.155 -77.12 135.245 -76.112 ;
      RECT 135.105 -76.885 135.245 -76.715 ;
      RECT 135.155 -75.698 135.245 -74.69 ;
      RECT 135.105 -75.095 135.245 -74.925 ;
      RECT 135.155 -73.89 135.245 -72.882 ;
      RECT 135.105 -73.655 135.245 -73.485 ;
      RECT 135.155 -72.468 135.245 -71.46 ;
      RECT 135.105 -71.865 135.245 -71.695 ;
      RECT 135.155 -70.66 135.245 -69.652 ;
      RECT 135.105 -70.425 135.245 -70.255 ;
      RECT 135.155 -69.238 135.245 -68.23 ;
      RECT 135.105 -68.635 135.245 -68.465 ;
      RECT 135.155 -67.43 135.245 -66.422 ;
      RECT 135.105 -67.195 135.245 -67.025 ;
      RECT 135.155 -66.008 135.245 -65 ;
      RECT 135.105 -65.405 135.245 -65.235 ;
      RECT 135.155 -64.2 135.245 -63.192 ;
      RECT 135.105 -63.965 135.245 -63.795 ;
      RECT 135.155 -62.778 135.245 -61.77 ;
      RECT 135.105 -62.175 135.245 -62.005 ;
      RECT 135.155 -60.97 135.245 -59.962 ;
      RECT 135.105 -60.735 135.245 -60.565 ;
      RECT 135.155 -59.548 135.245 -58.54 ;
      RECT 135.105 -58.945 135.245 -58.775 ;
      RECT 135.155 -57.74 135.245 -56.732 ;
      RECT 135.105 -57.505 135.245 -57.335 ;
      RECT 135.155 -56.318 135.245 -55.31 ;
      RECT 135.105 -55.715 135.245 -55.545 ;
      RECT 135.155 -54.51 135.245 -53.502 ;
      RECT 135.105 -54.275 135.245 -54.105 ;
      RECT 135.155 -53.088 135.245 -52.08 ;
      RECT 135.105 -52.485 135.245 -52.315 ;
      RECT 135.155 -51.28 135.245 -50.272 ;
      RECT 135.105 -51.045 135.245 -50.875 ;
      RECT 135.155 -49.858 135.245 -48.85 ;
      RECT 135.105 -49.255 135.245 -49.085 ;
      RECT 135.155 -48.05 135.245 -47.042 ;
      RECT 135.105 -47.815 135.245 -47.645 ;
      RECT 135.155 -46.628 135.245 -45.62 ;
      RECT 135.105 -46.025 135.245 -45.855 ;
      RECT 135.155 -44.82 135.245 -43.812 ;
      RECT 135.105 -44.585 135.245 -44.415 ;
      RECT 135.155 -43.398 135.245 -42.39 ;
      RECT 135.105 -42.795 135.245 -42.625 ;
      RECT 135.155 -41.59 135.245 -40.582 ;
      RECT 135.105 -41.355 135.245 -41.185 ;
      RECT 135.155 -40.168 135.245 -39.16 ;
      RECT 135.105 -39.565 135.245 -39.395 ;
      RECT 135.155 -38.36 135.245 -37.352 ;
      RECT 135.105 -38.125 135.245 -37.955 ;
      RECT 135.155 -36.938 135.245 -35.93 ;
      RECT 135.105 -36.335 135.245 -36.165 ;
      RECT 135.155 -35.13 135.245 -34.122 ;
      RECT 135.105 -34.895 135.245 -34.725 ;
      RECT 135.155 -33.708 135.245 -32.7 ;
      RECT 135.105 -33.105 135.245 -32.935 ;
      RECT 135.155 -31.9 135.245 -30.892 ;
      RECT 135.105 -31.665 135.245 -31.495 ;
      RECT 135.155 -30.478 135.245 -29.47 ;
      RECT 135.105 -29.875 135.245 -29.705 ;
      RECT 135.155 -28.67 135.245 -27.662 ;
      RECT 135.105 -28.435 135.245 -28.265 ;
      RECT 135.155 -27.248 135.245 -26.24 ;
      RECT 135.105 -26.645 135.245 -26.475 ;
      RECT 135.155 -25.44 135.245 -24.432 ;
      RECT 135.105 -25.205 135.245 -25.035 ;
      RECT 135.155 -24.018 135.245 -23.01 ;
      RECT 135.105 -23.415 135.245 -23.245 ;
      RECT 135.155 -22.21 135.245 -21.202 ;
      RECT 135.105 -21.975 135.245 -21.805 ;
      RECT 135.155 -20.788 135.245 -19.78 ;
      RECT 135.105 -20.185 135.245 -20.015 ;
      RECT 135.155 -18.98 135.245 -17.972 ;
      RECT 135.105 -18.745 135.245 -18.575 ;
      RECT 135.155 -17.558 135.245 -16.55 ;
      RECT 135.105 -16.955 135.245 -16.785 ;
      RECT 135.155 -15.75 135.245 -14.742 ;
      RECT 135.105 -15.515 135.245 -15.345 ;
      RECT 135.155 -14.328 135.245 -13.32 ;
      RECT 135.105 -13.725 135.245 -13.555 ;
      RECT 135.155 -12.52 135.245 -11.512 ;
      RECT 135.105 -12.285 135.245 -12.115 ;
      RECT 135.155 -11.098 135.245 -10.09 ;
      RECT 135.105 -10.495 135.245 -10.325 ;
      RECT 135.155 -9.29 135.245 -8.282 ;
      RECT 135.105 -9.055 135.245 -8.885 ;
      RECT 135.155 -7.868 135.245 -6.86 ;
      RECT 135.105 -7.265 135.245 -7.095 ;
      RECT 135.155 -6.06 135.245 -5.052 ;
      RECT 135.105 -5.825 135.245 -5.655 ;
      RECT 135.155 -4.638 135.245 -3.63 ;
      RECT 135.105 -4.035 135.245 -3.865 ;
      RECT 135.155 -2.83 135.245 -1.822 ;
      RECT 135.105 -2.595 135.245 -2.425 ;
      RECT 135.155 -1.408 135.245 -0.4 ;
      RECT 135.105 -0.805 135.245 -0.635 ;
      RECT 135.155 0.4 135.245 1.408 ;
      RECT 135.105 0.635 135.245 0.805 ;
      RECT 134.755 -101.538 134.845 -100.531 ;
      RECT 134.755 -101.225 134.895 -101.055 ;
      RECT 134.755 -99.729 134.845 -98.722 ;
      RECT 134.755 -99.205 134.895 -99.035 ;
      RECT 134.755 -98.308 134.845 -97.301 ;
      RECT 134.755 -97.995 134.895 -97.825 ;
      RECT 134.755 -96.499 134.845 -95.492 ;
      RECT 134.755 -95.975 134.895 -95.805 ;
      RECT 134.755 -95.078 134.845 -94.071 ;
      RECT 134.755 -94.765 134.895 -94.595 ;
      RECT 134.755 -93.269 134.845 -92.262 ;
      RECT 134.755 -92.745 134.895 -92.575 ;
      RECT 134.755 -91.848 134.845 -90.841 ;
      RECT 134.755 -91.535 134.895 -91.365 ;
      RECT 134.755 -90.039 134.845 -89.032 ;
      RECT 134.755 -89.515 134.895 -89.345 ;
      RECT 134.755 -88.618 134.845 -87.611 ;
      RECT 134.755 -88.305 134.895 -88.135 ;
      RECT 134.755 -86.809 134.845 -85.802 ;
      RECT 134.755 -86.285 134.895 -86.115 ;
      RECT 134.755 -85.388 134.845 -84.381 ;
      RECT 134.755 -85.075 134.895 -84.905 ;
      RECT 134.755 -83.579 134.845 -82.572 ;
      RECT 134.755 -83.055 134.895 -82.885 ;
      RECT 134.755 -82.158 134.845 -81.151 ;
      RECT 134.755 -81.845 134.895 -81.675 ;
      RECT 134.755 -80.349 134.845 -79.342 ;
      RECT 134.755 -79.825 134.895 -79.655 ;
      RECT 134.755 -78.928 134.845 -77.921 ;
      RECT 134.755 -78.615 134.895 -78.445 ;
      RECT 134.755 -77.119 134.845 -76.112 ;
      RECT 134.755 -76.595 134.895 -76.425 ;
      RECT 134.755 -75.698 134.845 -74.691 ;
      RECT 134.755 -75.385 134.895 -75.215 ;
      RECT 134.755 -73.889 134.845 -72.882 ;
      RECT 134.755 -73.365 134.895 -73.195 ;
      RECT 134.755 -72.468 134.845 -71.461 ;
      RECT 134.755 -72.155 134.895 -71.985 ;
      RECT 134.755 -70.659 134.845 -69.652 ;
      RECT 134.755 -70.135 134.895 -69.965 ;
      RECT 134.755 -69.238 134.845 -68.231 ;
      RECT 134.755 -68.925 134.895 -68.755 ;
      RECT 134.755 -67.429 134.845 -66.422 ;
      RECT 134.755 -66.905 134.895 -66.735 ;
      RECT 134.755 -66.008 134.845 -65.001 ;
      RECT 134.755 -65.695 134.895 -65.525 ;
      RECT 134.755 -64.199 134.845 -63.192 ;
      RECT 134.755 -63.675 134.895 -63.505 ;
      RECT 134.755 -62.778 134.845 -61.771 ;
      RECT 134.755 -62.465 134.895 -62.295 ;
      RECT 134.755 -60.969 134.845 -59.962 ;
      RECT 134.755 -60.445 134.895 -60.275 ;
      RECT 134.755 -59.548 134.845 -58.541 ;
      RECT 134.755 -59.235 134.895 -59.065 ;
      RECT 134.755 -57.739 134.845 -56.732 ;
      RECT 134.755 -57.215 134.895 -57.045 ;
      RECT 134.755 -56.318 134.845 -55.311 ;
      RECT 134.755 -56.005 134.895 -55.835 ;
      RECT 134.755 -54.509 134.845 -53.502 ;
      RECT 134.755 -53.985 134.895 -53.815 ;
      RECT 134.755 -53.088 134.845 -52.081 ;
      RECT 134.755 -52.775 134.895 -52.605 ;
      RECT 134.755 -51.279 134.845 -50.272 ;
      RECT 134.755 -50.755 134.895 -50.585 ;
      RECT 134.755 -49.858 134.845 -48.851 ;
      RECT 134.755 -49.545 134.895 -49.375 ;
      RECT 134.755 -48.049 134.845 -47.042 ;
      RECT 134.755 -47.525 134.895 -47.355 ;
      RECT 134.755 -46.628 134.845 -45.621 ;
      RECT 134.755 -46.315 134.895 -46.145 ;
      RECT 134.755 -44.819 134.845 -43.812 ;
      RECT 134.755 -44.295 134.895 -44.125 ;
      RECT 134.755 -43.398 134.845 -42.391 ;
      RECT 134.755 -43.085 134.895 -42.915 ;
      RECT 134.755 -41.589 134.845 -40.582 ;
      RECT 134.755 -41.065 134.895 -40.895 ;
      RECT 134.755 -40.168 134.845 -39.161 ;
      RECT 134.755 -39.855 134.895 -39.685 ;
      RECT 134.755 -38.359 134.845 -37.352 ;
      RECT 134.755 -37.835 134.895 -37.665 ;
      RECT 134.755 -36.938 134.845 -35.931 ;
      RECT 134.755 -36.625 134.895 -36.455 ;
      RECT 134.755 -35.129 134.845 -34.122 ;
      RECT 134.755 -34.605 134.895 -34.435 ;
      RECT 134.755 -33.708 134.845 -32.701 ;
      RECT 134.755 -33.395 134.895 -33.225 ;
      RECT 134.755 -31.899 134.845 -30.892 ;
      RECT 134.755 -31.375 134.895 -31.205 ;
      RECT 134.755 -30.478 134.845 -29.471 ;
      RECT 134.755 -30.165 134.895 -29.995 ;
      RECT 134.755 -28.669 134.845 -27.662 ;
      RECT 134.755 -28.145 134.895 -27.975 ;
      RECT 134.755 -27.248 134.845 -26.241 ;
      RECT 134.755 -26.935 134.895 -26.765 ;
      RECT 134.755 -25.439 134.845 -24.432 ;
      RECT 134.755 -24.915 134.895 -24.745 ;
      RECT 134.755 -24.018 134.845 -23.011 ;
      RECT 134.755 -23.705 134.895 -23.535 ;
      RECT 134.755 -22.209 134.845 -21.202 ;
      RECT 134.755 -21.685 134.895 -21.515 ;
      RECT 134.755 -20.788 134.845 -19.781 ;
      RECT 134.755 -20.475 134.895 -20.305 ;
      RECT 134.755 -18.979 134.845 -17.972 ;
      RECT 134.755 -18.455 134.895 -18.285 ;
      RECT 134.755 -17.558 134.845 -16.551 ;
      RECT 134.755 -17.245 134.895 -17.075 ;
      RECT 134.755 -15.749 134.845 -14.742 ;
      RECT 134.755 -15.225 134.895 -15.055 ;
      RECT 134.755 -14.328 134.845 -13.321 ;
      RECT 134.755 -14.015 134.895 -13.845 ;
      RECT 134.755 -12.519 134.845 -11.512 ;
      RECT 134.755 -11.995 134.895 -11.825 ;
      RECT 134.755 -11.098 134.845 -10.091 ;
      RECT 134.755 -10.785 134.895 -10.615 ;
      RECT 134.755 -9.289 134.845 -8.282 ;
      RECT 134.755 -8.765 134.895 -8.595 ;
      RECT 134.755 -7.868 134.845 -6.861 ;
      RECT 134.755 -7.555 134.895 -7.385 ;
      RECT 134.755 -6.059 134.845 -5.052 ;
      RECT 134.755 -5.535 134.895 -5.365 ;
      RECT 134.755 -4.638 134.845 -3.631 ;
      RECT 134.755 -4.325 134.895 -4.155 ;
      RECT 134.755 -2.829 134.845 -1.822 ;
      RECT 134.755 -2.305 134.895 -2.135 ;
      RECT 134.755 -1.408 134.845 -0.401 ;
      RECT 134.755 -1.095 134.895 -0.925 ;
      RECT 134.755 0.401 134.845 1.408 ;
      RECT 134.755 0.925 134.895 1.095 ;
      RECT 130.585 -108.935 134.365 -108.815 ;
      RECT 131.905 -109.475 132.005 -108.815 ;
      RECT 131.345 -109.475 131.445 -108.815 ;
      RECT 130.785 -109.475 130.885 -108.815 ;
      RECT 133.955 -101.538 134.045 -100.53 ;
      RECT 133.905 -100.935 134.045 -100.765 ;
      RECT 133.955 -99.73 134.045 -98.722 ;
      RECT 133.905 -99.495 134.045 -99.325 ;
      RECT 133.955 -98.308 134.045 -97.3 ;
      RECT 133.905 -97.705 134.045 -97.535 ;
      RECT 133.955 -96.5 134.045 -95.492 ;
      RECT 133.905 -96.265 134.045 -96.095 ;
      RECT 133.955 -95.078 134.045 -94.07 ;
      RECT 133.905 -94.475 134.045 -94.305 ;
      RECT 133.955 -93.27 134.045 -92.262 ;
      RECT 133.905 -93.035 134.045 -92.865 ;
      RECT 133.955 -91.848 134.045 -90.84 ;
      RECT 133.905 -91.245 134.045 -91.075 ;
      RECT 133.955 -90.04 134.045 -89.032 ;
      RECT 133.905 -89.805 134.045 -89.635 ;
      RECT 133.955 -88.618 134.045 -87.61 ;
      RECT 133.905 -88.015 134.045 -87.845 ;
      RECT 133.955 -86.81 134.045 -85.802 ;
      RECT 133.905 -86.575 134.045 -86.405 ;
      RECT 133.955 -85.388 134.045 -84.38 ;
      RECT 133.905 -84.785 134.045 -84.615 ;
      RECT 133.955 -83.58 134.045 -82.572 ;
      RECT 133.905 -83.345 134.045 -83.175 ;
      RECT 133.955 -82.158 134.045 -81.15 ;
      RECT 133.905 -81.555 134.045 -81.385 ;
      RECT 133.955 -80.35 134.045 -79.342 ;
      RECT 133.905 -80.115 134.045 -79.945 ;
      RECT 133.955 -78.928 134.045 -77.92 ;
      RECT 133.905 -78.325 134.045 -78.155 ;
      RECT 133.955 -77.12 134.045 -76.112 ;
      RECT 133.905 -76.885 134.045 -76.715 ;
      RECT 133.955 -75.698 134.045 -74.69 ;
      RECT 133.905 -75.095 134.045 -74.925 ;
      RECT 133.955 -73.89 134.045 -72.882 ;
      RECT 133.905 -73.655 134.045 -73.485 ;
      RECT 133.955 -72.468 134.045 -71.46 ;
      RECT 133.905 -71.865 134.045 -71.695 ;
      RECT 133.955 -70.66 134.045 -69.652 ;
      RECT 133.905 -70.425 134.045 -70.255 ;
      RECT 133.955 -69.238 134.045 -68.23 ;
      RECT 133.905 -68.635 134.045 -68.465 ;
      RECT 133.955 -67.43 134.045 -66.422 ;
      RECT 133.905 -67.195 134.045 -67.025 ;
      RECT 133.955 -66.008 134.045 -65 ;
      RECT 133.905 -65.405 134.045 -65.235 ;
      RECT 133.955 -64.2 134.045 -63.192 ;
      RECT 133.905 -63.965 134.045 -63.795 ;
      RECT 133.955 -62.778 134.045 -61.77 ;
      RECT 133.905 -62.175 134.045 -62.005 ;
      RECT 133.955 -60.97 134.045 -59.962 ;
      RECT 133.905 -60.735 134.045 -60.565 ;
      RECT 133.955 -59.548 134.045 -58.54 ;
      RECT 133.905 -58.945 134.045 -58.775 ;
      RECT 133.955 -57.74 134.045 -56.732 ;
      RECT 133.905 -57.505 134.045 -57.335 ;
      RECT 133.955 -56.318 134.045 -55.31 ;
      RECT 133.905 -55.715 134.045 -55.545 ;
      RECT 133.955 -54.51 134.045 -53.502 ;
      RECT 133.905 -54.275 134.045 -54.105 ;
      RECT 133.955 -53.088 134.045 -52.08 ;
      RECT 133.905 -52.485 134.045 -52.315 ;
      RECT 133.955 -51.28 134.045 -50.272 ;
      RECT 133.905 -51.045 134.045 -50.875 ;
      RECT 133.955 -49.858 134.045 -48.85 ;
      RECT 133.905 -49.255 134.045 -49.085 ;
      RECT 133.955 -48.05 134.045 -47.042 ;
      RECT 133.905 -47.815 134.045 -47.645 ;
      RECT 133.955 -46.628 134.045 -45.62 ;
      RECT 133.905 -46.025 134.045 -45.855 ;
      RECT 133.955 -44.82 134.045 -43.812 ;
      RECT 133.905 -44.585 134.045 -44.415 ;
      RECT 133.955 -43.398 134.045 -42.39 ;
      RECT 133.905 -42.795 134.045 -42.625 ;
      RECT 133.955 -41.59 134.045 -40.582 ;
      RECT 133.905 -41.355 134.045 -41.185 ;
      RECT 133.955 -40.168 134.045 -39.16 ;
      RECT 133.905 -39.565 134.045 -39.395 ;
      RECT 133.955 -38.36 134.045 -37.352 ;
      RECT 133.905 -38.125 134.045 -37.955 ;
      RECT 133.955 -36.938 134.045 -35.93 ;
      RECT 133.905 -36.335 134.045 -36.165 ;
      RECT 133.955 -35.13 134.045 -34.122 ;
      RECT 133.905 -34.895 134.045 -34.725 ;
      RECT 133.955 -33.708 134.045 -32.7 ;
      RECT 133.905 -33.105 134.045 -32.935 ;
      RECT 133.955 -31.9 134.045 -30.892 ;
      RECT 133.905 -31.665 134.045 -31.495 ;
      RECT 133.955 -30.478 134.045 -29.47 ;
      RECT 133.905 -29.875 134.045 -29.705 ;
      RECT 133.955 -28.67 134.045 -27.662 ;
      RECT 133.905 -28.435 134.045 -28.265 ;
      RECT 133.955 -27.248 134.045 -26.24 ;
      RECT 133.905 -26.645 134.045 -26.475 ;
      RECT 133.955 -25.44 134.045 -24.432 ;
      RECT 133.905 -25.205 134.045 -25.035 ;
      RECT 133.955 -24.018 134.045 -23.01 ;
      RECT 133.905 -23.415 134.045 -23.245 ;
      RECT 133.955 -22.21 134.045 -21.202 ;
      RECT 133.905 -21.975 134.045 -21.805 ;
      RECT 133.955 -20.788 134.045 -19.78 ;
      RECT 133.905 -20.185 134.045 -20.015 ;
      RECT 133.955 -18.98 134.045 -17.972 ;
      RECT 133.905 -18.745 134.045 -18.575 ;
      RECT 133.955 -17.558 134.045 -16.55 ;
      RECT 133.905 -16.955 134.045 -16.785 ;
      RECT 133.955 -15.75 134.045 -14.742 ;
      RECT 133.905 -15.515 134.045 -15.345 ;
      RECT 133.955 -14.328 134.045 -13.32 ;
      RECT 133.905 -13.725 134.045 -13.555 ;
      RECT 133.955 -12.52 134.045 -11.512 ;
      RECT 133.905 -12.285 134.045 -12.115 ;
      RECT 133.955 -11.098 134.045 -10.09 ;
      RECT 133.905 -10.495 134.045 -10.325 ;
      RECT 133.955 -9.29 134.045 -8.282 ;
      RECT 133.905 -9.055 134.045 -8.885 ;
      RECT 133.955 -7.868 134.045 -6.86 ;
      RECT 133.905 -7.265 134.045 -7.095 ;
      RECT 133.955 -6.06 134.045 -5.052 ;
      RECT 133.905 -5.825 134.045 -5.655 ;
      RECT 133.955 -4.638 134.045 -3.63 ;
      RECT 133.905 -4.035 134.045 -3.865 ;
      RECT 133.955 -2.83 134.045 -1.822 ;
      RECT 133.905 -2.595 134.045 -2.425 ;
      RECT 133.955 -1.408 134.045 -0.4 ;
      RECT 133.905 -0.805 134.045 -0.635 ;
      RECT 133.955 0.4 134.045 1.408 ;
      RECT 133.905 0.635 134.045 0.805 ;
      RECT 132.525 -111.685 134.005 -111.585 ;
      RECT 132.525 -112.195 132.625 -111.585 ;
      RECT 132.745 -109.15 134.005 -109.05 ;
      RECT 133.905 -109.475 134.005 -109.05 ;
      RECT 133.345 -109.475 133.445 -109.05 ;
      RECT 132.785 -109.475 132.885 -109.05 ;
      RECT 133.555 -101.538 133.645 -100.531 ;
      RECT 133.555 -101.225 133.695 -101.055 ;
      RECT 133.555 -99.729 133.645 -98.722 ;
      RECT 133.555 -99.205 133.695 -99.035 ;
      RECT 133.555 -98.308 133.645 -97.301 ;
      RECT 133.555 -97.995 133.695 -97.825 ;
      RECT 133.555 -96.499 133.645 -95.492 ;
      RECT 133.555 -95.975 133.695 -95.805 ;
      RECT 133.555 -95.078 133.645 -94.071 ;
      RECT 133.555 -94.765 133.695 -94.595 ;
      RECT 133.555 -93.269 133.645 -92.262 ;
      RECT 133.555 -92.745 133.695 -92.575 ;
      RECT 133.555 -91.848 133.645 -90.841 ;
      RECT 133.555 -91.535 133.695 -91.365 ;
      RECT 133.555 -90.039 133.645 -89.032 ;
      RECT 133.555 -89.515 133.695 -89.345 ;
      RECT 133.555 -88.618 133.645 -87.611 ;
      RECT 133.555 -88.305 133.695 -88.135 ;
      RECT 133.555 -86.809 133.645 -85.802 ;
      RECT 133.555 -86.285 133.695 -86.115 ;
      RECT 133.555 -85.388 133.645 -84.381 ;
      RECT 133.555 -85.075 133.695 -84.905 ;
      RECT 133.555 -83.579 133.645 -82.572 ;
      RECT 133.555 -83.055 133.695 -82.885 ;
      RECT 133.555 -82.158 133.645 -81.151 ;
      RECT 133.555 -81.845 133.695 -81.675 ;
      RECT 133.555 -80.349 133.645 -79.342 ;
      RECT 133.555 -79.825 133.695 -79.655 ;
      RECT 133.555 -78.928 133.645 -77.921 ;
      RECT 133.555 -78.615 133.695 -78.445 ;
      RECT 133.555 -77.119 133.645 -76.112 ;
      RECT 133.555 -76.595 133.695 -76.425 ;
      RECT 133.555 -75.698 133.645 -74.691 ;
      RECT 133.555 -75.385 133.695 -75.215 ;
      RECT 133.555 -73.889 133.645 -72.882 ;
      RECT 133.555 -73.365 133.695 -73.195 ;
      RECT 133.555 -72.468 133.645 -71.461 ;
      RECT 133.555 -72.155 133.695 -71.985 ;
      RECT 133.555 -70.659 133.645 -69.652 ;
      RECT 133.555 -70.135 133.695 -69.965 ;
      RECT 133.555 -69.238 133.645 -68.231 ;
      RECT 133.555 -68.925 133.695 -68.755 ;
      RECT 133.555 -67.429 133.645 -66.422 ;
      RECT 133.555 -66.905 133.695 -66.735 ;
      RECT 133.555 -66.008 133.645 -65.001 ;
      RECT 133.555 -65.695 133.695 -65.525 ;
      RECT 133.555 -64.199 133.645 -63.192 ;
      RECT 133.555 -63.675 133.695 -63.505 ;
      RECT 133.555 -62.778 133.645 -61.771 ;
      RECT 133.555 -62.465 133.695 -62.295 ;
      RECT 133.555 -60.969 133.645 -59.962 ;
      RECT 133.555 -60.445 133.695 -60.275 ;
      RECT 133.555 -59.548 133.645 -58.541 ;
      RECT 133.555 -59.235 133.695 -59.065 ;
      RECT 133.555 -57.739 133.645 -56.732 ;
      RECT 133.555 -57.215 133.695 -57.045 ;
      RECT 133.555 -56.318 133.645 -55.311 ;
      RECT 133.555 -56.005 133.695 -55.835 ;
      RECT 133.555 -54.509 133.645 -53.502 ;
      RECT 133.555 -53.985 133.695 -53.815 ;
      RECT 133.555 -53.088 133.645 -52.081 ;
      RECT 133.555 -52.775 133.695 -52.605 ;
      RECT 133.555 -51.279 133.645 -50.272 ;
      RECT 133.555 -50.755 133.695 -50.585 ;
      RECT 133.555 -49.858 133.645 -48.851 ;
      RECT 133.555 -49.545 133.695 -49.375 ;
      RECT 133.555 -48.049 133.645 -47.042 ;
      RECT 133.555 -47.525 133.695 -47.355 ;
      RECT 133.555 -46.628 133.645 -45.621 ;
      RECT 133.555 -46.315 133.695 -46.145 ;
      RECT 133.555 -44.819 133.645 -43.812 ;
      RECT 133.555 -44.295 133.695 -44.125 ;
      RECT 133.555 -43.398 133.645 -42.391 ;
      RECT 133.555 -43.085 133.695 -42.915 ;
      RECT 133.555 -41.589 133.645 -40.582 ;
      RECT 133.555 -41.065 133.695 -40.895 ;
      RECT 133.555 -40.168 133.645 -39.161 ;
      RECT 133.555 -39.855 133.695 -39.685 ;
      RECT 133.555 -38.359 133.645 -37.352 ;
      RECT 133.555 -37.835 133.695 -37.665 ;
      RECT 133.555 -36.938 133.645 -35.931 ;
      RECT 133.555 -36.625 133.695 -36.455 ;
      RECT 133.555 -35.129 133.645 -34.122 ;
      RECT 133.555 -34.605 133.695 -34.435 ;
      RECT 133.555 -33.708 133.645 -32.701 ;
      RECT 133.555 -33.395 133.695 -33.225 ;
      RECT 133.555 -31.899 133.645 -30.892 ;
      RECT 133.555 -31.375 133.695 -31.205 ;
      RECT 133.555 -30.478 133.645 -29.471 ;
      RECT 133.555 -30.165 133.695 -29.995 ;
      RECT 133.555 -28.669 133.645 -27.662 ;
      RECT 133.555 -28.145 133.695 -27.975 ;
      RECT 133.555 -27.248 133.645 -26.241 ;
      RECT 133.555 -26.935 133.695 -26.765 ;
      RECT 133.555 -25.439 133.645 -24.432 ;
      RECT 133.555 -24.915 133.695 -24.745 ;
      RECT 133.555 -24.018 133.645 -23.011 ;
      RECT 133.555 -23.705 133.695 -23.535 ;
      RECT 133.555 -22.209 133.645 -21.202 ;
      RECT 133.555 -21.685 133.695 -21.515 ;
      RECT 133.555 -20.788 133.645 -19.781 ;
      RECT 133.555 -20.475 133.695 -20.305 ;
      RECT 133.555 -18.979 133.645 -17.972 ;
      RECT 133.555 -18.455 133.695 -18.285 ;
      RECT 133.555 -17.558 133.645 -16.551 ;
      RECT 133.555 -17.245 133.695 -17.075 ;
      RECT 133.555 -15.749 133.645 -14.742 ;
      RECT 133.555 -15.225 133.695 -15.055 ;
      RECT 133.555 -14.328 133.645 -13.321 ;
      RECT 133.555 -14.015 133.695 -13.845 ;
      RECT 133.555 -12.519 133.645 -11.512 ;
      RECT 133.555 -11.995 133.695 -11.825 ;
      RECT 133.555 -11.098 133.645 -10.091 ;
      RECT 133.555 -10.785 133.695 -10.615 ;
      RECT 133.555 -9.289 133.645 -8.282 ;
      RECT 133.555 -8.765 133.695 -8.595 ;
      RECT 133.555 -7.868 133.645 -6.861 ;
      RECT 133.555 -7.555 133.695 -7.385 ;
      RECT 133.555 -6.059 133.645 -5.052 ;
      RECT 133.555 -5.535 133.695 -5.365 ;
      RECT 133.555 -4.638 133.645 -3.631 ;
      RECT 133.555 -4.325 133.695 -4.155 ;
      RECT 133.555 -2.829 133.645 -1.822 ;
      RECT 133.555 -2.305 133.695 -2.135 ;
      RECT 133.555 -1.408 133.645 -0.401 ;
      RECT 133.555 -1.095 133.695 -0.925 ;
      RECT 133.555 0.401 133.645 1.408 ;
      RECT 133.555 0.925 133.695 1.095 ;
      RECT 132.885 -111.495 133.055 -111.385 ;
      RECT 129.735 -111.495 133.055 -111.395 ;
      RECT 132.755 -101.538 132.845 -100.53 ;
      RECT 132.705 -100.935 132.845 -100.765 ;
      RECT 132.755 -99.73 132.845 -98.722 ;
      RECT 132.705 -99.495 132.845 -99.325 ;
      RECT 132.755 -98.308 132.845 -97.3 ;
      RECT 132.705 -97.705 132.845 -97.535 ;
      RECT 132.755 -96.5 132.845 -95.492 ;
      RECT 132.705 -96.265 132.845 -96.095 ;
      RECT 132.755 -95.078 132.845 -94.07 ;
      RECT 132.705 -94.475 132.845 -94.305 ;
      RECT 132.755 -93.27 132.845 -92.262 ;
      RECT 132.705 -93.035 132.845 -92.865 ;
      RECT 132.755 -91.848 132.845 -90.84 ;
      RECT 132.705 -91.245 132.845 -91.075 ;
      RECT 132.755 -90.04 132.845 -89.032 ;
      RECT 132.705 -89.805 132.845 -89.635 ;
      RECT 132.755 -88.618 132.845 -87.61 ;
      RECT 132.705 -88.015 132.845 -87.845 ;
      RECT 132.755 -86.81 132.845 -85.802 ;
      RECT 132.705 -86.575 132.845 -86.405 ;
      RECT 132.755 -85.388 132.845 -84.38 ;
      RECT 132.705 -84.785 132.845 -84.615 ;
      RECT 132.755 -83.58 132.845 -82.572 ;
      RECT 132.705 -83.345 132.845 -83.175 ;
      RECT 132.755 -82.158 132.845 -81.15 ;
      RECT 132.705 -81.555 132.845 -81.385 ;
      RECT 132.755 -80.35 132.845 -79.342 ;
      RECT 132.705 -80.115 132.845 -79.945 ;
      RECT 132.755 -78.928 132.845 -77.92 ;
      RECT 132.705 -78.325 132.845 -78.155 ;
      RECT 132.755 -77.12 132.845 -76.112 ;
      RECT 132.705 -76.885 132.845 -76.715 ;
      RECT 132.755 -75.698 132.845 -74.69 ;
      RECT 132.705 -75.095 132.845 -74.925 ;
      RECT 132.755 -73.89 132.845 -72.882 ;
      RECT 132.705 -73.655 132.845 -73.485 ;
      RECT 132.755 -72.468 132.845 -71.46 ;
      RECT 132.705 -71.865 132.845 -71.695 ;
      RECT 132.755 -70.66 132.845 -69.652 ;
      RECT 132.705 -70.425 132.845 -70.255 ;
      RECT 132.755 -69.238 132.845 -68.23 ;
      RECT 132.705 -68.635 132.845 -68.465 ;
      RECT 132.755 -67.43 132.845 -66.422 ;
      RECT 132.705 -67.195 132.845 -67.025 ;
      RECT 132.755 -66.008 132.845 -65 ;
      RECT 132.705 -65.405 132.845 -65.235 ;
      RECT 132.755 -64.2 132.845 -63.192 ;
      RECT 132.705 -63.965 132.845 -63.795 ;
      RECT 132.755 -62.778 132.845 -61.77 ;
      RECT 132.705 -62.175 132.845 -62.005 ;
      RECT 132.755 -60.97 132.845 -59.962 ;
      RECT 132.705 -60.735 132.845 -60.565 ;
      RECT 132.755 -59.548 132.845 -58.54 ;
      RECT 132.705 -58.945 132.845 -58.775 ;
      RECT 132.755 -57.74 132.845 -56.732 ;
      RECT 132.705 -57.505 132.845 -57.335 ;
      RECT 132.755 -56.318 132.845 -55.31 ;
      RECT 132.705 -55.715 132.845 -55.545 ;
      RECT 132.755 -54.51 132.845 -53.502 ;
      RECT 132.705 -54.275 132.845 -54.105 ;
      RECT 132.755 -53.088 132.845 -52.08 ;
      RECT 132.705 -52.485 132.845 -52.315 ;
      RECT 132.755 -51.28 132.845 -50.272 ;
      RECT 132.705 -51.045 132.845 -50.875 ;
      RECT 132.755 -49.858 132.845 -48.85 ;
      RECT 132.705 -49.255 132.845 -49.085 ;
      RECT 132.755 -48.05 132.845 -47.042 ;
      RECT 132.705 -47.815 132.845 -47.645 ;
      RECT 132.755 -46.628 132.845 -45.62 ;
      RECT 132.705 -46.025 132.845 -45.855 ;
      RECT 132.755 -44.82 132.845 -43.812 ;
      RECT 132.705 -44.585 132.845 -44.415 ;
      RECT 132.755 -43.398 132.845 -42.39 ;
      RECT 132.705 -42.795 132.845 -42.625 ;
      RECT 132.755 -41.59 132.845 -40.582 ;
      RECT 132.705 -41.355 132.845 -41.185 ;
      RECT 132.755 -40.168 132.845 -39.16 ;
      RECT 132.705 -39.565 132.845 -39.395 ;
      RECT 132.755 -38.36 132.845 -37.352 ;
      RECT 132.705 -38.125 132.845 -37.955 ;
      RECT 132.755 -36.938 132.845 -35.93 ;
      RECT 132.705 -36.335 132.845 -36.165 ;
      RECT 132.755 -35.13 132.845 -34.122 ;
      RECT 132.705 -34.895 132.845 -34.725 ;
      RECT 132.755 -33.708 132.845 -32.7 ;
      RECT 132.705 -33.105 132.845 -32.935 ;
      RECT 132.755 -31.9 132.845 -30.892 ;
      RECT 132.705 -31.665 132.845 -31.495 ;
      RECT 132.755 -30.478 132.845 -29.47 ;
      RECT 132.705 -29.875 132.845 -29.705 ;
      RECT 132.755 -28.67 132.845 -27.662 ;
      RECT 132.705 -28.435 132.845 -28.265 ;
      RECT 132.755 -27.248 132.845 -26.24 ;
      RECT 132.705 -26.645 132.845 -26.475 ;
      RECT 132.755 -25.44 132.845 -24.432 ;
      RECT 132.705 -25.205 132.845 -25.035 ;
      RECT 132.755 -24.018 132.845 -23.01 ;
      RECT 132.705 -23.415 132.845 -23.245 ;
      RECT 132.755 -22.21 132.845 -21.202 ;
      RECT 132.705 -21.975 132.845 -21.805 ;
      RECT 132.755 -20.788 132.845 -19.78 ;
      RECT 132.705 -20.185 132.845 -20.015 ;
      RECT 132.755 -18.98 132.845 -17.972 ;
      RECT 132.705 -18.745 132.845 -18.575 ;
      RECT 132.755 -17.558 132.845 -16.55 ;
      RECT 132.705 -16.955 132.845 -16.785 ;
      RECT 132.755 -15.75 132.845 -14.742 ;
      RECT 132.705 -15.515 132.845 -15.345 ;
      RECT 132.755 -14.328 132.845 -13.32 ;
      RECT 132.705 -13.725 132.845 -13.555 ;
      RECT 132.755 -12.52 132.845 -11.512 ;
      RECT 132.705 -12.285 132.845 -12.115 ;
      RECT 132.755 -11.098 132.845 -10.09 ;
      RECT 132.705 -10.495 132.845 -10.325 ;
      RECT 132.755 -9.29 132.845 -8.282 ;
      RECT 132.705 -9.055 132.845 -8.885 ;
      RECT 132.755 -7.868 132.845 -6.86 ;
      RECT 132.705 -7.265 132.845 -7.095 ;
      RECT 132.755 -6.06 132.845 -5.052 ;
      RECT 132.705 -5.825 132.845 -5.655 ;
      RECT 132.755 -4.638 132.845 -3.63 ;
      RECT 132.705 -4.035 132.845 -3.865 ;
      RECT 132.755 -2.83 132.845 -1.822 ;
      RECT 132.705 -2.595 132.845 -2.425 ;
      RECT 132.755 -1.408 132.845 -0.4 ;
      RECT 132.705 -0.805 132.845 -0.635 ;
      RECT 132.755 0.4 132.845 1.408 ;
      RECT 132.705 0.635 132.845 0.805 ;
      RECT 132.355 -101.538 132.445 -100.531 ;
      RECT 132.355 -101.225 132.495 -101.055 ;
      RECT 132.355 -99.729 132.445 -98.722 ;
      RECT 132.355 -99.205 132.495 -99.035 ;
      RECT 132.355 -98.308 132.445 -97.301 ;
      RECT 132.355 -97.995 132.495 -97.825 ;
      RECT 132.355 -96.499 132.445 -95.492 ;
      RECT 132.355 -95.975 132.495 -95.805 ;
      RECT 132.355 -95.078 132.445 -94.071 ;
      RECT 132.355 -94.765 132.495 -94.595 ;
      RECT 132.355 -93.269 132.445 -92.262 ;
      RECT 132.355 -92.745 132.495 -92.575 ;
      RECT 132.355 -91.848 132.445 -90.841 ;
      RECT 132.355 -91.535 132.495 -91.365 ;
      RECT 132.355 -90.039 132.445 -89.032 ;
      RECT 132.355 -89.515 132.495 -89.345 ;
      RECT 132.355 -88.618 132.445 -87.611 ;
      RECT 132.355 -88.305 132.495 -88.135 ;
      RECT 132.355 -86.809 132.445 -85.802 ;
      RECT 132.355 -86.285 132.495 -86.115 ;
      RECT 132.355 -85.388 132.445 -84.381 ;
      RECT 132.355 -85.075 132.495 -84.905 ;
      RECT 132.355 -83.579 132.445 -82.572 ;
      RECT 132.355 -83.055 132.495 -82.885 ;
      RECT 132.355 -82.158 132.445 -81.151 ;
      RECT 132.355 -81.845 132.495 -81.675 ;
      RECT 132.355 -80.349 132.445 -79.342 ;
      RECT 132.355 -79.825 132.495 -79.655 ;
      RECT 132.355 -78.928 132.445 -77.921 ;
      RECT 132.355 -78.615 132.495 -78.445 ;
      RECT 132.355 -77.119 132.445 -76.112 ;
      RECT 132.355 -76.595 132.495 -76.425 ;
      RECT 132.355 -75.698 132.445 -74.691 ;
      RECT 132.355 -75.385 132.495 -75.215 ;
      RECT 132.355 -73.889 132.445 -72.882 ;
      RECT 132.355 -73.365 132.495 -73.195 ;
      RECT 132.355 -72.468 132.445 -71.461 ;
      RECT 132.355 -72.155 132.495 -71.985 ;
      RECT 132.355 -70.659 132.445 -69.652 ;
      RECT 132.355 -70.135 132.495 -69.965 ;
      RECT 132.355 -69.238 132.445 -68.231 ;
      RECT 132.355 -68.925 132.495 -68.755 ;
      RECT 132.355 -67.429 132.445 -66.422 ;
      RECT 132.355 -66.905 132.495 -66.735 ;
      RECT 132.355 -66.008 132.445 -65.001 ;
      RECT 132.355 -65.695 132.495 -65.525 ;
      RECT 132.355 -64.199 132.445 -63.192 ;
      RECT 132.355 -63.675 132.495 -63.505 ;
      RECT 132.355 -62.778 132.445 -61.771 ;
      RECT 132.355 -62.465 132.495 -62.295 ;
      RECT 132.355 -60.969 132.445 -59.962 ;
      RECT 132.355 -60.445 132.495 -60.275 ;
      RECT 132.355 -59.548 132.445 -58.541 ;
      RECT 132.355 -59.235 132.495 -59.065 ;
      RECT 132.355 -57.739 132.445 -56.732 ;
      RECT 132.355 -57.215 132.495 -57.045 ;
      RECT 132.355 -56.318 132.445 -55.311 ;
      RECT 132.355 -56.005 132.495 -55.835 ;
      RECT 132.355 -54.509 132.445 -53.502 ;
      RECT 132.355 -53.985 132.495 -53.815 ;
      RECT 132.355 -53.088 132.445 -52.081 ;
      RECT 132.355 -52.775 132.495 -52.605 ;
      RECT 132.355 -51.279 132.445 -50.272 ;
      RECT 132.355 -50.755 132.495 -50.585 ;
      RECT 132.355 -49.858 132.445 -48.851 ;
      RECT 132.355 -49.545 132.495 -49.375 ;
      RECT 132.355 -48.049 132.445 -47.042 ;
      RECT 132.355 -47.525 132.495 -47.355 ;
      RECT 132.355 -46.628 132.445 -45.621 ;
      RECT 132.355 -46.315 132.495 -46.145 ;
      RECT 132.355 -44.819 132.445 -43.812 ;
      RECT 132.355 -44.295 132.495 -44.125 ;
      RECT 132.355 -43.398 132.445 -42.391 ;
      RECT 132.355 -43.085 132.495 -42.915 ;
      RECT 132.355 -41.589 132.445 -40.582 ;
      RECT 132.355 -41.065 132.495 -40.895 ;
      RECT 132.355 -40.168 132.445 -39.161 ;
      RECT 132.355 -39.855 132.495 -39.685 ;
      RECT 132.355 -38.359 132.445 -37.352 ;
      RECT 132.355 -37.835 132.495 -37.665 ;
      RECT 132.355 -36.938 132.445 -35.931 ;
      RECT 132.355 -36.625 132.495 -36.455 ;
      RECT 132.355 -35.129 132.445 -34.122 ;
      RECT 132.355 -34.605 132.495 -34.435 ;
      RECT 132.355 -33.708 132.445 -32.701 ;
      RECT 132.355 -33.395 132.495 -33.225 ;
      RECT 132.355 -31.899 132.445 -30.892 ;
      RECT 132.355 -31.375 132.495 -31.205 ;
      RECT 132.355 -30.478 132.445 -29.471 ;
      RECT 132.355 -30.165 132.495 -29.995 ;
      RECT 132.355 -28.669 132.445 -27.662 ;
      RECT 132.355 -28.145 132.495 -27.975 ;
      RECT 132.355 -27.248 132.445 -26.241 ;
      RECT 132.355 -26.935 132.495 -26.765 ;
      RECT 132.355 -25.439 132.445 -24.432 ;
      RECT 132.355 -24.915 132.495 -24.745 ;
      RECT 132.355 -24.018 132.445 -23.011 ;
      RECT 132.355 -23.705 132.495 -23.535 ;
      RECT 132.355 -22.209 132.445 -21.202 ;
      RECT 132.355 -21.685 132.495 -21.515 ;
      RECT 132.355 -20.788 132.445 -19.781 ;
      RECT 132.355 -20.475 132.495 -20.305 ;
      RECT 132.355 -18.979 132.445 -17.972 ;
      RECT 132.355 -18.455 132.495 -18.285 ;
      RECT 132.355 -17.558 132.445 -16.551 ;
      RECT 132.355 -17.245 132.495 -17.075 ;
      RECT 132.355 -15.749 132.445 -14.742 ;
      RECT 132.355 -15.225 132.495 -15.055 ;
      RECT 132.355 -14.328 132.445 -13.321 ;
      RECT 132.355 -14.015 132.495 -13.845 ;
      RECT 132.355 -12.519 132.445 -11.512 ;
      RECT 132.355 -11.995 132.495 -11.825 ;
      RECT 132.355 -11.098 132.445 -10.091 ;
      RECT 132.355 -10.785 132.495 -10.615 ;
      RECT 132.355 -9.289 132.445 -8.282 ;
      RECT 132.355 -8.765 132.495 -8.595 ;
      RECT 132.355 -7.868 132.445 -6.861 ;
      RECT 132.355 -7.555 132.495 -7.385 ;
      RECT 132.355 -6.059 132.445 -5.052 ;
      RECT 132.355 -5.535 132.495 -5.365 ;
      RECT 132.355 -4.638 132.445 -3.631 ;
      RECT 132.355 -4.325 132.495 -4.155 ;
      RECT 132.355 -2.829 132.445 -1.822 ;
      RECT 132.355 -2.305 132.495 -2.135 ;
      RECT 132.355 -1.408 132.445 -0.401 ;
      RECT 132.355 -1.095 132.495 -0.925 ;
      RECT 132.355 0.401 132.445 1.408 ;
      RECT 132.355 0.925 132.495 1.095 ;
      RECT 130.505 -111.685 131.985 -111.585 ;
      RECT 130.505 -112.055 130.605 -111.585 ;
      RECT 130.31 -114.395 131.885 -114.275 ;
      RECT 131.785 -114.895 131.885 -114.275 ;
      RECT 131.19 -114.895 131.29 -114.275 ;
      RECT 130.31 -114.85 130.41 -114.275 ;
      RECT 131.555 -101.538 131.645 -100.53 ;
      RECT 131.505 -100.935 131.645 -100.765 ;
      RECT 131.555 -99.73 131.645 -98.722 ;
      RECT 131.505 -99.495 131.645 -99.325 ;
      RECT 131.555 -98.308 131.645 -97.3 ;
      RECT 131.505 -97.705 131.645 -97.535 ;
      RECT 131.555 -96.5 131.645 -95.492 ;
      RECT 131.505 -96.265 131.645 -96.095 ;
      RECT 131.555 -95.078 131.645 -94.07 ;
      RECT 131.505 -94.475 131.645 -94.305 ;
      RECT 131.555 -93.27 131.645 -92.262 ;
      RECT 131.505 -93.035 131.645 -92.865 ;
      RECT 131.555 -91.848 131.645 -90.84 ;
      RECT 131.505 -91.245 131.645 -91.075 ;
      RECT 131.555 -90.04 131.645 -89.032 ;
      RECT 131.505 -89.805 131.645 -89.635 ;
      RECT 131.555 -88.618 131.645 -87.61 ;
      RECT 131.505 -88.015 131.645 -87.845 ;
      RECT 131.555 -86.81 131.645 -85.802 ;
      RECT 131.505 -86.575 131.645 -86.405 ;
      RECT 131.555 -85.388 131.645 -84.38 ;
      RECT 131.505 -84.785 131.645 -84.615 ;
      RECT 131.555 -83.58 131.645 -82.572 ;
      RECT 131.505 -83.345 131.645 -83.175 ;
      RECT 131.555 -82.158 131.645 -81.15 ;
      RECT 131.505 -81.555 131.645 -81.385 ;
      RECT 131.555 -80.35 131.645 -79.342 ;
      RECT 131.505 -80.115 131.645 -79.945 ;
      RECT 131.555 -78.928 131.645 -77.92 ;
      RECT 131.505 -78.325 131.645 -78.155 ;
      RECT 131.555 -77.12 131.645 -76.112 ;
      RECT 131.505 -76.885 131.645 -76.715 ;
      RECT 131.555 -75.698 131.645 -74.69 ;
      RECT 131.505 -75.095 131.645 -74.925 ;
      RECT 131.555 -73.89 131.645 -72.882 ;
      RECT 131.505 -73.655 131.645 -73.485 ;
      RECT 131.555 -72.468 131.645 -71.46 ;
      RECT 131.505 -71.865 131.645 -71.695 ;
      RECT 131.555 -70.66 131.645 -69.652 ;
      RECT 131.505 -70.425 131.645 -70.255 ;
      RECT 131.555 -69.238 131.645 -68.23 ;
      RECT 131.505 -68.635 131.645 -68.465 ;
      RECT 131.555 -67.43 131.645 -66.422 ;
      RECT 131.505 -67.195 131.645 -67.025 ;
      RECT 131.555 -66.008 131.645 -65 ;
      RECT 131.505 -65.405 131.645 -65.235 ;
      RECT 131.555 -64.2 131.645 -63.192 ;
      RECT 131.505 -63.965 131.645 -63.795 ;
      RECT 131.555 -62.778 131.645 -61.77 ;
      RECT 131.505 -62.175 131.645 -62.005 ;
      RECT 131.555 -60.97 131.645 -59.962 ;
      RECT 131.505 -60.735 131.645 -60.565 ;
      RECT 131.555 -59.548 131.645 -58.54 ;
      RECT 131.505 -58.945 131.645 -58.775 ;
      RECT 131.555 -57.74 131.645 -56.732 ;
      RECT 131.505 -57.505 131.645 -57.335 ;
      RECT 131.555 -56.318 131.645 -55.31 ;
      RECT 131.505 -55.715 131.645 -55.545 ;
      RECT 131.555 -54.51 131.645 -53.502 ;
      RECT 131.505 -54.275 131.645 -54.105 ;
      RECT 131.555 -53.088 131.645 -52.08 ;
      RECT 131.505 -52.485 131.645 -52.315 ;
      RECT 131.555 -51.28 131.645 -50.272 ;
      RECT 131.505 -51.045 131.645 -50.875 ;
      RECT 131.555 -49.858 131.645 -48.85 ;
      RECT 131.505 -49.255 131.645 -49.085 ;
      RECT 131.555 -48.05 131.645 -47.042 ;
      RECT 131.505 -47.815 131.645 -47.645 ;
      RECT 131.555 -46.628 131.645 -45.62 ;
      RECT 131.505 -46.025 131.645 -45.855 ;
      RECT 131.555 -44.82 131.645 -43.812 ;
      RECT 131.505 -44.585 131.645 -44.415 ;
      RECT 131.555 -43.398 131.645 -42.39 ;
      RECT 131.505 -42.795 131.645 -42.625 ;
      RECT 131.555 -41.59 131.645 -40.582 ;
      RECT 131.505 -41.355 131.645 -41.185 ;
      RECT 131.555 -40.168 131.645 -39.16 ;
      RECT 131.505 -39.565 131.645 -39.395 ;
      RECT 131.555 -38.36 131.645 -37.352 ;
      RECT 131.505 -38.125 131.645 -37.955 ;
      RECT 131.555 -36.938 131.645 -35.93 ;
      RECT 131.505 -36.335 131.645 -36.165 ;
      RECT 131.555 -35.13 131.645 -34.122 ;
      RECT 131.505 -34.895 131.645 -34.725 ;
      RECT 131.555 -33.708 131.645 -32.7 ;
      RECT 131.505 -33.105 131.645 -32.935 ;
      RECT 131.555 -31.9 131.645 -30.892 ;
      RECT 131.505 -31.665 131.645 -31.495 ;
      RECT 131.555 -30.478 131.645 -29.47 ;
      RECT 131.505 -29.875 131.645 -29.705 ;
      RECT 131.555 -28.67 131.645 -27.662 ;
      RECT 131.505 -28.435 131.645 -28.265 ;
      RECT 131.555 -27.248 131.645 -26.24 ;
      RECT 131.505 -26.645 131.645 -26.475 ;
      RECT 131.555 -25.44 131.645 -24.432 ;
      RECT 131.505 -25.205 131.645 -25.035 ;
      RECT 131.555 -24.018 131.645 -23.01 ;
      RECT 131.505 -23.415 131.645 -23.245 ;
      RECT 131.555 -22.21 131.645 -21.202 ;
      RECT 131.505 -21.975 131.645 -21.805 ;
      RECT 131.555 -20.788 131.645 -19.78 ;
      RECT 131.505 -20.185 131.645 -20.015 ;
      RECT 131.555 -18.98 131.645 -17.972 ;
      RECT 131.505 -18.745 131.645 -18.575 ;
      RECT 131.555 -17.558 131.645 -16.55 ;
      RECT 131.505 -16.955 131.645 -16.785 ;
      RECT 131.555 -15.75 131.645 -14.742 ;
      RECT 131.505 -15.515 131.645 -15.345 ;
      RECT 131.555 -14.328 131.645 -13.32 ;
      RECT 131.505 -13.725 131.645 -13.555 ;
      RECT 131.555 -12.52 131.645 -11.512 ;
      RECT 131.505 -12.285 131.645 -12.115 ;
      RECT 131.555 -11.098 131.645 -10.09 ;
      RECT 131.505 -10.495 131.645 -10.325 ;
      RECT 131.555 -9.29 131.645 -8.282 ;
      RECT 131.505 -9.055 131.645 -8.885 ;
      RECT 131.555 -7.868 131.645 -6.86 ;
      RECT 131.505 -7.265 131.645 -7.095 ;
      RECT 131.555 -6.06 131.645 -5.052 ;
      RECT 131.505 -5.825 131.645 -5.655 ;
      RECT 131.555 -4.638 131.645 -3.63 ;
      RECT 131.505 -4.035 131.645 -3.865 ;
      RECT 131.555 -2.83 131.645 -1.822 ;
      RECT 131.505 -2.595 131.645 -2.425 ;
      RECT 131.555 -1.408 131.645 -0.4 ;
      RECT 131.505 -0.805 131.645 -0.635 ;
      RECT 131.555 0.4 131.645 1.408 ;
      RECT 131.505 0.635 131.645 0.805 ;
      RECT 131.43 -114.685 131.605 -114.515 ;
      RECT 131.505 -114.895 131.605 -114.515 ;
      RECT 130.545 -113.555 130.645 -113.09 ;
      RECT 130.91 -113.555 131.01 -113.1 ;
      RECT 130.545 -113.555 131.39 -113.385 ;
      RECT 131.155 -101.538 131.245 -100.531 ;
      RECT 131.155 -101.225 131.295 -101.055 ;
      RECT 131.155 -99.729 131.245 -98.722 ;
      RECT 131.155 -99.205 131.295 -99.035 ;
      RECT 131.155 -98.308 131.245 -97.301 ;
      RECT 131.155 -97.995 131.295 -97.825 ;
      RECT 131.155 -96.499 131.245 -95.492 ;
      RECT 131.155 -95.975 131.295 -95.805 ;
      RECT 131.155 -95.078 131.245 -94.071 ;
      RECT 131.155 -94.765 131.295 -94.595 ;
      RECT 131.155 -93.269 131.245 -92.262 ;
      RECT 131.155 -92.745 131.295 -92.575 ;
      RECT 131.155 -91.848 131.245 -90.841 ;
      RECT 131.155 -91.535 131.295 -91.365 ;
      RECT 131.155 -90.039 131.245 -89.032 ;
      RECT 131.155 -89.515 131.295 -89.345 ;
      RECT 131.155 -88.618 131.245 -87.611 ;
      RECT 131.155 -88.305 131.295 -88.135 ;
      RECT 131.155 -86.809 131.245 -85.802 ;
      RECT 131.155 -86.285 131.295 -86.115 ;
      RECT 131.155 -85.388 131.245 -84.381 ;
      RECT 131.155 -85.075 131.295 -84.905 ;
      RECT 131.155 -83.579 131.245 -82.572 ;
      RECT 131.155 -83.055 131.295 -82.885 ;
      RECT 131.155 -82.158 131.245 -81.151 ;
      RECT 131.155 -81.845 131.295 -81.675 ;
      RECT 131.155 -80.349 131.245 -79.342 ;
      RECT 131.155 -79.825 131.295 -79.655 ;
      RECT 131.155 -78.928 131.245 -77.921 ;
      RECT 131.155 -78.615 131.295 -78.445 ;
      RECT 131.155 -77.119 131.245 -76.112 ;
      RECT 131.155 -76.595 131.295 -76.425 ;
      RECT 131.155 -75.698 131.245 -74.691 ;
      RECT 131.155 -75.385 131.295 -75.215 ;
      RECT 131.155 -73.889 131.245 -72.882 ;
      RECT 131.155 -73.365 131.295 -73.195 ;
      RECT 131.155 -72.468 131.245 -71.461 ;
      RECT 131.155 -72.155 131.295 -71.985 ;
      RECT 131.155 -70.659 131.245 -69.652 ;
      RECT 131.155 -70.135 131.295 -69.965 ;
      RECT 131.155 -69.238 131.245 -68.231 ;
      RECT 131.155 -68.925 131.295 -68.755 ;
      RECT 131.155 -67.429 131.245 -66.422 ;
      RECT 131.155 -66.905 131.295 -66.735 ;
      RECT 131.155 -66.008 131.245 -65.001 ;
      RECT 131.155 -65.695 131.295 -65.525 ;
      RECT 131.155 -64.199 131.245 -63.192 ;
      RECT 131.155 -63.675 131.295 -63.505 ;
      RECT 131.155 -62.778 131.245 -61.771 ;
      RECT 131.155 -62.465 131.295 -62.295 ;
      RECT 131.155 -60.969 131.245 -59.962 ;
      RECT 131.155 -60.445 131.295 -60.275 ;
      RECT 131.155 -59.548 131.245 -58.541 ;
      RECT 131.155 -59.235 131.295 -59.065 ;
      RECT 131.155 -57.739 131.245 -56.732 ;
      RECT 131.155 -57.215 131.295 -57.045 ;
      RECT 131.155 -56.318 131.245 -55.311 ;
      RECT 131.155 -56.005 131.295 -55.835 ;
      RECT 131.155 -54.509 131.245 -53.502 ;
      RECT 131.155 -53.985 131.295 -53.815 ;
      RECT 131.155 -53.088 131.245 -52.081 ;
      RECT 131.155 -52.775 131.295 -52.605 ;
      RECT 131.155 -51.279 131.245 -50.272 ;
      RECT 131.155 -50.755 131.295 -50.585 ;
      RECT 131.155 -49.858 131.245 -48.851 ;
      RECT 131.155 -49.545 131.295 -49.375 ;
      RECT 131.155 -48.049 131.245 -47.042 ;
      RECT 131.155 -47.525 131.295 -47.355 ;
      RECT 131.155 -46.628 131.245 -45.621 ;
      RECT 131.155 -46.315 131.295 -46.145 ;
      RECT 131.155 -44.819 131.245 -43.812 ;
      RECT 131.155 -44.295 131.295 -44.125 ;
      RECT 131.155 -43.398 131.245 -42.391 ;
      RECT 131.155 -43.085 131.295 -42.915 ;
      RECT 131.155 -41.589 131.245 -40.582 ;
      RECT 131.155 -41.065 131.295 -40.895 ;
      RECT 131.155 -40.168 131.245 -39.161 ;
      RECT 131.155 -39.855 131.295 -39.685 ;
      RECT 131.155 -38.359 131.245 -37.352 ;
      RECT 131.155 -37.835 131.295 -37.665 ;
      RECT 131.155 -36.938 131.245 -35.931 ;
      RECT 131.155 -36.625 131.295 -36.455 ;
      RECT 131.155 -35.129 131.245 -34.122 ;
      RECT 131.155 -34.605 131.295 -34.435 ;
      RECT 131.155 -33.708 131.245 -32.701 ;
      RECT 131.155 -33.395 131.295 -33.225 ;
      RECT 131.155 -31.899 131.245 -30.892 ;
      RECT 131.155 -31.375 131.295 -31.205 ;
      RECT 131.155 -30.478 131.245 -29.471 ;
      RECT 131.155 -30.165 131.295 -29.995 ;
      RECT 131.155 -28.669 131.245 -27.662 ;
      RECT 131.155 -28.145 131.295 -27.975 ;
      RECT 131.155 -27.248 131.245 -26.241 ;
      RECT 131.155 -26.935 131.295 -26.765 ;
      RECT 131.155 -25.439 131.245 -24.432 ;
      RECT 131.155 -24.915 131.295 -24.745 ;
      RECT 131.155 -24.018 131.245 -23.011 ;
      RECT 131.155 -23.705 131.295 -23.535 ;
      RECT 131.155 -22.209 131.245 -21.202 ;
      RECT 131.155 -21.685 131.295 -21.515 ;
      RECT 131.155 -20.788 131.245 -19.781 ;
      RECT 131.155 -20.475 131.295 -20.305 ;
      RECT 131.155 -18.979 131.245 -17.972 ;
      RECT 131.155 -18.455 131.295 -18.285 ;
      RECT 131.155 -17.558 131.245 -16.551 ;
      RECT 131.155 -17.245 131.295 -17.075 ;
      RECT 131.155 -15.749 131.245 -14.742 ;
      RECT 131.155 -15.225 131.295 -15.055 ;
      RECT 131.155 -14.328 131.245 -13.321 ;
      RECT 131.155 -14.015 131.295 -13.845 ;
      RECT 131.155 -12.519 131.245 -11.512 ;
      RECT 131.155 -11.995 131.295 -11.825 ;
      RECT 131.155 -11.098 131.245 -10.091 ;
      RECT 131.155 -10.785 131.295 -10.615 ;
      RECT 131.155 -9.289 131.245 -8.282 ;
      RECT 131.155 -8.765 131.295 -8.595 ;
      RECT 131.155 -7.868 131.245 -6.861 ;
      RECT 131.155 -7.555 131.295 -7.385 ;
      RECT 131.155 -6.059 131.245 -5.052 ;
      RECT 131.155 -5.535 131.295 -5.365 ;
      RECT 131.155 -4.638 131.245 -3.631 ;
      RECT 131.155 -4.325 131.295 -4.155 ;
      RECT 131.155 -2.829 131.245 -1.822 ;
      RECT 131.155 -2.305 131.295 -2.135 ;
      RECT 131.155 -1.408 131.245 -0.401 ;
      RECT 131.155 -1.095 131.295 -0.925 ;
      RECT 131.155 0.401 131.245 1.408 ;
      RECT 131.155 0.925 131.295 1.095 ;
      RECT 130.84 -114.685 131.01 -114.515 ;
      RECT 130.91 -114.895 131.01 -114.515 ;
      RECT 130.355 -101.538 130.445 -100.53 ;
      RECT 130.305 -100.935 130.445 -100.765 ;
      RECT 130.355 -99.73 130.445 -98.722 ;
      RECT 130.305 -99.495 130.445 -99.325 ;
      RECT 130.355 -98.308 130.445 -97.3 ;
      RECT 130.305 -97.705 130.445 -97.535 ;
      RECT 130.355 -96.5 130.445 -95.492 ;
      RECT 130.305 -96.265 130.445 -96.095 ;
      RECT 130.355 -95.078 130.445 -94.07 ;
      RECT 130.305 -94.475 130.445 -94.305 ;
      RECT 130.355 -93.27 130.445 -92.262 ;
      RECT 130.305 -93.035 130.445 -92.865 ;
      RECT 130.355 -91.848 130.445 -90.84 ;
      RECT 130.305 -91.245 130.445 -91.075 ;
      RECT 130.355 -90.04 130.445 -89.032 ;
      RECT 130.305 -89.805 130.445 -89.635 ;
      RECT 130.355 -88.618 130.445 -87.61 ;
      RECT 130.305 -88.015 130.445 -87.845 ;
      RECT 130.355 -86.81 130.445 -85.802 ;
      RECT 130.305 -86.575 130.445 -86.405 ;
      RECT 130.355 -85.388 130.445 -84.38 ;
      RECT 130.305 -84.785 130.445 -84.615 ;
      RECT 130.355 -83.58 130.445 -82.572 ;
      RECT 130.305 -83.345 130.445 -83.175 ;
      RECT 130.355 -82.158 130.445 -81.15 ;
      RECT 130.305 -81.555 130.445 -81.385 ;
      RECT 130.355 -80.35 130.445 -79.342 ;
      RECT 130.305 -80.115 130.445 -79.945 ;
      RECT 130.355 -78.928 130.445 -77.92 ;
      RECT 130.305 -78.325 130.445 -78.155 ;
      RECT 130.355 -77.12 130.445 -76.112 ;
      RECT 130.305 -76.885 130.445 -76.715 ;
      RECT 130.355 -75.698 130.445 -74.69 ;
      RECT 130.305 -75.095 130.445 -74.925 ;
      RECT 130.355 -73.89 130.445 -72.882 ;
      RECT 130.305 -73.655 130.445 -73.485 ;
      RECT 130.355 -72.468 130.445 -71.46 ;
      RECT 130.305 -71.865 130.445 -71.695 ;
      RECT 130.355 -70.66 130.445 -69.652 ;
      RECT 130.305 -70.425 130.445 -70.255 ;
      RECT 130.355 -69.238 130.445 -68.23 ;
      RECT 130.305 -68.635 130.445 -68.465 ;
      RECT 130.355 -67.43 130.445 -66.422 ;
      RECT 130.305 -67.195 130.445 -67.025 ;
      RECT 130.355 -66.008 130.445 -65 ;
      RECT 130.305 -65.405 130.445 -65.235 ;
      RECT 130.355 -64.2 130.445 -63.192 ;
      RECT 130.305 -63.965 130.445 -63.795 ;
      RECT 130.355 -62.778 130.445 -61.77 ;
      RECT 130.305 -62.175 130.445 -62.005 ;
      RECT 130.355 -60.97 130.445 -59.962 ;
      RECT 130.305 -60.735 130.445 -60.565 ;
      RECT 130.355 -59.548 130.445 -58.54 ;
      RECT 130.305 -58.945 130.445 -58.775 ;
      RECT 130.355 -57.74 130.445 -56.732 ;
      RECT 130.305 -57.505 130.445 -57.335 ;
      RECT 130.355 -56.318 130.445 -55.31 ;
      RECT 130.305 -55.715 130.445 -55.545 ;
      RECT 130.355 -54.51 130.445 -53.502 ;
      RECT 130.305 -54.275 130.445 -54.105 ;
      RECT 130.355 -53.088 130.445 -52.08 ;
      RECT 130.305 -52.485 130.445 -52.315 ;
      RECT 130.355 -51.28 130.445 -50.272 ;
      RECT 130.305 -51.045 130.445 -50.875 ;
      RECT 130.355 -49.858 130.445 -48.85 ;
      RECT 130.305 -49.255 130.445 -49.085 ;
      RECT 130.355 -48.05 130.445 -47.042 ;
      RECT 130.305 -47.815 130.445 -47.645 ;
      RECT 130.355 -46.628 130.445 -45.62 ;
      RECT 130.305 -46.025 130.445 -45.855 ;
      RECT 130.355 -44.82 130.445 -43.812 ;
      RECT 130.305 -44.585 130.445 -44.415 ;
      RECT 130.355 -43.398 130.445 -42.39 ;
      RECT 130.305 -42.795 130.445 -42.625 ;
      RECT 130.355 -41.59 130.445 -40.582 ;
      RECT 130.305 -41.355 130.445 -41.185 ;
      RECT 130.355 -40.168 130.445 -39.16 ;
      RECT 130.305 -39.565 130.445 -39.395 ;
      RECT 130.355 -38.36 130.445 -37.352 ;
      RECT 130.305 -38.125 130.445 -37.955 ;
      RECT 130.355 -36.938 130.445 -35.93 ;
      RECT 130.305 -36.335 130.445 -36.165 ;
      RECT 130.355 -35.13 130.445 -34.122 ;
      RECT 130.305 -34.895 130.445 -34.725 ;
      RECT 130.355 -33.708 130.445 -32.7 ;
      RECT 130.305 -33.105 130.445 -32.935 ;
      RECT 130.355 -31.9 130.445 -30.892 ;
      RECT 130.305 -31.665 130.445 -31.495 ;
      RECT 130.355 -30.478 130.445 -29.47 ;
      RECT 130.305 -29.875 130.445 -29.705 ;
      RECT 130.355 -28.67 130.445 -27.662 ;
      RECT 130.305 -28.435 130.445 -28.265 ;
      RECT 130.355 -27.248 130.445 -26.24 ;
      RECT 130.305 -26.645 130.445 -26.475 ;
      RECT 130.355 -25.44 130.445 -24.432 ;
      RECT 130.305 -25.205 130.445 -25.035 ;
      RECT 130.355 -24.018 130.445 -23.01 ;
      RECT 130.305 -23.415 130.445 -23.245 ;
      RECT 130.355 -22.21 130.445 -21.202 ;
      RECT 130.305 -21.975 130.445 -21.805 ;
      RECT 130.355 -20.788 130.445 -19.78 ;
      RECT 130.305 -20.185 130.445 -20.015 ;
      RECT 130.355 -18.98 130.445 -17.972 ;
      RECT 130.305 -18.745 130.445 -18.575 ;
      RECT 130.355 -17.558 130.445 -16.55 ;
      RECT 130.305 -16.955 130.445 -16.785 ;
      RECT 130.355 -15.75 130.445 -14.742 ;
      RECT 130.305 -15.515 130.445 -15.345 ;
      RECT 130.355 -14.328 130.445 -13.32 ;
      RECT 130.305 -13.725 130.445 -13.555 ;
      RECT 130.355 -12.52 130.445 -11.512 ;
      RECT 130.305 -12.285 130.445 -12.115 ;
      RECT 130.355 -11.098 130.445 -10.09 ;
      RECT 130.305 -10.495 130.445 -10.325 ;
      RECT 130.355 -9.29 130.445 -8.282 ;
      RECT 130.305 -9.055 130.445 -8.885 ;
      RECT 130.355 -7.868 130.445 -6.86 ;
      RECT 130.305 -7.265 130.445 -7.095 ;
      RECT 130.355 -6.06 130.445 -5.052 ;
      RECT 130.305 -5.825 130.445 -5.655 ;
      RECT 130.355 -4.638 130.445 -3.63 ;
      RECT 130.305 -4.035 130.445 -3.865 ;
      RECT 130.355 -2.83 130.445 -1.822 ;
      RECT 130.305 -2.595 130.445 -2.425 ;
      RECT 130.355 -1.408 130.445 -0.4 ;
      RECT 130.305 -0.805 130.445 -0.635 ;
      RECT 130.355 0.4 130.445 1.408 ;
      RECT 130.305 0.635 130.445 0.805 ;
      RECT 129.955 -101.538 130.045 -100.531 ;
      RECT 129.955 -101.225 130.095 -101.055 ;
      RECT 129.955 -99.729 130.045 -98.722 ;
      RECT 129.955 -99.205 130.095 -99.035 ;
      RECT 129.955 -98.308 130.045 -97.301 ;
      RECT 129.955 -97.995 130.095 -97.825 ;
      RECT 129.955 -96.499 130.045 -95.492 ;
      RECT 129.955 -95.975 130.095 -95.805 ;
      RECT 129.955 -95.078 130.045 -94.071 ;
      RECT 129.955 -94.765 130.095 -94.595 ;
      RECT 129.955 -93.269 130.045 -92.262 ;
      RECT 129.955 -92.745 130.095 -92.575 ;
      RECT 129.955 -91.848 130.045 -90.841 ;
      RECT 129.955 -91.535 130.095 -91.365 ;
      RECT 129.955 -90.039 130.045 -89.032 ;
      RECT 129.955 -89.515 130.095 -89.345 ;
      RECT 129.955 -88.618 130.045 -87.611 ;
      RECT 129.955 -88.305 130.095 -88.135 ;
      RECT 129.955 -86.809 130.045 -85.802 ;
      RECT 129.955 -86.285 130.095 -86.115 ;
      RECT 129.955 -85.388 130.045 -84.381 ;
      RECT 129.955 -85.075 130.095 -84.905 ;
      RECT 129.955 -83.579 130.045 -82.572 ;
      RECT 129.955 -83.055 130.095 -82.885 ;
      RECT 129.955 -82.158 130.045 -81.151 ;
      RECT 129.955 -81.845 130.095 -81.675 ;
      RECT 129.955 -80.349 130.045 -79.342 ;
      RECT 129.955 -79.825 130.095 -79.655 ;
      RECT 129.955 -78.928 130.045 -77.921 ;
      RECT 129.955 -78.615 130.095 -78.445 ;
      RECT 129.955 -77.119 130.045 -76.112 ;
      RECT 129.955 -76.595 130.095 -76.425 ;
      RECT 129.955 -75.698 130.045 -74.691 ;
      RECT 129.955 -75.385 130.095 -75.215 ;
      RECT 129.955 -73.889 130.045 -72.882 ;
      RECT 129.955 -73.365 130.095 -73.195 ;
      RECT 129.955 -72.468 130.045 -71.461 ;
      RECT 129.955 -72.155 130.095 -71.985 ;
      RECT 129.955 -70.659 130.045 -69.652 ;
      RECT 129.955 -70.135 130.095 -69.965 ;
      RECT 129.955 -69.238 130.045 -68.231 ;
      RECT 129.955 -68.925 130.095 -68.755 ;
      RECT 129.955 -67.429 130.045 -66.422 ;
      RECT 129.955 -66.905 130.095 -66.735 ;
      RECT 129.955 -66.008 130.045 -65.001 ;
      RECT 129.955 -65.695 130.095 -65.525 ;
      RECT 129.955 -64.199 130.045 -63.192 ;
      RECT 129.955 -63.675 130.095 -63.505 ;
      RECT 129.955 -62.778 130.045 -61.771 ;
      RECT 129.955 -62.465 130.095 -62.295 ;
      RECT 129.955 -60.969 130.045 -59.962 ;
      RECT 129.955 -60.445 130.095 -60.275 ;
      RECT 129.955 -59.548 130.045 -58.541 ;
      RECT 129.955 -59.235 130.095 -59.065 ;
      RECT 129.955 -57.739 130.045 -56.732 ;
      RECT 129.955 -57.215 130.095 -57.045 ;
      RECT 129.955 -56.318 130.045 -55.311 ;
      RECT 129.955 -56.005 130.095 -55.835 ;
      RECT 129.955 -54.509 130.045 -53.502 ;
      RECT 129.955 -53.985 130.095 -53.815 ;
      RECT 129.955 -53.088 130.045 -52.081 ;
      RECT 129.955 -52.775 130.095 -52.605 ;
      RECT 129.955 -51.279 130.045 -50.272 ;
      RECT 129.955 -50.755 130.095 -50.585 ;
      RECT 129.955 -49.858 130.045 -48.851 ;
      RECT 129.955 -49.545 130.095 -49.375 ;
      RECT 129.955 -48.049 130.045 -47.042 ;
      RECT 129.955 -47.525 130.095 -47.355 ;
      RECT 129.955 -46.628 130.045 -45.621 ;
      RECT 129.955 -46.315 130.095 -46.145 ;
      RECT 129.955 -44.819 130.045 -43.812 ;
      RECT 129.955 -44.295 130.095 -44.125 ;
      RECT 129.955 -43.398 130.045 -42.391 ;
      RECT 129.955 -43.085 130.095 -42.915 ;
      RECT 129.955 -41.589 130.045 -40.582 ;
      RECT 129.955 -41.065 130.095 -40.895 ;
      RECT 129.955 -40.168 130.045 -39.161 ;
      RECT 129.955 -39.855 130.095 -39.685 ;
      RECT 129.955 -38.359 130.045 -37.352 ;
      RECT 129.955 -37.835 130.095 -37.665 ;
      RECT 129.955 -36.938 130.045 -35.931 ;
      RECT 129.955 -36.625 130.095 -36.455 ;
      RECT 129.955 -35.129 130.045 -34.122 ;
      RECT 129.955 -34.605 130.095 -34.435 ;
      RECT 129.955 -33.708 130.045 -32.701 ;
      RECT 129.955 -33.395 130.095 -33.225 ;
      RECT 129.955 -31.899 130.045 -30.892 ;
      RECT 129.955 -31.375 130.095 -31.205 ;
      RECT 129.955 -30.478 130.045 -29.471 ;
      RECT 129.955 -30.165 130.095 -29.995 ;
      RECT 129.955 -28.669 130.045 -27.662 ;
      RECT 129.955 -28.145 130.095 -27.975 ;
      RECT 129.955 -27.248 130.045 -26.241 ;
      RECT 129.955 -26.935 130.095 -26.765 ;
      RECT 129.955 -25.439 130.045 -24.432 ;
      RECT 129.955 -24.915 130.095 -24.745 ;
      RECT 129.955 -24.018 130.045 -23.011 ;
      RECT 129.955 -23.705 130.095 -23.535 ;
      RECT 129.955 -22.209 130.045 -21.202 ;
      RECT 129.955 -21.685 130.095 -21.515 ;
      RECT 129.955 -20.788 130.045 -19.781 ;
      RECT 129.955 -20.475 130.095 -20.305 ;
      RECT 129.955 -18.979 130.045 -17.972 ;
      RECT 129.955 -18.455 130.095 -18.285 ;
      RECT 129.955 -17.558 130.045 -16.551 ;
      RECT 129.955 -17.245 130.095 -17.075 ;
      RECT 129.955 -15.749 130.045 -14.742 ;
      RECT 129.955 -15.225 130.095 -15.055 ;
      RECT 129.955 -14.328 130.045 -13.321 ;
      RECT 129.955 -14.015 130.095 -13.845 ;
      RECT 129.955 -12.519 130.045 -11.512 ;
      RECT 129.955 -11.995 130.095 -11.825 ;
      RECT 129.955 -11.098 130.045 -10.091 ;
      RECT 129.955 -10.785 130.095 -10.615 ;
      RECT 129.955 -9.289 130.045 -8.282 ;
      RECT 129.955 -8.765 130.095 -8.595 ;
      RECT 129.955 -7.868 130.045 -6.861 ;
      RECT 129.955 -7.555 130.095 -7.385 ;
      RECT 129.955 -6.059 130.045 -5.052 ;
      RECT 129.955 -5.535 130.095 -5.365 ;
      RECT 129.955 -4.638 130.045 -3.631 ;
      RECT 129.955 -4.325 130.095 -4.155 ;
      RECT 129.955 -2.829 130.045 -1.822 ;
      RECT 129.955 -2.305 130.095 -2.135 ;
      RECT 129.955 -1.408 130.045 -0.401 ;
      RECT 129.955 -1.095 130.095 -0.925 ;
      RECT 129.955 0.401 130.045 1.408 ;
      RECT 129.955 0.925 130.095 1.095 ;
      RECT 125.785 -108.935 129.565 -108.815 ;
      RECT 127.105 -109.475 127.205 -108.815 ;
      RECT 126.545 -109.475 126.645 -108.815 ;
      RECT 125.985 -109.475 126.085 -108.815 ;
      RECT 129.155 -101.538 129.245 -100.53 ;
      RECT 129.105 -100.935 129.245 -100.765 ;
      RECT 129.155 -99.73 129.245 -98.722 ;
      RECT 129.105 -99.495 129.245 -99.325 ;
      RECT 129.155 -98.308 129.245 -97.3 ;
      RECT 129.105 -97.705 129.245 -97.535 ;
      RECT 129.155 -96.5 129.245 -95.492 ;
      RECT 129.105 -96.265 129.245 -96.095 ;
      RECT 129.155 -95.078 129.245 -94.07 ;
      RECT 129.105 -94.475 129.245 -94.305 ;
      RECT 129.155 -93.27 129.245 -92.262 ;
      RECT 129.105 -93.035 129.245 -92.865 ;
      RECT 129.155 -91.848 129.245 -90.84 ;
      RECT 129.105 -91.245 129.245 -91.075 ;
      RECT 129.155 -90.04 129.245 -89.032 ;
      RECT 129.105 -89.805 129.245 -89.635 ;
      RECT 129.155 -88.618 129.245 -87.61 ;
      RECT 129.105 -88.015 129.245 -87.845 ;
      RECT 129.155 -86.81 129.245 -85.802 ;
      RECT 129.105 -86.575 129.245 -86.405 ;
      RECT 129.155 -85.388 129.245 -84.38 ;
      RECT 129.105 -84.785 129.245 -84.615 ;
      RECT 129.155 -83.58 129.245 -82.572 ;
      RECT 129.105 -83.345 129.245 -83.175 ;
      RECT 129.155 -82.158 129.245 -81.15 ;
      RECT 129.105 -81.555 129.245 -81.385 ;
      RECT 129.155 -80.35 129.245 -79.342 ;
      RECT 129.105 -80.115 129.245 -79.945 ;
      RECT 129.155 -78.928 129.245 -77.92 ;
      RECT 129.105 -78.325 129.245 -78.155 ;
      RECT 129.155 -77.12 129.245 -76.112 ;
      RECT 129.105 -76.885 129.245 -76.715 ;
      RECT 129.155 -75.698 129.245 -74.69 ;
      RECT 129.105 -75.095 129.245 -74.925 ;
      RECT 129.155 -73.89 129.245 -72.882 ;
      RECT 129.105 -73.655 129.245 -73.485 ;
      RECT 129.155 -72.468 129.245 -71.46 ;
      RECT 129.105 -71.865 129.245 -71.695 ;
      RECT 129.155 -70.66 129.245 -69.652 ;
      RECT 129.105 -70.425 129.245 -70.255 ;
      RECT 129.155 -69.238 129.245 -68.23 ;
      RECT 129.105 -68.635 129.245 -68.465 ;
      RECT 129.155 -67.43 129.245 -66.422 ;
      RECT 129.105 -67.195 129.245 -67.025 ;
      RECT 129.155 -66.008 129.245 -65 ;
      RECT 129.105 -65.405 129.245 -65.235 ;
      RECT 129.155 -64.2 129.245 -63.192 ;
      RECT 129.105 -63.965 129.245 -63.795 ;
      RECT 129.155 -62.778 129.245 -61.77 ;
      RECT 129.105 -62.175 129.245 -62.005 ;
      RECT 129.155 -60.97 129.245 -59.962 ;
      RECT 129.105 -60.735 129.245 -60.565 ;
      RECT 129.155 -59.548 129.245 -58.54 ;
      RECT 129.105 -58.945 129.245 -58.775 ;
      RECT 129.155 -57.74 129.245 -56.732 ;
      RECT 129.105 -57.505 129.245 -57.335 ;
      RECT 129.155 -56.318 129.245 -55.31 ;
      RECT 129.105 -55.715 129.245 -55.545 ;
      RECT 129.155 -54.51 129.245 -53.502 ;
      RECT 129.105 -54.275 129.245 -54.105 ;
      RECT 129.155 -53.088 129.245 -52.08 ;
      RECT 129.105 -52.485 129.245 -52.315 ;
      RECT 129.155 -51.28 129.245 -50.272 ;
      RECT 129.105 -51.045 129.245 -50.875 ;
      RECT 129.155 -49.858 129.245 -48.85 ;
      RECT 129.105 -49.255 129.245 -49.085 ;
      RECT 129.155 -48.05 129.245 -47.042 ;
      RECT 129.105 -47.815 129.245 -47.645 ;
      RECT 129.155 -46.628 129.245 -45.62 ;
      RECT 129.105 -46.025 129.245 -45.855 ;
      RECT 129.155 -44.82 129.245 -43.812 ;
      RECT 129.105 -44.585 129.245 -44.415 ;
      RECT 129.155 -43.398 129.245 -42.39 ;
      RECT 129.105 -42.795 129.245 -42.625 ;
      RECT 129.155 -41.59 129.245 -40.582 ;
      RECT 129.105 -41.355 129.245 -41.185 ;
      RECT 129.155 -40.168 129.245 -39.16 ;
      RECT 129.105 -39.565 129.245 -39.395 ;
      RECT 129.155 -38.36 129.245 -37.352 ;
      RECT 129.105 -38.125 129.245 -37.955 ;
      RECT 129.155 -36.938 129.245 -35.93 ;
      RECT 129.105 -36.335 129.245 -36.165 ;
      RECT 129.155 -35.13 129.245 -34.122 ;
      RECT 129.105 -34.895 129.245 -34.725 ;
      RECT 129.155 -33.708 129.245 -32.7 ;
      RECT 129.105 -33.105 129.245 -32.935 ;
      RECT 129.155 -31.9 129.245 -30.892 ;
      RECT 129.105 -31.665 129.245 -31.495 ;
      RECT 129.155 -30.478 129.245 -29.47 ;
      RECT 129.105 -29.875 129.245 -29.705 ;
      RECT 129.155 -28.67 129.245 -27.662 ;
      RECT 129.105 -28.435 129.245 -28.265 ;
      RECT 129.155 -27.248 129.245 -26.24 ;
      RECT 129.105 -26.645 129.245 -26.475 ;
      RECT 129.155 -25.44 129.245 -24.432 ;
      RECT 129.105 -25.205 129.245 -25.035 ;
      RECT 129.155 -24.018 129.245 -23.01 ;
      RECT 129.105 -23.415 129.245 -23.245 ;
      RECT 129.155 -22.21 129.245 -21.202 ;
      RECT 129.105 -21.975 129.245 -21.805 ;
      RECT 129.155 -20.788 129.245 -19.78 ;
      RECT 129.105 -20.185 129.245 -20.015 ;
      RECT 129.155 -18.98 129.245 -17.972 ;
      RECT 129.105 -18.745 129.245 -18.575 ;
      RECT 129.155 -17.558 129.245 -16.55 ;
      RECT 129.105 -16.955 129.245 -16.785 ;
      RECT 129.155 -15.75 129.245 -14.742 ;
      RECT 129.105 -15.515 129.245 -15.345 ;
      RECT 129.155 -14.328 129.245 -13.32 ;
      RECT 129.105 -13.725 129.245 -13.555 ;
      RECT 129.155 -12.52 129.245 -11.512 ;
      RECT 129.105 -12.285 129.245 -12.115 ;
      RECT 129.155 -11.098 129.245 -10.09 ;
      RECT 129.105 -10.495 129.245 -10.325 ;
      RECT 129.155 -9.29 129.245 -8.282 ;
      RECT 129.105 -9.055 129.245 -8.885 ;
      RECT 129.155 -7.868 129.245 -6.86 ;
      RECT 129.105 -7.265 129.245 -7.095 ;
      RECT 129.155 -6.06 129.245 -5.052 ;
      RECT 129.105 -5.825 129.245 -5.655 ;
      RECT 129.155 -4.638 129.245 -3.63 ;
      RECT 129.105 -4.035 129.245 -3.865 ;
      RECT 129.155 -2.83 129.245 -1.822 ;
      RECT 129.105 -2.595 129.245 -2.425 ;
      RECT 129.155 -1.408 129.245 -0.4 ;
      RECT 129.105 -0.805 129.245 -0.635 ;
      RECT 129.155 0.4 129.245 1.408 ;
      RECT 129.105 0.635 129.245 0.805 ;
      RECT 127.725 -111.685 129.205 -111.585 ;
      RECT 127.725 -112.195 127.825 -111.585 ;
      RECT 127.945 -109.15 129.205 -109.05 ;
      RECT 129.105 -109.475 129.205 -109.05 ;
      RECT 128.545 -109.475 128.645 -109.05 ;
      RECT 127.985 -109.475 128.085 -109.05 ;
      RECT 128.755 -101.538 128.845 -100.531 ;
      RECT 128.755 -101.225 128.895 -101.055 ;
      RECT 128.755 -99.729 128.845 -98.722 ;
      RECT 128.755 -99.205 128.895 -99.035 ;
      RECT 128.755 -98.308 128.845 -97.301 ;
      RECT 128.755 -97.995 128.895 -97.825 ;
      RECT 128.755 -96.499 128.845 -95.492 ;
      RECT 128.755 -95.975 128.895 -95.805 ;
      RECT 128.755 -95.078 128.845 -94.071 ;
      RECT 128.755 -94.765 128.895 -94.595 ;
      RECT 128.755 -93.269 128.845 -92.262 ;
      RECT 128.755 -92.745 128.895 -92.575 ;
      RECT 128.755 -91.848 128.845 -90.841 ;
      RECT 128.755 -91.535 128.895 -91.365 ;
      RECT 128.755 -90.039 128.845 -89.032 ;
      RECT 128.755 -89.515 128.895 -89.345 ;
      RECT 128.755 -88.618 128.845 -87.611 ;
      RECT 128.755 -88.305 128.895 -88.135 ;
      RECT 128.755 -86.809 128.845 -85.802 ;
      RECT 128.755 -86.285 128.895 -86.115 ;
      RECT 128.755 -85.388 128.845 -84.381 ;
      RECT 128.755 -85.075 128.895 -84.905 ;
      RECT 128.755 -83.579 128.845 -82.572 ;
      RECT 128.755 -83.055 128.895 -82.885 ;
      RECT 128.755 -82.158 128.845 -81.151 ;
      RECT 128.755 -81.845 128.895 -81.675 ;
      RECT 128.755 -80.349 128.845 -79.342 ;
      RECT 128.755 -79.825 128.895 -79.655 ;
      RECT 128.755 -78.928 128.845 -77.921 ;
      RECT 128.755 -78.615 128.895 -78.445 ;
      RECT 128.755 -77.119 128.845 -76.112 ;
      RECT 128.755 -76.595 128.895 -76.425 ;
      RECT 128.755 -75.698 128.845 -74.691 ;
      RECT 128.755 -75.385 128.895 -75.215 ;
      RECT 128.755 -73.889 128.845 -72.882 ;
      RECT 128.755 -73.365 128.895 -73.195 ;
      RECT 128.755 -72.468 128.845 -71.461 ;
      RECT 128.755 -72.155 128.895 -71.985 ;
      RECT 128.755 -70.659 128.845 -69.652 ;
      RECT 128.755 -70.135 128.895 -69.965 ;
      RECT 128.755 -69.238 128.845 -68.231 ;
      RECT 128.755 -68.925 128.895 -68.755 ;
      RECT 128.755 -67.429 128.845 -66.422 ;
      RECT 128.755 -66.905 128.895 -66.735 ;
      RECT 128.755 -66.008 128.845 -65.001 ;
      RECT 128.755 -65.695 128.895 -65.525 ;
      RECT 128.755 -64.199 128.845 -63.192 ;
      RECT 128.755 -63.675 128.895 -63.505 ;
      RECT 128.755 -62.778 128.845 -61.771 ;
      RECT 128.755 -62.465 128.895 -62.295 ;
      RECT 128.755 -60.969 128.845 -59.962 ;
      RECT 128.755 -60.445 128.895 -60.275 ;
      RECT 128.755 -59.548 128.845 -58.541 ;
      RECT 128.755 -59.235 128.895 -59.065 ;
      RECT 128.755 -57.739 128.845 -56.732 ;
      RECT 128.755 -57.215 128.895 -57.045 ;
      RECT 128.755 -56.318 128.845 -55.311 ;
      RECT 128.755 -56.005 128.895 -55.835 ;
      RECT 128.755 -54.509 128.845 -53.502 ;
      RECT 128.755 -53.985 128.895 -53.815 ;
      RECT 128.755 -53.088 128.845 -52.081 ;
      RECT 128.755 -52.775 128.895 -52.605 ;
      RECT 128.755 -51.279 128.845 -50.272 ;
      RECT 128.755 -50.755 128.895 -50.585 ;
      RECT 128.755 -49.858 128.845 -48.851 ;
      RECT 128.755 -49.545 128.895 -49.375 ;
      RECT 128.755 -48.049 128.845 -47.042 ;
      RECT 128.755 -47.525 128.895 -47.355 ;
      RECT 128.755 -46.628 128.845 -45.621 ;
      RECT 128.755 -46.315 128.895 -46.145 ;
      RECT 128.755 -44.819 128.845 -43.812 ;
      RECT 128.755 -44.295 128.895 -44.125 ;
      RECT 128.755 -43.398 128.845 -42.391 ;
      RECT 128.755 -43.085 128.895 -42.915 ;
      RECT 128.755 -41.589 128.845 -40.582 ;
      RECT 128.755 -41.065 128.895 -40.895 ;
      RECT 128.755 -40.168 128.845 -39.161 ;
      RECT 128.755 -39.855 128.895 -39.685 ;
      RECT 128.755 -38.359 128.845 -37.352 ;
      RECT 128.755 -37.835 128.895 -37.665 ;
      RECT 128.755 -36.938 128.845 -35.931 ;
      RECT 128.755 -36.625 128.895 -36.455 ;
      RECT 128.755 -35.129 128.845 -34.122 ;
      RECT 128.755 -34.605 128.895 -34.435 ;
      RECT 128.755 -33.708 128.845 -32.701 ;
      RECT 128.755 -33.395 128.895 -33.225 ;
      RECT 128.755 -31.899 128.845 -30.892 ;
      RECT 128.755 -31.375 128.895 -31.205 ;
      RECT 128.755 -30.478 128.845 -29.471 ;
      RECT 128.755 -30.165 128.895 -29.995 ;
      RECT 128.755 -28.669 128.845 -27.662 ;
      RECT 128.755 -28.145 128.895 -27.975 ;
      RECT 128.755 -27.248 128.845 -26.241 ;
      RECT 128.755 -26.935 128.895 -26.765 ;
      RECT 128.755 -25.439 128.845 -24.432 ;
      RECT 128.755 -24.915 128.895 -24.745 ;
      RECT 128.755 -24.018 128.845 -23.011 ;
      RECT 128.755 -23.705 128.895 -23.535 ;
      RECT 128.755 -22.209 128.845 -21.202 ;
      RECT 128.755 -21.685 128.895 -21.515 ;
      RECT 128.755 -20.788 128.845 -19.781 ;
      RECT 128.755 -20.475 128.895 -20.305 ;
      RECT 128.755 -18.979 128.845 -17.972 ;
      RECT 128.755 -18.455 128.895 -18.285 ;
      RECT 128.755 -17.558 128.845 -16.551 ;
      RECT 128.755 -17.245 128.895 -17.075 ;
      RECT 128.755 -15.749 128.845 -14.742 ;
      RECT 128.755 -15.225 128.895 -15.055 ;
      RECT 128.755 -14.328 128.845 -13.321 ;
      RECT 128.755 -14.015 128.895 -13.845 ;
      RECT 128.755 -12.519 128.845 -11.512 ;
      RECT 128.755 -11.995 128.895 -11.825 ;
      RECT 128.755 -11.098 128.845 -10.091 ;
      RECT 128.755 -10.785 128.895 -10.615 ;
      RECT 128.755 -9.289 128.845 -8.282 ;
      RECT 128.755 -8.765 128.895 -8.595 ;
      RECT 128.755 -7.868 128.845 -6.861 ;
      RECT 128.755 -7.555 128.895 -7.385 ;
      RECT 128.755 -6.059 128.845 -5.052 ;
      RECT 128.755 -5.535 128.895 -5.365 ;
      RECT 128.755 -4.638 128.845 -3.631 ;
      RECT 128.755 -4.325 128.895 -4.155 ;
      RECT 128.755 -2.829 128.845 -1.822 ;
      RECT 128.755 -2.305 128.895 -2.135 ;
      RECT 128.755 -1.408 128.845 -0.401 ;
      RECT 128.755 -1.095 128.895 -0.925 ;
      RECT 128.755 0.401 128.845 1.408 ;
      RECT 128.755 0.925 128.895 1.095 ;
      RECT 128.085 -111.495 128.255 -111.385 ;
      RECT 124.935 -111.495 128.255 -111.395 ;
      RECT 127.955 -101.538 128.045 -100.53 ;
      RECT 127.905 -100.935 128.045 -100.765 ;
      RECT 127.955 -99.73 128.045 -98.722 ;
      RECT 127.905 -99.495 128.045 -99.325 ;
      RECT 127.955 -98.308 128.045 -97.3 ;
      RECT 127.905 -97.705 128.045 -97.535 ;
      RECT 127.955 -96.5 128.045 -95.492 ;
      RECT 127.905 -96.265 128.045 -96.095 ;
      RECT 127.955 -95.078 128.045 -94.07 ;
      RECT 127.905 -94.475 128.045 -94.305 ;
      RECT 127.955 -93.27 128.045 -92.262 ;
      RECT 127.905 -93.035 128.045 -92.865 ;
      RECT 127.955 -91.848 128.045 -90.84 ;
      RECT 127.905 -91.245 128.045 -91.075 ;
      RECT 127.955 -90.04 128.045 -89.032 ;
      RECT 127.905 -89.805 128.045 -89.635 ;
      RECT 127.955 -88.618 128.045 -87.61 ;
      RECT 127.905 -88.015 128.045 -87.845 ;
      RECT 127.955 -86.81 128.045 -85.802 ;
      RECT 127.905 -86.575 128.045 -86.405 ;
      RECT 127.955 -85.388 128.045 -84.38 ;
      RECT 127.905 -84.785 128.045 -84.615 ;
      RECT 127.955 -83.58 128.045 -82.572 ;
      RECT 127.905 -83.345 128.045 -83.175 ;
      RECT 127.955 -82.158 128.045 -81.15 ;
      RECT 127.905 -81.555 128.045 -81.385 ;
      RECT 127.955 -80.35 128.045 -79.342 ;
      RECT 127.905 -80.115 128.045 -79.945 ;
      RECT 127.955 -78.928 128.045 -77.92 ;
      RECT 127.905 -78.325 128.045 -78.155 ;
      RECT 127.955 -77.12 128.045 -76.112 ;
      RECT 127.905 -76.885 128.045 -76.715 ;
      RECT 127.955 -75.698 128.045 -74.69 ;
      RECT 127.905 -75.095 128.045 -74.925 ;
      RECT 127.955 -73.89 128.045 -72.882 ;
      RECT 127.905 -73.655 128.045 -73.485 ;
      RECT 127.955 -72.468 128.045 -71.46 ;
      RECT 127.905 -71.865 128.045 -71.695 ;
      RECT 127.955 -70.66 128.045 -69.652 ;
      RECT 127.905 -70.425 128.045 -70.255 ;
      RECT 127.955 -69.238 128.045 -68.23 ;
      RECT 127.905 -68.635 128.045 -68.465 ;
      RECT 127.955 -67.43 128.045 -66.422 ;
      RECT 127.905 -67.195 128.045 -67.025 ;
      RECT 127.955 -66.008 128.045 -65 ;
      RECT 127.905 -65.405 128.045 -65.235 ;
      RECT 127.955 -64.2 128.045 -63.192 ;
      RECT 127.905 -63.965 128.045 -63.795 ;
      RECT 127.955 -62.778 128.045 -61.77 ;
      RECT 127.905 -62.175 128.045 -62.005 ;
      RECT 127.955 -60.97 128.045 -59.962 ;
      RECT 127.905 -60.735 128.045 -60.565 ;
      RECT 127.955 -59.548 128.045 -58.54 ;
      RECT 127.905 -58.945 128.045 -58.775 ;
      RECT 127.955 -57.74 128.045 -56.732 ;
      RECT 127.905 -57.505 128.045 -57.335 ;
      RECT 127.955 -56.318 128.045 -55.31 ;
      RECT 127.905 -55.715 128.045 -55.545 ;
      RECT 127.955 -54.51 128.045 -53.502 ;
      RECT 127.905 -54.275 128.045 -54.105 ;
      RECT 127.955 -53.088 128.045 -52.08 ;
      RECT 127.905 -52.485 128.045 -52.315 ;
      RECT 127.955 -51.28 128.045 -50.272 ;
      RECT 127.905 -51.045 128.045 -50.875 ;
      RECT 127.955 -49.858 128.045 -48.85 ;
      RECT 127.905 -49.255 128.045 -49.085 ;
      RECT 127.955 -48.05 128.045 -47.042 ;
      RECT 127.905 -47.815 128.045 -47.645 ;
      RECT 127.955 -46.628 128.045 -45.62 ;
      RECT 127.905 -46.025 128.045 -45.855 ;
      RECT 127.955 -44.82 128.045 -43.812 ;
      RECT 127.905 -44.585 128.045 -44.415 ;
      RECT 127.955 -43.398 128.045 -42.39 ;
      RECT 127.905 -42.795 128.045 -42.625 ;
      RECT 127.955 -41.59 128.045 -40.582 ;
      RECT 127.905 -41.355 128.045 -41.185 ;
      RECT 127.955 -40.168 128.045 -39.16 ;
      RECT 127.905 -39.565 128.045 -39.395 ;
      RECT 127.955 -38.36 128.045 -37.352 ;
      RECT 127.905 -38.125 128.045 -37.955 ;
      RECT 127.955 -36.938 128.045 -35.93 ;
      RECT 127.905 -36.335 128.045 -36.165 ;
      RECT 127.955 -35.13 128.045 -34.122 ;
      RECT 127.905 -34.895 128.045 -34.725 ;
      RECT 127.955 -33.708 128.045 -32.7 ;
      RECT 127.905 -33.105 128.045 -32.935 ;
      RECT 127.955 -31.9 128.045 -30.892 ;
      RECT 127.905 -31.665 128.045 -31.495 ;
      RECT 127.955 -30.478 128.045 -29.47 ;
      RECT 127.905 -29.875 128.045 -29.705 ;
      RECT 127.955 -28.67 128.045 -27.662 ;
      RECT 127.905 -28.435 128.045 -28.265 ;
      RECT 127.955 -27.248 128.045 -26.24 ;
      RECT 127.905 -26.645 128.045 -26.475 ;
      RECT 127.955 -25.44 128.045 -24.432 ;
      RECT 127.905 -25.205 128.045 -25.035 ;
      RECT 127.955 -24.018 128.045 -23.01 ;
      RECT 127.905 -23.415 128.045 -23.245 ;
      RECT 127.955 -22.21 128.045 -21.202 ;
      RECT 127.905 -21.975 128.045 -21.805 ;
      RECT 127.955 -20.788 128.045 -19.78 ;
      RECT 127.905 -20.185 128.045 -20.015 ;
      RECT 127.955 -18.98 128.045 -17.972 ;
      RECT 127.905 -18.745 128.045 -18.575 ;
      RECT 127.955 -17.558 128.045 -16.55 ;
      RECT 127.905 -16.955 128.045 -16.785 ;
      RECT 127.955 -15.75 128.045 -14.742 ;
      RECT 127.905 -15.515 128.045 -15.345 ;
      RECT 127.955 -14.328 128.045 -13.32 ;
      RECT 127.905 -13.725 128.045 -13.555 ;
      RECT 127.955 -12.52 128.045 -11.512 ;
      RECT 127.905 -12.285 128.045 -12.115 ;
      RECT 127.955 -11.098 128.045 -10.09 ;
      RECT 127.905 -10.495 128.045 -10.325 ;
      RECT 127.955 -9.29 128.045 -8.282 ;
      RECT 127.905 -9.055 128.045 -8.885 ;
      RECT 127.955 -7.868 128.045 -6.86 ;
      RECT 127.905 -7.265 128.045 -7.095 ;
      RECT 127.955 -6.06 128.045 -5.052 ;
      RECT 127.905 -5.825 128.045 -5.655 ;
      RECT 127.955 -4.638 128.045 -3.63 ;
      RECT 127.905 -4.035 128.045 -3.865 ;
      RECT 127.955 -2.83 128.045 -1.822 ;
      RECT 127.905 -2.595 128.045 -2.425 ;
      RECT 127.955 -1.408 128.045 -0.4 ;
      RECT 127.905 -0.805 128.045 -0.635 ;
      RECT 127.955 0.4 128.045 1.408 ;
      RECT 127.905 0.635 128.045 0.805 ;
      RECT 127.555 -101.538 127.645 -100.531 ;
      RECT 127.555 -101.225 127.695 -101.055 ;
      RECT 127.555 -99.729 127.645 -98.722 ;
      RECT 127.555 -99.205 127.695 -99.035 ;
      RECT 127.555 -98.308 127.645 -97.301 ;
      RECT 127.555 -97.995 127.695 -97.825 ;
      RECT 127.555 -96.499 127.645 -95.492 ;
      RECT 127.555 -95.975 127.695 -95.805 ;
      RECT 127.555 -95.078 127.645 -94.071 ;
      RECT 127.555 -94.765 127.695 -94.595 ;
      RECT 127.555 -93.269 127.645 -92.262 ;
      RECT 127.555 -92.745 127.695 -92.575 ;
      RECT 127.555 -91.848 127.645 -90.841 ;
      RECT 127.555 -91.535 127.695 -91.365 ;
      RECT 127.555 -90.039 127.645 -89.032 ;
      RECT 127.555 -89.515 127.695 -89.345 ;
      RECT 127.555 -88.618 127.645 -87.611 ;
      RECT 127.555 -88.305 127.695 -88.135 ;
      RECT 127.555 -86.809 127.645 -85.802 ;
      RECT 127.555 -86.285 127.695 -86.115 ;
      RECT 127.555 -85.388 127.645 -84.381 ;
      RECT 127.555 -85.075 127.695 -84.905 ;
      RECT 127.555 -83.579 127.645 -82.572 ;
      RECT 127.555 -83.055 127.695 -82.885 ;
      RECT 127.555 -82.158 127.645 -81.151 ;
      RECT 127.555 -81.845 127.695 -81.675 ;
      RECT 127.555 -80.349 127.645 -79.342 ;
      RECT 127.555 -79.825 127.695 -79.655 ;
      RECT 127.555 -78.928 127.645 -77.921 ;
      RECT 127.555 -78.615 127.695 -78.445 ;
      RECT 127.555 -77.119 127.645 -76.112 ;
      RECT 127.555 -76.595 127.695 -76.425 ;
      RECT 127.555 -75.698 127.645 -74.691 ;
      RECT 127.555 -75.385 127.695 -75.215 ;
      RECT 127.555 -73.889 127.645 -72.882 ;
      RECT 127.555 -73.365 127.695 -73.195 ;
      RECT 127.555 -72.468 127.645 -71.461 ;
      RECT 127.555 -72.155 127.695 -71.985 ;
      RECT 127.555 -70.659 127.645 -69.652 ;
      RECT 127.555 -70.135 127.695 -69.965 ;
      RECT 127.555 -69.238 127.645 -68.231 ;
      RECT 127.555 -68.925 127.695 -68.755 ;
      RECT 127.555 -67.429 127.645 -66.422 ;
      RECT 127.555 -66.905 127.695 -66.735 ;
      RECT 127.555 -66.008 127.645 -65.001 ;
      RECT 127.555 -65.695 127.695 -65.525 ;
      RECT 127.555 -64.199 127.645 -63.192 ;
      RECT 127.555 -63.675 127.695 -63.505 ;
      RECT 127.555 -62.778 127.645 -61.771 ;
      RECT 127.555 -62.465 127.695 -62.295 ;
      RECT 127.555 -60.969 127.645 -59.962 ;
      RECT 127.555 -60.445 127.695 -60.275 ;
      RECT 127.555 -59.548 127.645 -58.541 ;
      RECT 127.555 -59.235 127.695 -59.065 ;
      RECT 127.555 -57.739 127.645 -56.732 ;
      RECT 127.555 -57.215 127.695 -57.045 ;
      RECT 127.555 -56.318 127.645 -55.311 ;
      RECT 127.555 -56.005 127.695 -55.835 ;
      RECT 127.555 -54.509 127.645 -53.502 ;
      RECT 127.555 -53.985 127.695 -53.815 ;
      RECT 127.555 -53.088 127.645 -52.081 ;
      RECT 127.555 -52.775 127.695 -52.605 ;
      RECT 127.555 -51.279 127.645 -50.272 ;
      RECT 127.555 -50.755 127.695 -50.585 ;
      RECT 127.555 -49.858 127.645 -48.851 ;
      RECT 127.555 -49.545 127.695 -49.375 ;
      RECT 127.555 -48.049 127.645 -47.042 ;
      RECT 127.555 -47.525 127.695 -47.355 ;
      RECT 127.555 -46.628 127.645 -45.621 ;
      RECT 127.555 -46.315 127.695 -46.145 ;
      RECT 127.555 -44.819 127.645 -43.812 ;
      RECT 127.555 -44.295 127.695 -44.125 ;
      RECT 127.555 -43.398 127.645 -42.391 ;
      RECT 127.555 -43.085 127.695 -42.915 ;
      RECT 127.555 -41.589 127.645 -40.582 ;
      RECT 127.555 -41.065 127.695 -40.895 ;
      RECT 127.555 -40.168 127.645 -39.161 ;
      RECT 127.555 -39.855 127.695 -39.685 ;
      RECT 127.555 -38.359 127.645 -37.352 ;
      RECT 127.555 -37.835 127.695 -37.665 ;
      RECT 127.555 -36.938 127.645 -35.931 ;
      RECT 127.555 -36.625 127.695 -36.455 ;
      RECT 127.555 -35.129 127.645 -34.122 ;
      RECT 127.555 -34.605 127.695 -34.435 ;
      RECT 127.555 -33.708 127.645 -32.701 ;
      RECT 127.555 -33.395 127.695 -33.225 ;
      RECT 127.555 -31.899 127.645 -30.892 ;
      RECT 127.555 -31.375 127.695 -31.205 ;
      RECT 127.555 -30.478 127.645 -29.471 ;
      RECT 127.555 -30.165 127.695 -29.995 ;
      RECT 127.555 -28.669 127.645 -27.662 ;
      RECT 127.555 -28.145 127.695 -27.975 ;
      RECT 127.555 -27.248 127.645 -26.241 ;
      RECT 127.555 -26.935 127.695 -26.765 ;
      RECT 127.555 -25.439 127.645 -24.432 ;
      RECT 127.555 -24.915 127.695 -24.745 ;
      RECT 127.555 -24.018 127.645 -23.011 ;
      RECT 127.555 -23.705 127.695 -23.535 ;
      RECT 127.555 -22.209 127.645 -21.202 ;
      RECT 127.555 -21.685 127.695 -21.515 ;
      RECT 127.555 -20.788 127.645 -19.781 ;
      RECT 127.555 -20.475 127.695 -20.305 ;
      RECT 127.555 -18.979 127.645 -17.972 ;
      RECT 127.555 -18.455 127.695 -18.285 ;
      RECT 127.555 -17.558 127.645 -16.551 ;
      RECT 127.555 -17.245 127.695 -17.075 ;
      RECT 127.555 -15.749 127.645 -14.742 ;
      RECT 127.555 -15.225 127.695 -15.055 ;
      RECT 127.555 -14.328 127.645 -13.321 ;
      RECT 127.555 -14.015 127.695 -13.845 ;
      RECT 127.555 -12.519 127.645 -11.512 ;
      RECT 127.555 -11.995 127.695 -11.825 ;
      RECT 127.555 -11.098 127.645 -10.091 ;
      RECT 127.555 -10.785 127.695 -10.615 ;
      RECT 127.555 -9.289 127.645 -8.282 ;
      RECT 127.555 -8.765 127.695 -8.595 ;
      RECT 127.555 -7.868 127.645 -6.861 ;
      RECT 127.555 -7.555 127.695 -7.385 ;
      RECT 127.555 -6.059 127.645 -5.052 ;
      RECT 127.555 -5.535 127.695 -5.365 ;
      RECT 127.555 -4.638 127.645 -3.631 ;
      RECT 127.555 -4.325 127.695 -4.155 ;
      RECT 127.555 -2.829 127.645 -1.822 ;
      RECT 127.555 -2.305 127.695 -2.135 ;
      RECT 127.555 -1.408 127.645 -0.401 ;
      RECT 127.555 -1.095 127.695 -0.925 ;
      RECT 127.555 0.401 127.645 1.408 ;
      RECT 127.555 0.925 127.695 1.095 ;
      RECT 125.705 -111.685 127.185 -111.585 ;
      RECT 125.705 -112.055 125.805 -111.585 ;
      RECT 125.51 -114.395 127.085 -114.275 ;
      RECT 126.985 -114.895 127.085 -114.275 ;
      RECT 126.39 -114.895 126.49 -114.275 ;
      RECT 125.51 -114.85 125.61 -114.275 ;
      RECT 126.755 -101.538 126.845 -100.53 ;
      RECT 126.705 -100.935 126.845 -100.765 ;
      RECT 126.755 -99.73 126.845 -98.722 ;
      RECT 126.705 -99.495 126.845 -99.325 ;
      RECT 126.755 -98.308 126.845 -97.3 ;
      RECT 126.705 -97.705 126.845 -97.535 ;
      RECT 126.755 -96.5 126.845 -95.492 ;
      RECT 126.705 -96.265 126.845 -96.095 ;
      RECT 126.755 -95.078 126.845 -94.07 ;
      RECT 126.705 -94.475 126.845 -94.305 ;
      RECT 126.755 -93.27 126.845 -92.262 ;
      RECT 126.705 -93.035 126.845 -92.865 ;
      RECT 126.755 -91.848 126.845 -90.84 ;
      RECT 126.705 -91.245 126.845 -91.075 ;
      RECT 126.755 -90.04 126.845 -89.032 ;
      RECT 126.705 -89.805 126.845 -89.635 ;
      RECT 126.755 -88.618 126.845 -87.61 ;
      RECT 126.705 -88.015 126.845 -87.845 ;
      RECT 126.755 -86.81 126.845 -85.802 ;
      RECT 126.705 -86.575 126.845 -86.405 ;
      RECT 126.755 -85.388 126.845 -84.38 ;
      RECT 126.705 -84.785 126.845 -84.615 ;
      RECT 126.755 -83.58 126.845 -82.572 ;
      RECT 126.705 -83.345 126.845 -83.175 ;
      RECT 126.755 -82.158 126.845 -81.15 ;
      RECT 126.705 -81.555 126.845 -81.385 ;
      RECT 126.755 -80.35 126.845 -79.342 ;
      RECT 126.705 -80.115 126.845 -79.945 ;
      RECT 126.755 -78.928 126.845 -77.92 ;
      RECT 126.705 -78.325 126.845 -78.155 ;
      RECT 126.755 -77.12 126.845 -76.112 ;
      RECT 126.705 -76.885 126.845 -76.715 ;
      RECT 126.755 -75.698 126.845 -74.69 ;
      RECT 126.705 -75.095 126.845 -74.925 ;
      RECT 126.755 -73.89 126.845 -72.882 ;
      RECT 126.705 -73.655 126.845 -73.485 ;
      RECT 126.755 -72.468 126.845 -71.46 ;
      RECT 126.705 -71.865 126.845 -71.695 ;
      RECT 126.755 -70.66 126.845 -69.652 ;
      RECT 126.705 -70.425 126.845 -70.255 ;
      RECT 126.755 -69.238 126.845 -68.23 ;
      RECT 126.705 -68.635 126.845 -68.465 ;
      RECT 126.755 -67.43 126.845 -66.422 ;
      RECT 126.705 -67.195 126.845 -67.025 ;
      RECT 126.755 -66.008 126.845 -65 ;
      RECT 126.705 -65.405 126.845 -65.235 ;
      RECT 126.755 -64.2 126.845 -63.192 ;
      RECT 126.705 -63.965 126.845 -63.795 ;
      RECT 126.755 -62.778 126.845 -61.77 ;
      RECT 126.705 -62.175 126.845 -62.005 ;
      RECT 126.755 -60.97 126.845 -59.962 ;
      RECT 126.705 -60.735 126.845 -60.565 ;
      RECT 126.755 -59.548 126.845 -58.54 ;
      RECT 126.705 -58.945 126.845 -58.775 ;
      RECT 126.755 -57.74 126.845 -56.732 ;
      RECT 126.705 -57.505 126.845 -57.335 ;
      RECT 126.755 -56.318 126.845 -55.31 ;
      RECT 126.705 -55.715 126.845 -55.545 ;
      RECT 126.755 -54.51 126.845 -53.502 ;
      RECT 126.705 -54.275 126.845 -54.105 ;
      RECT 126.755 -53.088 126.845 -52.08 ;
      RECT 126.705 -52.485 126.845 -52.315 ;
      RECT 126.755 -51.28 126.845 -50.272 ;
      RECT 126.705 -51.045 126.845 -50.875 ;
      RECT 126.755 -49.858 126.845 -48.85 ;
      RECT 126.705 -49.255 126.845 -49.085 ;
      RECT 126.755 -48.05 126.845 -47.042 ;
      RECT 126.705 -47.815 126.845 -47.645 ;
      RECT 126.755 -46.628 126.845 -45.62 ;
      RECT 126.705 -46.025 126.845 -45.855 ;
      RECT 126.755 -44.82 126.845 -43.812 ;
      RECT 126.705 -44.585 126.845 -44.415 ;
      RECT 126.755 -43.398 126.845 -42.39 ;
      RECT 126.705 -42.795 126.845 -42.625 ;
      RECT 126.755 -41.59 126.845 -40.582 ;
      RECT 126.705 -41.355 126.845 -41.185 ;
      RECT 126.755 -40.168 126.845 -39.16 ;
      RECT 126.705 -39.565 126.845 -39.395 ;
      RECT 126.755 -38.36 126.845 -37.352 ;
      RECT 126.705 -38.125 126.845 -37.955 ;
      RECT 126.755 -36.938 126.845 -35.93 ;
      RECT 126.705 -36.335 126.845 -36.165 ;
      RECT 126.755 -35.13 126.845 -34.122 ;
      RECT 126.705 -34.895 126.845 -34.725 ;
      RECT 126.755 -33.708 126.845 -32.7 ;
      RECT 126.705 -33.105 126.845 -32.935 ;
      RECT 126.755 -31.9 126.845 -30.892 ;
      RECT 126.705 -31.665 126.845 -31.495 ;
      RECT 126.755 -30.478 126.845 -29.47 ;
      RECT 126.705 -29.875 126.845 -29.705 ;
      RECT 126.755 -28.67 126.845 -27.662 ;
      RECT 126.705 -28.435 126.845 -28.265 ;
      RECT 126.755 -27.248 126.845 -26.24 ;
      RECT 126.705 -26.645 126.845 -26.475 ;
      RECT 126.755 -25.44 126.845 -24.432 ;
      RECT 126.705 -25.205 126.845 -25.035 ;
      RECT 126.755 -24.018 126.845 -23.01 ;
      RECT 126.705 -23.415 126.845 -23.245 ;
      RECT 126.755 -22.21 126.845 -21.202 ;
      RECT 126.705 -21.975 126.845 -21.805 ;
      RECT 126.755 -20.788 126.845 -19.78 ;
      RECT 126.705 -20.185 126.845 -20.015 ;
      RECT 126.755 -18.98 126.845 -17.972 ;
      RECT 126.705 -18.745 126.845 -18.575 ;
      RECT 126.755 -17.558 126.845 -16.55 ;
      RECT 126.705 -16.955 126.845 -16.785 ;
      RECT 126.755 -15.75 126.845 -14.742 ;
      RECT 126.705 -15.515 126.845 -15.345 ;
      RECT 126.755 -14.328 126.845 -13.32 ;
      RECT 126.705 -13.725 126.845 -13.555 ;
      RECT 126.755 -12.52 126.845 -11.512 ;
      RECT 126.705 -12.285 126.845 -12.115 ;
      RECT 126.755 -11.098 126.845 -10.09 ;
      RECT 126.705 -10.495 126.845 -10.325 ;
      RECT 126.755 -9.29 126.845 -8.282 ;
      RECT 126.705 -9.055 126.845 -8.885 ;
      RECT 126.755 -7.868 126.845 -6.86 ;
      RECT 126.705 -7.265 126.845 -7.095 ;
      RECT 126.755 -6.06 126.845 -5.052 ;
      RECT 126.705 -5.825 126.845 -5.655 ;
      RECT 126.755 -4.638 126.845 -3.63 ;
      RECT 126.705 -4.035 126.845 -3.865 ;
      RECT 126.755 -2.83 126.845 -1.822 ;
      RECT 126.705 -2.595 126.845 -2.425 ;
      RECT 126.755 -1.408 126.845 -0.4 ;
      RECT 126.705 -0.805 126.845 -0.635 ;
      RECT 126.755 0.4 126.845 1.408 ;
      RECT 126.705 0.635 126.845 0.805 ;
      RECT 126.63 -114.685 126.805 -114.515 ;
      RECT 126.705 -114.895 126.805 -114.515 ;
      RECT 125.745 -113.555 125.845 -113.09 ;
      RECT 126.11 -113.555 126.21 -113.1 ;
      RECT 125.745 -113.555 126.59 -113.385 ;
      RECT 126.355 -101.538 126.445 -100.531 ;
      RECT 126.355 -101.225 126.495 -101.055 ;
      RECT 126.355 -99.729 126.445 -98.722 ;
      RECT 126.355 -99.205 126.495 -99.035 ;
      RECT 126.355 -98.308 126.445 -97.301 ;
      RECT 126.355 -97.995 126.495 -97.825 ;
      RECT 126.355 -96.499 126.445 -95.492 ;
      RECT 126.355 -95.975 126.495 -95.805 ;
      RECT 126.355 -95.078 126.445 -94.071 ;
      RECT 126.355 -94.765 126.495 -94.595 ;
      RECT 126.355 -93.269 126.445 -92.262 ;
      RECT 126.355 -92.745 126.495 -92.575 ;
      RECT 126.355 -91.848 126.445 -90.841 ;
      RECT 126.355 -91.535 126.495 -91.365 ;
      RECT 126.355 -90.039 126.445 -89.032 ;
      RECT 126.355 -89.515 126.495 -89.345 ;
      RECT 126.355 -88.618 126.445 -87.611 ;
      RECT 126.355 -88.305 126.495 -88.135 ;
      RECT 126.355 -86.809 126.445 -85.802 ;
      RECT 126.355 -86.285 126.495 -86.115 ;
      RECT 126.355 -85.388 126.445 -84.381 ;
      RECT 126.355 -85.075 126.495 -84.905 ;
      RECT 126.355 -83.579 126.445 -82.572 ;
      RECT 126.355 -83.055 126.495 -82.885 ;
      RECT 126.355 -82.158 126.445 -81.151 ;
      RECT 126.355 -81.845 126.495 -81.675 ;
      RECT 126.355 -80.349 126.445 -79.342 ;
      RECT 126.355 -79.825 126.495 -79.655 ;
      RECT 126.355 -78.928 126.445 -77.921 ;
      RECT 126.355 -78.615 126.495 -78.445 ;
      RECT 126.355 -77.119 126.445 -76.112 ;
      RECT 126.355 -76.595 126.495 -76.425 ;
      RECT 126.355 -75.698 126.445 -74.691 ;
      RECT 126.355 -75.385 126.495 -75.215 ;
      RECT 126.355 -73.889 126.445 -72.882 ;
      RECT 126.355 -73.365 126.495 -73.195 ;
      RECT 126.355 -72.468 126.445 -71.461 ;
      RECT 126.355 -72.155 126.495 -71.985 ;
      RECT 126.355 -70.659 126.445 -69.652 ;
      RECT 126.355 -70.135 126.495 -69.965 ;
      RECT 126.355 -69.238 126.445 -68.231 ;
      RECT 126.355 -68.925 126.495 -68.755 ;
      RECT 126.355 -67.429 126.445 -66.422 ;
      RECT 126.355 -66.905 126.495 -66.735 ;
      RECT 126.355 -66.008 126.445 -65.001 ;
      RECT 126.355 -65.695 126.495 -65.525 ;
      RECT 126.355 -64.199 126.445 -63.192 ;
      RECT 126.355 -63.675 126.495 -63.505 ;
      RECT 126.355 -62.778 126.445 -61.771 ;
      RECT 126.355 -62.465 126.495 -62.295 ;
      RECT 126.355 -60.969 126.445 -59.962 ;
      RECT 126.355 -60.445 126.495 -60.275 ;
      RECT 126.355 -59.548 126.445 -58.541 ;
      RECT 126.355 -59.235 126.495 -59.065 ;
      RECT 126.355 -57.739 126.445 -56.732 ;
      RECT 126.355 -57.215 126.495 -57.045 ;
      RECT 126.355 -56.318 126.445 -55.311 ;
      RECT 126.355 -56.005 126.495 -55.835 ;
      RECT 126.355 -54.509 126.445 -53.502 ;
      RECT 126.355 -53.985 126.495 -53.815 ;
      RECT 126.355 -53.088 126.445 -52.081 ;
      RECT 126.355 -52.775 126.495 -52.605 ;
      RECT 126.355 -51.279 126.445 -50.272 ;
      RECT 126.355 -50.755 126.495 -50.585 ;
      RECT 126.355 -49.858 126.445 -48.851 ;
      RECT 126.355 -49.545 126.495 -49.375 ;
      RECT 126.355 -48.049 126.445 -47.042 ;
      RECT 126.355 -47.525 126.495 -47.355 ;
      RECT 126.355 -46.628 126.445 -45.621 ;
      RECT 126.355 -46.315 126.495 -46.145 ;
      RECT 126.355 -44.819 126.445 -43.812 ;
      RECT 126.355 -44.295 126.495 -44.125 ;
      RECT 126.355 -43.398 126.445 -42.391 ;
      RECT 126.355 -43.085 126.495 -42.915 ;
      RECT 126.355 -41.589 126.445 -40.582 ;
      RECT 126.355 -41.065 126.495 -40.895 ;
      RECT 126.355 -40.168 126.445 -39.161 ;
      RECT 126.355 -39.855 126.495 -39.685 ;
      RECT 126.355 -38.359 126.445 -37.352 ;
      RECT 126.355 -37.835 126.495 -37.665 ;
      RECT 126.355 -36.938 126.445 -35.931 ;
      RECT 126.355 -36.625 126.495 -36.455 ;
      RECT 126.355 -35.129 126.445 -34.122 ;
      RECT 126.355 -34.605 126.495 -34.435 ;
      RECT 126.355 -33.708 126.445 -32.701 ;
      RECT 126.355 -33.395 126.495 -33.225 ;
      RECT 126.355 -31.899 126.445 -30.892 ;
      RECT 126.355 -31.375 126.495 -31.205 ;
      RECT 126.355 -30.478 126.445 -29.471 ;
      RECT 126.355 -30.165 126.495 -29.995 ;
      RECT 126.355 -28.669 126.445 -27.662 ;
      RECT 126.355 -28.145 126.495 -27.975 ;
      RECT 126.355 -27.248 126.445 -26.241 ;
      RECT 126.355 -26.935 126.495 -26.765 ;
      RECT 126.355 -25.439 126.445 -24.432 ;
      RECT 126.355 -24.915 126.495 -24.745 ;
      RECT 126.355 -24.018 126.445 -23.011 ;
      RECT 126.355 -23.705 126.495 -23.535 ;
      RECT 126.355 -22.209 126.445 -21.202 ;
      RECT 126.355 -21.685 126.495 -21.515 ;
      RECT 126.355 -20.788 126.445 -19.781 ;
      RECT 126.355 -20.475 126.495 -20.305 ;
      RECT 126.355 -18.979 126.445 -17.972 ;
      RECT 126.355 -18.455 126.495 -18.285 ;
      RECT 126.355 -17.558 126.445 -16.551 ;
      RECT 126.355 -17.245 126.495 -17.075 ;
      RECT 126.355 -15.749 126.445 -14.742 ;
      RECT 126.355 -15.225 126.495 -15.055 ;
      RECT 126.355 -14.328 126.445 -13.321 ;
      RECT 126.355 -14.015 126.495 -13.845 ;
      RECT 126.355 -12.519 126.445 -11.512 ;
      RECT 126.355 -11.995 126.495 -11.825 ;
      RECT 126.355 -11.098 126.445 -10.091 ;
      RECT 126.355 -10.785 126.495 -10.615 ;
      RECT 126.355 -9.289 126.445 -8.282 ;
      RECT 126.355 -8.765 126.495 -8.595 ;
      RECT 126.355 -7.868 126.445 -6.861 ;
      RECT 126.355 -7.555 126.495 -7.385 ;
      RECT 126.355 -6.059 126.445 -5.052 ;
      RECT 126.355 -5.535 126.495 -5.365 ;
      RECT 126.355 -4.638 126.445 -3.631 ;
      RECT 126.355 -4.325 126.495 -4.155 ;
      RECT 126.355 -2.829 126.445 -1.822 ;
      RECT 126.355 -2.305 126.495 -2.135 ;
      RECT 126.355 -1.408 126.445 -0.401 ;
      RECT 126.355 -1.095 126.495 -0.925 ;
      RECT 126.355 0.401 126.445 1.408 ;
      RECT 126.355 0.925 126.495 1.095 ;
      RECT 126.04 -114.685 126.21 -114.515 ;
      RECT 126.11 -114.895 126.21 -114.515 ;
      RECT 125.555 -101.538 125.645 -100.53 ;
      RECT 125.505 -100.935 125.645 -100.765 ;
      RECT 125.555 -99.73 125.645 -98.722 ;
      RECT 125.505 -99.495 125.645 -99.325 ;
      RECT 125.555 -98.308 125.645 -97.3 ;
      RECT 125.505 -97.705 125.645 -97.535 ;
      RECT 125.555 -96.5 125.645 -95.492 ;
      RECT 125.505 -96.265 125.645 -96.095 ;
      RECT 125.555 -95.078 125.645 -94.07 ;
      RECT 125.505 -94.475 125.645 -94.305 ;
      RECT 125.555 -93.27 125.645 -92.262 ;
      RECT 125.505 -93.035 125.645 -92.865 ;
      RECT 125.555 -91.848 125.645 -90.84 ;
      RECT 125.505 -91.245 125.645 -91.075 ;
      RECT 125.555 -90.04 125.645 -89.032 ;
      RECT 125.505 -89.805 125.645 -89.635 ;
      RECT 125.555 -88.618 125.645 -87.61 ;
      RECT 125.505 -88.015 125.645 -87.845 ;
      RECT 125.555 -86.81 125.645 -85.802 ;
      RECT 125.505 -86.575 125.645 -86.405 ;
      RECT 125.555 -85.388 125.645 -84.38 ;
      RECT 125.505 -84.785 125.645 -84.615 ;
      RECT 125.555 -83.58 125.645 -82.572 ;
      RECT 125.505 -83.345 125.645 -83.175 ;
      RECT 125.555 -82.158 125.645 -81.15 ;
      RECT 125.505 -81.555 125.645 -81.385 ;
      RECT 125.555 -80.35 125.645 -79.342 ;
      RECT 125.505 -80.115 125.645 -79.945 ;
      RECT 125.555 -78.928 125.645 -77.92 ;
      RECT 125.505 -78.325 125.645 -78.155 ;
      RECT 125.555 -77.12 125.645 -76.112 ;
      RECT 125.505 -76.885 125.645 -76.715 ;
      RECT 125.555 -75.698 125.645 -74.69 ;
      RECT 125.505 -75.095 125.645 -74.925 ;
      RECT 125.555 -73.89 125.645 -72.882 ;
      RECT 125.505 -73.655 125.645 -73.485 ;
      RECT 125.555 -72.468 125.645 -71.46 ;
      RECT 125.505 -71.865 125.645 -71.695 ;
      RECT 125.555 -70.66 125.645 -69.652 ;
      RECT 125.505 -70.425 125.645 -70.255 ;
      RECT 125.555 -69.238 125.645 -68.23 ;
      RECT 125.505 -68.635 125.645 -68.465 ;
      RECT 125.555 -67.43 125.645 -66.422 ;
      RECT 125.505 -67.195 125.645 -67.025 ;
      RECT 125.555 -66.008 125.645 -65 ;
      RECT 125.505 -65.405 125.645 -65.235 ;
      RECT 125.555 -64.2 125.645 -63.192 ;
      RECT 125.505 -63.965 125.645 -63.795 ;
      RECT 125.555 -62.778 125.645 -61.77 ;
      RECT 125.505 -62.175 125.645 -62.005 ;
      RECT 125.555 -60.97 125.645 -59.962 ;
      RECT 125.505 -60.735 125.645 -60.565 ;
      RECT 125.555 -59.548 125.645 -58.54 ;
      RECT 125.505 -58.945 125.645 -58.775 ;
      RECT 125.555 -57.74 125.645 -56.732 ;
      RECT 125.505 -57.505 125.645 -57.335 ;
      RECT 125.555 -56.318 125.645 -55.31 ;
      RECT 125.505 -55.715 125.645 -55.545 ;
      RECT 125.555 -54.51 125.645 -53.502 ;
      RECT 125.505 -54.275 125.645 -54.105 ;
      RECT 125.555 -53.088 125.645 -52.08 ;
      RECT 125.505 -52.485 125.645 -52.315 ;
      RECT 125.555 -51.28 125.645 -50.272 ;
      RECT 125.505 -51.045 125.645 -50.875 ;
      RECT 125.555 -49.858 125.645 -48.85 ;
      RECT 125.505 -49.255 125.645 -49.085 ;
      RECT 125.555 -48.05 125.645 -47.042 ;
      RECT 125.505 -47.815 125.645 -47.645 ;
      RECT 125.555 -46.628 125.645 -45.62 ;
      RECT 125.505 -46.025 125.645 -45.855 ;
      RECT 125.555 -44.82 125.645 -43.812 ;
      RECT 125.505 -44.585 125.645 -44.415 ;
      RECT 125.555 -43.398 125.645 -42.39 ;
      RECT 125.505 -42.795 125.645 -42.625 ;
      RECT 125.555 -41.59 125.645 -40.582 ;
      RECT 125.505 -41.355 125.645 -41.185 ;
      RECT 125.555 -40.168 125.645 -39.16 ;
      RECT 125.505 -39.565 125.645 -39.395 ;
      RECT 125.555 -38.36 125.645 -37.352 ;
      RECT 125.505 -38.125 125.645 -37.955 ;
      RECT 125.555 -36.938 125.645 -35.93 ;
      RECT 125.505 -36.335 125.645 -36.165 ;
      RECT 125.555 -35.13 125.645 -34.122 ;
      RECT 125.505 -34.895 125.645 -34.725 ;
      RECT 125.555 -33.708 125.645 -32.7 ;
      RECT 125.505 -33.105 125.645 -32.935 ;
      RECT 125.555 -31.9 125.645 -30.892 ;
      RECT 125.505 -31.665 125.645 -31.495 ;
      RECT 125.555 -30.478 125.645 -29.47 ;
      RECT 125.505 -29.875 125.645 -29.705 ;
      RECT 125.555 -28.67 125.645 -27.662 ;
      RECT 125.505 -28.435 125.645 -28.265 ;
      RECT 125.555 -27.248 125.645 -26.24 ;
      RECT 125.505 -26.645 125.645 -26.475 ;
      RECT 125.555 -25.44 125.645 -24.432 ;
      RECT 125.505 -25.205 125.645 -25.035 ;
      RECT 125.555 -24.018 125.645 -23.01 ;
      RECT 125.505 -23.415 125.645 -23.245 ;
      RECT 125.555 -22.21 125.645 -21.202 ;
      RECT 125.505 -21.975 125.645 -21.805 ;
      RECT 125.555 -20.788 125.645 -19.78 ;
      RECT 125.505 -20.185 125.645 -20.015 ;
      RECT 125.555 -18.98 125.645 -17.972 ;
      RECT 125.505 -18.745 125.645 -18.575 ;
      RECT 125.555 -17.558 125.645 -16.55 ;
      RECT 125.505 -16.955 125.645 -16.785 ;
      RECT 125.555 -15.75 125.645 -14.742 ;
      RECT 125.505 -15.515 125.645 -15.345 ;
      RECT 125.555 -14.328 125.645 -13.32 ;
      RECT 125.505 -13.725 125.645 -13.555 ;
      RECT 125.555 -12.52 125.645 -11.512 ;
      RECT 125.505 -12.285 125.645 -12.115 ;
      RECT 125.555 -11.098 125.645 -10.09 ;
      RECT 125.505 -10.495 125.645 -10.325 ;
      RECT 125.555 -9.29 125.645 -8.282 ;
      RECT 125.505 -9.055 125.645 -8.885 ;
      RECT 125.555 -7.868 125.645 -6.86 ;
      RECT 125.505 -7.265 125.645 -7.095 ;
      RECT 125.555 -6.06 125.645 -5.052 ;
      RECT 125.505 -5.825 125.645 -5.655 ;
      RECT 125.555 -4.638 125.645 -3.63 ;
      RECT 125.505 -4.035 125.645 -3.865 ;
      RECT 125.555 -2.83 125.645 -1.822 ;
      RECT 125.505 -2.595 125.645 -2.425 ;
      RECT 125.555 -1.408 125.645 -0.4 ;
      RECT 125.505 -0.805 125.645 -0.635 ;
      RECT 125.555 0.4 125.645 1.408 ;
      RECT 125.505 0.635 125.645 0.805 ;
      RECT 125.155 -101.538 125.245 -100.531 ;
      RECT 125.155 -101.225 125.295 -101.055 ;
      RECT 125.155 -99.729 125.245 -98.722 ;
      RECT 125.155 -99.205 125.295 -99.035 ;
      RECT 125.155 -98.308 125.245 -97.301 ;
      RECT 125.155 -97.995 125.295 -97.825 ;
      RECT 125.155 -96.499 125.245 -95.492 ;
      RECT 125.155 -95.975 125.295 -95.805 ;
      RECT 125.155 -95.078 125.245 -94.071 ;
      RECT 125.155 -94.765 125.295 -94.595 ;
      RECT 125.155 -93.269 125.245 -92.262 ;
      RECT 125.155 -92.745 125.295 -92.575 ;
      RECT 125.155 -91.848 125.245 -90.841 ;
      RECT 125.155 -91.535 125.295 -91.365 ;
      RECT 125.155 -90.039 125.245 -89.032 ;
      RECT 125.155 -89.515 125.295 -89.345 ;
      RECT 125.155 -88.618 125.245 -87.611 ;
      RECT 125.155 -88.305 125.295 -88.135 ;
      RECT 125.155 -86.809 125.245 -85.802 ;
      RECT 125.155 -86.285 125.295 -86.115 ;
      RECT 125.155 -85.388 125.245 -84.381 ;
      RECT 125.155 -85.075 125.295 -84.905 ;
      RECT 125.155 -83.579 125.245 -82.572 ;
      RECT 125.155 -83.055 125.295 -82.885 ;
      RECT 125.155 -82.158 125.245 -81.151 ;
      RECT 125.155 -81.845 125.295 -81.675 ;
      RECT 125.155 -80.349 125.245 -79.342 ;
      RECT 125.155 -79.825 125.295 -79.655 ;
      RECT 125.155 -78.928 125.245 -77.921 ;
      RECT 125.155 -78.615 125.295 -78.445 ;
      RECT 125.155 -77.119 125.245 -76.112 ;
      RECT 125.155 -76.595 125.295 -76.425 ;
      RECT 125.155 -75.698 125.245 -74.691 ;
      RECT 125.155 -75.385 125.295 -75.215 ;
      RECT 125.155 -73.889 125.245 -72.882 ;
      RECT 125.155 -73.365 125.295 -73.195 ;
      RECT 125.155 -72.468 125.245 -71.461 ;
      RECT 125.155 -72.155 125.295 -71.985 ;
      RECT 125.155 -70.659 125.245 -69.652 ;
      RECT 125.155 -70.135 125.295 -69.965 ;
      RECT 125.155 -69.238 125.245 -68.231 ;
      RECT 125.155 -68.925 125.295 -68.755 ;
      RECT 125.155 -67.429 125.245 -66.422 ;
      RECT 125.155 -66.905 125.295 -66.735 ;
      RECT 125.155 -66.008 125.245 -65.001 ;
      RECT 125.155 -65.695 125.295 -65.525 ;
      RECT 125.155 -64.199 125.245 -63.192 ;
      RECT 125.155 -63.675 125.295 -63.505 ;
      RECT 125.155 -62.778 125.245 -61.771 ;
      RECT 125.155 -62.465 125.295 -62.295 ;
      RECT 125.155 -60.969 125.245 -59.962 ;
      RECT 125.155 -60.445 125.295 -60.275 ;
      RECT 125.155 -59.548 125.245 -58.541 ;
      RECT 125.155 -59.235 125.295 -59.065 ;
      RECT 125.155 -57.739 125.245 -56.732 ;
      RECT 125.155 -57.215 125.295 -57.045 ;
      RECT 125.155 -56.318 125.245 -55.311 ;
      RECT 125.155 -56.005 125.295 -55.835 ;
      RECT 125.155 -54.509 125.245 -53.502 ;
      RECT 125.155 -53.985 125.295 -53.815 ;
      RECT 125.155 -53.088 125.245 -52.081 ;
      RECT 125.155 -52.775 125.295 -52.605 ;
      RECT 125.155 -51.279 125.245 -50.272 ;
      RECT 125.155 -50.755 125.295 -50.585 ;
      RECT 125.155 -49.858 125.245 -48.851 ;
      RECT 125.155 -49.545 125.295 -49.375 ;
      RECT 125.155 -48.049 125.245 -47.042 ;
      RECT 125.155 -47.525 125.295 -47.355 ;
      RECT 125.155 -46.628 125.245 -45.621 ;
      RECT 125.155 -46.315 125.295 -46.145 ;
      RECT 125.155 -44.819 125.245 -43.812 ;
      RECT 125.155 -44.295 125.295 -44.125 ;
      RECT 125.155 -43.398 125.245 -42.391 ;
      RECT 125.155 -43.085 125.295 -42.915 ;
      RECT 125.155 -41.589 125.245 -40.582 ;
      RECT 125.155 -41.065 125.295 -40.895 ;
      RECT 125.155 -40.168 125.245 -39.161 ;
      RECT 125.155 -39.855 125.295 -39.685 ;
      RECT 125.155 -38.359 125.245 -37.352 ;
      RECT 125.155 -37.835 125.295 -37.665 ;
      RECT 125.155 -36.938 125.245 -35.931 ;
      RECT 125.155 -36.625 125.295 -36.455 ;
      RECT 125.155 -35.129 125.245 -34.122 ;
      RECT 125.155 -34.605 125.295 -34.435 ;
      RECT 125.155 -33.708 125.245 -32.701 ;
      RECT 125.155 -33.395 125.295 -33.225 ;
      RECT 125.155 -31.899 125.245 -30.892 ;
      RECT 125.155 -31.375 125.295 -31.205 ;
      RECT 125.155 -30.478 125.245 -29.471 ;
      RECT 125.155 -30.165 125.295 -29.995 ;
      RECT 125.155 -28.669 125.245 -27.662 ;
      RECT 125.155 -28.145 125.295 -27.975 ;
      RECT 125.155 -27.248 125.245 -26.241 ;
      RECT 125.155 -26.935 125.295 -26.765 ;
      RECT 125.155 -25.439 125.245 -24.432 ;
      RECT 125.155 -24.915 125.295 -24.745 ;
      RECT 125.155 -24.018 125.245 -23.011 ;
      RECT 125.155 -23.705 125.295 -23.535 ;
      RECT 125.155 -22.209 125.245 -21.202 ;
      RECT 125.155 -21.685 125.295 -21.515 ;
      RECT 125.155 -20.788 125.245 -19.781 ;
      RECT 125.155 -20.475 125.295 -20.305 ;
      RECT 125.155 -18.979 125.245 -17.972 ;
      RECT 125.155 -18.455 125.295 -18.285 ;
      RECT 125.155 -17.558 125.245 -16.551 ;
      RECT 125.155 -17.245 125.295 -17.075 ;
      RECT 125.155 -15.749 125.245 -14.742 ;
      RECT 125.155 -15.225 125.295 -15.055 ;
      RECT 125.155 -14.328 125.245 -13.321 ;
      RECT 125.155 -14.015 125.295 -13.845 ;
      RECT 125.155 -12.519 125.245 -11.512 ;
      RECT 125.155 -11.995 125.295 -11.825 ;
      RECT 125.155 -11.098 125.245 -10.091 ;
      RECT 125.155 -10.785 125.295 -10.615 ;
      RECT 125.155 -9.289 125.245 -8.282 ;
      RECT 125.155 -8.765 125.295 -8.595 ;
      RECT 125.155 -7.868 125.245 -6.861 ;
      RECT 125.155 -7.555 125.295 -7.385 ;
      RECT 125.155 -6.059 125.245 -5.052 ;
      RECT 125.155 -5.535 125.295 -5.365 ;
      RECT 125.155 -4.638 125.245 -3.631 ;
      RECT 125.155 -4.325 125.295 -4.155 ;
      RECT 125.155 -2.829 125.245 -1.822 ;
      RECT 125.155 -2.305 125.295 -2.135 ;
      RECT 125.155 -1.408 125.245 -0.401 ;
      RECT 125.155 -1.095 125.295 -0.925 ;
      RECT 125.155 0.401 125.245 1.408 ;
      RECT 125.155 0.925 125.295 1.095 ;
      RECT 120.985 -108.935 124.765 -108.815 ;
      RECT 122.305 -109.475 122.405 -108.815 ;
      RECT 121.745 -109.475 121.845 -108.815 ;
      RECT 121.185 -109.475 121.285 -108.815 ;
      RECT 124.355 -101.538 124.445 -100.53 ;
      RECT 124.305 -100.935 124.445 -100.765 ;
      RECT 124.355 -99.73 124.445 -98.722 ;
      RECT 124.305 -99.495 124.445 -99.325 ;
      RECT 124.355 -98.308 124.445 -97.3 ;
      RECT 124.305 -97.705 124.445 -97.535 ;
      RECT 124.355 -96.5 124.445 -95.492 ;
      RECT 124.305 -96.265 124.445 -96.095 ;
      RECT 124.355 -95.078 124.445 -94.07 ;
      RECT 124.305 -94.475 124.445 -94.305 ;
      RECT 124.355 -93.27 124.445 -92.262 ;
      RECT 124.305 -93.035 124.445 -92.865 ;
      RECT 124.355 -91.848 124.445 -90.84 ;
      RECT 124.305 -91.245 124.445 -91.075 ;
      RECT 124.355 -90.04 124.445 -89.032 ;
      RECT 124.305 -89.805 124.445 -89.635 ;
      RECT 124.355 -88.618 124.445 -87.61 ;
      RECT 124.305 -88.015 124.445 -87.845 ;
      RECT 124.355 -86.81 124.445 -85.802 ;
      RECT 124.305 -86.575 124.445 -86.405 ;
      RECT 124.355 -85.388 124.445 -84.38 ;
      RECT 124.305 -84.785 124.445 -84.615 ;
      RECT 124.355 -83.58 124.445 -82.572 ;
      RECT 124.305 -83.345 124.445 -83.175 ;
      RECT 124.355 -82.158 124.445 -81.15 ;
      RECT 124.305 -81.555 124.445 -81.385 ;
      RECT 124.355 -80.35 124.445 -79.342 ;
      RECT 124.305 -80.115 124.445 -79.945 ;
      RECT 124.355 -78.928 124.445 -77.92 ;
      RECT 124.305 -78.325 124.445 -78.155 ;
      RECT 124.355 -77.12 124.445 -76.112 ;
      RECT 124.305 -76.885 124.445 -76.715 ;
      RECT 124.355 -75.698 124.445 -74.69 ;
      RECT 124.305 -75.095 124.445 -74.925 ;
      RECT 124.355 -73.89 124.445 -72.882 ;
      RECT 124.305 -73.655 124.445 -73.485 ;
      RECT 124.355 -72.468 124.445 -71.46 ;
      RECT 124.305 -71.865 124.445 -71.695 ;
      RECT 124.355 -70.66 124.445 -69.652 ;
      RECT 124.305 -70.425 124.445 -70.255 ;
      RECT 124.355 -69.238 124.445 -68.23 ;
      RECT 124.305 -68.635 124.445 -68.465 ;
      RECT 124.355 -67.43 124.445 -66.422 ;
      RECT 124.305 -67.195 124.445 -67.025 ;
      RECT 124.355 -66.008 124.445 -65 ;
      RECT 124.305 -65.405 124.445 -65.235 ;
      RECT 124.355 -64.2 124.445 -63.192 ;
      RECT 124.305 -63.965 124.445 -63.795 ;
      RECT 124.355 -62.778 124.445 -61.77 ;
      RECT 124.305 -62.175 124.445 -62.005 ;
      RECT 124.355 -60.97 124.445 -59.962 ;
      RECT 124.305 -60.735 124.445 -60.565 ;
      RECT 124.355 -59.548 124.445 -58.54 ;
      RECT 124.305 -58.945 124.445 -58.775 ;
      RECT 124.355 -57.74 124.445 -56.732 ;
      RECT 124.305 -57.505 124.445 -57.335 ;
      RECT 124.355 -56.318 124.445 -55.31 ;
      RECT 124.305 -55.715 124.445 -55.545 ;
      RECT 124.355 -54.51 124.445 -53.502 ;
      RECT 124.305 -54.275 124.445 -54.105 ;
      RECT 124.355 -53.088 124.445 -52.08 ;
      RECT 124.305 -52.485 124.445 -52.315 ;
      RECT 124.355 -51.28 124.445 -50.272 ;
      RECT 124.305 -51.045 124.445 -50.875 ;
      RECT 124.355 -49.858 124.445 -48.85 ;
      RECT 124.305 -49.255 124.445 -49.085 ;
      RECT 124.355 -48.05 124.445 -47.042 ;
      RECT 124.305 -47.815 124.445 -47.645 ;
      RECT 124.355 -46.628 124.445 -45.62 ;
      RECT 124.305 -46.025 124.445 -45.855 ;
      RECT 124.355 -44.82 124.445 -43.812 ;
      RECT 124.305 -44.585 124.445 -44.415 ;
      RECT 124.355 -43.398 124.445 -42.39 ;
      RECT 124.305 -42.795 124.445 -42.625 ;
      RECT 124.355 -41.59 124.445 -40.582 ;
      RECT 124.305 -41.355 124.445 -41.185 ;
      RECT 124.355 -40.168 124.445 -39.16 ;
      RECT 124.305 -39.565 124.445 -39.395 ;
      RECT 124.355 -38.36 124.445 -37.352 ;
      RECT 124.305 -38.125 124.445 -37.955 ;
      RECT 124.355 -36.938 124.445 -35.93 ;
      RECT 124.305 -36.335 124.445 -36.165 ;
      RECT 124.355 -35.13 124.445 -34.122 ;
      RECT 124.305 -34.895 124.445 -34.725 ;
      RECT 124.355 -33.708 124.445 -32.7 ;
      RECT 124.305 -33.105 124.445 -32.935 ;
      RECT 124.355 -31.9 124.445 -30.892 ;
      RECT 124.305 -31.665 124.445 -31.495 ;
      RECT 124.355 -30.478 124.445 -29.47 ;
      RECT 124.305 -29.875 124.445 -29.705 ;
      RECT 124.355 -28.67 124.445 -27.662 ;
      RECT 124.305 -28.435 124.445 -28.265 ;
      RECT 124.355 -27.248 124.445 -26.24 ;
      RECT 124.305 -26.645 124.445 -26.475 ;
      RECT 124.355 -25.44 124.445 -24.432 ;
      RECT 124.305 -25.205 124.445 -25.035 ;
      RECT 124.355 -24.018 124.445 -23.01 ;
      RECT 124.305 -23.415 124.445 -23.245 ;
      RECT 124.355 -22.21 124.445 -21.202 ;
      RECT 124.305 -21.975 124.445 -21.805 ;
      RECT 124.355 -20.788 124.445 -19.78 ;
      RECT 124.305 -20.185 124.445 -20.015 ;
      RECT 124.355 -18.98 124.445 -17.972 ;
      RECT 124.305 -18.745 124.445 -18.575 ;
      RECT 124.355 -17.558 124.445 -16.55 ;
      RECT 124.305 -16.955 124.445 -16.785 ;
      RECT 124.355 -15.75 124.445 -14.742 ;
      RECT 124.305 -15.515 124.445 -15.345 ;
      RECT 124.355 -14.328 124.445 -13.32 ;
      RECT 124.305 -13.725 124.445 -13.555 ;
      RECT 124.355 -12.52 124.445 -11.512 ;
      RECT 124.305 -12.285 124.445 -12.115 ;
      RECT 124.355 -11.098 124.445 -10.09 ;
      RECT 124.305 -10.495 124.445 -10.325 ;
      RECT 124.355 -9.29 124.445 -8.282 ;
      RECT 124.305 -9.055 124.445 -8.885 ;
      RECT 124.355 -7.868 124.445 -6.86 ;
      RECT 124.305 -7.265 124.445 -7.095 ;
      RECT 124.355 -6.06 124.445 -5.052 ;
      RECT 124.305 -5.825 124.445 -5.655 ;
      RECT 124.355 -4.638 124.445 -3.63 ;
      RECT 124.305 -4.035 124.445 -3.865 ;
      RECT 124.355 -2.83 124.445 -1.822 ;
      RECT 124.305 -2.595 124.445 -2.425 ;
      RECT 124.355 -1.408 124.445 -0.4 ;
      RECT 124.305 -0.805 124.445 -0.635 ;
      RECT 124.355 0.4 124.445 1.408 ;
      RECT 124.305 0.635 124.445 0.805 ;
      RECT 122.925 -111.685 124.405 -111.585 ;
      RECT 122.925 -112.195 123.025 -111.585 ;
      RECT 123.145 -109.15 124.405 -109.05 ;
      RECT 124.305 -109.475 124.405 -109.05 ;
      RECT 123.745 -109.475 123.845 -109.05 ;
      RECT 123.185 -109.475 123.285 -109.05 ;
      RECT 123.955 -101.538 124.045 -100.531 ;
      RECT 123.955 -101.225 124.095 -101.055 ;
      RECT 123.955 -99.729 124.045 -98.722 ;
      RECT 123.955 -99.205 124.095 -99.035 ;
      RECT 123.955 -98.308 124.045 -97.301 ;
      RECT 123.955 -97.995 124.095 -97.825 ;
      RECT 123.955 -96.499 124.045 -95.492 ;
      RECT 123.955 -95.975 124.095 -95.805 ;
      RECT 123.955 -95.078 124.045 -94.071 ;
      RECT 123.955 -94.765 124.095 -94.595 ;
      RECT 123.955 -93.269 124.045 -92.262 ;
      RECT 123.955 -92.745 124.095 -92.575 ;
      RECT 123.955 -91.848 124.045 -90.841 ;
      RECT 123.955 -91.535 124.095 -91.365 ;
      RECT 123.955 -90.039 124.045 -89.032 ;
      RECT 123.955 -89.515 124.095 -89.345 ;
      RECT 123.955 -88.618 124.045 -87.611 ;
      RECT 123.955 -88.305 124.095 -88.135 ;
      RECT 123.955 -86.809 124.045 -85.802 ;
      RECT 123.955 -86.285 124.095 -86.115 ;
      RECT 123.955 -85.388 124.045 -84.381 ;
      RECT 123.955 -85.075 124.095 -84.905 ;
      RECT 123.955 -83.579 124.045 -82.572 ;
      RECT 123.955 -83.055 124.095 -82.885 ;
      RECT 123.955 -82.158 124.045 -81.151 ;
      RECT 123.955 -81.845 124.095 -81.675 ;
      RECT 123.955 -80.349 124.045 -79.342 ;
      RECT 123.955 -79.825 124.095 -79.655 ;
      RECT 123.955 -78.928 124.045 -77.921 ;
      RECT 123.955 -78.615 124.095 -78.445 ;
      RECT 123.955 -77.119 124.045 -76.112 ;
      RECT 123.955 -76.595 124.095 -76.425 ;
      RECT 123.955 -75.698 124.045 -74.691 ;
      RECT 123.955 -75.385 124.095 -75.215 ;
      RECT 123.955 -73.889 124.045 -72.882 ;
      RECT 123.955 -73.365 124.095 -73.195 ;
      RECT 123.955 -72.468 124.045 -71.461 ;
      RECT 123.955 -72.155 124.095 -71.985 ;
      RECT 123.955 -70.659 124.045 -69.652 ;
      RECT 123.955 -70.135 124.095 -69.965 ;
      RECT 123.955 -69.238 124.045 -68.231 ;
      RECT 123.955 -68.925 124.095 -68.755 ;
      RECT 123.955 -67.429 124.045 -66.422 ;
      RECT 123.955 -66.905 124.095 -66.735 ;
      RECT 123.955 -66.008 124.045 -65.001 ;
      RECT 123.955 -65.695 124.095 -65.525 ;
      RECT 123.955 -64.199 124.045 -63.192 ;
      RECT 123.955 -63.675 124.095 -63.505 ;
      RECT 123.955 -62.778 124.045 -61.771 ;
      RECT 123.955 -62.465 124.095 -62.295 ;
      RECT 123.955 -60.969 124.045 -59.962 ;
      RECT 123.955 -60.445 124.095 -60.275 ;
      RECT 123.955 -59.548 124.045 -58.541 ;
      RECT 123.955 -59.235 124.095 -59.065 ;
      RECT 123.955 -57.739 124.045 -56.732 ;
      RECT 123.955 -57.215 124.095 -57.045 ;
      RECT 123.955 -56.318 124.045 -55.311 ;
      RECT 123.955 -56.005 124.095 -55.835 ;
      RECT 123.955 -54.509 124.045 -53.502 ;
      RECT 123.955 -53.985 124.095 -53.815 ;
      RECT 123.955 -53.088 124.045 -52.081 ;
      RECT 123.955 -52.775 124.095 -52.605 ;
      RECT 123.955 -51.279 124.045 -50.272 ;
      RECT 123.955 -50.755 124.095 -50.585 ;
      RECT 123.955 -49.858 124.045 -48.851 ;
      RECT 123.955 -49.545 124.095 -49.375 ;
      RECT 123.955 -48.049 124.045 -47.042 ;
      RECT 123.955 -47.525 124.095 -47.355 ;
      RECT 123.955 -46.628 124.045 -45.621 ;
      RECT 123.955 -46.315 124.095 -46.145 ;
      RECT 123.955 -44.819 124.045 -43.812 ;
      RECT 123.955 -44.295 124.095 -44.125 ;
      RECT 123.955 -43.398 124.045 -42.391 ;
      RECT 123.955 -43.085 124.095 -42.915 ;
      RECT 123.955 -41.589 124.045 -40.582 ;
      RECT 123.955 -41.065 124.095 -40.895 ;
      RECT 123.955 -40.168 124.045 -39.161 ;
      RECT 123.955 -39.855 124.095 -39.685 ;
      RECT 123.955 -38.359 124.045 -37.352 ;
      RECT 123.955 -37.835 124.095 -37.665 ;
      RECT 123.955 -36.938 124.045 -35.931 ;
      RECT 123.955 -36.625 124.095 -36.455 ;
      RECT 123.955 -35.129 124.045 -34.122 ;
      RECT 123.955 -34.605 124.095 -34.435 ;
      RECT 123.955 -33.708 124.045 -32.701 ;
      RECT 123.955 -33.395 124.095 -33.225 ;
      RECT 123.955 -31.899 124.045 -30.892 ;
      RECT 123.955 -31.375 124.095 -31.205 ;
      RECT 123.955 -30.478 124.045 -29.471 ;
      RECT 123.955 -30.165 124.095 -29.995 ;
      RECT 123.955 -28.669 124.045 -27.662 ;
      RECT 123.955 -28.145 124.095 -27.975 ;
      RECT 123.955 -27.248 124.045 -26.241 ;
      RECT 123.955 -26.935 124.095 -26.765 ;
      RECT 123.955 -25.439 124.045 -24.432 ;
      RECT 123.955 -24.915 124.095 -24.745 ;
      RECT 123.955 -24.018 124.045 -23.011 ;
      RECT 123.955 -23.705 124.095 -23.535 ;
      RECT 123.955 -22.209 124.045 -21.202 ;
      RECT 123.955 -21.685 124.095 -21.515 ;
      RECT 123.955 -20.788 124.045 -19.781 ;
      RECT 123.955 -20.475 124.095 -20.305 ;
      RECT 123.955 -18.979 124.045 -17.972 ;
      RECT 123.955 -18.455 124.095 -18.285 ;
      RECT 123.955 -17.558 124.045 -16.551 ;
      RECT 123.955 -17.245 124.095 -17.075 ;
      RECT 123.955 -15.749 124.045 -14.742 ;
      RECT 123.955 -15.225 124.095 -15.055 ;
      RECT 123.955 -14.328 124.045 -13.321 ;
      RECT 123.955 -14.015 124.095 -13.845 ;
      RECT 123.955 -12.519 124.045 -11.512 ;
      RECT 123.955 -11.995 124.095 -11.825 ;
      RECT 123.955 -11.098 124.045 -10.091 ;
      RECT 123.955 -10.785 124.095 -10.615 ;
      RECT 123.955 -9.289 124.045 -8.282 ;
      RECT 123.955 -8.765 124.095 -8.595 ;
      RECT 123.955 -7.868 124.045 -6.861 ;
      RECT 123.955 -7.555 124.095 -7.385 ;
      RECT 123.955 -6.059 124.045 -5.052 ;
      RECT 123.955 -5.535 124.095 -5.365 ;
      RECT 123.955 -4.638 124.045 -3.631 ;
      RECT 123.955 -4.325 124.095 -4.155 ;
      RECT 123.955 -2.829 124.045 -1.822 ;
      RECT 123.955 -2.305 124.095 -2.135 ;
      RECT 123.955 -1.408 124.045 -0.401 ;
      RECT 123.955 -1.095 124.095 -0.925 ;
      RECT 123.955 0.401 124.045 1.408 ;
      RECT 123.955 0.925 124.095 1.095 ;
      RECT 123.285 -111.495 123.455 -111.385 ;
      RECT 120.135 -111.495 123.455 -111.395 ;
      RECT 123.155 -101.538 123.245 -100.53 ;
      RECT 123.105 -100.935 123.245 -100.765 ;
      RECT 123.155 -99.73 123.245 -98.722 ;
      RECT 123.105 -99.495 123.245 -99.325 ;
      RECT 123.155 -98.308 123.245 -97.3 ;
      RECT 123.105 -97.705 123.245 -97.535 ;
      RECT 123.155 -96.5 123.245 -95.492 ;
      RECT 123.105 -96.265 123.245 -96.095 ;
      RECT 123.155 -95.078 123.245 -94.07 ;
      RECT 123.105 -94.475 123.245 -94.305 ;
      RECT 123.155 -93.27 123.245 -92.262 ;
      RECT 123.105 -93.035 123.245 -92.865 ;
      RECT 123.155 -91.848 123.245 -90.84 ;
      RECT 123.105 -91.245 123.245 -91.075 ;
      RECT 123.155 -90.04 123.245 -89.032 ;
      RECT 123.105 -89.805 123.245 -89.635 ;
      RECT 123.155 -88.618 123.245 -87.61 ;
      RECT 123.105 -88.015 123.245 -87.845 ;
      RECT 123.155 -86.81 123.245 -85.802 ;
      RECT 123.105 -86.575 123.245 -86.405 ;
      RECT 123.155 -85.388 123.245 -84.38 ;
      RECT 123.105 -84.785 123.245 -84.615 ;
      RECT 123.155 -83.58 123.245 -82.572 ;
      RECT 123.105 -83.345 123.245 -83.175 ;
      RECT 123.155 -82.158 123.245 -81.15 ;
      RECT 123.105 -81.555 123.245 -81.385 ;
      RECT 123.155 -80.35 123.245 -79.342 ;
      RECT 123.105 -80.115 123.245 -79.945 ;
      RECT 123.155 -78.928 123.245 -77.92 ;
      RECT 123.105 -78.325 123.245 -78.155 ;
      RECT 123.155 -77.12 123.245 -76.112 ;
      RECT 123.105 -76.885 123.245 -76.715 ;
      RECT 123.155 -75.698 123.245 -74.69 ;
      RECT 123.105 -75.095 123.245 -74.925 ;
      RECT 123.155 -73.89 123.245 -72.882 ;
      RECT 123.105 -73.655 123.245 -73.485 ;
      RECT 123.155 -72.468 123.245 -71.46 ;
      RECT 123.105 -71.865 123.245 -71.695 ;
      RECT 123.155 -70.66 123.245 -69.652 ;
      RECT 123.105 -70.425 123.245 -70.255 ;
      RECT 123.155 -69.238 123.245 -68.23 ;
      RECT 123.105 -68.635 123.245 -68.465 ;
      RECT 123.155 -67.43 123.245 -66.422 ;
      RECT 123.105 -67.195 123.245 -67.025 ;
      RECT 123.155 -66.008 123.245 -65 ;
      RECT 123.105 -65.405 123.245 -65.235 ;
      RECT 123.155 -64.2 123.245 -63.192 ;
      RECT 123.105 -63.965 123.245 -63.795 ;
      RECT 123.155 -62.778 123.245 -61.77 ;
      RECT 123.105 -62.175 123.245 -62.005 ;
      RECT 123.155 -60.97 123.245 -59.962 ;
      RECT 123.105 -60.735 123.245 -60.565 ;
      RECT 123.155 -59.548 123.245 -58.54 ;
      RECT 123.105 -58.945 123.245 -58.775 ;
      RECT 123.155 -57.74 123.245 -56.732 ;
      RECT 123.105 -57.505 123.245 -57.335 ;
      RECT 123.155 -56.318 123.245 -55.31 ;
      RECT 123.105 -55.715 123.245 -55.545 ;
      RECT 123.155 -54.51 123.245 -53.502 ;
      RECT 123.105 -54.275 123.245 -54.105 ;
      RECT 123.155 -53.088 123.245 -52.08 ;
      RECT 123.105 -52.485 123.245 -52.315 ;
      RECT 123.155 -51.28 123.245 -50.272 ;
      RECT 123.105 -51.045 123.245 -50.875 ;
      RECT 123.155 -49.858 123.245 -48.85 ;
      RECT 123.105 -49.255 123.245 -49.085 ;
      RECT 123.155 -48.05 123.245 -47.042 ;
      RECT 123.105 -47.815 123.245 -47.645 ;
      RECT 123.155 -46.628 123.245 -45.62 ;
      RECT 123.105 -46.025 123.245 -45.855 ;
      RECT 123.155 -44.82 123.245 -43.812 ;
      RECT 123.105 -44.585 123.245 -44.415 ;
      RECT 123.155 -43.398 123.245 -42.39 ;
      RECT 123.105 -42.795 123.245 -42.625 ;
      RECT 123.155 -41.59 123.245 -40.582 ;
      RECT 123.105 -41.355 123.245 -41.185 ;
      RECT 123.155 -40.168 123.245 -39.16 ;
      RECT 123.105 -39.565 123.245 -39.395 ;
      RECT 123.155 -38.36 123.245 -37.352 ;
      RECT 123.105 -38.125 123.245 -37.955 ;
      RECT 123.155 -36.938 123.245 -35.93 ;
      RECT 123.105 -36.335 123.245 -36.165 ;
      RECT 123.155 -35.13 123.245 -34.122 ;
      RECT 123.105 -34.895 123.245 -34.725 ;
      RECT 123.155 -33.708 123.245 -32.7 ;
      RECT 123.105 -33.105 123.245 -32.935 ;
      RECT 123.155 -31.9 123.245 -30.892 ;
      RECT 123.105 -31.665 123.245 -31.495 ;
      RECT 123.155 -30.478 123.245 -29.47 ;
      RECT 123.105 -29.875 123.245 -29.705 ;
      RECT 123.155 -28.67 123.245 -27.662 ;
      RECT 123.105 -28.435 123.245 -28.265 ;
      RECT 123.155 -27.248 123.245 -26.24 ;
      RECT 123.105 -26.645 123.245 -26.475 ;
      RECT 123.155 -25.44 123.245 -24.432 ;
      RECT 123.105 -25.205 123.245 -25.035 ;
      RECT 123.155 -24.018 123.245 -23.01 ;
      RECT 123.105 -23.415 123.245 -23.245 ;
      RECT 123.155 -22.21 123.245 -21.202 ;
      RECT 123.105 -21.975 123.245 -21.805 ;
      RECT 123.155 -20.788 123.245 -19.78 ;
      RECT 123.105 -20.185 123.245 -20.015 ;
      RECT 123.155 -18.98 123.245 -17.972 ;
      RECT 123.105 -18.745 123.245 -18.575 ;
      RECT 123.155 -17.558 123.245 -16.55 ;
      RECT 123.105 -16.955 123.245 -16.785 ;
      RECT 123.155 -15.75 123.245 -14.742 ;
      RECT 123.105 -15.515 123.245 -15.345 ;
      RECT 123.155 -14.328 123.245 -13.32 ;
      RECT 123.105 -13.725 123.245 -13.555 ;
      RECT 123.155 -12.52 123.245 -11.512 ;
      RECT 123.105 -12.285 123.245 -12.115 ;
      RECT 123.155 -11.098 123.245 -10.09 ;
      RECT 123.105 -10.495 123.245 -10.325 ;
      RECT 123.155 -9.29 123.245 -8.282 ;
      RECT 123.105 -9.055 123.245 -8.885 ;
      RECT 123.155 -7.868 123.245 -6.86 ;
      RECT 123.105 -7.265 123.245 -7.095 ;
      RECT 123.155 -6.06 123.245 -5.052 ;
      RECT 123.105 -5.825 123.245 -5.655 ;
      RECT 123.155 -4.638 123.245 -3.63 ;
      RECT 123.105 -4.035 123.245 -3.865 ;
      RECT 123.155 -2.83 123.245 -1.822 ;
      RECT 123.105 -2.595 123.245 -2.425 ;
      RECT 123.155 -1.408 123.245 -0.4 ;
      RECT 123.105 -0.805 123.245 -0.635 ;
      RECT 123.155 0.4 123.245 1.408 ;
      RECT 123.105 0.635 123.245 0.805 ;
      RECT 122.755 -101.538 122.845 -100.531 ;
      RECT 122.755 -101.225 122.895 -101.055 ;
      RECT 122.755 -99.729 122.845 -98.722 ;
      RECT 122.755 -99.205 122.895 -99.035 ;
      RECT 122.755 -98.308 122.845 -97.301 ;
      RECT 122.755 -97.995 122.895 -97.825 ;
      RECT 122.755 -96.499 122.845 -95.492 ;
      RECT 122.755 -95.975 122.895 -95.805 ;
      RECT 122.755 -95.078 122.845 -94.071 ;
      RECT 122.755 -94.765 122.895 -94.595 ;
      RECT 122.755 -93.269 122.845 -92.262 ;
      RECT 122.755 -92.745 122.895 -92.575 ;
      RECT 122.755 -91.848 122.845 -90.841 ;
      RECT 122.755 -91.535 122.895 -91.365 ;
      RECT 122.755 -90.039 122.845 -89.032 ;
      RECT 122.755 -89.515 122.895 -89.345 ;
      RECT 122.755 -88.618 122.845 -87.611 ;
      RECT 122.755 -88.305 122.895 -88.135 ;
      RECT 122.755 -86.809 122.845 -85.802 ;
      RECT 122.755 -86.285 122.895 -86.115 ;
      RECT 122.755 -85.388 122.845 -84.381 ;
      RECT 122.755 -85.075 122.895 -84.905 ;
      RECT 122.755 -83.579 122.845 -82.572 ;
      RECT 122.755 -83.055 122.895 -82.885 ;
      RECT 122.755 -82.158 122.845 -81.151 ;
      RECT 122.755 -81.845 122.895 -81.675 ;
      RECT 122.755 -80.349 122.845 -79.342 ;
      RECT 122.755 -79.825 122.895 -79.655 ;
      RECT 122.755 -78.928 122.845 -77.921 ;
      RECT 122.755 -78.615 122.895 -78.445 ;
      RECT 122.755 -77.119 122.845 -76.112 ;
      RECT 122.755 -76.595 122.895 -76.425 ;
      RECT 122.755 -75.698 122.845 -74.691 ;
      RECT 122.755 -75.385 122.895 -75.215 ;
      RECT 122.755 -73.889 122.845 -72.882 ;
      RECT 122.755 -73.365 122.895 -73.195 ;
      RECT 122.755 -72.468 122.845 -71.461 ;
      RECT 122.755 -72.155 122.895 -71.985 ;
      RECT 122.755 -70.659 122.845 -69.652 ;
      RECT 122.755 -70.135 122.895 -69.965 ;
      RECT 122.755 -69.238 122.845 -68.231 ;
      RECT 122.755 -68.925 122.895 -68.755 ;
      RECT 122.755 -67.429 122.845 -66.422 ;
      RECT 122.755 -66.905 122.895 -66.735 ;
      RECT 122.755 -66.008 122.845 -65.001 ;
      RECT 122.755 -65.695 122.895 -65.525 ;
      RECT 122.755 -64.199 122.845 -63.192 ;
      RECT 122.755 -63.675 122.895 -63.505 ;
      RECT 122.755 -62.778 122.845 -61.771 ;
      RECT 122.755 -62.465 122.895 -62.295 ;
      RECT 122.755 -60.969 122.845 -59.962 ;
      RECT 122.755 -60.445 122.895 -60.275 ;
      RECT 122.755 -59.548 122.845 -58.541 ;
      RECT 122.755 -59.235 122.895 -59.065 ;
      RECT 122.755 -57.739 122.845 -56.732 ;
      RECT 122.755 -57.215 122.895 -57.045 ;
      RECT 122.755 -56.318 122.845 -55.311 ;
      RECT 122.755 -56.005 122.895 -55.835 ;
      RECT 122.755 -54.509 122.845 -53.502 ;
      RECT 122.755 -53.985 122.895 -53.815 ;
      RECT 122.755 -53.088 122.845 -52.081 ;
      RECT 122.755 -52.775 122.895 -52.605 ;
      RECT 122.755 -51.279 122.845 -50.272 ;
      RECT 122.755 -50.755 122.895 -50.585 ;
      RECT 122.755 -49.858 122.845 -48.851 ;
      RECT 122.755 -49.545 122.895 -49.375 ;
      RECT 122.755 -48.049 122.845 -47.042 ;
      RECT 122.755 -47.525 122.895 -47.355 ;
      RECT 122.755 -46.628 122.845 -45.621 ;
      RECT 122.755 -46.315 122.895 -46.145 ;
      RECT 122.755 -44.819 122.845 -43.812 ;
      RECT 122.755 -44.295 122.895 -44.125 ;
      RECT 122.755 -43.398 122.845 -42.391 ;
      RECT 122.755 -43.085 122.895 -42.915 ;
      RECT 122.755 -41.589 122.845 -40.582 ;
      RECT 122.755 -41.065 122.895 -40.895 ;
      RECT 122.755 -40.168 122.845 -39.161 ;
      RECT 122.755 -39.855 122.895 -39.685 ;
      RECT 122.755 -38.359 122.845 -37.352 ;
      RECT 122.755 -37.835 122.895 -37.665 ;
      RECT 122.755 -36.938 122.845 -35.931 ;
      RECT 122.755 -36.625 122.895 -36.455 ;
      RECT 122.755 -35.129 122.845 -34.122 ;
      RECT 122.755 -34.605 122.895 -34.435 ;
      RECT 122.755 -33.708 122.845 -32.701 ;
      RECT 122.755 -33.395 122.895 -33.225 ;
      RECT 122.755 -31.899 122.845 -30.892 ;
      RECT 122.755 -31.375 122.895 -31.205 ;
      RECT 122.755 -30.478 122.845 -29.471 ;
      RECT 122.755 -30.165 122.895 -29.995 ;
      RECT 122.755 -28.669 122.845 -27.662 ;
      RECT 122.755 -28.145 122.895 -27.975 ;
      RECT 122.755 -27.248 122.845 -26.241 ;
      RECT 122.755 -26.935 122.895 -26.765 ;
      RECT 122.755 -25.439 122.845 -24.432 ;
      RECT 122.755 -24.915 122.895 -24.745 ;
      RECT 122.755 -24.018 122.845 -23.011 ;
      RECT 122.755 -23.705 122.895 -23.535 ;
      RECT 122.755 -22.209 122.845 -21.202 ;
      RECT 122.755 -21.685 122.895 -21.515 ;
      RECT 122.755 -20.788 122.845 -19.781 ;
      RECT 122.755 -20.475 122.895 -20.305 ;
      RECT 122.755 -18.979 122.845 -17.972 ;
      RECT 122.755 -18.455 122.895 -18.285 ;
      RECT 122.755 -17.558 122.845 -16.551 ;
      RECT 122.755 -17.245 122.895 -17.075 ;
      RECT 122.755 -15.749 122.845 -14.742 ;
      RECT 122.755 -15.225 122.895 -15.055 ;
      RECT 122.755 -14.328 122.845 -13.321 ;
      RECT 122.755 -14.015 122.895 -13.845 ;
      RECT 122.755 -12.519 122.845 -11.512 ;
      RECT 122.755 -11.995 122.895 -11.825 ;
      RECT 122.755 -11.098 122.845 -10.091 ;
      RECT 122.755 -10.785 122.895 -10.615 ;
      RECT 122.755 -9.289 122.845 -8.282 ;
      RECT 122.755 -8.765 122.895 -8.595 ;
      RECT 122.755 -7.868 122.845 -6.861 ;
      RECT 122.755 -7.555 122.895 -7.385 ;
      RECT 122.755 -6.059 122.845 -5.052 ;
      RECT 122.755 -5.535 122.895 -5.365 ;
      RECT 122.755 -4.638 122.845 -3.631 ;
      RECT 122.755 -4.325 122.895 -4.155 ;
      RECT 122.755 -2.829 122.845 -1.822 ;
      RECT 122.755 -2.305 122.895 -2.135 ;
      RECT 122.755 -1.408 122.845 -0.401 ;
      RECT 122.755 -1.095 122.895 -0.925 ;
      RECT 122.755 0.401 122.845 1.408 ;
      RECT 122.755 0.925 122.895 1.095 ;
      RECT 120.905 -111.685 122.385 -111.585 ;
      RECT 120.905 -112.055 121.005 -111.585 ;
      RECT 120.71 -114.395 122.285 -114.275 ;
      RECT 122.185 -114.895 122.285 -114.275 ;
      RECT 121.59 -114.895 121.69 -114.275 ;
      RECT 120.71 -114.85 120.81 -114.275 ;
      RECT 121.955 -101.538 122.045 -100.53 ;
      RECT 121.905 -100.935 122.045 -100.765 ;
      RECT 121.955 -99.73 122.045 -98.722 ;
      RECT 121.905 -99.495 122.045 -99.325 ;
      RECT 121.955 -98.308 122.045 -97.3 ;
      RECT 121.905 -97.705 122.045 -97.535 ;
      RECT 121.955 -96.5 122.045 -95.492 ;
      RECT 121.905 -96.265 122.045 -96.095 ;
      RECT 121.955 -95.078 122.045 -94.07 ;
      RECT 121.905 -94.475 122.045 -94.305 ;
      RECT 121.955 -93.27 122.045 -92.262 ;
      RECT 121.905 -93.035 122.045 -92.865 ;
      RECT 121.955 -91.848 122.045 -90.84 ;
      RECT 121.905 -91.245 122.045 -91.075 ;
      RECT 121.955 -90.04 122.045 -89.032 ;
      RECT 121.905 -89.805 122.045 -89.635 ;
      RECT 121.955 -88.618 122.045 -87.61 ;
      RECT 121.905 -88.015 122.045 -87.845 ;
      RECT 121.955 -86.81 122.045 -85.802 ;
      RECT 121.905 -86.575 122.045 -86.405 ;
      RECT 121.955 -85.388 122.045 -84.38 ;
      RECT 121.905 -84.785 122.045 -84.615 ;
      RECT 121.955 -83.58 122.045 -82.572 ;
      RECT 121.905 -83.345 122.045 -83.175 ;
      RECT 121.955 -82.158 122.045 -81.15 ;
      RECT 121.905 -81.555 122.045 -81.385 ;
      RECT 121.955 -80.35 122.045 -79.342 ;
      RECT 121.905 -80.115 122.045 -79.945 ;
      RECT 121.955 -78.928 122.045 -77.92 ;
      RECT 121.905 -78.325 122.045 -78.155 ;
      RECT 121.955 -77.12 122.045 -76.112 ;
      RECT 121.905 -76.885 122.045 -76.715 ;
      RECT 121.955 -75.698 122.045 -74.69 ;
      RECT 121.905 -75.095 122.045 -74.925 ;
      RECT 121.955 -73.89 122.045 -72.882 ;
      RECT 121.905 -73.655 122.045 -73.485 ;
      RECT 121.955 -72.468 122.045 -71.46 ;
      RECT 121.905 -71.865 122.045 -71.695 ;
      RECT 121.955 -70.66 122.045 -69.652 ;
      RECT 121.905 -70.425 122.045 -70.255 ;
      RECT 121.955 -69.238 122.045 -68.23 ;
      RECT 121.905 -68.635 122.045 -68.465 ;
      RECT 121.955 -67.43 122.045 -66.422 ;
      RECT 121.905 -67.195 122.045 -67.025 ;
      RECT 121.955 -66.008 122.045 -65 ;
      RECT 121.905 -65.405 122.045 -65.235 ;
      RECT 121.955 -64.2 122.045 -63.192 ;
      RECT 121.905 -63.965 122.045 -63.795 ;
      RECT 121.955 -62.778 122.045 -61.77 ;
      RECT 121.905 -62.175 122.045 -62.005 ;
      RECT 121.955 -60.97 122.045 -59.962 ;
      RECT 121.905 -60.735 122.045 -60.565 ;
      RECT 121.955 -59.548 122.045 -58.54 ;
      RECT 121.905 -58.945 122.045 -58.775 ;
      RECT 121.955 -57.74 122.045 -56.732 ;
      RECT 121.905 -57.505 122.045 -57.335 ;
      RECT 121.955 -56.318 122.045 -55.31 ;
      RECT 121.905 -55.715 122.045 -55.545 ;
      RECT 121.955 -54.51 122.045 -53.502 ;
      RECT 121.905 -54.275 122.045 -54.105 ;
      RECT 121.955 -53.088 122.045 -52.08 ;
      RECT 121.905 -52.485 122.045 -52.315 ;
      RECT 121.955 -51.28 122.045 -50.272 ;
      RECT 121.905 -51.045 122.045 -50.875 ;
      RECT 121.955 -49.858 122.045 -48.85 ;
      RECT 121.905 -49.255 122.045 -49.085 ;
      RECT 121.955 -48.05 122.045 -47.042 ;
      RECT 121.905 -47.815 122.045 -47.645 ;
      RECT 121.955 -46.628 122.045 -45.62 ;
      RECT 121.905 -46.025 122.045 -45.855 ;
      RECT 121.955 -44.82 122.045 -43.812 ;
      RECT 121.905 -44.585 122.045 -44.415 ;
      RECT 121.955 -43.398 122.045 -42.39 ;
      RECT 121.905 -42.795 122.045 -42.625 ;
      RECT 121.955 -41.59 122.045 -40.582 ;
      RECT 121.905 -41.355 122.045 -41.185 ;
      RECT 121.955 -40.168 122.045 -39.16 ;
      RECT 121.905 -39.565 122.045 -39.395 ;
      RECT 121.955 -38.36 122.045 -37.352 ;
      RECT 121.905 -38.125 122.045 -37.955 ;
      RECT 121.955 -36.938 122.045 -35.93 ;
      RECT 121.905 -36.335 122.045 -36.165 ;
      RECT 121.955 -35.13 122.045 -34.122 ;
      RECT 121.905 -34.895 122.045 -34.725 ;
      RECT 121.955 -33.708 122.045 -32.7 ;
      RECT 121.905 -33.105 122.045 -32.935 ;
      RECT 121.955 -31.9 122.045 -30.892 ;
      RECT 121.905 -31.665 122.045 -31.495 ;
      RECT 121.955 -30.478 122.045 -29.47 ;
      RECT 121.905 -29.875 122.045 -29.705 ;
      RECT 121.955 -28.67 122.045 -27.662 ;
      RECT 121.905 -28.435 122.045 -28.265 ;
      RECT 121.955 -27.248 122.045 -26.24 ;
      RECT 121.905 -26.645 122.045 -26.475 ;
      RECT 121.955 -25.44 122.045 -24.432 ;
      RECT 121.905 -25.205 122.045 -25.035 ;
      RECT 121.955 -24.018 122.045 -23.01 ;
      RECT 121.905 -23.415 122.045 -23.245 ;
      RECT 121.955 -22.21 122.045 -21.202 ;
      RECT 121.905 -21.975 122.045 -21.805 ;
      RECT 121.955 -20.788 122.045 -19.78 ;
      RECT 121.905 -20.185 122.045 -20.015 ;
      RECT 121.955 -18.98 122.045 -17.972 ;
      RECT 121.905 -18.745 122.045 -18.575 ;
      RECT 121.955 -17.558 122.045 -16.55 ;
      RECT 121.905 -16.955 122.045 -16.785 ;
      RECT 121.955 -15.75 122.045 -14.742 ;
      RECT 121.905 -15.515 122.045 -15.345 ;
      RECT 121.955 -14.328 122.045 -13.32 ;
      RECT 121.905 -13.725 122.045 -13.555 ;
      RECT 121.955 -12.52 122.045 -11.512 ;
      RECT 121.905 -12.285 122.045 -12.115 ;
      RECT 121.955 -11.098 122.045 -10.09 ;
      RECT 121.905 -10.495 122.045 -10.325 ;
      RECT 121.955 -9.29 122.045 -8.282 ;
      RECT 121.905 -9.055 122.045 -8.885 ;
      RECT 121.955 -7.868 122.045 -6.86 ;
      RECT 121.905 -7.265 122.045 -7.095 ;
      RECT 121.955 -6.06 122.045 -5.052 ;
      RECT 121.905 -5.825 122.045 -5.655 ;
      RECT 121.955 -4.638 122.045 -3.63 ;
      RECT 121.905 -4.035 122.045 -3.865 ;
      RECT 121.955 -2.83 122.045 -1.822 ;
      RECT 121.905 -2.595 122.045 -2.425 ;
      RECT 121.955 -1.408 122.045 -0.4 ;
      RECT 121.905 -0.805 122.045 -0.635 ;
      RECT 121.955 0.4 122.045 1.408 ;
      RECT 121.905 0.635 122.045 0.805 ;
      RECT 121.83 -114.685 122.005 -114.515 ;
      RECT 121.905 -114.895 122.005 -114.515 ;
      RECT 120.945 -113.555 121.045 -113.09 ;
      RECT 121.31 -113.555 121.41 -113.1 ;
      RECT 120.945 -113.555 121.79 -113.385 ;
      RECT 121.555 -101.538 121.645 -100.531 ;
      RECT 121.555 -101.225 121.695 -101.055 ;
      RECT 121.555 -99.729 121.645 -98.722 ;
      RECT 121.555 -99.205 121.695 -99.035 ;
      RECT 121.555 -98.308 121.645 -97.301 ;
      RECT 121.555 -97.995 121.695 -97.825 ;
      RECT 121.555 -96.499 121.645 -95.492 ;
      RECT 121.555 -95.975 121.695 -95.805 ;
      RECT 121.555 -95.078 121.645 -94.071 ;
      RECT 121.555 -94.765 121.695 -94.595 ;
      RECT 121.555 -93.269 121.645 -92.262 ;
      RECT 121.555 -92.745 121.695 -92.575 ;
      RECT 121.555 -91.848 121.645 -90.841 ;
      RECT 121.555 -91.535 121.695 -91.365 ;
      RECT 121.555 -90.039 121.645 -89.032 ;
      RECT 121.555 -89.515 121.695 -89.345 ;
      RECT 121.555 -88.618 121.645 -87.611 ;
      RECT 121.555 -88.305 121.695 -88.135 ;
      RECT 121.555 -86.809 121.645 -85.802 ;
      RECT 121.555 -86.285 121.695 -86.115 ;
      RECT 121.555 -85.388 121.645 -84.381 ;
      RECT 121.555 -85.075 121.695 -84.905 ;
      RECT 121.555 -83.579 121.645 -82.572 ;
      RECT 121.555 -83.055 121.695 -82.885 ;
      RECT 121.555 -82.158 121.645 -81.151 ;
      RECT 121.555 -81.845 121.695 -81.675 ;
      RECT 121.555 -80.349 121.645 -79.342 ;
      RECT 121.555 -79.825 121.695 -79.655 ;
      RECT 121.555 -78.928 121.645 -77.921 ;
      RECT 121.555 -78.615 121.695 -78.445 ;
      RECT 121.555 -77.119 121.645 -76.112 ;
      RECT 121.555 -76.595 121.695 -76.425 ;
      RECT 121.555 -75.698 121.645 -74.691 ;
      RECT 121.555 -75.385 121.695 -75.215 ;
      RECT 121.555 -73.889 121.645 -72.882 ;
      RECT 121.555 -73.365 121.695 -73.195 ;
      RECT 121.555 -72.468 121.645 -71.461 ;
      RECT 121.555 -72.155 121.695 -71.985 ;
      RECT 121.555 -70.659 121.645 -69.652 ;
      RECT 121.555 -70.135 121.695 -69.965 ;
      RECT 121.555 -69.238 121.645 -68.231 ;
      RECT 121.555 -68.925 121.695 -68.755 ;
      RECT 121.555 -67.429 121.645 -66.422 ;
      RECT 121.555 -66.905 121.695 -66.735 ;
      RECT 121.555 -66.008 121.645 -65.001 ;
      RECT 121.555 -65.695 121.695 -65.525 ;
      RECT 121.555 -64.199 121.645 -63.192 ;
      RECT 121.555 -63.675 121.695 -63.505 ;
      RECT 121.555 -62.778 121.645 -61.771 ;
      RECT 121.555 -62.465 121.695 -62.295 ;
      RECT 121.555 -60.969 121.645 -59.962 ;
      RECT 121.555 -60.445 121.695 -60.275 ;
      RECT 121.555 -59.548 121.645 -58.541 ;
      RECT 121.555 -59.235 121.695 -59.065 ;
      RECT 121.555 -57.739 121.645 -56.732 ;
      RECT 121.555 -57.215 121.695 -57.045 ;
      RECT 121.555 -56.318 121.645 -55.311 ;
      RECT 121.555 -56.005 121.695 -55.835 ;
      RECT 121.555 -54.509 121.645 -53.502 ;
      RECT 121.555 -53.985 121.695 -53.815 ;
      RECT 121.555 -53.088 121.645 -52.081 ;
      RECT 121.555 -52.775 121.695 -52.605 ;
      RECT 121.555 -51.279 121.645 -50.272 ;
      RECT 121.555 -50.755 121.695 -50.585 ;
      RECT 121.555 -49.858 121.645 -48.851 ;
      RECT 121.555 -49.545 121.695 -49.375 ;
      RECT 121.555 -48.049 121.645 -47.042 ;
      RECT 121.555 -47.525 121.695 -47.355 ;
      RECT 121.555 -46.628 121.645 -45.621 ;
      RECT 121.555 -46.315 121.695 -46.145 ;
      RECT 121.555 -44.819 121.645 -43.812 ;
      RECT 121.555 -44.295 121.695 -44.125 ;
      RECT 121.555 -43.398 121.645 -42.391 ;
      RECT 121.555 -43.085 121.695 -42.915 ;
      RECT 121.555 -41.589 121.645 -40.582 ;
      RECT 121.555 -41.065 121.695 -40.895 ;
      RECT 121.555 -40.168 121.645 -39.161 ;
      RECT 121.555 -39.855 121.695 -39.685 ;
      RECT 121.555 -38.359 121.645 -37.352 ;
      RECT 121.555 -37.835 121.695 -37.665 ;
      RECT 121.555 -36.938 121.645 -35.931 ;
      RECT 121.555 -36.625 121.695 -36.455 ;
      RECT 121.555 -35.129 121.645 -34.122 ;
      RECT 121.555 -34.605 121.695 -34.435 ;
      RECT 121.555 -33.708 121.645 -32.701 ;
      RECT 121.555 -33.395 121.695 -33.225 ;
      RECT 121.555 -31.899 121.645 -30.892 ;
      RECT 121.555 -31.375 121.695 -31.205 ;
      RECT 121.555 -30.478 121.645 -29.471 ;
      RECT 121.555 -30.165 121.695 -29.995 ;
      RECT 121.555 -28.669 121.645 -27.662 ;
      RECT 121.555 -28.145 121.695 -27.975 ;
      RECT 121.555 -27.248 121.645 -26.241 ;
      RECT 121.555 -26.935 121.695 -26.765 ;
      RECT 121.555 -25.439 121.645 -24.432 ;
      RECT 121.555 -24.915 121.695 -24.745 ;
      RECT 121.555 -24.018 121.645 -23.011 ;
      RECT 121.555 -23.705 121.695 -23.535 ;
      RECT 121.555 -22.209 121.645 -21.202 ;
      RECT 121.555 -21.685 121.695 -21.515 ;
      RECT 121.555 -20.788 121.645 -19.781 ;
      RECT 121.555 -20.475 121.695 -20.305 ;
      RECT 121.555 -18.979 121.645 -17.972 ;
      RECT 121.555 -18.455 121.695 -18.285 ;
      RECT 121.555 -17.558 121.645 -16.551 ;
      RECT 121.555 -17.245 121.695 -17.075 ;
      RECT 121.555 -15.749 121.645 -14.742 ;
      RECT 121.555 -15.225 121.695 -15.055 ;
      RECT 121.555 -14.328 121.645 -13.321 ;
      RECT 121.555 -14.015 121.695 -13.845 ;
      RECT 121.555 -12.519 121.645 -11.512 ;
      RECT 121.555 -11.995 121.695 -11.825 ;
      RECT 121.555 -11.098 121.645 -10.091 ;
      RECT 121.555 -10.785 121.695 -10.615 ;
      RECT 121.555 -9.289 121.645 -8.282 ;
      RECT 121.555 -8.765 121.695 -8.595 ;
      RECT 121.555 -7.868 121.645 -6.861 ;
      RECT 121.555 -7.555 121.695 -7.385 ;
      RECT 121.555 -6.059 121.645 -5.052 ;
      RECT 121.555 -5.535 121.695 -5.365 ;
      RECT 121.555 -4.638 121.645 -3.631 ;
      RECT 121.555 -4.325 121.695 -4.155 ;
      RECT 121.555 -2.829 121.645 -1.822 ;
      RECT 121.555 -2.305 121.695 -2.135 ;
      RECT 121.555 -1.408 121.645 -0.401 ;
      RECT 121.555 -1.095 121.695 -0.925 ;
      RECT 121.555 0.401 121.645 1.408 ;
      RECT 121.555 0.925 121.695 1.095 ;
      RECT 121.24 -114.685 121.41 -114.515 ;
      RECT 121.31 -114.895 121.41 -114.515 ;
      RECT 120.755 -101.538 120.845 -100.53 ;
      RECT 120.705 -100.935 120.845 -100.765 ;
      RECT 120.755 -99.73 120.845 -98.722 ;
      RECT 120.705 -99.495 120.845 -99.325 ;
      RECT 120.755 -98.308 120.845 -97.3 ;
      RECT 120.705 -97.705 120.845 -97.535 ;
      RECT 120.755 -96.5 120.845 -95.492 ;
      RECT 120.705 -96.265 120.845 -96.095 ;
      RECT 120.755 -95.078 120.845 -94.07 ;
      RECT 120.705 -94.475 120.845 -94.305 ;
      RECT 120.755 -93.27 120.845 -92.262 ;
      RECT 120.705 -93.035 120.845 -92.865 ;
      RECT 120.755 -91.848 120.845 -90.84 ;
      RECT 120.705 -91.245 120.845 -91.075 ;
      RECT 120.755 -90.04 120.845 -89.032 ;
      RECT 120.705 -89.805 120.845 -89.635 ;
      RECT 120.755 -88.618 120.845 -87.61 ;
      RECT 120.705 -88.015 120.845 -87.845 ;
      RECT 120.755 -86.81 120.845 -85.802 ;
      RECT 120.705 -86.575 120.845 -86.405 ;
      RECT 120.755 -85.388 120.845 -84.38 ;
      RECT 120.705 -84.785 120.845 -84.615 ;
      RECT 120.755 -83.58 120.845 -82.572 ;
      RECT 120.705 -83.345 120.845 -83.175 ;
      RECT 120.755 -82.158 120.845 -81.15 ;
      RECT 120.705 -81.555 120.845 -81.385 ;
      RECT 120.755 -80.35 120.845 -79.342 ;
      RECT 120.705 -80.115 120.845 -79.945 ;
      RECT 120.755 -78.928 120.845 -77.92 ;
      RECT 120.705 -78.325 120.845 -78.155 ;
      RECT 120.755 -77.12 120.845 -76.112 ;
      RECT 120.705 -76.885 120.845 -76.715 ;
      RECT 120.755 -75.698 120.845 -74.69 ;
      RECT 120.705 -75.095 120.845 -74.925 ;
      RECT 120.755 -73.89 120.845 -72.882 ;
      RECT 120.705 -73.655 120.845 -73.485 ;
      RECT 120.755 -72.468 120.845 -71.46 ;
      RECT 120.705 -71.865 120.845 -71.695 ;
      RECT 120.755 -70.66 120.845 -69.652 ;
      RECT 120.705 -70.425 120.845 -70.255 ;
      RECT 120.755 -69.238 120.845 -68.23 ;
      RECT 120.705 -68.635 120.845 -68.465 ;
      RECT 120.755 -67.43 120.845 -66.422 ;
      RECT 120.705 -67.195 120.845 -67.025 ;
      RECT 120.755 -66.008 120.845 -65 ;
      RECT 120.705 -65.405 120.845 -65.235 ;
      RECT 120.755 -64.2 120.845 -63.192 ;
      RECT 120.705 -63.965 120.845 -63.795 ;
      RECT 120.755 -62.778 120.845 -61.77 ;
      RECT 120.705 -62.175 120.845 -62.005 ;
      RECT 120.755 -60.97 120.845 -59.962 ;
      RECT 120.705 -60.735 120.845 -60.565 ;
      RECT 120.755 -59.548 120.845 -58.54 ;
      RECT 120.705 -58.945 120.845 -58.775 ;
      RECT 120.755 -57.74 120.845 -56.732 ;
      RECT 120.705 -57.505 120.845 -57.335 ;
      RECT 120.755 -56.318 120.845 -55.31 ;
      RECT 120.705 -55.715 120.845 -55.545 ;
      RECT 120.755 -54.51 120.845 -53.502 ;
      RECT 120.705 -54.275 120.845 -54.105 ;
      RECT 120.755 -53.088 120.845 -52.08 ;
      RECT 120.705 -52.485 120.845 -52.315 ;
      RECT 120.755 -51.28 120.845 -50.272 ;
      RECT 120.705 -51.045 120.845 -50.875 ;
      RECT 120.755 -49.858 120.845 -48.85 ;
      RECT 120.705 -49.255 120.845 -49.085 ;
      RECT 120.755 -48.05 120.845 -47.042 ;
      RECT 120.705 -47.815 120.845 -47.645 ;
      RECT 120.755 -46.628 120.845 -45.62 ;
      RECT 120.705 -46.025 120.845 -45.855 ;
      RECT 120.755 -44.82 120.845 -43.812 ;
      RECT 120.705 -44.585 120.845 -44.415 ;
      RECT 120.755 -43.398 120.845 -42.39 ;
      RECT 120.705 -42.795 120.845 -42.625 ;
      RECT 120.755 -41.59 120.845 -40.582 ;
      RECT 120.705 -41.355 120.845 -41.185 ;
      RECT 120.755 -40.168 120.845 -39.16 ;
      RECT 120.705 -39.565 120.845 -39.395 ;
      RECT 120.755 -38.36 120.845 -37.352 ;
      RECT 120.705 -38.125 120.845 -37.955 ;
      RECT 120.755 -36.938 120.845 -35.93 ;
      RECT 120.705 -36.335 120.845 -36.165 ;
      RECT 120.755 -35.13 120.845 -34.122 ;
      RECT 120.705 -34.895 120.845 -34.725 ;
      RECT 120.755 -33.708 120.845 -32.7 ;
      RECT 120.705 -33.105 120.845 -32.935 ;
      RECT 120.755 -31.9 120.845 -30.892 ;
      RECT 120.705 -31.665 120.845 -31.495 ;
      RECT 120.755 -30.478 120.845 -29.47 ;
      RECT 120.705 -29.875 120.845 -29.705 ;
      RECT 120.755 -28.67 120.845 -27.662 ;
      RECT 120.705 -28.435 120.845 -28.265 ;
      RECT 120.755 -27.248 120.845 -26.24 ;
      RECT 120.705 -26.645 120.845 -26.475 ;
      RECT 120.755 -25.44 120.845 -24.432 ;
      RECT 120.705 -25.205 120.845 -25.035 ;
      RECT 120.755 -24.018 120.845 -23.01 ;
      RECT 120.705 -23.415 120.845 -23.245 ;
      RECT 120.755 -22.21 120.845 -21.202 ;
      RECT 120.705 -21.975 120.845 -21.805 ;
      RECT 120.755 -20.788 120.845 -19.78 ;
      RECT 120.705 -20.185 120.845 -20.015 ;
      RECT 120.755 -18.98 120.845 -17.972 ;
      RECT 120.705 -18.745 120.845 -18.575 ;
      RECT 120.755 -17.558 120.845 -16.55 ;
      RECT 120.705 -16.955 120.845 -16.785 ;
      RECT 120.755 -15.75 120.845 -14.742 ;
      RECT 120.705 -15.515 120.845 -15.345 ;
      RECT 120.755 -14.328 120.845 -13.32 ;
      RECT 120.705 -13.725 120.845 -13.555 ;
      RECT 120.755 -12.52 120.845 -11.512 ;
      RECT 120.705 -12.285 120.845 -12.115 ;
      RECT 120.755 -11.098 120.845 -10.09 ;
      RECT 120.705 -10.495 120.845 -10.325 ;
      RECT 120.755 -9.29 120.845 -8.282 ;
      RECT 120.705 -9.055 120.845 -8.885 ;
      RECT 120.755 -7.868 120.845 -6.86 ;
      RECT 120.705 -7.265 120.845 -7.095 ;
      RECT 120.755 -6.06 120.845 -5.052 ;
      RECT 120.705 -5.825 120.845 -5.655 ;
      RECT 120.755 -4.638 120.845 -3.63 ;
      RECT 120.705 -4.035 120.845 -3.865 ;
      RECT 120.755 -2.83 120.845 -1.822 ;
      RECT 120.705 -2.595 120.845 -2.425 ;
      RECT 120.755 -1.408 120.845 -0.4 ;
      RECT 120.705 -0.805 120.845 -0.635 ;
      RECT 120.755 0.4 120.845 1.408 ;
      RECT 120.705 0.635 120.845 0.805 ;
      RECT 120.355 -101.538 120.445 -100.531 ;
      RECT 120.355 -101.225 120.495 -101.055 ;
      RECT 120.355 -99.729 120.445 -98.722 ;
      RECT 120.355 -99.205 120.495 -99.035 ;
      RECT 120.355 -98.308 120.445 -97.301 ;
      RECT 120.355 -97.995 120.495 -97.825 ;
      RECT 120.355 -96.499 120.445 -95.492 ;
      RECT 120.355 -95.975 120.495 -95.805 ;
      RECT 120.355 -95.078 120.445 -94.071 ;
      RECT 120.355 -94.765 120.495 -94.595 ;
      RECT 120.355 -93.269 120.445 -92.262 ;
      RECT 120.355 -92.745 120.495 -92.575 ;
      RECT 120.355 -91.848 120.445 -90.841 ;
      RECT 120.355 -91.535 120.495 -91.365 ;
      RECT 120.355 -90.039 120.445 -89.032 ;
      RECT 120.355 -89.515 120.495 -89.345 ;
      RECT 120.355 -88.618 120.445 -87.611 ;
      RECT 120.355 -88.305 120.495 -88.135 ;
      RECT 120.355 -86.809 120.445 -85.802 ;
      RECT 120.355 -86.285 120.495 -86.115 ;
      RECT 120.355 -85.388 120.445 -84.381 ;
      RECT 120.355 -85.075 120.495 -84.905 ;
      RECT 120.355 -83.579 120.445 -82.572 ;
      RECT 120.355 -83.055 120.495 -82.885 ;
      RECT 120.355 -82.158 120.445 -81.151 ;
      RECT 120.355 -81.845 120.495 -81.675 ;
      RECT 120.355 -80.349 120.445 -79.342 ;
      RECT 120.355 -79.825 120.495 -79.655 ;
      RECT 120.355 -78.928 120.445 -77.921 ;
      RECT 120.355 -78.615 120.495 -78.445 ;
      RECT 120.355 -77.119 120.445 -76.112 ;
      RECT 120.355 -76.595 120.495 -76.425 ;
      RECT 120.355 -75.698 120.445 -74.691 ;
      RECT 120.355 -75.385 120.495 -75.215 ;
      RECT 120.355 -73.889 120.445 -72.882 ;
      RECT 120.355 -73.365 120.495 -73.195 ;
      RECT 120.355 -72.468 120.445 -71.461 ;
      RECT 120.355 -72.155 120.495 -71.985 ;
      RECT 120.355 -70.659 120.445 -69.652 ;
      RECT 120.355 -70.135 120.495 -69.965 ;
      RECT 120.355 -69.238 120.445 -68.231 ;
      RECT 120.355 -68.925 120.495 -68.755 ;
      RECT 120.355 -67.429 120.445 -66.422 ;
      RECT 120.355 -66.905 120.495 -66.735 ;
      RECT 120.355 -66.008 120.445 -65.001 ;
      RECT 120.355 -65.695 120.495 -65.525 ;
      RECT 120.355 -64.199 120.445 -63.192 ;
      RECT 120.355 -63.675 120.495 -63.505 ;
      RECT 120.355 -62.778 120.445 -61.771 ;
      RECT 120.355 -62.465 120.495 -62.295 ;
      RECT 120.355 -60.969 120.445 -59.962 ;
      RECT 120.355 -60.445 120.495 -60.275 ;
      RECT 120.355 -59.548 120.445 -58.541 ;
      RECT 120.355 -59.235 120.495 -59.065 ;
      RECT 120.355 -57.739 120.445 -56.732 ;
      RECT 120.355 -57.215 120.495 -57.045 ;
      RECT 120.355 -56.318 120.445 -55.311 ;
      RECT 120.355 -56.005 120.495 -55.835 ;
      RECT 120.355 -54.509 120.445 -53.502 ;
      RECT 120.355 -53.985 120.495 -53.815 ;
      RECT 120.355 -53.088 120.445 -52.081 ;
      RECT 120.355 -52.775 120.495 -52.605 ;
      RECT 120.355 -51.279 120.445 -50.272 ;
      RECT 120.355 -50.755 120.495 -50.585 ;
      RECT 120.355 -49.858 120.445 -48.851 ;
      RECT 120.355 -49.545 120.495 -49.375 ;
      RECT 120.355 -48.049 120.445 -47.042 ;
      RECT 120.355 -47.525 120.495 -47.355 ;
      RECT 120.355 -46.628 120.445 -45.621 ;
      RECT 120.355 -46.315 120.495 -46.145 ;
      RECT 120.355 -44.819 120.445 -43.812 ;
      RECT 120.355 -44.295 120.495 -44.125 ;
      RECT 120.355 -43.398 120.445 -42.391 ;
      RECT 120.355 -43.085 120.495 -42.915 ;
      RECT 120.355 -41.589 120.445 -40.582 ;
      RECT 120.355 -41.065 120.495 -40.895 ;
      RECT 120.355 -40.168 120.445 -39.161 ;
      RECT 120.355 -39.855 120.495 -39.685 ;
      RECT 120.355 -38.359 120.445 -37.352 ;
      RECT 120.355 -37.835 120.495 -37.665 ;
      RECT 120.355 -36.938 120.445 -35.931 ;
      RECT 120.355 -36.625 120.495 -36.455 ;
      RECT 120.355 -35.129 120.445 -34.122 ;
      RECT 120.355 -34.605 120.495 -34.435 ;
      RECT 120.355 -33.708 120.445 -32.701 ;
      RECT 120.355 -33.395 120.495 -33.225 ;
      RECT 120.355 -31.899 120.445 -30.892 ;
      RECT 120.355 -31.375 120.495 -31.205 ;
      RECT 120.355 -30.478 120.445 -29.471 ;
      RECT 120.355 -30.165 120.495 -29.995 ;
      RECT 120.355 -28.669 120.445 -27.662 ;
      RECT 120.355 -28.145 120.495 -27.975 ;
      RECT 120.355 -27.248 120.445 -26.241 ;
      RECT 120.355 -26.935 120.495 -26.765 ;
      RECT 120.355 -25.439 120.445 -24.432 ;
      RECT 120.355 -24.915 120.495 -24.745 ;
      RECT 120.355 -24.018 120.445 -23.011 ;
      RECT 120.355 -23.705 120.495 -23.535 ;
      RECT 120.355 -22.209 120.445 -21.202 ;
      RECT 120.355 -21.685 120.495 -21.515 ;
      RECT 120.355 -20.788 120.445 -19.781 ;
      RECT 120.355 -20.475 120.495 -20.305 ;
      RECT 120.355 -18.979 120.445 -17.972 ;
      RECT 120.355 -18.455 120.495 -18.285 ;
      RECT 120.355 -17.558 120.445 -16.551 ;
      RECT 120.355 -17.245 120.495 -17.075 ;
      RECT 120.355 -15.749 120.445 -14.742 ;
      RECT 120.355 -15.225 120.495 -15.055 ;
      RECT 120.355 -14.328 120.445 -13.321 ;
      RECT 120.355 -14.015 120.495 -13.845 ;
      RECT 120.355 -12.519 120.445 -11.512 ;
      RECT 120.355 -11.995 120.495 -11.825 ;
      RECT 120.355 -11.098 120.445 -10.091 ;
      RECT 120.355 -10.785 120.495 -10.615 ;
      RECT 120.355 -9.289 120.445 -8.282 ;
      RECT 120.355 -8.765 120.495 -8.595 ;
      RECT 120.355 -7.868 120.445 -6.861 ;
      RECT 120.355 -7.555 120.495 -7.385 ;
      RECT 120.355 -6.059 120.445 -5.052 ;
      RECT 120.355 -5.535 120.495 -5.365 ;
      RECT 120.355 -4.638 120.445 -3.631 ;
      RECT 120.355 -4.325 120.495 -4.155 ;
      RECT 120.355 -2.829 120.445 -1.822 ;
      RECT 120.355 -2.305 120.495 -2.135 ;
      RECT 120.355 -1.408 120.445 -0.401 ;
      RECT 120.355 -1.095 120.495 -0.925 ;
      RECT 120.355 0.401 120.445 1.408 ;
      RECT 120.355 0.925 120.495 1.095 ;
      RECT 116.185 -108.935 119.965 -108.815 ;
      RECT 117.505 -109.475 117.605 -108.815 ;
      RECT 116.945 -109.475 117.045 -108.815 ;
      RECT 116.385 -109.475 116.485 -108.815 ;
      RECT 119.555 -101.538 119.645 -100.53 ;
      RECT 119.505 -100.935 119.645 -100.765 ;
      RECT 119.555 -99.73 119.645 -98.722 ;
      RECT 119.505 -99.495 119.645 -99.325 ;
      RECT 119.555 -98.308 119.645 -97.3 ;
      RECT 119.505 -97.705 119.645 -97.535 ;
      RECT 119.555 -96.5 119.645 -95.492 ;
      RECT 119.505 -96.265 119.645 -96.095 ;
      RECT 119.555 -95.078 119.645 -94.07 ;
      RECT 119.505 -94.475 119.645 -94.305 ;
      RECT 119.555 -93.27 119.645 -92.262 ;
      RECT 119.505 -93.035 119.645 -92.865 ;
      RECT 119.555 -91.848 119.645 -90.84 ;
      RECT 119.505 -91.245 119.645 -91.075 ;
      RECT 119.555 -90.04 119.645 -89.032 ;
      RECT 119.505 -89.805 119.645 -89.635 ;
      RECT 119.555 -88.618 119.645 -87.61 ;
      RECT 119.505 -88.015 119.645 -87.845 ;
      RECT 119.555 -86.81 119.645 -85.802 ;
      RECT 119.505 -86.575 119.645 -86.405 ;
      RECT 119.555 -85.388 119.645 -84.38 ;
      RECT 119.505 -84.785 119.645 -84.615 ;
      RECT 119.555 -83.58 119.645 -82.572 ;
      RECT 119.505 -83.345 119.645 -83.175 ;
      RECT 119.555 -82.158 119.645 -81.15 ;
      RECT 119.505 -81.555 119.645 -81.385 ;
      RECT 119.555 -80.35 119.645 -79.342 ;
      RECT 119.505 -80.115 119.645 -79.945 ;
      RECT 119.555 -78.928 119.645 -77.92 ;
      RECT 119.505 -78.325 119.645 -78.155 ;
      RECT 119.555 -77.12 119.645 -76.112 ;
      RECT 119.505 -76.885 119.645 -76.715 ;
      RECT 119.555 -75.698 119.645 -74.69 ;
      RECT 119.505 -75.095 119.645 -74.925 ;
      RECT 119.555 -73.89 119.645 -72.882 ;
      RECT 119.505 -73.655 119.645 -73.485 ;
      RECT 119.555 -72.468 119.645 -71.46 ;
      RECT 119.505 -71.865 119.645 -71.695 ;
      RECT 119.555 -70.66 119.645 -69.652 ;
      RECT 119.505 -70.425 119.645 -70.255 ;
      RECT 119.555 -69.238 119.645 -68.23 ;
      RECT 119.505 -68.635 119.645 -68.465 ;
      RECT 119.555 -67.43 119.645 -66.422 ;
      RECT 119.505 -67.195 119.645 -67.025 ;
      RECT 119.555 -66.008 119.645 -65 ;
      RECT 119.505 -65.405 119.645 -65.235 ;
      RECT 119.555 -64.2 119.645 -63.192 ;
      RECT 119.505 -63.965 119.645 -63.795 ;
      RECT 119.555 -62.778 119.645 -61.77 ;
      RECT 119.505 -62.175 119.645 -62.005 ;
      RECT 119.555 -60.97 119.645 -59.962 ;
      RECT 119.505 -60.735 119.645 -60.565 ;
      RECT 119.555 -59.548 119.645 -58.54 ;
      RECT 119.505 -58.945 119.645 -58.775 ;
      RECT 119.555 -57.74 119.645 -56.732 ;
      RECT 119.505 -57.505 119.645 -57.335 ;
      RECT 119.555 -56.318 119.645 -55.31 ;
      RECT 119.505 -55.715 119.645 -55.545 ;
      RECT 119.555 -54.51 119.645 -53.502 ;
      RECT 119.505 -54.275 119.645 -54.105 ;
      RECT 119.555 -53.088 119.645 -52.08 ;
      RECT 119.505 -52.485 119.645 -52.315 ;
      RECT 119.555 -51.28 119.645 -50.272 ;
      RECT 119.505 -51.045 119.645 -50.875 ;
      RECT 119.555 -49.858 119.645 -48.85 ;
      RECT 119.505 -49.255 119.645 -49.085 ;
      RECT 119.555 -48.05 119.645 -47.042 ;
      RECT 119.505 -47.815 119.645 -47.645 ;
      RECT 119.555 -46.628 119.645 -45.62 ;
      RECT 119.505 -46.025 119.645 -45.855 ;
      RECT 119.555 -44.82 119.645 -43.812 ;
      RECT 119.505 -44.585 119.645 -44.415 ;
      RECT 119.555 -43.398 119.645 -42.39 ;
      RECT 119.505 -42.795 119.645 -42.625 ;
      RECT 119.555 -41.59 119.645 -40.582 ;
      RECT 119.505 -41.355 119.645 -41.185 ;
      RECT 119.555 -40.168 119.645 -39.16 ;
      RECT 119.505 -39.565 119.645 -39.395 ;
      RECT 119.555 -38.36 119.645 -37.352 ;
      RECT 119.505 -38.125 119.645 -37.955 ;
      RECT 119.555 -36.938 119.645 -35.93 ;
      RECT 119.505 -36.335 119.645 -36.165 ;
      RECT 119.555 -35.13 119.645 -34.122 ;
      RECT 119.505 -34.895 119.645 -34.725 ;
      RECT 119.555 -33.708 119.645 -32.7 ;
      RECT 119.505 -33.105 119.645 -32.935 ;
      RECT 119.555 -31.9 119.645 -30.892 ;
      RECT 119.505 -31.665 119.645 -31.495 ;
      RECT 119.555 -30.478 119.645 -29.47 ;
      RECT 119.505 -29.875 119.645 -29.705 ;
      RECT 119.555 -28.67 119.645 -27.662 ;
      RECT 119.505 -28.435 119.645 -28.265 ;
      RECT 119.555 -27.248 119.645 -26.24 ;
      RECT 119.505 -26.645 119.645 -26.475 ;
      RECT 119.555 -25.44 119.645 -24.432 ;
      RECT 119.505 -25.205 119.645 -25.035 ;
      RECT 119.555 -24.018 119.645 -23.01 ;
      RECT 119.505 -23.415 119.645 -23.245 ;
      RECT 119.555 -22.21 119.645 -21.202 ;
      RECT 119.505 -21.975 119.645 -21.805 ;
      RECT 119.555 -20.788 119.645 -19.78 ;
      RECT 119.505 -20.185 119.645 -20.015 ;
      RECT 119.555 -18.98 119.645 -17.972 ;
      RECT 119.505 -18.745 119.645 -18.575 ;
      RECT 119.555 -17.558 119.645 -16.55 ;
      RECT 119.505 -16.955 119.645 -16.785 ;
      RECT 119.555 -15.75 119.645 -14.742 ;
      RECT 119.505 -15.515 119.645 -15.345 ;
      RECT 119.555 -14.328 119.645 -13.32 ;
      RECT 119.505 -13.725 119.645 -13.555 ;
      RECT 119.555 -12.52 119.645 -11.512 ;
      RECT 119.505 -12.285 119.645 -12.115 ;
      RECT 119.555 -11.098 119.645 -10.09 ;
      RECT 119.505 -10.495 119.645 -10.325 ;
      RECT 119.555 -9.29 119.645 -8.282 ;
      RECT 119.505 -9.055 119.645 -8.885 ;
      RECT 119.555 -7.868 119.645 -6.86 ;
      RECT 119.505 -7.265 119.645 -7.095 ;
      RECT 119.555 -6.06 119.645 -5.052 ;
      RECT 119.505 -5.825 119.645 -5.655 ;
      RECT 119.555 -4.638 119.645 -3.63 ;
      RECT 119.505 -4.035 119.645 -3.865 ;
      RECT 119.555 -2.83 119.645 -1.822 ;
      RECT 119.505 -2.595 119.645 -2.425 ;
      RECT 119.555 -1.408 119.645 -0.4 ;
      RECT 119.505 -0.805 119.645 -0.635 ;
      RECT 119.555 0.4 119.645 1.408 ;
      RECT 119.505 0.635 119.645 0.805 ;
      RECT 118.125 -111.685 119.605 -111.585 ;
      RECT 118.125 -112.195 118.225 -111.585 ;
      RECT 118.345 -109.15 119.605 -109.05 ;
      RECT 119.505 -109.475 119.605 -109.05 ;
      RECT 118.945 -109.475 119.045 -109.05 ;
      RECT 118.385 -109.475 118.485 -109.05 ;
      RECT 119.155 -101.538 119.245 -100.531 ;
      RECT 119.155 -101.225 119.295 -101.055 ;
      RECT 119.155 -99.729 119.245 -98.722 ;
      RECT 119.155 -99.205 119.295 -99.035 ;
      RECT 119.155 -98.308 119.245 -97.301 ;
      RECT 119.155 -97.995 119.295 -97.825 ;
      RECT 119.155 -96.499 119.245 -95.492 ;
      RECT 119.155 -95.975 119.295 -95.805 ;
      RECT 119.155 -95.078 119.245 -94.071 ;
      RECT 119.155 -94.765 119.295 -94.595 ;
      RECT 119.155 -93.269 119.245 -92.262 ;
      RECT 119.155 -92.745 119.295 -92.575 ;
      RECT 119.155 -91.848 119.245 -90.841 ;
      RECT 119.155 -91.535 119.295 -91.365 ;
      RECT 119.155 -90.039 119.245 -89.032 ;
      RECT 119.155 -89.515 119.295 -89.345 ;
      RECT 119.155 -88.618 119.245 -87.611 ;
      RECT 119.155 -88.305 119.295 -88.135 ;
      RECT 119.155 -86.809 119.245 -85.802 ;
      RECT 119.155 -86.285 119.295 -86.115 ;
      RECT 119.155 -85.388 119.245 -84.381 ;
      RECT 119.155 -85.075 119.295 -84.905 ;
      RECT 119.155 -83.579 119.245 -82.572 ;
      RECT 119.155 -83.055 119.295 -82.885 ;
      RECT 119.155 -82.158 119.245 -81.151 ;
      RECT 119.155 -81.845 119.295 -81.675 ;
      RECT 119.155 -80.349 119.245 -79.342 ;
      RECT 119.155 -79.825 119.295 -79.655 ;
      RECT 119.155 -78.928 119.245 -77.921 ;
      RECT 119.155 -78.615 119.295 -78.445 ;
      RECT 119.155 -77.119 119.245 -76.112 ;
      RECT 119.155 -76.595 119.295 -76.425 ;
      RECT 119.155 -75.698 119.245 -74.691 ;
      RECT 119.155 -75.385 119.295 -75.215 ;
      RECT 119.155 -73.889 119.245 -72.882 ;
      RECT 119.155 -73.365 119.295 -73.195 ;
      RECT 119.155 -72.468 119.245 -71.461 ;
      RECT 119.155 -72.155 119.295 -71.985 ;
      RECT 119.155 -70.659 119.245 -69.652 ;
      RECT 119.155 -70.135 119.295 -69.965 ;
      RECT 119.155 -69.238 119.245 -68.231 ;
      RECT 119.155 -68.925 119.295 -68.755 ;
      RECT 119.155 -67.429 119.245 -66.422 ;
      RECT 119.155 -66.905 119.295 -66.735 ;
      RECT 119.155 -66.008 119.245 -65.001 ;
      RECT 119.155 -65.695 119.295 -65.525 ;
      RECT 119.155 -64.199 119.245 -63.192 ;
      RECT 119.155 -63.675 119.295 -63.505 ;
      RECT 119.155 -62.778 119.245 -61.771 ;
      RECT 119.155 -62.465 119.295 -62.295 ;
      RECT 119.155 -60.969 119.245 -59.962 ;
      RECT 119.155 -60.445 119.295 -60.275 ;
      RECT 119.155 -59.548 119.245 -58.541 ;
      RECT 119.155 -59.235 119.295 -59.065 ;
      RECT 119.155 -57.739 119.245 -56.732 ;
      RECT 119.155 -57.215 119.295 -57.045 ;
      RECT 119.155 -56.318 119.245 -55.311 ;
      RECT 119.155 -56.005 119.295 -55.835 ;
      RECT 119.155 -54.509 119.245 -53.502 ;
      RECT 119.155 -53.985 119.295 -53.815 ;
      RECT 119.155 -53.088 119.245 -52.081 ;
      RECT 119.155 -52.775 119.295 -52.605 ;
      RECT 119.155 -51.279 119.245 -50.272 ;
      RECT 119.155 -50.755 119.295 -50.585 ;
      RECT 119.155 -49.858 119.245 -48.851 ;
      RECT 119.155 -49.545 119.295 -49.375 ;
      RECT 119.155 -48.049 119.245 -47.042 ;
      RECT 119.155 -47.525 119.295 -47.355 ;
      RECT 119.155 -46.628 119.245 -45.621 ;
      RECT 119.155 -46.315 119.295 -46.145 ;
      RECT 119.155 -44.819 119.245 -43.812 ;
      RECT 119.155 -44.295 119.295 -44.125 ;
      RECT 119.155 -43.398 119.245 -42.391 ;
      RECT 119.155 -43.085 119.295 -42.915 ;
      RECT 119.155 -41.589 119.245 -40.582 ;
      RECT 119.155 -41.065 119.295 -40.895 ;
      RECT 119.155 -40.168 119.245 -39.161 ;
      RECT 119.155 -39.855 119.295 -39.685 ;
      RECT 119.155 -38.359 119.245 -37.352 ;
      RECT 119.155 -37.835 119.295 -37.665 ;
      RECT 119.155 -36.938 119.245 -35.931 ;
      RECT 119.155 -36.625 119.295 -36.455 ;
      RECT 119.155 -35.129 119.245 -34.122 ;
      RECT 119.155 -34.605 119.295 -34.435 ;
      RECT 119.155 -33.708 119.245 -32.701 ;
      RECT 119.155 -33.395 119.295 -33.225 ;
      RECT 119.155 -31.899 119.245 -30.892 ;
      RECT 119.155 -31.375 119.295 -31.205 ;
      RECT 119.155 -30.478 119.245 -29.471 ;
      RECT 119.155 -30.165 119.295 -29.995 ;
      RECT 119.155 -28.669 119.245 -27.662 ;
      RECT 119.155 -28.145 119.295 -27.975 ;
      RECT 119.155 -27.248 119.245 -26.241 ;
      RECT 119.155 -26.935 119.295 -26.765 ;
      RECT 119.155 -25.439 119.245 -24.432 ;
      RECT 119.155 -24.915 119.295 -24.745 ;
      RECT 119.155 -24.018 119.245 -23.011 ;
      RECT 119.155 -23.705 119.295 -23.535 ;
      RECT 119.155 -22.209 119.245 -21.202 ;
      RECT 119.155 -21.685 119.295 -21.515 ;
      RECT 119.155 -20.788 119.245 -19.781 ;
      RECT 119.155 -20.475 119.295 -20.305 ;
      RECT 119.155 -18.979 119.245 -17.972 ;
      RECT 119.155 -18.455 119.295 -18.285 ;
      RECT 119.155 -17.558 119.245 -16.551 ;
      RECT 119.155 -17.245 119.295 -17.075 ;
      RECT 119.155 -15.749 119.245 -14.742 ;
      RECT 119.155 -15.225 119.295 -15.055 ;
      RECT 119.155 -14.328 119.245 -13.321 ;
      RECT 119.155 -14.015 119.295 -13.845 ;
      RECT 119.155 -12.519 119.245 -11.512 ;
      RECT 119.155 -11.995 119.295 -11.825 ;
      RECT 119.155 -11.098 119.245 -10.091 ;
      RECT 119.155 -10.785 119.295 -10.615 ;
      RECT 119.155 -9.289 119.245 -8.282 ;
      RECT 119.155 -8.765 119.295 -8.595 ;
      RECT 119.155 -7.868 119.245 -6.861 ;
      RECT 119.155 -7.555 119.295 -7.385 ;
      RECT 119.155 -6.059 119.245 -5.052 ;
      RECT 119.155 -5.535 119.295 -5.365 ;
      RECT 119.155 -4.638 119.245 -3.631 ;
      RECT 119.155 -4.325 119.295 -4.155 ;
      RECT 119.155 -2.829 119.245 -1.822 ;
      RECT 119.155 -2.305 119.295 -2.135 ;
      RECT 119.155 -1.408 119.245 -0.401 ;
      RECT 119.155 -1.095 119.295 -0.925 ;
      RECT 119.155 0.401 119.245 1.408 ;
      RECT 119.155 0.925 119.295 1.095 ;
      RECT 118.485 -111.495 118.655 -111.385 ;
      RECT 115.335 -111.495 118.655 -111.395 ;
      RECT 118.355 -101.538 118.445 -100.53 ;
      RECT 118.305 -100.935 118.445 -100.765 ;
      RECT 118.355 -99.73 118.445 -98.722 ;
      RECT 118.305 -99.495 118.445 -99.325 ;
      RECT 118.355 -98.308 118.445 -97.3 ;
      RECT 118.305 -97.705 118.445 -97.535 ;
      RECT 118.355 -96.5 118.445 -95.492 ;
      RECT 118.305 -96.265 118.445 -96.095 ;
      RECT 118.355 -95.078 118.445 -94.07 ;
      RECT 118.305 -94.475 118.445 -94.305 ;
      RECT 118.355 -93.27 118.445 -92.262 ;
      RECT 118.305 -93.035 118.445 -92.865 ;
      RECT 118.355 -91.848 118.445 -90.84 ;
      RECT 118.305 -91.245 118.445 -91.075 ;
      RECT 118.355 -90.04 118.445 -89.032 ;
      RECT 118.305 -89.805 118.445 -89.635 ;
      RECT 118.355 -88.618 118.445 -87.61 ;
      RECT 118.305 -88.015 118.445 -87.845 ;
      RECT 118.355 -86.81 118.445 -85.802 ;
      RECT 118.305 -86.575 118.445 -86.405 ;
      RECT 118.355 -85.388 118.445 -84.38 ;
      RECT 118.305 -84.785 118.445 -84.615 ;
      RECT 118.355 -83.58 118.445 -82.572 ;
      RECT 118.305 -83.345 118.445 -83.175 ;
      RECT 118.355 -82.158 118.445 -81.15 ;
      RECT 118.305 -81.555 118.445 -81.385 ;
      RECT 118.355 -80.35 118.445 -79.342 ;
      RECT 118.305 -80.115 118.445 -79.945 ;
      RECT 118.355 -78.928 118.445 -77.92 ;
      RECT 118.305 -78.325 118.445 -78.155 ;
      RECT 118.355 -77.12 118.445 -76.112 ;
      RECT 118.305 -76.885 118.445 -76.715 ;
      RECT 118.355 -75.698 118.445 -74.69 ;
      RECT 118.305 -75.095 118.445 -74.925 ;
      RECT 118.355 -73.89 118.445 -72.882 ;
      RECT 118.305 -73.655 118.445 -73.485 ;
      RECT 118.355 -72.468 118.445 -71.46 ;
      RECT 118.305 -71.865 118.445 -71.695 ;
      RECT 118.355 -70.66 118.445 -69.652 ;
      RECT 118.305 -70.425 118.445 -70.255 ;
      RECT 118.355 -69.238 118.445 -68.23 ;
      RECT 118.305 -68.635 118.445 -68.465 ;
      RECT 118.355 -67.43 118.445 -66.422 ;
      RECT 118.305 -67.195 118.445 -67.025 ;
      RECT 118.355 -66.008 118.445 -65 ;
      RECT 118.305 -65.405 118.445 -65.235 ;
      RECT 118.355 -64.2 118.445 -63.192 ;
      RECT 118.305 -63.965 118.445 -63.795 ;
      RECT 118.355 -62.778 118.445 -61.77 ;
      RECT 118.305 -62.175 118.445 -62.005 ;
      RECT 118.355 -60.97 118.445 -59.962 ;
      RECT 118.305 -60.735 118.445 -60.565 ;
      RECT 118.355 -59.548 118.445 -58.54 ;
      RECT 118.305 -58.945 118.445 -58.775 ;
      RECT 118.355 -57.74 118.445 -56.732 ;
      RECT 118.305 -57.505 118.445 -57.335 ;
      RECT 118.355 -56.318 118.445 -55.31 ;
      RECT 118.305 -55.715 118.445 -55.545 ;
      RECT 118.355 -54.51 118.445 -53.502 ;
      RECT 118.305 -54.275 118.445 -54.105 ;
      RECT 118.355 -53.088 118.445 -52.08 ;
      RECT 118.305 -52.485 118.445 -52.315 ;
      RECT 118.355 -51.28 118.445 -50.272 ;
      RECT 118.305 -51.045 118.445 -50.875 ;
      RECT 118.355 -49.858 118.445 -48.85 ;
      RECT 118.305 -49.255 118.445 -49.085 ;
      RECT 118.355 -48.05 118.445 -47.042 ;
      RECT 118.305 -47.815 118.445 -47.645 ;
      RECT 118.355 -46.628 118.445 -45.62 ;
      RECT 118.305 -46.025 118.445 -45.855 ;
      RECT 118.355 -44.82 118.445 -43.812 ;
      RECT 118.305 -44.585 118.445 -44.415 ;
      RECT 118.355 -43.398 118.445 -42.39 ;
      RECT 118.305 -42.795 118.445 -42.625 ;
      RECT 118.355 -41.59 118.445 -40.582 ;
      RECT 118.305 -41.355 118.445 -41.185 ;
      RECT 118.355 -40.168 118.445 -39.16 ;
      RECT 118.305 -39.565 118.445 -39.395 ;
      RECT 118.355 -38.36 118.445 -37.352 ;
      RECT 118.305 -38.125 118.445 -37.955 ;
      RECT 118.355 -36.938 118.445 -35.93 ;
      RECT 118.305 -36.335 118.445 -36.165 ;
      RECT 118.355 -35.13 118.445 -34.122 ;
      RECT 118.305 -34.895 118.445 -34.725 ;
      RECT 118.355 -33.708 118.445 -32.7 ;
      RECT 118.305 -33.105 118.445 -32.935 ;
      RECT 118.355 -31.9 118.445 -30.892 ;
      RECT 118.305 -31.665 118.445 -31.495 ;
      RECT 118.355 -30.478 118.445 -29.47 ;
      RECT 118.305 -29.875 118.445 -29.705 ;
      RECT 118.355 -28.67 118.445 -27.662 ;
      RECT 118.305 -28.435 118.445 -28.265 ;
      RECT 118.355 -27.248 118.445 -26.24 ;
      RECT 118.305 -26.645 118.445 -26.475 ;
      RECT 118.355 -25.44 118.445 -24.432 ;
      RECT 118.305 -25.205 118.445 -25.035 ;
      RECT 118.355 -24.018 118.445 -23.01 ;
      RECT 118.305 -23.415 118.445 -23.245 ;
      RECT 118.355 -22.21 118.445 -21.202 ;
      RECT 118.305 -21.975 118.445 -21.805 ;
      RECT 118.355 -20.788 118.445 -19.78 ;
      RECT 118.305 -20.185 118.445 -20.015 ;
      RECT 118.355 -18.98 118.445 -17.972 ;
      RECT 118.305 -18.745 118.445 -18.575 ;
      RECT 118.355 -17.558 118.445 -16.55 ;
      RECT 118.305 -16.955 118.445 -16.785 ;
      RECT 118.355 -15.75 118.445 -14.742 ;
      RECT 118.305 -15.515 118.445 -15.345 ;
      RECT 118.355 -14.328 118.445 -13.32 ;
      RECT 118.305 -13.725 118.445 -13.555 ;
      RECT 118.355 -12.52 118.445 -11.512 ;
      RECT 118.305 -12.285 118.445 -12.115 ;
      RECT 118.355 -11.098 118.445 -10.09 ;
      RECT 118.305 -10.495 118.445 -10.325 ;
      RECT 118.355 -9.29 118.445 -8.282 ;
      RECT 118.305 -9.055 118.445 -8.885 ;
      RECT 118.355 -7.868 118.445 -6.86 ;
      RECT 118.305 -7.265 118.445 -7.095 ;
      RECT 118.355 -6.06 118.445 -5.052 ;
      RECT 118.305 -5.825 118.445 -5.655 ;
      RECT 118.355 -4.638 118.445 -3.63 ;
      RECT 118.305 -4.035 118.445 -3.865 ;
      RECT 118.355 -2.83 118.445 -1.822 ;
      RECT 118.305 -2.595 118.445 -2.425 ;
      RECT 118.355 -1.408 118.445 -0.4 ;
      RECT 118.305 -0.805 118.445 -0.635 ;
      RECT 118.355 0.4 118.445 1.408 ;
      RECT 118.305 0.635 118.445 0.805 ;
      RECT 117.955 -101.538 118.045 -100.531 ;
      RECT 117.955 -101.225 118.095 -101.055 ;
      RECT 117.955 -99.729 118.045 -98.722 ;
      RECT 117.955 -99.205 118.095 -99.035 ;
      RECT 117.955 -98.308 118.045 -97.301 ;
      RECT 117.955 -97.995 118.095 -97.825 ;
      RECT 117.955 -96.499 118.045 -95.492 ;
      RECT 117.955 -95.975 118.095 -95.805 ;
      RECT 117.955 -95.078 118.045 -94.071 ;
      RECT 117.955 -94.765 118.095 -94.595 ;
      RECT 117.955 -93.269 118.045 -92.262 ;
      RECT 117.955 -92.745 118.095 -92.575 ;
      RECT 117.955 -91.848 118.045 -90.841 ;
      RECT 117.955 -91.535 118.095 -91.365 ;
      RECT 117.955 -90.039 118.045 -89.032 ;
      RECT 117.955 -89.515 118.095 -89.345 ;
      RECT 117.955 -88.618 118.045 -87.611 ;
      RECT 117.955 -88.305 118.095 -88.135 ;
      RECT 117.955 -86.809 118.045 -85.802 ;
      RECT 117.955 -86.285 118.095 -86.115 ;
      RECT 117.955 -85.388 118.045 -84.381 ;
      RECT 117.955 -85.075 118.095 -84.905 ;
      RECT 117.955 -83.579 118.045 -82.572 ;
      RECT 117.955 -83.055 118.095 -82.885 ;
      RECT 117.955 -82.158 118.045 -81.151 ;
      RECT 117.955 -81.845 118.095 -81.675 ;
      RECT 117.955 -80.349 118.045 -79.342 ;
      RECT 117.955 -79.825 118.095 -79.655 ;
      RECT 117.955 -78.928 118.045 -77.921 ;
      RECT 117.955 -78.615 118.095 -78.445 ;
      RECT 117.955 -77.119 118.045 -76.112 ;
      RECT 117.955 -76.595 118.095 -76.425 ;
      RECT 117.955 -75.698 118.045 -74.691 ;
      RECT 117.955 -75.385 118.095 -75.215 ;
      RECT 117.955 -73.889 118.045 -72.882 ;
      RECT 117.955 -73.365 118.095 -73.195 ;
      RECT 117.955 -72.468 118.045 -71.461 ;
      RECT 117.955 -72.155 118.095 -71.985 ;
      RECT 117.955 -70.659 118.045 -69.652 ;
      RECT 117.955 -70.135 118.095 -69.965 ;
      RECT 117.955 -69.238 118.045 -68.231 ;
      RECT 117.955 -68.925 118.095 -68.755 ;
      RECT 117.955 -67.429 118.045 -66.422 ;
      RECT 117.955 -66.905 118.095 -66.735 ;
      RECT 117.955 -66.008 118.045 -65.001 ;
      RECT 117.955 -65.695 118.095 -65.525 ;
      RECT 117.955 -64.199 118.045 -63.192 ;
      RECT 117.955 -63.675 118.095 -63.505 ;
      RECT 117.955 -62.778 118.045 -61.771 ;
      RECT 117.955 -62.465 118.095 -62.295 ;
      RECT 117.955 -60.969 118.045 -59.962 ;
      RECT 117.955 -60.445 118.095 -60.275 ;
      RECT 117.955 -59.548 118.045 -58.541 ;
      RECT 117.955 -59.235 118.095 -59.065 ;
      RECT 117.955 -57.739 118.045 -56.732 ;
      RECT 117.955 -57.215 118.095 -57.045 ;
      RECT 117.955 -56.318 118.045 -55.311 ;
      RECT 117.955 -56.005 118.095 -55.835 ;
      RECT 117.955 -54.509 118.045 -53.502 ;
      RECT 117.955 -53.985 118.095 -53.815 ;
      RECT 117.955 -53.088 118.045 -52.081 ;
      RECT 117.955 -52.775 118.095 -52.605 ;
      RECT 117.955 -51.279 118.045 -50.272 ;
      RECT 117.955 -50.755 118.095 -50.585 ;
      RECT 117.955 -49.858 118.045 -48.851 ;
      RECT 117.955 -49.545 118.095 -49.375 ;
      RECT 117.955 -48.049 118.045 -47.042 ;
      RECT 117.955 -47.525 118.095 -47.355 ;
      RECT 117.955 -46.628 118.045 -45.621 ;
      RECT 117.955 -46.315 118.095 -46.145 ;
      RECT 117.955 -44.819 118.045 -43.812 ;
      RECT 117.955 -44.295 118.095 -44.125 ;
      RECT 117.955 -43.398 118.045 -42.391 ;
      RECT 117.955 -43.085 118.095 -42.915 ;
      RECT 117.955 -41.589 118.045 -40.582 ;
      RECT 117.955 -41.065 118.095 -40.895 ;
      RECT 117.955 -40.168 118.045 -39.161 ;
      RECT 117.955 -39.855 118.095 -39.685 ;
      RECT 117.955 -38.359 118.045 -37.352 ;
      RECT 117.955 -37.835 118.095 -37.665 ;
      RECT 117.955 -36.938 118.045 -35.931 ;
      RECT 117.955 -36.625 118.095 -36.455 ;
      RECT 117.955 -35.129 118.045 -34.122 ;
      RECT 117.955 -34.605 118.095 -34.435 ;
      RECT 117.955 -33.708 118.045 -32.701 ;
      RECT 117.955 -33.395 118.095 -33.225 ;
      RECT 117.955 -31.899 118.045 -30.892 ;
      RECT 117.955 -31.375 118.095 -31.205 ;
      RECT 117.955 -30.478 118.045 -29.471 ;
      RECT 117.955 -30.165 118.095 -29.995 ;
      RECT 117.955 -28.669 118.045 -27.662 ;
      RECT 117.955 -28.145 118.095 -27.975 ;
      RECT 117.955 -27.248 118.045 -26.241 ;
      RECT 117.955 -26.935 118.095 -26.765 ;
      RECT 117.955 -25.439 118.045 -24.432 ;
      RECT 117.955 -24.915 118.095 -24.745 ;
      RECT 117.955 -24.018 118.045 -23.011 ;
      RECT 117.955 -23.705 118.095 -23.535 ;
      RECT 117.955 -22.209 118.045 -21.202 ;
      RECT 117.955 -21.685 118.095 -21.515 ;
      RECT 117.955 -20.788 118.045 -19.781 ;
      RECT 117.955 -20.475 118.095 -20.305 ;
      RECT 117.955 -18.979 118.045 -17.972 ;
      RECT 117.955 -18.455 118.095 -18.285 ;
      RECT 117.955 -17.558 118.045 -16.551 ;
      RECT 117.955 -17.245 118.095 -17.075 ;
      RECT 117.955 -15.749 118.045 -14.742 ;
      RECT 117.955 -15.225 118.095 -15.055 ;
      RECT 117.955 -14.328 118.045 -13.321 ;
      RECT 117.955 -14.015 118.095 -13.845 ;
      RECT 117.955 -12.519 118.045 -11.512 ;
      RECT 117.955 -11.995 118.095 -11.825 ;
      RECT 117.955 -11.098 118.045 -10.091 ;
      RECT 117.955 -10.785 118.095 -10.615 ;
      RECT 117.955 -9.289 118.045 -8.282 ;
      RECT 117.955 -8.765 118.095 -8.595 ;
      RECT 117.955 -7.868 118.045 -6.861 ;
      RECT 117.955 -7.555 118.095 -7.385 ;
      RECT 117.955 -6.059 118.045 -5.052 ;
      RECT 117.955 -5.535 118.095 -5.365 ;
      RECT 117.955 -4.638 118.045 -3.631 ;
      RECT 117.955 -4.325 118.095 -4.155 ;
      RECT 117.955 -2.829 118.045 -1.822 ;
      RECT 117.955 -2.305 118.095 -2.135 ;
      RECT 117.955 -1.408 118.045 -0.401 ;
      RECT 117.955 -1.095 118.095 -0.925 ;
      RECT 117.955 0.401 118.045 1.408 ;
      RECT 117.955 0.925 118.095 1.095 ;
      RECT 116.105 -111.685 117.585 -111.585 ;
      RECT 116.105 -112.055 116.205 -111.585 ;
      RECT 115.91 -114.395 117.485 -114.275 ;
      RECT 117.385 -114.895 117.485 -114.275 ;
      RECT 116.79 -114.895 116.89 -114.275 ;
      RECT 115.91 -114.85 116.01 -114.275 ;
      RECT 117.155 -101.538 117.245 -100.53 ;
      RECT 117.105 -100.935 117.245 -100.765 ;
      RECT 117.155 -99.73 117.245 -98.722 ;
      RECT 117.105 -99.495 117.245 -99.325 ;
      RECT 117.155 -98.308 117.245 -97.3 ;
      RECT 117.105 -97.705 117.245 -97.535 ;
      RECT 117.155 -96.5 117.245 -95.492 ;
      RECT 117.105 -96.265 117.245 -96.095 ;
      RECT 117.155 -95.078 117.245 -94.07 ;
      RECT 117.105 -94.475 117.245 -94.305 ;
      RECT 117.155 -93.27 117.245 -92.262 ;
      RECT 117.105 -93.035 117.245 -92.865 ;
      RECT 117.155 -91.848 117.245 -90.84 ;
      RECT 117.105 -91.245 117.245 -91.075 ;
      RECT 117.155 -90.04 117.245 -89.032 ;
      RECT 117.105 -89.805 117.245 -89.635 ;
      RECT 117.155 -88.618 117.245 -87.61 ;
      RECT 117.105 -88.015 117.245 -87.845 ;
      RECT 117.155 -86.81 117.245 -85.802 ;
      RECT 117.105 -86.575 117.245 -86.405 ;
      RECT 117.155 -85.388 117.245 -84.38 ;
      RECT 117.105 -84.785 117.245 -84.615 ;
      RECT 117.155 -83.58 117.245 -82.572 ;
      RECT 117.105 -83.345 117.245 -83.175 ;
      RECT 117.155 -82.158 117.245 -81.15 ;
      RECT 117.105 -81.555 117.245 -81.385 ;
      RECT 117.155 -80.35 117.245 -79.342 ;
      RECT 117.105 -80.115 117.245 -79.945 ;
      RECT 117.155 -78.928 117.245 -77.92 ;
      RECT 117.105 -78.325 117.245 -78.155 ;
      RECT 117.155 -77.12 117.245 -76.112 ;
      RECT 117.105 -76.885 117.245 -76.715 ;
      RECT 117.155 -75.698 117.245 -74.69 ;
      RECT 117.105 -75.095 117.245 -74.925 ;
      RECT 117.155 -73.89 117.245 -72.882 ;
      RECT 117.105 -73.655 117.245 -73.485 ;
      RECT 117.155 -72.468 117.245 -71.46 ;
      RECT 117.105 -71.865 117.245 -71.695 ;
      RECT 117.155 -70.66 117.245 -69.652 ;
      RECT 117.105 -70.425 117.245 -70.255 ;
      RECT 117.155 -69.238 117.245 -68.23 ;
      RECT 117.105 -68.635 117.245 -68.465 ;
      RECT 117.155 -67.43 117.245 -66.422 ;
      RECT 117.105 -67.195 117.245 -67.025 ;
      RECT 117.155 -66.008 117.245 -65 ;
      RECT 117.105 -65.405 117.245 -65.235 ;
      RECT 117.155 -64.2 117.245 -63.192 ;
      RECT 117.105 -63.965 117.245 -63.795 ;
      RECT 117.155 -62.778 117.245 -61.77 ;
      RECT 117.105 -62.175 117.245 -62.005 ;
      RECT 117.155 -60.97 117.245 -59.962 ;
      RECT 117.105 -60.735 117.245 -60.565 ;
      RECT 117.155 -59.548 117.245 -58.54 ;
      RECT 117.105 -58.945 117.245 -58.775 ;
      RECT 117.155 -57.74 117.245 -56.732 ;
      RECT 117.105 -57.505 117.245 -57.335 ;
      RECT 117.155 -56.318 117.245 -55.31 ;
      RECT 117.105 -55.715 117.245 -55.545 ;
      RECT 117.155 -54.51 117.245 -53.502 ;
      RECT 117.105 -54.275 117.245 -54.105 ;
      RECT 117.155 -53.088 117.245 -52.08 ;
      RECT 117.105 -52.485 117.245 -52.315 ;
      RECT 117.155 -51.28 117.245 -50.272 ;
      RECT 117.105 -51.045 117.245 -50.875 ;
      RECT 117.155 -49.858 117.245 -48.85 ;
      RECT 117.105 -49.255 117.245 -49.085 ;
      RECT 117.155 -48.05 117.245 -47.042 ;
      RECT 117.105 -47.815 117.245 -47.645 ;
      RECT 117.155 -46.628 117.245 -45.62 ;
      RECT 117.105 -46.025 117.245 -45.855 ;
      RECT 117.155 -44.82 117.245 -43.812 ;
      RECT 117.105 -44.585 117.245 -44.415 ;
      RECT 117.155 -43.398 117.245 -42.39 ;
      RECT 117.105 -42.795 117.245 -42.625 ;
      RECT 117.155 -41.59 117.245 -40.582 ;
      RECT 117.105 -41.355 117.245 -41.185 ;
      RECT 117.155 -40.168 117.245 -39.16 ;
      RECT 117.105 -39.565 117.245 -39.395 ;
      RECT 117.155 -38.36 117.245 -37.352 ;
      RECT 117.105 -38.125 117.245 -37.955 ;
      RECT 117.155 -36.938 117.245 -35.93 ;
      RECT 117.105 -36.335 117.245 -36.165 ;
      RECT 117.155 -35.13 117.245 -34.122 ;
      RECT 117.105 -34.895 117.245 -34.725 ;
      RECT 117.155 -33.708 117.245 -32.7 ;
      RECT 117.105 -33.105 117.245 -32.935 ;
      RECT 117.155 -31.9 117.245 -30.892 ;
      RECT 117.105 -31.665 117.245 -31.495 ;
      RECT 117.155 -30.478 117.245 -29.47 ;
      RECT 117.105 -29.875 117.245 -29.705 ;
      RECT 117.155 -28.67 117.245 -27.662 ;
      RECT 117.105 -28.435 117.245 -28.265 ;
      RECT 117.155 -27.248 117.245 -26.24 ;
      RECT 117.105 -26.645 117.245 -26.475 ;
      RECT 117.155 -25.44 117.245 -24.432 ;
      RECT 117.105 -25.205 117.245 -25.035 ;
      RECT 117.155 -24.018 117.245 -23.01 ;
      RECT 117.105 -23.415 117.245 -23.245 ;
      RECT 117.155 -22.21 117.245 -21.202 ;
      RECT 117.105 -21.975 117.245 -21.805 ;
      RECT 117.155 -20.788 117.245 -19.78 ;
      RECT 117.105 -20.185 117.245 -20.015 ;
      RECT 117.155 -18.98 117.245 -17.972 ;
      RECT 117.105 -18.745 117.245 -18.575 ;
      RECT 117.155 -17.558 117.245 -16.55 ;
      RECT 117.105 -16.955 117.245 -16.785 ;
      RECT 117.155 -15.75 117.245 -14.742 ;
      RECT 117.105 -15.515 117.245 -15.345 ;
      RECT 117.155 -14.328 117.245 -13.32 ;
      RECT 117.105 -13.725 117.245 -13.555 ;
      RECT 117.155 -12.52 117.245 -11.512 ;
      RECT 117.105 -12.285 117.245 -12.115 ;
      RECT 117.155 -11.098 117.245 -10.09 ;
      RECT 117.105 -10.495 117.245 -10.325 ;
      RECT 117.155 -9.29 117.245 -8.282 ;
      RECT 117.105 -9.055 117.245 -8.885 ;
      RECT 117.155 -7.868 117.245 -6.86 ;
      RECT 117.105 -7.265 117.245 -7.095 ;
      RECT 117.155 -6.06 117.245 -5.052 ;
      RECT 117.105 -5.825 117.245 -5.655 ;
      RECT 117.155 -4.638 117.245 -3.63 ;
      RECT 117.105 -4.035 117.245 -3.865 ;
      RECT 117.155 -2.83 117.245 -1.822 ;
      RECT 117.105 -2.595 117.245 -2.425 ;
      RECT 117.155 -1.408 117.245 -0.4 ;
      RECT 117.105 -0.805 117.245 -0.635 ;
      RECT 117.155 0.4 117.245 1.408 ;
      RECT 117.105 0.635 117.245 0.805 ;
      RECT 117.03 -114.685 117.205 -114.515 ;
      RECT 117.105 -114.895 117.205 -114.515 ;
      RECT 116.145 -113.555 116.245 -113.09 ;
      RECT 116.51 -113.555 116.61 -113.1 ;
      RECT 116.145 -113.555 116.99 -113.385 ;
      RECT 116.755 -101.538 116.845 -100.531 ;
      RECT 116.755 -101.225 116.895 -101.055 ;
      RECT 116.755 -99.729 116.845 -98.722 ;
      RECT 116.755 -99.205 116.895 -99.035 ;
      RECT 116.755 -98.308 116.845 -97.301 ;
      RECT 116.755 -97.995 116.895 -97.825 ;
      RECT 116.755 -96.499 116.845 -95.492 ;
      RECT 116.755 -95.975 116.895 -95.805 ;
      RECT 116.755 -95.078 116.845 -94.071 ;
      RECT 116.755 -94.765 116.895 -94.595 ;
      RECT 116.755 -93.269 116.845 -92.262 ;
      RECT 116.755 -92.745 116.895 -92.575 ;
      RECT 116.755 -91.848 116.845 -90.841 ;
      RECT 116.755 -91.535 116.895 -91.365 ;
      RECT 116.755 -90.039 116.845 -89.032 ;
      RECT 116.755 -89.515 116.895 -89.345 ;
      RECT 116.755 -88.618 116.845 -87.611 ;
      RECT 116.755 -88.305 116.895 -88.135 ;
      RECT 116.755 -86.809 116.845 -85.802 ;
      RECT 116.755 -86.285 116.895 -86.115 ;
      RECT 116.755 -85.388 116.845 -84.381 ;
      RECT 116.755 -85.075 116.895 -84.905 ;
      RECT 116.755 -83.579 116.845 -82.572 ;
      RECT 116.755 -83.055 116.895 -82.885 ;
      RECT 116.755 -82.158 116.845 -81.151 ;
      RECT 116.755 -81.845 116.895 -81.675 ;
      RECT 116.755 -80.349 116.845 -79.342 ;
      RECT 116.755 -79.825 116.895 -79.655 ;
      RECT 116.755 -78.928 116.845 -77.921 ;
      RECT 116.755 -78.615 116.895 -78.445 ;
      RECT 116.755 -77.119 116.845 -76.112 ;
      RECT 116.755 -76.595 116.895 -76.425 ;
      RECT 116.755 -75.698 116.845 -74.691 ;
      RECT 116.755 -75.385 116.895 -75.215 ;
      RECT 116.755 -73.889 116.845 -72.882 ;
      RECT 116.755 -73.365 116.895 -73.195 ;
      RECT 116.755 -72.468 116.845 -71.461 ;
      RECT 116.755 -72.155 116.895 -71.985 ;
      RECT 116.755 -70.659 116.845 -69.652 ;
      RECT 116.755 -70.135 116.895 -69.965 ;
      RECT 116.755 -69.238 116.845 -68.231 ;
      RECT 116.755 -68.925 116.895 -68.755 ;
      RECT 116.755 -67.429 116.845 -66.422 ;
      RECT 116.755 -66.905 116.895 -66.735 ;
      RECT 116.755 -66.008 116.845 -65.001 ;
      RECT 116.755 -65.695 116.895 -65.525 ;
      RECT 116.755 -64.199 116.845 -63.192 ;
      RECT 116.755 -63.675 116.895 -63.505 ;
      RECT 116.755 -62.778 116.845 -61.771 ;
      RECT 116.755 -62.465 116.895 -62.295 ;
      RECT 116.755 -60.969 116.845 -59.962 ;
      RECT 116.755 -60.445 116.895 -60.275 ;
      RECT 116.755 -59.548 116.845 -58.541 ;
      RECT 116.755 -59.235 116.895 -59.065 ;
      RECT 116.755 -57.739 116.845 -56.732 ;
      RECT 116.755 -57.215 116.895 -57.045 ;
      RECT 116.755 -56.318 116.845 -55.311 ;
      RECT 116.755 -56.005 116.895 -55.835 ;
      RECT 116.755 -54.509 116.845 -53.502 ;
      RECT 116.755 -53.985 116.895 -53.815 ;
      RECT 116.755 -53.088 116.845 -52.081 ;
      RECT 116.755 -52.775 116.895 -52.605 ;
      RECT 116.755 -51.279 116.845 -50.272 ;
      RECT 116.755 -50.755 116.895 -50.585 ;
      RECT 116.755 -49.858 116.845 -48.851 ;
      RECT 116.755 -49.545 116.895 -49.375 ;
      RECT 116.755 -48.049 116.845 -47.042 ;
      RECT 116.755 -47.525 116.895 -47.355 ;
      RECT 116.755 -46.628 116.845 -45.621 ;
      RECT 116.755 -46.315 116.895 -46.145 ;
      RECT 116.755 -44.819 116.845 -43.812 ;
      RECT 116.755 -44.295 116.895 -44.125 ;
      RECT 116.755 -43.398 116.845 -42.391 ;
      RECT 116.755 -43.085 116.895 -42.915 ;
      RECT 116.755 -41.589 116.845 -40.582 ;
      RECT 116.755 -41.065 116.895 -40.895 ;
      RECT 116.755 -40.168 116.845 -39.161 ;
      RECT 116.755 -39.855 116.895 -39.685 ;
      RECT 116.755 -38.359 116.845 -37.352 ;
      RECT 116.755 -37.835 116.895 -37.665 ;
      RECT 116.755 -36.938 116.845 -35.931 ;
      RECT 116.755 -36.625 116.895 -36.455 ;
      RECT 116.755 -35.129 116.845 -34.122 ;
      RECT 116.755 -34.605 116.895 -34.435 ;
      RECT 116.755 -33.708 116.845 -32.701 ;
      RECT 116.755 -33.395 116.895 -33.225 ;
      RECT 116.755 -31.899 116.845 -30.892 ;
      RECT 116.755 -31.375 116.895 -31.205 ;
      RECT 116.755 -30.478 116.845 -29.471 ;
      RECT 116.755 -30.165 116.895 -29.995 ;
      RECT 116.755 -28.669 116.845 -27.662 ;
      RECT 116.755 -28.145 116.895 -27.975 ;
      RECT 116.755 -27.248 116.845 -26.241 ;
      RECT 116.755 -26.935 116.895 -26.765 ;
      RECT 116.755 -25.439 116.845 -24.432 ;
      RECT 116.755 -24.915 116.895 -24.745 ;
      RECT 116.755 -24.018 116.845 -23.011 ;
      RECT 116.755 -23.705 116.895 -23.535 ;
      RECT 116.755 -22.209 116.845 -21.202 ;
      RECT 116.755 -21.685 116.895 -21.515 ;
      RECT 116.755 -20.788 116.845 -19.781 ;
      RECT 116.755 -20.475 116.895 -20.305 ;
      RECT 116.755 -18.979 116.845 -17.972 ;
      RECT 116.755 -18.455 116.895 -18.285 ;
      RECT 116.755 -17.558 116.845 -16.551 ;
      RECT 116.755 -17.245 116.895 -17.075 ;
      RECT 116.755 -15.749 116.845 -14.742 ;
      RECT 116.755 -15.225 116.895 -15.055 ;
      RECT 116.755 -14.328 116.845 -13.321 ;
      RECT 116.755 -14.015 116.895 -13.845 ;
      RECT 116.755 -12.519 116.845 -11.512 ;
      RECT 116.755 -11.995 116.895 -11.825 ;
      RECT 116.755 -11.098 116.845 -10.091 ;
      RECT 116.755 -10.785 116.895 -10.615 ;
      RECT 116.755 -9.289 116.845 -8.282 ;
      RECT 116.755 -8.765 116.895 -8.595 ;
      RECT 116.755 -7.868 116.845 -6.861 ;
      RECT 116.755 -7.555 116.895 -7.385 ;
      RECT 116.755 -6.059 116.845 -5.052 ;
      RECT 116.755 -5.535 116.895 -5.365 ;
      RECT 116.755 -4.638 116.845 -3.631 ;
      RECT 116.755 -4.325 116.895 -4.155 ;
      RECT 116.755 -2.829 116.845 -1.822 ;
      RECT 116.755 -2.305 116.895 -2.135 ;
      RECT 116.755 -1.408 116.845 -0.401 ;
      RECT 116.755 -1.095 116.895 -0.925 ;
      RECT 116.755 0.401 116.845 1.408 ;
      RECT 116.755 0.925 116.895 1.095 ;
      RECT 116.44 -114.685 116.61 -114.515 ;
      RECT 116.51 -114.895 116.61 -114.515 ;
      RECT 115.955 -101.538 116.045 -100.53 ;
      RECT 115.905 -100.935 116.045 -100.765 ;
      RECT 115.955 -99.73 116.045 -98.722 ;
      RECT 115.905 -99.495 116.045 -99.325 ;
      RECT 115.955 -98.308 116.045 -97.3 ;
      RECT 115.905 -97.705 116.045 -97.535 ;
      RECT 115.955 -96.5 116.045 -95.492 ;
      RECT 115.905 -96.265 116.045 -96.095 ;
      RECT 115.955 -95.078 116.045 -94.07 ;
      RECT 115.905 -94.475 116.045 -94.305 ;
      RECT 115.955 -93.27 116.045 -92.262 ;
      RECT 115.905 -93.035 116.045 -92.865 ;
      RECT 115.955 -91.848 116.045 -90.84 ;
      RECT 115.905 -91.245 116.045 -91.075 ;
      RECT 115.955 -90.04 116.045 -89.032 ;
      RECT 115.905 -89.805 116.045 -89.635 ;
      RECT 115.955 -88.618 116.045 -87.61 ;
      RECT 115.905 -88.015 116.045 -87.845 ;
      RECT 115.955 -86.81 116.045 -85.802 ;
      RECT 115.905 -86.575 116.045 -86.405 ;
      RECT 115.955 -85.388 116.045 -84.38 ;
      RECT 115.905 -84.785 116.045 -84.615 ;
      RECT 115.955 -83.58 116.045 -82.572 ;
      RECT 115.905 -83.345 116.045 -83.175 ;
      RECT 115.955 -82.158 116.045 -81.15 ;
      RECT 115.905 -81.555 116.045 -81.385 ;
      RECT 115.955 -80.35 116.045 -79.342 ;
      RECT 115.905 -80.115 116.045 -79.945 ;
      RECT 115.955 -78.928 116.045 -77.92 ;
      RECT 115.905 -78.325 116.045 -78.155 ;
      RECT 115.955 -77.12 116.045 -76.112 ;
      RECT 115.905 -76.885 116.045 -76.715 ;
      RECT 115.955 -75.698 116.045 -74.69 ;
      RECT 115.905 -75.095 116.045 -74.925 ;
      RECT 115.955 -73.89 116.045 -72.882 ;
      RECT 115.905 -73.655 116.045 -73.485 ;
      RECT 115.955 -72.468 116.045 -71.46 ;
      RECT 115.905 -71.865 116.045 -71.695 ;
      RECT 115.955 -70.66 116.045 -69.652 ;
      RECT 115.905 -70.425 116.045 -70.255 ;
      RECT 115.955 -69.238 116.045 -68.23 ;
      RECT 115.905 -68.635 116.045 -68.465 ;
      RECT 115.955 -67.43 116.045 -66.422 ;
      RECT 115.905 -67.195 116.045 -67.025 ;
      RECT 115.955 -66.008 116.045 -65 ;
      RECT 115.905 -65.405 116.045 -65.235 ;
      RECT 115.955 -64.2 116.045 -63.192 ;
      RECT 115.905 -63.965 116.045 -63.795 ;
      RECT 115.955 -62.778 116.045 -61.77 ;
      RECT 115.905 -62.175 116.045 -62.005 ;
      RECT 115.955 -60.97 116.045 -59.962 ;
      RECT 115.905 -60.735 116.045 -60.565 ;
      RECT 115.955 -59.548 116.045 -58.54 ;
      RECT 115.905 -58.945 116.045 -58.775 ;
      RECT 115.955 -57.74 116.045 -56.732 ;
      RECT 115.905 -57.505 116.045 -57.335 ;
      RECT 115.955 -56.318 116.045 -55.31 ;
      RECT 115.905 -55.715 116.045 -55.545 ;
      RECT 115.955 -54.51 116.045 -53.502 ;
      RECT 115.905 -54.275 116.045 -54.105 ;
      RECT 115.955 -53.088 116.045 -52.08 ;
      RECT 115.905 -52.485 116.045 -52.315 ;
      RECT 115.955 -51.28 116.045 -50.272 ;
      RECT 115.905 -51.045 116.045 -50.875 ;
      RECT 115.955 -49.858 116.045 -48.85 ;
      RECT 115.905 -49.255 116.045 -49.085 ;
      RECT 115.955 -48.05 116.045 -47.042 ;
      RECT 115.905 -47.815 116.045 -47.645 ;
      RECT 115.955 -46.628 116.045 -45.62 ;
      RECT 115.905 -46.025 116.045 -45.855 ;
      RECT 115.955 -44.82 116.045 -43.812 ;
      RECT 115.905 -44.585 116.045 -44.415 ;
      RECT 115.955 -43.398 116.045 -42.39 ;
      RECT 115.905 -42.795 116.045 -42.625 ;
      RECT 115.955 -41.59 116.045 -40.582 ;
      RECT 115.905 -41.355 116.045 -41.185 ;
      RECT 115.955 -40.168 116.045 -39.16 ;
      RECT 115.905 -39.565 116.045 -39.395 ;
      RECT 115.955 -38.36 116.045 -37.352 ;
      RECT 115.905 -38.125 116.045 -37.955 ;
      RECT 115.955 -36.938 116.045 -35.93 ;
      RECT 115.905 -36.335 116.045 -36.165 ;
      RECT 115.955 -35.13 116.045 -34.122 ;
      RECT 115.905 -34.895 116.045 -34.725 ;
      RECT 115.955 -33.708 116.045 -32.7 ;
      RECT 115.905 -33.105 116.045 -32.935 ;
      RECT 115.955 -31.9 116.045 -30.892 ;
      RECT 115.905 -31.665 116.045 -31.495 ;
      RECT 115.955 -30.478 116.045 -29.47 ;
      RECT 115.905 -29.875 116.045 -29.705 ;
      RECT 115.955 -28.67 116.045 -27.662 ;
      RECT 115.905 -28.435 116.045 -28.265 ;
      RECT 115.955 -27.248 116.045 -26.24 ;
      RECT 115.905 -26.645 116.045 -26.475 ;
      RECT 115.955 -25.44 116.045 -24.432 ;
      RECT 115.905 -25.205 116.045 -25.035 ;
      RECT 115.955 -24.018 116.045 -23.01 ;
      RECT 115.905 -23.415 116.045 -23.245 ;
      RECT 115.955 -22.21 116.045 -21.202 ;
      RECT 115.905 -21.975 116.045 -21.805 ;
      RECT 115.955 -20.788 116.045 -19.78 ;
      RECT 115.905 -20.185 116.045 -20.015 ;
      RECT 115.955 -18.98 116.045 -17.972 ;
      RECT 115.905 -18.745 116.045 -18.575 ;
      RECT 115.955 -17.558 116.045 -16.55 ;
      RECT 115.905 -16.955 116.045 -16.785 ;
      RECT 115.955 -15.75 116.045 -14.742 ;
      RECT 115.905 -15.515 116.045 -15.345 ;
      RECT 115.955 -14.328 116.045 -13.32 ;
      RECT 115.905 -13.725 116.045 -13.555 ;
      RECT 115.955 -12.52 116.045 -11.512 ;
      RECT 115.905 -12.285 116.045 -12.115 ;
      RECT 115.955 -11.098 116.045 -10.09 ;
      RECT 115.905 -10.495 116.045 -10.325 ;
      RECT 115.955 -9.29 116.045 -8.282 ;
      RECT 115.905 -9.055 116.045 -8.885 ;
      RECT 115.955 -7.868 116.045 -6.86 ;
      RECT 115.905 -7.265 116.045 -7.095 ;
      RECT 115.955 -6.06 116.045 -5.052 ;
      RECT 115.905 -5.825 116.045 -5.655 ;
      RECT 115.955 -4.638 116.045 -3.63 ;
      RECT 115.905 -4.035 116.045 -3.865 ;
      RECT 115.955 -2.83 116.045 -1.822 ;
      RECT 115.905 -2.595 116.045 -2.425 ;
      RECT 115.955 -1.408 116.045 -0.4 ;
      RECT 115.905 -0.805 116.045 -0.635 ;
      RECT 115.955 0.4 116.045 1.408 ;
      RECT 115.905 0.635 116.045 0.805 ;
      RECT 115.555 -101.538 115.645 -100.531 ;
      RECT 115.555 -101.225 115.695 -101.055 ;
      RECT 115.555 -99.729 115.645 -98.722 ;
      RECT 115.555 -99.205 115.695 -99.035 ;
      RECT 115.555 -98.308 115.645 -97.301 ;
      RECT 115.555 -97.995 115.695 -97.825 ;
      RECT 115.555 -96.499 115.645 -95.492 ;
      RECT 115.555 -95.975 115.695 -95.805 ;
      RECT 115.555 -95.078 115.645 -94.071 ;
      RECT 115.555 -94.765 115.695 -94.595 ;
      RECT 115.555 -93.269 115.645 -92.262 ;
      RECT 115.555 -92.745 115.695 -92.575 ;
      RECT 115.555 -91.848 115.645 -90.841 ;
      RECT 115.555 -91.535 115.695 -91.365 ;
      RECT 115.555 -90.039 115.645 -89.032 ;
      RECT 115.555 -89.515 115.695 -89.345 ;
      RECT 115.555 -88.618 115.645 -87.611 ;
      RECT 115.555 -88.305 115.695 -88.135 ;
      RECT 115.555 -86.809 115.645 -85.802 ;
      RECT 115.555 -86.285 115.695 -86.115 ;
      RECT 115.555 -85.388 115.645 -84.381 ;
      RECT 115.555 -85.075 115.695 -84.905 ;
      RECT 115.555 -83.579 115.645 -82.572 ;
      RECT 115.555 -83.055 115.695 -82.885 ;
      RECT 115.555 -82.158 115.645 -81.151 ;
      RECT 115.555 -81.845 115.695 -81.675 ;
      RECT 115.555 -80.349 115.645 -79.342 ;
      RECT 115.555 -79.825 115.695 -79.655 ;
      RECT 115.555 -78.928 115.645 -77.921 ;
      RECT 115.555 -78.615 115.695 -78.445 ;
      RECT 115.555 -77.119 115.645 -76.112 ;
      RECT 115.555 -76.595 115.695 -76.425 ;
      RECT 115.555 -75.698 115.645 -74.691 ;
      RECT 115.555 -75.385 115.695 -75.215 ;
      RECT 115.555 -73.889 115.645 -72.882 ;
      RECT 115.555 -73.365 115.695 -73.195 ;
      RECT 115.555 -72.468 115.645 -71.461 ;
      RECT 115.555 -72.155 115.695 -71.985 ;
      RECT 115.555 -70.659 115.645 -69.652 ;
      RECT 115.555 -70.135 115.695 -69.965 ;
      RECT 115.555 -69.238 115.645 -68.231 ;
      RECT 115.555 -68.925 115.695 -68.755 ;
      RECT 115.555 -67.429 115.645 -66.422 ;
      RECT 115.555 -66.905 115.695 -66.735 ;
      RECT 115.555 -66.008 115.645 -65.001 ;
      RECT 115.555 -65.695 115.695 -65.525 ;
      RECT 115.555 -64.199 115.645 -63.192 ;
      RECT 115.555 -63.675 115.695 -63.505 ;
      RECT 115.555 -62.778 115.645 -61.771 ;
      RECT 115.555 -62.465 115.695 -62.295 ;
      RECT 115.555 -60.969 115.645 -59.962 ;
      RECT 115.555 -60.445 115.695 -60.275 ;
      RECT 115.555 -59.548 115.645 -58.541 ;
      RECT 115.555 -59.235 115.695 -59.065 ;
      RECT 115.555 -57.739 115.645 -56.732 ;
      RECT 115.555 -57.215 115.695 -57.045 ;
      RECT 115.555 -56.318 115.645 -55.311 ;
      RECT 115.555 -56.005 115.695 -55.835 ;
      RECT 115.555 -54.509 115.645 -53.502 ;
      RECT 115.555 -53.985 115.695 -53.815 ;
      RECT 115.555 -53.088 115.645 -52.081 ;
      RECT 115.555 -52.775 115.695 -52.605 ;
      RECT 115.555 -51.279 115.645 -50.272 ;
      RECT 115.555 -50.755 115.695 -50.585 ;
      RECT 115.555 -49.858 115.645 -48.851 ;
      RECT 115.555 -49.545 115.695 -49.375 ;
      RECT 115.555 -48.049 115.645 -47.042 ;
      RECT 115.555 -47.525 115.695 -47.355 ;
      RECT 115.555 -46.628 115.645 -45.621 ;
      RECT 115.555 -46.315 115.695 -46.145 ;
      RECT 115.555 -44.819 115.645 -43.812 ;
      RECT 115.555 -44.295 115.695 -44.125 ;
      RECT 115.555 -43.398 115.645 -42.391 ;
      RECT 115.555 -43.085 115.695 -42.915 ;
      RECT 115.555 -41.589 115.645 -40.582 ;
      RECT 115.555 -41.065 115.695 -40.895 ;
      RECT 115.555 -40.168 115.645 -39.161 ;
      RECT 115.555 -39.855 115.695 -39.685 ;
      RECT 115.555 -38.359 115.645 -37.352 ;
      RECT 115.555 -37.835 115.695 -37.665 ;
      RECT 115.555 -36.938 115.645 -35.931 ;
      RECT 115.555 -36.625 115.695 -36.455 ;
      RECT 115.555 -35.129 115.645 -34.122 ;
      RECT 115.555 -34.605 115.695 -34.435 ;
      RECT 115.555 -33.708 115.645 -32.701 ;
      RECT 115.555 -33.395 115.695 -33.225 ;
      RECT 115.555 -31.899 115.645 -30.892 ;
      RECT 115.555 -31.375 115.695 -31.205 ;
      RECT 115.555 -30.478 115.645 -29.471 ;
      RECT 115.555 -30.165 115.695 -29.995 ;
      RECT 115.555 -28.669 115.645 -27.662 ;
      RECT 115.555 -28.145 115.695 -27.975 ;
      RECT 115.555 -27.248 115.645 -26.241 ;
      RECT 115.555 -26.935 115.695 -26.765 ;
      RECT 115.555 -25.439 115.645 -24.432 ;
      RECT 115.555 -24.915 115.695 -24.745 ;
      RECT 115.555 -24.018 115.645 -23.011 ;
      RECT 115.555 -23.705 115.695 -23.535 ;
      RECT 115.555 -22.209 115.645 -21.202 ;
      RECT 115.555 -21.685 115.695 -21.515 ;
      RECT 115.555 -20.788 115.645 -19.781 ;
      RECT 115.555 -20.475 115.695 -20.305 ;
      RECT 115.555 -18.979 115.645 -17.972 ;
      RECT 115.555 -18.455 115.695 -18.285 ;
      RECT 115.555 -17.558 115.645 -16.551 ;
      RECT 115.555 -17.245 115.695 -17.075 ;
      RECT 115.555 -15.749 115.645 -14.742 ;
      RECT 115.555 -15.225 115.695 -15.055 ;
      RECT 115.555 -14.328 115.645 -13.321 ;
      RECT 115.555 -14.015 115.695 -13.845 ;
      RECT 115.555 -12.519 115.645 -11.512 ;
      RECT 115.555 -11.995 115.695 -11.825 ;
      RECT 115.555 -11.098 115.645 -10.091 ;
      RECT 115.555 -10.785 115.695 -10.615 ;
      RECT 115.555 -9.289 115.645 -8.282 ;
      RECT 115.555 -8.765 115.695 -8.595 ;
      RECT 115.555 -7.868 115.645 -6.861 ;
      RECT 115.555 -7.555 115.695 -7.385 ;
      RECT 115.555 -6.059 115.645 -5.052 ;
      RECT 115.555 -5.535 115.695 -5.365 ;
      RECT 115.555 -4.638 115.645 -3.631 ;
      RECT 115.555 -4.325 115.695 -4.155 ;
      RECT 115.555 -2.829 115.645 -1.822 ;
      RECT 115.555 -2.305 115.695 -2.135 ;
      RECT 115.555 -1.408 115.645 -0.401 ;
      RECT 115.555 -1.095 115.695 -0.925 ;
      RECT 115.555 0.401 115.645 1.408 ;
      RECT 115.555 0.925 115.695 1.095 ;
      RECT 111.385 -108.935 115.165 -108.815 ;
      RECT 112.705 -109.475 112.805 -108.815 ;
      RECT 112.145 -109.475 112.245 -108.815 ;
      RECT 111.585 -109.475 111.685 -108.815 ;
      RECT 114.755 -101.538 114.845 -100.53 ;
      RECT 114.705 -100.935 114.845 -100.765 ;
      RECT 114.755 -99.73 114.845 -98.722 ;
      RECT 114.705 -99.495 114.845 -99.325 ;
      RECT 114.755 -98.308 114.845 -97.3 ;
      RECT 114.705 -97.705 114.845 -97.535 ;
      RECT 114.755 -96.5 114.845 -95.492 ;
      RECT 114.705 -96.265 114.845 -96.095 ;
      RECT 114.755 -95.078 114.845 -94.07 ;
      RECT 114.705 -94.475 114.845 -94.305 ;
      RECT 114.755 -93.27 114.845 -92.262 ;
      RECT 114.705 -93.035 114.845 -92.865 ;
      RECT 114.755 -91.848 114.845 -90.84 ;
      RECT 114.705 -91.245 114.845 -91.075 ;
      RECT 114.755 -90.04 114.845 -89.032 ;
      RECT 114.705 -89.805 114.845 -89.635 ;
      RECT 114.755 -88.618 114.845 -87.61 ;
      RECT 114.705 -88.015 114.845 -87.845 ;
      RECT 114.755 -86.81 114.845 -85.802 ;
      RECT 114.705 -86.575 114.845 -86.405 ;
      RECT 114.755 -85.388 114.845 -84.38 ;
      RECT 114.705 -84.785 114.845 -84.615 ;
      RECT 114.755 -83.58 114.845 -82.572 ;
      RECT 114.705 -83.345 114.845 -83.175 ;
      RECT 114.755 -82.158 114.845 -81.15 ;
      RECT 114.705 -81.555 114.845 -81.385 ;
      RECT 114.755 -80.35 114.845 -79.342 ;
      RECT 114.705 -80.115 114.845 -79.945 ;
      RECT 114.755 -78.928 114.845 -77.92 ;
      RECT 114.705 -78.325 114.845 -78.155 ;
      RECT 114.755 -77.12 114.845 -76.112 ;
      RECT 114.705 -76.885 114.845 -76.715 ;
      RECT 114.755 -75.698 114.845 -74.69 ;
      RECT 114.705 -75.095 114.845 -74.925 ;
      RECT 114.755 -73.89 114.845 -72.882 ;
      RECT 114.705 -73.655 114.845 -73.485 ;
      RECT 114.755 -72.468 114.845 -71.46 ;
      RECT 114.705 -71.865 114.845 -71.695 ;
      RECT 114.755 -70.66 114.845 -69.652 ;
      RECT 114.705 -70.425 114.845 -70.255 ;
      RECT 114.755 -69.238 114.845 -68.23 ;
      RECT 114.705 -68.635 114.845 -68.465 ;
      RECT 114.755 -67.43 114.845 -66.422 ;
      RECT 114.705 -67.195 114.845 -67.025 ;
      RECT 114.755 -66.008 114.845 -65 ;
      RECT 114.705 -65.405 114.845 -65.235 ;
      RECT 114.755 -64.2 114.845 -63.192 ;
      RECT 114.705 -63.965 114.845 -63.795 ;
      RECT 114.755 -62.778 114.845 -61.77 ;
      RECT 114.705 -62.175 114.845 -62.005 ;
      RECT 114.755 -60.97 114.845 -59.962 ;
      RECT 114.705 -60.735 114.845 -60.565 ;
      RECT 114.755 -59.548 114.845 -58.54 ;
      RECT 114.705 -58.945 114.845 -58.775 ;
      RECT 114.755 -57.74 114.845 -56.732 ;
      RECT 114.705 -57.505 114.845 -57.335 ;
      RECT 114.755 -56.318 114.845 -55.31 ;
      RECT 114.705 -55.715 114.845 -55.545 ;
      RECT 114.755 -54.51 114.845 -53.502 ;
      RECT 114.705 -54.275 114.845 -54.105 ;
      RECT 114.755 -53.088 114.845 -52.08 ;
      RECT 114.705 -52.485 114.845 -52.315 ;
      RECT 114.755 -51.28 114.845 -50.272 ;
      RECT 114.705 -51.045 114.845 -50.875 ;
      RECT 114.755 -49.858 114.845 -48.85 ;
      RECT 114.705 -49.255 114.845 -49.085 ;
      RECT 114.755 -48.05 114.845 -47.042 ;
      RECT 114.705 -47.815 114.845 -47.645 ;
      RECT 114.755 -46.628 114.845 -45.62 ;
      RECT 114.705 -46.025 114.845 -45.855 ;
      RECT 114.755 -44.82 114.845 -43.812 ;
      RECT 114.705 -44.585 114.845 -44.415 ;
      RECT 114.755 -43.398 114.845 -42.39 ;
      RECT 114.705 -42.795 114.845 -42.625 ;
      RECT 114.755 -41.59 114.845 -40.582 ;
      RECT 114.705 -41.355 114.845 -41.185 ;
      RECT 114.755 -40.168 114.845 -39.16 ;
      RECT 114.705 -39.565 114.845 -39.395 ;
      RECT 114.755 -38.36 114.845 -37.352 ;
      RECT 114.705 -38.125 114.845 -37.955 ;
      RECT 114.755 -36.938 114.845 -35.93 ;
      RECT 114.705 -36.335 114.845 -36.165 ;
      RECT 114.755 -35.13 114.845 -34.122 ;
      RECT 114.705 -34.895 114.845 -34.725 ;
      RECT 114.755 -33.708 114.845 -32.7 ;
      RECT 114.705 -33.105 114.845 -32.935 ;
      RECT 114.755 -31.9 114.845 -30.892 ;
      RECT 114.705 -31.665 114.845 -31.495 ;
      RECT 114.755 -30.478 114.845 -29.47 ;
      RECT 114.705 -29.875 114.845 -29.705 ;
      RECT 114.755 -28.67 114.845 -27.662 ;
      RECT 114.705 -28.435 114.845 -28.265 ;
      RECT 114.755 -27.248 114.845 -26.24 ;
      RECT 114.705 -26.645 114.845 -26.475 ;
      RECT 114.755 -25.44 114.845 -24.432 ;
      RECT 114.705 -25.205 114.845 -25.035 ;
      RECT 114.755 -24.018 114.845 -23.01 ;
      RECT 114.705 -23.415 114.845 -23.245 ;
      RECT 114.755 -22.21 114.845 -21.202 ;
      RECT 114.705 -21.975 114.845 -21.805 ;
      RECT 114.755 -20.788 114.845 -19.78 ;
      RECT 114.705 -20.185 114.845 -20.015 ;
      RECT 114.755 -18.98 114.845 -17.972 ;
      RECT 114.705 -18.745 114.845 -18.575 ;
      RECT 114.755 -17.558 114.845 -16.55 ;
      RECT 114.705 -16.955 114.845 -16.785 ;
      RECT 114.755 -15.75 114.845 -14.742 ;
      RECT 114.705 -15.515 114.845 -15.345 ;
      RECT 114.755 -14.328 114.845 -13.32 ;
      RECT 114.705 -13.725 114.845 -13.555 ;
      RECT 114.755 -12.52 114.845 -11.512 ;
      RECT 114.705 -12.285 114.845 -12.115 ;
      RECT 114.755 -11.098 114.845 -10.09 ;
      RECT 114.705 -10.495 114.845 -10.325 ;
      RECT 114.755 -9.29 114.845 -8.282 ;
      RECT 114.705 -9.055 114.845 -8.885 ;
      RECT 114.755 -7.868 114.845 -6.86 ;
      RECT 114.705 -7.265 114.845 -7.095 ;
      RECT 114.755 -6.06 114.845 -5.052 ;
      RECT 114.705 -5.825 114.845 -5.655 ;
      RECT 114.755 -4.638 114.845 -3.63 ;
      RECT 114.705 -4.035 114.845 -3.865 ;
      RECT 114.755 -2.83 114.845 -1.822 ;
      RECT 114.705 -2.595 114.845 -2.425 ;
      RECT 114.755 -1.408 114.845 -0.4 ;
      RECT 114.705 -0.805 114.845 -0.635 ;
      RECT 114.755 0.4 114.845 1.408 ;
      RECT 114.705 0.635 114.845 0.805 ;
      RECT 113.325 -111.685 114.805 -111.585 ;
      RECT 113.325 -112.195 113.425 -111.585 ;
      RECT 113.545 -109.15 114.805 -109.05 ;
      RECT 114.705 -109.475 114.805 -109.05 ;
      RECT 114.145 -109.475 114.245 -109.05 ;
      RECT 113.585 -109.475 113.685 -109.05 ;
      RECT 114.355 -101.538 114.445 -100.531 ;
      RECT 114.355 -101.225 114.495 -101.055 ;
      RECT 114.355 -99.729 114.445 -98.722 ;
      RECT 114.355 -99.205 114.495 -99.035 ;
      RECT 114.355 -98.308 114.445 -97.301 ;
      RECT 114.355 -97.995 114.495 -97.825 ;
      RECT 114.355 -96.499 114.445 -95.492 ;
      RECT 114.355 -95.975 114.495 -95.805 ;
      RECT 114.355 -95.078 114.445 -94.071 ;
      RECT 114.355 -94.765 114.495 -94.595 ;
      RECT 114.355 -93.269 114.445 -92.262 ;
      RECT 114.355 -92.745 114.495 -92.575 ;
      RECT 114.355 -91.848 114.445 -90.841 ;
      RECT 114.355 -91.535 114.495 -91.365 ;
      RECT 114.355 -90.039 114.445 -89.032 ;
      RECT 114.355 -89.515 114.495 -89.345 ;
      RECT 114.355 -88.618 114.445 -87.611 ;
      RECT 114.355 -88.305 114.495 -88.135 ;
      RECT 114.355 -86.809 114.445 -85.802 ;
      RECT 114.355 -86.285 114.495 -86.115 ;
      RECT 114.355 -85.388 114.445 -84.381 ;
      RECT 114.355 -85.075 114.495 -84.905 ;
      RECT 114.355 -83.579 114.445 -82.572 ;
      RECT 114.355 -83.055 114.495 -82.885 ;
      RECT 114.355 -82.158 114.445 -81.151 ;
      RECT 114.355 -81.845 114.495 -81.675 ;
      RECT 114.355 -80.349 114.445 -79.342 ;
      RECT 114.355 -79.825 114.495 -79.655 ;
      RECT 114.355 -78.928 114.445 -77.921 ;
      RECT 114.355 -78.615 114.495 -78.445 ;
      RECT 114.355 -77.119 114.445 -76.112 ;
      RECT 114.355 -76.595 114.495 -76.425 ;
      RECT 114.355 -75.698 114.445 -74.691 ;
      RECT 114.355 -75.385 114.495 -75.215 ;
      RECT 114.355 -73.889 114.445 -72.882 ;
      RECT 114.355 -73.365 114.495 -73.195 ;
      RECT 114.355 -72.468 114.445 -71.461 ;
      RECT 114.355 -72.155 114.495 -71.985 ;
      RECT 114.355 -70.659 114.445 -69.652 ;
      RECT 114.355 -70.135 114.495 -69.965 ;
      RECT 114.355 -69.238 114.445 -68.231 ;
      RECT 114.355 -68.925 114.495 -68.755 ;
      RECT 114.355 -67.429 114.445 -66.422 ;
      RECT 114.355 -66.905 114.495 -66.735 ;
      RECT 114.355 -66.008 114.445 -65.001 ;
      RECT 114.355 -65.695 114.495 -65.525 ;
      RECT 114.355 -64.199 114.445 -63.192 ;
      RECT 114.355 -63.675 114.495 -63.505 ;
      RECT 114.355 -62.778 114.445 -61.771 ;
      RECT 114.355 -62.465 114.495 -62.295 ;
      RECT 114.355 -60.969 114.445 -59.962 ;
      RECT 114.355 -60.445 114.495 -60.275 ;
      RECT 114.355 -59.548 114.445 -58.541 ;
      RECT 114.355 -59.235 114.495 -59.065 ;
      RECT 114.355 -57.739 114.445 -56.732 ;
      RECT 114.355 -57.215 114.495 -57.045 ;
      RECT 114.355 -56.318 114.445 -55.311 ;
      RECT 114.355 -56.005 114.495 -55.835 ;
      RECT 114.355 -54.509 114.445 -53.502 ;
      RECT 114.355 -53.985 114.495 -53.815 ;
      RECT 114.355 -53.088 114.445 -52.081 ;
      RECT 114.355 -52.775 114.495 -52.605 ;
      RECT 114.355 -51.279 114.445 -50.272 ;
      RECT 114.355 -50.755 114.495 -50.585 ;
      RECT 114.355 -49.858 114.445 -48.851 ;
      RECT 114.355 -49.545 114.495 -49.375 ;
      RECT 114.355 -48.049 114.445 -47.042 ;
      RECT 114.355 -47.525 114.495 -47.355 ;
      RECT 114.355 -46.628 114.445 -45.621 ;
      RECT 114.355 -46.315 114.495 -46.145 ;
      RECT 114.355 -44.819 114.445 -43.812 ;
      RECT 114.355 -44.295 114.495 -44.125 ;
      RECT 114.355 -43.398 114.445 -42.391 ;
      RECT 114.355 -43.085 114.495 -42.915 ;
      RECT 114.355 -41.589 114.445 -40.582 ;
      RECT 114.355 -41.065 114.495 -40.895 ;
      RECT 114.355 -40.168 114.445 -39.161 ;
      RECT 114.355 -39.855 114.495 -39.685 ;
      RECT 114.355 -38.359 114.445 -37.352 ;
      RECT 114.355 -37.835 114.495 -37.665 ;
      RECT 114.355 -36.938 114.445 -35.931 ;
      RECT 114.355 -36.625 114.495 -36.455 ;
      RECT 114.355 -35.129 114.445 -34.122 ;
      RECT 114.355 -34.605 114.495 -34.435 ;
      RECT 114.355 -33.708 114.445 -32.701 ;
      RECT 114.355 -33.395 114.495 -33.225 ;
      RECT 114.355 -31.899 114.445 -30.892 ;
      RECT 114.355 -31.375 114.495 -31.205 ;
      RECT 114.355 -30.478 114.445 -29.471 ;
      RECT 114.355 -30.165 114.495 -29.995 ;
      RECT 114.355 -28.669 114.445 -27.662 ;
      RECT 114.355 -28.145 114.495 -27.975 ;
      RECT 114.355 -27.248 114.445 -26.241 ;
      RECT 114.355 -26.935 114.495 -26.765 ;
      RECT 114.355 -25.439 114.445 -24.432 ;
      RECT 114.355 -24.915 114.495 -24.745 ;
      RECT 114.355 -24.018 114.445 -23.011 ;
      RECT 114.355 -23.705 114.495 -23.535 ;
      RECT 114.355 -22.209 114.445 -21.202 ;
      RECT 114.355 -21.685 114.495 -21.515 ;
      RECT 114.355 -20.788 114.445 -19.781 ;
      RECT 114.355 -20.475 114.495 -20.305 ;
      RECT 114.355 -18.979 114.445 -17.972 ;
      RECT 114.355 -18.455 114.495 -18.285 ;
      RECT 114.355 -17.558 114.445 -16.551 ;
      RECT 114.355 -17.245 114.495 -17.075 ;
      RECT 114.355 -15.749 114.445 -14.742 ;
      RECT 114.355 -15.225 114.495 -15.055 ;
      RECT 114.355 -14.328 114.445 -13.321 ;
      RECT 114.355 -14.015 114.495 -13.845 ;
      RECT 114.355 -12.519 114.445 -11.512 ;
      RECT 114.355 -11.995 114.495 -11.825 ;
      RECT 114.355 -11.098 114.445 -10.091 ;
      RECT 114.355 -10.785 114.495 -10.615 ;
      RECT 114.355 -9.289 114.445 -8.282 ;
      RECT 114.355 -8.765 114.495 -8.595 ;
      RECT 114.355 -7.868 114.445 -6.861 ;
      RECT 114.355 -7.555 114.495 -7.385 ;
      RECT 114.355 -6.059 114.445 -5.052 ;
      RECT 114.355 -5.535 114.495 -5.365 ;
      RECT 114.355 -4.638 114.445 -3.631 ;
      RECT 114.355 -4.325 114.495 -4.155 ;
      RECT 114.355 -2.829 114.445 -1.822 ;
      RECT 114.355 -2.305 114.495 -2.135 ;
      RECT 114.355 -1.408 114.445 -0.401 ;
      RECT 114.355 -1.095 114.495 -0.925 ;
      RECT 114.355 0.401 114.445 1.408 ;
      RECT 114.355 0.925 114.495 1.095 ;
      RECT 113.685 -111.495 113.855 -111.385 ;
      RECT 110.535 -111.495 113.855 -111.395 ;
      RECT 113.555 -101.538 113.645 -100.53 ;
      RECT 113.505 -100.935 113.645 -100.765 ;
      RECT 113.555 -99.73 113.645 -98.722 ;
      RECT 113.505 -99.495 113.645 -99.325 ;
      RECT 113.555 -98.308 113.645 -97.3 ;
      RECT 113.505 -97.705 113.645 -97.535 ;
      RECT 113.555 -96.5 113.645 -95.492 ;
      RECT 113.505 -96.265 113.645 -96.095 ;
      RECT 113.555 -95.078 113.645 -94.07 ;
      RECT 113.505 -94.475 113.645 -94.305 ;
      RECT 113.555 -93.27 113.645 -92.262 ;
      RECT 113.505 -93.035 113.645 -92.865 ;
      RECT 113.555 -91.848 113.645 -90.84 ;
      RECT 113.505 -91.245 113.645 -91.075 ;
      RECT 113.555 -90.04 113.645 -89.032 ;
      RECT 113.505 -89.805 113.645 -89.635 ;
      RECT 113.555 -88.618 113.645 -87.61 ;
      RECT 113.505 -88.015 113.645 -87.845 ;
      RECT 113.555 -86.81 113.645 -85.802 ;
      RECT 113.505 -86.575 113.645 -86.405 ;
      RECT 113.555 -85.388 113.645 -84.38 ;
      RECT 113.505 -84.785 113.645 -84.615 ;
      RECT 113.555 -83.58 113.645 -82.572 ;
      RECT 113.505 -83.345 113.645 -83.175 ;
      RECT 113.555 -82.158 113.645 -81.15 ;
      RECT 113.505 -81.555 113.645 -81.385 ;
      RECT 113.555 -80.35 113.645 -79.342 ;
      RECT 113.505 -80.115 113.645 -79.945 ;
      RECT 113.555 -78.928 113.645 -77.92 ;
      RECT 113.505 -78.325 113.645 -78.155 ;
      RECT 113.555 -77.12 113.645 -76.112 ;
      RECT 113.505 -76.885 113.645 -76.715 ;
      RECT 113.555 -75.698 113.645 -74.69 ;
      RECT 113.505 -75.095 113.645 -74.925 ;
      RECT 113.555 -73.89 113.645 -72.882 ;
      RECT 113.505 -73.655 113.645 -73.485 ;
      RECT 113.555 -72.468 113.645 -71.46 ;
      RECT 113.505 -71.865 113.645 -71.695 ;
      RECT 113.555 -70.66 113.645 -69.652 ;
      RECT 113.505 -70.425 113.645 -70.255 ;
      RECT 113.555 -69.238 113.645 -68.23 ;
      RECT 113.505 -68.635 113.645 -68.465 ;
      RECT 113.555 -67.43 113.645 -66.422 ;
      RECT 113.505 -67.195 113.645 -67.025 ;
      RECT 113.555 -66.008 113.645 -65 ;
      RECT 113.505 -65.405 113.645 -65.235 ;
      RECT 113.555 -64.2 113.645 -63.192 ;
      RECT 113.505 -63.965 113.645 -63.795 ;
      RECT 113.555 -62.778 113.645 -61.77 ;
      RECT 113.505 -62.175 113.645 -62.005 ;
      RECT 113.555 -60.97 113.645 -59.962 ;
      RECT 113.505 -60.735 113.645 -60.565 ;
      RECT 113.555 -59.548 113.645 -58.54 ;
      RECT 113.505 -58.945 113.645 -58.775 ;
      RECT 113.555 -57.74 113.645 -56.732 ;
      RECT 113.505 -57.505 113.645 -57.335 ;
      RECT 113.555 -56.318 113.645 -55.31 ;
      RECT 113.505 -55.715 113.645 -55.545 ;
      RECT 113.555 -54.51 113.645 -53.502 ;
      RECT 113.505 -54.275 113.645 -54.105 ;
      RECT 113.555 -53.088 113.645 -52.08 ;
      RECT 113.505 -52.485 113.645 -52.315 ;
      RECT 113.555 -51.28 113.645 -50.272 ;
      RECT 113.505 -51.045 113.645 -50.875 ;
      RECT 113.555 -49.858 113.645 -48.85 ;
      RECT 113.505 -49.255 113.645 -49.085 ;
      RECT 113.555 -48.05 113.645 -47.042 ;
      RECT 113.505 -47.815 113.645 -47.645 ;
      RECT 113.555 -46.628 113.645 -45.62 ;
      RECT 113.505 -46.025 113.645 -45.855 ;
      RECT 113.555 -44.82 113.645 -43.812 ;
      RECT 113.505 -44.585 113.645 -44.415 ;
      RECT 113.555 -43.398 113.645 -42.39 ;
      RECT 113.505 -42.795 113.645 -42.625 ;
      RECT 113.555 -41.59 113.645 -40.582 ;
      RECT 113.505 -41.355 113.645 -41.185 ;
      RECT 113.555 -40.168 113.645 -39.16 ;
      RECT 113.505 -39.565 113.645 -39.395 ;
      RECT 113.555 -38.36 113.645 -37.352 ;
      RECT 113.505 -38.125 113.645 -37.955 ;
      RECT 113.555 -36.938 113.645 -35.93 ;
      RECT 113.505 -36.335 113.645 -36.165 ;
      RECT 113.555 -35.13 113.645 -34.122 ;
      RECT 113.505 -34.895 113.645 -34.725 ;
      RECT 113.555 -33.708 113.645 -32.7 ;
      RECT 113.505 -33.105 113.645 -32.935 ;
      RECT 113.555 -31.9 113.645 -30.892 ;
      RECT 113.505 -31.665 113.645 -31.495 ;
      RECT 113.555 -30.478 113.645 -29.47 ;
      RECT 113.505 -29.875 113.645 -29.705 ;
      RECT 113.555 -28.67 113.645 -27.662 ;
      RECT 113.505 -28.435 113.645 -28.265 ;
      RECT 113.555 -27.248 113.645 -26.24 ;
      RECT 113.505 -26.645 113.645 -26.475 ;
      RECT 113.555 -25.44 113.645 -24.432 ;
      RECT 113.505 -25.205 113.645 -25.035 ;
      RECT 113.555 -24.018 113.645 -23.01 ;
      RECT 113.505 -23.415 113.645 -23.245 ;
      RECT 113.555 -22.21 113.645 -21.202 ;
      RECT 113.505 -21.975 113.645 -21.805 ;
      RECT 113.555 -20.788 113.645 -19.78 ;
      RECT 113.505 -20.185 113.645 -20.015 ;
      RECT 113.555 -18.98 113.645 -17.972 ;
      RECT 113.505 -18.745 113.645 -18.575 ;
      RECT 113.555 -17.558 113.645 -16.55 ;
      RECT 113.505 -16.955 113.645 -16.785 ;
      RECT 113.555 -15.75 113.645 -14.742 ;
      RECT 113.505 -15.515 113.645 -15.345 ;
      RECT 113.555 -14.328 113.645 -13.32 ;
      RECT 113.505 -13.725 113.645 -13.555 ;
      RECT 113.555 -12.52 113.645 -11.512 ;
      RECT 113.505 -12.285 113.645 -12.115 ;
      RECT 113.555 -11.098 113.645 -10.09 ;
      RECT 113.505 -10.495 113.645 -10.325 ;
      RECT 113.555 -9.29 113.645 -8.282 ;
      RECT 113.505 -9.055 113.645 -8.885 ;
      RECT 113.555 -7.868 113.645 -6.86 ;
      RECT 113.505 -7.265 113.645 -7.095 ;
      RECT 113.555 -6.06 113.645 -5.052 ;
      RECT 113.505 -5.825 113.645 -5.655 ;
      RECT 113.555 -4.638 113.645 -3.63 ;
      RECT 113.505 -4.035 113.645 -3.865 ;
      RECT 113.555 -2.83 113.645 -1.822 ;
      RECT 113.505 -2.595 113.645 -2.425 ;
      RECT 113.555 -1.408 113.645 -0.4 ;
      RECT 113.505 -0.805 113.645 -0.635 ;
      RECT 113.555 0.4 113.645 1.408 ;
      RECT 113.505 0.635 113.645 0.805 ;
      RECT 113.155 -101.538 113.245 -100.531 ;
      RECT 113.155 -101.225 113.295 -101.055 ;
      RECT 113.155 -99.729 113.245 -98.722 ;
      RECT 113.155 -99.205 113.295 -99.035 ;
      RECT 113.155 -98.308 113.245 -97.301 ;
      RECT 113.155 -97.995 113.295 -97.825 ;
      RECT 113.155 -96.499 113.245 -95.492 ;
      RECT 113.155 -95.975 113.295 -95.805 ;
      RECT 113.155 -95.078 113.245 -94.071 ;
      RECT 113.155 -94.765 113.295 -94.595 ;
      RECT 113.155 -93.269 113.245 -92.262 ;
      RECT 113.155 -92.745 113.295 -92.575 ;
      RECT 113.155 -91.848 113.245 -90.841 ;
      RECT 113.155 -91.535 113.295 -91.365 ;
      RECT 113.155 -90.039 113.245 -89.032 ;
      RECT 113.155 -89.515 113.295 -89.345 ;
      RECT 113.155 -88.618 113.245 -87.611 ;
      RECT 113.155 -88.305 113.295 -88.135 ;
      RECT 113.155 -86.809 113.245 -85.802 ;
      RECT 113.155 -86.285 113.295 -86.115 ;
      RECT 113.155 -85.388 113.245 -84.381 ;
      RECT 113.155 -85.075 113.295 -84.905 ;
      RECT 113.155 -83.579 113.245 -82.572 ;
      RECT 113.155 -83.055 113.295 -82.885 ;
      RECT 113.155 -82.158 113.245 -81.151 ;
      RECT 113.155 -81.845 113.295 -81.675 ;
      RECT 113.155 -80.349 113.245 -79.342 ;
      RECT 113.155 -79.825 113.295 -79.655 ;
      RECT 113.155 -78.928 113.245 -77.921 ;
      RECT 113.155 -78.615 113.295 -78.445 ;
      RECT 113.155 -77.119 113.245 -76.112 ;
      RECT 113.155 -76.595 113.295 -76.425 ;
      RECT 113.155 -75.698 113.245 -74.691 ;
      RECT 113.155 -75.385 113.295 -75.215 ;
      RECT 113.155 -73.889 113.245 -72.882 ;
      RECT 113.155 -73.365 113.295 -73.195 ;
      RECT 113.155 -72.468 113.245 -71.461 ;
      RECT 113.155 -72.155 113.295 -71.985 ;
      RECT 113.155 -70.659 113.245 -69.652 ;
      RECT 113.155 -70.135 113.295 -69.965 ;
      RECT 113.155 -69.238 113.245 -68.231 ;
      RECT 113.155 -68.925 113.295 -68.755 ;
      RECT 113.155 -67.429 113.245 -66.422 ;
      RECT 113.155 -66.905 113.295 -66.735 ;
      RECT 113.155 -66.008 113.245 -65.001 ;
      RECT 113.155 -65.695 113.295 -65.525 ;
      RECT 113.155 -64.199 113.245 -63.192 ;
      RECT 113.155 -63.675 113.295 -63.505 ;
      RECT 113.155 -62.778 113.245 -61.771 ;
      RECT 113.155 -62.465 113.295 -62.295 ;
      RECT 113.155 -60.969 113.245 -59.962 ;
      RECT 113.155 -60.445 113.295 -60.275 ;
      RECT 113.155 -59.548 113.245 -58.541 ;
      RECT 113.155 -59.235 113.295 -59.065 ;
      RECT 113.155 -57.739 113.245 -56.732 ;
      RECT 113.155 -57.215 113.295 -57.045 ;
      RECT 113.155 -56.318 113.245 -55.311 ;
      RECT 113.155 -56.005 113.295 -55.835 ;
      RECT 113.155 -54.509 113.245 -53.502 ;
      RECT 113.155 -53.985 113.295 -53.815 ;
      RECT 113.155 -53.088 113.245 -52.081 ;
      RECT 113.155 -52.775 113.295 -52.605 ;
      RECT 113.155 -51.279 113.245 -50.272 ;
      RECT 113.155 -50.755 113.295 -50.585 ;
      RECT 113.155 -49.858 113.245 -48.851 ;
      RECT 113.155 -49.545 113.295 -49.375 ;
      RECT 113.155 -48.049 113.245 -47.042 ;
      RECT 113.155 -47.525 113.295 -47.355 ;
      RECT 113.155 -46.628 113.245 -45.621 ;
      RECT 113.155 -46.315 113.295 -46.145 ;
      RECT 113.155 -44.819 113.245 -43.812 ;
      RECT 113.155 -44.295 113.295 -44.125 ;
      RECT 113.155 -43.398 113.245 -42.391 ;
      RECT 113.155 -43.085 113.295 -42.915 ;
      RECT 113.155 -41.589 113.245 -40.582 ;
      RECT 113.155 -41.065 113.295 -40.895 ;
      RECT 113.155 -40.168 113.245 -39.161 ;
      RECT 113.155 -39.855 113.295 -39.685 ;
      RECT 113.155 -38.359 113.245 -37.352 ;
      RECT 113.155 -37.835 113.295 -37.665 ;
      RECT 113.155 -36.938 113.245 -35.931 ;
      RECT 113.155 -36.625 113.295 -36.455 ;
      RECT 113.155 -35.129 113.245 -34.122 ;
      RECT 113.155 -34.605 113.295 -34.435 ;
      RECT 113.155 -33.708 113.245 -32.701 ;
      RECT 113.155 -33.395 113.295 -33.225 ;
      RECT 113.155 -31.899 113.245 -30.892 ;
      RECT 113.155 -31.375 113.295 -31.205 ;
      RECT 113.155 -30.478 113.245 -29.471 ;
      RECT 113.155 -30.165 113.295 -29.995 ;
      RECT 113.155 -28.669 113.245 -27.662 ;
      RECT 113.155 -28.145 113.295 -27.975 ;
      RECT 113.155 -27.248 113.245 -26.241 ;
      RECT 113.155 -26.935 113.295 -26.765 ;
      RECT 113.155 -25.439 113.245 -24.432 ;
      RECT 113.155 -24.915 113.295 -24.745 ;
      RECT 113.155 -24.018 113.245 -23.011 ;
      RECT 113.155 -23.705 113.295 -23.535 ;
      RECT 113.155 -22.209 113.245 -21.202 ;
      RECT 113.155 -21.685 113.295 -21.515 ;
      RECT 113.155 -20.788 113.245 -19.781 ;
      RECT 113.155 -20.475 113.295 -20.305 ;
      RECT 113.155 -18.979 113.245 -17.972 ;
      RECT 113.155 -18.455 113.295 -18.285 ;
      RECT 113.155 -17.558 113.245 -16.551 ;
      RECT 113.155 -17.245 113.295 -17.075 ;
      RECT 113.155 -15.749 113.245 -14.742 ;
      RECT 113.155 -15.225 113.295 -15.055 ;
      RECT 113.155 -14.328 113.245 -13.321 ;
      RECT 113.155 -14.015 113.295 -13.845 ;
      RECT 113.155 -12.519 113.245 -11.512 ;
      RECT 113.155 -11.995 113.295 -11.825 ;
      RECT 113.155 -11.098 113.245 -10.091 ;
      RECT 113.155 -10.785 113.295 -10.615 ;
      RECT 113.155 -9.289 113.245 -8.282 ;
      RECT 113.155 -8.765 113.295 -8.595 ;
      RECT 113.155 -7.868 113.245 -6.861 ;
      RECT 113.155 -7.555 113.295 -7.385 ;
      RECT 113.155 -6.059 113.245 -5.052 ;
      RECT 113.155 -5.535 113.295 -5.365 ;
      RECT 113.155 -4.638 113.245 -3.631 ;
      RECT 113.155 -4.325 113.295 -4.155 ;
      RECT 113.155 -2.829 113.245 -1.822 ;
      RECT 113.155 -2.305 113.295 -2.135 ;
      RECT 113.155 -1.408 113.245 -0.401 ;
      RECT 113.155 -1.095 113.295 -0.925 ;
      RECT 113.155 0.401 113.245 1.408 ;
      RECT 113.155 0.925 113.295 1.095 ;
      RECT 111.305 -111.685 112.785 -111.585 ;
      RECT 111.305 -112.055 111.405 -111.585 ;
      RECT 111.11 -114.395 112.685 -114.275 ;
      RECT 112.585 -114.895 112.685 -114.275 ;
      RECT 111.99 -114.895 112.09 -114.275 ;
      RECT 111.11 -114.85 111.21 -114.275 ;
      RECT 112.355 -101.538 112.445 -100.53 ;
      RECT 112.305 -100.935 112.445 -100.765 ;
      RECT 112.355 -99.73 112.445 -98.722 ;
      RECT 112.305 -99.495 112.445 -99.325 ;
      RECT 112.355 -98.308 112.445 -97.3 ;
      RECT 112.305 -97.705 112.445 -97.535 ;
      RECT 112.355 -96.5 112.445 -95.492 ;
      RECT 112.305 -96.265 112.445 -96.095 ;
      RECT 112.355 -95.078 112.445 -94.07 ;
      RECT 112.305 -94.475 112.445 -94.305 ;
      RECT 112.355 -93.27 112.445 -92.262 ;
      RECT 112.305 -93.035 112.445 -92.865 ;
      RECT 112.355 -91.848 112.445 -90.84 ;
      RECT 112.305 -91.245 112.445 -91.075 ;
      RECT 112.355 -90.04 112.445 -89.032 ;
      RECT 112.305 -89.805 112.445 -89.635 ;
      RECT 112.355 -88.618 112.445 -87.61 ;
      RECT 112.305 -88.015 112.445 -87.845 ;
      RECT 112.355 -86.81 112.445 -85.802 ;
      RECT 112.305 -86.575 112.445 -86.405 ;
      RECT 112.355 -85.388 112.445 -84.38 ;
      RECT 112.305 -84.785 112.445 -84.615 ;
      RECT 112.355 -83.58 112.445 -82.572 ;
      RECT 112.305 -83.345 112.445 -83.175 ;
      RECT 112.355 -82.158 112.445 -81.15 ;
      RECT 112.305 -81.555 112.445 -81.385 ;
      RECT 112.355 -80.35 112.445 -79.342 ;
      RECT 112.305 -80.115 112.445 -79.945 ;
      RECT 112.355 -78.928 112.445 -77.92 ;
      RECT 112.305 -78.325 112.445 -78.155 ;
      RECT 112.355 -77.12 112.445 -76.112 ;
      RECT 112.305 -76.885 112.445 -76.715 ;
      RECT 112.355 -75.698 112.445 -74.69 ;
      RECT 112.305 -75.095 112.445 -74.925 ;
      RECT 112.355 -73.89 112.445 -72.882 ;
      RECT 112.305 -73.655 112.445 -73.485 ;
      RECT 112.355 -72.468 112.445 -71.46 ;
      RECT 112.305 -71.865 112.445 -71.695 ;
      RECT 112.355 -70.66 112.445 -69.652 ;
      RECT 112.305 -70.425 112.445 -70.255 ;
      RECT 112.355 -69.238 112.445 -68.23 ;
      RECT 112.305 -68.635 112.445 -68.465 ;
      RECT 112.355 -67.43 112.445 -66.422 ;
      RECT 112.305 -67.195 112.445 -67.025 ;
      RECT 112.355 -66.008 112.445 -65 ;
      RECT 112.305 -65.405 112.445 -65.235 ;
      RECT 112.355 -64.2 112.445 -63.192 ;
      RECT 112.305 -63.965 112.445 -63.795 ;
      RECT 112.355 -62.778 112.445 -61.77 ;
      RECT 112.305 -62.175 112.445 -62.005 ;
      RECT 112.355 -60.97 112.445 -59.962 ;
      RECT 112.305 -60.735 112.445 -60.565 ;
      RECT 112.355 -59.548 112.445 -58.54 ;
      RECT 112.305 -58.945 112.445 -58.775 ;
      RECT 112.355 -57.74 112.445 -56.732 ;
      RECT 112.305 -57.505 112.445 -57.335 ;
      RECT 112.355 -56.318 112.445 -55.31 ;
      RECT 112.305 -55.715 112.445 -55.545 ;
      RECT 112.355 -54.51 112.445 -53.502 ;
      RECT 112.305 -54.275 112.445 -54.105 ;
      RECT 112.355 -53.088 112.445 -52.08 ;
      RECT 112.305 -52.485 112.445 -52.315 ;
      RECT 112.355 -51.28 112.445 -50.272 ;
      RECT 112.305 -51.045 112.445 -50.875 ;
      RECT 112.355 -49.858 112.445 -48.85 ;
      RECT 112.305 -49.255 112.445 -49.085 ;
      RECT 112.355 -48.05 112.445 -47.042 ;
      RECT 112.305 -47.815 112.445 -47.645 ;
      RECT 112.355 -46.628 112.445 -45.62 ;
      RECT 112.305 -46.025 112.445 -45.855 ;
      RECT 112.355 -44.82 112.445 -43.812 ;
      RECT 112.305 -44.585 112.445 -44.415 ;
      RECT 112.355 -43.398 112.445 -42.39 ;
      RECT 112.305 -42.795 112.445 -42.625 ;
      RECT 112.355 -41.59 112.445 -40.582 ;
      RECT 112.305 -41.355 112.445 -41.185 ;
      RECT 112.355 -40.168 112.445 -39.16 ;
      RECT 112.305 -39.565 112.445 -39.395 ;
      RECT 112.355 -38.36 112.445 -37.352 ;
      RECT 112.305 -38.125 112.445 -37.955 ;
      RECT 112.355 -36.938 112.445 -35.93 ;
      RECT 112.305 -36.335 112.445 -36.165 ;
      RECT 112.355 -35.13 112.445 -34.122 ;
      RECT 112.305 -34.895 112.445 -34.725 ;
      RECT 112.355 -33.708 112.445 -32.7 ;
      RECT 112.305 -33.105 112.445 -32.935 ;
      RECT 112.355 -31.9 112.445 -30.892 ;
      RECT 112.305 -31.665 112.445 -31.495 ;
      RECT 112.355 -30.478 112.445 -29.47 ;
      RECT 112.305 -29.875 112.445 -29.705 ;
      RECT 112.355 -28.67 112.445 -27.662 ;
      RECT 112.305 -28.435 112.445 -28.265 ;
      RECT 112.355 -27.248 112.445 -26.24 ;
      RECT 112.305 -26.645 112.445 -26.475 ;
      RECT 112.355 -25.44 112.445 -24.432 ;
      RECT 112.305 -25.205 112.445 -25.035 ;
      RECT 112.355 -24.018 112.445 -23.01 ;
      RECT 112.305 -23.415 112.445 -23.245 ;
      RECT 112.355 -22.21 112.445 -21.202 ;
      RECT 112.305 -21.975 112.445 -21.805 ;
      RECT 112.355 -20.788 112.445 -19.78 ;
      RECT 112.305 -20.185 112.445 -20.015 ;
      RECT 112.355 -18.98 112.445 -17.972 ;
      RECT 112.305 -18.745 112.445 -18.575 ;
      RECT 112.355 -17.558 112.445 -16.55 ;
      RECT 112.305 -16.955 112.445 -16.785 ;
      RECT 112.355 -15.75 112.445 -14.742 ;
      RECT 112.305 -15.515 112.445 -15.345 ;
      RECT 112.355 -14.328 112.445 -13.32 ;
      RECT 112.305 -13.725 112.445 -13.555 ;
      RECT 112.355 -12.52 112.445 -11.512 ;
      RECT 112.305 -12.285 112.445 -12.115 ;
      RECT 112.355 -11.098 112.445 -10.09 ;
      RECT 112.305 -10.495 112.445 -10.325 ;
      RECT 112.355 -9.29 112.445 -8.282 ;
      RECT 112.305 -9.055 112.445 -8.885 ;
      RECT 112.355 -7.868 112.445 -6.86 ;
      RECT 112.305 -7.265 112.445 -7.095 ;
      RECT 112.355 -6.06 112.445 -5.052 ;
      RECT 112.305 -5.825 112.445 -5.655 ;
      RECT 112.355 -4.638 112.445 -3.63 ;
      RECT 112.305 -4.035 112.445 -3.865 ;
      RECT 112.355 -2.83 112.445 -1.822 ;
      RECT 112.305 -2.595 112.445 -2.425 ;
      RECT 112.355 -1.408 112.445 -0.4 ;
      RECT 112.305 -0.805 112.445 -0.635 ;
      RECT 112.355 0.4 112.445 1.408 ;
      RECT 112.305 0.635 112.445 0.805 ;
      RECT 112.23 -114.685 112.405 -114.515 ;
      RECT 112.305 -114.895 112.405 -114.515 ;
      RECT 111.345 -113.555 111.445 -113.09 ;
      RECT 111.71 -113.555 111.81 -113.1 ;
      RECT 111.345 -113.555 112.19 -113.385 ;
      RECT 111.955 -101.538 112.045 -100.531 ;
      RECT 111.955 -101.225 112.095 -101.055 ;
      RECT 111.955 -99.729 112.045 -98.722 ;
      RECT 111.955 -99.205 112.095 -99.035 ;
      RECT 111.955 -98.308 112.045 -97.301 ;
      RECT 111.955 -97.995 112.095 -97.825 ;
      RECT 111.955 -96.499 112.045 -95.492 ;
      RECT 111.955 -95.975 112.095 -95.805 ;
      RECT 111.955 -95.078 112.045 -94.071 ;
      RECT 111.955 -94.765 112.095 -94.595 ;
      RECT 111.955 -93.269 112.045 -92.262 ;
      RECT 111.955 -92.745 112.095 -92.575 ;
      RECT 111.955 -91.848 112.045 -90.841 ;
      RECT 111.955 -91.535 112.095 -91.365 ;
      RECT 111.955 -90.039 112.045 -89.032 ;
      RECT 111.955 -89.515 112.095 -89.345 ;
      RECT 111.955 -88.618 112.045 -87.611 ;
      RECT 111.955 -88.305 112.095 -88.135 ;
      RECT 111.955 -86.809 112.045 -85.802 ;
      RECT 111.955 -86.285 112.095 -86.115 ;
      RECT 111.955 -85.388 112.045 -84.381 ;
      RECT 111.955 -85.075 112.095 -84.905 ;
      RECT 111.955 -83.579 112.045 -82.572 ;
      RECT 111.955 -83.055 112.095 -82.885 ;
      RECT 111.955 -82.158 112.045 -81.151 ;
      RECT 111.955 -81.845 112.095 -81.675 ;
      RECT 111.955 -80.349 112.045 -79.342 ;
      RECT 111.955 -79.825 112.095 -79.655 ;
      RECT 111.955 -78.928 112.045 -77.921 ;
      RECT 111.955 -78.615 112.095 -78.445 ;
      RECT 111.955 -77.119 112.045 -76.112 ;
      RECT 111.955 -76.595 112.095 -76.425 ;
      RECT 111.955 -75.698 112.045 -74.691 ;
      RECT 111.955 -75.385 112.095 -75.215 ;
      RECT 111.955 -73.889 112.045 -72.882 ;
      RECT 111.955 -73.365 112.095 -73.195 ;
      RECT 111.955 -72.468 112.045 -71.461 ;
      RECT 111.955 -72.155 112.095 -71.985 ;
      RECT 111.955 -70.659 112.045 -69.652 ;
      RECT 111.955 -70.135 112.095 -69.965 ;
      RECT 111.955 -69.238 112.045 -68.231 ;
      RECT 111.955 -68.925 112.095 -68.755 ;
      RECT 111.955 -67.429 112.045 -66.422 ;
      RECT 111.955 -66.905 112.095 -66.735 ;
      RECT 111.955 -66.008 112.045 -65.001 ;
      RECT 111.955 -65.695 112.095 -65.525 ;
      RECT 111.955 -64.199 112.045 -63.192 ;
      RECT 111.955 -63.675 112.095 -63.505 ;
      RECT 111.955 -62.778 112.045 -61.771 ;
      RECT 111.955 -62.465 112.095 -62.295 ;
      RECT 111.955 -60.969 112.045 -59.962 ;
      RECT 111.955 -60.445 112.095 -60.275 ;
      RECT 111.955 -59.548 112.045 -58.541 ;
      RECT 111.955 -59.235 112.095 -59.065 ;
      RECT 111.955 -57.739 112.045 -56.732 ;
      RECT 111.955 -57.215 112.095 -57.045 ;
      RECT 111.955 -56.318 112.045 -55.311 ;
      RECT 111.955 -56.005 112.095 -55.835 ;
      RECT 111.955 -54.509 112.045 -53.502 ;
      RECT 111.955 -53.985 112.095 -53.815 ;
      RECT 111.955 -53.088 112.045 -52.081 ;
      RECT 111.955 -52.775 112.095 -52.605 ;
      RECT 111.955 -51.279 112.045 -50.272 ;
      RECT 111.955 -50.755 112.095 -50.585 ;
      RECT 111.955 -49.858 112.045 -48.851 ;
      RECT 111.955 -49.545 112.095 -49.375 ;
      RECT 111.955 -48.049 112.045 -47.042 ;
      RECT 111.955 -47.525 112.095 -47.355 ;
      RECT 111.955 -46.628 112.045 -45.621 ;
      RECT 111.955 -46.315 112.095 -46.145 ;
      RECT 111.955 -44.819 112.045 -43.812 ;
      RECT 111.955 -44.295 112.095 -44.125 ;
      RECT 111.955 -43.398 112.045 -42.391 ;
      RECT 111.955 -43.085 112.095 -42.915 ;
      RECT 111.955 -41.589 112.045 -40.582 ;
      RECT 111.955 -41.065 112.095 -40.895 ;
      RECT 111.955 -40.168 112.045 -39.161 ;
      RECT 111.955 -39.855 112.095 -39.685 ;
      RECT 111.955 -38.359 112.045 -37.352 ;
      RECT 111.955 -37.835 112.095 -37.665 ;
      RECT 111.955 -36.938 112.045 -35.931 ;
      RECT 111.955 -36.625 112.095 -36.455 ;
      RECT 111.955 -35.129 112.045 -34.122 ;
      RECT 111.955 -34.605 112.095 -34.435 ;
      RECT 111.955 -33.708 112.045 -32.701 ;
      RECT 111.955 -33.395 112.095 -33.225 ;
      RECT 111.955 -31.899 112.045 -30.892 ;
      RECT 111.955 -31.375 112.095 -31.205 ;
      RECT 111.955 -30.478 112.045 -29.471 ;
      RECT 111.955 -30.165 112.095 -29.995 ;
      RECT 111.955 -28.669 112.045 -27.662 ;
      RECT 111.955 -28.145 112.095 -27.975 ;
      RECT 111.955 -27.248 112.045 -26.241 ;
      RECT 111.955 -26.935 112.095 -26.765 ;
      RECT 111.955 -25.439 112.045 -24.432 ;
      RECT 111.955 -24.915 112.095 -24.745 ;
      RECT 111.955 -24.018 112.045 -23.011 ;
      RECT 111.955 -23.705 112.095 -23.535 ;
      RECT 111.955 -22.209 112.045 -21.202 ;
      RECT 111.955 -21.685 112.095 -21.515 ;
      RECT 111.955 -20.788 112.045 -19.781 ;
      RECT 111.955 -20.475 112.095 -20.305 ;
      RECT 111.955 -18.979 112.045 -17.972 ;
      RECT 111.955 -18.455 112.095 -18.285 ;
      RECT 111.955 -17.558 112.045 -16.551 ;
      RECT 111.955 -17.245 112.095 -17.075 ;
      RECT 111.955 -15.749 112.045 -14.742 ;
      RECT 111.955 -15.225 112.095 -15.055 ;
      RECT 111.955 -14.328 112.045 -13.321 ;
      RECT 111.955 -14.015 112.095 -13.845 ;
      RECT 111.955 -12.519 112.045 -11.512 ;
      RECT 111.955 -11.995 112.095 -11.825 ;
      RECT 111.955 -11.098 112.045 -10.091 ;
      RECT 111.955 -10.785 112.095 -10.615 ;
      RECT 111.955 -9.289 112.045 -8.282 ;
      RECT 111.955 -8.765 112.095 -8.595 ;
      RECT 111.955 -7.868 112.045 -6.861 ;
      RECT 111.955 -7.555 112.095 -7.385 ;
      RECT 111.955 -6.059 112.045 -5.052 ;
      RECT 111.955 -5.535 112.095 -5.365 ;
      RECT 111.955 -4.638 112.045 -3.631 ;
      RECT 111.955 -4.325 112.095 -4.155 ;
      RECT 111.955 -2.829 112.045 -1.822 ;
      RECT 111.955 -2.305 112.095 -2.135 ;
      RECT 111.955 -1.408 112.045 -0.401 ;
      RECT 111.955 -1.095 112.095 -0.925 ;
      RECT 111.955 0.401 112.045 1.408 ;
      RECT 111.955 0.925 112.095 1.095 ;
      RECT 111.64 -114.685 111.81 -114.515 ;
      RECT 111.71 -114.895 111.81 -114.515 ;
      RECT 111.155 -101.538 111.245 -100.53 ;
      RECT 111.105 -100.935 111.245 -100.765 ;
      RECT 111.155 -99.73 111.245 -98.722 ;
      RECT 111.105 -99.495 111.245 -99.325 ;
      RECT 111.155 -98.308 111.245 -97.3 ;
      RECT 111.105 -97.705 111.245 -97.535 ;
      RECT 111.155 -96.5 111.245 -95.492 ;
      RECT 111.105 -96.265 111.245 -96.095 ;
      RECT 111.155 -95.078 111.245 -94.07 ;
      RECT 111.105 -94.475 111.245 -94.305 ;
      RECT 111.155 -93.27 111.245 -92.262 ;
      RECT 111.105 -93.035 111.245 -92.865 ;
      RECT 111.155 -91.848 111.245 -90.84 ;
      RECT 111.105 -91.245 111.245 -91.075 ;
      RECT 111.155 -90.04 111.245 -89.032 ;
      RECT 111.105 -89.805 111.245 -89.635 ;
      RECT 111.155 -88.618 111.245 -87.61 ;
      RECT 111.105 -88.015 111.245 -87.845 ;
      RECT 111.155 -86.81 111.245 -85.802 ;
      RECT 111.105 -86.575 111.245 -86.405 ;
      RECT 111.155 -85.388 111.245 -84.38 ;
      RECT 111.105 -84.785 111.245 -84.615 ;
      RECT 111.155 -83.58 111.245 -82.572 ;
      RECT 111.105 -83.345 111.245 -83.175 ;
      RECT 111.155 -82.158 111.245 -81.15 ;
      RECT 111.105 -81.555 111.245 -81.385 ;
      RECT 111.155 -80.35 111.245 -79.342 ;
      RECT 111.105 -80.115 111.245 -79.945 ;
      RECT 111.155 -78.928 111.245 -77.92 ;
      RECT 111.105 -78.325 111.245 -78.155 ;
      RECT 111.155 -77.12 111.245 -76.112 ;
      RECT 111.105 -76.885 111.245 -76.715 ;
      RECT 111.155 -75.698 111.245 -74.69 ;
      RECT 111.105 -75.095 111.245 -74.925 ;
      RECT 111.155 -73.89 111.245 -72.882 ;
      RECT 111.105 -73.655 111.245 -73.485 ;
      RECT 111.155 -72.468 111.245 -71.46 ;
      RECT 111.105 -71.865 111.245 -71.695 ;
      RECT 111.155 -70.66 111.245 -69.652 ;
      RECT 111.105 -70.425 111.245 -70.255 ;
      RECT 111.155 -69.238 111.245 -68.23 ;
      RECT 111.105 -68.635 111.245 -68.465 ;
      RECT 111.155 -67.43 111.245 -66.422 ;
      RECT 111.105 -67.195 111.245 -67.025 ;
      RECT 111.155 -66.008 111.245 -65 ;
      RECT 111.105 -65.405 111.245 -65.235 ;
      RECT 111.155 -64.2 111.245 -63.192 ;
      RECT 111.105 -63.965 111.245 -63.795 ;
      RECT 111.155 -62.778 111.245 -61.77 ;
      RECT 111.105 -62.175 111.245 -62.005 ;
      RECT 111.155 -60.97 111.245 -59.962 ;
      RECT 111.105 -60.735 111.245 -60.565 ;
      RECT 111.155 -59.548 111.245 -58.54 ;
      RECT 111.105 -58.945 111.245 -58.775 ;
      RECT 111.155 -57.74 111.245 -56.732 ;
      RECT 111.105 -57.505 111.245 -57.335 ;
      RECT 111.155 -56.318 111.245 -55.31 ;
      RECT 111.105 -55.715 111.245 -55.545 ;
      RECT 111.155 -54.51 111.245 -53.502 ;
      RECT 111.105 -54.275 111.245 -54.105 ;
      RECT 111.155 -53.088 111.245 -52.08 ;
      RECT 111.105 -52.485 111.245 -52.315 ;
      RECT 111.155 -51.28 111.245 -50.272 ;
      RECT 111.105 -51.045 111.245 -50.875 ;
      RECT 111.155 -49.858 111.245 -48.85 ;
      RECT 111.105 -49.255 111.245 -49.085 ;
      RECT 111.155 -48.05 111.245 -47.042 ;
      RECT 111.105 -47.815 111.245 -47.645 ;
      RECT 111.155 -46.628 111.245 -45.62 ;
      RECT 111.105 -46.025 111.245 -45.855 ;
      RECT 111.155 -44.82 111.245 -43.812 ;
      RECT 111.105 -44.585 111.245 -44.415 ;
      RECT 111.155 -43.398 111.245 -42.39 ;
      RECT 111.105 -42.795 111.245 -42.625 ;
      RECT 111.155 -41.59 111.245 -40.582 ;
      RECT 111.105 -41.355 111.245 -41.185 ;
      RECT 111.155 -40.168 111.245 -39.16 ;
      RECT 111.105 -39.565 111.245 -39.395 ;
      RECT 111.155 -38.36 111.245 -37.352 ;
      RECT 111.105 -38.125 111.245 -37.955 ;
      RECT 111.155 -36.938 111.245 -35.93 ;
      RECT 111.105 -36.335 111.245 -36.165 ;
      RECT 111.155 -35.13 111.245 -34.122 ;
      RECT 111.105 -34.895 111.245 -34.725 ;
      RECT 111.155 -33.708 111.245 -32.7 ;
      RECT 111.105 -33.105 111.245 -32.935 ;
      RECT 111.155 -31.9 111.245 -30.892 ;
      RECT 111.105 -31.665 111.245 -31.495 ;
      RECT 111.155 -30.478 111.245 -29.47 ;
      RECT 111.105 -29.875 111.245 -29.705 ;
      RECT 111.155 -28.67 111.245 -27.662 ;
      RECT 111.105 -28.435 111.245 -28.265 ;
      RECT 111.155 -27.248 111.245 -26.24 ;
      RECT 111.105 -26.645 111.245 -26.475 ;
      RECT 111.155 -25.44 111.245 -24.432 ;
      RECT 111.105 -25.205 111.245 -25.035 ;
      RECT 111.155 -24.018 111.245 -23.01 ;
      RECT 111.105 -23.415 111.245 -23.245 ;
      RECT 111.155 -22.21 111.245 -21.202 ;
      RECT 111.105 -21.975 111.245 -21.805 ;
      RECT 111.155 -20.788 111.245 -19.78 ;
      RECT 111.105 -20.185 111.245 -20.015 ;
      RECT 111.155 -18.98 111.245 -17.972 ;
      RECT 111.105 -18.745 111.245 -18.575 ;
      RECT 111.155 -17.558 111.245 -16.55 ;
      RECT 111.105 -16.955 111.245 -16.785 ;
      RECT 111.155 -15.75 111.245 -14.742 ;
      RECT 111.105 -15.515 111.245 -15.345 ;
      RECT 111.155 -14.328 111.245 -13.32 ;
      RECT 111.105 -13.725 111.245 -13.555 ;
      RECT 111.155 -12.52 111.245 -11.512 ;
      RECT 111.105 -12.285 111.245 -12.115 ;
      RECT 111.155 -11.098 111.245 -10.09 ;
      RECT 111.105 -10.495 111.245 -10.325 ;
      RECT 111.155 -9.29 111.245 -8.282 ;
      RECT 111.105 -9.055 111.245 -8.885 ;
      RECT 111.155 -7.868 111.245 -6.86 ;
      RECT 111.105 -7.265 111.245 -7.095 ;
      RECT 111.155 -6.06 111.245 -5.052 ;
      RECT 111.105 -5.825 111.245 -5.655 ;
      RECT 111.155 -4.638 111.245 -3.63 ;
      RECT 111.105 -4.035 111.245 -3.865 ;
      RECT 111.155 -2.83 111.245 -1.822 ;
      RECT 111.105 -2.595 111.245 -2.425 ;
      RECT 111.155 -1.408 111.245 -0.4 ;
      RECT 111.105 -0.805 111.245 -0.635 ;
      RECT 111.155 0.4 111.245 1.408 ;
      RECT 111.105 0.635 111.245 0.805 ;
      RECT 110.755 -101.538 110.845 -100.531 ;
      RECT 110.755 -101.225 110.895 -101.055 ;
      RECT 110.755 -99.729 110.845 -98.722 ;
      RECT 110.755 -99.205 110.895 -99.035 ;
      RECT 110.755 -98.308 110.845 -97.301 ;
      RECT 110.755 -97.995 110.895 -97.825 ;
      RECT 110.755 -96.499 110.845 -95.492 ;
      RECT 110.755 -95.975 110.895 -95.805 ;
      RECT 110.755 -95.078 110.845 -94.071 ;
      RECT 110.755 -94.765 110.895 -94.595 ;
      RECT 110.755 -93.269 110.845 -92.262 ;
      RECT 110.755 -92.745 110.895 -92.575 ;
      RECT 110.755 -91.848 110.845 -90.841 ;
      RECT 110.755 -91.535 110.895 -91.365 ;
      RECT 110.755 -90.039 110.845 -89.032 ;
      RECT 110.755 -89.515 110.895 -89.345 ;
      RECT 110.755 -88.618 110.845 -87.611 ;
      RECT 110.755 -88.305 110.895 -88.135 ;
      RECT 110.755 -86.809 110.845 -85.802 ;
      RECT 110.755 -86.285 110.895 -86.115 ;
      RECT 110.755 -85.388 110.845 -84.381 ;
      RECT 110.755 -85.075 110.895 -84.905 ;
      RECT 110.755 -83.579 110.845 -82.572 ;
      RECT 110.755 -83.055 110.895 -82.885 ;
      RECT 110.755 -82.158 110.845 -81.151 ;
      RECT 110.755 -81.845 110.895 -81.675 ;
      RECT 110.755 -80.349 110.845 -79.342 ;
      RECT 110.755 -79.825 110.895 -79.655 ;
      RECT 110.755 -78.928 110.845 -77.921 ;
      RECT 110.755 -78.615 110.895 -78.445 ;
      RECT 110.755 -77.119 110.845 -76.112 ;
      RECT 110.755 -76.595 110.895 -76.425 ;
      RECT 110.755 -75.698 110.845 -74.691 ;
      RECT 110.755 -75.385 110.895 -75.215 ;
      RECT 110.755 -73.889 110.845 -72.882 ;
      RECT 110.755 -73.365 110.895 -73.195 ;
      RECT 110.755 -72.468 110.845 -71.461 ;
      RECT 110.755 -72.155 110.895 -71.985 ;
      RECT 110.755 -70.659 110.845 -69.652 ;
      RECT 110.755 -70.135 110.895 -69.965 ;
      RECT 110.755 -69.238 110.845 -68.231 ;
      RECT 110.755 -68.925 110.895 -68.755 ;
      RECT 110.755 -67.429 110.845 -66.422 ;
      RECT 110.755 -66.905 110.895 -66.735 ;
      RECT 110.755 -66.008 110.845 -65.001 ;
      RECT 110.755 -65.695 110.895 -65.525 ;
      RECT 110.755 -64.199 110.845 -63.192 ;
      RECT 110.755 -63.675 110.895 -63.505 ;
      RECT 110.755 -62.778 110.845 -61.771 ;
      RECT 110.755 -62.465 110.895 -62.295 ;
      RECT 110.755 -60.969 110.845 -59.962 ;
      RECT 110.755 -60.445 110.895 -60.275 ;
      RECT 110.755 -59.548 110.845 -58.541 ;
      RECT 110.755 -59.235 110.895 -59.065 ;
      RECT 110.755 -57.739 110.845 -56.732 ;
      RECT 110.755 -57.215 110.895 -57.045 ;
      RECT 110.755 -56.318 110.845 -55.311 ;
      RECT 110.755 -56.005 110.895 -55.835 ;
      RECT 110.755 -54.509 110.845 -53.502 ;
      RECT 110.755 -53.985 110.895 -53.815 ;
      RECT 110.755 -53.088 110.845 -52.081 ;
      RECT 110.755 -52.775 110.895 -52.605 ;
      RECT 110.755 -51.279 110.845 -50.272 ;
      RECT 110.755 -50.755 110.895 -50.585 ;
      RECT 110.755 -49.858 110.845 -48.851 ;
      RECT 110.755 -49.545 110.895 -49.375 ;
      RECT 110.755 -48.049 110.845 -47.042 ;
      RECT 110.755 -47.525 110.895 -47.355 ;
      RECT 110.755 -46.628 110.845 -45.621 ;
      RECT 110.755 -46.315 110.895 -46.145 ;
      RECT 110.755 -44.819 110.845 -43.812 ;
      RECT 110.755 -44.295 110.895 -44.125 ;
      RECT 110.755 -43.398 110.845 -42.391 ;
      RECT 110.755 -43.085 110.895 -42.915 ;
      RECT 110.755 -41.589 110.845 -40.582 ;
      RECT 110.755 -41.065 110.895 -40.895 ;
      RECT 110.755 -40.168 110.845 -39.161 ;
      RECT 110.755 -39.855 110.895 -39.685 ;
      RECT 110.755 -38.359 110.845 -37.352 ;
      RECT 110.755 -37.835 110.895 -37.665 ;
      RECT 110.755 -36.938 110.845 -35.931 ;
      RECT 110.755 -36.625 110.895 -36.455 ;
      RECT 110.755 -35.129 110.845 -34.122 ;
      RECT 110.755 -34.605 110.895 -34.435 ;
      RECT 110.755 -33.708 110.845 -32.701 ;
      RECT 110.755 -33.395 110.895 -33.225 ;
      RECT 110.755 -31.899 110.845 -30.892 ;
      RECT 110.755 -31.375 110.895 -31.205 ;
      RECT 110.755 -30.478 110.845 -29.471 ;
      RECT 110.755 -30.165 110.895 -29.995 ;
      RECT 110.755 -28.669 110.845 -27.662 ;
      RECT 110.755 -28.145 110.895 -27.975 ;
      RECT 110.755 -27.248 110.845 -26.241 ;
      RECT 110.755 -26.935 110.895 -26.765 ;
      RECT 110.755 -25.439 110.845 -24.432 ;
      RECT 110.755 -24.915 110.895 -24.745 ;
      RECT 110.755 -24.018 110.845 -23.011 ;
      RECT 110.755 -23.705 110.895 -23.535 ;
      RECT 110.755 -22.209 110.845 -21.202 ;
      RECT 110.755 -21.685 110.895 -21.515 ;
      RECT 110.755 -20.788 110.845 -19.781 ;
      RECT 110.755 -20.475 110.895 -20.305 ;
      RECT 110.755 -18.979 110.845 -17.972 ;
      RECT 110.755 -18.455 110.895 -18.285 ;
      RECT 110.755 -17.558 110.845 -16.551 ;
      RECT 110.755 -17.245 110.895 -17.075 ;
      RECT 110.755 -15.749 110.845 -14.742 ;
      RECT 110.755 -15.225 110.895 -15.055 ;
      RECT 110.755 -14.328 110.845 -13.321 ;
      RECT 110.755 -14.015 110.895 -13.845 ;
      RECT 110.755 -12.519 110.845 -11.512 ;
      RECT 110.755 -11.995 110.895 -11.825 ;
      RECT 110.755 -11.098 110.845 -10.091 ;
      RECT 110.755 -10.785 110.895 -10.615 ;
      RECT 110.755 -9.289 110.845 -8.282 ;
      RECT 110.755 -8.765 110.895 -8.595 ;
      RECT 110.755 -7.868 110.845 -6.861 ;
      RECT 110.755 -7.555 110.895 -7.385 ;
      RECT 110.755 -6.059 110.845 -5.052 ;
      RECT 110.755 -5.535 110.895 -5.365 ;
      RECT 110.755 -4.638 110.845 -3.631 ;
      RECT 110.755 -4.325 110.895 -4.155 ;
      RECT 110.755 -2.829 110.845 -1.822 ;
      RECT 110.755 -2.305 110.895 -2.135 ;
      RECT 110.755 -1.408 110.845 -0.401 ;
      RECT 110.755 -1.095 110.895 -0.925 ;
      RECT 110.755 0.401 110.845 1.408 ;
      RECT 110.755 0.925 110.895 1.095 ;
      RECT 106.585 -108.935 110.365 -108.815 ;
      RECT 107.905 -109.475 108.005 -108.815 ;
      RECT 107.345 -109.475 107.445 -108.815 ;
      RECT 106.785 -109.475 106.885 -108.815 ;
      RECT 109.955 -101.538 110.045 -100.53 ;
      RECT 109.905 -100.935 110.045 -100.765 ;
      RECT 109.955 -99.73 110.045 -98.722 ;
      RECT 109.905 -99.495 110.045 -99.325 ;
      RECT 109.955 -98.308 110.045 -97.3 ;
      RECT 109.905 -97.705 110.045 -97.535 ;
      RECT 109.955 -96.5 110.045 -95.492 ;
      RECT 109.905 -96.265 110.045 -96.095 ;
      RECT 109.955 -95.078 110.045 -94.07 ;
      RECT 109.905 -94.475 110.045 -94.305 ;
      RECT 109.955 -93.27 110.045 -92.262 ;
      RECT 109.905 -93.035 110.045 -92.865 ;
      RECT 109.955 -91.848 110.045 -90.84 ;
      RECT 109.905 -91.245 110.045 -91.075 ;
      RECT 109.955 -90.04 110.045 -89.032 ;
      RECT 109.905 -89.805 110.045 -89.635 ;
      RECT 109.955 -88.618 110.045 -87.61 ;
      RECT 109.905 -88.015 110.045 -87.845 ;
      RECT 109.955 -86.81 110.045 -85.802 ;
      RECT 109.905 -86.575 110.045 -86.405 ;
      RECT 109.955 -85.388 110.045 -84.38 ;
      RECT 109.905 -84.785 110.045 -84.615 ;
      RECT 109.955 -83.58 110.045 -82.572 ;
      RECT 109.905 -83.345 110.045 -83.175 ;
      RECT 109.955 -82.158 110.045 -81.15 ;
      RECT 109.905 -81.555 110.045 -81.385 ;
      RECT 109.955 -80.35 110.045 -79.342 ;
      RECT 109.905 -80.115 110.045 -79.945 ;
      RECT 109.955 -78.928 110.045 -77.92 ;
      RECT 109.905 -78.325 110.045 -78.155 ;
      RECT 109.955 -77.12 110.045 -76.112 ;
      RECT 109.905 -76.885 110.045 -76.715 ;
      RECT 109.955 -75.698 110.045 -74.69 ;
      RECT 109.905 -75.095 110.045 -74.925 ;
      RECT 109.955 -73.89 110.045 -72.882 ;
      RECT 109.905 -73.655 110.045 -73.485 ;
      RECT 109.955 -72.468 110.045 -71.46 ;
      RECT 109.905 -71.865 110.045 -71.695 ;
      RECT 109.955 -70.66 110.045 -69.652 ;
      RECT 109.905 -70.425 110.045 -70.255 ;
      RECT 109.955 -69.238 110.045 -68.23 ;
      RECT 109.905 -68.635 110.045 -68.465 ;
      RECT 109.955 -67.43 110.045 -66.422 ;
      RECT 109.905 -67.195 110.045 -67.025 ;
      RECT 109.955 -66.008 110.045 -65 ;
      RECT 109.905 -65.405 110.045 -65.235 ;
      RECT 109.955 -64.2 110.045 -63.192 ;
      RECT 109.905 -63.965 110.045 -63.795 ;
      RECT 109.955 -62.778 110.045 -61.77 ;
      RECT 109.905 -62.175 110.045 -62.005 ;
      RECT 109.955 -60.97 110.045 -59.962 ;
      RECT 109.905 -60.735 110.045 -60.565 ;
      RECT 109.955 -59.548 110.045 -58.54 ;
      RECT 109.905 -58.945 110.045 -58.775 ;
      RECT 109.955 -57.74 110.045 -56.732 ;
      RECT 109.905 -57.505 110.045 -57.335 ;
      RECT 109.955 -56.318 110.045 -55.31 ;
      RECT 109.905 -55.715 110.045 -55.545 ;
      RECT 109.955 -54.51 110.045 -53.502 ;
      RECT 109.905 -54.275 110.045 -54.105 ;
      RECT 109.955 -53.088 110.045 -52.08 ;
      RECT 109.905 -52.485 110.045 -52.315 ;
      RECT 109.955 -51.28 110.045 -50.272 ;
      RECT 109.905 -51.045 110.045 -50.875 ;
      RECT 109.955 -49.858 110.045 -48.85 ;
      RECT 109.905 -49.255 110.045 -49.085 ;
      RECT 109.955 -48.05 110.045 -47.042 ;
      RECT 109.905 -47.815 110.045 -47.645 ;
      RECT 109.955 -46.628 110.045 -45.62 ;
      RECT 109.905 -46.025 110.045 -45.855 ;
      RECT 109.955 -44.82 110.045 -43.812 ;
      RECT 109.905 -44.585 110.045 -44.415 ;
      RECT 109.955 -43.398 110.045 -42.39 ;
      RECT 109.905 -42.795 110.045 -42.625 ;
      RECT 109.955 -41.59 110.045 -40.582 ;
      RECT 109.905 -41.355 110.045 -41.185 ;
      RECT 109.955 -40.168 110.045 -39.16 ;
      RECT 109.905 -39.565 110.045 -39.395 ;
      RECT 109.955 -38.36 110.045 -37.352 ;
      RECT 109.905 -38.125 110.045 -37.955 ;
      RECT 109.955 -36.938 110.045 -35.93 ;
      RECT 109.905 -36.335 110.045 -36.165 ;
      RECT 109.955 -35.13 110.045 -34.122 ;
      RECT 109.905 -34.895 110.045 -34.725 ;
      RECT 109.955 -33.708 110.045 -32.7 ;
      RECT 109.905 -33.105 110.045 -32.935 ;
      RECT 109.955 -31.9 110.045 -30.892 ;
      RECT 109.905 -31.665 110.045 -31.495 ;
      RECT 109.955 -30.478 110.045 -29.47 ;
      RECT 109.905 -29.875 110.045 -29.705 ;
      RECT 109.955 -28.67 110.045 -27.662 ;
      RECT 109.905 -28.435 110.045 -28.265 ;
      RECT 109.955 -27.248 110.045 -26.24 ;
      RECT 109.905 -26.645 110.045 -26.475 ;
      RECT 109.955 -25.44 110.045 -24.432 ;
      RECT 109.905 -25.205 110.045 -25.035 ;
      RECT 109.955 -24.018 110.045 -23.01 ;
      RECT 109.905 -23.415 110.045 -23.245 ;
      RECT 109.955 -22.21 110.045 -21.202 ;
      RECT 109.905 -21.975 110.045 -21.805 ;
      RECT 109.955 -20.788 110.045 -19.78 ;
      RECT 109.905 -20.185 110.045 -20.015 ;
      RECT 109.955 -18.98 110.045 -17.972 ;
      RECT 109.905 -18.745 110.045 -18.575 ;
      RECT 109.955 -17.558 110.045 -16.55 ;
      RECT 109.905 -16.955 110.045 -16.785 ;
      RECT 109.955 -15.75 110.045 -14.742 ;
      RECT 109.905 -15.515 110.045 -15.345 ;
      RECT 109.955 -14.328 110.045 -13.32 ;
      RECT 109.905 -13.725 110.045 -13.555 ;
      RECT 109.955 -12.52 110.045 -11.512 ;
      RECT 109.905 -12.285 110.045 -12.115 ;
      RECT 109.955 -11.098 110.045 -10.09 ;
      RECT 109.905 -10.495 110.045 -10.325 ;
      RECT 109.955 -9.29 110.045 -8.282 ;
      RECT 109.905 -9.055 110.045 -8.885 ;
      RECT 109.955 -7.868 110.045 -6.86 ;
      RECT 109.905 -7.265 110.045 -7.095 ;
      RECT 109.955 -6.06 110.045 -5.052 ;
      RECT 109.905 -5.825 110.045 -5.655 ;
      RECT 109.955 -4.638 110.045 -3.63 ;
      RECT 109.905 -4.035 110.045 -3.865 ;
      RECT 109.955 -2.83 110.045 -1.822 ;
      RECT 109.905 -2.595 110.045 -2.425 ;
      RECT 109.955 -1.408 110.045 -0.4 ;
      RECT 109.905 -0.805 110.045 -0.635 ;
      RECT 109.955 0.4 110.045 1.408 ;
      RECT 109.905 0.635 110.045 0.805 ;
      RECT 108.525 -111.685 110.005 -111.585 ;
      RECT 108.525 -112.195 108.625 -111.585 ;
      RECT 108.745 -109.15 110.005 -109.05 ;
      RECT 109.905 -109.475 110.005 -109.05 ;
      RECT 109.345 -109.475 109.445 -109.05 ;
      RECT 108.785 -109.475 108.885 -109.05 ;
      RECT 109.555 -101.538 109.645 -100.531 ;
      RECT 109.555 -101.225 109.695 -101.055 ;
      RECT 109.555 -99.729 109.645 -98.722 ;
      RECT 109.555 -99.205 109.695 -99.035 ;
      RECT 109.555 -98.308 109.645 -97.301 ;
      RECT 109.555 -97.995 109.695 -97.825 ;
      RECT 109.555 -96.499 109.645 -95.492 ;
      RECT 109.555 -95.975 109.695 -95.805 ;
      RECT 109.555 -95.078 109.645 -94.071 ;
      RECT 109.555 -94.765 109.695 -94.595 ;
      RECT 109.555 -93.269 109.645 -92.262 ;
      RECT 109.555 -92.745 109.695 -92.575 ;
      RECT 109.555 -91.848 109.645 -90.841 ;
      RECT 109.555 -91.535 109.695 -91.365 ;
      RECT 109.555 -90.039 109.645 -89.032 ;
      RECT 109.555 -89.515 109.695 -89.345 ;
      RECT 109.555 -88.618 109.645 -87.611 ;
      RECT 109.555 -88.305 109.695 -88.135 ;
      RECT 109.555 -86.809 109.645 -85.802 ;
      RECT 109.555 -86.285 109.695 -86.115 ;
      RECT 109.555 -85.388 109.645 -84.381 ;
      RECT 109.555 -85.075 109.695 -84.905 ;
      RECT 109.555 -83.579 109.645 -82.572 ;
      RECT 109.555 -83.055 109.695 -82.885 ;
      RECT 109.555 -82.158 109.645 -81.151 ;
      RECT 109.555 -81.845 109.695 -81.675 ;
      RECT 109.555 -80.349 109.645 -79.342 ;
      RECT 109.555 -79.825 109.695 -79.655 ;
      RECT 109.555 -78.928 109.645 -77.921 ;
      RECT 109.555 -78.615 109.695 -78.445 ;
      RECT 109.555 -77.119 109.645 -76.112 ;
      RECT 109.555 -76.595 109.695 -76.425 ;
      RECT 109.555 -75.698 109.645 -74.691 ;
      RECT 109.555 -75.385 109.695 -75.215 ;
      RECT 109.555 -73.889 109.645 -72.882 ;
      RECT 109.555 -73.365 109.695 -73.195 ;
      RECT 109.555 -72.468 109.645 -71.461 ;
      RECT 109.555 -72.155 109.695 -71.985 ;
      RECT 109.555 -70.659 109.645 -69.652 ;
      RECT 109.555 -70.135 109.695 -69.965 ;
      RECT 109.555 -69.238 109.645 -68.231 ;
      RECT 109.555 -68.925 109.695 -68.755 ;
      RECT 109.555 -67.429 109.645 -66.422 ;
      RECT 109.555 -66.905 109.695 -66.735 ;
      RECT 109.555 -66.008 109.645 -65.001 ;
      RECT 109.555 -65.695 109.695 -65.525 ;
      RECT 109.555 -64.199 109.645 -63.192 ;
      RECT 109.555 -63.675 109.695 -63.505 ;
      RECT 109.555 -62.778 109.645 -61.771 ;
      RECT 109.555 -62.465 109.695 -62.295 ;
      RECT 109.555 -60.969 109.645 -59.962 ;
      RECT 109.555 -60.445 109.695 -60.275 ;
      RECT 109.555 -59.548 109.645 -58.541 ;
      RECT 109.555 -59.235 109.695 -59.065 ;
      RECT 109.555 -57.739 109.645 -56.732 ;
      RECT 109.555 -57.215 109.695 -57.045 ;
      RECT 109.555 -56.318 109.645 -55.311 ;
      RECT 109.555 -56.005 109.695 -55.835 ;
      RECT 109.555 -54.509 109.645 -53.502 ;
      RECT 109.555 -53.985 109.695 -53.815 ;
      RECT 109.555 -53.088 109.645 -52.081 ;
      RECT 109.555 -52.775 109.695 -52.605 ;
      RECT 109.555 -51.279 109.645 -50.272 ;
      RECT 109.555 -50.755 109.695 -50.585 ;
      RECT 109.555 -49.858 109.645 -48.851 ;
      RECT 109.555 -49.545 109.695 -49.375 ;
      RECT 109.555 -48.049 109.645 -47.042 ;
      RECT 109.555 -47.525 109.695 -47.355 ;
      RECT 109.555 -46.628 109.645 -45.621 ;
      RECT 109.555 -46.315 109.695 -46.145 ;
      RECT 109.555 -44.819 109.645 -43.812 ;
      RECT 109.555 -44.295 109.695 -44.125 ;
      RECT 109.555 -43.398 109.645 -42.391 ;
      RECT 109.555 -43.085 109.695 -42.915 ;
      RECT 109.555 -41.589 109.645 -40.582 ;
      RECT 109.555 -41.065 109.695 -40.895 ;
      RECT 109.555 -40.168 109.645 -39.161 ;
      RECT 109.555 -39.855 109.695 -39.685 ;
      RECT 109.555 -38.359 109.645 -37.352 ;
      RECT 109.555 -37.835 109.695 -37.665 ;
      RECT 109.555 -36.938 109.645 -35.931 ;
      RECT 109.555 -36.625 109.695 -36.455 ;
      RECT 109.555 -35.129 109.645 -34.122 ;
      RECT 109.555 -34.605 109.695 -34.435 ;
      RECT 109.555 -33.708 109.645 -32.701 ;
      RECT 109.555 -33.395 109.695 -33.225 ;
      RECT 109.555 -31.899 109.645 -30.892 ;
      RECT 109.555 -31.375 109.695 -31.205 ;
      RECT 109.555 -30.478 109.645 -29.471 ;
      RECT 109.555 -30.165 109.695 -29.995 ;
      RECT 109.555 -28.669 109.645 -27.662 ;
      RECT 109.555 -28.145 109.695 -27.975 ;
      RECT 109.555 -27.248 109.645 -26.241 ;
      RECT 109.555 -26.935 109.695 -26.765 ;
      RECT 109.555 -25.439 109.645 -24.432 ;
      RECT 109.555 -24.915 109.695 -24.745 ;
      RECT 109.555 -24.018 109.645 -23.011 ;
      RECT 109.555 -23.705 109.695 -23.535 ;
      RECT 109.555 -22.209 109.645 -21.202 ;
      RECT 109.555 -21.685 109.695 -21.515 ;
      RECT 109.555 -20.788 109.645 -19.781 ;
      RECT 109.555 -20.475 109.695 -20.305 ;
      RECT 109.555 -18.979 109.645 -17.972 ;
      RECT 109.555 -18.455 109.695 -18.285 ;
      RECT 109.555 -17.558 109.645 -16.551 ;
      RECT 109.555 -17.245 109.695 -17.075 ;
      RECT 109.555 -15.749 109.645 -14.742 ;
      RECT 109.555 -15.225 109.695 -15.055 ;
      RECT 109.555 -14.328 109.645 -13.321 ;
      RECT 109.555 -14.015 109.695 -13.845 ;
      RECT 109.555 -12.519 109.645 -11.512 ;
      RECT 109.555 -11.995 109.695 -11.825 ;
      RECT 109.555 -11.098 109.645 -10.091 ;
      RECT 109.555 -10.785 109.695 -10.615 ;
      RECT 109.555 -9.289 109.645 -8.282 ;
      RECT 109.555 -8.765 109.695 -8.595 ;
      RECT 109.555 -7.868 109.645 -6.861 ;
      RECT 109.555 -7.555 109.695 -7.385 ;
      RECT 109.555 -6.059 109.645 -5.052 ;
      RECT 109.555 -5.535 109.695 -5.365 ;
      RECT 109.555 -4.638 109.645 -3.631 ;
      RECT 109.555 -4.325 109.695 -4.155 ;
      RECT 109.555 -2.829 109.645 -1.822 ;
      RECT 109.555 -2.305 109.695 -2.135 ;
      RECT 109.555 -1.408 109.645 -0.401 ;
      RECT 109.555 -1.095 109.695 -0.925 ;
      RECT 109.555 0.401 109.645 1.408 ;
      RECT 109.555 0.925 109.695 1.095 ;
      RECT 108.885 -111.495 109.055 -111.385 ;
      RECT 105.735 -111.495 109.055 -111.395 ;
      RECT 108.755 -101.538 108.845 -100.53 ;
      RECT 108.705 -100.935 108.845 -100.765 ;
      RECT 108.755 -99.73 108.845 -98.722 ;
      RECT 108.705 -99.495 108.845 -99.325 ;
      RECT 108.755 -98.308 108.845 -97.3 ;
      RECT 108.705 -97.705 108.845 -97.535 ;
      RECT 108.755 -96.5 108.845 -95.492 ;
      RECT 108.705 -96.265 108.845 -96.095 ;
      RECT 108.755 -95.078 108.845 -94.07 ;
      RECT 108.705 -94.475 108.845 -94.305 ;
      RECT 108.755 -93.27 108.845 -92.262 ;
      RECT 108.705 -93.035 108.845 -92.865 ;
      RECT 108.755 -91.848 108.845 -90.84 ;
      RECT 108.705 -91.245 108.845 -91.075 ;
      RECT 108.755 -90.04 108.845 -89.032 ;
      RECT 108.705 -89.805 108.845 -89.635 ;
      RECT 108.755 -88.618 108.845 -87.61 ;
      RECT 108.705 -88.015 108.845 -87.845 ;
      RECT 108.755 -86.81 108.845 -85.802 ;
      RECT 108.705 -86.575 108.845 -86.405 ;
      RECT 108.755 -85.388 108.845 -84.38 ;
      RECT 108.705 -84.785 108.845 -84.615 ;
      RECT 108.755 -83.58 108.845 -82.572 ;
      RECT 108.705 -83.345 108.845 -83.175 ;
      RECT 108.755 -82.158 108.845 -81.15 ;
      RECT 108.705 -81.555 108.845 -81.385 ;
      RECT 108.755 -80.35 108.845 -79.342 ;
      RECT 108.705 -80.115 108.845 -79.945 ;
      RECT 108.755 -78.928 108.845 -77.92 ;
      RECT 108.705 -78.325 108.845 -78.155 ;
      RECT 108.755 -77.12 108.845 -76.112 ;
      RECT 108.705 -76.885 108.845 -76.715 ;
      RECT 108.755 -75.698 108.845 -74.69 ;
      RECT 108.705 -75.095 108.845 -74.925 ;
      RECT 108.755 -73.89 108.845 -72.882 ;
      RECT 108.705 -73.655 108.845 -73.485 ;
      RECT 108.755 -72.468 108.845 -71.46 ;
      RECT 108.705 -71.865 108.845 -71.695 ;
      RECT 108.755 -70.66 108.845 -69.652 ;
      RECT 108.705 -70.425 108.845 -70.255 ;
      RECT 108.755 -69.238 108.845 -68.23 ;
      RECT 108.705 -68.635 108.845 -68.465 ;
      RECT 108.755 -67.43 108.845 -66.422 ;
      RECT 108.705 -67.195 108.845 -67.025 ;
      RECT 108.755 -66.008 108.845 -65 ;
      RECT 108.705 -65.405 108.845 -65.235 ;
      RECT 108.755 -64.2 108.845 -63.192 ;
      RECT 108.705 -63.965 108.845 -63.795 ;
      RECT 108.755 -62.778 108.845 -61.77 ;
      RECT 108.705 -62.175 108.845 -62.005 ;
      RECT 108.755 -60.97 108.845 -59.962 ;
      RECT 108.705 -60.735 108.845 -60.565 ;
      RECT 108.755 -59.548 108.845 -58.54 ;
      RECT 108.705 -58.945 108.845 -58.775 ;
      RECT 108.755 -57.74 108.845 -56.732 ;
      RECT 108.705 -57.505 108.845 -57.335 ;
      RECT 108.755 -56.318 108.845 -55.31 ;
      RECT 108.705 -55.715 108.845 -55.545 ;
      RECT 108.755 -54.51 108.845 -53.502 ;
      RECT 108.705 -54.275 108.845 -54.105 ;
      RECT 108.755 -53.088 108.845 -52.08 ;
      RECT 108.705 -52.485 108.845 -52.315 ;
      RECT 108.755 -51.28 108.845 -50.272 ;
      RECT 108.705 -51.045 108.845 -50.875 ;
      RECT 108.755 -49.858 108.845 -48.85 ;
      RECT 108.705 -49.255 108.845 -49.085 ;
      RECT 108.755 -48.05 108.845 -47.042 ;
      RECT 108.705 -47.815 108.845 -47.645 ;
      RECT 108.755 -46.628 108.845 -45.62 ;
      RECT 108.705 -46.025 108.845 -45.855 ;
      RECT 108.755 -44.82 108.845 -43.812 ;
      RECT 108.705 -44.585 108.845 -44.415 ;
      RECT 108.755 -43.398 108.845 -42.39 ;
      RECT 108.705 -42.795 108.845 -42.625 ;
      RECT 108.755 -41.59 108.845 -40.582 ;
      RECT 108.705 -41.355 108.845 -41.185 ;
      RECT 108.755 -40.168 108.845 -39.16 ;
      RECT 108.705 -39.565 108.845 -39.395 ;
      RECT 108.755 -38.36 108.845 -37.352 ;
      RECT 108.705 -38.125 108.845 -37.955 ;
      RECT 108.755 -36.938 108.845 -35.93 ;
      RECT 108.705 -36.335 108.845 -36.165 ;
      RECT 108.755 -35.13 108.845 -34.122 ;
      RECT 108.705 -34.895 108.845 -34.725 ;
      RECT 108.755 -33.708 108.845 -32.7 ;
      RECT 108.705 -33.105 108.845 -32.935 ;
      RECT 108.755 -31.9 108.845 -30.892 ;
      RECT 108.705 -31.665 108.845 -31.495 ;
      RECT 108.755 -30.478 108.845 -29.47 ;
      RECT 108.705 -29.875 108.845 -29.705 ;
      RECT 108.755 -28.67 108.845 -27.662 ;
      RECT 108.705 -28.435 108.845 -28.265 ;
      RECT 108.755 -27.248 108.845 -26.24 ;
      RECT 108.705 -26.645 108.845 -26.475 ;
      RECT 108.755 -25.44 108.845 -24.432 ;
      RECT 108.705 -25.205 108.845 -25.035 ;
      RECT 108.755 -24.018 108.845 -23.01 ;
      RECT 108.705 -23.415 108.845 -23.245 ;
      RECT 108.755 -22.21 108.845 -21.202 ;
      RECT 108.705 -21.975 108.845 -21.805 ;
      RECT 108.755 -20.788 108.845 -19.78 ;
      RECT 108.705 -20.185 108.845 -20.015 ;
      RECT 108.755 -18.98 108.845 -17.972 ;
      RECT 108.705 -18.745 108.845 -18.575 ;
      RECT 108.755 -17.558 108.845 -16.55 ;
      RECT 108.705 -16.955 108.845 -16.785 ;
      RECT 108.755 -15.75 108.845 -14.742 ;
      RECT 108.705 -15.515 108.845 -15.345 ;
      RECT 108.755 -14.328 108.845 -13.32 ;
      RECT 108.705 -13.725 108.845 -13.555 ;
      RECT 108.755 -12.52 108.845 -11.512 ;
      RECT 108.705 -12.285 108.845 -12.115 ;
      RECT 108.755 -11.098 108.845 -10.09 ;
      RECT 108.705 -10.495 108.845 -10.325 ;
      RECT 108.755 -9.29 108.845 -8.282 ;
      RECT 108.705 -9.055 108.845 -8.885 ;
      RECT 108.755 -7.868 108.845 -6.86 ;
      RECT 108.705 -7.265 108.845 -7.095 ;
      RECT 108.755 -6.06 108.845 -5.052 ;
      RECT 108.705 -5.825 108.845 -5.655 ;
      RECT 108.755 -4.638 108.845 -3.63 ;
      RECT 108.705 -4.035 108.845 -3.865 ;
      RECT 108.755 -2.83 108.845 -1.822 ;
      RECT 108.705 -2.595 108.845 -2.425 ;
      RECT 108.755 -1.408 108.845 -0.4 ;
      RECT 108.705 -0.805 108.845 -0.635 ;
      RECT 108.755 0.4 108.845 1.408 ;
      RECT 108.705 0.635 108.845 0.805 ;
      RECT 108.355 -101.538 108.445 -100.531 ;
      RECT 108.355 -101.225 108.495 -101.055 ;
      RECT 108.355 -99.729 108.445 -98.722 ;
      RECT 108.355 -99.205 108.495 -99.035 ;
      RECT 108.355 -98.308 108.445 -97.301 ;
      RECT 108.355 -97.995 108.495 -97.825 ;
      RECT 108.355 -96.499 108.445 -95.492 ;
      RECT 108.355 -95.975 108.495 -95.805 ;
      RECT 108.355 -95.078 108.445 -94.071 ;
      RECT 108.355 -94.765 108.495 -94.595 ;
      RECT 108.355 -93.269 108.445 -92.262 ;
      RECT 108.355 -92.745 108.495 -92.575 ;
      RECT 108.355 -91.848 108.445 -90.841 ;
      RECT 108.355 -91.535 108.495 -91.365 ;
      RECT 108.355 -90.039 108.445 -89.032 ;
      RECT 108.355 -89.515 108.495 -89.345 ;
      RECT 108.355 -88.618 108.445 -87.611 ;
      RECT 108.355 -88.305 108.495 -88.135 ;
      RECT 108.355 -86.809 108.445 -85.802 ;
      RECT 108.355 -86.285 108.495 -86.115 ;
      RECT 108.355 -85.388 108.445 -84.381 ;
      RECT 108.355 -85.075 108.495 -84.905 ;
      RECT 108.355 -83.579 108.445 -82.572 ;
      RECT 108.355 -83.055 108.495 -82.885 ;
      RECT 108.355 -82.158 108.445 -81.151 ;
      RECT 108.355 -81.845 108.495 -81.675 ;
      RECT 108.355 -80.349 108.445 -79.342 ;
      RECT 108.355 -79.825 108.495 -79.655 ;
      RECT 108.355 -78.928 108.445 -77.921 ;
      RECT 108.355 -78.615 108.495 -78.445 ;
      RECT 108.355 -77.119 108.445 -76.112 ;
      RECT 108.355 -76.595 108.495 -76.425 ;
      RECT 108.355 -75.698 108.445 -74.691 ;
      RECT 108.355 -75.385 108.495 -75.215 ;
      RECT 108.355 -73.889 108.445 -72.882 ;
      RECT 108.355 -73.365 108.495 -73.195 ;
      RECT 108.355 -72.468 108.445 -71.461 ;
      RECT 108.355 -72.155 108.495 -71.985 ;
      RECT 108.355 -70.659 108.445 -69.652 ;
      RECT 108.355 -70.135 108.495 -69.965 ;
      RECT 108.355 -69.238 108.445 -68.231 ;
      RECT 108.355 -68.925 108.495 -68.755 ;
      RECT 108.355 -67.429 108.445 -66.422 ;
      RECT 108.355 -66.905 108.495 -66.735 ;
      RECT 108.355 -66.008 108.445 -65.001 ;
      RECT 108.355 -65.695 108.495 -65.525 ;
      RECT 108.355 -64.199 108.445 -63.192 ;
      RECT 108.355 -63.675 108.495 -63.505 ;
      RECT 108.355 -62.778 108.445 -61.771 ;
      RECT 108.355 -62.465 108.495 -62.295 ;
      RECT 108.355 -60.969 108.445 -59.962 ;
      RECT 108.355 -60.445 108.495 -60.275 ;
      RECT 108.355 -59.548 108.445 -58.541 ;
      RECT 108.355 -59.235 108.495 -59.065 ;
      RECT 108.355 -57.739 108.445 -56.732 ;
      RECT 108.355 -57.215 108.495 -57.045 ;
      RECT 108.355 -56.318 108.445 -55.311 ;
      RECT 108.355 -56.005 108.495 -55.835 ;
      RECT 108.355 -54.509 108.445 -53.502 ;
      RECT 108.355 -53.985 108.495 -53.815 ;
      RECT 108.355 -53.088 108.445 -52.081 ;
      RECT 108.355 -52.775 108.495 -52.605 ;
      RECT 108.355 -51.279 108.445 -50.272 ;
      RECT 108.355 -50.755 108.495 -50.585 ;
      RECT 108.355 -49.858 108.445 -48.851 ;
      RECT 108.355 -49.545 108.495 -49.375 ;
      RECT 108.355 -48.049 108.445 -47.042 ;
      RECT 108.355 -47.525 108.495 -47.355 ;
      RECT 108.355 -46.628 108.445 -45.621 ;
      RECT 108.355 -46.315 108.495 -46.145 ;
      RECT 108.355 -44.819 108.445 -43.812 ;
      RECT 108.355 -44.295 108.495 -44.125 ;
      RECT 108.355 -43.398 108.445 -42.391 ;
      RECT 108.355 -43.085 108.495 -42.915 ;
      RECT 108.355 -41.589 108.445 -40.582 ;
      RECT 108.355 -41.065 108.495 -40.895 ;
      RECT 108.355 -40.168 108.445 -39.161 ;
      RECT 108.355 -39.855 108.495 -39.685 ;
      RECT 108.355 -38.359 108.445 -37.352 ;
      RECT 108.355 -37.835 108.495 -37.665 ;
      RECT 108.355 -36.938 108.445 -35.931 ;
      RECT 108.355 -36.625 108.495 -36.455 ;
      RECT 108.355 -35.129 108.445 -34.122 ;
      RECT 108.355 -34.605 108.495 -34.435 ;
      RECT 108.355 -33.708 108.445 -32.701 ;
      RECT 108.355 -33.395 108.495 -33.225 ;
      RECT 108.355 -31.899 108.445 -30.892 ;
      RECT 108.355 -31.375 108.495 -31.205 ;
      RECT 108.355 -30.478 108.445 -29.471 ;
      RECT 108.355 -30.165 108.495 -29.995 ;
      RECT 108.355 -28.669 108.445 -27.662 ;
      RECT 108.355 -28.145 108.495 -27.975 ;
      RECT 108.355 -27.248 108.445 -26.241 ;
      RECT 108.355 -26.935 108.495 -26.765 ;
      RECT 108.355 -25.439 108.445 -24.432 ;
      RECT 108.355 -24.915 108.495 -24.745 ;
      RECT 108.355 -24.018 108.445 -23.011 ;
      RECT 108.355 -23.705 108.495 -23.535 ;
      RECT 108.355 -22.209 108.445 -21.202 ;
      RECT 108.355 -21.685 108.495 -21.515 ;
      RECT 108.355 -20.788 108.445 -19.781 ;
      RECT 108.355 -20.475 108.495 -20.305 ;
      RECT 108.355 -18.979 108.445 -17.972 ;
      RECT 108.355 -18.455 108.495 -18.285 ;
      RECT 108.355 -17.558 108.445 -16.551 ;
      RECT 108.355 -17.245 108.495 -17.075 ;
      RECT 108.355 -15.749 108.445 -14.742 ;
      RECT 108.355 -15.225 108.495 -15.055 ;
      RECT 108.355 -14.328 108.445 -13.321 ;
      RECT 108.355 -14.015 108.495 -13.845 ;
      RECT 108.355 -12.519 108.445 -11.512 ;
      RECT 108.355 -11.995 108.495 -11.825 ;
      RECT 108.355 -11.098 108.445 -10.091 ;
      RECT 108.355 -10.785 108.495 -10.615 ;
      RECT 108.355 -9.289 108.445 -8.282 ;
      RECT 108.355 -8.765 108.495 -8.595 ;
      RECT 108.355 -7.868 108.445 -6.861 ;
      RECT 108.355 -7.555 108.495 -7.385 ;
      RECT 108.355 -6.059 108.445 -5.052 ;
      RECT 108.355 -5.535 108.495 -5.365 ;
      RECT 108.355 -4.638 108.445 -3.631 ;
      RECT 108.355 -4.325 108.495 -4.155 ;
      RECT 108.355 -2.829 108.445 -1.822 ;
      RECT 108.355 -2.305 108.495 -2.135 ;
      RECT 108.355 -1.408 108.445 -0.401 ;
      RECT 108.355 -1.095 108.495 -0.925 ;
      RECT 108.355 0.401 108.445 1.408 ;
      RECT 108.355 0.925 108.495 1.095 ;
      RECT 106.505 -111.685 107.985 -111.585 ;
      RECT 106.505 -112.055 106.605 -111.585 ;
      RECT 106.31 -114.395 107.885 -114.275 ;
      RECT 107.785 -114.895 107.885 -114.275 ;
      RECT 107.19 -114.895 107.29 -114.275 ;
      RECT 106.31 -114.85 106.41 -114.275 ;
      RECT 107.555 -101.538 107.645 -100.53 ;
      RECT 107.505 -100.935 107.645 -100.765 ;
      RECT 107.555 -99.73 107.645 -98.722 ;
      RECT 107.505 -99.495 107.645 -99.325 ;
      RECT 107.555 -98.308 107.645 -97.3 ;
      RECT 107.505 -97.705 107.645 -97.535 ;
      RECT 107.555 -96.5 107.645 -95.492 ;
      RECT 107.505 -96.265 107.645 -96.095 ;
      RECT 107.555 -95.078 107.645 -94.07 ;
      RECT 107.505 -94.475 107.645 -94.305 ;
      RECT 107.555 -93.27 107.645 -92.262 ;
      RECT 107.505 -93.035 107.645 -92.865 ;
      RECT 107.555 -91.848 107.645 -90.84 ;
      RECT 107.505 -91.245 107.645 -91.075 ;
      RECT 107.555 -90.04 107.645 -89.032 ;
      RECT 107.505 -89.805 107.645 -89.635 ;
      RECT 107.555 -88.618 107.645 -87.61 ;
      RECT 107.505 -88.015 107.645 -87.845 ;
      RECT 107.555 -86.81 107.645 -85.802 ;
      RECT 107.505 -86.575 107.645 -86.405 ;
      RECT 107.555 -85.388 107.645 -84.38 ;
      RECT 107.505 -84.785 107.645 -84.615 ;
      RECT 107.555 -83.58 107.645 -82.572 ;
      RECT 107.505 -83.345 107.645 -83.175 ;
      RECT 107.555 -82.158 107.645 -81.15 ;
      RECT 107.505 -81.555 107.645 -81.385 ;
      RECT 107.555 -80.35 107.645 -79.342 ;
      RECT 107.505 -80.115 107.645 -79.945 ;
      RECT 107.555 -78.928 107.645 -77.92 ;
      RECT 107.505 -78.325 107.645 -78.155 ;
      RECT 107.555 -77.12 107.645 -76.112 ;
      RECT 107.505 -76.885 107.645 -76.715 ;
      RECT 107.555 -75.698 107.645 -74.69 ;
      RECT 107.505 -75.095 107.645 -74.925 ;
      RECT 107.555 -73.89 107.645 -72.882 ;
      RECT 107.505 -73.655 107.645 -73.485 ;
      RECT 107.555 -72.468 107.645 -71.46 ;
      RECT 107.505 -71.865 107.645 -71.695 ;
      RECT 107.555 -70.66 107.645 -69.652 ;
      RECT 107.505 -70.425 107.645 -70.255 ;
      RECT 107.555 -69.238 107.645 -68.23 ;
      RECT 107.505 -68.635 107.645 -68.465 ;
      RECT 107.555 -67.43 107.645 -66.422 ;
      RECT 107.505 -67.195 107.645 -67.025 ;
      RECT 107.555 -66.008 107.645 -65 ;
      RECT 107.505 -65.405 107.645 -65.235 ;
      RECT 107.555 -64.2 107.645 -63.192 ;
      RECT 107.505 -63.965 107.645 -63.795 ;
      RECT 107.555 -62.778 107.645 -61.77 ;
      RECT 107.505 -62.175 107.645 -62.005 ;
      RECT 107.555 -60.97 107.645 -59.962 ;
      RECT 107.505 -60.735 107.645 -60.565 ;
      RECT 107.555 -59.548 107.645 -58.54 ;
      RECT 107.505 -58.945 107.645 -58.775 ;
      RECT 107.555 -57.74 107.645 -56.732 ;
      RECT 107.505 -57.505 107.645 -57.335 ;
      RECT 107.555 -56.318 107.645 -55.31 ;
      RECT 107.505 -55.715 107.645 -55.545 ;
      RECT 107.555 -54.51 107.645 -53.502 ;
      RECT 107.505 -54.275 107.645 -54.105 ;
      RECT 107.555 -53.088 107.645 -52.08 ;
      RECT 107.505 -52.485 107.645 -52.315 ;
      RECT 107.555 -51.28 107.645 -50.272 ;
      RECT 107.505 -51.045 107.645 -50.875 ;
      RECT 107.555 -49.858 107.645 -48.85 ;
      RECT 107.505 -49.255 107.645 -49.085 ;
      RECT 107.555 -48.05 107.645 -47.042 ;
      RECT 107.505 -47.815 107.645 -47.645 ;
      RECT 107.555 -46.628 107.645 -45.62 ;
      RECT 107.505 -46.025 107.645 -45.855 ;
      RECT 107.555 -44.82 107.645 -43.812 ;
      RECT 107.505 -44.585 107.645 -44.415 ;
      RECT 107.555 -43.398 107.645 -42.39 ;
      RECT 107.505 -42.795 107.645 -42.625 ;
      RECT 107.555 -41.59 107.645 -40.582 ;
      RECT 107.505 -41.355 107.645 -41.185 ;
      RECT 107.555 -40.168 107.645 -39.16 ;
      RECT 107.505 -39.565 107.645 -39.395 ;
      RECT 107.555 -38.36 107.645 -37.352 ;
      RECT 107.505 -38.125 107.645 -37.955 ;
      RECT 107.555 -36.938 107.645 -35.93 ;
      RECT 107.505 -36.335 107.645 -36.165 ;
      RECT 107.555 -35.13 107.645 -34.122 ;
      RECT 107.505 -34.895 107.645 -34.725 ;
      RECT 107.555 -33.708 107.645 -32.7 ;
      RECT 107.505 -33.105 107.645 -32.935 ;
      RECT 107.555 -31.9 107.645 -30.892 ;
      RECT 107.505 -31.665 107.645 -31.495 ;
      RECT 107.555 -30.478 107.645 -29.47 ;
      RECT 107.505 -29.875 107.645 -29.705 ;
      RECT 107.555 -28.67 107.645 -27.662 ;
      RECT 107.505 -28.435 107.645 -28.265 ;
      RECT 107.555 -27.248 107.645 -26.24 ;
      RECT 107.505 -26.645 107.645 -26.475 ;
      RECT 107.555 -25.44 107.645 -24.432 ;
      RECT 107.505 -25.205 107.645 -25.035 ;
      RECT 107.555 -24.018 107.645 -23.01 ;
      RECT 107.505 -23.415 107.645 -23.245 ;
      RECT 107.555 -22.21 107.645 -21.202 ;
      RECT 107.505 -21.975 107.645 -21.805 ;
      RECT 107.555 -20.788 107.645 -19.78 ;
      RECT 107.505 -20.185 107.645 -20.015 ;
      RECT 107.555 -18.98 107.645 -17.972 ;
      RECT 107.505 -18.745 107.645 -18.575 ;
      RECT 107.555 -17.558 107.645 -16.55 ;
      RECT 107.505 -16.955 107.645 -16.785 ;
      RECT 107.555 -15.75 107.645 -14.742 ;
      RECT 107.505 -15.515 107.645 -15.345 ;
      RECT 107.555 -14.328 107.645 -13.32 ;
      RECT 107.505 -13.725 107.645 -13.555 ;
      RECT 107.555 -12.52 107.645 -11.512 ;
      RECT 107.505 -12.285 107.645 -12.115 ;
      RECT 107.555 -11.098 107.645 -10.09 ;
      RECT 107.505 -10.495 107.645 -10.325 ;
      RECT 107.555 -9.29 107.645 -8.282 ;
      RECT 107.505 -9.055 107.645 -8.885 ;
      RECT 107.555 -7.868 107.645 -6.86 ;
      RECT 107.505 -7.265 107.645 -7.095 ;
      RECT 107.555 -6.06 107.645 -5.052 ;
      RECT 107.505 -5.825 107.645 -5.655 ;
      RECT 107.555 -4.638 107.645 -3.63 ;
      RECT 107.505 -4.035 107.645 -3.865 ;
      RECT 107.555 -2.83 107.645 -1.822 ;
      RECT 107.505 -2.595 107.645 -2.425 ;
      RECT 107.555 -1.408 107.645 -0.4 ;
      RECT 107.505 -0.805 107.645 -0.635 ;
      RECT 107.555 0.4 107.645 1.408 ;
      RECT 107.505 0.635 107.645 0.805 ;
      RECT 107.43 -114.685 107.605 -114.515 ;
      RECT 107.505 -114.895 107.605 -114.515 ;
      RECT 106.545 -113.555 106.645 -113.09 ;
      RECT 106.91 -113.555 107.01 -113.1 ;
      RECT 106.545 -113.555 107.39 -113.385 ;
      RECT 107.155 -101.538 107.245 -100.531 ;
      RECT 107.155 -101.225 107.295 -101.055 ;
      RECT 107.155 -99.729 107.245 -98.722 ;
      RECT 107.155 -99.205 107.295 -99.035 ;
      RECT 107.155 -98.308 107.245 -97.301 ;
      RECT 107.155 -97.995 107.295 -97.825 ;
      RECT 107.155 -96.499 107.245 -95.492 ;
      RECT 107.155 -95.975 107.295 -95.805 ;
      RECT 107.155 -95.078 107.245 -94.071 ;
      RECT 107.155 -94.765 107.295 -94.595 ;
      RECT 107.155 -93.269 107.245 -92.262 ;
      RECT 107.155 -92.745 107.295 -92.575 ;
      RECT 107.155 -91.848 107.245 -90.841 ;
      RECT 107.155 -91.535 107.295 -91.365 ;
      RECT 107.155 -90.039 107.245 -89.032 ;
      RECT 107.155 -89.515 107.295 -89.345 ;
      RECT 107.155 -88.618 107.245 -87.611 ;
      RECT 107.155 -88.305 107.295 -88.135 ;
      RECT 107.155 -86.809 107.245 -85.802 ;
      RECT 107.155 -86.285 107.295 -86.115 ;
      RECT 107.155 -85.388 107.245 -84.381 ;
      RECT 107.155 -85.075 107.295 -84.905 ;
      RECT 107.155 -83.579 107.245 -82.572 ;
      RECT 107.155 -83.055 107.295 -82.885 ;
      RECT 107.155 -82.158 107.245 -81.151 ;
      RECT 107.155 -81.845 107.295 -81.675 ;
      RECT 107.155 -80.349 107.245 -79.342 ;
      RECT 107.155 -79.825 107.295 -79.655 ;
      RECT 107.155 -78.928 107.245 -77.921 ;
      RECT 107.155 -78.615 107.295 -78.445 ;
      RECT 107.155 -77.119 107.245 -76.112 ;
      RECT 107.155 -76.595 107.295 -76.425 ;
      RECT 107.155 -75.698 107.245 -74.691 ;
      RECT 107.155 -75.385 107.295 -75.215 ;
      RECT 107.155 -73.889 107.245 -72.882 ;
      RECT 107.155 -73.365 107.295 -73.195 ;
      RECT 107.155 -72.468 107.245 -71.461 ;
      RECT 107.155 -72.155 107.295 -71.985 ;
      RECT 107.155 -70.659 107.245 -69.652 ;
      RECT 107.155 -70.135 107.295 -69.965 ;
      RECT 107.155 -69.238 107.245 -68.231 ;
      RECT 107.155 -68.925 107.295 -68.755 ;
      RECT 107.155 -67.429 107.245 -66.422 ;
      RECT 107.155 -66.905 107.295 -66.735 ;
      RECT 107.155 -66.008 107.245 -65.001 ;
      RECT 107.155 -65.695 107.295 -65.525 ;
      RECT 107.155 -64.199 107.245 -63.192 ;
      RECT 107.155 -63.675 107.295 -63.505 ;
      RECT 107.155 -62.778 107.245 -61.771 ;
      RECT 107.155 -62.465 107.295 -62.295 ;
      RECT 107.155 -60.969 107.245 -59.962 ;
      RECT 107.155 -60.445 107.295 -60.275 ;
      RECT 107.155 -59.548 107.245 -58.541 ;
      RECT 107.155 -59.235 107.295 -59.065 ;
      RECT 107.155 -57.739 107.245 -56.732 ;
      RECT 107.155 -57.215 107.295 -57.045 ;
      RECT 107.155 -56.318 107.245 -55.311 ;
      RECT 107.155 -56.005 107.295 -55.835 ;
      RECT 107.155 -54.509 107.245 -53.502 ;
      RECT 107.155 -53.985 107.295 -53.815 ;
      RECT 107.155 -53.088 107.245 -52.081 ;
      RECT 107.155 -52.775 107.295 -52.605 ;
      RECT 107.155 -51.279 107.245 -50.272 ;
      RECT 107.155 -50.755 107.295 -50.585 ;
      RECT 107.155 -49.858 107.245 -48.851 ;
      RECT 107.155 -49.545 107.295 -49.375 ;
      RECT 107.155 -48.049 107.245 -47.042 ;
      RECT 107.155 -47.525 107.295 -47.355 ;
      RECT 107.155 -46.628 107.245 -45.621 ;
      RECT 107.155 -46.315 107.295 -46.145 ;
      RECT 107.155 -44.819 107.245 -43.812 ;
      RECT 107.155 -44.295 107.295 -44.125 ;
      RECT 107.155 -43.398 107.245 -42.391 ;
      RECT 107.155 -43.085 107.295 -42.915 ;
      RECT 107.155 -41.589 107.245 -40.582 ;
      RECT 107.155 -41.065 107.295 -40.895 ;
      RECT 107.155 -40.168 107.245 -39.161 ;
      RECT 107.155 -39.855 107.295 -39.685 ;
      RECT 107.155 -38.359 107.245 -37.352 ;
      RECT 107.155 -37.835 107.295 -37.665 ;
      RECT 107.155 -36.938 107.245 -35.931 ;
      RECT 107.155 -36.625 107.295 -36.455 ;
      RECT 107.155 -35.129 107.245 -34.122 ;
      RECT 107.155 -34.605 107.295 -34.435 ;
      RECT 107.155 -33.708 107.245 -32.701 ;
      RECT 107.155 -33.395 107.295 -33.225 ;
      RECT 107.155 -31.899 107.245 -30.892 ;
      RECT 107.155 -31.375 107.295 -31.205 ;
      RECT 107.155 -30.478 107.245 -29.471 ;
      RECT 107.155 -30.165 107.295 -29.995 ;
      RECT 107.155 -28.669 107.245 -27.662 ;
      RECT 107.155 -28.145 107.295 -27.975 ;
      RECT 107.155 -27.248 107.245 -26.241 ;
      RECT 107.155 -26.935 107.295 -26.765 ;
      RECT 107.155 -25.439 107.245 -24.432 ;
      RECT 107.155 -24.915 107.295 -24.745 ;
      RECT 107.155 -24.018 107.245 -23.011 ;
      RECT 107.155 -23.705 107.295 -23.535 ;
      RECT 107.155 -22.209 107.245 -21.202 ;
      RECT 107.155 -21.685 107.295 -21.515 ;
      RECT 107.155 -20.788 107.245 -19.781 ;
      RECT 107.155 -20.475 107.295 -20.305 ;
      RECT 107.155 -18.979 107.245 -17.972 ;
      RECT 107.155 -18.455 107.295 -18.285 ;
      RECT 107.155 -17.558 107.245 -16.551 ;
      RECT 107.155 -17.245 107.295 -17.075 ;
      RECT 107.155 -15.749 107.245 -14.742 ;
      RECT 107.155 -15.225 107.295 -15.055 ;
      RECT 107.155 -14.328 107.245 -13.321 ;
      RECT 107.155 -14.015 107.295 -13.845 ;
      RECT 107.155 -12.519 107.245 -11.512 ;
      RECT 107.155 -11.995 107.295 -11.825 ;
      RECT 107.155 -11.098 107.245 -10.091 ;
      RECT 107.155 -10.785 107.295 -10.615 ;
      RECT 107.155 -9.289 107.245 -8.282 ;
      RECT 107.155 -8.765 107.295 -8.595 ;
      RECT 107.155 -7.868 107.245 -6.861 ;
      RECT 107.155 -7.555 107.295 -7.385 ;
      RECT 107.155 -6.059 107.245 -5.052 ;
      RECT 107.155 -5.535 107.295 -5.365 ;
      RECT 107.155 -4.638 107.245 -3.631 ;
      RECT 107.155 -4.325 107.295 -4.155 ;
      RECT 107.155 -2.829 107.245 -1.822 ;
      RECT 107.155 -2.305 107.295 -2.135 ;
      RECT 107.155 -1.408 107.245 -0.401 ;
      RECT 107.155 -1.095 107.295 -0.925 ;
      RECT 107.155 0.401 107.245 1.408 ;
      RECT 107.155 0.925 107.295 1.095 ;
      RECT 106.84 -114.685 107.01 -114.515 ;
      RECT 106.91 -114.895 107.01 -114.515 ;
      RECT 106.355 -101.538 106.445 -100.53 ;
      RECT 106.305 -100.935 106.445 -100.765 ;
      RECT 106.355 -99.73 106.445 -98.722 ;
      RECT 106.305 -99.495 106.445 -99.325 ;
      RECT 106.355 -98.308 106.445 -97.3 ;
      RECT 106.305 -97.705 106.445 -97.535 ;
      RECT 106.355 -96.5 106.445 -95.492 ;
      RECT 106.305 -96.265 106.445 -96.095 ;
      RECT 106.355 -95.078 106.445 -94.07 ;
      RECT 106.305 -94.475 106.445 -94.305 ;
      RECT 106.355 -93.27 106.445 -92.262 ;
      RECT 106.305 -93.035 106.445 -92.865 ;
      RECT 106.355 -91.848 106.445 -90.84 ;
      RECT 106.305 -91.245 106.445 -91.075 ;
      RECT 106.355 -90.04 106.445 -89.032 ;
      RECT 106.305 -89.805 106.445 -89.635 ;
      RECT 106.355 -88.618 106.445 -87.61 ;
      RECT 106.305 -88.015 106.445 -87.845 ;
      RECT 106.355 -86.81 106.445 -85.802 ;
      RECT 106.305 -86.575 106.445 -86.405 ;
      RECT 106.355 -85.388 106.445 -84.38 ;
      RECT 106.305 -84.785 106.445 -84.615 ;
      RECT 106.355 -83.58 106.445 -82.572 ;
      RECT 106.305 -83.345 106.445 -83.175 ;
      RECT 106.355 -82.158 106.445 -81.15 ;
      RECT 106.305 -81.555 106.445 -81.385 ;
      RECT 106.355 -80.35 106.445 -79.342 ;
      RECT 106.305 -80.115 106.445 -79.945 ;
      RECT 106.355 -78.928 106.445 -77.92 ;
      RECT 106.305 -78.325 106.445 -78.155 ;
      RECT 106.355 -77.12 106.445 -76.112 ;
      RECT 106.305 -76.885 106.445 -76.715 ;
      RECT 106.355 -75.698 106.445 -74.69 ;
      RECT 106.305 -75.095 106.445 -74.925 ;
      RECT 106.355 -73.89 106.445 -72.882 ;
      RECT 106.305 -73.655 106.445 -73.485 ;
      RECT 106.355 -72.468 106.445 -71.46 ;
      RECT 106.305 -71.865 106.445 -71.695 ;
      RECT 106.355 -70.66 106.445 -69.652 ;
      RECT 106.305 -70.425 106.445 -70.255 ;
      RECT 106.355 -69.238 106.445 -68.23 ;
      RECT 106.305 -68.635 106.445 -68.465 ;
      RECT 106.355 -67.43 106.445 -66.422 ;
      RECT 106.305 -67.195 106.445 -67.025 ;
      RECT 106.355 -66.008 106.445 -65 ;
      RECT 106.305 -65.405 106.445 -65.235 ;
      RECT 106.355 -64.2 106.445 -63.192 ;
      RECT 106.305 -63.965 106.445 -63.795 ;
      RECT 106.355 -62.778 106.445 -61.77 ;
      RECT 106.305 -62.175 106.445 -62.005 ;
      RECT 106.355 -60.97 106.445 -59.962 ;
      RECT 106.305 -60.735 106.445 -60.565 ;
      RECT 106.355 -59.548 106.445 -58.54 ;
      RECT 106.305 -58.945 106.445 -58.775 ;
      RECT 106.355 -57.74 106.445 -56.732 ;
      RECT 106.305 -57.505 106.445 -57.335 ;
      RECT 106.355 -56.318 106.445 -55.31 ;
      RECT 106.305 -55.715 106.445 -55.545 ;
      RECT 106.355 -54.51 106.445 -53.502 ;
      RECT 106.305 -54.275 106.445 -54.105 ;
      RECT 106.355 -53.088 106.445 -52.08 ;
      RECT 106.305 -52.485 106.445 -52.315 ;
      RECT 106.355 -51.28 106.445 -50.272 ;
      RECT 106.305 -51.045 106.445 -50.875 ;
      RECT 106.355 -49.858 106.445 -48.85 ;
      RECT 106.305 -49.255 106.445 -49.085 ;
      RECT 106.355 -48.05 106.445 -47.042 ;
      RECT 106.305 -47.815 106.445 -47.645 ;
      RECT 106.355 -46.628 106.445 -45.62 ;
      RECT 106.305 -46.025 106.445 -45.855 ;
      RECT 106.355 -44.82 106.445 -43.812 ;
      RECT 106.305 -44.585 106.445 -44.415 ;
      RECT 106.355 -43.398 106.445 -42.39 ;
      RECT 106.305 -42.795 106.445 -42.625 ;
      RECT 106.355 -41.59 106.445 -40.582 ;
      RECT 106.305 -41.355 106.445 -41.185 ;
      RECT 106.355 -40.168 106.445 -39.16 ;
      RECT 106.305 -39.565 106.445 -39.395 ;
      RECT 106.355 -38.36 106.445 -37.352 ;
      RECT 106.305 -38.125 106.445 -37.955 ;
      RECT 106.355 -36.938 106.445 -35.93 ;
      RECT 106.305 -36.335 106.445 -36.165 ;
      RECT 106.355 -35.13 106.445 -34.122 ;
      RECT 106.305 -34.895 106.445 -34.725 ;
      RECT 106.355 -33.708 106.445 -32.7 ;
      RECT 106.305 -33.105 106.445 -32.935 ;
      RECT 106.355 -31.9 106.445 -30.892 ;
      RECT 106.305 -31.665 106.445 -31.495 ;
      RECT 106.355 -30.478 106.445 -29.47 ;
      RECT 106.305 -29.875 106.445 -29.705 ;
      RECT 106.355 -28.67 106.445 -27.662 ;
      RECT 106.305 -28.435 106.445 -28.265 ;
      RECT 106.355 -27.248 106.445 -26.24 ;
      RECT 106.305 -26.645 106.445 -26.475 ;
      RECT 106.355 -25.44 106.445 -24.432 ;
      RECT 106.305 -25.205 106.445 -25.035 ;
      RECT 106.355 -24.018 106.445 -23.01 ;
      RECT 106.305 -23.415 106.445 -23.245 ;
      RECT 106.355 -22.21 106.445 -21.202 ;
      RECT 106.305 -21.975 106.445 -21.805 ;
      RECT 106.355 -20.788 106.445 -19.78 ;
      RECT 106.305 -20.185 106.445 -20.015 ;
      RECT 106.355 -18.98 106.445 -17.972 ;
      RECT 106.305 -18.745 106.445 -18.575 ;
      RECT 106.355 -17.558 106.445 -16.55 ;
      RECT 106.305 -16.955 106.445 -16.785 ;
      RECT 106.355 -15.75 106.445 -14.742 ;
      RECT 106.305 -15.515 106.445 -15.345 ;
      RECT 106.355 -14.328 106.445 -13.32 ;
      RECT 106.305 -13.725 106.445 -13.555 ;
      RECT 106.355 -12.52 106.445 -11.512 ;
      RECT 106.305 -12.285 106.445 -12.115 ;
      RECT 106.355 -11.098 106.445 -10.09 ;
      RECT 106.305 -10.495 106.445 -10.325 ;
      RECT 106.355 -9.29 106.445 -8.282 ;
      RECT 106.305 -9.055 106.445 -8.885 ;
      RECT 106.355 -7.868 106.445 -6.86 ;
      RECT 106.305 -7.265 106.445 -7.095 ;
      RECT 106.355 -6.06 106.445 -5.052 ;
      RECT 106.305 -5.825 106.445 -5.655 ;
      RECT 106.355 -4.638 106.445 -3.63 ;
      RECT 106.305 -4.035 106.445 -3.865 ;
      RECT 106.355 -2.83 106.445 -1.822 ;
      RECT 106.305 -2.595 106.445 -2.425 ;
      RECT 106.355 -1.408 106.445 -0.4 ;
      RECT 106.305 -0.805 106.445 -0.635 ;
      RECT 106.355 0.4 106.445 1.408 ;
      RECT 106.305 0.635 106.445 0.805 ;
      RECT 105.955 -101.538 106.045 -100.531 ;
      RECT 105.955 -101.225 106.095 -101.055 ;
      RECT 105.955 -99.729 106.045 -98.722 ;
      RECT 105.955 -99.205 106.095 -99.035 ;
      RECT 105.955 -98.308 106.045 -97.301 ;
      RECT 105.955 -97.995 106.095 -97.825 ;
      RECT 105.955 -96.499 106.045 -95.492 ;
      RECT 105.955 -95.975 106.095 -95.805 ;
      RECT 105.955 -95.078 106.045 -94.071 ;
      RECT 105.955 -94.765 106.095 -94.595 ;
      RECT 105.955 -93.269 106.045 -92.262 ;
      RECT 105.955 -92.745 106.095 -92.575 ;
      RECT 105.955 -91.848 106.045 -90.841 ;
      RECT 105.955 -91.535 106.095 -91.365 ;
      RECT 105.955 -90.039 106.045 -89.032 ;
      RECT 105.955 -89.515 106.095 -89.345 ;
      RECT 105.955 -88.618 106.045 -87.611 ;
      RECT 105.955 -88.305 106.095 -88.135 ;
      RECT 105.955 -86.809 106.045 -85.802 ;
      RECT 105.955 -86.285 106.095 -86.115 ;
      RECT 105.955 -85.388 106.045 -84.381 ;
      RECT 105.955 -85.075 106.095 -84.905 ;
      RECT 105.955 -83.579 106.045 -82.572 ;
      RECT 105.955 -83.055 106.095 -82.885 ;
      RECT 105.955 -82.158 106.045 -81.151 ;
      RECT 105.955 -81.845 106.095 -81.675 ;
      RECT 105.955 -80.349 106.045 -79.342 ;
      RECT 105.955 -79.825 106.095 -79.655 ;
      RECT 105.955 -78.928 106.045 -77.921 ;
      RECT 105.955 -78.615 106.095 -78.445 ;
      RECT 105.955 -77.119 106.045 -76.112 ;
      RECT 105.955 -76.595 106.095 -76.425 ;
      RECT 105.955 -75.698 106.045 -74.691 ;
      RECT 105.955 -75.385 106.095 -75.215 ;
      RECT 105.955 -73.889 106.045 -72.882 ;
      RECT 105.955 -73.365 106.095 -73.195 ;
      RECT 105.955 -72.468 106.045 -71.461 ;
      RECT 105.955 -72.155 106.095 -71.985 ;
      RECT 105.955 -70.659 106.045 -69.652 ;
      RECT 105.955 -70.135 106.095 -69.965 ;
      RECT 105.955 -69.238 106.045 -68.231 ;
      RECT 105.955 -68.925 106.095 -68.755 ;
      RECT 105.955 -67.429 106.045 -66.422 ;
      RECT 105.955 -66.905 106.095 -66.735 ;
      RECT 105.955 -66.008 106.045 -65.001 ;
      RECT 105.955 -65.695 106.095 -65.525 ;
      RECT 105.955 -64.199 106.045 -63.192 ;
      RECT 105.955 -63.675 106.095 -63.505 ;
      RECT 105.955 -62.778 106.045 -61.771 ;
      RECT 105.955 -62.465 106.095 -62.295 ;
      RECT 105.955 -60.969 106.045 -59.962 ;
      RECT 105.955 -60.445 106.095 -60.275 ;
      RECT 105.955 -59.548 106.045 -58.541 ;
      RECT 105.955 -59.235 106.095 -59.065 ;
      RECT 105.955 -57.739 106.045 -56.732 ;
      RECT 105.955 -57.215 106.095 -57.045 ;
      RECT 105.955 -56.318 106.045 -55.311 ;
      RECT 105.955 -56.005 106.095 -55.835 ;
      RECT 105.955 -54.509 106.045 -53.502 ;
      RECT 105.955 -53.985 106.095 -53.815 ;
      RECT 105.955 -53.088 106.045 -52.081 ;
      RECT 105.955 -52.775 106.095 -52.605 ;
      RECT 105.955 -51.279 106.045 -50.272 ;
      RECT 105.955 -50.755 106.095 -50.585 ;
      RECT 105.955 -49.858 106.045 -48.851 ;
      RECT 105.955 -49.545 106.095 -49.375 ;
      RECT 105.955 -48.049 106.045 -47.042 ;
      RECT 105.955 -47.525 106.095 -47.355 ;
      RECT 105.955 -46.628 106.045 -45.621 ;
      RECT 105.955 -46.315 106.095 -46.145 ;
      RECT 105.955 -44.819 106.045 -43.812 ;
      RECT 105.955 -44.295 106.095 -44.125 ;
      RECT 105.955 -43.398 106.045 -42.391 ;
      RECT 105.955 -43.085 106.095 -42.915 ;
      RECT 105.955 -41.589 106.045 -40.582 ;
      RECT 105.955 -41.065 106.095 -40.895 ;
      RECT 105.955 -40.168 106.045 -39.161 ;
      RECT 105.955 -39.855 106.095 -39.685 ;
      RECT 105.955 -38.359 106.045 -37.352 ;
      RECT 105.955 -37.835 106.095 -37.665 ;
      RECT 105.955 -36.938 106.045 -35.931 ;
      RECT 105.955 -36.625 106.095 -36.455 ;
      RECT 105.955 -35.129 106.045 -34.122 ;
      RECT 105.955 -34.605 106.095 -34.435 ;
      RECT 105.955 -33.708 106.045 -32.701 ;
      RECT 105.955 -33.395 106.095 -33.225 ;
      RECT 105.955 -31.899 106.045 -30.892 ;
      RECT 105.955 -31.375 106.095 -31.205 ;
      RECT 105.955 -30.478 106.045 -29.471 ;
      RECT 105.955 -30.165 106.095 -29.995 ;
      RECT 105.955 -28.669 106.045 -27.662 ;
      RECT 105.955 -28.145 106.095 -27.975 ;
      RECT 105.955 -27.248 106.045 -26.241 ;
      RECT 105.955 -26.935 106.095 -26.765 ;
      RECT 105.955 -25.439 106.045 -24.432 ;
      RECT 105.955 -24.915 106.095 -24.745 ;
      RECT 105.955 -24.018 106.045 -23.011 ;
      RECT 105.955 -23.705 106.095 -23.535 ;
      RECT 105.955 -22.209 106.045 -21.202 ;
      RECT 105.955 -21.685 106.095 -21.515 ;
      RECT 105.955 -20.788 106.045 -19.781 ;
      RECT 105.955 -20.475 106.095 -20.305 ;
      RECT 105.955 -18.979 106.045 -17.972 ;
      RECT 105.955 -18.455 106.095 -18.285 ;
      RECT 105.955 -17.558 106.045 -16.551 ;
      RECT 105.955 -17.245 106.095 -17.075 ;
      RECT 105.955 -15.749 106.045 -14.742 ;
      RECT 105.955 -15.225 106.095 -15.055 ;
      RECT 105.955 -14.328 106.045 -13.321 ;
      RECT 105.955 -14.015 106.095 -13.845 ;
      RECT 105.955 -12.519 106.045 -11.512 ;
      RECT 105.955 -11.995 106.095 -11.825 ;
      RECT 105.955 -11.098 106.045 -10.091 ;
      RECT 105.955 -10.785 106.095 -10.615 ;
      RECT 105.955 -9.289 106.045 -8.282 ;
      RECT 105.955 -8.765 106.095 -8.595 ;
      RECT 105.955 -7.868 106.045 -6.861 ;
      RECT 105.955 -7.555 106.095 -7.385 ;
      RECT 105.955 -6.059 106.045 -5.052 ;
      RECT 105.955 -5.535 106.095 -5.365 ;
      RECT 105.955 -4.638 106.045 -3.631 ;
      RECT 105.955 -4.325 106.095 -4.155 ;
      RECT 105.955 -2.829 106.045 -1.822 ;
      RECT 105.955 -2.305 106.095 -2.135 ;
      RECT 105.955 -1.408 106.045 -0.401 ;
      RECT 105.955 -1.095 106.095 -0.925 ;
      RECT 105.955 0.401 106.045 1.408 ;
      RECT 105.955 0.925 106.095 1.095 ;
      RECT 101.785 -108.935 105.565 -108.815 ;
      RECT 103.105 -109.475 103.205 -108.815 ;
      RECT 102.545 -109.475 102.645 -108.815 ;
      RECT 101.985 -109.475 102.085 -108.815 ;
      RECT 105.155 -101.538 105.245 -100.53 ;
      RECT 105.105 -100.935 105.245 -100.765 ;
      RECT 105.155 -99.73 105.245 -98.722 ;
      RECT 105.105 -99.495 105.245 -99.325 ;
      RECT 105.155 -98.308 105.245 -97.3 ;
      RECT 105.105 -97.705 105.245 -97.535 ;
      RECT 105.155 -96.5 105.245 -95.492 ;
      RECT 105.105 -96.265 105.245 -96.095 ;
      RECT 105.155 -95.078 105.245 -94.07 ;
      RECT 105.105 -94.475 105.245 -94.305 ;
      RECT 105.155 -93.27 105.245 -92.262 ;
      RECT 105.105 -93.035 105.245 -92.865 ;
      RECT 105.155 -91.848 105.245 -90.84 ;
      RECT 105.105 -91.245 105.245 -91.075 ;
      RECT 105.155 -90.04 105.245 -89.032 ;
      RECT 105.105 -89.805 105.245 -89.635 ;
      RECT 105.155 -88.618 105.245 -87.61 ;
      RECT 105.105 -88.015 105.245 -87.845 ;
      RECT 105.155 -86.81 105.245 -85.802 ;
      RECT 105.105 -86.575 105.245 -86.405 ;
      RECT 105.155 -85.388 105.245 -84.38 ;
      RECT 105.105 -84.785 105.245 -84.615 ;
      RECT 105.155 -83.58 105.245 -82.572 ;
      RECT 105.105 -83.345 105.245 -83.175 ;
      RECT 105.155 -82.158 105.245 -81.15 ;
      RECT 105.105 -81.555 105.245 -81.385 ;
      RECT 105.155 -80.35 105.245 -79.342 ;
      RECT 105.105 -80.115 105.245 -79.945 ;
      RECT 105.155 -78.928 105.245 -77.92 ;
      RECT 105.105 -78.325 105.245 -78.155 ;
      RECT 105.155 -77.12 105.245 -76.112 ;
      RECT 105.105 -76.885 105.245 -76.715 ;
      RECT 105.155 -75.698 105.245 -74.69 ;
      RECT 105.105 -75.095 105.245 -74.925 ;
      RECT 105.155 -73.89 105.245 -72.882 ;
      RECT 105.105 -73.655 105.245 -73.485 ;
      RECT 105.155 -72.468 105.245 -71.46 ;
      RECT 105.105 -71.865 105.245 -71.695 ;
      RECT 105.155 -70.66 105.245 -69.652 ;
      RECT 105.105 -70.425 105.245 -70.255 ;
      RECT 105.155 -69.238 105.245 -68.23 ;
      RECT 105.105 -68.635 105.245 -68.465 ;
      RECT 105.155 -67.43 105.245 -66.422 ;
      RECT 105.105 -67.195 105.245 -67.025 ;
      RECT 105.155 -66.008 105.245 -65 ;
      RECT 105.105 -65.405 105.245 -65.235 ;
      RECT 105.155 -64.2 105.245 -63.192 ;
      RECT 105.105 -63.965 105.245 -63.795 ;
      RECT 105.155 -62.778 105.245 -61.77 ;
      RECT 105.105 -62.175 105.245 -62.005 ;
      RECT 105.155 -60.97 105.245 -59.962 ;
      RECT 105.105 -60.735 105.245 -60.565 ;
      RECT 105.155 -59.548 105.245 -58.54 ;
      RECT 105.105 -58.945 105.245 -58.775 ;
      RECT 105.155 -57.74 105.245 -56.732 ;
      RECT 105.105 -57.505 105.245 -57.335 ;
      RECT 105.155 -56.318 105.245 -55.31 ;
      RECT 105.105 -55.715 105.245 -55.545 ;
      RECT 105.155 -54.51 105.245 -53.502 ;
      RECT 105.105 -54.275 105.245 -54.105 ;
      RECT 105.155 -53.088 105.245 -52.08 ;
      RECT 105.105 -52.485 105.245 -52.315 ;
      RECT 105.155 -51.28 105.245 -50.272 ;
      RECT 105.105 -51.045 105.245 -50.875 ;
      RECT 105.155 -49.858 105.245 -48.85 ;
      RECT 105.105 -49.255 105.245 -49.085 ;
      RECT 105.155 -48.05 105.245 -47.042 ;
      RECT 105.105 -47.815 105.245 -47.645 ;
      RECT 105.155 -46.628 105.245 -45.62 ;
      RECT 105.105 -46.025 105.245 -45.855 ;
      RECT 105.155 -44.82 105.245 -43.812 ;
      RECT 105.105 -44.585 105.245 -44.415 ;
      RECT 105.155 -43.398 105.245 -42.39 ;
      RECT 105.105 -42.795 105.245 -42.625 ;
      RECT 105.155 -41.59 105.245 -40.582 ;
      RECT 105.105 -41.355 105.245 -41.185 ;
      RECT 105.155 -40.168 105.245 -39.16 ;
      RECT 105.105 -39.565 105.245 -39.395 ;
      RECT 105.155 -38.36 105.245 -37.352 ;
      RECT 105.105 -38.125 105.245 -37.955 ;
      RECT 105.155 -36.938 105.245 -35.93 ;
      RECT 105.105 -36.335 105.245 -36.165 ;
      RECT 105.155 -35.13 105.245 -34.122 ;
      RECT 105.105 -34.895 105.245 -34.725 ;
      RECT 105.155 -33.708 105.245 -32.7 ;
      RECT 105.105 -33.105 105.245 -32.935 ;
      RECT 105.155 -31.9 105.245 -30.892 ;
      RECT 105.105 -31.665 105.245 -31.495 ;
      RECT 105.155 -30.478 105.245 -29.47 ;
      RECT 105.105 -29.875 105.245 -29.705 ;
      RECT 105.155 -28.67 105.245 -27.662 ;
      RECT 105.105 -28.435 105.245 -28.265 ;
      RECT 105.155 -27.248 105.245 -26.24 ;
      RECT 105.105 -26.645 105.245 -26.475 ;
      RECT 105.155 -25.44 105.245 -24.432 ;
      RECT 105.105 -25.205 105.245 -25.035 ;
      RECT 105.155 -24.018 105.245 -23.01 ;
      RECT 105.105 -23.415 105.245 -23.245 ;
      RECT 105.155 -22.21 105.245 -21.202 ;
      RECT 105.105 -21.975 105.245 -21.805 ;
      RECT 105.155 -20.788 105.245 -19.78 ;
      RECT 105.105 -20.185 105.245 -20.015 ;
      RECT 105.155 -18.98 105.245 -17.972 ;
      RECT 105.105 -18.745 105.245 -18.575 ;
      RECT 105.155 -17.558 105.245 -16.55 ;
      RECT 105.105 -16.955 105.245 -16.785 ;
      RECT 105.155 -15.75 105.245 -14.742 ;
      RECT 105.105 -15.515 105.245 -15.345 ;
      RECT 105.155 -14.328 105.245 -13.32 ;
      RECT 105.105 -13.725 105.245 -13.555 ;
      RECT 105.155 -12.52 105.245 -11.512 ;
      RECT 105.105 -12.285 105.245 -12.115 ;
      RECT 105.155 -11.098 105.245 -10.09 ;
      RECT 105.105 -10.495 105.245 -10.325 ;
      RECT 105.155 -9.29 105.245 -8.282 ;
      RECT 105.105 -9.055 105.245 -8.885 ;
      RECT 105.155 -7.868 105.245 -6.86 ;
      RECT 105.105 -7.265 105.245 -7.095 ;
      RECT 105.155 -6.06 105.245 -5.052 ;
      RECT 105.105 -5.825 105.245 -5.655 ;
      RECT 105.155 -4.638 105.245 -3.63 ;
      RECT 105.105 -4.035 105.245 -3.865 ;
      RECT 105.155 -2.83 105.245 -1.822 ;
      RECT 105.105 -2.595 105.245 -2.425 ;
      RECT 105.155 -1.408 105.245 -0.4 ;
      RECT 105.105 -0.805 105.245 -0.635 ;
      RECT 105.155 0.4 105.245 1.408 ;
      RECT 105.105 0.635 105.245 0.805 ;
      RECT 103.725 -111.685 105.205 -111.585 ;
      RECT 103.725 -112.195 103.825 -111.585 ;
      RECT 103.945 -109.15 105.205 -109.05 ;
      RECT 105.105 -109.475 105.205 -109.05 ;
      RECT 104.545 -109.475 104.645 -109.05 ;
      RECT 103.985 -109.475 104.085 -109.05 ;
      RECT 104.755 -101.538 104.845 -100.531 ;
      RECT 104.755 -101.225 104.895 -101.055 ;
      RECT 104.755 -99.729 104.845 -98.722 ;
      RECT 104.755 -99.205 104.895 -99.035 ;
      RECT 104.755 -98.308 104.845 -97.301 ;
      RECT 104.755 -97.995 104.895 -97.825 ;
      RECT 104.755 -96.499 104.845 -95.492 ;
      RECT 104.755 -95.975 104.895 -95.805 ;
      RECT 104.755 -95.078 104.845 -94.071 ;
      RECT 104.755 -94.765 104.895 -94.595 ;
      RECT 104.755 -93.269 104.845 -92.262 ;
      RECT 104.755 -92.745 104.895 -92.575 ;
      RECT 104.755 -91.848 104.845 -90.841 ;
      RECT 104.755 -91.535 104.895 -91.365 ;
      RECT 104.755 -90.039 104.845 -89.032 ;
      RECT 104.755 -89.515 104.895 -89.345 ;
      RECT 104.755 -88.618 104.845 -87.611 ;
      RECT 104.755 -88.305 104.895 -88.135 ;
      RECT 104.755 -86.809 104.845 -85.802 ;
      RECT 104.755 -86.285 104.895 -86.115 ;
      RECT 104.755 -85.388 104.845 -84.381 ;
      RECT 104.755 -85.075 104.895 -84.905 ;
      RECT 104.755 -83.579 104.845 -82.572 ;
      RECT 104.755 -83.055 104.895 -82.885 ;
      RECT 104.755 -82.158 104.845 -81.151 ;
      RECT 104.755 -81.845 104.895 -81.675 ;
      RECT 104.755 -80.349 104.845 -79.342 ;
      RECT 104.755 -79.825 104.895 -79.655 ;
      RECT 104.755 -78.928 104.845 -77.921 ;
      RECT 104.755 -78.615 104.895 -78.445 ;
      RECT 104.755 -77.119 104.845 -76.112 ;
      RECT 104.755 -76.595 104.895 -76.425 ;
      RECT 104.755 -75.698 104.845 -74.691 ;
      RECT 104.755 -75.385 104.895 -75.215 ;
      RECT 104.755 -73.889 104.845 -72.882 ;
      RECT 104.755 -73.365 104.895 -73.195 ;
      RECT 104.755 -72.468 104.845 -71.461 ;
      RECT 104.755 -72.155 104.895 -71.985 ;
      RECT 104.755 -70.659 104.845 -69.652 ;
      RECT 104.755 -70.135 104.895 -69.965 ;
      RECT 104.755 -69.238 104.845 -68.231 ;
      RECT 104.755 -68.925 104.895 -68.755 ;
      RECT 104.755 -67.429 104.845 -66.422 ;
      RECT 104.755 -66.905 104.895 -66.735 ;
      RECT 104.755 -66.008 104.845 -65.001 ;
      RECT 104.755 -65.695 104.895 -65.525 ;
      RECT 104.755 -64.199 104.845 -63.192 ;
      RECT 104.755 -63.675 104.895 -63.505 ;
      RECT 104.755 -62.778 104.845 -61.771 ;
      RECT 104.755 -62.465 104.895 -62.295 ;
      RECT 104.755 -60.969 104.845 -59.962 ;
      RECT 104.755 -60.445 104.895 -60.275 ;
      RECT 104.755 -59.548 104.845 -58.541 ;
      RECT 104.755 -59.235 104.895 -59.065 ;
      RECT 104.755 -57.739 104.845 -56.732 ;
      RECT 104.755 -57.215 104.895 -57.045 ;
      RECT 104.755 -56.318 104.845 -55.311 ;
      RECT 104.755 -56.005 104.895 -55.835 ;
      RECT 104.755 -54.509 104.845 -53.502 ;
      RECT 104.755 -53.985 104.895 -53.815 ;
      RECT 104.755 -53.088 104.845 -52.081 ;
      RECT 104.755 -52.775 104.895 -52.605 ;
      RECT 104.755 -51.279 104.845 -50.272 ;
      RECT 104.755 -50.755 104.895 -50.585 ;
      RECT 104.755 -49.858 104.845 -48.851 ;
      RECT 104.755 -49.545 104.895 -49.375 ;
      RECT 104.755 -48.049 104.845 -47.042 ;
      RECT 104.755 -47.525 104.895 -47.355 ;
      RECT 104.755 -46.628 104.845 -45.621 ;
      RECT 104.755 -46.315 104.895 -46.145 ;
      RECT 104.755 -44.819 104.845 -43.812 ;
      RECT 104.755 -44.295 104.895 -44.125 ;
      RECT 104.755 -43.398 104.845 -42.391 ;
      RECT 104.755 -43.085 104.895 -42.915 ;
      RECT 104.755 -41.589 104.845 -40.582 ;
      RECT 104.755 -41.065 104.895 -40.895 ;
      RECT 104.755 -40.168 104.845 -39.161 ;
      RECT 104.755 -39.855 104.895 -39.685 ;
      RECT 104.755 -38.359 104.845 -37.352 ;
      RECT 104.755 -37.835 104.895 -37.665 ;
      RECT 104.755 -36.938 104.845 -35.931 ;
      RECT 104.755 -36.625 104.895 -36.455 ;
      RECT 104.755 -35.129 104.845 -34.122 ;
      RECT 104.755 -34.605 104.895 -34.435 ;
      RECT 104.755 -33.708 104.845 -32.701 ;
      RECT 104.755 -33.395 104.895 -33.225 ;
      RECT 104.755 -31.899 104.845 -30.892 ;
      RECT 104.755 -31.375 104.895 -31.205 ;
      RECT 104.755 -30.478 104.845 -29.471 ;
      RECT 104.755 -30.165 104.895 -29.995 ;
      RECT 104.755 -28.669 104.845 -27.662 ;
      RECT 104.755 -28.145 104.895 -27.975 ;
      RECT 104.755 -27.248 104.845 -26.241 ;
      RECT 104.755 -26.935 104.895 -26.765 ;
      RECT 104.755 -25.439 104.845 -24.432 ;
      RECT 104.755 -24.915 104.895 -24.745 ;
      RECT 104.755 -24.018 104.845 -23.011 ;
      RECT 104.755 -23.705 104.895 -23.535 ;
      RECT 104.755 -22.209 104.845 -21.202 ;
      RECT 104.755 -21.685 104.895 -21.515 ;
      RECT 104.755 -20.788 104.845 -19.781 ;
      RECT 104.755 -20.475 104.895 -20.305 ;
      RECT 104.755 -18.979 104.845 -17.972 ;
      RECT 104.755 -18.455 104.895 -18.285 ;
      RECT 104.755 -17.558 104.845 -16.551 ;
      RECT 104.755 -17.245 104.895 -17.075 ;
      RECT 104.755 -15.749 104.845 -14.742 ;
      RECT 104.755 -15.225 104.895 -15.055 ;
      RECT 104.755 -14.328 104.845 -13.321 ;
      RECT 104.755 -14.015 104.895 -13.845 ;
      RECT 104.755 -12.519 104.845 -11.512 ;
      RECT 104.755 -11.995 104.895 -11.825 ;
      RECT 104.755 -11.098 104.845 -10.091 ;
      RECT 104.755 -10.785 104.895 -10.615 ;
      RECT 104.755 -9.289 104.845 -8.282 ;
      RECT 104.755 -8.765 104.895 -8.595 ;
      RECT 104.755 -7.868 104.845 -6.861 ;
      RECT 104.755 -7.555 104.895 -7.385 ;
      RECT 104.755 -6.059 104.845 -5.052 ;
      RECT 104.755 -5.535 104.895 -5.365 ;
      RECT 104.755 -4.638 104.845 -3.631 ;
      RECT 104.755 -4.325 104.895 -4.155 ;
      RECT 104.755 -2.829 104.845 -1.822 ;
      RECT 104.755 -2.305 104.895 -2.135 ;
      RECT 104.755 -1.408 104.845 -0.401 ;
      RECT 104.755 -1.095 104.895 -0.925 ;
      RECT 104.755 0.401 104.845 1.408 ;
      RECT 104.755 0.925 104.895 1.095 ;
      RECT 104.085 -111.495 104.255 -111.385 ;
      RECT 100.935 -111.495 104.255 -111.395 ;
      RECT 103.955 -101.538 104.045 -100.53 ;
      RECT 103.905 -100.935 104.045 -100.765 ;
      RECT 103.955 -99.73 104.045 -98.722 ;
      RECT 103.905 -99.495 104.045 -99.325 ;
      RECT 103.955 -98.308 104.045 -97.3 ;
      RECT 103.905 -97.705 104.045 -97.535 ;
      RECT 103.955 -96.5 104.045 -95.492 ;
      RECT 103.905 -96.265 104.045 -96.095 ;
      RECT 103.955 -95.078 104.045 -94.07 ;
      RECT 103.905 -94.475 104.045 -94.305 ;
      RECT 103.955 -93.27 104.045 -92.262 ;
      RECT 103.905 -93.035 104.045 -92.865 ;
      RECT 103.955 -91.848 104.045 -90.84 ;
      RECT 103.905 -91.245 104.045 -91.075 ;
      RECT 103.955 -90.04 104.045 -89.032 ;
      RECT 103.905 -89.805 104.045 -89.635 ;
      RECT 103.955 -88.618 104.045 -87.61 ;
      RECT 103.905 -88.015 104.045 -87.845 ;
      RECT 103.955 -86.81 104.045 -85.802 ;
      RECT 103.905 -86.575 104.045 -86.405 ;
      RECT 103.955 -85.388 104.045 -84.38 ;
      RECT 103.905 -84.785 104.045 -84.615 ;
      RECT 103.955 -83.58 104.045 -82.572 ;
      RECT 103.905 -83.345 104.045 -83.175 ;
      RECT 103.955 -82.158 104.045 -81.15 ;
      RECT 103.905 -81.555 104.045 -81.385 ;
      RECT 103.955 -80.35 104.045 -79.342 ;
      RECT 103.905 -80.115 104.045 -79.945 ;
      RECT 103.955 -78.928 104.045 -77.92 ;
      RECT 103.905 -78.325 104.045 -78.155 ;
      RECT 103.955 -77.12 104.045 -76.112 ;
      RECT 103.905 -76.885 104.045 -76.715 ;
      RECT 103.955 -75.698 104.045 -74.69 ;
      RECT 103.905 -75.095 104.045 -74.925 ;
      RECT 103.955 -73.89 104.045 -72.882 ;
      RECT 103.905 -73.655 104.045 -73.485 ;
      RECT 103.955 -72.468 104.045 -71.46 ;
      RECT 103.905 -71.865 104.045 -71.695 ;
      RECT 103.955 -70.66 104.045 -69.652 ;
      RECT 103.905 -70.425 104.045 -70.255 ;
      RECT 103.955 -69.238 104.045 -68.23 ;
      RECT 103.905 -68.635 104.045 -68.465 ;
      RECT 103.955 -67.43 104.045 -66.422 ;
      RECT 103.905 -67.195 104.045 -67.025 ;
      RECT 103.955 -66.008 104.045 -65 ;
      RECT 103.905 -65.405 104.045 -65.235 ;
      RECT 103.955 -64.2 104.045 -63.192 ;
      RECT 103.905 -63.965 104.045 -63.795 ;
      RECT 103.955 -62.778 104.045 -61.77 ;
      RECT 103.905 -62.175 104.045 -62.005 ;
      RECT 103.955 -60.97 104.045 -59.962 ;
      RECT 103.905 -60.735 104.045 -60.565 ;
      RECT 103.955 -59.548 104.045 -58.54 ;
      RECT 103.905 -58.945 104.045 -58.775 ;
      RECT 103.955 -57.74 104.045 -56.732 ;
      RECT 103.905 -57.505 104.045 -57.335 ;
      RECT 103.955 -56.318 104.045 -55.31 ;
      RECT 103.905 -55.715 104.045 -55.545 ;
      RECT 103.955 -54.51 104.045 -53.502 ;
      RECT 103.905 -54.275 104.045 -54.105 ;
      RECT 103.955 -53.088 104.045 -52.08 ;
      RECT 103.905 -52.485 104.045 -52.315 ;
      RECT 103.955 -51.28 104.045 -50.272 ;
      RECT 103.905 -51.045 104.045 -50.875 ;
      RECT 103.955 -49.858 104.045 -48.85 ;
      RECT 103.905 -49.255 104.045 -49.085 ;
      RECT 103.955 -48.05 104.045 -47.042 ;
      RECT 103.905 -47.815 104.045 -47.645 ;
      RECT 103.955 -46.628 104.045 -45.62 ;
      RECT 103.905 -46.025 104.045 -45.855 ;
      RECT 103.955 -44.82 104.045 -43.812 ;
      RECT 103.905 -44.585 104.045 -44.415 ;
      RECT 103.955 -43.398 104.045 -42.39 ;
      RECT 103.905 -42.795 104.045 -42.625 ;
      RECT 103.955 -41.59 104.045 -40.582 ;
      RECT 103.905 -41.355 104.045 -41.185 ;
      RECT 103.955 -40.168 104.045 -39.16 ;
      RECT 103.905 -39.565 104.045 -39.395 ;
      RECT 103.955 -38.36 104.045 -37.352 ;
      RECT 103.905 -38.125 104.045 -37.955 ;
      RECT 103.955 -36.938 104.045 -35.93 ;
      RECT 103.905 -36.335 104.045 -36.165 ;
      RECT 103.955 -35.13 104.045 -34.122 ;
      RECT 103.905 -34.895 104.045 -34.725 ;
      RECT 103.955 -33.708 104.045 -32.7 ;
      RECT 103.905 -33.105 104.045 -32.935 ;
      RECT 103.955 -31.9 104.045 -30.892 ;
      RECT 103.905 -31.665 104.045 -31.495 ;
      RECT 103.955 -30.478 104.045 -29.47 ;
      RECT 103.905 -29.875 104.045 -29.705 ;
      RECT 103.955 -28.67 104.045 -27.662 ;
      RECT 103.905 -28.435 104.045 -28.265 ;
      RECT 103.955 -27.248 104.045 -26.24 ;
      RECT 103.905 -26.645 104.045 -26.475 ;
      RECT 103.955 -25.44 104.045 -24.432 ;
      RECT 103.905 -25.205 104.045 -25.035 ;
      RECT 103.955 -24.018 104.045 -23.01 ;
      RECT 103.905 -23.415 104.045 -23.245 ;
      RECT 103.955 -22.21 104.045 -21.202 ;
      RECT 103.905 -21.975 104.045 -21.805 ;
      RECT 103.955 -20.788 104.045 -19.78 ;
      RECT 103.905 -20.185 104.045 -20.015 ;
      RECT 103.955 -18.98 104.045 -17.972 ;
      RECT 103.905 -18.745 104.045 -18.575 ;
      RECT 103.955 -17.558 104.045 -16.55 ;
      RECT 103.905 -16.955 104.045 -16.785 ;
      RECT 103.955 -15.75 104.045 -14.742 ;
      RECT 103.905 -15.515 104.045 -15.345 ;
      RECT 103.955 -14.328 104.045 -13.32 ;
      RECT 103.905 -13.725 104.045 -13.555 ;
      RECT 103.955 -12.52 104.045 -11.512 ;
      RECT 103.905 -12.285 104.045 -12.115 ;
      RECT 103.955 -11.098 104.045 -10.09 ;
      RECT 103.905 -10.495 104.045 -10.325 ;
      RECT 103.955 -9.29 104.045 -8.282 ;
      RECT 103.905 -9.055 104.045 -8.885 ;
      RECT 103.955 -7.868 104.045 -6.86 ;
      RECT 103.905 -7.265 104.045 -7.095 ;
      RECT 103.955 -6.06 104.045 -5.052 ;
      RECT 103.905 -5.825 104.045 -5.655 ;
      RECT 103.955 -4.638 104.045 -3.63 ;
      RECT 103.905 -4.035 104.045 -3.865 ;
      RECT 103.955 -2.83 104.045 -1.822 ;
      RECT 103.905 -2.595 104.045 -2.425 ;
      RECT 103.955 -1.408 104.045 -0.4 ;
      RECT 103.905 -0.805 104.045 -0.635 ;
      RECT 103.955 0.4 104.045 1.408 ;
      RECT 103.905 0.635 104.045 0.805 ;
      RECT 103.555 -101.538 103.645 -100.531 ;
      RECT 103.555 -101.225 103.695 -101.055 ;
      RECT 103.555 -99.729 103.645 -98.722 ;
      RECT 103.555 -99.205 103.695 -99.035 ;
      RECT 103.555 -98.308 103.645 -97.301 ;
      RECT 103.555 -97.995 103.695 -97.825 ;
      RECT 103.555 -96.499 103.645 -95.492 ;
      RECT 103.555 -95.975 103.695 -95.805 ;
      RECT 103.555 -95.078 103.645 -94.071 ;
      RECT 103.555 -94.765 103.695 -94.595 ;
      RECT 103.555 -93.269 103.645 -92.262 ;
      RECT 103.555 -92.745 103.695 -92.575 ;
      RECT 103.555 -91.848 103.645 -90.841 ;
      RECT 103.555 -91.535 103.695 -91.365 ;
      RECT 103.555 -90.039 103.645 -89.032 ;
      RECT 103.555 -89.515 103.695 -89.345 ;
      RECT 103.555 -88.618 103.645 -87.611 ;
      RECT 103.555 -88.305 103.695 -88.135 ;
      RECT 103.555 -86.809 103.645 -85.802 ;
      RECT 103.555 -86.285 103.695 -86.115 ;
      RECT 103.555 -85.388 103.645 -84.381 ;
      RECT 103.555 -85.075 103.695 -84.905 ;
      RECT 103.555 -83.579 103.645 -82.572 ;
      RECT 103.555 -83.055 103.695 -82.885 ;
      RECT 103.555 -82.158 103.645 -81.151 ;
      RECT 103.555 -81.845 103.695 -81.675 ;
      RECT 103.555 -80.349 103.645 -79.342 ;
      RECT 103.555 -79.825 103.695 -79.655 ;
      RECT 103.555 -78.928 103.645 -77.921 ;
      RECT 103.555 -78.615 103.695 -78.445 ;
      RECT 103.555 -77.119 103.645 -76.112 ;
      RECT 103.555 -76.595 103.695 -76.425 ;
      RECT 103.555 -75.698 103.645 -74.691 ;
      RECT 103.555 -75.385 103.695 -75.215 ;
      RECT 103.555 -73.889 103.645 -72.882 ;
      RECT 103.555 -73.365 103.695 -73.195 ;
      RECT 103.555 -72.468 103.645 -71.461 ;
      RECT 103.555 -72.155 103.695 -71.985 ;
      RECT 103.555 -70.659 103.645 -69.652 ;
      RECT 103.555 -70.135 103.695 -69.965 ;
      RECT 103.555 -69.238 103.645 -68.231 ;
      RECT 103.555 -68.925 103.695 -68.755 ;
      RECT 103.555 -67.429 103.645 -66.422 ;
      RECT 103.555 -66.905 103.695 -66.735 ;
      RECT 103.555 -66.008 103.645 -65.001 ;
      RECT 103.555 -65.695 103.695 -65.525 ;
      RECT 103.555 -64.199 103.645 -63.192 ;
      RECT 103.555 -63.675 103.695 -63.505 ;
      RECT 103.555 -62.778 103.645 -61.771 ;
      RECT 103.555 -62.465 103.695 -62.295 ;
      RECT 103.555 -60.969 103.645 -59.962 ;
      RECT 103.555 -60.445 103.695 -60.275 ;
      RECT 103.555 -59.548 103.645 -58.541 ;
      RECT 103.555 -59.235 103.695 -59.065 ;
      RECT 103.555 -57.739 103.645 -56.732 ;
      RECT 103.555 -57.215 103.695 -57.045 ;
      RECT 103.555 -56.318 103.645 -55.311 ;
      RECT 103.555 -56.005 103.695 -55.835 ;
      RECT 103.555 -54.509 103.645 -53.502 ;
      RECT 103.555 -53.985 103.695 -53.815 ;
      RECT 103.555 -53.088 103.645 -52.081 ;
      RECT 103.555 -52.775 103.695 -52.605 ;
      RECT 103.555 -51.279 103.645 -50.272 ;
      RECT 103.555 -50.755 103.695 -50.585 ;
      RECT 103.555 -49.858 103.645 -48.851 ;
      RECT 103.555 -49.545 103.695 -49.375 ;
      RECT 103.555 -48.049 103.645 -47.042 ;
      RECT 103.555 -47.525 103.695 -47.355 ;
      RECT 103.555 -46.628 103.645 -45.621 ;
      RECT 103.555 -46.315 103.695 -46.145 ;
      RECT 103.555 -44.819 103.645 -43.812 ;
      RECT 103.555 -44.295 103.695 -44.125 ;
      RECT 103.555 -43.398 103.645 -42.391 ;
      RECT 103.555 -43.085 103.695 -42.915 ;
      RECT 103.555 -41.589 103.645 -40.582 ;
      RECT 103.555 -41.065 103.695 -40.895 ;
      RECT 103.555 -40.168 103.645 -39.161 ;
      RECT 103.555 -39.855 103.695 -39.685 ;
      RECT 103.555 -38.359 103.645 -37.352 ;
      RECT 103.555 -37.835 103.695 -37.665 ;
      RECT 103.555 -36.938 103.645 -35.931 ;
      RECT 103.555 -36.625 103.695 -36.455 ;
      RECT 103.555 -35.129 103.645 -34.122 ;
      RECT 103.555 -34.605 103.695 -34.435 ;
      RECT 103.555 -33.708 103.645 -32.701 ;
      RECT 103.555 -33.395 103.695 -33.225 ;
      RECT 103.555 -31.899 103.645 -30.892 ;
      RECT 103.555 -31.375 103.695 -31.205 ;
      RECT 103.555 -30.478 103.645 -29.471 ;
      RECT 103.555 -30.165 103.695 -29.995 ;
      RECT 103.555 -28.669 103.645 -27.662 ;
      RECT 103.555 -28.145 103.695 -27.975 ;
      RECT 103.555 -27.248 103.645 -26.241 ;
      RECT 103.555 -26.935 103.695 -26.765 ;
      RECT 103.555 -25.439 103.645 -24.432 ;
      RECT 103.555 -24.915 103.695 -24.745 ;
      RECT 103.555 -24.018 103.645 -23.011 ;
      RECT 103.555 -23.705 103.695 -23.535 ;
      RECT 103.555 -22.209 103.645 -21.202 ;
      RECT 103.555 -21.685 103.695 -21.515 ;
      RECT 103.555 -20.788 103.645 -19.781 ;
      RECT 103.555 -20.475 103.695 -20.305 ;
      RECT 103.555 -18.979 103.645 -17.972 ;
      RECT 103.555 -18.455 103.695 -18.285 ;
      RECT 103.555 -17.558 103.645 -16.551 ;
      RECT 103.555 -17.245 103.695 -17.075 ;
      RECT 103.555 -15.749 103.645 -14.742 ;
      RECT 103.555 -15.225 103.695 -15.055 ;
      RECT 103.555 -14.328 103.645 -13.321 ;
      RECT 103.555 -14.015 103.695 -13.845 ;
      RECT 103.555 -12.519 103.645 -11.512 ;
      RECT 103.555 -11.995 103.695 -11.825 ;
      RECT 103.555 -11.098 103.645 -10.091 ;
      RECT 103.555 -10.785 103.695 -10.615 ;
      RECT 103.555 -9.289 103.645 -8.282 ;
      RECT 103.555 -8.765 103.695 -8.595 ;
      RECT 103.555 -7.868 103.645 -6.861 ;
      RECT 103.555 -7.555 103.695 -7.385 ;
      RECT 103.555 -6.059 103.645 -5.052 ;
      RECT 103.555 -5.535 103.695 -5.365 ;
      RECT 103.555 -4.638 103.645 -3.631 ;
      RECT 103.555 -4.325 103.695 -4.155 ;
      RECT 103.555 -2.829 103.645 -1.822 ;
      RECT 103.555 -2.305 103.695 -2.135 ;
      RECT 103.555 -1.408 103.645 -0.401 ;
      RECT 103.555 -1.095 103.695 -0.925 ;
      RECT 103.555 0.401 103.645 1.408 ;
      RECT 103.555 0.925 103.695 1.095 ;
      RECT 101.705 -111.685 103.185 -111.585 ;
      RECT 101.705 -112.055 101.805 -111.585 ;
      RECT 101.51 -114.395 103.085 -114.275 ;
      RECT 102.985 -114.895 103.085 -114.275 ;
      RECT 102.39 -114.895 102.49 -114.275 ;
      RECT 101.51 -114.85 101.61 -114.275 ;
      RECT 102.755 -101.538 102.845 -100.53 ;
      RECT 102.705 -100.935 102.845 -100.765 ;
      RECT 102.755 -99.73 102.845 -98.722 ;
      RECT 102.705 -99.495 102.845 -99.325 ;
      RECT 102.755 -98.308 102.845 -97.3 ;
      RECT 102.705 -97.705 102.845 -97.535 ;
      RECT 102.755 -96.5 102.845 -95.492 ;
      RECT 102.705 -96.265 102.845 -96.095 ;
      RECT 102.755 -95.078 102.845 -94.07 ;
      RECT 102.705 -94.475 102.845 -94.305 ;
      RECT 102.755 -93.27 102.845 -92.262 ;
      RECT 102.705 -93.035 102.845 -92.865 ;
      RECT 102.755 -91.848 102.845 -90.84 ;
      RECT 102.705 -91.245 102.845 -91.075 ;
      RECT 102.755 -90.04 102.845 -89.032 ;
      RECT 102.705 -89.805 102.845 -89.635 ;
      RECT 102.755 -88.618 102.845 -87.61 ;
      RECT 102.705 -88.015 102.845 -87.845 ;
      RECT 102.755 -86.81 102.845 -85.802 ;
      RECT 102.705 -86.575 102.845 -86.405 ;
      RECT 102.755 -85.388 102.845 -84.38 ;
      RECT 102.705 -84.785 102.845 -84.615 ;
      RECT 102.755 -83.58 102.845 -82.572 ;
      RECT 102.705 -83.345 102.845 -83.175 ;
      RECT 102.755 -82.158 102.845 -81.15 ;
      RECT 102.705 -81.555 102.845 -81.385 ;
      RECT 102.755 -80.35 102.845 -79.342 ;
      RECT 102.705 -80.115 102.845 -79.945 ;
      RECT 102.755 -78.928 102.845 -77.92 ;
      RECT 102.705 -78.325 102.845 -78.155 ;
      RECT 102.755 -77.12 102.845 -76.112 ;
      RECT 102.705 -76.885 102.845 -76.715 ;
      RECT 102.755 -75.698 102.845 -74.69 ;
      RECT 102.705 -75.095 102.845 -74.925 ;
      RECT 102.755 -73.89 102.845 -72.882 ;
      RECT 102.705 -73.655 102.845 -73.485 ;
      RECT 102.755 -72.468 102.845 -71.46 ;
      RECT 102.705 -71.865 102.845 -71.695 ;
      RECT 102.755 -70.66 102.845 -69.652 ;
      RECT 102.705 -70.425 102.845 -70.255 ;
      RECT 102.755 -69.238 102.845 -68.23 ;
      RECT 102.705 -68.635 102.845 -68.465 ;
      RECT 102.755 -67.43 102.845 -66.422 ;
      RECT 102.705 -67.195 102.845 -67.025 ;
      RECT 102.755 -66.008 102.845 -65 ;
      RECT 102.705 -65.405 102.845 -65.235 ;
      RECT 102.755 -64.2 102.845 -63.192 ;
      RECT 102.705 -63.965 102.845 -63.795 ;
      RECT 102.755 -62.778 102.845 -61.77 ;
      RECT 102.705 -62.175 102.845 -62.005 ;
      RECT 102.755 -60.97 102.845 -59.962 ;
      RECT 102.705 -60.735 102.845 -60.565 ;
      RECT 102.755 -59.548 102.845 -58.54 ;
      RECT 102.705 -58.945 102.845 -58.775 ;
      RECT 102.755 -57.74 102.845 -56.732 ;
      RECT 102.705 -57.505 102.845 -57.335 ;
      RECT 102.755 -56.318 102.845 -55.31 ;
      RECT 102.705 -55.715 102.845 -55.545 ;
      RECT 102.755 -54.51 102.845 -53.502 ;
      RECT 102.705 -54.275 102.845 -54.105 ;
      RECT 102.755 -53.088 102.845 -52.08 ;
      RECT 102.705 -52.485 102.845 -52.315 ;
      RECT 102.755 -51.28 102.845 -50.272 ;
      RECT 102.705 -51.045 102.845 -50.875 ;
      RECT 102.755 -49.858 102.845 -48.85 ;
      RECT 102.705 -49.255 102.845 -49.085 ;
      RECT 102.755 -48.05 102.845 -47.042 ;
      RECT 102.705 -47.815 102.845 -47.645 ;
      RECT 102.755 -46.628 102.845 -45.62 ;
      RECT 102.705 -46.025 102.845 -45.855 ;
      RECT 102.755 -44.82 102.845 -43.812 ;
      RECT 102.705 -44.585 102.845 -44.415 ;
      RECT 102.755 -43.398 102.845 -42.39 ;
      RECT 102.705 -42.795 102.845 -42.625 ;
      RECT 102.755 -41.59 102.845 -40.582 ;
      RECT 102.705 -41.355 102.845 -41.185 ;
      RECT 102.755 -40.168 102.845 -39.16 ;
      RECT 102.705 -39.565 102.845 -39.395 ;
      RECT 102.755 -38.36 102.845 -37.352 ;
      RECT 102.705 -38.125 102.845 -37.955 ;
      RECT 102.755 -36.938 102.845 -35.93 ;
      RECT 102.705 -36.335 102.845 -36.165 ;
      RECT 102.755 -35.13 102.845 -34.122 ;
      RECT 102.705 -34.895 102.845 -34.725 ;
      RECT 102.755 -33.708 102.845 -32.7 ;
      RECT 102.705 -33.105 102.845 -32.935 ;
      RECT 102.755 -31.9 102.845 -30.892 ;
      RECT 102.705 -31.665 102.845 -31.495 ;
      RECT 102.755 -30.478 102.845 -29.47 ;
      RECT 102.705 -29.875 102.845 -29.705 ;
      RECT 102.755 -28.67 102.845 -27.662 ;
      RECT 102.705 -28.435 102.845 -28.265 ;
      RECT 102.755 -27.248 102.845 -26.24 ;
      RECT 102.705 -26.645 102.845 -26.475 ;
      RECT 102.755 -25.44 102.845 -24.432 ;
      RECT 102.705 -25.205 102.845 -25.035 ;
      RECT 102.755 -24.018 102.845 -23.01 ;
      RECT 102.705 -23.415 102.845 -23.245 ;
      RECT 102.755 -22.21 102.845 -21.202 ;
      RECT 102.705 -21.975 102.845 -21.805 ;
      RECT 102.755 -20.788 102.845 -19.78 ;
      RECT 102.705 -20.185 102.845 -20.015 ;
      RECT 102.755 -18.98 102.845 -17.972 ;
      RECT 102.705 -18.745 102.845 -18.575 ;
      RECT 102.755 -17.558 102.845 -16.55 ;
      RECT 102.705 -16.955 102.845 -16.785 ;
      RECT 102.755 -15.75 102.845 -14.742 ;
      RECT 102.705 -15.515 102.845 -15.345 ;
      RECT 102.755 -14.328 102.845 -13.32 ;
      RECT 102.705 -13.725 102.845 -13.555 ;
      RECT 102.755 -12.52 102.845 -11.512 ;
      RECT 102.705 -12.285 102.845 -12.115 ;
      RECT 102.755 -11.098 102.845 -10.09 ;
      RECT 102.705 -10.495 102.845 -10.325 ;
      RECT 102.755 -9.29 102.845 -8.282 ;
      RECT 102.705 -9.055 102.845 -8.885 ;
      RECT 102.755 -7.868 102.845 -6.86 ;
      RECT 102.705 -7.265 102.845 -7.095 ;
      RECT 102.755 -6.06 102.845 -5.052 ;
      RECT 102.705 -5.825 102.845 -5.655 ;
      RECT 102.755 -4.638 102.845 -3.63 ;
      RECT 102.705 -4.035 102.845 -3.865 ;
      RECT 102.755 -2.83 102.845 -1.822 ;
      RECT 102.705 -2.595 102.845 -2.425 ;
      RECT 102.755 -1.408 102.845 -0.4 ;
      RECT 102.705 -0.805 102.845 -0.635 ;
      RECT 102.755 0.4 102.845 1.408 ;
      RECT 102.705 0.635 102.845 0.805 ;
      RECT 102.63 -114.685 102.805 -114.515 ;
      RECT 102.705 -114.895 102.805 -114.515 ;
      RECT 101.745 -113.555 101.845 -113.09 ;
      RECT 102.11 -113.555 102.21 -113.1 ;
      RECT 101.745 -113.555 102.59 -113.385 ;
      RECT 102.355 -101.538 102.445 -100.531 ;
      RECT 102.355 -101.225 102.495 -101.055 ;
      RECT 102.355 -99.729 102.445 -98.722 ;
      RECT 102.355 -99.205 102.495 -99.035 ;
      RECT 102.355 -98.308 102.445 -97.301 ;
      RECT 102.355 -97.995 102.495 -97.825 ;
      RECT 102.355 -96.499 102.445 -95.492 ;
      RECT 102.355 -95.975 102.495 -95.805 ;
      RECT 102.355 -95.078 102.445 -94.071 ;
      RECT 102.355 -94.765 102.495 -94.595 ;
      RECT 102.355 -93.269 102.445 -92.262 ;
      RECT 102.355 -92.745 102.495 -92.575 ;
      RECT 102.355 -91.848 102.445 -90.841 ;
      RECT 102.355 -91.535 102.495 -91.365 ;
      RECT 102.355 -90.039 102.445 -89.032 ;
      RECT 102.355 -89.515 102.495 -89.345 ;
      RECT 102.355 -88.618 102.445 -87.611 ;
      RECT 102.355 -88.305 102.495 -88.135 ;
      RECT 102.355 -86.809 102.445 -85.802 ;
      RECT 102.355 -86.285 102.495 -86.115 ;
      RECT 102.355 -85.388 102.445 -84.381 ;
      RECT 102.355 -85.075 102.495 -84.905 ;
      RECT 102.355 -83.579 102.445 -82.572 ;
      RECT 102.355 -83.055 102.495 -82.885 ;
      RECT 102.355 -82.158 102.445 -81.151 ;
      RECT 102.355 -81.845 102.495 -81.675 ;
      RECT 102.355 -80.349 102.445 -79.342 ;
      RECT 102.355 -79.825 102.495 -79.655 ;
      RECT 102.355 -78.928 102.445 -77.921 ;
      RECT 102.355 -78.615 102.495 -78.445 ;
      RECT 102.355 -77.119 102.445 -76.112 ;
      RECT 102.355 -76.595 102.495 -76.425 ;
      RECT 102.355 -75.698 102.445 -74.691 ;
      RECT 102.355 -75.385 102.495 -75.215 ;
      RECT 102.355 -73.889 102.445 -72.882 ;
      RECT 102.355 -73.365 102.495 -73.195 ;
      RECT 102.355 -72.468 102.445 -71.461 ;
      RECT 102.355 -72.155 102.495 -71.985 ;
      RECT 102.355 -70.659 102.445 -69.652 ;
      RECT 102.355 -70.135 102.495 -69.965 ;
      RECT 102.355 -69.238 102.445 -68.231 ;
      RECT 102.355 -68.925 102.495 -68.755 ;
      RECT 102.355 -67.429 102.445 -66.422 ;
      RECT 102.355 -66.905 102.495 -66.735 ;
      RECT 102.355 -66.008 102.445 -65.001 ;
      RECT 102.355 -65.695 102.495 -65.525 ;
      RECT 102.355 -64.199 102.445 -63.192 ;
      RECT 102.355 -63.675 102.495 -63.505 ;
      RECT 102.355 -62.778 102.445 -61.771 ;
      RECT 102.355 -62.465 102.495 -62.295 ;
      RECT 102.355 -60.969 102.445 -59.962 ;
      RECT 102.355 -60.445 102.495 -60.275 ;
      RECT 102.355 -59.548 102.445 -58.541 ;
      RECT 102.355 -59.235 102.495 -59.065 ;
      RECT 102.355 -57.739 102.445 -56.732 ;
      RECT 102.355 -57.215 102.495 -57.045 ;
      RECT 102.355 -56.318 102.445 -55.311 ;
      RECT 102.355 -56.005 102.495 -55.835 ;
      RECT 102.355 -54.509 102.445 -53.502 ;
      RECT 102.355 -53.985 102.495 -53.815 ;
      RECT 102.355 -53.088 102.445 -52.081 ;
      RECT 102.355 -52.775 102.495 -52.605 ;
      RECT 102.355 -51.279 102.445 -50.272 ;
      RECT 102.355 -50.755 102.495 -50.585 ;
      RECT 102.355 -49.858 102.445 -48.851 ;
      RECT 102.355 -49.545 102.495 -49.375 ;
      RECT 102.355 -48.049 102.445 -47.042 ;
      RECT 102.355 -47.525 102.495 -47.355 ;
      RECT 102.355 -46.628 102.445 -45.621 ;
      RECT 102.355 -46.315 102.495 -46.145 ;
      RECT 102.355 -44.819 102.445 -43.812 ;
      RECT 102.355 -44.295 102.495 -44.125 ;
      RECT 102.355 -43.398 102.445 -42.391 ;
      RECT 102.355 -43.085 102.495 -42.915 ;
      RECT 102.355 -41.589 102.445 -40.582 ;
      RECT 102.355 -41.065 102.495 -40.895 ;
      RECT 102.355 -40.168 102.445 -39.161 ;
      RECT 102.355 -39.855 102.495 -39.685 ;
      RECT 102.355 -38.359 102.445 -37.352 ;
      RECT 102.355 -37.835 102.495 -37.665 ;
      RECT 102.355 -36.938 102.445 -35.931 ;
      RECT 102.355 -36.625 102.495 -36.455 ;
      RECT 102.355 -35.129 102.445 -34.122 ;
      RECT 102.355 -34.605 102.495 -34.435 ;
      RECT 102.355 -33.708 102.445 -32.701 ;
      RECT 102.355 -33.395 102.495 -33.225 ;
      RECT 102.355 -31.899 102.445 -30.892 ;
      RECT 102.355 -31.375 102.495 -31.205 ;
      RECT 102.355 -30.478 102.445 -29.471 ;
      RECT 102.355 -30.165 102.495 -29.995 ;
      RECT 102.355 -28.669 102.445 -27.662 ;
      RECT 102.355 -28.145 102.495 -27.975 ;
      RECT 102.355 -27.248 102.445 -26.241 ;
      RECT 102.355 -26.935 102.495 -26.765 ;
      RECT 102.355 -25.439 102.445 -24.432 ;
      RECT 102.355 -24.915 102.495 -24.745 ;
      RECT 102.355 -24.018 102.445 -23.011 ;
      RECT 102.355 -23.705 102.495 -23.535 ;
      RECT 102.355 -22.209 102.445 -21.202 ;
      RECT 102.355 -21.685 102.495 -21.515 ;
      RECT 102.355 -20.788 102.445 -19.781 ;
      RECT 102.355 -20.475 102.495 -20.305 ;
      RECT 102.355 -18.979 102.445 -17.972 ;
      RECT 102.355 -18.455 102.495 -18.285 ;
      RECT 102.355 -17.558 102.445 -16.551 ;
      RECT 102.355 -17.245 102.495 -17.075 ;
      RECT 102.355 -15.749 102.445 -14.742 ;
      RECT 102.355 -15.225 102.495 -15.055 ;
      RECT 102.355 -14.328 102.445 -13.321 ;
      RECT 102.355 -14.015 102.495 -13.845 ;
      RECT 102.355 -12.519 102.445 -11.512 ;
      RECT 102.355 -11.995 102.495 -11.825 ;
      RECT 102.355 -11.098 102.445 -10.091 ;
      RECT 102.355 -10.785 102.495 -10.615 ;
      RECT 102.355 -9.289 102.445 -8.282 ;
      RECT 102.355 -8.765 102.495 -8.595 ;
      RECT 102.355 -7.868 102.445 -6.861 ;
      RECT 102.355 -7.555 102.495 -7.385 ;
      RECT 102.355 -6.059 102.445 -5.052 ;
      RECT 102.355 -5.535 102.495 -5.365 ;
      RECT 102.355 -4.638 102.445 -3.631 ;
      RECT 102.355 -4.325 102.495 -4.155 ;
      RECT 102.355 -2.829 102.445 -1.822 ;
      RECT 102.355 -2.305 102.495 -2.135 ;
      RECT 102.355 -1.408 102.445 -0.401 ;
      RECT 102.355 -1.095 102.495 -0.925 ;
      RECT 102.355 0.401 102.445 1.408 ;
      RECT 102.355 0.925 102.495 1.095 ;
      RECT 102.04 -114.685 102.21 -114.515 ;
      RECT 102.11 -114.895 102.21 -114.515 ;
      RECT 101.555 -101.538 101.645 -100.53 ;
      RECT 101.505 -100.935 101.645 -100.765 ;
      RECT 101.555 -99.73 101.645 -98.722 ;
      RECT 101.505 -99.495 101.645 -99.325 ;
      RECT 101.555 -98.308 101.645 -97.3 ;
      RECT 101.505 -97.705 101.645 -97.535 ;
      RECT 101.555 -96.5 101.645 -95.492 ;
      RECT 101.505 -96.265 101.645 -96.095 ;
      RECT 101.555 -95.078 101.645 -94.07 ;
      RECT 101.505 -94.475 101.645 -94.305 ;
      RECT 101.555 -93.27 101.645 -92.262 ;
      RECT 101.505 -93.035 101.645 -92.865 ;
      RECT 101.555 -91.848 101.645 -90.84 ;
      RECT 101.505 -91.245 101.645 -91.075 ;
      RECT 101.555 -90.04 101.645 -89.032 ;
      RECT 101.505 -89.805 101.645 -89.635 ;
      RECT 101.555 -88.618 101.645 -87.61 ;
      RECT 101.505 -88.015 101.645 -87.845 ;
      RECT 101.555 -86.81 101.645 -85.802 ;
      RECT 101.505 -86.575 101.645 -86.405 ;
      RECT 101.555 -85.388 101.645 -84.38 ;
      RECT 101.505 -84.785 101.645 -84.615 ;
      RECT 101.555 -83.58 101.645 -82.572 ;
      RECT 101.505 -83.345 101.645 -83.175 ;
      RECT 101.555 -82.158 101.645 -81.15 ;
      RECT 101.505 -81.555 101.645 -81.385 ;
      RECT 101.555 -80.35 101.645 -79.342 ;
      RECT 101.505 -80.115 101.645 -79.945 ;
      RECT 101.555 -78.928 101.645 -77.92 ;
      RECT 101.505 -78.325 101.645 -78.155 ;
      RECT 101.555 -77.12 101.645 -76.112 ;
      RECT 101.505 -76.885 101.645 -76.715 ;
      RECT 101.555 -75.698 101.645 -74.69 ;
      RECT 101.505 -75.095 101.645 -74.925 ;
      RECT 101.555 -73.89 101.645 -72.882 ;
      RECT 101.505 -73.655 101.645 -73.485 ;
      RECT 101.555 -72.468 101.645 -71.46 ;
      RECT 101.505 -71.865 101.645 -71.695 ;
      RECT 101.555 -70.66 101.645 -69.652 ;
      RECT 101.505 -70.425 101.645 -70.255 ;
      RECT 101.555 -69.238 101.645 -68.23 ;
      RECT 101.505 -68.635 101.645 -68.465 ;
      RECT 101.555 -67.43 101.645 -66.422 ;
      RECT 101.505 -67.195 101.645 -67.025 ;
      RECT 101.555 -66.008 101.645 -65 ;
      RECT 101.505 -65.405 101.645 -65.235 ;
      RECT 101.555 -64.2 101.645 -63.192 ;
      RECT 101.505 -63.965 101.645 -63.795 ;
      RECT 101.555 -62.778 101.645 -61.77 ;
      RECT 101.505 -62.175 101.645 -62.005 ;
      RECT 101.555 -60.97 101.645 -59.962 ;
      RECT 101.505 -60.735 101.645 -60.565 ;
      RECT 101.555 -59.548 101.645 -58.54 ;
      RECT 101.505 -58.945 101.645 -58.775 ;
      RECT 101.555 -57.74 101.645 -56.732 ;
      RECT 101.505 -57.505 101.645 -57.335 ;
      RECT 101.555 -56.318 101.645 -55.31 ;
      RECT 101.505 -55.715 101.645 -55.545 ;
      RECT 101.555 -54.51 101.645 -53.502 ;
      RECT 101.505 -54.275 101.645 -54.105 ;
      RECT 101.555 -53.088 101.645 -52.08 ;
      RECT 101.505 -52.485 101.645 -52.315 ;
      RECT 101.555 -51.28 101.645 -50.272 ;
      RECT 101.505 -51.045 101.645 -50.875 ;
      RECT 101.555 -49.858 101.645 -48.85 ;
      RECT 101.505 -49.255 101.645 -49.085 ;
      RECT 101.555 -48.05 101.645 -47.042 ;
      RECT 101.505 -47.815 101.645 -47.645 ;
      RECT 101.555 -46.628 101.645 -45.62 ;
      RECT 101.505 -46.025 101.645 -45.855 ;
      RECT 101.555 -44.82 101.645 -43.812 ;
      RECT 101.505 -44.585 101.645 -44.415 ;
      RECT 101.555 -43.398 101.645 -42.39 ;
      RECT 101.505 -42.795 101.645 -42.625 ;
      RECT 101.555 -41.59 101.645 -40.582 ;
      RECT 101.505 -41.355 101.645 -41.185 ;
      RECT 101.555 -40.168 101.645 -39.16 ;
      RECT 101.505 -39.565 101.645 -39.395 ;
      RECT 101.555 -38.36 101.645 -37.352 ;
      RECT 101.505 -38.125 101.645 -37.955 ;
      RECT 101.555 -36.938 101.645 -35.93 ;
      RECT 101.505 -36.335 101.645 -36.165 ;
      RECT 101.555 -35.13 101.645 -34.122 ;
      RECT 101.505 -34.895 101.645 -34.725 ;
      RECT 101.555 -33.708 101.645 -32.7 ;
      RECT 101.505 -33.105 101.645 -32.935 ;
      RECT 101.555 -31.9 101.645 -30.892 ;
      RECT 101.505 -31.665 101.645 -31.495 ;
      RECT 101.555 -30.478 101.645 -29.47 ;
      RECT 101.505 -29.875 101.645 -29.705 ;
      RECT 101.555 -28.67 101.645 -27.662 ;
      RECT 101.505 -28.435 101.645 -28.265 ;
      RECT 101.555 -27.248 101.645 -26.24 ;
      RECT 101.505 -26.645 101.645 -26.475 ;
      RECT 101.555 -25.44 101.645 -24.432 ;
      RECT 101.505 -25.205 101.645 -25.035 ;
      RECT 101.555 -24.018 101.645 -23.01 ;
      RECT 101.505 -23.415 101.645 -23.245 ;
      RECT 101.555 -22.21 101.645 -21.202 ;
      RECT 101.505 -21.975 101.645 -21.805 ;
      RECT 101.555 -20.788 101.645 -19.78 ;
      RECT 101.505 -20.185 101.645 -20.015 ;
      RECT 101.555 -18.98 101.645 -17.972 ;
      RECT 101.505 -18.745 101.645 -18.575 ;
      RECT 101.555 -17.558 101.645 -16.55 ;
      RECT 101.505 -16.955 101.645 -16.785 ;
      RECT 101.555 -15.75 101.645 -14.742 ;
      RECT 101.505 -15.515 101.645 -15.345 ;
      RECT 101.555 -14.328 101.645 -13.32 ;
      RECT 101.505 -13.725 101.645 -13.555 ;
      RECT 101.555 -12.52 101.645 -11.512 ;
      RECT 101.505 -12.285 101.645 -12.115 ;
      RECT 101.555 -11.098 101.645 -10.09 ;
      RECT 101.505 -10.495 101.645 -10.325 ;
      RECT 101.555 -9.29 101.645 -8.282 ;
      RECT 101.505 -9.055 101.645 -8.885 ;
      RECT 101.555 -7.868 101.645 -6.86 ;
      RECT 101.505 -7.265 101.645 -7.095 ;
      RECT 101.555 -6.06 101.645 -5.052 ;
      RECT 101.505 -5.825 101.645 -5.655 ;
      RECT 101.555 -4.638 101.645 -3.63 ;
      RECT 101.505 -4.035 101.645 -3.865 ;
      RECT 101.555 -2.83 101.645 -1.822 ;
      RECT 101.505 -2.595 101.645 -2.425 ;
      RECT 101.555 -1.408 101.645 -0.4 ;
      RECT 101.505 -0.805 101.645 -0.635 ;
      RECT 101.555 0.4 101.645 1.408 ;
      RECT 101.505 0.635 101.645 0.805 ;
      RECT 101.155 -101.538 101.245 -100.531 ;
      RECT 101.155 -101.225 101.295 -101.055 ;
      RECT 101.155 -99.729 101.245 -98.722 ;
      RECT 101.155 -99.205 101.295 -99.035 ;
      RECT 101.155 -98.308 101.245 -97.301 ;
      RECT 101.155 -97.995 101.295 -97.825 ;
      RECT 101.155 -96.499 101.245 -95.492 ;
      RECT 101.155 -95.975 101.295 -95.805 ;
      RECT 101.155 -95.078 101.245 -94.071 ;
      RECT 101.155 -94.765 101.295 -94.595 ;
      RECT 101.155 -93.269 101.245 -92.262 ;
      RECT 101.155 -92.745 101.295 -92.575 ;
      RECT 101.155 -91.848 101.245 -90.841 ;
      RECT 101.155 -91.535 101.295 -91.365 ;
      RECT 101.155 -90.039 101.245 -89.032 ;
      RECT 101.155 -89.515 101.295 -89.345 ;
      RECT 101.155 -88.618 101.245 -87.611 ;
      RECT 101.155 -88.305 101.295 -88.135 ;
      RECT 101.155 -86.809 101.245 -85.802 ;
      RECT 101.155 -86.285 101.295 -86.115 ;
      RECT 101.155 -85.388 101.245 -84.381 ;
      RECT 101.155 -85.075 101.295 -84.905 ;
      RECT 101.155 -83.579 101.245 -82.572 ;
      RECT 101.155 -83.055 101.295 -82.885 ;
      RECT 101.155 -82.158 101.245 -81.151 ;
      RECT 101.155 -81.845 101.295 -81.675 ;
      RECT 101.155 -80.349 101.245 -79.342 ;
      RECT 101.155 -79.825 101.295 -79.655 ;
      RECT 101.155 -78.928 101.245 -77.921 ;
      RECT 101.155 -78.615 101.295 -78.445 ;
      RECT 101.155 -77.119 101.245 -76.112 ;
      RECT 101.155 -76.595 101.295 -76.425 ;
      RECT 101.155 -75.698 101.245 -74.691 ;
      RECT 101.155 -75.385 101.295 -75.215 ;
      RECT 101.155 -73.889 101.245 -72.882 ;
      RECT 101.155 -73.365 101.295 -73.195 ;
      RECT 101.155 -72.468 101.245 -71.461 ;
      RECT 101.155 -72.155 101.295 -71.985 ;
      RECT 101.155 -70.659 101.245 -69.652 ;
      RECT 101.155 -70.135 101.295 -69.965 ;
      RECT 101.155 -69.238 101.245 -68.231 ;
      RECT 101.155 -68.925 101.295 -68.755 ;
      RECT 101.155 -67.429 101.245 -66.422 ;
      RECT 101.155 -66.905 101.295 -66.735 ;
      RECT 101.155 -66.008 101.245 -65.001 ;
      RECT 101.155 -65.695 101.295 -65.525 ;
      RECT 101.155 -64.199 101.245 -63.192 ;
      RECT 101.155 -63.675 101.295 -63.505 ;
      RECT 101.155 -62.778 101.245 -61.771 ;
      RECT 101.155 -62.465 101.295 -62.295 ;
      RECT 101.155 -60.969 101.245 -59.962 ;
      RECT 101.155 -60.445 101.295 -60.275 ;
      RECT 101.155 -59.548 101.245 -58.541 ;
      RECT 101.155 -59.235 101.295 -59.065 ;
      RECT 101.155 -57.739 101.245 -56.732 ;
      RECT 101.155 -57.215 101.295 -57.045 ;
      RECT 101.155 -56.318 101.245 -55.311 ;
      RECT 101.155 -56.005 101.295 -55.835 ;
      RECT 101.155 -54.509 101.245 -53.502 ;
      RECT 101.155 -53.985 101.295 -53.815 ;
      RECT 101.155 -53.088 101.245 -52.081 ;
      RECT 101.155 -52.775 101.295 -52.605 ;
      RECT 101.155 -51.279 101.245 -50.272 ;
      RECT 101.155 -50.755 101.295 -50.585 ;
      RECT 101.155 -49.858 101.245 -48.851 ;
      RECT 101.155 -49.545 101.295 -49.375 ;
      RECT 101.155 -48.049 101.245 -47.042 ;
      RECT 101.155 -47.525 101.295 -47.355 ;
      RECT 101.155 -46.628 101.245 -45.621 ;
      RECT 101.155 -46.315 101.295 -46.145 ;
      RECT 101.155 -44.819 101.245 -43.812 ;
      RECT 101.155 -44.295 101.295 -44.125 ;
      RECT 101.155 -43.398 101.245 -42.391 ;
      RECT 101.155 -43.085 101.295 -42.915 ;
      RECT 101.155 -41.589 101.245 -40.582 ;
      RECT 101.155 -41.065 101.295 -40.895 ;
      RECT 101.155 -40.168 101.245 -39.161 ;
      RECT 101.155 -39.855 101.295 -39.685 ;
      RECT 101.155 -38.359 101.245 -37.352 ;
      RECT 101.155 -37.835 101.295 -37.665 ;
      RECT 101.155 -36.938 101.245 -35.931 ;
      RECT 101.155 -36.625 101.295 -36.455 ;
      RECT 101.155 -35.129 101.245 -34.122 ;
      RECT 101.155 -34.605 101.295 -34.435 ;
      RECT 101.155 -33.708 101.245 -32.701 ;
      RECT 101.155 -33.395 101.295 -33.225 ;
      RECT 101.155 -31.899 101.245 -30.892 ;
      RECT 101.155 -31.375 101.295 -31.205 ;
      RECT 101.155 -30.478 101.245 -29.471 ;
      RECT 101.155 -30.165 101.295 -29.995 ;
      RECT 101.155 -28.669 101.245 -27.662 ;
      RECT 101.155 -28.145 101.295 -27.975 ;
      RECT 101.155 -27.248 101.245 -26.241 ;
      RECT 101.155 -26.935 101.295 -26.765 ;
      RECT 101.155 -25.439 101.245 -24.432 ;
      RECT 101.155 -24.915 101.295 -24.745 ;
      RECT 101.155 -24.018 101.245 -23.011 ;
      RECT 101.155 -23.705 101.295 -23.535 ;
      RECT 101.155 -22.209 101.245 -21.202 ;
      RECT 101.155 -21.685 101.295 -21.515 ;
      RECT 101.155 -20.788 101.245 -19.781 ;
      RECT 101.155 -20.475 101.295 -20.305 ;
      RECT 101.155 -18.979 101.245 -17.972 ;
      RECT 101.155 -18.455 101.295 -18.285 ;
      RECT 101.155 -17.558 101.245 -16.551 ;
      RECT 101.155 -17.245 101.295 -17.075 ;
      RECT 101.155 -15.749 101.245 -14.742 ;
      RECT 101.155 -15.225 101.295 -15.055 ;
      RECT 101.155 -14.328 101.245 -13.321 ;
      RECT 101.155 -14.015 101.295 -13.845 ;
      RECT 101.155 -12.519 101.245 -11.512 ;
      RECT 101.155 -11.995 101.295 -11.825 ;
      RECT 101.155 -11.098 101.245 -10.091 ;
      RECT 101.155 -10.785 101.295 -10.615 ;
      RECT 101.155 -9.289 101.245 -8.282 ;
      RECT 101.155 -8.765 101.295 -8.595 ;
      RECT 101.155 -7.868 101.245 -6.861 ;
      RECT 101.155 -7.555 101.295 -7.385 ;
      RECT 101.155 -6.059 101.245 -5.052 ;
      RECT 101.155 -5.535 101.295 -5.365 ;
      RECT 101.155 -4.638 101.245 -3.631 ;
      RECT 101.155 -4.325 101.295 -4.155 ;
      RECT 101.155 -2.829 101.245 -1.822 ;
      RECT 101.155 -2.305 101.295 -2.135 ;
      RECT 101.155 -1.408 101.245 -0.401 ;
      RECT 101.155 -1.095 101.295 -0.925 ;
      RECT 101.155 0.401 101.245 1.408 ;
      RECT 101.155 0.925 101.295 1.095 ;
      RECT 96.985 -108.935 100.765 -108.815 ;
      RECT 98.305 -109.475 98.405 -108.815 ;
      RECT 97.745 -109.475 97.845 -108.815 ;
      RECT 97.185 -109.475 97.285 -108.815 ;
      RECT 100.355 -101.538 100.445 -100.53 ;
      RECT 100.305 -100.935 100.445 -100.765 ;
      RECT 100.355 -99.73 100.445 -98.722 ;
      RECT 100.305 -99.495 100.445 -99.325 ;
      RECT 100.355 -98.308 100.445 -97.3 ;
      RECT 100.305 -97.705 100.445 -97.535 ;
      RECT 100.355 -96.5 100.445 -95.492 ;
      RECT 100.305 -96.265 100.445 -96.095 ;
      RECT 100.355 -95.078 100.445 -94.07 ;
      RECT 100.305 -94.475 100.445 -94.305 ;
      RECT 100.355 -93.27 100.445 -92.262 ;
      RECT 100.305 -93.035 100.445 -92.865 ;
      RECT 100.355 -91.848 100.445 -90.84 ;
      RECT 100.305 -91.245 100.445 -91.075 ;
      RECT 100.355 -90.04 100.445 -89.032 ;
      RECT 100.305 -89.805 100.445 -89.635 ;
      RECT 100.355 -88.618 100.445 -87.61 ;
      RECT 100.305 -88.015 100.445 -87.845 ;
      RECT 100.355 -86.81 100.445 -85.802 ;
      RECT 100.305 -86.575 100.445 -86.405 ;
      RECT 100.355 -85.388 100.445 -84.38 ;
      RECT 100.305 -84.785 100.445 -84.615 ;
      RECT 100.355 -83.58 100.445 -82.572 ;
      RECT 100.305 -83.345 100.445 -83.175 ;
      RECT 100.355 -82.158 100.445 -81.15 ;
      RECT 100.305 -81.555 100.445 -81.385 ;
      RECT 100.355 -80.35 100.445 -79.342 ;
      RECT 100.305 -80.115 100.445 -79.945 ;
      RECT 100.355 -78.928 100.445 -77.92 ;
      RECT 100.305 -78.325 100.445 -78.155 ;
      RECT 100.355 -77.12 100.445 -76.112 ;
      RECT 100.305 -76.885 100.445 -76.715 ;
      RECT 100.355 -75.698 100.445 -74.69 ;
      RECT 100.305 -75.095 100.445 -74.925 ;
      RECT 100.355 -73.89 100.445 -72.882 ;
      RECT 100.305 -73.655 100.445 -73.485 ;
      RECT 100.355 -72.468 100.445 -71.46 ;
      RECT 100.305 -71.865 100.445 -71.695 ;
      RECT 100.355 -70.66 100.445 -69.652 ;
      RECT 100.305 -70.425 100.445 -70.255 ;
      RECT 100.355 -69.238 100.445 -68.23 ;
      RECT 100.305 -68.635 100.445 -68.465 ;
      RECT 100.355 -67.43 100.445 -66.422 ;
      RECT 100.305 -67.195 100.445 -67.025 ;
      RECT 100.355 -66.008 100.445 -65 ;
      RECT 100.305 -65.405 100.445 -65.235 ;
      RECT 100.355 -64.2 100.445 -63.192 ;
      RECT 100.305 -63.965 100.445 -63.795 ;
      RECT 100.355 -62.778 100.445 -61.77 ;
      RECT 100.305 -62.175 100.445 -62.005 ;
      RECT 100.355 -60.97 100.445 -59.962 ;
      RECT 100.305 -60.735 100.445 -60.565 ;
      RECT 100.355 -59.548 100.445 -58.54 ;
      RECT 100.305 -58.945 100.445 -58.775 ;
      RECT 100.355 -57.74 100.445 -56.732 ;
      RECT 100.305 -57.505 100.445 -57.335 ;
      RECT 100.355 -56.318 100.445 -55.31 ;
      RECT 100.305 -55.715 100.445 -55.545 ;
      RECT 100.355 -54.51 100.445 -53.502 ;
      RECT 100.305 -54.275 100.445 -54.105 ;
      RECT 100.355 -53.088 100.445 -52.08 ;
      RECT 100.305 -52.485 100.445 -52.315 ;
      RECT 100.355 -51.28 100.445 -50.272 ;
      RECT 100.305 -51.045 100.445 -50.875 ;
      RECT 100.355 -49.858 100.445 -48.85 ;
      RECT 100.305 -49.255 100.445 -49.085 ;
      RECT 100.355 -48.05 100.445 -47.042 ;
      RECT 100.305 -47.815 100.445 -47.645 ;
      RECT 100.355 -46.628 100.445 -45.62 ;
      RECT 100.305 -46.025 100.445 -45.855 ;
      RECT 100.355 -44.82 100.445 -43.812 ;
      RECT 100.305 -44.585 100.445 -44.415 ;
      RECT 100.355 -43.398 100.445 -42.39 ;
      RECT 100.305 -42.795 100.445 -42.625 ;
      RECT 100.355 -41.59 100.445 -40.582 ;
      RECT 100.305 -41.355 100.445 -41.185 ;
      RECT 100.355 -40.168 100.445 -39.16 ;
      RECT 100.305 -39.565 100.445 -39.395 ;
      RECT 100.355 -38.36 100.445 -37.352 ;
      RECT 100.305 -38.125 100.445 -37.955 ;
      RECT 100.355 -36.938 100.445 -35.93 ;
      RECT 100.305 -36.335 100.445 -36.165 ;
      RECT 100.355 -35.13 100.445 -34.122 ;
      RECT 100.305 -34.895 100.445 -34.725 ;
      RECT 100.355 -33.708 100.445 -32.7 ;
      RECT 100.305 -33.105 100.445 -32.935 ;
      RECT 100.355 -31.9 100.445 -30.892 ;
      RECT 100.305 -31.665 100.445 -31.495 ;
      RECT 100.355 -30.478 100.445 -29.47 ;
      RECT 100.305 -29.875 100.445 -29.705 ;
      RECT 100.355 -28.67 100.445 -27.662 ;
      RECT 100.305 -28.435 100.445 -28.265 ;
      RECT 100.355 -27.248 100.445 -26.24 ;
      RECT 100.305 -26.645 100.445 -26.475 ;
      RECT 100.355 -25.44 100.445 -24.432 ;
      RECT 100.305 -25.205 100.445 -25.035 ;
      RECT 100.355 -24.018 100.445 -23.01 ;
      RECT 100.305 -23.415 100.445 -23.245 ;
      RECT 100.355 -22.21 100.445 -21.202 ;
      RECT 100.305 -21.975 100.445 -21.805 ;
      RECT 100.355 -20.788 100.445 -19.78 ;
      RECT 100.305 -20.185 100.445 -20.015 ;
      RECT 100.355 -18.98 100.445 -17.972 ;
      RECT 100.305 -18.745 100.445 -18.575 ;
      RECT 100.355 -17.558 100.445 -16.55 ;
      RECT 100.305 -16.955 100.445 -16.785 ;
      RECT 100.355 -15.75 100.445 -14.742 ;
      RECT 100.305 -15.515 100.445 -15.345 ;
      RECT 100.355 -14.328 100.445 -13.32 ;
      RECT 100.305 -13.725 100.445 -13.555 ;
      RECT 100.355 -12.52 100.445 -11.512 ;
      RECT 100.305 -12.285 100.445 -12.115 ;
      RECT 100.355 -11.098 100.445 -10.09 ;
      RECT 100.305 -10.495 100.445 -10.325 ;
      RECT 100.355 -9.29 100.445 -8.282 ;
      RECT 100.305 -9.055 100.445 -8.885 ;
      RECT 100.355 -7.868 100.445 -6.86 ;
      RECT 100.305 -7.265 100.445 -7.095 ;
      RECT 100.355 -6.06 100.445 -5.052 ;
      RECT 100.305 -5.825 100.445 -5.655 ;
      RECT 100.355 -4.638 100.445 -3.63 ;
      RECT 100.305 -4.035 100.445 -3.865 ;
      RECT 100.355 -2.83 100.445 -1.822 ;
      RECT 100.305 -2.595 100.445 -2.425 ;
      RECT 100.355 -1.408 100.445 -0.4 ;
      RECT 100.305 -0.805 100.445 -0.635 ;
      RECT 100.355 0.4 100.445 1.408 ;
      RECT 100.305 0.635 100.445 0.805 ;
      RECT 98.925 -111.685 100.405 -111.585 ;
      RECT 98.925 -112.195 99.025 -111.585 ;
      RECT 99.145 -109.15 100.405 -109.05 ;
      RECT 100.305 -109.475 100.405 -109.05 ;
      RECT 99.745 -109.475 99.845 -109.05 ;
      RECT 99.185 -109.475 99.285 -109.05 ;
      RECT 99.955 -101.538 100.045 -100.531 ;
      RECT 99.955 -101.225 100.095 -101.055 ;
      RECT 99.955 -99.729 100.045 -98.722 ;
      RECT 99.955 -99.205 100.095 -99.035 ;
      RECT 99.955 -98.308 100.045 -97.301 ;
      RECT 99.955 -97.995 100.095 -97.825 ;
      RECT 99.955 -96.499 100.045 -95.492 ;
      RECT 99.955 -95.975 100.095 -95.805 ;
      RECT 99.955 -95.078 100.045 -94.071 ;
      RECT 99.955 -94.765 100.095 -94.595 ;
      RECT 99.955 -93.269 100.045 -92.262 ;
      RECT 99.955 -92.745 100.095 -92.575 ;
      RECT 99.955 -91.848 100.045 -90.841 ;
      RECT 99.955 -91.535 100.095 -91.365 ;
      RECT 99.955 -90.039 100.045 -89.032 ;
      RECT 99.955 -89.515 100.095 -89.345 ;
      RECT 99.955 -88.618 100.045 -87.611 ;
      RECT 99.955 -88.305 100.095 -88.135 ;
      RECT 99.955 -86.809 100.045 -85.802 ;
      RECT 99.955 -86.285 100.095 -86.115 ;
      RECT 99.955 -85.388 100.045 -84.381 ;
      RECT 99.955 -85.075 100.095 -84.905 ;
      RECT 99.955 -83.579 100.045 -82.572 ;
      RECT 99.955 -83.055 100.095 -82.885 ;
      RECT 99.955 -82.158 100.045 -81.151 ;
      RECT 99.955 -81.845 100.095 -81.675 ;
      RECT 99.955 -80.349 100.045 -79.342 ;
      RECT 99.955 -79.825 100.095 -79.655 ;
      RECT 99.955 -78.928 100.045 -77.921 ;
      RECT 99.955 -78.615 100.095 -78.445 ;
      RECT 99.955 -77.119 100.045 -76.112 ;
      RECT 99.955 -76.595 100.095 -76.425 ;
      RECT 99.955 -75.698 100.045 -74.691 ;
      RECT 99.955 -75.385 100.095 -75.215 ;
      RECT 99.955 -73.889 100.045 -72.882 ;
      RECT 99.955 -73.365 100.095 -73.195 ;
      RECT 99.955 -72.468 100.045 -71.461 ;
      RECT 99.955 -72.155 100.095 -71.985 ;
      RECT 99.955 -70.659 100.045 -69.652 ;
      RECT 99.955 -70.135 100.095 -69.965 ;
      RECT 99.955 -69.238 100.045 -68.231 ;
      RECT 99.955 -68.925 100.095 -68.755 ;
      RECT 99.955 -67.429 100.045 -66.422 ;
      RECT 99.955 -66.905 100.095 -66.735 ;
      RECT 99.955 -66.008 100.045 -65.001 ;
      RECT 99.955 -65.695 100.095 -65.525 ;
      RECT 99.955 -64.199 100.045 -63.192 ;
      RECT 99.955 -63.675 100.095 -63.505 ;
      RECT 99.955 -62.778 100.045 -61.771 ;
      RECT 99.955 -62.465 100.095 -62.295 ;
      RECT 99.955 -60.969 100.045 -59.962 ;
      RECT 99.955 -60.445 100.095 -60.275 ;
      RECT 99.955 -59.548 100.045 -58.541 ;
      RECT 99.955 -59.235 100.095 -59.065 ;
      RECT 99.955 -57.739 100.045 -56.732 ;
      RECT 99.955 -57.215 100.095 -57.045 ;
      RECT 99.955 -56.318 100.045 -55.311 ;
      RECT 99.955 -56.005 100.095 -55.835 ;
      RECT 99.955 -54.509 100.045 -53.502 ;
      RECT 99.955 -53.985 100.095 -53.815 ;
      RECT 99.955 -53.088 100.045 -52.081 ;
      RECT 99.955 -52.775 100.095 -52.605 ;
      RECT 99.955 -51.279 100.045 -50.272 ;
      RECT 99.955 -50.755 100.095 -50.585 ;
      RECT 99.955 -49.858 100.045 -48.851 ;
      RECT 99.955 -49.545 100.095 -49.375 ;
      RECT 99.955 -48.049 100.045 -47.042 ;
      RECT 99.955 -47.525 100.095 -47.355 ;
      RECT 99.955 -46.628 100.045 -45.621 ;
      RECT 99.955 -46.315 100.095 -46.145 ;
      RECT 99.955 -44.819 100.045 -43.812 ;
      RECT 99.955 -44.295 100.095 -44.125 ;
      RECT 99.955 -43.398 100.045 -42.391 ;
      RECT 99.955 -43.085 100.095 -42.915 ;
      RECT 99.955 -41.589 100.045 -40.582 ;
      RECT 99.955 -41.065 100.095 -40.895 ;
      RECT 99.955 -40.168 100.045 -39.161 ;
      RECT 99.955 -39.855 100.095 -39.685 ;
      RECT 99.955 -38.359 100.045 -37.352 ;
      RECT 99.955 -37.835 100.095 -37.665 ;
      RECT 99.955 -36.938 100.045 -35.931 ;
      RECT 99.955 -36.625 100.095 -36.455 ;
      RECT 99.955 -35.129 100.045 -34.122 ;
      RECT 99.955 -34.605 100.095 -34.435 ;
      RECT 99.955 -33.708 100.045 -32.701 ;
      RECT 99.955 -33.395 100.095 -33.225 ;
      RECT 99.955 -31.899 100.045 -30.892 ;
      RECT 99.955 -31.375 100.095 -31.205 ;
      RECT 99.955 -30.478 100.045 -29.471 ;
      RECT 99.955 -30.165 100.095 -29.995 ;
      RECT 99.955 -28.669 100.045 -27.662 ;
      RECT 99.955 -28.145 100.095 -27.975 ;
      RECT 99.955 -27.248 100.045 -26.241 ;
      RECT 99.955 -26.935 100.095 -26.765 ;
      RECT 99.955 -25.439 100.045 -24.432 ;
      RECT 99.955 -24.915 100.095 -24.745 ;
      RECT 99.955 -24.018 100.045 -23.011 ;
      RECT 99.955 -23.705 100.095 -23.535 ;
      RECT 99.955 -22.209 100.045 -21.202 ;
      RECT 99.955 -21.685 100.095 -21.515 ;
      RECT 99.955 -20.788 100.045 -19.781 ;
      RECT 99.955 -20.475 100.095 -20.305 ;
      RECT 99.955 -18.979 100.045 -17.972 ;
      RECT 99.955 -18.455 100.095 -18.285 ;
      RECT 99.955 -17.558 100.045 -16.551 ;
      RECT 99.955 -17.245 100.095 -17.075 ;
      RECT 99.955 -15.749 100.045 -14.742 ;
      RECT 99.955 -15.225 100.095 -15.055 ;
      RECT 99.955 -14.328 100.045 -13.321 ;
      RECT 99.955 -14.015 100.095 -13.845 ;
      RECT 99.955 -12.519 100.045 -11.512 ;
      RECT 99.955 -11.995 100.095 -11.825 ;
      RECT 99.955 -11.098 100.045 -10.091 ;
      RECT 99.955 -10.785 100.095 -10.615 ;
      RECT 99.955 -9.289 100.045 -8.282 ;
      RECT 99.955 -8.765 100.095 -8.595 ;
      RECT 99.955 -7.868 100.045 -6.861 ;
      RECT 99.955 -7.555 100.095 -7.385 ;
      RECT 99.955 -6.059 100.045 -5.052 ;
      RECT 99.955 -5.535 100.095 -5.365 ;
      RECT 99.955 -4.638 100.045 -3.631 ;
      RECT 99.955 -4.325 100.095 -4.155 ;
      RECT 99.955 -2.829 100.045 -1.822 ;
      RECT 99.955 -2.305 100.095 -2.135 ;
      RECT 99.955 -1.408 100.045 -0.401 ;
      RECT 99.955 -1.095 100.095 -0.925 ;
      RECT 99.955 0.401 100.045 1.408 ;
      RECT 99.955 0.925 100.095 1.095 ;
      RECT 99.285 -111.495 99.455 -111.385 ;
      RECT 96.135 -111.495 99.455 -111.395 ;
      RECT 99.155 -101.538 99.245 -100.53 ;
      RECT 99.105 -100.935 99.245 -100.765 ;
      RECT 99.155 -99.73 99.245 -98.722 ;
      RECT 99.105 -99.495 99.245 -99.325 ;
      RECT 99.155 -98.308 99.245 -97.3 ;
      RECT 99.105 -97.705 99.245 -97.535 ;
      RECT 99.155 -96.5 99.245 -95.492 ;
      RECT 99.105 -96.265 99.245 -96.095 ;
      RECT 99.155 -95.078 99.245 -94.07 ;
      RECT 99.105 -94.475 99.245 -94.305 ;
      RECT 99.155 -93.27 99.245 -92.262 ;
      RECT 99.105 -93.035 99.245 -92.865 ;
      RECT 99.155 -91.848 99.245 -90.84 ;
      RECT 99.105 -91.245 99.245 -91.075 ;
      RECT 99.155 -90.04 99.245 -89.032 ;
      RECT 99.105 -89.805 99.245 -89.635 ;
      RECT 99.155 -88.618 99.245 -87.61 ;
      RECT 99.105 -88.015 99.245 -87.845 ;
      RECT 99.155 -86.81 99.245 -85.802 ;
      RECT 99.105 -86.575 99.245 -86.405 ;
      RECT 99.155 -85.388 99.245 -84.38 ;
      RECT 99.105 -84.785 99.245 -84.615 ;
      RECT 99.155 -83.58 99.245 -82.572 ;
      RECT 99.105 -83.345 99.245 -83.175 ;
      RECT 99.155 -82.158 99.245 -81.15 ;
      RECT 99.105 -81.555 99.245 -81.385 ;
      RECT 99.155 -80.35 99.245 -79.342 ;
      RECT 99.105 -80.115 99.245 -79.945 ;
      RECT 99.155 -78.928 99.245 -77.92 ;
      RECT 99.105 -78.325 99.245 -78.155 ;
      RECT 99.155 -77.12 99.245 -76.112 ;
      RECT 99.105 -76.885 99.245 -76.715 ;
      RECT 99.155 -75.698 99.245 -74.69 ;
      RECT 99.105 -75.095 99.245 -74.925 ;
      RECT 99.155 -73.89 99.245 -72.882 ;
      RECT 99.105 -73.655 99.245 -73.485 ;
      RECT 99.155 -72.468 99.245 -71.46 ;
      RECT 99.105 -71.865 99.245 -71.695 ;
      RECT 99.155 -70.66 99.245 -69.652 ;
      RECT 99.105 -70.425 99.245 -70.255 ;
      RECT 99.155 -69.238 99.245 -68.23 ;
      RECT 99.105 -68.635 99.245 -68.465 ;
      RECT 99.155 -67.43 99.245 -66.422 ;
      RECT 99.105 -67.195 99.245 -67.025 ;
      RECT 99.155 -66.008 99.245 -65 ;
      RECT 99.105 -65.405 99.245 -65.235 ;
      RECT 99.155 -64.2 99.245 -63.192 ;
      RECT 99.105 -63.965 99.245 -63.795 ;
      RECT 99.155 -62.778 99.245 -61.77 ;
      RECT 99.105 -62.175 99.245 -62.005 ;
      RECT 99.155 -60.97 99.245 -59.962 ;
      RECT 99.105 -60.735 99.245 -60.565 ;
      RECT 99.155 -59.548 99.245 -58.54 ;
      RECT 99.105 -58.945 99.245 -58.775 ;
      RECT 99.155 -57.74 99.245 -56.732 ;
      RECT 99.105 -57.505 99.245 -57.335 ;
      RECT 99.155 -56.318 99.245 -55.31 ;
      RECT 99.105 -55.715 99.245 -55.545 ;
      RECT 99.155 -54.51 99.245 -53.502 ;
      RECT 99.105 -54.275 99.245 -54.105 ;
      RECT 99.155 -53.088 99.245 -52.08 ;
      RECT 99.105 -52.485 99.245 -52.315 ;
      RECT 99.155 -51.28 99.245 -50.272 ;
      RECT 99.105 -51.045 99.245 -50.875 ;
      RECT 99.155 -49.858 99.245 -48.85 ;
      RECT 99.105 -49.255 99.245 -49.085 ;
      RECT 99.155 -48.05 99.245 -47.042 ;
      RECT 99.105 -47.815 99.245 -47.645 ;
      RECT 99.155 -46.628 99.245 -45.62 ;
      RECT 99.105 -46.025 99.245 -45.855 ;
      RECT 99.155 -44.82 99.245 -43.812 ;
      RECT 99.105 -44.585 99.245 -44.415 ;
      RECT 99.155 -43.398 99.245 -42.39 ;
      RECT 99.105 -42.795 99.245 -42.625 ;
      RECT 99.155 -41.59 99.245 -40.582 ;
      RECT 99.105 -41.355 99.245 -41.185 ;
      RECT 99.155 -40.168 99.245 -39.16 ;
      RECT 99.105 -39.565 99.245 -39.395 ;
      RECT 99.155 -38.36 99.245 -37.352 ;
      RECT 99.105 -38.125 99.245 -37.955 ;
      RECT 99.155 -36.938 99.245 -35.93 ;
      RECT 99.105 -36.335 99.245 -36.165 ;
      RECT 99.155 -35.13 99.245 -34.122 ;
      RECT 99.105 -34.895 99.245 -34.725 ;
      RECT 99.155 -33.708 99.245 -32.7 ;
      RECT 99.105 -33.105 99.245 -32.935 ;
      RECT 99.155 -31.9 99.245 -30.892 ;
      RECT 99.105 -31.665 99.245 -31.495 ;
      RECT 99.155 -30.478 99.245 -29.47 ;
      RECT 99.105 -29.875 99.245 -29.705 ;
      RECT 99.155 -28.67 99.245 -27.662 ;
      RECT 99.105 -28.435 99.245 -28.265 ;
      RECT 99.155 -27.248 99.245 -26.24 ;
      RECT 99.105 -26.645 99.245 -26.475 ;
      RECT 99.155 -25.44 99.245 -24.432 ;
      RECT 99.105 -25.205 99.245 -25.035 ;
      RECT 99.155 -24.018 99.245 -23.01 ;
      RECT 99.105 -23.415 99.245 -23.245 ;
      RECT 99.155 -22.21 99.245 -21.202 ;
      RECT 99.105 -21.975 99.245 -21.805 ;
      RECT 99.155 -20.788 99.245 -19.78 ;
      RECT 99.105 -20.185 99.245 -20.015 ;
      RECT 99.155 -18.98 99.245 -17.972 ;
      RECT 99.105 -18.745 99.245 -18.575 ;
      RECT 99.155 -17.558 99.245 -16.55 ;
      RECT 99.105 -16.955 99.245 -16.785 ;
      RECT 99.155 -15.75 99.245 -14.742 ;
      RECT 99.105 -15.515 99.245 -15.345 ;
      RECT 99.155 -14.328 99.245 -13.32 ;
      RECT 99.105 -13.725 99.245 -13.555 ;
      RECT 99.155 -12.52 99.245 -11.512 ;
      RECT 99.105 -12.285 99.245 -12.115 ;
      RECT 99.155 -11.098 99.245 -10.09 ;
      RECT 99.105 -10.495 99.245 -10.325 ;
      RECT 99.155 -9.29 99.245 -8.282 ;
      RECT 99.105 -9.055 99.245 -8.885 ;
      RECT 99.155 -7.868 99.245 -6.86 ;
      RECT 99.105 -7.265 99.245 -7.095 ;
      RECT 99.155 -6.06 99.245 -5.052 ;
      RECT 99.105 -5.825 99.245 -5.655 ;
      RECT 99.155 -4.638 99.245 -3.63 ;
      RECT 99.105 -4.035 99.245 -3.865 ;
      RECT 99.155 -2.83 99.245 -1.822 ;
      RECT 99.105 -2.595 99.245 -2.425 ;
      RECT 99.155 -1.408 99.245 -0.4 ;
      RECT 99.105 -0.805 99.245 -0.635 ;
      RECT 99.155 0.4 99.245 1.408 ;
      RECT 99.105 0.635 99.245 0.805 ;
      RECT 98.755 -101.538 98.845 -100.531 ;
      RECT 98.755 -101.225 98.895 -101.055 ;
      RECT 98.755 -99.729 98.845 -98.722 ;
      RECT 98.755 -99.205 98.895 -99.035 ;
      RECT 98.755 -98.308 98.845 -97.301 ;
      RECT 98.755 -97.995 98.895 -97.825 ;
      RECT 98.755 -96.499 98.845 -95.492 ;
      RECT 98.755 -95.975 98.895 -95.805 ;
      RECT 98.755 -95.078 98.845 -94.071 ;
      RECT 98.755 -94.765 98.895 -94.595 ;
      RECT 98.755 -93.269 98.845 -92.262 ;
      RECT 98.755 -92.745 98.895 -92.575 ;
      RECT 98.755 -91.848 98.845 -90.841 ;
      RECT 98.755 -91.535 98.895 -91.365 ;
      RECT 98.755 -90.039 98.845 -89.032 ;
      RECT 98.755 -89.515 98.895 -89.345 ;
      RECT 98.755 -88.618 98.845 -87.611 ;
      RECT 98.755 -88.305 98.895 -88.135 ;
      RECT 98.755 -86.809 98.845 -85.802 ;
      RECT 98.755 -86.285 98.895 -86.115 ;
      RECT 98.755 -85.388 98.845 -84.381 ;
      RECT 98.755 -85.075 98.895 -84.905 ;
      RECT 98.755 -83.579 98.845 -82.572 ;
      RECT 98.755 -83.055 98.895 -82.885 ;
      RECT 98.755 -82.158 98.845 -81.151 ;
      RECT 98.755 -81.845 98.895 -81.675 ;
      RECT 98.755 -80.349 98.845 -79.342 ;
      RECT 98.755 -79.825 98.895 -79.655 ;
      RECT 98.755 -78.928 98.845 -77.921 ;
      RECT 98.755 -78.615 98.895 -78.445 ;
      RECT 98.755 -77.119 98.845 -76.112 ;
      RECT 98.755 -76.595 98.895 -76.425 ;
      RECT 98.755 -75.698 98.845 -74.691 ;
      RECT 98.755 -75.385 98.895 -75.215 ;
      RECT 98.755 -73.889 98.845 -72.882 ;
      RECT 98.755 -73.365 98.895 -73.195 ;
      RECT 98.755 -72.468 98.845 -71.461 ;
      RECT 98.755 -72.155 98.895 -71.985 ;
      RECT 98.755 -70.659 98.845 -69.652 ;
      RECT 98.755 -70.135 98.895 -69.965 ;
      RECT 98.755 -69.238 98.845 -68.231 ;
      RECT 98.755 -68.925 98.895 -68.755 ;
      RECT 98.755 -67.429 98.845 -66.422 ;
      RECT 98.755 -66.905 98.895 -66.735 ;
      RECT 98.755 -66.008 98.845 -65.001 ;
      RECT 98.755 -65.695 98.895 -65.525 ;
      RECT 98.755 -64.199 98.845 -63.192 ;
      RECT 98.755 -63.675 98.895 -63.505 ;
      RECT 98.755 -62.778 98.845 -61.771 ;
      RECT 98.755 -62.465 98.895 -62.295 ;
      RECT 98.755 -60.969 98.845 -59.962 ;
      RECT 98.755 -60.445 98.895 -60.275 ;
      RECT 98.755 -59.548 98.845 -58.541 ;
      RECT 98.755 -59.235 98.895 -59.065 ;
      RECT 98.755 -57.739 98.845 -56.732 ;
      RECT 98.755 -57.215 98.895 -57.045 ;
      RECT 98.755 -56.318 98.845 -55.311 ;
      RECT 98.755 -56.005 98.895 -55.835 ;
      RECT 98.755 -54.509 98.845 -53.502 ;
      RECT 98.755 -53.985 98.895 -53.815 ;
      RECT 98.755 -53.088 98.845 -52.081 ;
      RECT 98.755 -52.775 98.895 -52.605 ;
      RECT 98.755 -51.279 98.845 -50.272 ;
      RECT 98.755 -50.755 98.895 -50.585 ;
      RECT 98.755 -49.858 98.845 -48.851 ;
      RECT 98.755 -49.545 98.895 -49.375 ;
      RECT 98.755 -48.049 98.845 -47.042 ;
      RECT 98.755 -47.525 98.895 -47.355 ;
      RECT 98.755 -46.628 98.845 -45.621 ;
      RECT 98.755 -46.315 98.895 -46.145 ;
      RECT 98.755 -44.819 98.845 -43.812 ;
      RECT 98.755 -44.295 98.895 -44.125 ;
      RECT 98.755 -43.398 98.845 -42.391 ;
      RECT 98.755 -43.085 98.895 -42.915 ;
      RECT 98.755 -41.589 98.845 -40.582 ;
      RECT 98.755 -41.065 98.895 -40.895 ;
      RECT 98.755 -40.168 98.845 -39.161 ;
      RECT 98.755 -39.855 98.895 -39.685 ;
      RECT 98.755 -38.359 98.845 -37.352 ;
      RECT 98.755 -37.835 98.895 -37.665 ;
      RECT 98.755 -36.938 98.845 -35.931 ;
      RECT 98.755 -36.625 98.895 -36.455 ;
      RECT 98.755 -35.129 98.845 -34.122 ;
      RECT 98.755 -34.605 98.895 -34.435 ;
      RECT 98.755 -33.708 98.845 -32.701 ;
      RECT 98.755 -33.395 98.895 -33.225 ;
      RECT 98.755 -31.899 98.845 -30.892 ;
      RECT 98.755 -31.375 98.895 -31.205 ;
      RECT 98.755 -30.478 98.845 -29.471 ;
      RECT 98.755 -30.165 98.895 -29.995 ;
      RECT 98.755 -28.669 98.845 -27.662 ;
      RECT 98.755 -28.145 98.895 -27.975 ;
      RECT 98.755 -27.248 98.845 -26.241 ;
      RECT 98.755 -26.935 98.895 -26.765 ;
      RECT 98.755 -25.439 98.845 -24.432 ;
      RECT 98.755 -24.915 98.895 -24.745 ;
      RECT 98.755 -24.018 98.845 -23.011 ;
      RECT 98.755 -23.705 98.895 -23.535 ;
      RECT 98.755 -22.209 98.845 -21.202 ;
      RECT 98.755 -21.685 98.895 -21.515 ;
      RECT 98.755 -20.788 98.845 -19.781 ;
      RECT 98.755 -20.475 98.895 -20.305 ;
      RECT 98.755 -18.979 98.845 -17.972 ;
      RECT 98.755 -18.455 98.895 -18.285 ;
      RECT 98.755 -17.558 98.845 -16.551 ;
      RECT 98.755 -17.245 98.895 -17.075 ;
      RECT 98.755 -15.749 98.845 -14.742 ;
      RECT 98.755 -15.225 98.895 -15.055 ;
      RECT 98.755 -14.328 98.845 -13.321 ;
      RECT 98.755 -14.015 98.895 -13.845 ;
      RECT 98.755 -12.519 98.845 -11.512 ;
      RECT 98.755 -11.995 98.895 -11.825 ;
      RECT 98.755 -11.098 98.845 -10.091 ;
      RECT 98.755 -10.785 98.895 -10.615 ;
      RECT 98.755 -9.289 98.845 -8.282 ;
      RECT 98.755 -8.765 98.895 -8.595 ;
      RECT 98.755 -7.868 98.845 -6.861 ;
      RECT 98.755 -7.555 98.895 -7.385 ;
      RECT 98.755 -6.059 98.845 -5.052 ;
      RECT 98.755 -5.535 98.895 -5.365 ;
      RECT 98.755 -4.638 98.845 -3.631 ;
      RECT 98.755 -4.325 98.895 -4.155 ;
      RECT 98.755 -2.829 98.845 -1.822 ;
      RECT 98.755 -2.305 98.895 -2.135 ;
      RECT 98.755 -1.408 98.845 -0.401 ;
      RECT 98.755 -1.095 98.895 -0.925 ;
      RECT 98.755 0.401 98.845 1.408 ;
      RECT 98.755 0.925 98.895 1.095 ;
      RECT 96.905 -111.685 98.385 -111.585 ;
      RECT 96.905 -112.055 97.005 -111.585 ;
      RECT 96.71 -114.395 98.285 -114.275 ;
      RECT 98.185 -114.895 98.285 -114.275 ;
      RECT 97.59 -114.895 97.69 -114.275 ;
      RECT 96.71 -114.85 96.81 -114.275 ;
      RECT 97.955 -101.538 98.045 -100.53 ;
      RECT 97.905 -100.935 98.045 -100.765 ;
      RECT 97.955 -99.73 98.045 -98.722 ;
      RECT 97.905 -99.495 98.045 -99.325 ;
      RECT 97.955 -98.308 98.045 -97.3 ;
      RECT 97.905 -97.705 98.045 -97.535 ;
      RECT 97.955 -96.5 98.045 -95.492 ;
      RECT 97.905 -96.265 98.045 -96.095 ;
      RECT 97.955 -95.078 98.045 -94.07 ;
      RECT 97.905 -94.475 98.045 -94.305 ;
      RECT 97.955 -93.27 98.045 -92.262 ;
      RECT 97.905 -93.035 98.045 -92.865 ;
      RECT 97.955 -91.848 98.045 -90.84 ;
      RECT 97.905 -91.245 98.045 -91.075 ;
      RECT 97.955 -90.04 98.045 -89.032 ;
      RECT 97.905 -89.805 98.045 -89.635 ;
      RECT 97.955 -88.618 98.045 -87.61 ;
      RECT 97.905 -88.015 98.045 -87.845 ;
      RECT 97.955 -86.81 98.045 -85.802 ;
      RECT 97.905 -86.575 98.045 -86.405 ;
      RECT 97.955 -85.388 98.045 -84.38 ;
      RECT 97.905 -84.785 98.045 -84.615 ;
      RECT 97.955 -83.58 98.045 -82.572 ;
      RECT 97.905 -83.345 98.045 -83.175 ;
      RECT 97.955 -82.158 98.045 -81.15 ;
      RECT 97.905 -81.555 98.045 -81.385 ;
      RECT 97.955 -80.35 98.045 -79.342 ;
      RECT 97.905 -80.115 98.045 -79.945 ;
      RECT 97.955 -78.928 98.045 -77.92 ;
      RECT 97.905 -78.325 98.045 -78.155 ;
      RECT 97.955 -77.12 98.045 -76.112 ;
      RECT 97.905 -76.885 98.045 -76.715 ;
      RECT 97.955 -75.698 98.045 -74.69 ;
      RECT 97.905 -75.095 98.045 -74.925 ;
      RECT 97.955 -73.89 98.045 -72.882 ;
      RECT 97.905 -73.655 98.045 -73.485 ;
      RECT 97.955 -72.468 98.045 -71.46 ;
      RECT 97.905 -71.865 98.045 -71.695 ;
      RECT 97.955 -70.66 98.045 -69.652 ;
      RECT 97.905 -70.425 98.045 -70.255 ;
      RECT 97.955 -69.238 98.045 -68.23 ;
      RECT 97.905 -68.635 98.045 -68.465 ;
      RECT 97.955 -67.43 98.045 -66.422 ;
      RECT 97.905 -67.195 98.045 -67.025 ;
      RECT 97.955 -66.008 98.045 -65 ;
      RECT 97.905 -65.405 98.045 -65.235 ;
      RECT 97.955 -64.2 98.045 -63.192 ;
      RECT 97.905 -63.965 98.045 -63.795 ;
      RECT 97.955 -62.778 98.045 -61.77 ;
      RECT 97.905 -62.175 98.045 -62.005 ;
      RECT 97.955 -60.97 98.045 -59.962 ;
      RECT 97.905 -60.735 98.045 -60.565 ;
      RECT 97.955 -59.548 98.045 -58.54 ;
      RECT 97.905 -58.945 98.045 -58.775 ;
      RECT 97.955 -57.74 98.045 -56.732 ;
      RECT 97.905 -57.505 98.045 -57.335 ;
      RECT 97.955 -56.318 98.045 -55.31 ;
      RECT 97.905 -55.715 98.045 -55.545 ;
      RECT 97.955 -54.51 98.045 -53.502 ;
      RECT 97.905 -54.275 98.045 -54.105 ;
      RECT 97.955 -53.088 98.045 -52.08 ;
      RECT 97.905 -52.485 98.045 -52.315 ;
      RECT 97.955 -51.28 98.045 -50.272 ;
      RECT 97.905 -51.045 98.045 -50.875 ;
      RECT 97.955 -49.858 98.045 -48.85 ;
      RECT 97.905 -49.255 98.045 -49.085 ;
      RECT 97.955 -48.05 98.045 -47.042 ;
      RECT 97.905 -47.815 98.045 -47.645 ;
      RECT 97.955 -46.628 98.045 -45.62 ;
      RECT 97.905 -46.025 98.045 -45.855 ;
      RECT 97.955 -44.82 98.045 -43.812 ;
      RECT 97.905 -44.585 98.045 -44.415 ;
      RECT 97.955 -43.398 98.045 -42.39 ;
      RECT 97.905 -42.795 98.045 -42.625 ;
      RECT 97.955 -41.59 98.045 -40.582 ;
      RECT 97.905 -41.355 98.045 -41.185 ;
      RECT 97.955 -40.168 98.045 -39.16 ;
      RECT 97.905 -39.565 98.045 -39.395 ;
      RECT 97.955 -38.36 98.045 -37.352 ;
      RECT 97.905 -38.125 98.045 -37.955 ;
      RECT 97.955 -36.938 98.045 -35.93 ;
      RECT 97.905 -36.335 98.045 -36.165 ;
      RECT 97.955 -35.13 98.045 -34.122 ;
      RECT 97.905 -34.895 98.045 -34.725 ;
      RECT 97.955 -33.708 98.045 -32.7 ;
      RECT 97.905 -33.105 98.045 -32.935 ;
      RECT 97.955 -31.9 98.045 -30.892 ;
      RECT 97.905 -31.665 98.045 -31.495 ;
      RECT 97.955 -30.478 98.045 -29.47 ;
      RECT 97.905 -29.875 98.045 -29.705 ;
      RECT 97.955 -28.67 98.045 -27.662 ;
      RECT 97.905 -28.435 98.045 -28.265 ;
      RECT 97.955 -27.248 98.045 -26.24 ;
      RECT 97.905 -26.645 98.045 -26.475 ;
      RECT 97.955 -25.44 98.045 -24.432 ;
      RECT 97.905 -25.205 98.045 -25.035 ;
      RECT 97.955 -24.018 98.045 -23.01 ;
      RECT 97.905 -23.415 98.045 -23.245 ;
      RECT 97.955 -22.21 98.045 -21.202 ;
      RECT 97.905 -21.975 98.045 -21.805 ;
      RECT 97.955 -20.788 98.045 -19.78 ;
      RECT 97.905 -20.185 98.045 -20.015 ;
      RECT 97.955 -18.98 98.045 -17.972 ;
      RECT 97.905 -18.745 98.045 -18.575 ;
      RECT 97.955 -17.558 98.045 -16.55 ;
      RECT 97.905 -16.955 98.045 -16.785 ;
      RECT 97.955 -15.75 98.045 -14.742 ;
      RECT 97.905 -15.515 98.045 -15.345 ;
      RECT 97.955 -14.328 98.045 -13.32 ;
      RECT 97.905 -13.725 98.045 -13.555 ;
      RECT 97.955 -12.52 98.045 -11.512 ;
      RECT 97.905 -12.285 98.045 -12.115 ;
      RECT 97.955 -11.098 98.045 -10.09 ;
      RECT 97.905 -10.495 98.045 -10.325 ;
      RECT 97.955 -9.29 98.045 -8.282 ;
      RECT 97.905 -9.055 98.045 -8.885 ;
      RECT 97.955 -7.868 98.045 -6.86 ;
      RECT 97.905 -7.265 98.045 -7.095 ;
      RECT 97.955 -6.06 98.045 -5.052 ;
      RECT 97.905 -5.825 98.045 -5.655 ;
      RECT 97.955 -4.638 98.045 -3.63 ;
      RECT 97.905 -4.035 98.045 -3.865 ;
      RECT 97.955 -2.83 98.045 -1.822 ;
      RECT 97.905 -2.595 98.045 -2.425 ;
      RECT 97.955 -1.408 98.045 -0.4 ;
      RECT 97.905 -0.805 98.045 -0.635 ;
      RECT 97.955 0.4 98.045 1.408 ;
      RECT 97.905 0.635 98.045 0.805 ;
      RECT 97.83 -114.685 98.005 -114.515 ;
      RECT 97.905 -114.895 98.005 -114.515 ;
      RECT 96.945 -113.555 97.045 -113.09 ;
      RECT 97.31 -113.555 97.41 -113.1 ;
      RECT 96.945 -113.555 97.79 -113.385 ;
      RECT 97.555 -101.538 97.645 -100.531 ;
      RECT 97.555 -101.225 97.695 -101.055 ;
      RECT 97.555 -99.729 97.645 -98.722 ;
      RECT 97.555 -99.205 97.695 -99.035 ;
      RECT 97.555 -98.308 97.645 -97.301 ;
      RECT 97.555 -97.995 97.695 -97.825 ;
      RECT 97.555 -96.499 97.645 -95.492 ;
      RECT 97.555 -95.975 97.695 -95.805 ;
      RECT 97.555 -95.078 97.645 -94.071 ;
      RECT 97.555 -94.765 97.695 -94.595 ;
      RECT 97.555 -93.269 97.645 -92.262 ;
      RECT 97.555 -92.745 97.695 -92.575 ;
      RECT 97.555 -91.848 97.645 -90.841 ;
      RECT 97.555 -91.535 97.695 -91.365 ;
      RECT 97.555 -90.039 97.645 -89.032 ;
      RECT 97.555 -89.515 97.695 -89.345 ;
      RECT 97.555 -88.618 97.645 -87.611 ;
      RECT 97.555 -88.305 97.695 -88.135 ;
      RECT 97.555 -86.809 97.645 -85.802 ;
      RECT 97.555 -86.285 97.695 -86.115 ;
      RECT 97.555 -85.388 97.645 -84.381 ;
      RECT 97.555 -85.075 97.695 -84.905 ;
      RECT 97.555 -83.579 97.645 -82.572 ;
      RECT 97.555 -83.055 97.695 -82.885 ;
      RECT 97.555 -82.158 97.645 -81.151 ;
      RECT 97.555 -81.845 97.695 -81.675 ;
      RECT 97.555 -80.349 97.645 -79.342 ;
      RECT 97.555 -79.825 97.695 -79.655 ;
      RECT 97.555 -78.928 97.645 -77.921 ;
      RECT 97.555 -78.615 97.695 -78.445 ;
      RECT 97.555 -77.119 97.645 -76.112 ;
      RECT 97.555 -76.595 97.695 -76.425 ;
      RECT 97.555 -75.698 97.645 -74.691 ;
      RECT 97.555 -75.385 97.695 -75.215 ;
      RECT 97.555 -73.889 97.645 -72.882 ;
      RECT 97.555 -73.365 97.695 -73.195 ;
      RECT 97.555 -72.468 97.645 -71.461 ;
      RECT 97.555 -72.155 97.695 -71.985 ;
      RECT 97.555 -70.659 97.645 -69.652 ;
      RECT 97.555 -70.135 97.695 -69.965 ;
      RECT 97.555 -69.238 97.645 -68.231 ;
      RECT 97.555 -68.925 97.695 -68.755 ;
      RECT 97.555 -67.429 97.645 -66.422 ;
      RECT 97.555 -66.905 97.695 -66.735 ;
      RECT 97.555 -66.008 97.645 -65.001 ;
      RECT 97.555 -65.695 97.695 -65.525 ;
      RECT 97.555 -64.199 97.645 -63.192 ;
      RECT 97.555 -63.675 97.695 -63.505 ;
      RECT 97.555 -62.778 97.645 -61.771 ;
      RECT 97.555 -62.465 97.695 -62.295 ;
      RECT 97.555 -60.969 97.645 -59.962 ;
      RECT 97.555 -60.445 97.695 -60.275 ;
      RECT 97.555 -59.548 97.645 -58.541 ;
      RECT 97.555 -59.235 97.695 -59.065 ;
      RECT 97.555 -57.739 97.645 -56.732 ;
      RECT 97.555 -57.215 97.695 -57.045 ;
      RECT 97.555 -56.318 97.645 -55.311 ;
      RECT 97.555 -56.005 97.695 -55.835 ;
      RECT 97.555 -54.509 97.645 -53.502 ;
      RECT 97.555 -53.985 97.695 -53.815 ;
      RECT 97.555 -53.088 97.645 -52.081 ;
      RECT 97.555 -52.775 97.695 -52.605 ;
      RECT 97.555 -51.279 97.645 -50.272 ;
      RECT 97.555 -50.755 97.695 -50.585 ;
      RECT 97.555 -49.858 97.645 -48.851 ;
      RECT 97.555 -49.545 97.695 -49.375 ;
      RECT 97.555 -48.049 97.645 -47.042 ;
      RECT 97.555 -47.525 97.695 -47.355 ;
      RECT 97.555 -46.628 97.645 -45.621 ;
      RECT 97.555 -46.315 97.695 -46.145 ;
      RECT 97.555 -44.819 97.645 -43.812 ;
      RECT 97.555 -44.295 97.695 -44.125 ;
      RECT 97.555 -43.398 97.645 -42.391 ;
      RECT 97.555 -43.085 97.695 -42.915 ;
      RECT 97.555 -41.589 97.645 -40.582 ;
      RECT 97.555 -41.065 97.695 -40.895 ;
      RECT 97.555 -40.168 97.645 -39.161 ;
      RECT 97.555 -39.855 97.695 -39.685 ;
      RECT 97.555 -38.359 97.645 -37.352 ;
      RECT 97.555 -37.835 97.695 -37.665 ;
      RECT 97.555 -36.938 97.645 -35.931 ;
      RECT 97.555 -36.625 97.695 -36.455 ;
      RECT 97.555 -35.129 97.645 -34.122 ;
      RECT 97.555 -34.605 97.695 -34.435 ;
      RECT 97.555 -33.708 97.645 -32.701 ;
      RECT 97.555 -33.395 97.695 -33.225 ;
      RECT 97.555 -31.899 97.645 -30.892 ;
      RECT 97.555 -31.375 97.695 -31.205 ;
      RECT 97.555 -30.478 97.645 -29.471 ;
      RECT 97.555 -30.165 97.695 -29.995 ;
      RECT 97.555 -28.669 97.645 -27.662 ;
      RECT 97.555 -28.145 97.695 -27.975 ;
      RECT 97.555 -27.248 97.645 -26.241 ;
      RECT 97.555 -26.935 97.695 -26.765 ;
      RECT 97.555 -25.439 97.645 -24.432 ;
      RECT 97.555 -24.915 97.695 -24.745 ;
      RECT 97.555 -24.018 97.645 -23.011 ;
      RECT 97.555 -23.705 97.695 -23.535 ;
      RECT 97.555 -22.209 97.645 -21.202 ;
      RECT 97.555 -21.685 97.695 -21.515 ;
      RECT 97.555 -20.788 97.645 -19.781 ;
      RECT 97.555 -20.475 97.695 -20.305 ;
      RECT 97.555 -18.979 97.645 -17.972 ;
      RECT 97.555 -18.455 97.695 -18.285 ;
      RECT 97.555 -17.558 97.645 -16.551 ;
      RECT 97.555 -17.245 97.695 -17.075 ;
      RECT 97.555 -15.749 97.645 -14.742 ;
      RECT 97.555 -15.225 97.695 -15.055 ;
      RECT 97.555 -14.328 97.645 -13.321 ;
      RECT 97.555 -14.015 97.695 -13.845 ;
      RECT 97.555 -12.519 97.645 -11.512 ;
      RECT 97.555 -11.995 97.695 -11.825 ;
      RECT 97.555 -11.098 97.645 -10.091 ;
      RECT 97.555 -10.785 97.695 -10.615 ;
      RECT 97.555 -9.289 97.645 -8.282 ;
      RECT 97.555 -8.765 97.695 -8.595 ;
      RECT 97.555 -7.868 97.645 -6.861 ;
      RECT 97.555 -7.555 97.695 -7.385 ;
      RECT 97.555 -6.059 97.645 -5.052 ;
      RECT 97.555 -5.535 97.695 -5.365 ;
      RECT 97.555 -4.638 97.645 -3.631 ;
      RECT 97.555 -4.325 97.695 -4.155 ;
      RECT 97.555 -2.829 97.645 -1.822 ;
      RECT 97.555 -2.305 97.695 -2.135 ;
      RECT 97.555 -1.408 97.645 -0.401 ;
      RECT 97.555 -1.095 97.695 -0.925 ;
      RECT 97.555 0.401 97.645 1.408 ;
      RECT 97.555 0.925 97.695 1.095 ;
      RECT 97.24 -114.685 97.41 -114.515 ;
      RECT 97.31 -114.895 97.41 -114.515 ;
      RECT 96.755 -101.538 96.845 -100.53 ;
      RECT 96.705 -100.935 96.845 -100.765 ;
      RECT 96.755 -99.73 96.845 -98.722 ;
      RECT 96.705 -99.495 96.845 -99.325 ;
      RECT 96.755 -98.308 96.845 -97.3 ;
      RECT 96.705 -97.705 96.845 -97.535 ;
      RECT 96.755 -96.5 96.845 -95.492 ;
      RECT 96.705 -96.265 96.845 -96.095 ;
      RECT 96.755 -95.078 96.845 -94.07 ;
      RECT 96.705 -94.475 96.845 -94.305 ;
      RECT 96.755 -93.27 96.845 -92.262 ;
      RECT 96.705 -93.035 96.845 -92.865 ;
      RECT 96.755 -91.848 96.845 -90.84 ;
      RECT 96.705 -91.245 96.845 -91.075 ;
      RECT 96.755 -90.04 96.845 -89.032 ;
      RECT 96.705 -89.805 96.845 -89.635 ;
      RECT 96.755 -88.618 96.845 -87.61 ;
      RECT 96.705 -88.015 96.845 -87.845 ;
      RECT 96.755 -86.81 96.845 -85.802 ;
      RECT 96.705 -86.575 96.845 -86.405 ;
      RECT 96.755 -85.388 96.845 -84.38 ;
      RECT 96.705 -84.785 96.845 -84.615 ;
      RECT 96.755 -83.58 96.845 -82.572 ;
      RECT 96.705 -83.345 96.845 -83.175 ;
      RECT 96.755 -82.158 96.845 -81.15 ;
      RECT 96.705 -81.555 96.845 -81.385 ;
      RECT 96.755 -80.35 96.845 -79.342 ;
      RECT 96.705 -80.115 96.845 -79.945 ;
      RECT 96.755 -78.928 96.845 -77.92 ;
      RECT 96.705 -78.325 96.845 -78.155 ;
      RECT 96.755 -77.12 96.845 -76.112 ;
      RECT 96.705 -76.885 96.845 -76.715 ;
      RECT 96.755 -75.698 96.845 -74.69 ;
      RECT 96.705 -75.095 96.845 -74.925 ;
      RECT 96.755 -73.89 96.845 -72.882 ;
      RECT 96.705 -73.655 96.845 -73.485 ;
      RECT 96.755 -72.468 96.845 -71.46 ;
      RECT 96.705 -71.865 96.845 -71.695 ;
      RECT 96.755 -70.66 96.845 -69.652 ;
      RECT 96.705 -70.425 96.845 -70.255 ;
      RECT 96.755 -69.238 96.845 -68.23 ;
      RECT 96.705 -68.635 96.845 -68.465 ;
      RECT 96.755 -67.43 96.845 -66.422 ;
      RECT 96.705 -67.195 96.845 -67.025 ;
      RECT 96.755 -66.008 96.845 -65 ;
      RECT 96.705 -65.405 96.845 -65.235 ;
      RECT 96.755 -64.2 96.845 -63.192 ;
      RECT 96.705 -63.965 96.845 -63.795 ;
      RECT 96.755 -62.778 96.845 -61.77 ;
      RECT 96.705 -62.175 96.845 -62.005 ;
      RECT 96.755 -60.97 96.845 -59.962 ;
      RECT 96.705 -60.735 96.845 -60.565 ;
      RECT 96.755 -59.548 96.845 -58.54 ;
      RECT 96.705 -58.945 96.845 -58.775 ;
      RECT 96.755 -57.74 96.845 -56.732 ;
      RECT 96.705 -57.505 96.845 -57.335 ;
      RECT 96.755 -56.318 96.845 -55.31 ;
      RECT 96.705 -55.715 96.845 -55.545 ;
      RECT 96.755 -54.51 96.845 -53.502 ;
      RECT 96.705 -54.275 96.845 -54.105 ;
      RECT 96.755 -53.088 96.845 -52.08 ;
      RECT 96.705 -52.485 96.845 -52.315 ;
      RECT 96.755 -51.28 96.845 -50.272 ;
      RECT 96.705 -51.045 96.845 -50.875 ;
      RECT 96.755 -49.858 96.845 -48.85 ;
      RECT 96.705 -49.255 96.845 -49.085 ;
      RECT 96.755 -48.05 96.845 -47.042 ;
      RECT 96.705 -47.815 96.845 -47.645 ;
      RECT 96.755 -46.628 96.845 -45.62 ;
      RECT 96.705 -46.025 96.845 -45.855 ;
      RECT 96.755 -44.82 96.845 -43.812 ;
      RECT 96.705 -44.585 96.845 -44.415 ;
      RECT 96.755 -43.398 96.845 -42.39 ;
      RECT 96.705 -42.795 96.845 -42.625 ;
      RECT 96.755 -41.59 96.845 -40.582 ;
      RECT 96.705 -41.355 96.845 -41.185 ;
      RECT 96.755 -40.168 96.845 -39.16 ;
      RECT 96.705 -39.565 96.845 -39.395 ;
      RECT 96.755 -38.36 96.845 -37.352 ;
      RECT 96.705 -38.125 96.845 -37.955 ;
      RECT 96.755 -36.938 96.845 -35.93 ;
      RECT 96.705 -36.335 96.845 -36.165 ;
      RECT 96.755 -35.13 96.845 -34.122 ;
      RECT 96.705 -34.895 96.845 -34.725 ;
      RECT 96.755 -33.708 96.845 -32.7 ;
      RECT 96.705 -33.105 96.845 -32.935 ;
      RECT 96.755 -31.9 96.845 -30.892 ;
      RECT 96.705 -31.665 96.845 -31.495 ;
      RECT 96.755 -30.478 96.845 -29.47 ;
      RECT 96.705 -29.875 96.845 -29.705 ;
      RECT 96.755 -28.67 96.845 -27.662 ;
      RECT 96.705 -28.435 96.845 -28.265 ;
      RECT 96.755 -27.248 96.845 -26.24 ;
      RECT 96.705 -26.645 96.845 -26.475 ;
      RECT 96.755 -25.44 96.845 -24.432 ;
      RECT 96.705 -25.205 96.845 -25.035 ;
      RECT 96.755 -24.018 96.845 -23.01 ;
      RECT 96.705 -23.415 96.845 -23.245 ;
      RECT 96.755 -22.21 96.845 -21.202 ;
      RECT 96.705 -21.975 96.845 -21.805 ;
      RECT 96.755 -20.788 96.845 -19.78 ;
      RECT 96.705 -20.185 96.845 -20.015 ;
      RECT 96.755 -18.98 96.845 -17.972 ;
      RECT 96.705 -18.745 96.845 -18.575 ;
      RECT 96.755 -17.558 96.845 -16.55 ;
      RECT 96.705 -16.955 96.845 -16.785 ;
      RECT 96.755 -15.75 96.845 -14.742 ;
      RECT 96.705 -15.515 96.845 -15.345 ;
      RECT 96.755 -14.328 96.845 -13.32 ;
      RECT 96.705 -13.725 96.845 -13.555 ;
      RECT 96.755 -12.52 96.845 -11.512 ;
      RECT 96.705 -12.285 96.845 -12.115 ;
      RECT 96.755 -11.098 96.845 -10.09 ;
      RECT 96.705 -10.495 96.845 -10.325 ;
      RECT 96.755 -9.29 96.845 -8.282 ;
      RECT 96.705 -9.055 96.845 -8.885 ;
      RECT 96.755 -7.868 96.845 -6.86 ;
      RECT 96.705 -7.265 96.845 -7.095 ;
      RECT 96.755 -6.06 96.845 -5.052 ;
      RECT 96.705 -5.825 96.845 -5.655 ;
      RECT 96.755 -4.638 96.845 -3.63 ;
      RECT 96.705 -4.035 96.845 -3.865 ;
      RECT 96.755 -2.83 96.845 -1.822 ;
      RECT 96.705 -2.595 96.845 -2.425 ;
      RECT 96.755 -1.408 96.845 -0.4 ;
      RECT 96.705 -0.805 96.845 -0.635 ;
      RECT 96.755 0.4 96.845 1.408 ;
      RECT 96.705 0.635 96.845 0.805 ;
      RECT 96.355 -101.538 96.445 -100.531 ;
      RECT 96.355 -101.225 96.495 -101.055 ;
      RECT 96.355 -99.729 96.445 -98.722 ;
      RECT 96.355 -99.205 96.495 -99.035 ;
      RECT 96.355 -98.308 96.445 -97.301 ;
      RECT 96.355 -97.995 96.495 -97.825 ;
      RECT 96.355 -96.499 96.445 -95.492 ;
      RECT 96.355 -95.975 96.495 -95.805 ;
      RECT 96.355 -95.078 96.445 -94.071 ;
      RECT 96.355 -94.765 96.495 -94.595 ;
      RECT 96.355 -93.269 96.445 -92.262 ;
      RECT 96.355 -92.745 96.495 -92.575 ;
      RECT 96.355 -91.848 96.445 -90.841 ;
      RECT 96.355 -91.535 96.495 -91.365 ;
      RECT 96.355 -90.039 96.445 -89.032 ;
      RECT 96.355 -89.515 96.495 -89.345 ;
      RECT 96.355 -88.618 96.445 -87.611 ;
      RECT 96.355 -88.305 96.495 -88.135 ;
      RECT 96.355 -86.809 96.445 -85.802 ;
      RECT 96.355 -86.285 96.495 -86.115 ;
      RECT 96.355 -85.388 96.445 -84.381 ;
      RECT 96.355 -85.075 96.495 -84.905 ;
      RECT 96.355 -83.579 96.445 -82.572 ;
      RECT 96.355 -83.055 96.495 -82.885 ;
      RECT 96.355 -82.158 96.445 -81.151 ;
      RECT 96.355 -81.845 96.495 -81.675 ;
      RECT 96.355 -80.349 96.445 -79.342 ;
      RECT 96.355 -79.825 96.495 -79.655 ;
      RECT 96.355 -78.928 96.445 -77.921 ;
      RECT 96.355 -78.615 96.495 -78.445 ;
      RECT 96.355 -77.119 96.445 -76.112 ;
      RECT 96.355 -76.595 96.495 -76.425 ;
      RECT 96.355 -75.698 96.445 -74.691 ;
      RECT 96.355 -75.385 96.495 -75.215 ;
      RECT 96.355 -73.889 96.445 -72.882 ;
      RECT 96.355 -73.365 96.495 -73.195 ;
      RECT 96.355 -72.468 96.445 -71.461 ;
      RECT 96.355 -72.155 96.495 -71.985 ;
      RECT 96.355 -70.659 96.445 -69.652 ;
      RECT 96.355 -70.135 96.495 -69.965 ;
      RECT 96.355 -69.238 96.445 -68.231 ;
      RECT 96.355 -68.925 96.495 -68.755 ;
      RECT 96.355 -67.429 96.445 -66.422 ;
      RECT 96.355 -66.905 96.495 -66.735 ;
      RECT 96.355 -66.008 96.445 -65.001 ;
      RECT 96.355 -65.695 96.495 -65.525 ;
      RECT 96.355 -64.199 96.445 -63.192 ;
      RECT 96.355 -63.675 96.495 -63.505 ;
      RECT 96.355 -62.778 96.445 -61.771 ;
      RECT 96.355 -62.465 96.495 -62.295 ;
      RECT 96.355 -60.969 96.445 -59.962 ;
      RECT 96.355 -60.445 96.495 -60.275 ;
      RECT 96.355 -59.548 96.445 -58.541 ;
      RECT 96.355 -59.235 96.495 -59.065 ;
      RECT 96.355 -57.739 96.445 -56.732 ;
      RECT 96.355 -57.215 96.495 -57.045 ;
      RECT 96.355 -56.318 96.445 -55.311 ;
      RECT 96.355 -56.005 96.495 -55.835 ;
      RECT 96.355 -54.509 96.445 -53.502 ;
      RECT 96.355 -53.985 96.495 -53.815 ;
      RECT 96.355 -53.088 96.445 -52.081 ;
      RECT 96.355 -52.775 96.495 -52.605 ;
      RECT 96.355 -51.279 96.445 -50.272 ;
      RECT 96.355 -50.755 96.495 -50.585 ;
      RECT 96.355 -49.858 96.445 -48.851 ;
      RECT 96.355 -49.545 96.495 -49.375 ;
      RECT 96.355 -48.049 96.445 -47.042 ;
      RECT 96.355 -47.525 96.495 -47.355 ;
      RECT 96.355 -46.628 96.445 -45.621 ;
      RECT 96.355 -46.315 96.495 -46.145 ;
      RECT 96.355 -44.819 96.445 -43.812 ;
      RECT 96.355 -44.295 96.495 -44.125 ;
      RECT 96.355 -43.398 96.445 -42.391 ;
      RECT 96.355 -43.085 96.495 -42.915 ;
      RECT 96.355 -41.589 96.445 -40.582 ;
      RECT 96.355 -41.065 96.495 -40.895 ;
      RECT 96.355 -40.168 96.445 -39.161 ;
      RECT 96.355 -39.855 96.495 -39.685 ;
      RECT 96.355 -38.359 96.445 -37.352 ;
      RECT 96.355 -37.835 96.495 -37.665 ;
      RECT 96.355 -36.938 96.445 -35.931 ;
      RECT 96.355 -36.625 96.495 -36.455 ;
      RECT 96.355 -35.129 96.445 -34.122 ;
      RECT 96.355 -34.605 96.495 -34.435 ;
      RECT 96.355 -33.708 96.445 -32.701 ;
      RECT 96.355 -33.395 96.495 -33.225 ;
      RECT 96.355 -31.899 96.445 -30.892 ;
      RECT 96.355 -31.375 96.495 -31.205 ;
      RECT 96.355 -30.478 96.445 -29.471 ;
      RECT 96.355 -30.165 96.495 -29.995 ;
      RECT 96.355 -28.669 96.445 -27.662 ;
      RECT 96.355 -28.145 96.495 -27.975 ;
      RECT 96.355 -27.248 96.445 -26.241 ;
      RECT 96.355 -26.935 96.495 -26.765 ;
      RECT 96.355 -25.439 96.445 -24.432 ;
      RECT 96.355 -24.915 96.495 -24.745 ;
      RECT 96.355 -24.018 96.445 -23.011 ;
      RECT 96.355 -23.705 96.495 -23.535 ;
      RECT 96.355 -22.209 96.445 -21.202 ;
      RECT 96.355 -21.685 96.495 -21.515 ;
      RECT 96.355 -20.788 96.445 -19.781 ;
      RECT 96.355 -20.475 96.495 -20.305 ;
      RECT 96.355 -18.979 96.445 -17.972 ;
      RECT 96.355 -18.455 96.495 -18.285 ;
      RECT 96.355 -17.558 96.445 -16.551 ;
      RECT 96.355 -17.245 96.495 -17.075 ;
      RECT 96.355 -15.749 96.445 -14.742 ;
      RECT 96.355 -15.225 96.495 -15.055 ;
      RECT 96.355 -14.328 96.445 -13.321 ;
      RECT 96.355 -14.015 96.495 -13.845 ;
      RECT 96.355 -12.519 96.445 -11.512 ;
      RECT 96.355 -11.995 96.495 -11.825 ;
      RECT 96.355 -11.098 96.445 -10.091 ;
      RECT 96.355 -10.785 96.495 -10.615 ;
      RECT 96.355 -9.289 96.445 -8.282 ;
      RECT 96.355 -8.765 96.495 -8.595 ;
      RECT 96.355 -7.868 96.445 -6.861 ;
      RECT 96.355 -7.555 96.495 -7.385 ;
      RECT 96.355 -6.059 96.445 -5.052 ;
      RECT 96.355 -5.535 96.495 -5.365 ;
      RECT 96.355 -4.638 96.445 -3.631 ;
      RECT 96.355 -4.325 96.495 -4.155 ;
      RECT 96.355 -2.829 96.445 -1.822 ;
      RECT 96.355 -2.305 96.495 -2.135 ;
      RECT 96.355 -1.408 96.445 -0.401 ;
      RECT 96.355 -1.095 96.495 -0.925 ;
      RECT 96.355 0.401 96.445 1.408 ;
      RECT 96.355 0.925 96.495 1.095 ;
      RECT 92.185 -108.935 95.965 -108.815 ;
      RECT 93.505 -109.475 93.605 -108.815 ;
      RECT 92.945 -109.475 93.045 -108.815 ;
      RECT 92.385 -109.475 92.485 -108.815 ;
      RECT 95.555 -101.538 95.645 -100.53 ;
      RECT 95.505 -100.935 95.645 -100.765 ;
      RECT 95.555 -99.73 95.645 -98.722 ;
      RECT 95.505 -99.495 95.645 -99.325 ;
      RECT 95.555 -98.308 95.645 -97.3 ;
      RECT 95.505 -97.705 95.645 -97.535 ;
      RECT 95.555 -96.5 95.645 -95.492 ;
      RECT 95.505 -96.265 95.645 -96.095 ;
      RECT 95.555 -95.078 95.645 -94.07 ;
      RECT 95.505 -94.475 95.645 -94.305 ;
      RECT 95.555 -93.27 95.645 -92.262 ;
      RECT 95.505 -93.035 95.645 -92.865 ;
      RECT 95.555 -91.848 95.645 -90.84 ;
      RECT 95.505 -91.245 95.645 -91.075 ;
      RECT 95.555 -90.04 95.645 -89.032 ;
      RECT 95.505 -89.805 95.645 -89.635 ;
      RECT 95.555 -88.618 95.645 -87.61 ;
      RECT 95.505 -88.015 95.645 -87.845 ;
      RECT 95.555 -86.81 95.645 -85.802 ;
      RECT 95.505 -86.575 95.645 -86.405 ;
      RECT 95.555 -85.388 95.645 -84.38 ;
      RECT 95.505 -84.785 95.645 -84.615 ;
      RECT 95.555 -83.58 95.645 -82.572 ;
      RECT 95.505 -83.345 95.645 -83.175 ;
      RECT 95.555 -82.158 95.645 -81.15 ;
      RECT 95.505 -81.555 95.645 -81.385 ;
      RECT 95.555 -80.35 95.645 -79.342 ;
      RECT 95.505 -80.115 95.645 -79.945 ;
      RECT 95.555 -78.928 95.645 -77.92 ;
      RECT 95.505 -78.325 95.645 -78.155 ;
      RECT 95.555 -77.12 95.645 -76.112 ;
      RECT 95.505 -76.885 95.645 -76.715 ;
      RECT 95.555 -75.698 95.645 -74.69 ;
      RECT 95.505 -75.095 95.645 -74.925 ;
      RECT 95.555 -73.89 95.645 -72.882 ;
      RECT 95.505 -73.655 95.645 -73.485 ;
      RECT 95.555 -72.468 95.645 -71.46 ;
      RECT 95.505 -71.865 95.645 -71.695 ;
      RECT 95.555 -70.66 95.645 -69.652 ;
      RECT 95.505 -70.425 95.645 -70.255 ;
      RECT 95.555 -69.238 95.645 -68.23 ;
      RECT 95.505 -68.635 95.645 -68.465 ;
      RECT 95.555 -67.43 95.645 -66.422 ;
      RECT 95.505 -67.195 95.645 -67.025 ;
      RECT 95.555 -66.008 95.645 -65 ;
      RECT 95.505 -65.405 95.645 -65.235 ;
      RECT 95.555 -64.2 95.645 -63.192 ;
      RECT 95.505 -63.965 95.645 -63.795 ;
      RECT 95.555 -62.778 95.645 -61.77 ;
      RECT 95.505 -62.175 95.645 -62.005 ;
      RECT 95.555 -60.97 95.645 -59.962 ;
      RECT 95.505 -60.735 95.645 -60.565 ;
      RECT 95.555 -59.548 95.645 -58.54 ;
      RECT 95.505 -58.945 95.645 -58.775 ;
      RECT 95.555 -57.74 95.645 -56.732 ;
      RECT 95.505 -57.505 95.645 -57.335 ;
      RECT 95.555 -56.318 95.645 -55.31 ;
      RECT 95.505 -55.715 95.645 -55.545 ;
      RECT 95.555 -54.51 95.645 -53.502 ;
      RECT 95.505 -54.275 95.645 -54.105 ;
      RECT 95.555 -53.088 95.645 -52.08 ;
      RECT 95.505 -52.485 95.645 -52.315 ;
      RECT 95.555 -51.28 95.645 -50.272 ;
      RECT 95.505 -51.045 95.645 -50.875 ;
      RECT 95.555 -49.858 95.645 -48.85 ;
      RECT 95.505 -49.255 95.645 -49.085 ;
      RECT 95.555 -48.05 95.645 -47.042 ;
      RECT 95.505 -47.815 95.645 -47.645 ;
      RECT 95.555 -46.628 95.645 -45.62 ;
      RECT 95.505 -46.025 95.645 -45.855 ;
      RECT 95.555 -44.82 95.645 -43.812 ;
      RECT 95.505 -44.585 95.645 -44.415 ;
      RECT 95.555 -43.398 95.645 -42.39 ;
      RECT 95.505 -42.795 95.645 -42.625 ;
      RECT 95.555 -41.59 95.645 -40.582 ;
      RECT 95.505 -41.355 95.645 -41.185 ;
      RECT 95.555 -40.168 95.645 -39.16 ;
      RECT 95.505 -39.565 95.645 -39.395 ;
      RECT 95.555 -38.36 95.645 -37.352 ;
      RECT 95.505 -38.125 95.645 -37.955 ;
      RECT 95.555 -36.938 95.645 -35.93 ;
      RECT 95.505 -36.335 95.645 -36.165 ;
      RECT 95.555 -35.13 95.645 -34.122 ;
      RECT 95.505 -34.895 95.645 -34.725 ;
      RECT 95.555 -33.708 95.645 -32.7 ;
      RECT 95.505 -33.105 95.645 -32.935 ;
      RECT 95.555 -31.9 95.645 -30.892 ;
      RECT 95.505 -31.665 95.645 -31.495 ;
      RECT 95.555 -30.478 95.645 -29.47 ;
      RECT 95.505 -29.875 95.645 -29.705 ;
      RECT 95.555 -28.67 95.645 -27.662 ;
      RECT 95.505 -28.435 95.645 -28.265 ;
      RECT 95.555 -27.248 95.645 -26.24 ;
      RECT 95.505 -26.645 95.645 -26.475 ;
      RECT 95.555 -25.44 95.645 -24.432 ;
      RECT 95.505 -25.205 95.645 -25.035 ;
      RECT 95.555 -24.018 95.645 -23.01 ;
      RECT 95.505 -23.415 95.645 -23.245 ;
      RECT 95.555 -22.21 95.645 -21.202 ;
      RECT 95.505 -21.975 95.645 -21.805 ;
      RECT 95.555 -20.788 95.645 -19.78 ;
      RECT 95.505 -20.185 95.645 -20.015 ;
      RECT 95.555 -18.98 95.645 -17.972 ;
      RECT 95.505 -18.745 95.645 -18.575 ;
      RECT 95.555 -17.558 95.645 -16.55 ;
      RECT 95.505 -16.955 95.645 -16.785 ;
      RECT 95.555 -15.75 95.645 -14.742 ;
      RECT 95.505 -15.515 95.645 -15.345 ;
      RECT 95.555 -14.328 95.645 -13.32 ;
      RECT 95.505 -13.725 95.645 -13.555 ;
      RECT 95.555 -12.52 95.645 -11.512 ;
      RECT 95.505 -12.285 95.645 -12.115 ;
      RECT 95.555 -11.098 95.645 -10.09 ;
      RECT 95.505 -10.495 95.645 -10.325 ;
      RECT 95.555 -9.29 95.645 -8.282 ;
      RECT 95.505 -9.055 95.645 -8.885 ;
      RECT 95.555 -7.868 95.645 -6.86 ;
      RECT 95.505 -7.265 95.645 -7.095 ;
      RECT 95.555 -6.06 95.645 -5.052 ;
      RECT 95.505 -5.825 95.645 -5.655 ;
      RECT 95.555 -4.638 95.645 -3.63 ;
      RECT 95.505 -4.035 95.645 -3.865 ;
      RECT 95.555 -2.83 95.645 -1.822 ;
      RECT 95.505 -2.595 95.645 -2.425 ;
      RECT 95.555 -1.408 95.645 -0.4 ;
      RECT 95.505 -0.805 95.645 -0.635 ;
      RECT 95.555 0.4 95.645 1.408 ;
      RECT 95.505 0.635 95.645 0.805 ;
      RECT 94.125 -111.685 95.605 -111.585 ;
      RECT 94.125 -112.195 94.225 -111.585 ;
      RECT 94.345 -109.15 95.605 -109.05 ;
      RECT 95.505 -109.475 95.605 -109.05 ;
      RECT 94.945 -109.475 95.045 -109.05 ;
      RECT 94.385 -109.475 94.485 -109.05 ;
      RECT 95.155 -101.538 95.245 -100.531 ;
      RECT 95.155 -101.225 95.295 -101.055 ;
      RECT 95.155 -99.729 95.245 -98.722 ;
      RECT 95.155 -99.205 95.295 -99.035 ;
      RECT 95.155 -98.308 95.245 -97.301 ;
      RECT 95.155 -97.995 95.295 -97.825 ;
      RECT 95.155 -96.499 95.245 -95.492 ;
      RECT 95.155 -95.975 95.295 -95.805 ;
      RECT 95.155 -95.078 95.245 -94.071 ;
      RECT 95.155 -94.765 95.295 -94.595 ;
      RECT 95.155 -93.269 95.245 -92.262 ;
      RECT 95.155 -92.745 95.295 -92.575 ;
      RECT 95.155 -91.848 95.245 -90.841 ;
      RECT 95.155 -91.535 95.295 -91.365 ;
      RECT 95.155 -90.039 95.245 -89.032 ;
      RECT 95.155 -89.515 95.295 -89.345 ;
      RECT 95.155 -88.618 95.245 -87.611 ;
      RECT 95.155 -88.305 95.295 -88.135 ;
      RECT 95.155 -86.809 95.245 -85.802 ;
      RECT 95.155 -86.285 95.295 -86.115 ;
      RECT 95.155 -85.388 95.245 -84.381 ;
      RECT 95.155 -85.075 95.295 -84.905 ;
      RECT 95.155 -83.579 95.245 -82.572 ;
      RECT 95.155 -83.055 95.295 -82.885 ;
      RECT 95.155 -82.158 95.245 -81.151 ;
      RECT 95.155 -81.845 95.295 -81.675 ;
      RECT 95.155 -80.349 95.245 -79.342 ;
      RECT 95.155 -79.825 95.295 -79.655 ;
      RECT 95.155 -78.928 95.245 -77.921 ;
      RECT 95.155 -78.615 95.295 -78.445 ;
      RECT 95.155 -77.119 95.245 -76.112 ;
      RECT 95.155 -76.595 95.295 -76.425 ;
      RECT 95.155 -75.698 95.245 -74.691 ;
      RECT 95.155 -75.385 95.295 -75.215 ;
      RECT 95.155 -73.889 95.245 -72.882 ;
      RECT 95.155 -73.365 95.295 -73.195 ;
      RECT 95.155 -72.468 95.245 -71.461 ;
      RECT 95.155 -72.155 95.295 -71.985 ;
      RECT 95.155 -70.659 95.245 -69.652 ;
      RECT 95.155 -70.135 95.295 -69.965 ;
      RECT 95.155 -69.238 95.245 -68.231 ;
      RECT 95.155 -68.925 95.295 -68.755 ;
      RECT 95.155 -67.429 95.245 -66.422 ;
      RECT 95.155 -66.905 95.295 -66.735 ;
      RECT 95.155 -66.008 95.245 -65.001 ;
      RECT 95.155 -65.695 95.295 -65.525 ;
      RECT 95.155 -64.199 95.245 -63.192 ;
      RECT 95.155 -63.675 95.295 -63.505 ;
      RECT 95.155 -62.778 95.245 -61.771 ;
      RECT 95.155 -62.465 95.295 -62.295 ;
      RECT 95.155 -60.969 95.245 -59.962 ;
      RECT 95.155 -60.445 95.295 -60.275 ;
      RECT 95.155 -59.548 95.245 -58.541 ;
      RECT 95.155 -59.235 95.295 -59.065 ;
      RECT 95.155 -57.739 95.245 -56.732 ;
      RECT 95.155 -57.215 95.295 -57.045 ;
      RECT 95.155 -56.318 95.245 -55.311 ;
      RECT 95.155 -56.005 95.295 -55.835 ;
      RECT 95.155 -54.509 95.245 -53.502 ;
      RECT 95.155 -53.985 95.295 -53.815 ;
      RECT 95.155 -53.088 95.245 -52.081 ;
      RECT 95.155 -52.775 95.295 -52.605 ;
      RECT 95.155 -51.279 95.245 -50.272 ;
      RECT 95.155 -50.755 95.295 -50.585 ;
      RECT 95.155 -49.858 95.245 -48.851 ;
      RECT 95.155 -49.545 95.295 -49.375 ;
      RECT 95.155 -48.049 95.245 -47.042 ;
      RECT 95.155 -47.525 95.295 -47.355 ;
      RECT 95.155 -46.628 95.245 -45.621 ;
      RECT 95.155 -46.315 95.295 -46.145 ;
      RECT 95.155 -44.819 95.245 -43.812 ;
      RECT 95.155 -44.295 95.295 -44.125 ;
      RECT 95.155 -43.398 95.245 -42.391 ;
      RECT 95.155 -43.085 95.295 -42.915 ;
      RECT 95.155 -41.589 95.245 -40.582 ;
      RECT 95.155 -41.065 95.295 -40.895 ;
      RECT 95.155 -40.168 95.245 -39.161 ;
      RECT 95.155 -39.855 95.295 -39.685 ;
      RECT 95.155 -38.359 95.245 -37.352 ;
      RECT 95.155 -37.835 95.295 -37.665 ;
      RECT 95.155 -36.938 95.245 -35.931 ;
      RECT 95.155 -36.625 95.295 -36.455 ;
      RECT 95.155 -35.129 95.245 -34.122 ;
      RECT 95.155 -34.605 95.295 -34.435 ;
      RECT 95.155 -33.708 95.245 -32.701 ;
      RECT 95.155 -33.395 95.295 -33.225 ;
      RECT 95.155 -31.899 95.245 -30.892 ;
      RECT 95.155 -31.375 95.295 -31.205 ;
      RECT 95.155 -30.478 95.245 -29.471 ;
      RECT 95.155 -30.165 95.295 -29.995 ;
      RECT 95.155 -28.669 95.245 -27.662 ;
      RECT 95.155 -28.145 95.295 -27.975 ;
      RECT 95.155 -27.248 95.245 -26.241 ;
      RECT 95.155 -26.935 95.295 -26.765 ;
      RECT 95.155 -25.439 95.245 -24.432 ;
      RECT 95.155 -24.915 95.295 -24.745 ;
      RECT 95.155 -24.018 95.245 -23.011 ;
      RECT 95.155 -23.705 95.295 -23.535 ;
      RECT 95.155 -22.209 95.245 -21.202 ;
      RECT 95.155 -21.685 95.295 -21.515 ;
      RECT 95.155 -20.788 95.245 -19.781 ;
      RECT 95.155 -20.475 95.295 -20.305 ;
      RECT 95.155 -18.979 95.245 -17.972 ;
      RECT 95.155 -18.455 95.295 -18.285 ;
      RECT 95.155 -17.558 95.245 -16.551 ;
      RECT 95.155 -17.245 95.295 -17.075 ;
      RECT 95.155 -15.749 95.245 -14.742 ;
      RECT 95.155 -15.225 95.295 -15.055 ;
      RECT 95.155 -14.328 95.245 -13.321 ;
      RECT 95.155 -14.015 95.295 -13.845 ;
      RECT 95.155 -12.519 95.245 -11.512 ;
      RECT 95.155 -11.995 95.295 -11.825 ;
      RECT 95.155 -11.098 95.245 -10.091 ;
      RECT 95.155 -10.785 95.295 -10.615 ;
      RECT 95.155 -9.289 95.245 -8.282 ;
      RECT 95.155 -8.765 95.295 -8.595 ;
      RECT 95.155 -7.868 95.245 -6.861 ;
      RECT 95.155 -7.555 95.295 -7.385 ;
      RECT 95.155 -6.059 95.245 -5.052 ;
      RECT 95.155 -5.535 95.295 -5.365 ;
      RECT 95.155 -4.638 95.245 -3.631 ;
      RECT 95.155 -4.325 95.295 -4.155 ;
      RECT 95.155 -2.829 95.245 -1.822 ;
      RECT 95.155 -2.305 95.295 -2.135 ;
      RECT 95.155 -1.408 95.245 -0.401 ;
      RECT 95.155 -1.095 95.295 -0.925 ;
      RECT 95.155 0.401 95.245 1.408 ;
      RECT 95.155 0.925 95.295 1.095 ;
      RECT 94.485 -111.495 94.655 -111.385 ;
      RECT 91.335 -111.495 94.655 -111.395 ;
      RECT 94.355 -101.538 94.445 -100.53 ;
      RECT 94.305 -100.935 94.445 -100.765 ;
      RECT 94.355 -99.73 94.445 -98.722 ;
      RECT 94.305 -99.495 94.445 -99.325 ;
      RECT 94.355 -98.308 94.445 -97.3 ;
      RECT 94.305 -97.705 94.445 -97.535 ;
      RECT 94.355 -96.5 94.445 -95.492 ;
      RECT 94.305 -96.265 94.445 -96.095 ;
      RECT 94.355 -95.078 94.445 -94.07 ;
      RECT 94.305 -94.475 94.445 -94.305 ;
      RECT 94.355 -93.27 94.445 -92.262 ;
      RECT 94.305 -93.035 94.445 -92.865 ;
      RECT 94.355 -91.848 94.445 -90.84 ;
      RECT 94.305 -91.245 94.445 -91.075 ;
      RECT 94.355 -90.04 94.445 -89.032 ;
      RECT 94.305 -89.805 94.445 -89.635 ;
      RECT 94.355 -88.618 94.445 -87.61 ;
      RECT 94.305 -88.015 94.445 -87.845 ;
      RECT 94.355 -86.81 94.445 -85.802 ;
      RECT 94.305 -86.575 94.445 -86.405 ;
      RECT 94.355 -85.388 94.445 -84.38 ;
      RECT 94.305 -84.785 94.445 -84.615 ;
      RECT 94.355 -83.58 94.445 -82.572 ;
      RECT 94.305 -83.345 94.445 -83.175 ;
      RECT 94.355 -82.158 94.445 -81.15 ;
      RECT 94.305 -81.555 94.445 -81.385 ;
      RECT 94.355 -80.35 94.445 -79.342 ;
      RECT 94.305 -80.115 94.445 -79.945 ;
      RECT 94.355 -78.928 94.445 -77.92 ;
      RECT 94.305 -78.325 94.445 -78.155 ;
      RECT 94.355 -77.12 94.445 -76.112 ;
      RECT 94.305 -76.885 94.445 -76.715 ;
      RECT 94.355 -75.698 94.445 -74.69 ;
      RECT 94.305 -75.095 94.445 -74.925 ;
      RECT 94.355 -73.89 94.445 -72.882 ;
      RECT 94.305 -73.655 94.445 -73.485 ;
      RECT 94.355 -72.468 94.445 -71.46 ;
      RECT 94.305 -71.865 94.445 -71.695 ;
      RECT 94.355 -70.66 94.445 -69.652 ;
      RECT 94.305 -70.425 94.445 -70.255 ;
      RECT 94.355 -69.238 94.445 -68.23 ;
      RECT 94.305 -68.635 94.445 -68.465 ;
      RECT 94.355 -67.43 94.445 -66.422 ;
      RECT 94.305 -67.195 94.445 -67.025 ;
      RECT 94.355 -66.008 94.445 -65 ;
      RECT 94.305 -65.405 94.445 -65.235 ;
      RECT 94.355 -64.2 94.445 -63.192 ;
      RECT 94.305 -63.965 94.445 -63.795 ;
      RECT 94.355 -62.778 94.445 -61.77 ;
      RECT 94.305 -62.175 94.445 -62.005 ;
      RECT 94.355 -60.97 94.445 -59.962 ;
      RECT 94.305 -60.735 94.445 -60.565 ;
      RECT 94.355 -59.548 94.445 -58.54 ;
      RECT 94.305 -58.945 94.445 -58.775 ;
      RECT 94.355 -57.74 94.445 -56.732 ;
      RECT 94.305 -57.505 94.445 -57.335 ;
      RECT 94.355 -56.318 94.445 -55.31 ;
      RECT 94.305 -55.715 94.445 -55.545 ;
      RECT 94.355 -54.51 94.445 -53.502 ;
      RECT 94.305 -54.275 94.445 -54.105 ;
      RECT 94.355 -53.088 94.445 -52.08 ;
      RECT 94.305 -52.485 94.445 -52.315 ;
      RECT 94.355 -51.28 94.445 -50.272 ;
      RECT 94.305 -51.045 94.445 -50.875 ;
      RECT 94.355 -49.858 94.445 -48.85 ;
      RECT 94.305 -49.255 94.445 -49.085 ;
      RECT 94.355 -48.05 94.445 -47.042 ;
      RECT 94.305 -47.815 94.445 -47.645 ;
      RECT 94.355 -46.628 94.445 -45.62 ;
      RECT 94.305 -46.025 94.445 -45.855 ;
      RECT 94.355 -44.82 94.445 -43.812 ;
      RECT 94.305 -44.585 94.445 -44.415 ;
      RECT 94.355 -43.398 94.445 -42.39 ;
      RECT 94.305 -42.795 94.445 -42.625 ;
      RECT 94.355 -41.59 94.445 -40.582 ;
      RECT 94.305 -41.355 94.445 -41.185 ;
      RECT 94.355 -40.168 94.445 -39.16 ;
      RECT 94.305 -39.565 94.445 -39.395 ;
      RECT 94.355 -38.36 94.445 -37.352 ;
      RECT 94.305 -38.125 94.445 -37.955 ;
      RECT 94.355 -36.938 94.445 -35.93 ;
      RECT 94.305 -36.335 94.445 -36.165 ;
      RECT 94.355 -35.13 94.445 -34.122 ;
      RECT 94.305 -34.895 94.445 -34.725 ;
      RECT 94.355 -33.708 94.445 -32.7 ;
      RECT 94.305 -33.105 94.445 -32.935 ;
      RECT 94.355 -31.9 94.445 -30.892 ;
      RECT 94.305 -31.665 94.445 -31.495 ;
      RECT 94.355 -30.478 94.445 -29.47 ;
      RECT 94.305 -29.875 94.445 -29.705 ;
      RECT 94.355 -28.67 94.445 -27.662 ;
      RECT 94.305 -28.435 94.445 -28.265 ;
      RECT 94.355 -27.248 94.445 -26.24 ;
      RECT 94.305 -26.645 94.445 -26.475 ;
      RECT 94.355 -25.44 94.445 -24.432 ;
      RECT 94.305 -25.205 94.445 -25.035 ;
      RECT 94.355 -24.018 94.445 -23.01 ;
      RECT 94.305 -23.415 94.445 -23.245 ;
      RECT 94.355 -22.21 94.445 -21.202 ;
      RECT 94.305 -21.975 94.445 -21.805 ;
      RECT 94.355 -20.788 94.445 -19.78 ;
      RECT 94.305 -20.185 94.445 -20.015 ;
      RECT 94.355 -18.98 94.445 -17.972 ;
      RECT 94.305 -18.745 94.445 -18.575 ;
      RECT 94.355 -17.558 94.445 -16.55 ;
      RECT 94.305 -16.955 94.445 -16.785 ;
      RECT 94.355 -15.75 94.445 -14.742 ;
      RECT 94.305 -15.515 94.445 -15.345 ;
      RECT 94.355 -14.328 94.445 -13.32 ;
      RECT 94.305 -13.725 94.445 -13.555 ;
      RECT 94.355 -12.52 94.445 -11.512 ;
      RECT 94.305 -12.285 94.445 -12.115 ;
      RECT 94.355 -11.098 94.445 -10.09 ;
      RECT 94.305 -10.495 94.445 -10.325 ;
      RECT 94.355 -9.29 94.445 -8.282 ;
      RECT 94.305 -9.055 94.445 -8.885 ;
      RECT 94.355 -7.868 94.445 -6.86 ;
      RECT 94.305 -7.265 94.445 -7.095 ;
      RECT 94.355 -6.06 94.445 -5.052 ;
      RECT 94.305 -5.825 94.445 -5.655 ;
      RECT 94.355 -4.638 94.445 -3.63 ;
      RECT 94.305 -4.035 94.445 -3.865 ;
      RECT 94.355 -2.83 94.445 -1.822 ;
      RECT 94.305 -2.595 94.445 -2.425 ;
      RECT 94.355 -1.408 94.445 -0.4 ;
      RECT 94.305 -0.805 94.445 -0.635 ;
      RECT 94.355 0.4 94.445 1.408 ;
      RECT 94.305 0.635 94.445 0.805 ;
      RECT 93.955 -101.538 94.045 -100.531 ;
      RECT 93.955 -101.225 94.095 -101.055 ;
      RECT 93.955 -99.729 94.045 -98.722 ;
      RECT 93.955 -99.205 94.095 -99.035 ;
      RECT 93.955 -98.308 94.045 -97.301 ;
      RECT 93.955 -97.995 94.095 -97.825 ;
      RECT 93.955 -96.499 94.045 -95.492 ;
      RECT 93.955 -95.975 94.095 -95.805 ;
      RECT 93.955 -95.078 94.045 -94.071 ;
      RECT 93.955 -94.765 94.095 -94.595 ;
      RECT 93.955 -93.269 94.045 -92.262 ;
      RECT 93.955 -92.745 94.095 -92.575 ;
      RECT 93.955 -91.848 94.045 -90.841 ;
      RECT 93.955 -91.535 94.095 -91.365 ;
      RECT 93.955 -90.039 94.045 -89.032 ;
      RECT 93.955 -89.515 94.095 -89.345 ;
      RECT 93.955 -88.618 94.045 -87.611 ;
      RECT 93.955 -88.305 94.095 -88.135 ;
      RECT 93.955 -86.809 94.045 -85.802 ;
      RECT 93.955 -86.285 94.095 -86.115 ;
      RECT 93.955 -85.388 94.045 -84.381 ;
      RECT 93.955 -85.075 94.095 -84.905 ;
      RECT 93.955 -83.579 94.045 -82.572 ;
      RECT 93.955 -83.055 94.095 -82.885 ;
      RECT 93.955 -82.158 94.045 -81.151 ;
      RECT 93.955 -81.845 94.095 -81.675 ;
      RECT 93.955 -80.349 94.045 -79.342 ;
      RECT 93.955 -79.825 94.095 -79.655 ;
      RECT 93.955 -78.928 94.045 -77.921 ;
      RECT 93.955 -78.615 94.095 -78.445 ;
      RECT 93.955 -77.119 94.045 -76.112 ;
      RECT 93.955 -76.595 94.095 -76.425 ;
      RECT 93.955 -75.698 94.045 -74.691 ;
      RECT 93.955 -75.385 94.095 -75.215 ;
      RECT 93.955 -73.889 94.045 -72.882 ;
      RECT 93.955 -73.365 94.095 -73.195 ;
      RECT 93.955 -72.468 94.045 -71.461 ;
      RECT 93.955 -72.155 94.095 -71.985 ;
      RECT 93.955 -70.659 94.045 -69.652 ;
      RECT 93.955 -70.135 94.095 -69.965 ;
      RECT 93.955 -69.238 94.045 -68.231 ;
      RECT 93.955 -68.925 94.095 -68.755 ;
      RECT 93.955 -67.429 94.045 -66.422 ;
      RECT 93.955 -66.905 94.095 -66.735 ;
      RECT 93.955 -66.008 94.045 -65.001 ;
      RECT 93.955 -65.695 94.095 -65.525 ;
      RECT 93.955 -64.199 94.045 -63.192 ;
      RECT 93.955 -63.675 94.095 -63.505 ;
      RECT 93.955 -62.778 94.045 -61.771 ;
      RECT 93.955 -62.465 94.095 -62.295 ;
      RECT 93.955 -60.969 94.045 -59.962 ;
      RECT 93.955 -60.445 94.095 -60.275 ;
      RECT 93.955 -59.548 94.045 -58.541 ;
      RECT 93.955 -59.235 94.095 -59.065 ;
      RECT 93.955 -57.739 94.045 -56.732 ;
      RECT 93.955 -57.215 94.095 -57.045 ;
      RECT 93.955 -56.318 94.045 -55.311 ;
      RECT 93.955 -56.005 94.095 -55.835 ;
      RECT 93.955 -54.509 94.045 -53.502 ;
      RECT 93.955 -53.985 94.095 -53.815 ;
      RECT 93.955 -53.088 94.045 -52.081 ;
      RECT 93.955 -52.775 94.095 -52.605 ;
      RECT 93.955 -51.279 94.045 -50.272 ;
      RECT 93.955 -50.755 94.095 -50.585 ;
      RECT 93.955 -49.858 94.045 -48.851 ;
      RECT 93.955 -49.545 94.095 -49.375 ;
      RECT 93.955 -48.049 94.045 -47.042 ;
      RECT 93.955 -47.525 94.095 -47.355 ;
      RECT 93.955 -46.628 94.045 -45.621 ;
      RECT 93.955 -46.315 94.095 -46.145 ;
      RECT 93.955 -44.819 94.045 -43.812 ;
      RECT 93.955 -44.295 94.095 -44.125 ;
      RECT 93.955 -43.398 94.045 -42.391 ;
      RECT 93.955 -43.085 94.095 -42.915 ;
      RECT 93.955 -41.589 94.045 -40.582 ;
      RECT 93.955 -41.065 94.095 -40.895 ;
      RECT 93.955 -40.168 94.045 -39.161 ;
      RECT 93.955 -39.855 94.095 -39.685 ;
      RECT 93.955 -38.359 94.045 -37.352 ;
      RECT 93.955 -37.835 94.095 -37.665 ;
      RECT 93.955 -36.938 94.045 -35.931 ;
      RECT 93.955 -36.625 94.095 -36.455 ;
      RECT 93.955 -35.129 94.045 -34.122 ;
      RECT 93.955 -34.605 94.095 -34.435 ;
      RECT 93.955 -33.708 94.045 -32.701 ;
      RECT 93.955 -33.395 94.095 -33.225 ;
      RECT 93.955 -31.899 94.045 -30.892 ;
      RECT 93.955 -31.375 94.095 -31.205 ;
      RECT 93.955 -30.478 94.045 -29.471 ;
      RECT 93.955 -30.165 94.095 -29.995 ;
      RECT 93.955 -28.669 94.045 -27.662 ;
      RECT 93.955 -28.145 94.095 -27.975 ;
      RECT 93.955 -27.248 94.045 -26.241 ;
      RECT 93.955 -26.935 94.095 -26.765 ;
      RECT 93.955 -25.439 94.045 -24.432 ;
      RECT 93.955 -24.915 94.095 -24.745 ;
      RECT 93.955 -24.018 94.045 -23.011 ;
      RECT 93.955 -23.705 94.095 -23.535 ;
      RECT 93.955 -22.209 94.045 -21.202 ;
      RECT 93.955 -21.685 94.095 -21.515 ;
      RECT 93.955 -20.788 94.045 -19.781 ;
      RECT 93.955 -20.475 94.095 -20.305 ;
      RECT 93.955 -18.979 94.045 -17.972 ;
      RECT 93.955 -18.455 94.095 -18.285 ;
      RECT 93.955 -17.558 94.045 -16.551 ;
      RECT 93.955 -17.245 94.095 -17.075 ;
      RECT 93.955 -15.749 94.045 -14.742 ;
      RECT 93.955 -15.225 94.095 -15.055 ;
      RECT 93.955 -14.328 94.045 -13.321 ;
      RECT 93.955 -14.015 94.095 -13.845 ;
      RECT 93.955 -12.519 94.045 -11.512 ;
      RECT 93.955 -11.995 94.095 -11.825 ;
      RECT 93.955 -11.098 94.045 -10.091 ;
      RECT 93.955 -10.785 94.095 -10.615 ;
      RECT 93.955 -9.289 94.045 -8.282 ;
      RECT 93.955 -8.765 94.095 -8.595 ;
      RECT 93.955 -7.868 94.045 -6.861 ;
      RECT 93.955 -7.555 94.095 -7.385 ;
      RECT 93.955 -6.059 94.045 -5.052 ;
      RECT 93.955 -5.535 94.095 -5.365 ;
      RECT 93.955 -4.638 94.045 -3.631 ;
      RECT 93.955 -4.325 94.095 -4.155 ;
      RECT 93.955 -2.829 94.045 -1.822 ;
      RECT 93.955 -2.305 94.095 -2.135 ;
      RECT 93.955 -1.408 94.045 -0.401 ;
      RECT 93.955 -1.095 94.095 -0.925 ;
      RECT 93.955 0.401 94.045 1.408 ;
      RECT 93.955 0.925 94.095 1.095 ;
      RECT 92.105 -111.685 93.585 -111.585 ;
      RECT 92.105 -112.055 92.205 -111.585 ;
      RECT 91.91 -114.395 93.485 -114.275 ;
      RECT 93.385 -114.895 93.485 -114.275 ;
      RECT 92.79 -114.895 92.89 -114.275 ;
      RECT 91.91 -114.85 92.01 -114.275 ;
      RECT 93.155 -101.538 93.245 -100.53 ;
      RECT 93.105 -100.935 93.245 -100.765 ;
      RECT 93.155 -99.73 93.245 -98.722 ;
      RECT 93.105 -99.495 93.245 -99.325 ;
      RECT 93.155 -98.308 93.245 -97.3 ;
      RECT 93.105 -97.705 93.245 -97.535 ;
      RECT 93.155 -96.5 93.245 -95.492 ;
      RECT 93.105 -96.265 93.245 -96.095 ;
      RECT 93.155 -95.078 93.245 -94.07 ;
      RECT 93.105 -94.475 93.245 -94.305 ;
      RECT 93.155 -93.27 93.245 -92.262 ;
      RECT 93.105 -93.035 93.245 -92.865 ;
      RECT 93.155 -91.848 93.245 -90.84 ;
      RECT 93.105 -91.245 93.245 -91.075 ;
      RECT 93.155 -90.04 93.245 -89.032 ;
      RECT 93.105 -89.805 93.245 -89.635 ;
      RECT 93.155 -88.618 93.245 -87.61 ;
      RECT 93.105 -88.015 93.245 -87.845 ;
      RECT 93.155 -86.81 93.245 -85.802 ;
      RECT 93.105 -86.575 93.245 -86.405 ;
      RECT 93.155 -85.388 93.245 -84.38 ;
      RECT 93.105 -84.785 93.245 -84.615 ;
      RECT 93.155 -83.58 93.245 -82.572 ;
      RECT 93.105 -83.345 93.245 -83.175 ;
      RECT 93.155 -82.158 93.245 -81.15 ;
      RECT 93.105 -81.555 93.245 -81.385 ;
      RECT 93.155 -80.35 93.245 -79.342 ;
      RECT 93.105 -80.115 93.245 -79.945 ;
      RECT 93.155 -78.928 93.245 -77.92 ;
      RECT 93.105 -78.325 93.245 -78.155 ;
      RECT 93.155 -77.12 93.245 -76.112 ;
      RECT 93.105 -76.885 93.245 -76.715 ;
      RECT 93.155 -75.698 93.245 -74.69 ;
      RECT 93.105 -75.095 93.245 -74.925 ;
      RECT 93.155 -73.89 93.245 -72.882 ;
      RECT 93.105 -73.655 93.245 -73.485 ;
      RECT 93.155 -72.468 93.245 -71.46 ;
      RECT 93.105 -71.865 93.245 -71.695 ;
      RECT 93.155 -70.66 93.245 -69.652 ;
      RECT 93.105 -70.425 93.245 -70.255 ;
      RECT 93.155 -69.238 93.245 -68.23 ;
      RECT 93.105 -68.635 93.245 -68.465 ;
      RECT 93.155 -67.43 93.245 -66.422 ;
      RECT 93.105 -67.195 93.245 -67.025 ;
      RECT 93.155 -66.008 93.245 -65 ;
      RECT 93.105 -65.405 93.245 -65.235 ;
      RECT 93.155 -64.2 93.245 -63.192 ;
      RECT 93.105 -63.965 93.245 -63.795 ;
      RECT 93.155 -62.778 93.245 -61.77 ;
      RECT 93.105 -62.175 93.245 -62.005 ;
      RECT 93.155 -60.97 93.245 -59.962 ;
      RECT 93.105 -60.735 93.245 -60.565 ;
      RECT 93.155 -59.548 93.245 -58.54 ;
      RECT 93.105 -58.945 93.245 -58.775 ;
      RECT 93.155 -57.74 93.245 -56.732 ;
      RECT 93.105 -57.505 93.245 -57.335 ;
      RECT 93.155 -56.318 93.245 -55.31 ;
      RECT 93.105 -55.715 93.245 -55.545 ;
      RECT 93.155 -54.51 93.245 -53.502 ;
      RECT 93.105 -54.275 93.245 -54.105 ;
      RECT 93.155 -53.088 93.245 -52.08 ;
      RECT 93.105 -52.485 93.245 -52.315 ;
      RECT 93.155 -51.28 93.245 -50.272 ;
      RECT 93.105 -51.045 93.245 -50.875 ;
      RECT 93.155 -49.858 93.245 -48.85 ;
      RECT 93.105 -49.255 93.245 -49.085 ;
      RECT 93.155 -48.05 93.245 -47.042 ;
      RECT 93.105 -47.815 93.245 -47.645 ;
      RECT 93.155 -46.628 93.245 -45.62 ;
      RECT 93.105 -46.025 93.245 -45.855 ;
      RECT 93.155 -44.82 93.245 -43.812 ;
      RECT 93.105 -44.585 93.245 -44.415 ;
      RECT 93.155 -43.398 93.245 -42.39 ;
      RECT 93.105 -42.795 93.245 -42.625 ;
      RECT 93.155 -41.59 93.245 -40.582 ;
      RECT 93.105 -41.355 93.245 -41.185 ;
      RECT 93.155 -40.168 93.245 -39.16 ;
      RECT 93.105 -39.565 93.245 -39.395 ;
      RECT 93.155 -38.36 93.245 -37.352 ;
      RECT 93.105 -38.125 93.245 -37.955 ;
      RECT 93.155 -36.938 93.245 -35.93 ;
      RECT 93.105 -36.335 93.245 -36.165 ;
      RECT 93.155 -35.13 93.245 -34.122 ;
      RECT 93.105 -34.895 93.245 -34.725 ;
      RECT 93.155 -33.708 93.245 -32.7 ;
      RECT 93.105 -33.105 93.245 -32.935 ;
      RECT 93.155 -31.9 93.245 -30.892 ;
      RECT 93.105 -31.665 93.245 -31.495 ;
      RECT 93.155 -30.478 93.245 -29.47 ;
      RECT 93.105 -29.875 93.245 -29.705 ;
      RECT 93.155 -28.67 93.245 -27.662 ;
      RECT 93.105 -28.435 93.245 -28.265 ;
      RECT 93.155 -27.248 93.245 -26.24 ;
      RECT 93.105 -26.645 93.245 -26.475 ;
      RECT 93.155 -25.44 93.245 -24.432 ;
      RECT 93.105 -25.205 93.245 -25.035 ;
      RECT 93.155 -24.018 93.245 -23.01 ;
      RECT 93.105 -23.415 93.245 -23.245 ;
      RECT 93.155 -22.21 93.245 -21.202 ;
      RECT 93.105 -21.975 93.245 -21.805 ;
      RECT 93.155 -20.788 93.245 -19.78 ;
      RECT 93.105 -20.185 93.245 -20.015 ;
      RECT 93.155 -18.98 93.245 -17.972 ;
      RECT 93.105 -18.745 93.245 -18.575 ;
      RECT 93.155 -17.558 93.245 -16.55 ;
      RECT 93.105 -16.955 93.245 -16.785 ;
      RECT 93.155 -15.75 93.245 -14.742 ;
      RECT 93.105 -15.515 93.245 -15.345 ;
      RECT 93.155 -14.328 93.245 -13.32 ;
      RECT 93.105 -13.725 93.245 -13.555 ;
      RECT 93.155 -12.52 93.245 -11.512 ;
      RECT 93.105 -12.285 93.245 -12.115 ;
      RECT 93.155 -11.098 93.245 -10.09 ;
      RECT 93.105 -10.495 93.245 -10.325 ;
      RECT 93.155 -9.29 93.245 -8.282 ;
      RECT 93.105 -9.055 93.245 -8.885 ;
      RECT 93.155 -7.868 93.245 -6.86 ;
      RECT 93.105 -7.265 93.245 -7.095 ;
      RECT 93.155 -6.06 93.245 -5.052 ;
      RECT 93.105 -5.825 93.245 -5.655 ;
      RECT 93.155 -4.638 93.245 -3.63 ;
      RECT 93.105 -4.035 93.245 -3.865 ;
      RECT 93.155 -2.83 93.245 -1.822 ;
      RECT 93.105 -2.595 93.245 -2.425 ;
      RECT 93.155 -1.408 93.245 -0.4 ;
      RECT 93.105 -0.805 93.245 -0.635 ;
      RECT 93.155 0.4 93.245 1.408 ;
      RECT 93.105 0.635 93.245 0.805 ;
      RECT 93.03 -114.685 93.205 -114.515 ;
      RECT 93.105 -114.895 93.205 -114.515 ;
      RECT 92.145 -113.555 92.245 -113.09 ;
      RECT 92.51 -113.555 92.61 -113.1 ;
      RECT 92.145 -113.555 92.99 -113.385 ;
      RECT 92.755 -101.538 92.845 -100.531 ;
      RECT 92.755 -101.225 92.895 -101.055 ;
      RECT 92.755 -99.729 92.845 -98.722 ;
      RECT 92.755 -99.205 92.895 -99.035 ;
      RECT 92.755 -98.308 92.845 -97.301 ;
      RECT 92.755 -97.995 92.895 -97.825 ;
      RECT 92.755 -96.499 92.845 -95.492 ;
      RECT 92.755 -95.975 92.895 -95.805 ;
      RECT 92.755 -95.078 92.845 -94.071 ;
      RECT 92.755 -94.765 92.895 -94.595 ;
      RECT 92.755 -93.269 92.845 -92.262 ;
      RECT 92.755 -92.745 92.895 -92.575 ;
      RECT 92.755 -91.848 92.845 -90.841 ;
      RECT 92.755 -91.535 92.895 -91.365 ;
      RECT 92.755 -90.039 92.845 -89.032 ;
      RECT 92.755 -89.515 92.895 -89.345 ;
      RECT 92.755 -88.618 92.845 -87.611 ;
      RECT 92.755 -88.305 92.895 -88.135 ;
      RECT 92.755 -86.809 92.845 -85.802 ;
      RECT 92.755 -86.285 92.895 -86.115 ;
      RECT 92.755 -85.388 92.845 -84.381 ;
      RECT 92.755 -85.075 92.895 -84.905 ;
      RECT 92.755 -83.579 92.845 -82.572 ;
      RECT 92.755 -83.055 92.895 -82.885 ;
      RECT 92.755 -82.158 92.845 -81.151 ;
      RECT 92.755 -81.845 92.895 -81.675 ;
      RECT 92.755 -80.349 92.845 -79.342 ;
      RECT 92.755 -79.825 92.895 -79.655 ;
      RECT 92.755 -78.928 92.845 -77.921 ;
      RECT 92.755 -78.615 92.895 -78.445 ;
      RECT 92.755 -77.119 92.845 -76.112 ;
      RECT 92.755 -76.595 92.895 -76.425 ;
      RECT 92.755 -75.698 92.845 -74.691 ;
      RECT 92.755 -75.385 92.895 -75.215 ;
      RECT 92.755 -73.889 92.845 -72.882 ;
      RECT 92.755 -73.365 92.895 -73.195 ;
      RECT 92.755 -72.468 92.845 -71.461 ;
      RECT 92.755 -72.155 92.895 -71.985 ;
      RECT 92.755 -70.659 92.845 -69.652 ;
      RECT 92.755 -70.135 92.895 -69.965 ;
      RECT 92.755 -69.238 92.845 -68.231 ;
      RECT 92.755 -68.925 92.895 -68.755 ;
      RECT 92.755 -67.429 92.845 -66.422 ;
      RECT 92.755 -66.905 92.895 -66.735 ;
      RECT 92.755 -66.008 92.845 -65.001 ;
      RECT 92.755 -65.695 92.895 -65.525 ;
      RECT 92.755 -64.199 92.845 -63.192 ;
      RECT 92.755 -63.675 92.895 -63.505 ;
      RECT 92.755 -62.778 92.845 -61.771 ;
      RECT 92.755 -62.465 92.895 -62.295 ;
      RECT 92.755 -60.969 92.845 -59.962 ;
      RECT 92.755 -60.445 92.895 -60.275 ;
      RECT 92.755 -59.548 92.845 -58.541 ;
      RECT 92.755 -59.235 92.895 -59.065 ;
      RECT 92.755 -57.739 92.845 -56.732 ;
      RECT 92.755 -57.215 92.895 -57.045 ;
      RECT 92.755 -56.318 92.845 -55.311 ;
      RECT 92.755 -56.005 92.895 -55.835 ;
      RECT 92.755 -54.509 92.845 -53.502 ;
      RECT 92.755 -53.985 92.895 -53.815 ;
      RECT 92.755 -53.088 92.845 -52.081 ;
      RECT 92.755 -52.775 92.895 -52.605 ;
      RECT 92.755 -51.279 92.845 -50.272 ;
      RECT 92.755 -50.755 92.895 -50.585 ;
      RECT 92.755 -49.858 92.845 -48.851 ;
      RECT 92.755 -49.545 92.895 -49.375 ;
      RECT 92.755 -48.049 92.845 -47.042 ;
      RECT 92.755 -47.525 92.895 -47.355 ;
      RECT 92.755 -46.628 92.845 -45.621 ;
      RECT 92.755 -46.315 92.895 -46.145 ;
      RECT 92.755 -44.819 92.845 -43.812 ;
      RECT 92.755 -44.295 92.895 -44.125 ;
      RECT 92.755 -43.398 92.845 -42.391 ;
      RECT 92.755 -43.085 92.895 -42.915 ;
      RECT 92.755 -41.589 92.845 -40.582 ;
      RECT 92.755 -41.065 92.895 -40.895 ;
      RECT 92.755 -40.168 92.845 -39.161 ;
      RECT 92.755 -39.855 92.895 -39.685 ;
      RECT 92.755 -38.359 92.845 -37.352 ;
      RECT 92.755 -37.835 92.895 -37.665 ;
      RECT 92.755 -36.938 92.845 -35.931 ;
      RECT 92.755 -36.625 92.895 -36.455 ;
      RECT 92.755 -35.129 92.845 -34.122 ;
      RECT 92.755 -34.605 92.895 -34.435 ;
      RECT 92.755 -33.708 92.845 -32.701 ;
      RECT 92.755 -33.395 92.895 -33.225 ;
      RECT 92.755 -31.899 92.845 -30.892 ;
      RECT 92.755 -31.375 92.895 -31.205 ;
      RECT 92.755 -30.478 92.845 -29.471 ;
      RECT 92.755 -30.165 92.895 -29.995 ;
      RECT 92.755 -28.669 92.845 -27.662 ;
      RECT 92.755 -28.145 92.895 -27.975 ;
      RECT 92.755 -27.248 92.845 -26.241 ;
      RECT 92.755 -26.935 92.895 -26.765 ;
      RECT 92.755 -25.439 92.845 -24.432 ;
      RECT 92.755 -24.915 92.895 -24.745 ;
      RECT 92.755 -24.018 92.845 -23.011 ;
      RECT 92.755 -23.705 92.895 -23.535 ;
      RECT 92.755 -22.209 92.845 -21.202 ;
      RECT 92.755 -21.685 92.895 -21.515 ;
      RECT 92.755 -20.788 92.845 -19.781 ;
      RECT 92.755 -20.475 92.895 -20.305 ;
      RECT 92.755 -18.979 92.845 -17.972 ;
      RECT 92.755 -18.455 92.895 -18.285 ;
      RECT 92.755 -17.558 92.845 -16.551 ;
      RECT 92.755 -17.245 92.895 -17.075 ;
      RECT 92.755 -15.749 92.845 -14.742 ;
      RECT 92.755 -15.225 92.895 -15.055 ;
      RECT 92.755 -14.328 92.845 -13.321 ;
      RECT 92.755 -14.015 92.895 -13.845 ;
      RECT 92.755 -12.519 92.845 -11.512 ;
      RECT 92.755 -11.995 92.895 -11.825 ;
      RECT 92.755 -11.098 92.845 -10.091 ;
      RECT 92.755 -10.785 92.895 -10.615 ;
      RECT 92.755 -9.289 92.845 -8.282 ;
      RECT 92.755 -8.765 92.895 -8.595 ;
      RECT 92.755 -7.868 92.845 -6.861 ;
      RECT 92.755 -7.555 92.895 -7.385 ;
      RECT 92.755 -6.059 92.845 -5.052 ;
      RECT 92.755 -5.535 92.895 -5.365 ;
      RECT 92.755 -4.638 92.845 -3.631 ;
      RECT 92.755 -4.325 92.895 -4.155 ;
      RECT 92.755 -2.829 92.845 -1.822 ;
      RECT 92.755 -2.305 92.895 -2.135 ;
      RECT 92.755 -1.408 92.845 -0.401 ;
      RECT 92.755 -1.095 92.895 -0.925 ;
      RECT 92.755 0.401 92.845 1.408 ;
      RECT 92.755 0.925 92.895 1.095 ;
      RECT 92.44 -114.685 92.61 -114.515 ;
      RECT 92.51 -114.895 92.61 -114.515 ;
      RECT 91.955 -101.538 92.045 -100.53 ;
      RECT 91.905 -100.935 92.045 -100.765 ;
      RECT 91.955 -99.73 92.045 -98.722 ;
      RECT 91.905 -99.495 92.045 -99.325 ;
      RECT 91.955 -98.308 92.045 -97.3 ;
      RECT 91.905 -97.705 92.045 -97.535 ;
      RECT 91.955 -96.5 92.045 -95.492 ;
      RECT 91.905 -96.265 92.045 -96.095 ;
      RECT 91.955 -95.078 92.045 -94.07 ;
      RECT 91.905 -94.475 92.045 -94.305 ;
      RECT 91.955 -93.27 92.045 -92.262 ;
      RECT 91.905 -93.035 92.045 -92.865 ;
      RECT 91.955 -91.848 92.045 -90.84 ;
      RECT 91.905 -91.245 92.045 -91.075 ;
      RECT 91.955 -90.04 92.045 -89.032 ;
      RECT 91.905 -89.805 92.045 -89.635 ;
      RECT 91.955 -88.618 92.045 -87.61 ;
      RECT 91.905 -88.015 92.045 -87.845 ;
      RECT 91.955 -86.81 92.045 -85.802 ;
      RECT 91.905 -86.575 92.045 -86.405 ;
      RECT 91.955 -85.388 92.045 -84.38 ;
      RECT 91.905 -84.785 92.045 -84.615 ;
      RECT 91.955 -83.58 92.045 -82.572 ;
      RECT 91.905 -83.345 92.045 -83.175 ;
      RECT 91.955 -82.158 92.045 -81.15 ;
      RECT 91.905 -81.555 92.045 -81.385 ;
      RECT 91.955 -80.35 92.045 -79.342 ;
      RECT 91.905 -80.115 92.045 -79.945 ;
      RECT 91.955 -78.928 92.045 -77.92 ;
      RECT 91.905 -78.325 92.045 -78.155 ;
      RECT 91.955 -77.12 92.045 -76.112 ;
      RECT 91.905 -76.885 92.045 -76.715 ;
      RECT 91.955 -75.698 92.045 -74.69 ;
      RECT 91.905 -75.095 92.045 -74.925 ;
      RECT 91.955 -73.89 92.045 -72.882 ;
      RECT 91.905 -73.655 92.045 -73.485 ;
      RECT 91.955 -72.468 92.045 -71.46 ;
      RECT 91.905 -71.865 92.045 -71.695 ;
      RECT 91.955 -70.66 92.045 -69.652 ;
      RECT 91.905 -70.425 92.045 -70.255 ;
      RECT 91.955 -69.238 92.045 -68.23 ;
      RECT 91.905 -68.635 92.045 -68.465 ;
      RECT 91.955 -67.43 92.045 -66.422 ;
      RECT 91.905 -67.195 92.045 -67.025 ;
      RECT 91.955 -66.008 92.045 -65 ;
      RECT 91.905 -65.405 92.045 -65.235 ;
      RECT 91.955 -64.2 92.045 -63.192 ;
      RECT 91.905 -63.965 92.045 -63.795 ;
      RECT 91.955 -62.778 92.045 -61.77 ;
      RECT 91.905 -62.175 92.045 -62.005 ;
      RECT 91.955 -60.97 92.045 -59.962 ;
      RECT 91.905 -60.735 92.045 -60.565 ;
      RECT 91.955 -59.548 92.045 -58.54 ;
      RECT 91.905 -58.945 92.045 -58.775 ;
      RECT 91.955 -57.74 92.045 -56.732 ;
      RECT 91.905 -57.505 92.045 -57.335 ;
      RECT 91.955 -56.318 92.045 -55.31 ;
      RECT 91.905 -55.715 92.045 -55.545 ;
      RECT 91.955 -54.51 92.045 -53.502 ;
      RECT 91.905 -54.275 92.045 -54.105 ;
      RECT 91.955 -53.088 92.045 -52.08 ;
      RECT 91.905 -52.485 92.045 -52.315 ;
      RECT 91.955 -51.28 92.045 -50.272 ;
      RECT 91.905 -51.045 92.045 -50.875 ;
      RECT 91.955 -49.858 92.045 -48.85 ;
      RECT 91.905 -49.255 92.045 -49.085 ;
      RECT 91.955 -48.05 92.045 -47.042 ;
      RECT 91.905 -47.815 92.045 -47.645 ;
      RECT 91.955 -46.628 92.045 -45.62 ;
      RECT 91.905 -46.025 92.045 -45.855 ;
      RECT 91.955 -44.82 92.045 -43.812 ;
      RECT 91.905 -44.585 92.045 -44.415 ;
      RECT 91.955 -43.398 92.045 -42.39 ;
      RECT 91.905 -42.795 92.045 -42.625 ;
      RECT 91.955 -41.59 92.045 -40.582 ;
      RECT 91.905 -41.355 92.045 -41.185 ;
      RECT 91.955 -40.168 92.045 -39.16 ;
      RECT 91.905 -39.565 92.045 -39.395 ;
      RECT 91.955 -38.36 92.045 -37.352 ;
      RECT 91.905 -38.125 92.045 -37.955 ;
      RECT 91.955 -36.938 92.045 -35.93 ;
      RECT 91.905 -36.335 92.045 -36.165 ;
      RECT 91.955 -35.13 92.045 -34.122 ;
      RECT 91.905 -34.895 92.045 -34.725 ;
      RECT 91.955 -33.708 92.045 -32.7 ;
      RECT 91.905 -33.105 92.045 -32.935 ;
      RECT 91.955 -31.9 92.045 -30.892 ;
      RECT 91.905 -31.665 92.045 -31.495 ;
      RECT 91.955 -30.478 92.045 -29.47 ;
      RECT 91.905 -29.875 92.045 -29.705 ;
      RECT 91.955 -28.67 92.045 -27.662 ;
      RECT 91.905 -28.435 92.045 -28.265 ;
      RECT 91.955 -27.248 92.045 -26.24 ;
      RECT 91.905 -26.645 92.045 -26.475 ;
      RECT 91.955 -25.44 92.045 -24.432 ;
      RECT 91.905 -25.205 92.045 -25.035 ;
      RECT 91.955 -24.018 92.045 -23.01 ;
      RECT 91.905 -23.415 92.045 -23.245 ;
      RECT 91.955 -22.21 92.045 -21.202 ;
      RECT 91.905 -21.975 92.045 -21.805 ;
      RECT 91.955 -20.788 92.045 -19.78 ;
      RECT 91.905 -20.185 92.045 -20.015 ;
      RECT 91.955 -18.98 92.045 -17.972 ;
      RECT 91.905 -18.745 92.045 -18.575 ;
      RECT 91.955 -17.558 92.045 -16.55 ;
      RECT 91.905 -16.955 92.045 -16.785 ;
      RECT 91.955 -15.75 92.045 -14.742 ;
      RECT 91.905 -15.515 92.045 -15.345 ;
      RECT 91.955 -14.328 92.045 -13.32 ;
      RECT 91.905 -13.725 92.045 -13.555 ;
      RECT 91.955 -12.52 92.045 -11.512 ;
      RECT 91.905 -12.285 92.045 -12.115 ;
      RECT 91.955 -11.098 92.045 -10.09 ;
      RECT 91.905 -10.495 92.045 -10.325 ;
      RECT 91.955 -9.29 92.045 -8.282 ;
      RECT 91.905 -9.055 92.045 -8.885 ;
      RECT 91.955 -7.868 92.045 -6.86 ;
      RECT 91.905 -7.265 92.045 -7.095 ;
      RECT 91.955 -6.06 92.045 -5.052 ;
      RECT 91.905 -5.825 92.045 -5.655 ;
      RECT 91.955 -4.638 92.045 -3.63 ;
      RECT 91.905 -4.035 92.045 -3.865 ;
      RECT 91.955 -2.83 92.045 -1.822 ;
      RECT 91.905 -2.595 92.045 -2.425 ;
      RECT 91.955 -1.408 92.045 -0.4 ;
      RECT 91.905 -0.805 92.045 -0.635 ;
      RECT 91.955 0.4 92.045 1.408 ;
      RECT 91.905 0.635 92.045 0.805 ;
      RECT 91.555 -101.538 91.645 -100.531 ;
      RECT 91.555 -101.225 91.695 -101.055 ;
      RECT 91.555 -99.729 91.645 -98.722 ;
      RECT 91.555 -99.205 91.695 -99.035 ;
      RECT 91.555 -98.308 91.645 -97.301 ;
      RECT 91.555 -97.995 91.695 -97.825 ;
      RECT 91.555 -96.499 91.645 -95.492 ;
      RECT 91.555 -95.975 91.695 -95.805 ;
      RECT 91.555 -95.078 91.645 -94.071 ;
      RECT 91.555 -94.765 91.695 -94.595 ;
      RECT 91.555 -93.269 91.645 -92.262 ;
      RECT 91.555 -92.745 91.695 -92.575 ;
      RECT 91.555 -91.848 91.645 -90.841 ;
      RECT 91.555 -91.535 91.695 -91.365 ;
      RECT 91.555 -90.039 91.645 -89.032 ;
      RECT 91.555 -89.515 91.695 -89.345 ;
      RECT 91.555 -88.618 91.645 -87.611 ;
      RECT 91.555 -88.305 91.695 -88.135 ;
      RECT 91.555 -86.809 91.645 -85.802 ;
      RECT 91.555 -86.285 91.695 -86.115 ;
      RECT 91.555 -85.388 91.645 -84.381 ;
      RECT 91.555 -85.075 91.695 -84.905 ;
      RECT 91.555 -83.579 91.645 -82.572 ;
      RECT 91.555 -83.055 91.695 -82.885 ;
      RECT 91.555 -82.158 91.645 -81.151 ;
      RECT 91.555 -81.845 91.695 -81.675 ;
      RECT 91.555 -80.349 91.645 -79.342 ;
      RECT 91.555 -79.825 91.695 -79.655 ;
      RECT 91.555 -78.928 91.645 -77.921 ;
      RECT 91.555 -78.615 91.695 -78.445 ;
      RECT 91.555 -77.119 91.645 -76.112 ;
      RECT 91.555 -76.595 91.695 -76.425 ;
      RECT 91.555 -75.698 91.645 -74.691 ;
      RECT 91.555 -75.385 91.695 -75.215 ;
      RECT 91.555 -73.889 91.645 -72.882 ;
      RECT 91.555 -73.365 91.695 -73.195 ;
      RECT 91.555 -72.468 91.645 -71.461 ;
      RECT 91.555 -72.155 91.695 -71.985 ;
      RECT 91.555 -70.659 91.645 -69.652 ;
      RECT 91.555 -70.135 91.695 -69.965 ;
      RECT 91.555 -69.238 91.645 -68.231 ;
      RECT 91.555 -68.925 91.695 -68.755 ;
      RECT 91.555 -67.429 91.645 -66.422 ;
      RECT 91.555 -66.905 91.695 -66.735 ;
      RECT 91.555 -66.008 91.645 -65.001 ;
      RECT 91.555 -65.695 91.695 -65.525 ;
      RECT 91.555 -64.199 91.645 -63.192 ;
      RECT 91.555 -63.675 91.695 -63.505 ;
      RECT 91.555 -62.778 91.645 -61.771 ;
      RECT 91.555 -62.465 91.695 -62.295 ;
      RECT 91.555 -60.969 91.645 -59.962 ;
      RECT 91.555 -60.445 91.695 -60.275 ;
      RECT 91.555 -59.548 91.645 -58.541 ;
      RECT 91.555 -59.235 91.695 -59.065 ;
      RECT 91.555 -57.739 91.645 -56.732 ;
      RECT 91.555 -57.215 91.695 -57.045 ;
      RECT 91.555 -56.318 91.645 -55.311 ;
      RECT 91.555 -56.005 91.695 -55.835 ;
      RECT 91.555 -54.509 91.645 -53.502 ;
      RECT 91.555 -53.985 91.695 -53.815 ;
      RECT 91.555 -53.088 91.645 -52.081 ;
      RECT 91.555 -52.775 91.695 -52.605 ;
      RECT 91.555 -51.279 91.645 -50.272 ;
      RECT 91.555 -50.755 91.695 -50.585 ;
      RECT 91.555 -49.858 91.645 -48.851 ;
      RECT 91.555 -49.545 91.695 -49.375 ;
      RECT 91.555 -48.049 91.645 -47.042 ;
      RECT 91.555 -47.525 91.695 -47.355 ;
      RECT 91.555 -46.628 91.645 -45.621 ;
      RECT 91.555 -46.315 91.695 -46.145 ;
      RECT 91.555 -44.819 91.645 -43.812 ;
      RECT 91.555 -44.295 91.695 -44.125 ;
      RECT 91.555 -43.398 91.645 -42.391 ;
      RECT 91.555 -43.085 91.695 -42.915 ;
      RECT 91.555 -41.589 91.645 -40.582 ;
      RECT 91.555 -41.065 91.695 -40.895 ;
      RECT 91.555 -40.168 91.645 -39.161 ;
      RECT 91.555 -39.855 91.695 -39.685 ;
      RECT 91.555 -38.359 91.645 -37.352 ;
      RECT 91.555 -37.835 91.695 -37.665 ;
      RECT 91.555 -36.938 91.645 -35.931 ;
      RECT 91.555 -36.625 91.695 -36.455 ;
      RECT 91.555 -35.129 91.645 -34.122 ;
      RECT 91.555 -34.605 91.695 -34.435 ;
      RECT 91.555 -33.708 91.645 -32.701 ;
      RECT 91.555 -33.395 91.695 -33.225 ;
      RECT 91.555 -31.899 91.645 -30.892 ;
      RECT 91.555 -31.375 91.695 -31.205 ;
      RECT 91.555 -30.478 91.645 -29.471 ;
      RECT 91.555 -30.165 91.695 -29.995 ;
      RECT 91.555 -28.669 91.645 -27.662 ;
      RECT 91.555 -28.145 91.695 -27.975 ;
      RECT 91.555 -27.248 91.645 -26.241 ;
      RECT 91.555 -26.935 91.695 -26.765 ;
      RECT 91.555 -25.439 91.645 -24.432 ;
      RECT 91.555 -24.915 91.695 -24.745 ;
      RECT 91.555 -24.018 91.645 -23.011 ;
      RECT 91.555 -23.705 91.695 -23.535 ;
      RECT 91.555 -22.209 91.645 -21.202 ;
      RECT 91.555 -21.685 91.695 -21.515 ;
      RECT 91.555 -20.788 91.645 -19.781 ;
      RECT 91.555 -20.475 91.695 -20.305 ;
      RECT 91.555 -18.979 91.645 -17.972 ;
      RECT 91.555 -18.455 91.695 -18.285 ;
      RECT 91.555 -17.558 91.645 -16.551 ;
      RECT 91.555 -17.245 91.695 -17.075 ;
      RECT 91.555 -15.749 91.645 -14.742 ;
      RECT 91.555 -15.225 91.695 -15.055 ;
      RECT 91.555 -14.328 91.645 -13.321 ;
      RECT 91.555 -14.015 91.695 -13.845 ;
      RECT 91.555 -12.519 91.645 -11.512 ;
      RECT 91.555 -11.995 91.695 -11.825 ;
      RECT 91.555 -11.098 91.645 -10.091 ;
      RECT 91.555 -10.785 91.695 -10.615 ;
      RECT 91.555 -9.289 91.645 -8.282 ;
      RECT 91.555 -8.765 91.695 -8.595 ;
      RECT 91.555 -7.868 91.645 -6.861 ;
      RECT 91.555 -7.555 91.695 -7.385 ;
      RECT 91.555 -6.059 91.645 -5.052 ;
      RECT 91.555 -5.535 91.695 -5.365 ;
      RECT 91.555 -4.638 91.645 -3.631 ;
      RECT 91.555 -4.325 91.695 -4.155 ;
      RECT 91.555 -2.829 91.645 -1.822 ;
      RECT 91.555 -2.305 91.695 -2.135 ;
      RECT 91.555 -1.408 91.645 -0.401 ;
      RECT 91.555 -1.095 91.695 -0.925 ;
      RECT 91.555 0.401 91.645 1.408 ;
      RECT 91.555 0.925 91.695 1.095 ;
      RECT 87.385 -108.935 91.165 -108.815 ;
      RECT 88.705 -109.475 88.805 -108.815 ;
      RECT 88.145 -109.475 88.245 -108.815 ;
      RECT 87.585 -109.475 87.685 -108.815 ;
      RECT 90.755 -101.538 90.845 -100.53 ;
      RECT 90.705 -100.935 90.845 -100.765 ;
      RECT 90.755 -99.73 90.845 -98.722 ;
      RECT 90.705 -99.495 90.845 -99.325 ;
      RECT 90.755 -98.308 90.845 -97.3 ;
      RECT 90.705 -97.705 90.845 -97.535 ;
      RECT 90.755 -96.5 90.845 -95.492 ;
      RECT 90.705 -96.265 90.845 -96.095 ;
      RECT 90.755 -95.078 90.845 -94.07 ;
      RECT 90.705 -94.475 90.845 -94.305 ;
      RECT 90.755 -93.27 90.845 -92.262 ;
      RECT 90.705 -93.035 90.845 -92.865 ;
      RECT 90.755 -91.848 90.845 -90.84 ;
      RECT 90.705 -91.245 90.845 -91.075 ;
      RECT 90.755 -90.04 90.845 -89.032 ;
      RECT 90.705 -89.805 90.845 -89.635 ;
      RECT 90.755 -88.618 90.845 -87.61 ;
      RECT 90.705 -88.015 90.845 -87.845 ;
      RECT 90.755 -86.81 90.845 -85.802 ;
      RECT 90.705 -86.575 90.845 -86.405 ;
      RECT 90.755 -85.388 90.845 -84.38 ;
      RECT 90.705 -84.785 90.845 -84.615 ;
      RECT 90.755 -83.58 90.845 -82.572 ;
      RECT 90.705 -83.345 90.845 -83.175 ;
      RECT 90.755 -82.158 90.845 -81.15 ;
      RECT 90.705 -81.555 90.845 -81.385 ;
      RECT 90.755 -80.35 90.845 -79.342 ;
      RECT 90.705 -80.115 90.845 -79.945 ;
      RECT 90.755 -78.928 90.845 -77.92 ;
      RECT 90.705 -78.325 90.845 -78.155 ;
      RECT 90.755 -77.12 90.845 -76.112 ;
      RECT 90.705 -76.885 90.845 -76.715 ;
      RECT 90.755 -75.698 90.845 -74.69 ;
      RECT 90.705 -75.095 90.845 -74.925 ;
      RECT 90.755 -73.89 90.845 -72.882 ;
      RECT 90.705 -73.655 90.845 -73.485 ;
      RECT 90.755 -72.468 90.845 -71.46 ;
      RECT 90.705 -71.865 90.845 -71.695 ;
      RECT 90.755 -70.66 90.845 -69.652 ;
      RECT 90.705 -70.425 90.845 -70.255 ;
      RECT 90.755 -69.238 90.845 -68.23 ;
      RECT 90.705 -68.635 90.845 -68.465 ;
      RECT 90.755 -67.43 90.845 -66.422 ;
      RECT 90.705 -67.195 90.845 -67.025 ;
      RECT 90.755 -66.008 90.845 -65 ;
      RECT 90.705 -65.405 90.845 -65.235 ;
      RECT 90.755 -64.2 90.845 -63.192 ;
      RECT 90.705 -63.965 90.845 -63.795 ;
      RECT 90.755 -62.778 90.845 -61.77 ;
      RECT 90.705 -62.175 90.845 -62.005 ;
      RECT 90.755 -60.97 90.845 -59.962 ;
      RECT 90.705 -60.735 90.845 -60.565 ;
      RECT 90.755 -59.548 90.845 -58.54 ;
      RECT 90.705 -58.945 90.845 -58.775 ;
      RECT 90.755 -57.74 90.845 -56.732 ;
      RECT 90.705 -57.505 90.845 -57.335 ;
      RECT 90.755 -56.318 90.845 -55.31 ;
      RECT 90.705 -55.715 90.845 -55.545 ;
      RECT 90.755 -54.51 90.845 -53.502 ;
      RECT 90.705 -54.275 90.845 -54.105 ;
      RECT 90.755 -53.088 90.845 -52.08 ;
      RECT 90.705 -52.485 90.845 -52.315 ;
      RECT 90.755 -51.28 90.845 -50.272 ;
      RECT 90.705 -51.045 90.845 -50.875 ;
      RECT 90.755 -49.858 90.845 -48.85 ;
      RECT 90.705 -49.255 90.845 -49.085 ;
      RECT 90.755 -48.05 90.845 -47.042 ;
      RECT 90.705 -47.815 90.845 -47.645 ;
      RECT 90.755 -46.628 90.845 -45.62 ;
      RECT 90.705 -46.025 90.845 -45.855 ;
      RECT 90.755 -44.82 90.845 -43.812 ;
      RECT 90.705 -44.585 90.845 -44.415 ;
      RECT 90.755 -43.398 90.845 -42.39 ;
      RECT 90.705 -42.795 90.845 -42.625 ;
      RECT 90.755 -41.59 90.845 -40.582 ;
      RECT 90.705 -41.355 90.845 -41.185 ;
      RECT 90.755 -40.168 90.845 -39.16 ;
      RECT 90.705 -39.565 90.845 -39.395 ;
      RECT 90.755 -38.36 90.845 -37.352 ;
      RECT 90.705 -38.125 90.845 -37.955 ;
      RECT 90.755 -36.938 90.845 -35.93 ;
      RECT 90.705 -36.335 90.845 -36.165 ;
      RECT 90.755 -35.13 90.845 -34.122 ;
      RECT 90.705 -34.895 90.845 -34.725 ;
      RECT 90.755 -33.708 90.845 -32.7 ;
      RECT 90.705 -33.105 90.845 -32.935 ;
      RECT 90.755 -31.9 90.845 -30.892 ;
      RECT 90.705 -31.665 90.845 -31.495 ;
      RECT 90.755 -30.478 90.845 -29.47 ;
      RECT 90.705 -29.875 90.845 -29.705 ;
      RECT 90.755 -28.67 90.845 -27.662 ;
      RECT 90.705 -28.435 90.845 -28.265 ;
      RECT 90.755 -27.248 90.845 -26.24 ;
      RECT 90.705 -26.645 90.845 -26.475 ;
      RECT 90.755 -25.44 90.845 -24.432 ;
      RECT 90.705 -25.205 90.845 -25.035 ;
      RECT 90.755 -24.018 90.845 -23.01 ;
      RECT 90.705 -23.415 90.845 -23.245 ;
      RECT 90.755 -22.21 90.845 -21.202 ;
      RECT 90.705 -21.975 90.845 -21.805 ;
      RECT 90.755 -20.788 90.845 -19.78 ;
      RECT 90.705 -20.185 90.845 -20.015 ;
      RECT 90.755 -18.98 90.845 -17.972 ;
      RECT 90.705 -18.745 90.845 -18.575 ;
      RECT 90.755 -17.558 90.845 -16.55 ;
      RECT 90.705 -16.955 90.845 -16.785 ;
      RECT 90.755 -15.75 90.845 -14.742 ;
      RECT 90.705 -15.515 90.845 -15.345 ;
      RECT 90.755 -14.328 90.845 -13.32 ;
      RECT 90.705 -13.725 90.845 -13.555 ;
      RECT 90.755 -12.52 90.845 -11.512 ;
      RECT 90.705 -12.285 90.845 -12.115 ;
      RECT 90.755 -11.098 90.845 -10.09 ;
      RECT 90.705 -10.495 90.845 -10.325 ;
      RECT 90.755 -9.29 90.845 -8.282 ;
      RECT 90.705 -9.055 90.845 -8.885 ;
      RECT 90.755 -7.868 90.845 -6.86 ;
      RECT 90.705 -7.265 90.845 -7.095 ;
      RECT 90.755 -6.06 90.845 -5.052 ;
      RECT 90.705 -5.825 90.845 -5.655 ;
      RECT 90.755 -4.638 90.845 -3.63 ;
      RECT 90.705 -4.035 90.845 -3.865 ;
      RECT 90.755 -2.83 90.845 -1.822 ;
      RECT 90.705 -2.595 90.845 -2.425 ;
      RECT 90.755 -1.408 90.845 -0.4 ;
      RECT 90.705 -0.805 90.845 -0.635 ;
      RECT 90.755 0.4 90.845 1.408 ;
      RECT 90.705 0.635 90.845 0.805 ;
      RECT 89.325 -111.685 90.805 -111.585 ;
      RECT 89.325 -112.195 89.425 -111.585 ;
      RECT 89.545 -109.15 90.805 -109.05 ;
      RECT 90.705 -109.475 90.805 -109.05 ;
      RECT 90.145 -109.475 90.245 -109.05 ;
      RECT 89.585 -109.475 89.685 -109.05 ;
      RECT 90.355 -101.538 90.445 -100.531 ;
      RECT 90.355 -101.225 90.495 -101.055 ;
      RECT 90.355 -99.729 90.445 -98.722 ;
      RECT 90.355 -99.205 90.495 -99.035 ;
      RECT 90.355 -98.308 90.445 -97.301 ;
      RECT 90.355 -97.995 90.495 -97.825 ;
      RECT 90.355 -96.499 90.445 -95.492 ;
      RECT 90.355 -95.975 90.495 -95.805 ;
      RECT 90.355 -95.078 90.445 -94.071 ;
      RECT 90.355 -94.765 90.495 -94.595 ;
      RECT 90.355 -93.269 90.445 -92.262 ;
      RECT 90.355 -92.745 90.495 -92.575 ;
      RECT 90.355 -91.848 90.445 -90.841 ;
      RECT 90.355 -91.535 90.495 -91.365 ;
      RECT 90.355 -90.039 90.445 -89.032 ;
      RECT 90.355 -89.515 90.495 -89.345 ;
      RECT 90.355 -88.618 90.445 -87.611 ;
      RECT 90.355 -88.305 90.495 -88.135 ;
      RECT 90.355 -86.809 90.445 -85.802 ;
      RECT 90.355 -86.285 90.495 -86.115 ;
      RECT 90.355 -85.388 90.445 -84.381 ;
      RECT 90.355 -85.075 90.495 -84.905 ;
      RECT 90.355 -83.579 90.445 -82.572 ;
      RECT 90.355 -83.055 90.495 -82.885 ;
      RECT 90.355 -82.158 90.445 -81.151 ;
      RECT 90.355 -81.845 90.495 -81.675 ;
      RECT 90.355 -80.349 90.445 -79.342 ;
      RECT 90.355 -79.825 90.495 -79.655 ;
      RECT 90.355 -78.928 90.445 -77.921 ;
      RECT 90.355 -78.615 90.495 -78.445 ;
      RECT 90.355 -77.119 90.445 -76.112 ;
      RECT 90.355 -76.595 90.495 -76.425 ;
      RECT 90.355 -75.698 90.445 -74.691 ;
      RECT 90.355 -75.385 90.495 -75.215 ;
      RECT 90.355 -73.889 90.445 -72.882 ;
      RECT 90.355 -73.365 90.495 -73.195 ;
      RECT 90.355 -72.468 90.445 -71.461 ;
      RECT 90.355 -72.155 90.495 -71.985 ;
      RECT 90.355 -70.659 90.445 -69.652 ;
      RECT 90.355 -70.135 90.495 -69.965 ;
      RECT 90.355 -69.238 90.445 -68.231 ;
      RECT 90.355 -68.925 90.495 -68.755 ;
      RECT 90.355 -67.429 90.445 -66.422 ;
      RECT 90.355 -66.905 90.495 -66.735 ;
      RECT 90.355 -66.008 90.445 -65.001 ;
      RECT 90.355 -65.695 90.495 -65.525 ;
      RECT 90.355 -64.199 90.445 -63.192 ;
      RECT 90.355 -63.675 90.495 -63.505 ;
      RECT 90.355 -62.778 90.445 -61.771 ;
      RECT 90.355 -62.465 90.495 -62.295 ;
      RECT 90.355 -60.969 90.445 -59.962 ;
      RECT 90.355 -60.445 90.495 -60.275 ;
      RECT 90.355 -59.548 90.445 -58.541 ;
      RECT 90.355 -59.235 90.495 -59.065 ;
      RECT 90.355 -57.739 90.445 -56.732 ;
      RECT 90.355 -57.215 90.495 -57.045 ;
      RECT 90.355 -56.318 90.445 -55.311 ;
      RECT 90.355 -56.005 90.495 -55.835 ;
      RECT 90.355 -54.509 90.445 -53.502 ;
      RECT 90.355 -53.985 90.495 -53.815 ;
      RECT 90.355 -53.088 90.445 -52.081 ;
      RECT 90.355 -52.775 90.495 -52.605 ;
      RECT 90.355 -51.279 90.445 -50.272 ;
      RECT 90.355 -50.755 90.495 -50.585 ;
      RECT 90.355 -49.858 90.445 -48.851 ;
      RECT 90.355 -49.545 90.495 -49.375 ;
      RECT 90.355 -48.049 90.445 -47.042 ;
      RECT 90.355 -47.525 90.495 -47.355 ;
      RECT 90.355 -46.628 90.445 -45.621 ;
      RECT 90.355 -46.315 90.495 -46.145 ;
      RECT 90.355 -44.819 90.445 -43.812 ;
      RECT 90.355 -44.295 90.495 -44.125 ;
      RECT 90.355 -43.398 90.445 -42.391 ;
      RECT 90.355 -43.085 90.495 -42.915 ;
      RECT 90.355 -41.589 90.445 -40.582 ;
      RECT 90.355 -41.065 90.495 -40.895 ;
      RECT 90.355 -40.168 90.445 -39.161 ;
      RECT 90.355 -39.855 90.495 -39.685 ;
      RECT 90.355 -38.359 90.445 -37.352 ;
      RECT 90.355 -37.835 90.495 -37.665 ;
      RECT 90.355 -36.938 90.445 -35.931 ;
      RECT 90.355 -36.625 90.495 -36.455 ;
      RECT 90.355 -35.129 90.445 -34.122 ;
      RECT 90.355 -34.605 90.495 -34.435 ;
      RECT 90.355 -33.708 90.445 -32.701 ;
      RECT 90.355 -33.395 90.495 -33.225 ;
      RECT 90.355 -31.899 90.445 -30.892 ;
      RECT 90.355 -31.375 90.495 -31.205 ;
      RECT 90.355 -30.478 90.445 -29.471 ;
      RECT 90.355 -30.165 90.495 -29.995 ;
      RECT 90.355 -28.669 90.445 -27.662 ;
      RECT 90.355 -28.145 90.495 -27.975 ;
      RECT 90.355 -27.248 90.445 -26.241 ;
      RECT 90.355 -26.935 90.495 -26.765 ;
      RECT 90.355 -25.439 90.445 -24.432 ;
      RECT 90.355 -24.915 90.495 -24.745 ;
      RECT 90.355 -24.018 90.445 -23.011 ;
      RECT 90.355 -23.705 90.495 -23.535 ;
      RECT 90.355 -22.209 90.445 -21.202 ;
      RECT 90.355 -21.685 90.495 -21.515 ;
      RECT 90.355 -20.788 90.445 -19.781 ;
      RECT 90.355 -20.475 90.495 -20.305 ;
      RECT 90.355 -18.979 90.445 -17.972 ;
      RECT 90.355 -18.455 90.495 -18.285 ;
      RECT 90.355 -17.558 90.445 -16.551 ;
      RECT 90.355 -17.245 90.495 -17.075 ;
      RECT 90.355 -15.749 90.445 -14.742 ;
      RECT 90.355 -15.225 90.495 -15.055 ;
      RECT 90.355 -14.328 90.445 -13.321 ;
      RECT 90.355 -14.015 90.495 -13.845 ;
      RECT 90.355 -12.519 90.445 -11.512 ;
      RECT 90.355 -11.995 90.495 -11.825 ;
      RECT 90.355 -11.098 90.445 -10.091 ;
      RECT 90.355 -10.785 90.495 -10.615 ;
      RECT 90.355 -9.289 90.445 -8.282 ;
      RECT 90.355 -8.765 90.495 -8.595 ;
      RECT 90.355 -7.868 90.445 -6.861 ;
      RECT 90.355 -7.555 90.495 -7.385 ;
      RECT 90.355 -6.059 90.445 -5.052 ;
      RECT 90.355 -5.535 90.495 -5.365 ;
      RECT 90.355 -4.638 90.445 -3.631 ;
      RECT 90.355 -4.325 90.495 -4.155 ;
      RECT 90.355 -2.829 90.445 -1.822 ;
      RECT 90.355 -2.305 90.495 -2.135 ;
      RECT 90.355 -1.408 90.445 -0.401 ;
      RECT 90.355 -1.095 90.495 -0.925 ;
      RECT 90.355 0.401 90.445 1.408 ;
      RECT 90.355 0.925 90.495 1.095 ;
      RECT 89.685 -111.495 89.855 -111.385 ;
      RECT 86.535 -111.495 89.855 -111.395 ;
      RECT 89.555 -101.538 89.645 -100.53 ;
      RECT 89.505 -100.935 89.645 -100.765 ;
      RECT 89.555 -99.73 89.645 -98.722 ;
      RECT 89.505 -99.495 89.645 -99.325 ;
      RECT 89.555 -98.308 89.645 -97.3 ;
      RECT 89.505 -97.705 89.645 -97.535 ;
      RECT 89.555 -96.5 89.645 -95.492 ;
      RECT 89.505 -96.265 89.645 -96.095 ;
      RECT 89.555 -95.078 89.645 -94.07 ;
      RECT 89.505 -94.475 89.645 -94.305 ;
      RECT 89.555 -93.27 89.645 -92.262 ;
      RECT 89.505 -93.035 89.645 -92.865 ;
      RECT 89.555 -91.848 89.645 -90.84 ;
      RECT 89.505 -91.245 89.645 -91.075 ;
      RECT 89.555 -90.04 89.645 -89.032 ;
      RECT 89.505 -89.805 89.645 -89.635 ;
      RECT 89.555 -88.618 89.645 -87.61 ;
      RECT 89.505 -88.015 89.645 -87.845 ;
      RECT 89.555 -86.81 89.645 -85.802 ;
      RECT 89.505 -86.575 89.645 -86.405 ;
      RECT 89.555 -85.388 89.645 -84.38 ;
      RECT 89.505 -84.785 89.645 -84.615 ;
      RECT 89.555 -83.58 89.645 -82.572 ;
      RECT 89.505 -83.345 89.645 -83.175 ;
      RECT 89.555 -82.158 89.645 -81.15 ;
      RECT 89.505 -81.555 89.645 -81.385 ;
      RECT 89.555 -80.35 89.645 -79.342 ;
      RECT 89.505 -80.115 89.645 -79.945 ;
      RECT 89.555 -78.928 89.645 -77.92 ;
      RECT 89.505 -78.325 89.645 -78.155 ;
      RECT 89.555 -77.12 89.645 -76.112 ;
      RECT 89.505 -76.885 89.645 -76.715 ;
      RECT 89.555 -75.698 89.645 -74.69 ;
      RECT 89.505 -75.095 89.645 -74.925 ;
      RECT 89.555 -73.89 89.645 -72.882 ;
      RECT 89.505 -73.655 89.645 -73.485 ;
      RECT 89.555 -72.468 89.645 -71.46 ;
      RECT 89.505 -71.865 89.645 -71.695 ;
      RECT 89.555 -70.66 89.645 -69.652 ;
      RECT 89.505 -70.425 89.645 -70.255 ;
      RECT 89.555 -69.238 89.645 -68.23 ;
      RECT 89.505 -68.635 89.645 -68.465 ;
      RECT 89.555 -67.43 89.645 -66.422 ;
      RECT 89.505 -67.195 89.645 -67.025 ;
      RECT 89.555 -66.008 89.645 -65 ;
      RECT 89.505 -65.405 89.645 -65.235 ;
      RECT 89.555 -64.2 89.645 -63.192 ;
      RECT 89.505 -63.965 89.645 -63.795 ;
      RECT 89.555 -62.778 89.645 -61.77 ;
      RECT 89.505 -62.175 89.645 -62.005 ;
      RECT 89.555 -60.97 89.645 -59.962 ;
      RECT 89.505 -60.735 89.645 -60.565 ;
      RECT 89.555 -59.548 89.645 -58.54 ;
      RECT 89.505 -58.945 89.645 -58.775 ;
      RECT 89.555 -57.74 89.645 -56.732 ;
      RECT 89.505 -57.505 89.645 -57.335 ;
      RECT 89.555 -56.318 89.645 -55.31 ;
      RECT 89.505 -55.715 89.645 -55.545 ;
      RECT 89.555 -54.51 89.645 -53.502 ;
      RECT 89.505 -54.275 89.645 -54.105 ;
      RECT 89.555 -53.088 89.645 -52.08 ;
      RECT 89.505 -52.485 89.645 -52.315 ;
      RECT 89.555 -51.28 89.645 -50.272 ;
      RECT 89.505 -51.045 89.645 -50.875 ;
      RECT 89.555 -49.858 89.645 -48.85 ;
      RECT 89.505 -49.255 89.645 -49.085 ;
      RECT 89.555 -48.05 89.645 -47.042 ;
      RECT 89.505 -47.815 89.645 -47.645 ;
      RECT 89.555 -46.628 89.645 -45.62 ;
      RECT 89.505 -46.025 89.645 -45.855 ;
      RECT 89.555 -44.82 89.645 -43.812 ;
      RECT 89.505 -44.585 89.645 -44.415 ;
      RECT 89.555 -43.398 89.645 -42.39 ;
      RECT 89.505 -42.795 89.645 -42.625 ;
      RECT 89.555 -41.59 89.645 -40.582 ;
      RECT 89.505 -41.355 89.645 -41.185 ;
      RECT 89.555 -40.168 89.645 -39.16 ;
      RECT 89.505 -39.565 89.645 -39.395 ;
      RECT 89.555 -38.36 89.645 -37.352 ;
      RECT 89.505 -38.125 89.645 -37.955 ;
      RECT 89.555 -36.938 89.645 -35.93 ;
      RECT 89.505 -36.335 89.645 -36.165 ;
      RECT 89.555 -35.13 89.645 -34.122 ;
      RECT 89.505 -34.895 89.645 -34.725 ;
      RECT 89.555 -33.708 89.645 -32.7 ;
      RECT 89.505 -33.105 89.645 -32.935 ;
      RECT 89.555 -31.9 89.645 -30.892 ;
      RECT 89.505 -31.665 89.645 -31.495 ;
      RECT 89.555 -30.478 89.645 -29.47 ;
      RECT 89.505 -29.875 89.645 -29.705 ;
      RECT 89.555 -28.67 89.645 -27.662 ;
      RECT 89.505 -28.435 89.645 -28.265 ;
      RECT 89.555 -27.248 89.645 -26.24 ;
      RECT 89.505 -26.645 89.645 -26.475 ;
      RECT 89.555 -25.44 89.645 -24.432 ;
      RECT 89.505 -25.205 89.645 -25.035 ;
      RECT 89.555 -24.018 89.645 -23.01 ;
      RECT 89.505 -23.415 89.645 -23.245 ;
      RECT 89.555 -22.21 89.645 -21.202 ;
      RECT 89.505 -21.975 89.645 -21.805 ;
      RECT 89.555 -20.788 89.645 -19.78 ;
      RECT 89.505 -20.185 89.645 -20.015 ;
      RECT 89.555 -18.98 89.645 -17.972 ;
      RECT 89.505 -18.745 89.645 -18.575 ;
      RECT 89.555 -17.558 89.645 -16.55 ;
      RECT 89.505 -16.955 89.645 -16.785 ;
      RECT 89.555 -15.75 89.645 -14.742 ;
      RECT 89.505 -15.515 89.645 -15.345 ;
      RECT 89.555 -14.328 89.645 -13.32 ;
      RECT 89.505 -13.725 89.645 -13.555 ;
      RECT 89.555 -12.52 89.645 -11.512 ;
      RECT 89.505 -12.285 89.645 -12.115 ;
      RECT 89.555 -11.098 89.645 -10.09 ;
      RECT 89.505 -10.495 89.645 -10.325 ;
      RECT 89.555 -9.29 89.645 -8.282 ;
      RECT 89.505 -9.055 89.645 -8.885 ;
      RECT 89.555 -7.868 89.645 -6.86 ;
      RECT 89.505 -7.265 89.645 -7.095 ;
      RECT 89.555 -6.06 89.645 -5.052 ;
      RECT 89.505 -5.825 89.645 -5.655 ;
      RECT 89.555 -4.638 89.645 -3.63 ;
      RECT 89.505 -4.035 89.645 -3.865 ;
      RECT 89.555 -2.83 89.645 -1.822 ;
      RECT 89.505 -2.595 89.645 -2.425 ;
      RECT 89.555 -1.408 89.645 -0.4 ;
      RECT 89.505 -0.805 89.645 -0.635 ;
      RECT 89.555 0.4 89.645 1.408 ;
      RECT 89.505 0.635 89.645 0.805 ;
      RECT 89.155 -101.538 89.245 -100.531 ;
      RECT 89.155 -101.225 89.295 -101.055 ;
      RECT 89.155 -99.729 89.245 -98.722 ;
      RECT 89.155 -99.205 89.295 -99.035 ;
      RECT 89.155 -98.308 89.245 -97.301 ;
      RECT 89.155 -97.995 89.295 -97.825 ;
      RECT 89.155 -96.499 89.245 -95.492 ;
      RECT 89.155 -95.975 89.295 -95.805 ;
      RECT 89.155 -95.078 89.245 -94.071 ;
      RECT 89.155 -94.765 89.295 -94.595 ;
      RECT 89.155 -93.269 89.245 -92.262 ;
      RECT 89.155 -92.745 89.295 -92.575 ;
      RECT 89.155 -91.848 89.245 -90.841 ;
      RECT 89.155 -91.535 89.295 -91.365 ;
      RECT 89.155 -90.039 89.245 -89.032 ;
      RECT 89.155 -89.515 89.295 -89.345 ;
      RECT 89.155 -88.618 89.245 -87.611 ;
      RECT 89.155 -88.305 89.295 -88.135 ;
      RECT 89.155 -86.809 89.245 -85.802 ;
      RECT 89.155 -86.285 89.295 -86.115 ;
      RECT 89.155 -85.388 89.245 -84.381 ;
      RECT 89.155 -85.075 89.295 -84.905 ;
      RECT 89.155 -83.579 89.245 -82.572 ;
      RECT 89.155 -83.055 89.295 -82.885 ;
      RECT 89.155 -82.158 89.245 -81.151 ;
      RECT 89.155 -81.845 89.295 -81.675 ;
      RECT 89.155 -80.349 89.245 -79.342 ;
      RECT 89.155 -79.825 89.295 -79.655 ;
      RECT 89.155 -78.928 89.245 -77.921 ;
      RECT 89.155 -78.615 89.295 -78.445 ;
      RECT 89.155 -77.119 89.245 -76.112 ;
      RECT 89.155 -76.595 89.295 -76.425 ;
      RECT 89.155 -75.698 89.245 -74.691 ;
      RECT 89.155 -75.385 89.295 -75.215 ;
      RECT 89.155 -73.889 89.245 -72.882 ;
      RECT 89.155 -73.365 89.295 -73.195 ;
      RECT 89.155 -72.468 89.245 -71.461 ;
      RECT 89.155 -72.155 89.295 -71.985 ;
      RECT 89.155 -70.659 89.245 -69.652 ;
      RECT 89.155 -70.135 89.295 -69.965 ;
      RECT 89.155 -69.238 89.245 -68.231 ;
      RECT 89.155 -68.925 89.295 -68.755 ;
      RECT 89.155 -67.429 89.245 -66.422 ;
      RECT 89.155 -66.905 89.295 -66.735 ;
      RECT 89.155 -66.008 89.245 -65.001 ;
      RECT 89.155 -65.695 89.295 -65.525 ;
      RECT 89.155 -64.199 89.245 -63.192 ;
      RECT 89.155 -63.675 89.295 -63.505 ;
      RECT 89.155 -62.778 89.245 -61.771 ;
      RECT 89.155 -62.465 89.295 -62.295 ;
      RECT 89.155 -60.969 89.245 -59.962 ;
      RECT 89.155 -60.445 89.295 -60.275 ;
      RECT 89.155 -59.548 89.245 -58.541 ;
      RECT 89.155 -59.235 89.295 -59.065 ;
      RECT 89.155 -57.739 89.245 -56.732 ;
      RECT 89.155 -57.215 89.295 -57.045 ;
      RECT 89.155 -56.318 89.245 -55.311 ;
      RECT 89.155 -56.005 89.295 -55.835 ;
      RECT 89.155 -54.509 89.245 -53.502 ;
      RECT 89.155 -53.985 89.295 -53.815 ;
      RECT 89.155 -53.088 89.245 -52.081 ;
      RECT 89.155 -52.775 89.295 -52.605 ;
      RECT 89.155 -51.279 89.245 -50.272 ;
      RECT 89.155 -50.755 89.295 -50.585 ;
      RECT 89.155 -49.858 89.245 -48.851 ;
      RECT 89.155 -49.545 89.295 -49.375 ;
      RECT 89.155 -48.049 89.245 -47.042 ;
      RECT 89.155 -47.525 89.295 -47.355 ;
      RECT 89.155 -46.628 89.245 -45.621 ;
      RECT 89.155 -46.315 89.295 -46.145 ;
      RECT 89.155 -44.819 89.245 -43.812 ;
      RECT 89.155 -44.295 89.295 -44.125 ;
      RECT 89.155 -43.398 89.245 -42.391 ;
      RECT 89.155 -43.085 89.295 -42.915 ;
      RECT 89.155 -41.589 89.245 -40.582 ;
      RECT 89.155 -41.065 89.295 -40.895 ;
      RECT 89.155 -40.168 89.245 -39.161 ;
      RECT 89.155 -39.855 89.295 -39.685 ;
      RECT 89.155 -38.359 89.245 -37.352 ;
      RECT 89.155 -37.835 89.295 -37.665 ;
      RECT 89.155 -36.938 89.245 -35.931 ;
      RECT 89.155 -36.625 89.295 -36.455 ;
      RECT 89.155 -35.129 89.245 -34.122 ;
      RECT 89.155 -34.605 89.295 -34.435 ;
      RECT 89.155 -33.708 89.245 -32.701 ;
      RECT 89.155 -33.395 89.295 -33.225 ;
      RECT 89.155 -31.899 89.245 -30.892 ;
      RECT 89.155 -31.375 89.295 -31.205 ;
      RECT 89.155 -30.478 89.245 -29.471 ;
      RECT 89.155 -30.165 89.295 -29.995 ;
      RECT 89.155 -28.669 89.245 -27.662 ;
      RECT 89.155 -28.145 89.295 -27.975 ;
      RECT 89.155 -27.248 89.245 -26.241 ;
      RECT 89.155 -26.935 89.295 -26.765 ;
      RECT 89.155 -25.439 89.245 -24.432 ;
      RECT 89.155 -24.915 89.295 -24.745 ;
      RECT 89.155 -24.018 89.245 -23.011 ;
      RECT 89.155 -23.705 89.295 -23.535 ;
      RECT 89.155 -22.209 89.245 -21.202 ;
      RECT 89.155 -21.685 89.295 -21.515 ;
      RECT 89.155 -20.788 89.245 -19.781 ;
      RECT 89.155 -20.475 89.295 -20.305 ;
      RECT 89.155 -18.979 89.245 -17.972 ;
      RECT 89.155 -18.455 89.295 -18.285 ;
      RECT 89.155 -17.558 89.245 -16.551 ;
      RECT 89.155 -17.245 89.295 -17.075 ;
      RECT 89.155 -15.749 89.245 -14.742 ;
      RECT 89.155 -15.225 89.295 -15.055 ;
      RECT 89.155 -14.328 89.245 -13.321 ;
      RECT 89.155 -14.015 89.295 -13.845 ;
      RECT 89.155 -12.519 89.245 -11.512 ;
      RECT 89.155 -11.995 89.295 -11.825 ;
      RECT 89.155 -11.098 89.245 -10.091 ;
      RECT 89.155 -10.785 89.295 -10.615 ;
      RECT 89.155 -9.289 89.245 -8.282 ;
      RECT 89.155 -8.765 89.295 -8.595 ;
      RECT 89.155 -7.868 89.245 -6.861 ;
      RECT 89.155 -7.555 89.295 -7.385 ;
      RECT 89.155 -6.059 89.245 -5.052 ;
      RECT 89.155 -5.535 89.295 -5.365 ;
      RECT 89.155 -4.638 89.245 -3.631 ;
      RECT 89.155 -4.325 89.295 -4.155 ;
      RECT 89.155 -2.829 89.245 -1.822 ;
      RECT 89.155 -2.305 89.295 -2.135 ;
      RECT 89.155 -1.408 89.245 -0.401 ;
      RECT 89.155 -1.095 89.295 -0.925 ;
      RECT 89.155 0.401 89.245 1.408 ;
      RECT 89.155 0.925 89.295 1.095 ;
      RECT 87.305 -111.685 88.785 -111.585 ;
      RECT 87.305 -112.055 87.405 -111.585 ;
      RECT 87.11 -114.395 88.685 -114.275 ;
      RECT 88.585 -114.895 88.685 -114.275 ;
      RECT 87.99 -114.895 88.09 -114.275 ;
      RECT 87.11 -114.85 87.21 -114.275 ;
      RECT 88.355 -101.538 88.445 -100.53 ;
      RECT 88.305 -100.935 88.445 -100.765 ;
      RECT 88.355 -99.73 88.445 -98.722 ;
      RECT 88.305 -99.495 88.445 -99.325 ;
      RECT 88.355 -98.308 88.445 -97.3 ;
      RECT 88.305 -97.705 88.445 -97.535 ;
      RECT 88.355 -96.5 88.445 -95.492 ;
      RECT 88.305 -96.265 88.445 -96.095 ;
      RECT 88.355 -95.078 88.445 -94.07 ;
      RECT 88.305 -94.475 88.445 -94.305 ;
      RECT 88.355 -93.27 88.445 -92.262 ;
      RECT 88.305 -93.035 88.445 -92.865 ;
      RECT 88.355 -91.848 88.445 -90.84 ;
      RECT 88.305 -91.245 88.445 -91.075 ;
      RECT 88.355 -90.04 88.445 -89.032 ;
      RECT 88.305 -89.805 88.445 -89.635 ;
      RECT 88.355 -88.618 88.445 -87.61 ;
      RECT 88.305 -88.015 88.445 -87.845 ;
      RECT 88.355 -86.81 88.445 -85.802 ;
      RECT 88.305 -86.575 88.445 -86.405 ;
      RECT 88.355 -85.388 88.445 -84.38 ;
      RECT 88.305 -84.785 88.445 -84.615 ;
      RECT 88.355 -83.58 88.445 -82.572 ;
      RECT 88.305 -83.345 88.445 -83.175 ;
      RECT 88.355 -82.158 88.445 -81.15 ;
      RECT 88.305 -81.555 88.445 -81.385 ;
      RECT 88.355 -80.35 88.445 -79.342 ;
      RECT 88.305 -80.115 88.445 -79.945 ;
      RECT 88.355 -78.928 88.445 -77.92 ;
      RECT 88.305 -78.325 88.445 -78.155 ;
      RECT 88.355 -77.12 88.445 -76.112 ;
      RECT 88.305 -76.885 88.445 -76.715 ;
      RECT 88.355 -75.698 88.445 -74.69 ;
      RECT 88.305 -75.095 88.445 -74.925 ;
      RECT 88.355 -73.89 88.445 -72.882 ;
      RECT 88.305 -73.655 88.445 -73.485 ;
      RECT 88.355 -72.468 88.445 -71.46 ;
      RECT 88.305 -71.865 88.445 -71.695 ;
      RECT 88.355 -70.66 88.445 -69.652 ;
      RECT 88.305 -70.425 88.445 -70.255 ;
      RECT 88.355 -69.238 88.445 -68.23 ;
      RECT 88.305 -68.635 88.445 -68.465 ;
      RECT 88.355 -67.43 88.445 -66.422 ;
      RECT 88.305 -67.195 88.445 -67.025 ;
      RECT 88.355 -66.008 88.445 -65 ;
      RECT 88.305 -65.405 88.445 -65.235 ;
      RECT 88.355 -64.2 88.445 -63.192 ;
      RECT 88.305 -63.965 88.445 -63.795 ;
      RECT 88.355 -62.778 88.445 -61.77 ;
      RECT 88.305 -62.175 88.445 -62.005 ;
      RECT 88.355 -60.97 88.445 -59.962 ;
      RECT 88.305 -60.735 88.445 -60.565 ;
      RECT 88.355 -59.548 88.445 -58.54 ;
      RECT 88.305 -58.945 88.445 -58.775 ;
      RECT 88.355 -57.74 88.445 -56.732 ;
      RECT 88.305 -57.505 88.445 -57.335 ;
      RECT 88.355 -56.318 88.445 -55.31 ;
      RECT 88.305 -55.715 88.445 -55.545 ;
      RECT 88.355 -54.51 88.445 -53.502 ;
      RECT 88.305 -54.275 88.445 -54.105 ;
      RECT 88.355 -53.088 88.445 -52.08 ;
      RECT 88.305 -52.485 88.445 -52.315 ;
      RECT 88.355 -51.28 88.445 -50.272 ;
      RECT 88.305 -51.045 88.445 -50.875 ;
      RECT 88.355 -49.858 88.445 -48.85 ;
      RECT 88.305 -49.255 88.445 -49.085 ;
      RECT 88.355 -48.05 88.445 -47.042 ;
      RECT 88.305 -47.815 88.445 -47.645 ;
      RECT 88.355 -46.628 88.445 -45.62 ;
      RECT 88.305 -46.025 88.445 -45.855 ;
      RECT 88.355 -44.82 88.445 -43.812 ;
      RECT 88.305 -44.585 88.445 -44.415 ;
      RECT 88.355 -43.398 88.445 -42.39 ;
      RECT 88.305 -42.795 88.445 -42.625 ;
      RECT 88.355 -41.59 88.445 -40.582 ;
      RECT 88.305 -41.355 88.445 -41.185 ;
      RECT 88.355 -40.168 88.445 -39.16 ;
      RECT 88.305 -39.565 88.445 -39.395 ;
      RECT 88.355 -38.36 88.445 -37.352 ;
      RECT 88.305 -38.125 88.445 -37.955 ;
      RECT 88.355 -36.938 88.445 -35.93 ;
      RECT 88.305 -36.335 88.445 -36.165 ;
      RECT 88.355 -35.13 88.445 -34.122 ;
      RECT 88.305 -34.895 88.445 -34.725 ;
      RECT 88.355 -33.708 88.445 -32.7 ;
      RECT 88.305 -33.105 88.445 -32.935 ;
      RECT 88.355 -31.9 88.445 -30.892 ;
      RECT 88.305 -31.665 88.445 -31.495 ;
      RECT 88.355 -30.478 88.445 -29.47 ;
      RECT 88.305 -29.875 88.445 -29.705 ;
      RECT 88.355 -28.67 88.445 -27.662 ;
      RECT 88.305 -28.435 88.445 -28.265 ;
      RECT 88.355 -27.248 88.445 -26.24 ;
      RECT 88.305 -26.645 88.445 -26.475 ;
      RECT 88.355 -25.44 88.445 -24.432 ;
      RECT 88.305 -25.205 88.445 -25.035 ;
      RECT 88.355 -24.018 88.445 -23.01 ;
      RECT 88.305 -23.415 88.445 -23.245 ;
      RECT 88.355 -22.21 88.445 -21.202 ;
      RECT 88.305 -21.975 88.445 -21.805 ;
      RECT 88.355 -20.788 88.445 -19.78 ;
      RECT 88.305 -20.185 88.445 -20.015 ;
      RECT 88.355 -18.98 88.445 -17.972 ;
      RECT 88.305 -18.745 88.445 -18.575 ;
      RECT 88.355 -17.558 88.445 -16.55 ;
      RECT 88.305 -16.955 88.445 -16.785 ;
      RECT 88.355 -15.75 88.445 -14.742 ;
      RECT 88.305 -15.515 88.445 -15.345 ;
      RECT 88.355 -14.328 88.445 -13.32 ;
      RECT 88.305 -13.725 88.445 -13.555 ;
      RECT 88.355 -12.52 88.445 -11.512 ;
      RECT 88.305 -12.285 88.445 -12.115 ;
      RECT 88.355 -11.098 88.445 -10.09 ;
      RECT 88.305 -10.495 88.445 -10.325 ;
      RECT 88.355 -9.29 88.445 -8.282 ;
      RECT 88.305 -9.055 88.445 -8.885 ;
      RECT 88.355 -7.868 88.445 -6.86 ;
      RECT 88.305 -7.265 88.445 -7.095 ;
      RECT 88.355 -6.06 88.445 -5.052 ;
      RECT 88.305 -5.825 88.445 -5.655 ;
      RECT 88.355 -4.638 88.445 -3.63 ;
      RECT 88.305 -4.035 88.445 -3.865 ;
      RECT 88.355 -2.83 88.445 -1.822 ;
      RECT 88.305 -2.595 88.445 -2.425 ;
      RECT 88.355 -1.408 88.445 -0.4 ;
      RECT 88.305 -0.805 88.445 -0.635 ;
      RECT 88.355 0.4 88.445 1.408 ;
      RECT 88.305 0.635 88.445 0.805 ;
      RECT 88.23 -114.685 88.405 -114.515 ;
      RECT 88.305 -114.895 88.405 -114.515 ;
      RECT 87.345 -113.555 87.445 -113.09 ;
      RECT 87.71 -113.555 87.81 -113.1 ;
      RECT 87.345 -113.555 88.19 -113.385 ;
      RECT 87.955 -101.538 88.045 -100.531 ;
      RECT 87.955 -101.225 88.095 -101.055 ;
      RECT 87.955 -99.729 88.045 -98.722 ;
      RECT 87.955 -99.205 88.095 -99.035 ;
      RECT 87.955 -98.308 88.045 -97.301 ;
      RECT 87.955 -97.995 88.095 -97.825 ;
      RECT 87.955 -96.499 88.045 -95.492 ;
      RECT 87.955 -95.975 88.095 -95.805 ;
      RECT 87.955 -95.078 88.045 -94.071 ;
      RECT 87.955 -94.765 88.095 -94.595 ;
      RECT 87.955 -93.269 88.045 -92.262 ;
      RECT 87.955 -92.745 88.095 -92.575 ;
      RECT 87.955 -91.848 88.045 -90.841 ;
      RECT 87.955 -91.535 88.095 -91.365 ;
      RECT 87.955 -90.039 88.045 -89.032 ;
      RECT 87.955 -89.515 88.095 -89.345 ;
      RECT 87.955 -88.618 88.045 -87.611 ;
      RECT 87.955 -88.305 88.095 -88.135 ;
      RECT 87.955 -86.809 88.045 -85.802 ;
      RECT 87.955 -86.285 88.095 -86.115 ;
      RECT 87.955 -85.388 88.045 -84.381 ;
      RECT 87.955 -85.075 88.095 -84.905 ;
      RECT 87.955 -83.579 88.045 -82.572 ;
      RECT 87.955 -83.055 88.095 -82.885 ;
      RECT 87.955 -82.158 88.045 -81.151 ;
      RECT 87.955 -81.845 88.095 -81.675 ;
      RECT 87.955 -80.349 88.045 -79.342 ;
      RECT 87.955 -79.825 88.095 -79.655 ;
      RECT 87.955 -78.928 88.045 -77.921 ;
      RECT 87.955 -78.615 88.095 -78.445 ;
      RECT 87.955 -77.119 88.045 -76.112 ;
      RECT 87.955 -76.595 88.095 -76.425 ;
      RECT 87.955 -75.698 88.045 -74.691 ;
      RECT 87.955 -75.385 88.095 -75.215 ;
      RECT 87.955 -73.889 88.045 -72.882 ;
      RECT 87.955 -73.365 88.095 -73.195 ;
      RECT 87.955 -72.468 88.045 -71.461 ;
      RECT 87.955 -72.155 88.095 -71.985 ;
      RECT 87.955 -70.659 88.045 -69.652 ;
      RECT 87.955 -70.135 88.095 -69.965 ;
      RECT 87.955 -69.238 88.045 -68.231 ;
      RECT 87.955 -68.925 88.095 -68.755 ;
      RECT 87.955 -67.429 88.045 -66.422 ;
      RECT 87.955 -66.905 88.095 -66.735 ;
      RECT 87.955 -66.008 88.045 -65.001 ;
      RECT 87.955 -65.695 88.095 -65.525 ;
      RECT 87.955 -64.199 88.045 -63.192 ;
      RECT 87.955 -63.675 88.095 -63.505 ;
      RECT 87.955 -62.778 88.045 -61.771 ;
      RECT 87.955 -62.465 88.095 -62.295 ;
      RECT 87.955 -60.969 88.045 -59.962 ;
      RECT 87.955 -60.445 88.095 -60.275 ;
      RECT 87.955 -59.548 88.045 -58.541 ;
      RECT 87.955 -59.235 88.095 -59.065 ;
      RECT 87.955 -57.739 88.045 -56.732 ;
      RECT 87.955 -57.215 88.095 -57.045 ;
      RECT 87.955 -56.318 88.045 -55.311 ;
      RECT 87.955 -56.005 88.095 -55.835 ;
      RECT 87.955 -54.509 88.045 -53.502 ;
      RECT 87.955 -53.985 88.095 -53.815 ;
      RECT 87.955 -53.088 88.045 -52.081 ;
      RECT 87.955 -52.775 88.095 -52.605 ;
      RECT 87.955 -51.279 88.045 -50.272 ;
      RECT 87.955 -50.755 88.095 -50.585 ;
      RECT 87.955 -49.858 88.045 -48.851 ;
      RECT 87.955 -49.545 88.095 -49.375 ;
      RECT 87.955 -48.049 88.045 -47.042 ;
      RECT 87.955 -47.525 88.095 -47.355 ;
      RECT 87.955 -46.628 88.045 -45.621 ;
      RECT 87.955 -46.315 88.095 -46.145 ;
      RECT 87.955 -44.819 88.045 -43.812 ;
      RECT 87.955 -44.295 88.095 -44.125 ;
      RECT 87.955 -43.398 88.045 -42.391 ;
      RECT 87.955 -43.085 88.095 -42.915 ;
      RECT 87.955 -41.589 88.045 -40.582 ;
      RECT 87.955 -41.065 88.095 -40.895 ;
      RECT 87.955 -40.168 88.045 -39.161 ;
      RECT 87.955 -39.855 88.095 -39.685 ;
      RECT 87.955 -38.359 88.045 -37.352 ;
      RECT 87.955 -37.835 88.095 -37.665 ;
      RECT 87.955 -36.938 88.045 -35.931 ;
      RECT 87.955 -36.625 88.095 -36.455 ;
      RECT 87.955 -35.129 88.045 -34.122 ;
      RECT 87.955 -34.605 88.095 -34.435 ;
      RECT 87.955 -33.708 88.045 -32.701 ;
      RECT 87.955 -33.395 88.095 -33.225 ;
      RECT 87.955 -31.899 88.045 -30.892 ;
      RECT 87.955 -31.375 88.095 -31.205 ;
      RECT 87.955 -30.478 88.045 -29.471 ;
      RECT 87.955 -30.165 88.095 -29.995 ;
      RECT 87.955 -28.669 88.045 -27.662 ;
      RECT 87.955 -28.145 88.095 -27.975 ;
      RECT 87.955 -27.248 88.045 -26.241 ;
      RECT 87.955 -26.935 88.095 -26.765 ;
      RECT 87.955 -25.439 88.045 -24.432 ;
      RECT 87.955 -24.915 88.095 -24.745 ;
      RECT 87.955 -24.018 88.045 -23.011 ;
      RECT 87.955 -23.705 88.095 -23.535 ;
      RECT 87.955 -22.209 88.045 -21.202 ;
      RECT 87.955 -21.685 88.095 -21.515 ;
      RECT 87.955 -20.788 88.045 -19.781 ;
      RECT 87.955 -20.475 88.095 -20.305 ;
      RECT 87.955 -18.979 88.045 -17.972 ;
      RECT 87.955 -18.455 88.095 -18.285 ;
      RECT 87.955 -17.558 88.045 -16.551 ;
      RECT 87.955 -17.245 88.095 -17.075 ;
      RECT 87.955 -15.749 88.045 -14.742 ;
      RECT 87.955 -15.225 88.095 -15.055 ;
      RECT 87.955 -14.328 88.045 -13.321 ;
      RECT 87.955 -14.015 88.095 -13.845 ;
      RECT 87.955 -12.519 88.045 -11.512 ;
      RECT 87.955 -11.995 88.095 -11.825 ;
      RECT 87.955 -11.098 88.045 -10.091 ;
      RECT 87.955 -10.785 88.095 -10.615 ;
      RECT 87.955 -9.289 88.045 -8.282 ;
      RECT 87.955 -8.765 88.095 -8.595 ;
      RECT 87.955 -7.868 88.045 -6.861 ;
      RECT 87.955 -7.555 88.095 -7.385 ;
      RECT 87.955 -6.059 88.045 -5.052 ;
      RECT 87.955 -5.535 88.095 -5.365 ;
      RECT 87.955 -4.638 88.045 -3.631 ;
      RECT 87.955 -4.325 88.095 -4.155 ;
      RECT 87.955 -2.829 88.045 -1.822 ;
      RECT 87.955 -2.305 88.095 -2.135 ;
      RECT 87.955 -1.408 88.045 -0.401 ;
      RECT 87.955 -1.095 88.095 -0.925 ;
      RECT 87.955 0.401 88.045 1.408 ;
      RECT 87.955 0.925 88.095 1.095 ;
      RECT 87.64 -114.685 87.81 -114.515 ;
      RECT 87.71 -114.895 87.81 -114.515 ;
      RECT 87.155 -101.538 87.245 -100.53 ;
      RECT 87.105 -100.935 87.245 -100.765 ;
      RECT 87.155 -99.73 87.245 -98.722 ;
      RECT 87.105 -99.495 87.245 -99.325 ;
      RECT 87.155 -98.308 87.245 -97.3 ;
      RECT 87.105 -97.705 87.245 -97.535 ;
      RECT 87.155 -96.5 87.245 -95.492 ;
      RECT 87.105 -96.265 87.245 -96.095 ;
      RECT 87.155 -95.078 87.245 -94.07 ;
      RECT 87.105 -94.475 87.245 -94.305 ;
      RECT 87.155 -93.27 87.245 -92.262 ;
      RECT 87.105 -93.035 87.245 -92.865 ;
      RECT 87.155 -91.848 87.245 -90.84 ;
      RECT 87.105 -91.245 87.245 -91.075 ;
      RECT 87.155 -90.04 87.245 -89.032 ;
      RECT 87.105 -89.805 87.245 -89.635 ;
      RECT 87.155 -88.618 87.245 -87.61 ;
      RECT 87.105 -88.015 87.245 -87.845 ;
      RECT 87.155 -86.81 87.245 -85.802 ;
      RECT 87.105 -86.575 87.245 -86.405 ;
      RECT 87.155 -85.388 87.245 -84.38 ;
      RECT 87.105 -84.785 87.245 -84.615 ;
      RECT 87.155 -83.58 87.245 -82.572 ;
      RECT 87.105 -83.345 87.245 -83.175 ;
      RECT 87.155 -82.158 87.245 -81.15 ;
      RECT 87.105 -81.555 87.245 -81.385 ;
      RECT 87.155 -80.35 87.245 -79.342 ;
      RECT 87.105 -80.115 87.245 -79.945 ;
      RECT 87.155 -78.928 87.245 -77.92 ;
      RECT 87.105 -78.325 87.245 -78.155 ;
      RECT 87.155 -77.12 87.245 -76.112 ;
      RECT 87.105 -76.885 87.245 -76.715 ;
      RECT 87.155 -75.698 87.245 -74.69 ;
      RECT 87.105 -75.095 87.245 -74.925 ;
      RECT 87.155 -73.89 87.245 -72.882 ;
      RECT 87.105 -73.655 87.245 -73.485 ;
      RECT 87.155 -72.468 87.245 -71.46 ;
      RECT 87.105 -71.865 87.245 -71.695 ;
      RECT 87.155 -70.66 87.245 -69.652 ;
      RECT 87.105 -70.425 87.245 -70.255 ;
      RECT 87.155 -69.238 87.245 -68.23 ;
      RECT 87.105 -68.635 87.245 -68.465 ;
      RECT 87.155 -67.43 87.245 -66.422 ;
      RECT 87.105 -67.195 87.245 -67.025 ;
      RECT 87.155 -66.008 87.245 -65 ;
      RECT 87.105 -65.405 87.245 -65.235 ;
      RECT 87.155 -64.2 87.245 -63.192 ;
      RECT 87.105 -63.965 87.245 -63.795 ;
      RECT 87.155 -62.778 87.245 -61.77 ;
      RECT 87.105 -62.175 87.245 -62.005 ;
      RECT 87.155 -60.97 87.245 -59.962 ;
      RECT 87.105 -60.735 87.245 -60.565 ;
      RECT 87.155 -59.548 87.245 -58.54 ;
      RECT 87.105 -58.945 87.245 -58.775 ;
      RECT 87.155 -57.74 87.245 -56.732 ;
      RECT 87.105 -57.505 87.245 -57.335 ;
      RECT 87.155 -56.318 87.245 -55.31 ;
      RECT 87.105 -55.715 87.245 -55.545 ;
      RECT 87.155 -54.51 87.245 -53.502 ;
      RECT 87.105 -54.275 87.245 -54.105 ;
      RECT 87.155 -53.088 87.245 -52.08 ;
      RECT 87.105 -52.485 87.245 -52.315 ;
      RECT 87.155 -51.28 87.245 -50.272 ;
      RECT 87.105 -51.045 87.245 -50.875 ;
      RECT 87.155 -49.858 87.245 -48.85 ;
      RECT 87.105 -49.255 87.245 -49.085 ;
      RECT 87.155 -48.05 87.245 -47.042 ;
      RECT 87.105 -47.815 87.245 -47.645 ;
      RECT 87.155 -46.628 87.245 -45.62 ;
      RECT 87.105 -46.025 87.245 -45.855 ;
      RECT 87.155 -44.82 87.245 -43.812 ;
      RECT 87.105 -44.585 87.245 -44.415 ;
      RECT 87.155 -43.398 87.245 -42.39 ;
      RECT 87.105 -42.795 87.245 -42.625 ;
      RECT 87.155 -41.59 87.245 -40.582 ;
      RECT 87.105 -41.355 87.245 -41.185 ;
      RECT 87.155 -40.168 87.245 -39.16 ;
      RECT 87.105 -39.565 87.245 -39.395 ;
      RECT 87.155 -38.36 87.245 -37.352 ;
      RECT 87.105 -38.125 87.245 -37.955 ;
      RECT 87.155 -36.938 87.245 -35.93 ;
      RECT 87.105 -36.335 87.245 -36.165 ;
      RECT 87.155 -35.13 87.245 -34.122 ;
      RECT 87.105 -34.895 87.245 -34.725 ;
      RECT 87.155 -33.708 87.245 -32.7 ;
      RECT 87.105 -33.105 87.245 -32.935 ;
      RECT 87.155 -31.9 87.245 -30.892 ;
      RECT 87.105 -31.665 87.245 -31.495 ;
      RECT 87.155 -30.478 87.245 -29.47 ;
      RECT 87.105 -29.875 87.245 -29.705 ;
      RECT 87.155 -28.67 87.245 -27.662 ;
      RECT 87.105 -28.435 87.245 -28.265 ;
      RECT 87.155 -27.248 87.245 -26.24 ;
      RECT 87.105 -26.645 87.245 -26.475 ;
      RECT 87.155 -25.44 87.245 -24.432 ;
      RECT 87.105 -25.205 87.245 -25.035 ;
      RECT 87.155 -24.018 87.245 -23.01 ;
      RECT 87.105 -23.415 87.245 -23.245 ;
      RECT 87.155 -22.21 87.245 -21.202 ;
      RECT 87.105 -21.975 87.245 -21.805 ;
      RECT 87.155 -20.788 87.245 -19.78 ;
      RECT 87.105 -20.185 87.245 -20.015 ;
      RECT 87.155 -18.98 87.245 -17.972 ;
      RECT 87.105 -18.745 87.245 -18.575 ;
      RECT 87.155 -17.558 87.245 -16.55 ;
      RECT 87.105 -16.955 87.245 -16.785 ;
      RECT 87.155 -15.75 87.245 -14.742 ;
      RECT 87.105 -15.515 87.245 -15.345 ;
      RECT 87.155 -14.328 87.245 -13.32 ;
      RECT 87.105 -13.725 87.245 -13.555 ;
      RECT 87.155 -12.52 87.245 -11.512 ;
      RECT 87.105 -12.285 87.245 -12.115 ;
      RECT 87.155 -11.098 87.245 -10.09 ;
      RECT 87.105 -10.495 87.245 -10.325 ;
      RECT 87.155 -9.29 87.245 -8.282 ;
      RECT 87.105 -9.055 87.245 -8.885 ;
      RECT 87.155 -7.868 87.245 -6.86 ;
      RECT 87.105 -7.265 87.245 -7.095 ;
      RECT 87.155 -6.06 87.245 -5.052 ;
      RECT 87.105 -5.825 87.245 -5.655 ;
      RECT 87.155 -4.638 87.245 -3.63 ;
      RECT 87.105 -4.035 87.245 -3.865 ;
      RECT 87.155 -2.83 87.245 -1.822 ;
      RECT 87.105 -2.595 87.245 -2.425 ;
      RECT 87.155 -1.408 87.245 -0.4 ;
      RECT 87.105 -0.805 87.245 -0.635 ;
      RECT 87.155 0.4 87.245 1.408 ;
      RECT 87.105 0.635 87.245 0.805 ;
      RECT 86.755 -101.538 86.845 -100.531 ;
      RECT 86.755 -101.225 86.895 -101.055 ;
      RECT 86.755 -99.729 86.845 -98.722 ;
      RECT 86.755 -99.205 86.895 -99.035 ;
      RECT 86.755 -98.308 86.845 -97.301 ;
      RECT 86.755 -97.995 86.895 -97.825 ;
      RECT 86.755 -96.499 86.845 -95.492 ;
      RECT 86.755 -95.975 86.895 -95.805 ;
      RECT 86.755 -95.078 86.845 -94.071 ;
      RECT 86.755 -94.765 86.895 -94.595 ;
      RECT 86.755 -93.269 86.845 -92.262 ;
      RECT 86.755 -92.745 86.895 -92.575 ;
      RECT 86.755 -91.848 86.845 -90.841 ;
      RECT 86.755 -91.535 86.895 -91.365 ;
      RECT 86.755 -90.039 86.845 -89.032 ;
      RECT 86.755 -89.515 86.895 -89.345 ;
      RECT 86.755 -88.618 86.845 -87.611 ;
      RECT 86.755 -88.305 86.895 -88.135 ;
      RECT 86.755 -86.809 86.845 -85.802 ;
      RECT 86.755 -86.285 86.895 -86.115 ;
      RECT 86.755 -85.388 86.845 -84.381 ;
      RECT 86.755 -85.075 86.895 -84.905 ;
      RECT 86.755 -83.579 86.845 -82.572 ;
      RECT 86.755 -83.055 86.895 -82.885 ;
      RECT 86.755 -82.158 86.845 -81.151 ;
      RECT 86.755 -81.845 86.895 -81.675 ;
      RECT 86.755 -80.349 86.845 -79.342 ;
      RECT 86.755 -79.825 86.895 -79.655 ;
      RECT 86.755 -78.928 86.845 -77.921 ;
      RECT 86.755 -78.615 86.895 -78.445 ;
      RECT 86.755 -77.119 86.845 -76.112 ;
      RECT 86.755 -76.595 86.895 -76.425 ;
      RECT 86.755 -75.698 86.845 -74.691 ;
      RECT 86.755 -75.385 86.895 -75.215 ;
      RECT 86.755 -73.889 86.845 -72.882 ;
      RECT 86.755 -73.365 86.895 -73.195 ;
      RECT 86.755 -72.468 86.845 -71.461 ;
      RECT 86.755 -72.155 86.895 -71.985 ;
      RECT 86.755 -70.659 86.845 -69.652 ;
      RECT 86.755 -70.135 86.895 -69.965 ;
      RECT 86.755 -69.238 86.845 -68.231 ;
      RECT 86.755 -68.925 86.895 -68.755 ;
      RECT 86.755 -67.429 86.845 -66.422 ;
      RECT 86.755 -66.905 86.895 -66.735 ;
      RECT 86.755 -66.008 86.845 -65.001 ;
      RECT 86.755 -65.695 86.895 -65.525 ;
      RECT 86.755 -64.199 86.845 -63.192 ;
      RECT 86.755 -63.675 86.895 -63.505 ;
      RECT 86.755 -62.778 86.845 -61.771 ;
      RECT 86.755 -62.465 86.895 -62.295 ;
      RECT 86.755 -60.969 86.845 -59.962 ;
      RECT 86.755 -60.445 86.895 -60.275 ;
      RECT 86.755 -59.548 86.845 -58.541 ;
      RECT 86.755 -59.235 86.895 -59.065 ;
      RECT 86.755 -57.739 86.845 -56.732 ;
      RECT 86.755 -57.215 86.895 -57.045 ;
      RECT 86.755 -56.318 86.845 -55.311 ;
      RECT 86.755 -56.005 86.895 -55.835 ;
      RECT 86.755 -54.509 86.845 -53.502 ;
      RECT 86.755 -53.985 86.895 -53.815 ;
      RECT 86.755 -53.088 86.845 -52.081 ;
      RECT 86.755 -52.775 86.895 -52.605 ;
      RECT 86.755 -51.279 86.845 -50.272 ;
      RECT 86.755 -50.755 86.895 -50.585 ;
      RECT 86.755 -49.858 86.845 -48.851 ;
      RECT 86.755 -49.545 86.895 -49.375 ;
      RECT 86.755 -48.049 86.845 -47.042 ;
      RECT 86.755 -47.525 86.895 -47.355 ;
      RECT 86.755 -46.628 86.845 -45.621 ;
      RECT 86.755 -46.315 86.895 -46.145 ;
      RECT 86.755 -44.819 86.845 -43.812 ;
      RECT 86.755 -44.295 86.895 -44.125 ;
      RECT 86.755 -43.398 86.845 -42.391 ;
      RECT 86.755 -43.085 86.895 -42.915 ;
      RECT 86.755 -41.589 86.845 -40.582 ;
      RECT 86.755 -41.065 86.895 -40.895 ;
      RECT 86.755 -40.168 86.845 -39.161 ;
      RECT 86.755 -39.855 86.895 -39.685 ;
      RECT 86.755 -38.359 86.845 -37.352 ;
      RECT 86.755 -37.835 86.895 -37.665 ;
      RECT 86.755 -36.938 86.845 -35.931 ;
      RECT 86.755 -36.625 86.895 -36.455 ;
      RECT 86.755 -35.129 86.845 -34.122 ;
      RECT 86.755 -34.605 86.895 -34.435 ;
      RECT 86.755 -33.708 86.845 -32.701 ;
      RECT 86.755 -33.395 86.895 -33.225 ;
      RECT 86.755 -31.899 86.845 -30.892 ;
      RECT 86.755 -31.375 86.895 -31.205 ;
      RECT 86.755 -30.478 86.845 -29.471 ;
      RECT 86.755 -30.165 86.895 -29.995 ;
      RECT 86.755 -28.669 86.845 -27.662 ;
      RECT 86.755 -28.145 86.895 -27.975 ;
      RECT 86.755 -27.248 86.845 -26.241 ;
      RECT 86.755 -26.935 86.895 -26.765 ;
      RECT 86.755 -25.439 86.845 -24.432 ;
      RECT 86.755 -24.915 86.895 -24.745 ;
      RECT 86.755 -24.018 86.845 -23.011 ;
      RECT 86.755 -23.705 86.895 -23.535 ;
      RECT 86.755 -22.209 86.845 -21.202 ;
      RECT 86.755 -21.685 86.895 -21.515 ;
      RECT 86.755 -20.788 86.845 -19.781 ;
      RECT 86.755 -20.475 86.895 -20.305 ;
      RECT 86.755 -18.979 86.845 -17.972 ;
      RECT 86.755 -18.455 86.895 -18.285 ;
      RECT 86.755 -17.558 86.845 -16.551 ;
      RECT 86.755 -17.245 86.895 -17.075 ;
      RECT 86.755 -15.749 86.845 -14.742 ;
      RECT 86.755 -15.225 86.895 -15.055 ;
      RECT 86.755 -14.328 86.845 -13.321 ;
      RECT 86.755 -14.015 86.895 -13.845 ;
      RECT 86.755 -12.519 86.845 -11.512 ;
      RECT 86.755 -11.995 86.895 -11.825 ;
      RECT 86.755 -11.098 86.845 -10.091 ;
      RECT 86.755 -10.785 86.895 -10.615 ;
      RECT 86.755 -9.289 86.845 -8.282 ;
      RECT 86.755 -8.765 86.895 -8.595 ;
      RECT 86.755 -7.868 86.845 -6.861 ;
      RECT 86.755 -7.555 86.895 -7.385 ;
      RECT 86.755 -6.059 86.845 -5.052 ;
      RECT 86.755 -5.535 86.895 -5.365 ;
      RECT 86.755 -4.638 86.845 -3.631 ;
      RECT 86.755 -4.325 86.895 -4.155 ;
      RECT 86.755 -2.829 86.845 -1.822 ;
      RECT 86.755 -2.305 86.895 -2.135 ;
      RECT 86.755 -1.408 86.845 -0.401 ;
      RECT 86.755 -1.095 86.895 -0.925 ;
      RECT 86.755 0.401 86.845 1.408 ;
      RECT 86.755 0.925 86.895 1.095 ;
      RECT 82.585 -108.935 86.365 -108.815 ;
      RECT 83.905 -109.475 84.005 -108.815 ;
      RECT 83.345 -109.475 83.445 -108.815 ;
      RECT 82.785 -109.475 82.885 -108.815 ;
      RECT 85.955 -101.538 86.045 -100.53 ;
      RECT 85.905 -100.935 86.045 -100.765 ;
      RECT 85.955 -99.73 86.045 -98.722 ;
      RECT 85.905 -99.495 86.045 -99.325 ;
      RECT 85.955 -98.308 86.045 -97.3 ;
      RECT 85.905 -97.705 86.045 -97.535 ;
      RECT 85.955 -96.5 86.045 -95.492 ;
      RECT 85.905 -96.265 86.045 -96.095 ;
      RECT 85.955 -95.078 86.045 -94.07 ;
      RECT 85.905 -94.475 86.045 -94.305 ;
      RECT 85.955 -93.27 86.045 -92.262 ;
      RECT 85.905 -93.035 86.045 -92.865 ;
      RECT 85.955 -91.848 86.045 -90.84 ;
      RECT 85.905 -91.245 86.045 -91.075 ;
      RECT 85.955 -90.04 86.045 -89.032 ;
      RECT 85.905 -89.805 86.045 -89.635 ;
      RECT 85.955 -88.618 86.045 -87.61 ;
      RECT 85.905 -88.015 86.045 -87.845 ;
      RECT 85.955 -86.81 86.045 -85.802 ;
      RECT 85.905 -86.575 86.045 -86.405 ;
      RECT 85.955 -85.388 86.045 -84.38 ;
      RECT 85.905 -84.785 86.045 -84.615 ;
      RECT 85.955 -83.58 86.045 -82.572 ;
      RECT 85.905 -83.345 86.045 -83.175 ;
      RECT 85.955 -82.158 86.045 -81.15 ;
      RECT 85.905 -81.555 86.045 -81.385 ;
      RECT 85.955 -80.35 86.045 -79.342 ;
      RECT 85.905 -80.115 86.045 -79.945 ;
      RECT 85.955 -78.928 86.045 -77.92 ;
      RECT 85.905 -78.325 86.045 -78.155 ;
      RECT 85.955 -77.12 86.045 -76.112 ;
      RECT 85.905 -76.885 86.045 -76.715 ;
      RECT 85.955 -75.698 86.045 -74.69 ;
      RECT 85.905 -75.095 86.045 -74.925 ;
      RECT 85.955 -73.89 86.045 -72.882 ;
      RECT 85.905 -73.655 86.045 -73.485 ;
      RECT 85.955 -72.468 86.045 -71.46 ;
      RECT 85.905 -71.865 86.045 -71.695 ;
      RECT 85.955 -70.66 86.045 -69.652 ;
      RECT 85.905 -70.425 86.045 -70.255 ;
      RECT 85.955 -69.238 86.045 -68.23 ;
      RECT 85.905 -68.635 86.045 -68.465 ;
      RECT 85.955 -67.43 86.045 -66.422 ;
      RECT 85.905 -67.195 86.045 -67.025 ;
      RECT 85.955 -66.008 86.045 -65 ;
      RECT 85.905 -65.405 86.045 -65.235 ;
      RECT 85.955 -64.2 86.045 -63.192 ;
      RECT 85.905 -63.965 86.045 -63.795 ;
      RECT 85.955 -62.778 86.045 -61.77 ;
      RECT 85.905 -62.175 86.045 -62.005 ;
      RECT 85.955 -60.97 86.045 -59.962 ;
      RECT 85.905 -60.735 86.045 -60.565 ;
      RECT 85.955 -59.548 86.045 -58.54 ;
      RECT 85.905 -58.945 86.045 -58.775 ;
      RECT 85.955 -57.74 86.045 -56.732 ;
      RECT 85.905 -57.505 86.045 -57.335 ;
      RECT 85.955 -56.318 86.045 -55.31 ;
      RECT 85.905 -55.715 86.045 -55.545 ;
      RECT 85.955 -54.51 86.045 -53.502 ;
      RECT 85.905 -54.275 86.045 -54.105 ;
      RECT 85.955 -53.088 86.045 -52.08 ;
      RECT 85.905 -52.485 86.045 -52.315 ;
      RECT 85.955 -51.28 86.045 -50.272 ;
      RECT 85.905 -51.045 86.045 -50.875 ;
      RECT 85.955 -49.858 86.045 -48.85 ;
      RECT 85.905 -49.255 86.045 -49.085 ;
      RECT 85.955 -48.05 86.045 -47.042 ;
      RECT 85.905 -47.815 86.045 -47.645 ;
      RECT 85.955 -46.628 86.045 -45.62 ;
      RECT 85.905 -46.025 86.045 -45.855 ;
      RECT 85.955 -44.82 86.045 -43.812 ;
      RECT 85.905 -44.585 86.045 -44.415 ;
      RECT 85.955 -43.398 86.045 -42.39 ;
      RECT 85.905 -42.795 86.045 -42.625 ;
      RECT 85.955 -41.59 86.045 -40.582 ;
      RECT 85.905 -41.355 86.045 -41.185 ;
      RECT 85.955 -40.168 86.045 -39.16 ;
      RECT 85.905 -39.565 86.045 -39.395 ;
      RECT 85.955 -38.36 86.045 -37.352 ;
      RECT 85.905 -38.125 86.045 -37.955 ;
      RECT 85.955 -36.938 86.045 -35.93 ;
      RECT 85.905 -36.335 86.045 -36.165 ;
      RECT 85.955 -35.13 86.045 -34.122 ;
      RECT 85.905 -34.895 86.045 -34.725 ;
      RECT 85.955 -33.708 86.045 -32.7 ;
      RECT 85.905 -33.105 86.045 -32.935 ;
      RECT 85.955 -31.9 86.045 -30.892 ;
      RECT 85.905 -31.665 86.045 -31.495 ;
      RECT 85.955 -30.478 86.045 -29.47 ;
      RECT 85.905 -29.875 86.045 -29.705 ;
      RECT 85.955 -28.67 86.045 -27.662 ;
      RECT 85.905 -28.435 86.045 -28.265 ;
      RECT 85.955 -27.248 86.045 -26.24 ;
      RECT 85.905 -26.645 86.045 -26.475 ;
      RECT 85.955 -25.44 86.045 -24.432 ;
      RECT 85.905 -25.205 86.045 -25.035 ;
      RECT 85.955 -24.018 86.045 -23.01 ;
      RECT 85.905 -23.415 86.045 -23.245 ;
      RECT 85.955 -22.21 86.045 -21.202 ;
      RECT 85.905 -21.975 86.045 -21.805 ;
      RECT 85.955 -20.788 86.045 -19.78 ;
      RECT 85.905 -20.185 86.045 -20.015 ;
      RECT 85.955 -18.98 86.045 -17.972 ;
      RECT 85.905 -18.745 86.045 -18.575 ;
      RECT 85.955 -17.558 86.045 -16.55 ;
      RECT 85.905 -16.955 86.045 -16.785 ;
      RECT 85.955 -15.75 86.045 -14.742 ;
      RECT 85.905 -15.515 86.045 -15.345 ;
      RECT 85.955 -14.328 86.045 -13.32 ;
      RECT 85.905 -13.725 86.045 -13.555 ;
      RECT 85.955 -12.52 86.045 -11.512 ;
      RECT 85.905 -12.285 86.045 -12.115 ;
      RECT 85.955 -11.098 86.045 -10.09 ;
      RECT 85.905 -10.495 86.045 -10.325 ;
      RECT 85.955 -9.29 86.045 -8.282 ;
      RECT 85.905 -9.055 86.045 -8.885 ;
      RECT 85.955 -7.868 86.045 -6.86 ;
      RECT 85.905 -7.265 86.045 -7.095 ;
      RECT 85.955 -6.06 86.045 -5.052 ;
      RECT 85.905 -5.825 86.045 -5.655 ;
      RECT 85.955 -4.638 86.045 -3.63 ;
      RECT 85.905 -4.035 86.045 -3.865 ;
      RECT 85.955 -2.83 86.045 -1.822 ;
      RECT 85.905 -2.595 86.045 -2.425 ;
      RECT 85.955 -1.408 86.045 -0.4 ;
      RECT 85.905 -0.805 86.045 -0.635 ;
      RECT 85.955 0.4 86.045 1.408 ;
      RECT 85.905 0.635 86.045 0.805 ;
      RECT 84.525 -111.685 86.005 -111.585 ;
      RECT 84.525 -112.195 84.625 -111.585 ;
      RECT 84.745 -109.15 86.005 -109.05 ;
      RECT 85.905 -109.475 86.005 -109.05 ;
      RECT 85.345 -109.475 85.445 -109.05 ;
      RECT 84.785 -109.475 84.885 -109.05 ;
      RECT 85.555 -101.538 85.645 -100.531 ;
      RECT 85.555 -101.225 85.695 -101.055 ;
      RECT 85.555 -99.729 85.645 -98.722 ;
      RECT 85.555 -99.205 85.695 -99.035 ;
      RECT 85.555 -98.308 85.645 -97.301 ;
      RECT 85.555 -97.995 85.695 -97.825 ;
      RECT 85.555 -96.499 85.645 -95.492 ;
      RECT 85.555 -95.975 85.695 -95.805 ;
      RECT 85.555 -95.078 85.645 -94.071 ;
      RECT 85.555 -94.765 85.695 -94.595 ;
      RECT 85.555 -93.269 85.645 -92.262 ;
      RECT 85.555 -92.745 85.695 -92.575 ;
      RECT 85.555 -91.848 85.645 -90.841 ;
      RECT 85.555 -91.535 85.695 -91.365 ;
      RECT 85.555 -90.039 85.645 -89.032 ;
      RECT 85.555 -89.515 85.695 -89.345 ;
      RECT 85.555 -88.618 85.645 -87.611 ;
      RECT 85.555 -88.305 85.695 -88.135 ;
      RECT 85.555 -86.809 85.645 -85.802 ;
      RECT 85.555 -86.285 85.695 -86.115 ;
      RECT 85.555 -85.388 85.645 -84.381 ;
      RECT 85.555 -85.075 85.695 -84.905 ;
      RECT 85.555 -83.579 85.645 -82.572 ;
      RECT 85.555 -83.055 85.695 -82.885 ;
      RECT 85.555 -82.158 85.645 -81.151 ;
      RECT 85.555 -81.845 85.695 -81.675 ;
      RECT 85.555 -80.349 85.645 -79.342 ;
      RECT 85.555 -79.825 85.695 -79.655 ;
      RECT 85.555 -78.928 85.645 -77.921 ;
      RECT 85.555 -78.615 85.695 -78.445 ;
      RECT 85.555 -77.119 85.645 -76.112 ;
      RECT 85.555 -76.595 85.695 -76.425 ;
      RECT 85.555 -75.698 85.645 -74.691 ;
      RECT 85.555 -75.385 85.695 -75.215 ;
      RECT 85.555 -73.889 85.645 -72.882 ;
      RECT 85.555 -73.365 85.695 -73.195 ;
      RECT 85.555 -72.468 85.645 -71.461 ;
      RECT 85.555 -72.155 85.695 -71.985 ;
      RECT 85.555 -70.659 85.645 -69.652 ;
      RECT 85.555 -70.135 85.695 -69.965 ;
      RECT 85.555 -69.238 85.645 -68.231 ;
      RECT 85.555 -68.925 85.695 -68.755 ;
      RECT 85.555 -67.429 85.645 -66.422 ;
      RECT 85.555 -66.905 85.695 -66.735 ;
      RECT 85.555 -66.008 85.645 -65.001 ;
      RECT 85.555 -65.695 85.695 -65.525 ;
      RECT 85.555 -64.199 85.645 -63.192 ;
      RECT 85.555 -63.675 85.695 -63.505 ;
      RECT 85.555 -62.778 85.645 -61.771 ;
      RECT 85.555 -62.465 85.695 -62.295 ;
      RECT 85.555 -60.969 85.645 -59.962 ;
      RECT 85.555 -60.445 85.695 -60.275 ;
      RECT 85.555 -59.548 85.645 -58.541 ;
      RECT 85.555 -59.235 85.695 -59.065 ;
      RECT 85.555 -57.739 85.645 -56.732 ;
      RECT 85.555 -57.215 85.695 -57.045 ;
      RECT 85.555 -56.318 85.645 -55.311 ;
      RECT 85.555 -56.005 85.695 -55.835 ;
      RECT 85.555 -54.509 85.645 -53.502 ;
      RECT 85.555 -53.985 85.695 -53.815 ;
      RECT 85.555 -53.088 85.645 -52.081 ;
      RECT 85.555 -52.775 85.695 -52.605 ;
      RECT 85.555 -51.279 85.645 -50.272 ;
      RECT 85.555 -50.755 85.695 -50.585 ;
      RECT 85.555 -49.858 85.645 -48.851 ;
      RECT 85.555 -49.545 85.695 -49.375 ;
      RECT 85.555 -48.049 85.645 -47.042 ;
      RECT 85.555 -47.525 85.695 -47.355 ;
      RECT 85.555 -46.628 85.645 -45.621 ;
      RECT 85.555 -46.315 85.695 -46.145 ;
      RECT 85.555 -44.819 85.645 -43.812 ;
      RECT 85.555 -44.295 85.695 -44.125 ;
      RECT 85.555 -43.398 85.645 -42.391 ;
      RECT 85.555 -43.085 85.695 -42.915 ;
      RECT 85.555 -41.589 85.645 -40.582 ;
      RECT 85.555 -41.065 85.695 -40.895 ;
      RECT 85.555 -40.168 85.645 -39.161 ;
      RECT 85.555 -39.855 85.695 -39.685 ;
      RECT 85.555 -38.359 85.645 -37.352 ;
      RECT 85.555 -37.835 85.695 -37.665 ;
      RECT 85.555 -36.938 85.645 -35.931 ;
      RECT 85.555 -36.625 85.695 -36.455 ;
      RECT 85.555 -35.129 85.645 -34.122 ;
      RECT 85.555 -34.605 85.695 -34.435 ;
      RECT 85.555 -33.708 85.645 -32.701 ;
      RECT 85.555 -33.395 85.695 -33.225 ;
      RECT 85.555 -31.899 85.645 -30.892 ;
      RECT 85.555 -31.375 85.695 -31.205 ;
      RECT 85.555 -30.478 85.645 -29.471 ;
      RECT 85.555 -30.165 85.695 -29.995 ;
      RECT 85.555 -28.669 85.645 -27.662 ;
      RECT 85.555 -28.145 85.695 -27.975 ;
      RECT 85.555 -27.248 85.645 -26.241 ;
      RECT 85.555 -26.935 85.695 -26.765 ;
      RECT 85.555 -25.439 85.645 -24.432 ;
      RECT 85.555 -24.915 85.695 -24.745 ;
      RECT 85.555 -24.018 85.645 -23.011 ;
      RECT 85.555 -23.705 85.695 -23.535 ;
      RECT 85.555 -22.209 85.645 -21.202 ;
      RECT 85.555 -21.685 85.695 -21.515 ;
      RECT 85.555 -20.788 85.645 -19.781 ;
      RECT 85.555 -20.475 85.695 -20.305 ;
      RECT 85.555 -18.979 85.645 -17.972 ;
      RECT 85.555 -18.455 85.695 -18.285 ;
      RECT 85.555 -17.558 85.645 -16.551 ;
      RECT 85.555 -17.245 85.695 -17.075 ;
      RECT 85.555 -15.749 85.645 -14.742 ;
      RECT 85.555 -15.225 85.695 -15.055 ;
      RECT 85.555 -14.328 85.645 -13.321 ;
      RECT 85.555 -14.015 85.695 -13.845 ;
      RECT 85.555 -12.519 85.645 -11.512 ;
      RECT 85.555 -11.995 85.695 -11.825 ;
      RECT 85.555 -11.098 85.645 -10.091 ;
      RECT 85.555 -10.785 85.695 -10.615 ;
      RECT 85.555 -9.289 85.645 -8.282 ;
      RECT 85.555 -8.765 85.695 -8.595 ;
      RECT 85.555 -7.868 85.645 -6.861 ;
      RECT 85.555 -7.555 85.695 -7.385 ;
      RECT 85.555 -6.059 85.645 -5.052 ;
      RECT 85.555 -5.535 85.695 -5.365 ;
      RECT 85.555 -4.638 85.645 -3.631 ;
      RECT 85.555 -4.325 85.695 -4.155 ;
      RECT 85.555 -2.829 85.645 -1.822 ;
      RECT 85.555 -2.305 85.695 -2.135 ;
      RECT 85.555 -1.408 85.645 -0.401 ;
      RECT 85.555 -1.095 85.695 -0.925 ;
      RECT 85.555 0.401 85.645 1.408 ;
      RECT 85.555 0.925 85.695 1.095 ;
      RECT 84.885 -111.495 85.055 -111.385 ;
      RECT 81.735 -111.495 85.055 -111.395 ;
      RECT 84.755 -101.538 84.845 -100.53 ;
      RECT 84.705 -100.935 84.845 -100.765 ;
      RECT 84.755 -99.73 84.845 -98.722 ;
      RECT 84.705 -99.495 84.845 -99.325 ;
      RECT 84.755 -98.308 84.845 -97.3 ;
      RECT 84.705 -97.705 84.845 -97.535 ;
      RECT 84.755 -96.5 84.845 -95.492 ;
      RECT 84.705 -96.265 84.845 -96.095 ;
      RECT 84.755 -95.078 84.845 -94.07 ;
      RECT 84.705 -94.475 84.845 -94.305 ;
      RECT 84.755 -93.27 84.845 -92.262 ;
      RECT 84.705 -93.035 84.845 -92.865 ;
      RECT 84.755 -91.848 84.845 -90.84 ;
      RECT 84.705 -91.245 84.845 -91.075 ;
      RECT 84.755 -90.04 84.845 -89.032 ;
      RECT 84.705 -89.805 84.845 -89.635 ;
      RECT 84.755 -88.618 84.845 -87.61 ;
      RECT 84.705 -88.015 84.845 -87.845 ;
      RECT 84.755 -86.81 84.845 -85.802 ;
      RECT 84.705 -86.575 84.845 -86.405 ;
      RECT 84.755 -85.388 84.845 -84.38 ;
      RECT 84.705 -84.785 84.845 -84.615 ;
      RECT 84.755 -83.58 84.845 -82.572 ;
      RECT 84.705 -83.345 84.845 -83.175 ;
      RECT 84.755 -82.158 84.845 -81.15 ;
      RECT 84.705 -81.555 84.845 -81.385 ;
      RECT 84.755 -80.35 84.845 -79.342 ;
      RECT 84.705 -80.115 84.845 -79.945 ;
      RECT 84.755 -78.928 84.845 -77.92 ;
      RECT 84.705 -78.325 84.845 -78.155 ;
      RECT 84.755 -77.12 84.845 -76.112 ;
      RECT 84.705 -76.885 84.845 -76.715 ;
      RECT 84.755 -75.698 84.845 -74.69 ;
      RECT 84.705 -75.095 84.845 -74.925 ;
      RECT 84.755 -73.89 84.845 -72.882 ;
      RECT 84.705 -73.655 84.845 -73.485 ;
      RECT 84.755 -72.468 84.845 -71.46 ;
      RECT 84.705 -71.865 84.845 -71.695 ;
      RECT 84.755 -70.66 84.845 -69.652 ;
      RECT 84.705 -70.425 84.845 -70.255 ;
      RECT 84.755 -69.238 84.845 -68.23 ;
      RECT 84.705 -68.635 84.845 -68.465 ;
      RECT 84.755 -67.43 84.845 -66.422 ;
      RECT 84.705 -67.195 84.845 -67.025 ;
      RECT 84.755 -66.008 84.845 -65 ;
      RECT 84.705 -65.405 84.845 -65.235 ;
      RECT 84.755 -64.2 84.845 -63.192 ;
      RECT 84.705 -63.965 84.845 -63.795 ;
      RECT 84.755 -62.778 84.845 -61.77 ;
      RECT 84.705 -62.175 84.845 -62.005 ;
      RECT 84.755 -60.97 84.845 -59.962 ;
      RECT 84.705 -60.735 84.845 -60.565 ;
      RECT 84.755 -59.548 84.845 -58.54 ;
      RECT 84.705 -58.945 84.845 -58.775 ;
      RECT 84.755 -57.74 84.845 -56.732 ;
      RECT 84.705 -57.505 84.845 -57.335 ;
      RECT 84.755 -56.318 84.845 -55.31 ;
      RECT 84.705 -55.715 84.845 -55.545 ;
      RECT 84.755 -54.51 84.845 -53.502 ;
      RECT 84.705 -54.275 84.845 -54.105 ;
      RECT 84.755 -53.088 84.845 -52.08 ;
      RECT 84.705 -52.485 84.845 -52.315 ;
      RECT 84.755 -51.28 84.845 -50.272 ;
      RECT 84.705 -51.045 84.845 -50.875 ;
      RECT 84.755 -49.858 84.845 -48.85 ;
      RECT 84.705 -49.255 84.845 -49.085 ;
      RECT 84.755 -48.05 84.845 -47.042 ;
      RECT 84.705 -47.815 84.845 -47.645 ;
      RECT 84.755 -46.628 84.845 -45.62 ;
      RECT 84.705 -46.025 84.845 -45.855 ;
      RECT 84.755 -44.82 84.845 -43.812 ;
      RECT 84.705 -44.585 84.845 -44.415 ;
      RECT 84.755 -43.398 84.845 -42.39 ;
      RECT 84.705 -42.795 84.845 -42.625 ;
      RECT 84.755 -41.59 84.845 -40.582 ;
      RECT 84.705 -41.355 84.845 -41.185 ;
      RECT 84.755 -40.168 84.845 -39.16 ;
      RECT 84.705 -39.565 84.845 -39.395 ;
      RECT 84.755 -38.36 84.845 -37.352 ;
      RECT 84.705 -38.125 84.845 -37.955 ;
      RECT 84.755 -36.938 84.845 -35.93 ;
      RECT 84.705 -36.335 84.845 -36.165 ;
      RECT 84.755 -35.13 84.845 -34.122 ;
      RECT 84.705 -34.895 84.845 -34.725 ;
      RECT 84.755 -33.708 84.845 -32.7 ;
      RECT 84.705 -33.105 84.845 -32.935 ;
      RECT 84.755 -31.9 84.845 -30.892 ;
      RECT 84.705 -31.665 84.845 -31.495 ;
      RECT 84.755 -30.478 84.845 -29.47 ;
      RECT 84.705 -29.875 84.845 -29.705 ;
      RECT 84.755 -28.67 84.845 -27.662 ;
      RECT 84.705 -28.435 84.845 -28.265 ;
      RECT 84.755 -27.248 84.845 -26.24 ;
      RECT 84.705 -26.645 84.845 -26.475 ;
      RECT 84.755 -25.44 84.845 -24.432 ;
      RECT 84.705 -25.205 84.845 -25.035 ;
      RECT 84.755 -24.018 84.845 -23.01 ;
      RECT 84.705 -23.415 84.845 -23.245 ;
      RECT 84.755 -22.21 84.845 -21.202 ;
      RECT 84.705 -21.975 84.845 -21.805 ;
      RECT 84.755 -20.788 84.845 -19.78 ;
      RECT 84.705 -20.185 84.845 -20.015 ;
      RECT 84.755 -18.98 84.845 -17.972 ;
      RECT 84.705 -18.745 84.845 -18.575 ;
      RECT 84.755 -17.558 84.845 -16.55 ;
      RECT 84.705 -16.955 84.845 -16.785 ;
      RECT 84.755 -15.75 84.845 -14.742 ;
      RECT 84.705 -15.515 84.845 -15.345 ;
      RECT 84.755 -14.328 84.845 -13.32 ;
      RECT 84.705 -13.725 84.845 -13.555 ;
      RECT 84.755 -12.52 84.845 -11.512 ;
      RECT 84.705 -12.285 84.845 -12.115 ;
      RECT 84.755 -11.098 84.845 -10.09 ;
      RECT 84.705 -10.495 84.845 -10.325 ;
      RECT 84.755 -9.29 84.845 -8.282 ;
      RECT 84.705 -9.055 84.845 -8.885 ;
      RECT 84.755 -7.868 84.845 -6.86 ;
      RECT 84.705 -7.265 84.845 -7.095 ;
      RECT 84.755 -6.06 84.845 -5.052 ;
      RECT 84.705 -5.825 84.845 -5.655 ;
      RECT 84.755 -4.638 84.845 -3.63 ;
      RECT 84.705 -4.035 84.845 -3.865 ;
      RECT 84.755 -2.83 84.845 -1.822 ;
      RECT 84.705 -2.595 84.845 -2.425 ;
      RECT 84.755 -1.408 84.845 -0.4 ;
      RECT 84.705 -0.805 84.845 -0.635 ;
      RECT 84.755 0.4 84.845 1.408 ;
      RECT 84.705 0.635 84.845 0.805 ;
      RECT 84.355 -101.538 84.445 -100.531 ;
      RECT 84.355 -101.225 84.495 -101.055 ;
      RECT 84.355 -99.729 84.445 -98.722 ;
      RECT 84.355 -99.205 84.495 -99.035 ;
      RECT 84.355 -98.308 84.445 -97.301 ;
      RECT 84.355 -97.995 84.495 -97.825 ;
      RECT 84.355 -96.499 84.445 -95.492 ;
      RECT 84.355 -95.975 84.495 -95.805 ;
      RECT 84.355 -95.078 84.445 -94.071 ;
      RECT 84.355 -94.765 84.495 -94.595 ;
      RECT 84.355 -93.269 84.445 -92.262 ;
      RECT 84.355 -92.745 84.495 -92.575 ;
      RECT 84.355 -91.848 84.445 -90.841 ;
      RECT 84.355 -91.535 84.495 -91.365 ;
      RECT 84.355 -90.039 84.445 -89.032 ;
      RECT 84.355 -89.515 84.495 -89.345 ;
      RECT 84.355 -88.618 84.445 -87.611 ;
      RECT 84.355 -88.305 84.495 -88.135 ;
      RECT 84.355 -86.809 84.445 -85.802 ;
      RECT 84.355 -86.285 84.495 -86.115 ;
      RECT 84.355 -85.388 84.445 -84.381 ;
      RECT 84.355 -85.075 84.495 -84.905 ;
      RECT 84.355 -83.579 84.445 -82.572 ;
      RECT 84.355 -83.055 84.495 -82.885 ;
      RECT 84.355 -82.158 84.445 -81.151 ;
      RECT 84.355 -81.845 84.495 -81.675 ;
      RECT 84.355 -80.349 84.445 -79.342 ;
      RECT 84.355 -79.825 84.495 -79.655 ;
      RECT 84.355 -78.928 84.445 -77.921 ;
      RECT 84.355 -78.615 84.495 -78.445 ;
      RECT 84.355 -77.119 84.445 -76.112 ;
      RECT 84.355 -76.595 84.495 -76.425 ;
      RECT 84.355 -75.698 84.445 -74.691 ;
      RECT 84.355 -75.385 84.495 -75.215 ;
      RECT 84.355 -73.889 84.445 -72.882 ;
      RECT 84.355 -73.365 84.495 -73.195 ;
      RECT 84.355 -72.468 84.445 -71.461 ;
      RECT 84.355 -72.155 84.495 -71.985 ;
      RECT 84.355 -70.659 84.445 -69.652 ;
      RECT 84.355 -70.135 84.495 -69.965 ;
      RECT 84.355 -69.238 84.445 -68.231 ;
      RECT 84.355 -68.925 84.495 -68.755 ;
      RECT 84.355 -67.429 84.445 -66.422 ;
      RECT 84.355 -66.905 84.495 -66.735 ;
      RECT 84.355 -66.008 84.445 -65.001 ;
      RECT 84.355 -65.695 84.495 -65.525 ;
      RECT 84.355 -64.199 84.445 -63.192 ;
      RECT 84.355 -63.675 84.495 -63.505 ;
      RECT 84.355 -62.778 84.445 -61.771 ;
      RECT 84.355 -62.465 84.495 -62.295 ;
      RECT 84.355 -60.969 84.445 -59.962 ;
      RECT 84.355 -60.445 84.495 -60.275 ;
      RECT 84.355 -59.548 84.445 -58.541 ;
      RECT 84.355 -59.235 84.495 -59.065 ;
      RECT 84.355 -57.739 84.445 -56.732 ;
      RECT 84.355 -57.215 84.495 -57.045 ;
      RECT 84.355 -56.318 84.445 -55.311 ;
      RECT 84.355 -56.005 84.495 -55.835 ;
      RECT 84.355 -54.509 84.445 -53.502 ;
      RECT 84.355 -53.985 84.495 -53.815 ;
      RECT 84.355 -53.088 84.445 -52.081 ;
      RECT 84.355 -52.775 84.495 -52.605 ;
      RECT 84.355 -51.279 84.445 -50.272 ;
      RECT 84.355 -50.755 84.495 -50.585 ;
      RECT 84.355 -49.858 84.445 -48.851 ;
      RECT 84.355 -49.545 84.495 -49.375 ;
      RECT 84.355 -48.049 84.445 -47.042 ;
      RECT 84.355 -47.525 84.495 -47.355 ;
      RECT 84.355 -46.628 84.445 -45.621 ;
      RECT 84.355 -46.315 84.495 -46.145 ;
      RECT 84.355 -44.819 84.445 -43.812 ;
      RECT 84.355 -44.295 84.495 -44.125 ;
      RECT 84.355 -43.398 84.445 -42.391 ;
      RECT 84.355 -43.085 84.495 -42.915 ;
      RECT 84.355 -41.589 84.445 -40.582 ;
      RECT 84.355 -41.065 84.495 -40.895 ;
      RECT 84.355 -40.168 84.445 -39.161 ;
      RECT 84.355 -39.855 84.495 -39.685 ;
      RECT 84.355 -38.359 84.445 -37.352 ;
      RECT 84.355 -37.835 84.495 -37.665 ;
      RECT 84.355 -36.938 84.445 -35.931 ;
      RECT 84.355 -36.625 84.495 -36.455 ;
      RECT 84.355 -35.129 84.445 -34.122 ;
      RECT 84.355 -34.605 84.495 -34.435 ;
      RECT 84.355 -33.708 84.445 -32.701 ;
      RECT 84.355 -33.395 84.495 -33.225 ;
      RECT 84.355 -31.899 84.445 -30.892 ;
      RECT 84.355 -31.375 84.495 -31.205 ;
      RECT 84.355 -30.478 84.445 -29.471 ;
      RECT 84.355 -30.165 84.495 -29.995 ;
      RECT 84.355 -28.669 84.445 -27.662 ;
      RECT 84.355 -28.145 84.495 -27.975 ;
      RECT 84.355 -27.248 84.445 -26.241 ;
      RECT 84.355 -26.935 84.495 -26.765 ;
      RECT 84.355 -25.439 84.445 -24.432 ;
      RECT 84.355 -24.915 84.495 -24.745 ;
      RECT 84.355 -24.018 84.445 -23.011 ;
      RECT 84.355 -23.705 84.495 -23.535 ;
      RECT 84.355 -22.209 84.445 -21.202 ;
      RECT 84.355 -21.685 84.495 -21.515 ;
      RECT 84.355 -20.788 84.445 -19.781 ;
      RECT 84.355 -20.475 84.495 -20.305 ;
      RECT 84.355 -18.979 84.445 -17.972 ;
      RECT 84.355 -18.455 84.495 -18.285 ;
      RECT 84.355 -17.558 84.445 -16.551 ;
      RECT 84.355 -17.245 84.495 -17.075 ;
      RECT 84.355 -15.749 84.445 -14.742 ;
      RECT 84.355 -15.225 84.495 -15.055 ;
      RECT 84.355 -14.328 84.445 -13.321 ;
      RECT 84.355 -14.015 84.495 -13.845 ;
      RECT 84.355 -12.519 84.445 -11.512 ;
      RECT 84.355 -11.995 84.495 -11.825 ;
      RECT 84.355 -11.098 84.445 -10.091 ;
      RECT 84.355 -10.785 84.495 -10.615 ;
      RECT 84.355 -9.289 84.445 -8.282 ;
      RECT 84.355 -8.765 84.495 -8.595 ;
      RECT 84.355 -7.868 84.445 -6.861 ;
      RECT 84.355 -7.555 84.495 -7.385 ;
      RECT 84.355 -6.059 84.445 -5.052 ;
      RECT 84.355 -5.535 84.495 -5.365 ;
      RECT 84.355 -4.638 84.445 -3.631 ;
      RECT 84.355 -4.325 84.495 -4.155 ;
      RECT 84.355 -2.829 84.445 -1.822 ;
      RECT 84.355 -2.305 84.495 -2.135 ;
      RECT 84.355 -1.408 84.445 -0.401 ;
      RECT 84.355 -1.095 84.495 -0.925 ;
      RECT 84.355 0.401 84.445 1.408 ;
      RECT 84.355 0.925 84.495 1.095 ;
      RECT 82.505 -111.685 83.985 -111.585 ;
      RECT 82.505 -112.055 82.605 -111.585 ;
      RECT 82.31 -114.395 83.885 -114.275 ;
      RECT 83.785 -114.895 83.885 -114.275 ;
      RECT 83.19 -114.895 83.29 -114.275 ;
      RECT 82.31 -114.85 82.41 -114.275 ;
      RECT 83.555 -101.538 83.645 -100.53 ;
      RECT 83.505 -100.935 83.645 -100.765 ;
      RECT 83.555 -99.73 83.645 -98.722 ;
      RECT 83.505 -99.495 83.645 -99.325 ;
      RECT 83.555 -98.308 83.645 -97.3 ;
      RECT 83.505 -97.705 83.645 -97.535 ;
      RECT 83.555 -96.5 83.645 -95.492 ;
      RECT 83.505 -96.265 83.645 -96.095 ;
      RECT 83.555 -95.078 83.645 -94.07 ;
      RECT 83.505 -94.475 83.645 -94.305 ;
      RECT 83.555 -93.27 83.645 -92.262 ;
      RECT 83.505 -93.035 83.645 -92.865 ;
      RECT 83.555 -91.848 83.645 -90.84 ;
      RECT 83.505 -91.245 83.645 -91.075 ;
      RECT 83.555 -90.04 83.645 -89.032 ;
      RECT 83.505 -89.805 83.645 -89.635 ;
      RECT 83.555 -88.618 83.645 -87.61 ;
      RECT 83.505 -88.015 83.645 -87.845 ;
      RECT 83.555 -86.81 83.645 -85.802 ;
      RECT 83.505 -86.575 83.645 -86.405 ;
      RECT 83.555 -85.388 83.645 -84.38 ;
      RECT 83.505 -84.785 83.645 -84.615 ;
      RECT 83.555 -83.58 83.645 -82.572 ;
      RECT 83.505 -83.345 83.645 -83.175 ;
      RECT 83.555 -82.158 83.645 -81.15 ;
      RECT 83.505 -81.555 83.645 -81.385 ;
      RECT 83.555 -80.35 83.645 -79.342 ;
      RECT 83.505 -80.115 83.645 -79.945 ;
      RECT 83.555 -78.928 83.645 -77.92 ;
      RECT 83.505 -78.325 83.645 -78.155 ;
      RECT 83.555 -77.12 83.645 -76.112 ;
      RECT 83.505 -76.885 83.645 -76.715 ;
      RECT 83.555 -75.698 83.645 -74.69 ;
      RECT 83.505 -75.095 83.645 -74.925 ;
      RECT 83.555 -73.89 83.645 -72.882 ;
      RECT 83.505 -73.655 83.645 -73.485 ;
      RECT 83.555 -72.468 83.645 -71.46 ;
      RECT 83.505 -71.865 83.645 -71.695 ;
      RECT 83.555 -70.66 83.645 -69.652 ;
      RECT 83.505 -70.425 83.645 -70.255 ;
      RECT 83.555 -69.238 83.645 -68.23 ;
      RECT 83.505 -68.635 83.645 -68.465 ;
      RECT 83.555 -67.43 83.645 -66.422 ;
      RECT 83.505 -67.195 83.645 -67.025 ;
      RECT 83.555 -66.008 83.645 -65 ;
      RECT 83.505 -65.405 83.645 -65.235 ;
      RECT 83.555 -64.2 83.645 -63.192 ;
      RECT 83.505 -63.965 83.645 -63.795 ;
      RECT 83.555 -62.778 83.645 -61.77 ;
      RECT 83.505 -62.175 83.645 -62.005 ;
      RECT 83.555 -60.97 83.645 -59.962 ;
      RECT 83.505 -60.735 83.645 -60.565 ;
      RECT 83.555 -59.548 83.645 -58.54 ;
      RECT 83.505 -58.945 83.645 -58.775 ;
      RECT 83.555 -57.74 83.645 -56.732 ;
      RECT 83.505 -57.505 83.645 -57.335 ;
      RECT 83.555 -56.318 83.645 -55.31 ;
      RECT 83.505 -55.715 83.645 -55.545 ;
      RECT 83.555 -54.51 83.645 -53.502 ;
      RECT 83.505 -54.275 83.645 -54.105 ;
      RECT 83.555 -53.088 83.645 -52.08 ;
      RECT 83.505 -52.485 83.645 -52.315 ;
      RECT 83.555 -51.28 83.645 -50.272 ;
      RECT 83.505 -51.045 83.645 -50.875 ;
      RECT 83.555 -49.858 83.645 -48.85 ;
      RECT 83.505 -49.255 83.645 -49.085 ;
      RECT 83.555 -48.05 83.645 -47.042 ;
      RECT 83.505 -47.815 83.645 -47.645 ;
      RECT 83.555 -46.628 83.645 -45.62 ;
      RECT 83.505 -46.025 83.645 -45.855 ;
      RECT 83.555 -44.82 83.645 -43.812 ;
      RECT 83.505 -44.585 83.645 -44.415 ;
      RECT 83.555 -43.398 83.645 -42.39 ;
      RECT 83.505 -42.795 83.645 -42.625 ;
      RECT 83.555 -41.59 83.645 -40.582 ;
      RECT 83.505 -41.355 83.645 -41.185 ;
      RECT 83.555 -40.168 83.645 -39.16 ;
      RECT 83.505 -39.565 83.645 -39.395 ;
      RECT 83.555 -38.36 83.645 -37.352 ;
      RECT 83.505 -38.125 83.645 -37.955 ;
      RECT 83.555 -36.938 83.645 -35.93 ;
      RECT 83.505 -36.335 83.645 -36.165 ;
      RECT 83.555 -35.13 83.645 -34.122 ;
      RECT 83.505 -34.895 83.645 -34.725 ;
      RECT 83.555 -33.708 83.645 -32.7 ;
      RECT 83.505 -33.105 83.645 -32.935 ;
      RECT 83.555 -31.9 83.645 -30.892 ;
      RECT 83.505 -31.665 83.645 -31.495 ;
      RECT 83.555 -30.478 83.645 -29.47 ;
      RECT 83.505 -29.875 83.645 -29.705 ;
      RECT 83.555 -28.67 83.645 -27.662 ;
      RECT 83.505 -28.435 83.645 -28.265 ;
      RECT 83.555 -27.248 83.645 -26.24 ;
      RECT 83.505 -26.645 83.645 -26.475 ;
      RECT 83.555 -25.44 83.645 -24.432 ;
      RECT 83.505 -25.205 83.645 -25.035 ;
      RECT 83.555 -24.018 83.645 -23.01 ;
      RECT 83.505 -23.415 83.645 -23.245 ;
      RECT 83.555 -22.21 83.645 -21.202 ;
      RECT 83.505 -21.975 83.645 -21.805 ;
      RECT 83.555 -20.788 83.645 -19.78 ;
      RECT 83.505 -20.185 83.645 -20.015 ;
      RECT 83.555 -18.98 83.645 -17.972 ;
      RECT 83.505 -18.745 83.645 -18.575 ;
      RECT 83.555 -17.558 83.645 -16.55 ;
      RECT 83.505 -16.955 83.645 -16.785 ;
      RECT 83.555 -15.75 83.645 -14.742 ;
      RECT 83.505 -15.515 83.645 -15.345 ;
      RECT 83.555 -14.328 83.645 -13.32 ;
      RECT 83.505 -13.725 83.645 -13.555 ;
      RECT 83.555 -12.52 83.645 -11.512 ;
      RECT 83.505 -12.285 83.645 -12.115 ;
      RECT 83.555 -11.098 83.645 -10.09 ;
      RECT 83.505 -10.495 83.645 -10.325 ;
      RECT 83.555 -9.29 83.645 -8.282 ;
      RECT 83.505 -9.055 83.645 -8.885 ;
      RECT 83.555 -7.868 83.645 -6.86 ;
      RECT 83.505 -7.265 83.645 -7.095 ;
      RECT 83.555 -6.06 83.645 -5.052 ;
      RECT 83.505 -5.825 83.645 -5.655 ;
      RECT 83.555 -4.638 83.645 -3.63 ;
      RECT 83.505 -4.035 83.645 -3.865 ;
      RECT 83.555 -2.83 83.645 -1.822 ;
      RECT 83.505 -2.595 83.645 -2.425 ;
      RECT 83.555 -1.408 83.645 -0.4 ;
      RECT 83.505 -0.805 83.645 -0.635 ;
      RECT 83.555 0.4 83.645 1.408 ;
      RECT 83.505 0.635 83.645 0.805 ;
      RECT 83.43 -114.685 83.605 -114.515 ;
      RECT 83.505 -114.895 83.605 -114.515 ;
      RECT 82.545 -113.555 82.645 -113.09 ;
      RECT 82.91 -113.555 83.01 -113.1 ;
      RECT 82.545 -113.555 83.39 -113.385 ;
      RECT 83.155 -101.538 83.245 -100.531 ;
      RECT 83.155 -101.225 83.295 -101.055 ;
      RECT 83.155 -99.729 83.245 -98.722 ;
      RECT 83.155 -99.205 83.295 -99.035 ;
      RECT 83.155 -98.308 83.245 -97.301 ;
      RECT 83.155 -97.995 83.295 -97.825 ;
      RECT 83.155 -96.499 83.245 -95.492 ;
      RECT 83.155 -95.975 83.295 -95.805 ;
      RECT 83.155 -95.078 83.245 -94.071 ;
      RECT 83.155 -94.765 83.295 -94.595 ;
      RECT 83.155 -93.269 83.245 -92.262 ;
      RECT 83.155 -92.745 83.295 -92.575 ;
      RECT 83.155 -91.848 83.245 -90.841 ;
      RECT 83.155 -91.535 83.295 -91.365 ;
      RECT 83.155 -90.039 83.245 -89.032 ;
      RECT 83.155 -89.515 83.295 -89.345 ;
      RECT 83.155 -88.618 83.245 -87.611 ;
      RECT 83.155 -88.305 83.295 -88.135 ;
      RECT 83.155 -86.809 83.245 -85.802 ;
      RECT 83.155 -86.285 83.295 -86.115 ;
      RECT 83.155 -85.388 83.245 -84.381 ;
      RECT 83.155 -85.075 83.295 -84.905 ;
      RECT 83.155 -83.579 83.245 -82.572 ;
      RECT 83.155 -83.055 83.295 -82.885 ;
      RECT 83.155 -82.158 83.245 -81.151 ;
      RECT 83.155 -81.845 83.295 -81.675 ;
      RECT 83.155 -80.349 83.245 -79.342 ;
      RECT 83.155 -79.825 83.295 -79.655 ;
      RECT 83.155 -78.928 83.245 -77.921 ;
      RECT 83.155 -78.615 83.295 -78.445 ;
      RECT 83.155 -77.119 83.245 -76.112 ;
      RECT 83.155 -76.595 83.295 -76.425 ;
      RECT 83.155 -75.698 83.245 -74.691 ;
      RECT 83.155 -75.385 83.295 -75.215 ;
      RECT 83.155 -73.889 83.245 -72.882 ;
      RECT 83.155 -73.365 83.295 -73.195 ;
      RECT 83.155 -72.468 83.245 -71.461 ;
      RECT 83.155 -72.155 83.295 -71.985 ;
      RECT 83.155 -70.659 83.245 -69.652 ;
      RECT 83.155 -70.135 83.295 -69.965 ;
      RECT 83.155 -69.238 83.245 -68.231 ;
      RECT 83.155 -68.925 83.295 -68.755 ;
      RECT 83.155 -67.429 83.245 -66.422 ;
      RECT 83.155 -66.905 83.295 -66.735 ;
      RECT 83.155 -66.008 83.245 -65.001 ;
      RECT 83.155 -65.695 83.295 -65.525 ;
      RECT 83.155 -64.199 83.245 -63.192 ;
      RECT 83.155 -63.675 83.295 -63.505 ;
      RECT 83.155 -62.778 83.245 -61.771 ;
      RECT 83.155 -62.465 83.295 -62.295 ;
      RECT 83.155 -60.969 83.245 -59.962 ;
      RECT 83.155 -60.445 83.295 -60.275 ;
      RECT 83.155 -59.548 83.245 -58.541 ;
      RECT 83.155 -59.235 83.295 -59.065 ;
      RECT 83.155 -57.739 83.245 -56.732 ;
      RECT 83.155 -57.215 83.295 -57.045 ;
      RECT 83.155 -56.318 83.245 -55.311 ;
      RECT 83.155 -56.005 83.295 -55.835 ;
      RECT 83.155 -54.509 83.245 -53.502 ;
      RECT 83.155 -53.985 83.295 -53.815 ;
      RECT 83.155 -53.088 83.245 -52.081 ;
      RECT 83.155 -52.775 83.295 -52.605 ;
      RECT 83.155 -51.279 83.245 -50.272 ;
      RECT 83.155 -50.755 83.295 -50.585 ;
      RECT 83.155 -49.858 83.245 -48.851 ;
      RECT 83.155 -49.545 83.295 -49.375 ;
      RECT 83.155 -48.049 83.245 -47.042 ;
      RECT 83.155 -47.525 83.295 -47.355 ;
      RECT 83.155 -46.628 83.245 -45.621 ;
      RECT 83.155 -46.315 83.295 -46.145 ;
      RECT 83.155 -44.819 83.245 -43.812 ;
      RECT 83.155 -44.295 83.295 -44.125 ;
      RECT 83.155 -43.398 83.245 -42.391 ;
      RECT 83.155 -43.085 83.295 -42.915 ;
      RECT 83.155 -41.589 83.245 -40.582 ;
      RECT 83.155 -41.065 83.295 -40.895 ;
      RECT 83.155 -40.168 83.245 -39.161 ;
      RECT 83.155 -39.855 83.295 -39.685 ;
      RECT 83.155 -38.359 83.245 -37.352 ;
      RECT 83.155 -37.835 83.295 -37.665 ;
      RECT 83.155 -36.938 83.245 -35.931 ;
      RECT 83.155 -36.625 83.295 -36.455 ;
      RECT 83.155 -35.129 83.245 -34.122 ;
      RECT 83.155 -34.605 83.295 -34.435 ;
      RECT 83.155 -33.708 83.245 -32.701 ;
      RECT 83.155 -33.395 83.295 -33.225 ;
      RECT 83.155 -31.899 83.245 -30.892 ;
      RECT 83.155 -31.375 83.295 -31.205 ;
      RECT 83.155 -30.478 83.245 -29.471 ;
      RECT 83.155 -30.165 83.295 -29.995 ;
      RECT 83.155 -28.669 83.245 -27.662 ;
      RECT 83.155 -28.145 83.295 -27.975 ;
      RECT 83.155 -27.248 83.245 -26.241 ;
      RECT 83.155 -26.935 83.295 -26.765 ;
      RECT 83.155 -25.439 83.245 -24.432 ;
      RECT 83.155 -24.915 83.295 -24.745 ;
      RECT 83.155 -24.018 83.245 -23.011 ;
      RECT 83.155 -23.705 83.295 -23.535 ;
      RECT 83.155 -22.209 83.245 -21.202 ;
      RECT 83.155 -21.685 83.295 -21.515 ;
      RECT 83.155 -20.788 83.245 -19.781 ;
      RECT 83.155 -20.475 83.295 -20.305 ;
      RECT 83.155 -18.979 83.245 -17.972 ;
      RECT 83.155 -18.455 83.295 -18.285 ;
      RECT 83.155 -17.558 83.245 -16.551 ;
      RECT 83.155 -17.245 83.295 -17.075 ;
      RECT 83.155 -15.749 83.245 -14.742 ;
      RECT 83.155 -15.225 83.295 -15.055 ;
      RECT 83.155 -14.328 83.245 -13.321 ;
      RECT 83.155 -14.015 83.295 -13.845 ;
      RECT 83.155 -12.519 83.245 -11.512 ;
      RECT 83.155 -11.995 83.295 -11.825 ;
      RECT 83.155 -11.098 83.245 -10.091 ;
      RECT 83.155 -10.785 83.295 -10.615 ;
      RECT 83.155 -9.289 83.245 -8.282 ;
      RECT 83.155 -8.765 83.295 -8.595 ;
      RECT 83.155 -7.868 83.245 -6.861 ;
      RECT 83.155 -7.555 83.295 -7.385 ;
      RECT 83.155 -6.059 83.245 -5.052 ;
      RECT 83.155 -5.535 83.295 -5.365 ;
      RECT 83.155 -4.638 83.245 -3.631 ;
      RECT 83.155 -4.325 83.295 -4.155 ;
      RECT 83.155 -2.829 83.245 -1.822 ;
      RECT 83.155 -2.305 83.295 -2.135 ;
      RECT 83.155 -1.408 83.245 -0.401 ;
      RECT 83.155 -1.095 83.295 -0.925 ;
      RECT 83.155 0.401 83.245 1.408 ;
      RECT 83.155 0.925 83.295 1.095 ;
      RECT 82.84 -114.685 83.01 -114.515 ;
      RECT 82.91 -114.895 83.01 -114.515 ;
      RECT 82.355 -101.538 82.445 -100.53 ;
      RECT 82.305 -100.935 82.445 -100.765 ;
      RECT 82.355 -99.73 82.445 -98.722 ;
      RECT 82.305 -99.495 82.445 -99.325 ;
      RECT 82.355 -98.308 82.445 -97.3 ;
      RECT 82.305 -97.705 82.445 -97.535 ;
      RECT 82.355 -96.5 82.445 -95.492 ;
      RECT 82.305 -96.265 82.445 -96.095 ;
      RECT 82.355 -95.078 82.445 -94.07 ;
      RECT 82.305 -94.475 82.445 -94.305 ;
      RECT 82.355 -93.27 82.445 -92.262 ;
      RECT 82.305 -93.035 82.445 -92.865 ;
      RECT 82.355 -91.848 82.445 -90.84 ;
      RECT 82.305 -91.245 82.445 -91.075 ;
      RECT 82.355 -90.04 82.445 -89.032 ;
      RECT 82.305 -89.805 82.445 -89.635 ;
      RECT 82.355 -88.618 82.445 -87.61 ;
      RECT 82.305 -88.015 82.445 -87.845 ;
      RECT 82.355 -86.81 82.445 -85.802 ;
      RECT 82.305 -86.575 82.445 -86.405 ;
      RECT 82.355 -85.388 82.445 -84.38 ;
      RECT 82.305 -84.785 82.445 -84.615 ;
      RECT 82.355 -83.58 82.445 -82.572 ;
      RECT 82.305 -83.345 82.445 -83.175 ;
      RECT 82.355 -82.158 82.445 -81.15 ;
      RECT 82.305 -81.555 82.445 -81.385 ;
      RECT 82.355 -80.35 82.445 -79.342 ;
      RECT 82.305 -80.115 82.445 -79.945 ;
      RECT 82.355 -78.928 82.445 -77.92 ;
      RECT 82.305 -78.325 82.445 -78.155 ;
      RECT 82.355 -77.12 82.445 -76.112 ;
      RECT 82.305 -76.885 82.445 -76.715 ;
      RECT 82.355 -75.698 82.445 -74.69 ;
      RECT 82.305 -75.095 82.445 -74.925 ;
      RECT 82.355 -73.89 82.445 -72.882 ;
      RECT 82.305 -73.655 82.445 -73.485 ;
      RECT 82.355 -72.468 82.445 -71.46 ;
      RECT 82.305 -71.865 82.445 -71.695 ;
      RECT 82.355 -70.66 82.445 -69.652 ;
      RECT 82.305 -70.425 82.445 -70.255 ;
      RECT 82.355 -69.238 82.445 -68.23 ;
      RECT 82.305 -68.635 82.445 -68.465 ;
      RECT 82.355 -67.43 82.445 -66.422 ;
      RECT 82.305 -67.195 82.445 -67.025 ;
      RECT 82.355 -66.008 82.445 -65 ;
      RECT 82.305 -65.405 82.445 -65.235 ;
      RECT 82.355 -64.2 82.445 -63.192 ;
      RECT 82.305 -63.965 82.445 -63.795 ;
      RECT 82.355 -62.778 82.445 -61.77 ;
      RECT 82.305 -62.175 82.445 -62.005 ;
      RECT 82.355 -60.97 82.445 -59.962 ;
      RECT 82.305 -60.735 82.445 -60.565 ;
      RECT 82.355 -59.548 82.445 -58.54 ;
      RECT 82.305 -58.945 82.445 -58.775 ;
      RECT 82.355 -57.74 82.445 -56.732 ;
      RECT 82.305 -57.505 82.445 -57.335 ;
      RECT 82.355 -56.318 82.445 -55.31 ;
      RECT 82.305 -55.715 82.445 -55.545 ;
      RECT 82.355 -54.51 82.445 -53.502 ;
      RECT 82.305 -54.275 82.445 -54.105 ;
      RECT 82.355 -53.088 82.445 -52.08 ;
      RECT 82.305 -52.485 82.445 -52.315 ;
      RECT 82.355 -51.28 82.445 -50.272 ;
      RECT 82.305 -51.045 82.445 -50.875 ;
      RECT 82.355 -49.858 82.445 -48.85 ;
      RECT 82.305 -49.255 82.445 -49.085 ;
      RECT 82.355 -48.05 82.445 -47.042 ;
      RECT 82.305 -47.815 82.445 -47.645 ;
      RECT 82.355 -46.628 82.445 -45.62 ;
      RECT 82.305 -46.025 82.445 -45.855 ;
      RECT 82.355 -44.82 82.445 -43.812 ;
      RECT 82.305 -44.585 82.445 -44.415 ;
      RECT 82.355 -43.398 82.445 -42.39 ;
      RECT 82.305 -42.795 82.445 -42.625 ;
      RECT 82.355 -41.59 82.445 -40.582 ;
      RECT 82.305 -41.355 82.445 -41.185 ;
      RECT 82.355 -40.168 82.445 -39.16 ;
      RECT 82.305 -39.565 82.445 -39.395 ;
      RECT 82.355 -38.36 82.445 -37.352 ;
      RECT 82.305 -38.125 82.445 -37.955 ;
      RECT 82.355 -36.938 82.445 -35.93 ;
      RECT 82.305 -36.335 82.445 -36.165 ;
      RECT 82.355 -35.13 82.445 -34.122 ;
      RECT 82.305 -34.895 82.445 -34.725 ;
      RECT 82.355 -33.708 82.445 -32.7 ;
      RECT 82.305 -33.105 82.445 -32.935 ;
      RECT 82.355 -31.9 82.445 -30.892 ;
      RECT 82.305 -31.665 82.445 -31.495 ;
      RECT 82.355 -30.478 82.445 -29.47 ;
      RECT 82.305 -29.875 82.445 -29.705 ;
      RECT 82.355 -28.67 82.445 -27.662 ;
      RECT 82.305 -28.435 82.445 -28.265 ;
      RECT 82.355 -27.248 82.445 -26.24 ;
      RECT 82.305 -26.645 82.445 -26.475 ;
      RECT 82.355 -25.44 82.445 -24.432 ;
      RECT 82.305 -25.205 82.445 -25.035 ;
      RECT 82.355 -24.018 82.445 -23.01 ;
      RECT 82.305 -23.415 82.445 -23.245 ;
      RECT 82.355 -22.21 82.445 -21.202 ;
      RECT 82.305 -21.975 82.445 -21.805 ;
      RECT 82.355 -20.788 82.445 -19.78 ;
      RECT 82.305 -20.185 82.445 -20.015 ;
      RECT 82.355 -18.98 82.445 -17.972 ;
      RECT 82.305 -18.745 82.445 -18.575 ;
      RECT 82.355 -17.558 82.445 -16.55 ;
      RECT 82.305 -16.955 82.445 -16.785 ;
      RECT 82.355 -15.75 82.445 -14.742 ;
      RECT 82.305 -15.515 82.445 -15.345 ;
      RECT 82.355 -14.328 82.445 -13.32 ;
      RECT 82.305 -13.725 82.445 -13.555 ;
      RECT 82.355 -12.52 82.445 -11.512 ;
      RECT 82.305 -12.285 82.445 -12.115 ;
      RECT 82.355 -11.098 82.445 -10.09 ;
      RECT 82.305 -10.495 82.445 -10.325 ;
      RECT 82.355 -9.29 82.445 -8.282 ;
      RECT 82.305 -9.055 82.445 -8.885 ;
      RECT 82.355 -7.868 82.445 -6.86 ;
      RECT 82.305 -7.265 82.445 -7.095 ;
      RECT 82.355 -6.06 82.445 -5.052 ;
      RECT 82.305 -5.825 82.445 -5.655 ;
      RECT 82.355 -4.638 82.445 -3.63 ;
      RECT 82.305 -4.035 82.445 -3.865 ;
      RECT 82.355 -2.83 82.445 -1.822 ;
      RECT 82.305 -2.595 82.445 -2.425 ;
      RECT 82.355 -1.408 82.445 -0.4 ;
      RECT 82.305 -0.805 82.445 -0.635 ;
      RECT 82.355 0.4 82.445 1.408 ;
      RECT 82.305 0.635 82.445 0.805 ;
      RECT 81.955 -101.538 82.045 -100.531 ;
      RECT 81.955 -101.225 82.095 -101.055 ;
      RECT 81.955 -99.729 82.045 -98.722 ;
      RECT 81.955 -99.205 82.095 -99.035 ;
      RECT 81.955 -98.308 82.045 -97.301 ;
      RECT 81.955 -97.995 82.095 -97.825 ;
      RECT 81.955 -96.499 82.045 -95.492 ;
      RECT 81.955 -95.975 82.095 -95.805 ;
      RECT 81.955 -95.078 82.045 -94.071 ;
      RECT 81.955 -94.765 82.095 -94.595 ;
      RECT 81.955 -93.269 82.045 -92.262 ;
      RECT 81.955 -92.745 82.095 -92.575 ;
      RECT 81.955 -91.848 82.045 -90.841 ;
      RECT 81.955 -91.535 82.095 -91.365 ;
      RECT 81.955 -90.039 82.045 -89.032 ;
      RECT 81.955 -89.515 82.095 -89.345 ;
      RECT 81.955 -88.618 82.045 -87.611 ;
      RECT 81.955 -88.305 82.095 -88.135 ;
      RECT 81.955 -86.809 82.045 -85.802 ;
      RECT 81.955 -86.285 82.095 -86.115 ;
      RECT 81.955 -85.388 82.045 -84.381 ;
      RECT 81.955 -85.075 82.095 -84.905 ;
      RECT 81.955 -83.579 82.045 -82.572 ;
      RECT 81.955 -83.055 82.095 -82.885 ;
      RECT 81.955 -82.158 82.045 -81.151 ;
      RECT 81.955 -81.845 82.095 -81.675 ;
      RECT 81.955 -80.349 82.045 -79.342 ;
      RECT 81.955 -79.825 82.095 -79.655 ;
      RECT 81.955 -78.928 82.045 -77.921 ;
      RECT 81.955 -78.615 82.095 -78.445 ;
      RECT 81.955 -77.119 82.045 -76.112 ;
      RECT 81.955 -76.595 82.095 -76.425 ;
      RECT 81.955 -75.698 82.045 -74.691 ;
      RECT 81.955 -75.385 82.095 -75.215 ;
      RECT 81.955 -73.889 82.045 -72.882 ;
      RECT 81.955 -73.365 82.095 -73.195 ;
      RECT 81.955 -72.468 82.045 -71.461 ;
      RECT 81.955 -72.155 82.095 -71.985 ;
      RECT 81.955 -70.659 82.045 -69.652 ;
      RECT 81.955 -70.135 82.095 -69.965 ;
      RECT 81.955 -69.238 82.045 -68.231 ;
      RECT 81.955 -68.925 82.095 -68.755 ;
      RECT 81.955 -67.429 82.045 -66.422 ;
      RECT 81.955 -66.905 82.095 -66.735 ;
      RECT 81.955 -66.008 82.045 -65.001 ;
      RECT 81.955 -65.695 82.095 -65.525 ;
      RECT 81.955 -64.199 82.045 -63.192 ;
      RECT 81.955 -63.675 82.095 -63.505 ;
      RECT 81.955 -62.778 82.045 -61.771 ;
      RECT 81.955 -62.465 82.095 -62.295 ;
      RECT 81.955 -60.969 82.045 -59.962 ;
      RECT 81.955 -60.445 82.095 -60.275 ;
      RECT 81.955 -59.548 82.045 -58.541 ;
      RECT 81.955 -59.235 82.095 -59.065 ;
      RECT 81.955 -57.739 82.045 -56.732 ;
      RECT 81.955 -57.215 82.095 -57.045 ;
      RECT 81.955 -56.318 82.045 -55.311 ;
      RECT 81.955 -56.005 82.095 -55.835 ;
      RECT 81.955 -54.509 82.045 -53.502 ;
      RECT 81.955 -53.985 82.095 -53.815 ;
      RECT 81.955 -53.088 82.045 -52.081 ;
      RECT 81.955 -52.775 82.095 -52.605 ;
      RECT 81.955 -51.279 82.045 -50.272 ;
      RECT 81.955 -50.755 82.095 -50.585 ;
      RECT 81.955 -49.858 82.045 -48.851 ;
      RECT 81.955 -49.545 82.095 -49.375 ;
      RECT 81.955 -48.049 82.045 -47.042 ;
      RECT 81.955 -47.525 82.095 -47.355 ;
      RECT 81.955 -46.628 82.045 -45.621 ;
      RECT 81.955 -46.315 82.095 -46.145 ;
      RECT 81.955 -44.819 82.045 -43.812 ;
      RECT 81.955 -44.295 82.095 -44.125 ;
      RECT 81.955 -43.398 82.045 -42.391 ;
      RECT 81.955 -43.085 82.095 -42.915 ;
      RECT 81.955 -41.589 82.045 -40.582 ;
      RECT 81.955 -41.065 82.095 -40.895 ;
      RECT 81.955 -40.168 82.045 -39.161 ;
      RECT 81.955 -39.855 82.095 -39.685 ;
      RECT 81.955 -38.359 82.045 -37.352 ;
      RECT 81.955 -37.835 82.095 -37.665 ;
      RECT 81.955 -36.938 82.045 -35.931 ;
      RECT 81.955 -36.625 82.095 -36.455 ;
      RECT 81.955 -35.129 82.045 -34.122 ;
      RECT 81.955 -34.605 82.095 -34.435 ;
      RECT 81.955 -33.708 82.045 -32.701 ;
      RECT 81.955 -33.395 82.095 -33.225 ;
      RECT 81.955 -31.899 82.045 -30.892 ;
      RECT 81.955 -31.375 82.095 -31.205 ;
      RECT 81.955 -30.478 82.045 -29.471 ;
      RECT 81.955 -30.165 82.095 -29.995 ;
      RECT 81.955 -28.669 82.045 -27.662 ;
      RECT 81.955 -28.145 82.095 -27.975 ;
      RECT 81.955 -27.248 82.045 -26.241 ;
      RECT 81.955 -26.935 82.095 -26.765 ;
      RECT 81.955 -25.439 82.045 -24.432 ;
      RECT 81.955 -24.915 82.095 -24.745 ;
      RECT 81.955 -24.018 82.045 -23.011 ;
      RECT 81.955 -23.705 82.095 -23.535 ;
      RECT 81.955 -22.209 82.045 -21.202 ;
      RECT 81.955 -21.685 82.095 -21.515 ;
      RECT 81.955 -20.788 82.045 -19.781 ;
      RECT 81.955 -20.475 82.095 -20.305 ;
      RECT 81.955 -18.979 82.045 -17.972 ;
      RECT 81.955 -18.455 82.095 -18.285 ;
      RECT 81.955 -17.558 82.045 -16.551 ;
      RECT 81.955 -17.245 82.095 -17.075 ;
      RECT 81.955 -15.749 82.045 -14.742 ;
      RECT 81.955 -15.225 82.095 -15.055 ;
      RECT 81.955 -14.328 82.045 -13.321 ;
      RECT 81.955 -14.015 82.095 -13.845 ;
      RECT 81.955 -12.519 82.045 -11.512 ;
      RECT 81.955 -11.995 82.095 -11.825 ;
      RECT 81.955 -11.098 82.045 -10.091 ;
      RECT 81.955 -10.785 82.095 -10.615 ;
      RECT 81.955 -9.289 82.045 -8.282 ;
      RECT 81.955 -8.765 82.095 -8.595 ;
      RECT 81.955 -7.868 82.045 -6.861 ;
      RECT 81.955 -7.555 82.095 -7.385 ;
      RECT 81.955 -6.059 82.045 -5.052 ;
      RECT 81.955 -5.535 82.095 -5.365 ;
      RECT 81.955 -4.638 82.045 -3.631 ;
      RECT 81.955 -4.325 82.095 -4.155 ;
      RECT 81.955 -2.829 82.045 -1.822 ;
      RECT 81.955 -2.305 82.095 -2.135 ;
      RECT 81.955 -1.408 82.045 -0.401 ;
      RECT 81.955 -1.095 82.095 -0.925 ;
      RECT 81.955 0.401 82.045 1.408 ;
      RECT 81.955 0.925 82.095 1.095 ;
      RECT 77.785 -108.935 81.565 -108.815 ;
      RECT 79.105 -109.475 79.205 -108.815 ;
      RECT 78.545 -109.475 78.645 -108.815 ;
      RECT 77.985 -109.475 78.085 -108.815 ;
      RECT 81.155 -101.538 81.245 -100.53 ;
      RECT 81.105 -100.935 81.245 -100.765 ;
      RECT 81.155 -99.73 81.245 -98.722 ;
      RECT 81.105 -99.495 81.245 -99.325 ;
      RECT 81.155 -98.308 81.245 -97.3 ;
      RECT 81.105 -97.705 81.245 -97.535 ;
      RECT 81.155 -96.5 81.245 -95.492 ;
      RECT 81.105 -96.265 81.245 -96.095 ;
      RECT 81.155 -95.078 81.245 -94.07 ;
      RECT 81.105 -94.475 81.245 -94.305 ;
      RECT 81.155 -93.27 81.245 -92.262 ;
      RECT 81.105 -93.035 81.245 -92.865 ;
      RECT 81.155 -91.848 81.245 -90.84 ;
      RECT 81.105 -91.245 81.245 -91.075 ;
      RECT 81.155 -90.04 81.245 -89.032 ;
      RECT 81.105 -89.805 81.245 -89.635 ;
      RECT 81.155 -88.618 81.245 -87.61 ;
      RECT 81.105 -88.015 81.245 -87.845 ;
      RECT 81.155 -86.81 81.245 -85.802 ;
      RECT 81.105 -86.575 81.245 -86.405 ;
      RECT 81.155 -85.388 81.245 -84.38 ;
      RECT 81.105 -84.785 81.245 -84.615 ;
      RECT 81.155 -83.58 81.245 -82.572 ;
      RECT 81.105 -83.345 81.245 -83.175 ;
      RECT 81.155 -82.158 81.245 -81.15 ;
      RECT 81.105 -81.555 81.245 -81.385 ;
      RECT 81.155 -80.35 81.245 -79.342 ;
      RECT 81.105 -80.115 81.245 -79.945 ;
      RECT 81.155 -78.928 81.245 -77.92 ;
      RECT 81.105 -78.325 81.245 -78.155 ;
      RECT 81.155 -77.12 81.245 -76.112 ;
      RECT 81.105 -76.885 81.245 -76.715 ;
      RECT 81.155 -75.698 81.245 -74.69 ;
      RECT 81.105 -75.095 81.245 -74.925 ;
      RECT 81.155 -73.89 81.245 -72.882 ;
      RECT 81.105 -73.655 81.245 -73.485 ;
      RECT 81.155 -72.468 81.245 -71.46 ;
      RECT 81.105 -71.865 81.245 -71.695 ;
      RECT 81.155 -70.66 81.245 -69.652 ;
      RECT 81.105 -70.425 81.245 -70.255 ;
      RECT 81.155 -69.238 81.245 -68.23 ;
      RECT 81.105 -68.635 81.245 -68.465 ;
      RECT 81.155 -67.43 81.245 -66.422 ;
      RECT 81.105 -67.195 81.245 -67.025 ;
      RECT 81.155 -66.008 81.245 -65 ;
      RECT 81.105 -65.405 81.245 -65.235 ;
      RECT 81.155 -64.2 81.245 -63.192 ;
      RECT 81.105 -63.965 81.245 -63.795 ;
      RECT 81.155 -62.778 81.245 -61.77 ;
      RECT 81.105 -62.175 81.245 -62.005 ;
      RECT 81.155 -60.97 81.245 -59.962 ;
      RECT 81.105 -60.735 81.245 -60.565 ;
      RECT 81.155 -59.548 81.245 -58.54 ;
      RECT 81.105 -58.945 81.245 -58.775 ;
      RECT 81.155 -57.74 81.245 -56.732 ;
      RECT 81.105 -57.505 81.245 -57.335 ;
      RECT 81.155 -56.318 81.245 -55.31 ;
      RECT 81.105 -55.715 81.245 -55.545 ;
      RECT 81.155 -54.51 81.245 -53.502 ;
      RECT 81.105 -54.275 81.245 -54.105 ;
      RECT 81.155 -53.088 81.245 -52.08 ;
      RECT 81.105 -52.485 81.245 -52.315 ;
      RECT 81.155 -51.28 81.245 -50.272 ;
      RECT 81.105 -51.045 81.245 -50.875 ;
      RECT 81.155 -49.858 81.245 -48.85 ;
      RECT 81.105 -49.255 81.245 -49.085 ;
      RECT 81.155 -48.05 81.245 -47.042 ;
      RECT 81.105 -47.815 81.245 -47.645 ;
      RECT 81.155 -46.628 81.245 -45.62 ;
      RECT 81.105 -46.025 81.245 -45.855 ;
      RECT 81.155 -44.82 81.245 -43.812 ;
      RECT 81.105 -44.585 81.245 -44.415 ;
      RECT 81.155 -43.398 81.245 -42.39 ;
      RECT 81.105 -42.795 81.245 -42.625 ;
      RECT 81.155 -41.59 81.245 -40.582 ;
      RECT 81.105 -41.355 81.245 -41.185 ;
      RECT 81.155 -40.168 81.245 -39.16 ;
      RECT 81.105 -39.565 81.245 -39.395 ;
      RECT 81.155 -38.36 81.245 -37.352 ;
      RECT 81.105 -38.125 81.245 -37.955 ;
      RECT 81.155 -36.938 81.245 -35.93 ;
      RECT 81.105 -36.335 81.245 -36.165 ;
      RECT 81.155 -35.13 81.245 -34.122 ;
      RECT 81.105 -34.895 81.245 -34.725 ;
      RECT 81.155 -33.708 81.245 -32.7 ;
      RECT 81.105 -33.105 81.245 -32.935 ;
      RECT 81.155 -31.9 81.245 -30.892 ;
      RECT 81.105 -31.665 81.245 -31.495 ;
      RECT 81.155 -30.478 81.245 -29.47 ;
      RECT 81.105 -29.875 81.245 -29.705 ;
      RECT 81.155 -28.67 81.245 -27.662 ;
      RECT 81.105 -28.435 81.245 -28.265 ;
      RECT 81.155 -27.248 81.245 -26.24 ;
      RECT 81.105 -26.645 81.245 -26.475 ;
      RECT 81.155 -25.44 81.245 -24.432 ;
      RECT 81.105 -25.205 81.245 -25.035 ;
      RECT 81.155 -24.018 81.245 -23.01 ;
      RECT 81.105 -23.415 81.245 -23.245 ;
      RECT 81.155 -22.21 81.245 -21.202 ;
      RECT 81.105 -21.975 81.245 -21.805 ;
      RECT 81.155 -20.788 81.245 -19.78 ;
      RECT 81.105 -20.185 81.245 -20.015 ;
      RECT 81.155 -18.98 81.245 -17.972 ;
      RECT 81.105 -18.745 81.245 -18.575 ;
      RECT 81.155 -17.558 81.245 -16.55 ;
      RECT 81.105 -16.955 81.245 -16.785 ;
      RECT 81.155 -15.75 81.245 -14.742 ;
      RECT 81.105 -15.515 81.245 -15.345 ;
      RECT 81.155 -14.328 81.245 -13.32 ;
      RECT 81.105 -13.725 81.245 -13.555 ;
      RECT 81.155 -12.52 81.245 -11.512 ;
      RECT 81.105 -12.285 81.245 -12.115 ;
      RECT 81.155 -11.098 81.245 -10.09 ;
      RECT 81.105 -10.495 81.245 -10.325 ;
      RECT 81.155 -9.29 81.245 -8.282 ;
      RECT 81.105 -9.055 81.245 -8.885 ;
      RECT 81.155 -7.868 81.245 -6.86 ;
      RECT 81.105 -7.265 81.245 -7.095 ;
      RECT 81.155 -6.06 81.245 -5.052 ;
      RECT 81.105 -5.825 81.245 -5.655 ;
      RECT 81.155 -4.638 81.245 -3.63 ;
      RECT 81.105 -4.035 81.245 -3.865 ;
      RECT 81.155 -2.83 81.245 -1.822 ;
      RECT 81.105 -2.595 81.245 -2.425 ;
      RECT 81.155 -1.408 81.245 -0.4 ;
      RECT 81.105 -0.805 81.245 -0.635 ;
      RECT 81.155 0.4 81.245 1.408 ;
      RECT 81.105 0.635 81.245 0.805 ;
      RECT 79.725 -111.685 81.205 -111.585 ;
      RECT 79.725 -112.195 79.825 -111.585 ;
      RECT 79.945 -109.15 81.205 -109.05 ;
      RECT 81.105 -109.475 81.205 -109.05 ;
      RECT 80.545 -109.475 80.645 -109.05 ;
      RECT 79.985 -109.475 80.085 -109.05 ;
      RECT 80.755 -101.538 80.845 -100.531 ;
      RECT 80.755 -101.225 80.895 -101.055 ;
      RECT 80.755 -99.729 80.845 -98.722 ;
      RECT 80.755 -99.205 80.895 -99.035 ;
      RECT 80.755 -98.308 80.845 -97.301 ;
      RECT 80.755 -97.995 80.895 -97.825 ;
      RECT 80.755 -96.499 80.845 -95.492 ;
      RECT 80.755 -95.975 80.895 -95.805 ;
      RECT 80.755 -95.078 80.845 -94.071 ;
      RECT 80.755 -94.765 80.895 -94.595 ;
      RECT 80.755 -93.269 80.845 -92.262 ;
      RECT 80.755 -92.745 80.895 -92.575 ;
      RECT 80.755 -91.848 80.845 -90.841 ;
      RECT 80.755 -91.535 80.895 -91.365 ;
      RECT 80.755 -90.039 80.845 -89.032 ;
      RECT 80.755 -89.515 80.895 -89.345 ;
      RECT 80.755 -88.618 80.845 -87.611 ;
      RECT 80.755 -88.305 80.895 -88.135 ;
      RECT 80.755 -86.809 80.845 -85.802 ;
      RECT 80.755 -86.285 80.895 -86.115 ;
      RECT 80.755 -85.388 80.845 -84.381 ;
      RECT 80.755 -85.075 80.895 -84.905 ;
      RECT 80.755 -83.579 80.845 -82.572 ;
      RECT 80.755 -83.055 80.895 -82.885 ;
      RECT 80.755 -82.158 80.845 -81.151 ;
      RECT 80.755 -81.845 80.895 -81.675 ;
      RECT 80.755 -80.349 80.845 -79.342 ;
      RECT 80.755 -79.825 80.895 -79.655 ;
      RECT 80.755 -78.928 80.845 -77.921 ;
      RECT 80.755 -78.615 80.895 -78.445 ;
      RECT 80.755 -77.119 80.845 -76.112 ;
      RECT 80.755 -76.595 80.895 -76.425 ;
      RECT 80.755 -75.698 80.845 -74.691 ;
      RECT 80.755 -75.385 80.895 -75.215 ;
      RECT 80.755 -73.889 80.845 -72.882 ;
      RECT 80.755 -73.365 80.895 -73.195 ;
      RECT 80.755 -72.468 80.845 -71.461 ;
      RECT 80.755 -72.155 80.895 -71.985 ;
      RECT 80.755 -70.659 80.845 -69.652 ;
      RECT 80.755 -70.135 80.895 -69.965 ;
      RECT 80.755 -69.238 80.845 -68.231 ;
      RECT 80.755 -68.925 80.895 -68.755 ;
      RECT 80.755 -67.429 80.845 -66.422 ;
      RECT 80.755 -66.905 80.895 -66.735 ;
      RECT 80.755 -66.008 80.845 -65.001 ;
      RECT 80.755 -65.695 80.895 -65.525 ;
      RECT 80.755 -64.199 80.845 -63.192 ;
      RECT 80.755 -63.675 80.895 -63.505 ;
      RECT 80.755 -62.778 80.845 -61.771 ;
      RECT 80.755 -62.465 80.895 -62.295 ;
      RECT 80.755 -60.969 80.845 -59.962 ;
      RECT 80.755 -60.445 80.895 -60.275 ;
      RECT 80.755 -59.548 80.845 -58.541 ;
      RECT 80.755 -59.235 80.895 -59.065 ;
      RECT 80.755 -57.739 80.845 -56.732 ;
      RECT 80.755 -57.215 80.895 -57.045 ;
      RECT 80.755 -56.318 80.845 -55.311 ;
      RECT 80.755 -56.005 80.895 -55.835 ;
      RECT 80.755 -54.509 80.845 -53.502 ;
      RECT 80.755 -53.985 80.895 -53.815 ;
      RECT 80.755 -53.088 80.845 -52.081 ;
      RECT 80.755 -52.775 80.895 -52.605 ;
      RECT 80.755 -51.279 80.845 -50.272 ;
      RECT 80.755 -50.755 80.895 -50.585 ;
      RECT 80.755 -49.858 80.845 -48.851 ;
      RECT 80.755 -49.545 80.895 -49.375 ;
      RECT 80.755 -48.049 80.845 -47.042 ;
      RECT 80.755 -47.525 80.895 -47.355 ;
      RECT 80.755 -46.628 80.845 -45.621 ;
      RECT 80.755 -46.315 80.895 -46.145 ;
      RECT 80.755 -44.819 80.845 -43.812 ;
      RECT 80.755 -44.295 80.895 -44.125 ;
      RECT 80.755 -43.398 80.845 -42.391 ;
      RECT 80.755 -43.085 80.895 -42.915 ;
      RECT 80.755 -41.589 80.845 -40.582 ;
      RECT 80.755 -41.065 80.895 -40.895 ;
      RECT 80.755 -40.168 80.845 -39.161 ;
      RECT 80.755 -39.855 80.895 -39.685 ;
      RECT 80.755 -38.359 80.845 -37.352 ;
      RECT 80.755 -37.835 80.895 -37.665 ;
      RECT 80.755 -36.938 80.845 -35.931 ;
      RECT 80.755 -36.625 80.895 -36.455 ;
      RECT 80.755 -35.129 80.845 -34.122 ;
      RECT 80.755 -34.605 80.895 -34.435 ;
      RECT 80.755 -33.708 80.845 -32.701 ;
      RECT 80.755 -33.395 80.895 -33.225 ;
      RECT 80.755 -31.899 80.845 -30.892 ;
      RECT 80.755 -31.375 80.895 -31.205 ;
      RECT 80.755 -30.478 80.845 -29.471 ;
      RECT 80.755 -30.165 80.895 -29.995 ;
      RECT 80.755 -28.669 80.845 -27.662 ;
      RECT 80.755 -28.145 80.895 -27.975 ;
      RECT 80.755 -27.248 80.845 -26.241 ;
      RECT 80.755 -26.935 80.895 -26.765 ;
      RECT 80.755 -25.439 80.845 -24.432 ;
      RECT 80.755 -24.915 80.895 -24.745 ;
      RECT 80.755 -24.018 80.845 -23.011 ;
      RECT 80.755 -23.705 80.895 -23.535 ;
      RECT 80.755 -22.209 80.845 -21.202 ;
      RECT 80.755 -21.685 80.895 -21.515 ;
      RECT 80.755 -20.788 80.845 -19.781 ;
      RECT 80.755 -20.475 80.895 -20.305 ;
      RECT 80.755 -18.979 80.845 -17.972 ;
      RECT 80.755 -18.455 80.895 -18.285 ;
      RECT 80.755 -17.558 80.845 -16.551 ;
      RECT 80.755 -17.245 80.895 -17.075 ;
      RECT 80.755 -15.749 80.845 -14.742 ;
      RECT 80.755 -15.225 80.895 -15.055 ;
      RECT 80.755 -14.328 80.845 -13.321 ;
      RECT 80.755 -14.015 80.895 -13.845 ;
      RECT 80.755 -12.519 80.845 -11.512 ;
      RECT 80.755 -11.995 80.895 -11.825 ;
      RECT 80.755 -11.098 80.845 -10.091 ;
      RECT 80.755 -10.785 80.895 -10.615 ;
      RECT 80.755 -9.289 80.845 -8.282 ;
      RECT 80.755 -8.765 80.895 -8.595 ;
      RECT 80.755 -7.868 80.845 -6.861 ;
      RECT 80.755 -7.555 80.895 -7.385 ;
      RECT 80.755 -6.059 80.845 -5.052 ;
      RECT 80.755 -5.535 80.895 -5.365 ;
      RECT 80.755 -4.638 80.845 -3.631 ;
      RECT 80.755 -4.325 80.895 -4.155 ;
      RECT 80.755 -2.829 80.845 -1.822 ;
      RECT 80.755 -2.305 80.895 -2.135 ;
      RECT 80.755 -1.408 80.845 -0.401 ;
      RECT 80.755 -1.095 80.895 -0.925 ;
      RECT 80.755 0.401 80.845 1.408 ;
      RECT 80.755 0.925 80.895 1.095 ;
      RECT 80.085 -111.495 80.255 -111.385 ;
      RECT 76.935 -111.495 80.255 -111.395 ;
      RECT 79.955 -101.538 80.045 -100.53 ;
      RECT 79.905 -100.935 80.045 -100.765 ;
      RECT 79.955 -99.73 80.045 -98.722 ;
      RECT 79.905 -99.495 80.045 -99.325 ;
      RECT 79.955 -98.308 80.045 -97.3 ;
      RECT 79.905 -97.705 80.045 -97.535 ;
      RECT 79.955 -96.5 80.045 -95.492 ;
      RECT 79.905 -96.265 80.045 -96.095 ;
      RECT 79.955 -95.078 80.045 -94.07 ;
      RECT 79.905 -94.475 80.045 -94.305 ;
      RECT 79.955 -93.27 80.045 -92.262 ;
      RECT 79.905 -93.035 80.045 -92.865 ;
      RECT 79.955 -91.848 80.045 -90.84 ;
      RECT 79.905 -91.245 80.045 -91.075 ;
      RECT 79.955 -90.04 80.045 -89.032 ;
      RECT 79.905 -89.805 80.045 -89.635 ;
      RECT 79.955 -88.618 80.045 -87.61 ;
      RECT 79.905 -88.015 80.045 -87.845 ;
      RECT 79.955 -86.81 80.045 -85.802 ;
      RECT 79.905 -86.575 80.045 -86.405 ;
      RECT 79.955 -85.388 80.045 -84.38 ;
      RECT 79.905 -84.785 80.045 -84.615 ;
      RECT 79.955 -83.58 80.045 -82.572 ;
      RECT 79.905 -83.345 80.045 -83.175 ;
      RECT 79.955 -82.158 80.045 -81.15 ;
      RECT 79.905 -81.555 80.045 -81.385 ;
      RECT 79.955 -80.35 80.045 -79.342 ;
      RECT 79.905 -80.115 80.045 -79.945 ;
      RECT 79.955 -78.928 80.045 -77.92 ;
      RECT 79.905 -78.325 80.045 -78.155 ;
      RECT 79.955 -77.12 80.045 -76.112 ;
      RECT 79.905 -76.885 80.045 -76.715 ;
      RECT 79.955 -75.698 80.045 -74.69 ;
      RECT 79.905 -75.095 80.045 -74.925 ;
      RECT 79.955 -73.89 80.045 -72.882 ;
      RECT 79.905 -73.655 80.045 -73.485 ;
      RECT 79.955 -72.468 80.045 -71.46 ;
      RECT 79.905 -71.865 80.045 -71.695 ;
      RECT 79.955 -70.66 80.045 -69.652 ;
      RECT 79.905 -70.425 80.045 -70.255 ;
      RECT 79.955 -69.238 80.045 -68.23 ;
      RECT 79.905 -68.635 80.045 -68.465 ;
      RECT 79.955 -67.43 80.045 -66.422 ;
      RECT 79.905 -67.195 80.045 -67.025 ;
      RECT 79.955 -66.008 80.045 -65 ;
      RECT 79.905 -65.405 80.045 -65.235 ;
      RECT 79.955 -64.2 80.045 -63.192 ;
      RECT 79.905 -63.965 80.045 -63.795 ;
      RECT 79.955 -62.778 80.045 -61.77 ;
      RECT 79.905 -62.175 80.045 -62.005 ;
      RECT 79.955 -60.97 80.045 -59.962 ;
      RECT 79.905 -60.735 80.045 -60.565 ;
      RECT 79.955 -59.548 80.045 -58.54 ;
      RECT 79.905 -58.945 80.045 -58.775 ;
      RECT 79.955 -57.74 80.045 -56.732 ;
      RECT 79.905 -57.505 80.045 -57.335 ;
      RECT 79.955 -56.318 80.045 -55.31 ;
      RECT 79.905 -55.715 80.045 -55.545 ;
      RECT 79.955 -54.51 80.045 -53.502 ;
      RECT 79.905 -54.275 80.045 -54.105 ;
      RECT 79.955 -53.088 80.045 -52.08 ;
      RECT 79.905 -52.485 80.045 -52.315 ;
      RECT 79.955 -51.28 80.045 -50.272 ;
      RECT 79.905 -51.045 80.045 -50.875 ;
      RECT 79.955 -49.858 80.045 -48.85 ;
      RECT 79.905 -49.255 80.045 -49.085 ;
      RECT 79.955 -48.05 80.045 -47.042 ;
      RECT 79.905 -47.815 80.045 -47.645 ;
      RECT 79.955 -46.628 80.045 -45.62 ;
      RECT 79.905 -46.025 80.045 -45.855 ;
      RECT 79.955 -44.82 80.045 -43.812 ;
      RECT 79.905 -44.585 80.045 -44.415 ;
      RECT 79.955 -43.398 80.045 -42.39 ;
      RECT 79.905 -42.795 80.045 -42.625 ;
      RECT 79.955 -41.59 80.045 -40.582 ;
      RECT 79.905 -41.355 80.045 -41.185 ;
      RECT 79.955 -40.168 80.045 -39.16 ;
      RECT 79.905 -39.565 80.045 -39.395 ;
      RECT 79.955 -38.36 80.045 -37.352 ;
      RECT 79.905 -38.125 80.045 -37.955 ;
      RECT 79.955 -36.938 80.045 -35.93 ;
      RECT 79.905 -36.335 80.045 -36.165 ;
      RECT 79.955 -35.13 80.045 -34.122 ;
      RECT 79.905 -34.895 80.045 -34.725 ;
      RECT 79.955 -33.708 80.045 -32.7 ;
      RECT 79.905 -33.105 80.045 -32.935 ;
      RECT 79.955 -31.9 80.045 -30.892 ;
      RECT 79.905 -31.665 80.045 -31.495 ;
      RECT 79.955 -30.478 80.045 -29.47 ;
      RECT 79.905 -29.875 80.045 -29.705 ;
      RECT 79.955 -28.67 80.045 -27.662 ;
      RECT 79.905 -28.435 80.045 -28.265 ;
      RECT 79.955 -27.248 80.045 -26.24 ;
      RECT 79.905 -26.645 80.045 -26.475 ;
      RECT 79.955 -25.44 80.045 -24.432 ;
      RECT 79.905 -25.205 80.045 -25.035 ;
      RECT 79.955 -24.018 80.045 -23.01 ;
      RECT 79.905 -23.415 80.045 -23.245 ;
      RECT 79.955 -22.21 80.045 -21.202 ;
      RECT 79.905 -21.975 80.045 -21.805 ;
      RECT 79.955 -20.788 80.045 -19.78 ;
      RECT 79.905 -20.185 80.045 -20.015 ;
      RECT 79.955 -18.98 80.045 -17.972 ;
      RECT 79.905 -18.745 80.045 -18.575 ;
      RECT 79.955 -17.558 80.045 -16.55 ;
      RECT 79.905 -16.955 80.045 -16.785 ;
      RECT 79.955 -15.75 80.045 -14.742 ;
      RECT 79.905 -15.515 80.045 -15.345 ;
      RECT 79.955 -14.328 80.045 -13.32 ;
      RECT 79.905 -13.725 80.045 -13.555 ;
      RECT 79.955 -12.52 80.045 -11.512 ;
      RECT 79.905 -12.285 80.045 -12.115 ;
      RECT 79.955 -11.098 80.045 -10.09 ;
      RECT 79.905 -10.495 80.045 -10.325 ;
      RECT 79.955 -9.29 80.045 -8.282 ;
      RECT 79.905 -9.055 80.045 -8.885 ;
      RECT 79.955 -7.868 80.045 -6.86 ;
      RECT 79.905 -7.265 80.045 -7.095 ;
      RECT 79.955 -6.06 80.045 -5.052 ;
      RECT 79.905 -5.825 80.045 -5.655 ;
      RECT 79.955 -4.638 80.045 -3.63 ;
      RECT 79.905 -4.035 80.045 -3.865 ;
      RECT 79.955 -2.83 80.045 -1.822 ;
      RECT 79.905 -2.595 80.045 -2.425 ;
      RECT 79.955 -1.408 80.045 -0.4 ;
      RECT 79.905 -0.805 80.045 -0.635 ;
      RECT 79.955 0.4 80.045 1.408 ;
      RECT 79.905 0.635 80.045 0.805 ;
      RECT 79.555 -101.538 79.645 -100.531 ;
      RECT 79.555 -101.225 79.695 -101.055 ;
      RECT 79.555 -99.729 79.645 -98.722 ;
      RECT 79.555 -99.205 79.695 -99.035 ;
      RECT 79.555 -98.308 79.645 -97.301 ;
      RECT 79.555 -97.995 79.695 -97.825 ;
      RECT 79.555 -96.499 79.645 -95.492 ;
      RECT 79.555 -95.975 79.695 -95.805 ;
      RECT 79.555 -95.078 79.645 -94.071 ;
      RECT 79.555 -94.765 79.695 -94.595 ;
      RECT 79.555 -93.269 79.645 -92.262 ;
      RECT 79.555 -92.745 79.695 -92.575 ;
      RECT 79.555 -91.848 79.645 -90.841 ;
      RECT 79.555 -91.535 79.695 -91.365 ;
      RECT 79.555 -90.039 79.645 -89.032 ;
      RECT 79.555 -89.515 79.695 -89.345 ;
      RECT 79.555 -88.618 79.645 -87.611 ;
      RECT 79.555 -88.305 79.695 -88.135 ;
      RECT 79.555 -86.809 79.645 -85.802 ;
      RECT 79.555 -86.285 79.695 -86.115 ;
      RECT 79.555 -85.388 79.645 -84.381 ;
      RECT 79.555 -85.075 79.695 -84.905 ;
      RECT 79.555 -83.579 79.645 -82.572 ;
      RECT 79.555 -83.055 79.695 -82.885 ;
      RECT 79.555 -82.158 79.645 -81.151 ;
      RECT 79.555 -81.845 79.695 -81.675 ;
      RECT 79.555 -80.349 79.645 -79.342 ;
      RECT 79.555 -79.825 79.695 -79.655 ;
      RECT 79.555 -78.928 79.645 -77.921 ;
      RECT 79.555 -78.615 79.695 -78.445 ;
      RECT 79.555 -77.119 79.645 -76.112 ;
      RECT 79.555 -76.595 79.695 -76.425 ;
      RECT 79.555 -75.698 79.645 -74.691 ;
      RECT 79.555 -75.385 79.695 -75.215 ;
      RECT 79.555 -73.889 79.645 -72.882 ;
      RECT 79.555 -73.365 79.695 -73.195 ;
      RECT 79.555 -72.468 79.645 -71.461 ;
      RECT 79.555 -72.155 79.695 -71.985 ;
      RECT 79.555 -70.659 79.645 -69.652 ;
      RECT 79.555 -70.135 79.695 -69.965 ;
      RECT 79.555 -69.238 79.645 -68.231 ;
      RECT 79.555 -68.925 79.695 -68.755 ;
      RECT 79.555 -67.429 79.645 -66.422 ;
      RECT 79.555 -66.905 79.695 -66.735 ;
      RECT 79.555 -66.008 79.645 -65.001 ;
      RECT 79.555 -65.695 79.695 -65.525 ;
      RECT 79.555 -64.199 79.645 -63.192 ;
      RECT 79.555 -63.675 79.695 -63.505 ;
      RECT 79.555 -62.778 79.645 -61.771 ;
      RECT 79.555 -62.465 79.695 -62.295 ;
      RECT 79.555 -60.969 79.645 -59.962 ;
      RECT 79.555 -60.445 79.695 -60.275 ;
      RECT 79.555 -59.548 79.645 -58.541 ;
      RECT 79.555 -59.235 79.695 -59.065 ;
      RECT 79.555 -57.739 79.645 -56.732 ;
      RECT 79.555 -57.215 79.695 -57.045 ;
      RECT 79.555 -56.318 79.645 -55.311 ;
      RECT 79.555 -56.005 79.695 -55.835 ;
      RECT 79.555 -54.509 79.645 -53.502 ;
      RECT 79.555 -53.985 79.695 -53.815 ;
      RECT 79.555 -53.088 79.645 -52.081 ;
      RECT 79.555 -52.775 79.695 -52.605 ;
      RECT 79.555 -51.279 79.645 -50.272 ;
      RECT 79.555 -50.755 79.695 -50.585 ;
      RECT 79.555 -49.858 79.645 -48.851 ;
      RECT 79.555 -49.545 79.695 -49.375 ;
      RECT 79.555 -48.049 79.645 -47.042 ;
      RECT 79.555 -47.525 79.695 -47.355 ;
      RECT 79.555 -46.628 79.645 -45.621 ;
      RECT 79.555 -46.315 79.695 -46.145 ;
      RECT 79.555 -44.819 79.645 -43.812 ;
      RECT 79.555 -44.295 79.695 -44.125 ;
      RECT 79.555 -43.398 79.645 -42.391 ;
      RECT 79.555 -43.085 79.695 -42.915 ;
      RECT 79.555 -41.589 79.645 -40.582 ;
      RECT 79.555 -41.065 79.695 -40.895 ;
      RECT 79.555 -40.168 79.645 -39.161 ;
      RECT 79.555 -39.855 79.695 -39.685 ;
      RECT 79.555 -38.359 79.645 -37.352 ;
      RECT 79.555 -37.835 79.695 -37.665 ;
      RECT 79.555 -36.938 79.645 -35.931 ;
      RECT 79.555 -36.625 79.695 -36.455 ;
      RECT 79.555 -35.129 79.645 -34.122 ;
      RECT 79.555 -34.605 79.695 -34.435 ;
      RECT 79.555 -33.708 79.645 -32.701 ;
      RECT 79.555 -33.395 79.695 -33.225 ;
      RECT 79.555 -31.899 79.645 -30.892 ;
      RECT 79.555 -31.375 79.695 -31.205 ;
      RECT 79.555 -30.478 79.645 -29.471 ;
      RECT 79.555 -30.165 79.695 -29.995 ;
      RECT 79.555 -28.669 79.645 -27.662 ;
      RECT 79.555 -28.145 79.695 -27.975 ;
      RECT 79.555 -27.248 79.645 -26.241 ;
      RECT 79.555 -26.935 79.695 -26.765 ;
      RECT 79.555 -25.439 79.645 -24.432 ;
      RECT 79.555 -24.915 79.695 -24.745 ;
      RECT 79.555 -24.018 79.645 -23.011 ;
      RECT 79.555 -23.705 79.695 -23.535 ;
      RECT 79.555 -22.209 79.645 -21.202 ;
      RECT 79.555 -21.685 79.695 -21.515 ;
      RECT 79.555 -20.788 79.645 -19.781 ;
      RECT 79.555 -20.475 79.695 -20.305 ;
      RECT 79.555 -18.979 79.645 -17.972 ;
      RECT 79.555 -18.455 79.695 -18.285 ;
      RECT 79.555 -17.558 79.645 -16.551 ;
      RECT 79.555 -17.245 79.695 -17.075 ;
      RECT 79.555 -15.749 79.645 -14.742 ;
      RECT 79.555 -15.225 79.695 -15.055 ;
      RECT 79.555 -14.328 79.645 -13.321 ;
      RECT 79.555 -14.015 79.695 -13.845 ;
      RECT 79.555 -12.519 79.645 -11.512 ;
      RECT 79.555 -11.995 79.695 -11.825 ;
      RECT 79.555 -11.098 79.645 -10.091 ;
      RECT 79.555 -10.785 79.695 -10.615 ;
      RECT 79.555 -9.289 79.645 -8.282 ;
      RECT 79.555 -8.765 79.695 -8.595 ;
      RECT 79.555 -7.868 79.645 -6.861 ;
      RECT 79.555 -7.555 79.695 -7.385 ;
      RECT 79.555 -6.059 79.645 -5.052 ;
      RECT 79.555 -5.535 79.695 -5.365 ;
      RECT 79.555 -4.638 79.645 -3.631 ;
      RECT 79.555 -4.325 79.695 -4.155 ;
      RECT 79.555 -2.829 79.645 -1.822 ;
      RECT 79.555 -2.305 79.695 -2.135 ;
      RECT 79.555 -1.408 79.645 -0.401 ;
      RECT 79.555 -1.095 79.695 -0.925 ;
      RECT 79.555 0.401 79.645 1.408 ;
      RECT 79.555 0.925 79.695 1.095 ;
      RECT 77.705 -111.685 79.185 -111.585 ;
      RECT 77.705 -112.055 77.805 -111.585 ;
      RECT 77.51 -114.395 79.085 -114.275 ;
      RECT 78.985 -114.895 79.085 -114.275 ;
      RECT 78.39 -114.895 78.49 -114.275 ;
      RECT 77.51 -114.85 77.61 -114.275 ;
      RECT 78.755 -101.538 78.845 -100.53 ;
      RECT 78.705 -100.935 78.845 -100.765 ;
      RECT 78.755 -99.73 78.845 -98.722 ;
      RECT 78.705 -99.495 78.845 -99.325 ;
      RECT 78.755 -98.308 78.845 -97.3 ;
      RECT 78.705 -97.705 78.845 -97.535 ;
      RECT 78.755 -96.5 78.845 -95.492 ;
      RECT 78.705 -96.265 78.845 -96.095 ;
      RECT 78.755 -95.078 78.845 -94.07 ;
      RECT 78.705 -94.475 78.845 -94.305 ;
      RECT 78.755 -93.27 78.845 -92.262 ;
      RECT 78.705 -93.035 78.845 -92.865 ;
      RECT 78.755 -91.848 78.845 -90.84 ;
      RECT 78.705 -91.245 78.845 -91.075 ;
      RECT 78.755 -90.04 78.845 -89.032 ;
      RECT 78.705 -89.805 78.845 -89.635 ;
      RECT 78.755 -88.618 78.845 -87.61 ;
      RECT 78.705 -88.015 78.845 -87.845 ;
      RECT 78.755 -86.81 78.845 -85.802 ;
      RECT 78.705 -86.575 78.845 -86.405 ;
      RECT 78.755 -85.388 78.845 -84.38 ;
      RECT 78.705 -84.785 78.845 -84.615 ;
      RECT 78.755 -83.58 78.845 -82.572 ;
      RECT 78.705 -83.345 78.845 -83.175 ;
      RECT 78.755 -82.158 78.845 -81.15 ;
      RECT 78.705 -81.555 78.845 -81.385 ;
      RECT 78.755 -80.35 78.845 -79.342 ;
      RECT 78.705 -80.115 78.845 -79.945 ;
      RECT 78.755 -78.928 78.845 -77.92 ;
      RECT 78.705 -78.325 78.845 -78.155 ;
      RECT 78.755 -77.12 78.845 -76.112 ;
      RECT 78.705 -76.885 78.845 -76.715 ;
      RECT 78.755 -75.698 78.845 -74.69 ;
      RECT 78.705 -75.095 78.845 -74.925 ;
      RECT 78.755 -73.89 78.845 -72.882 ;
      RECT 78.705 -73.655 78.845 -73.485 ;
      RECT 78.755 -72.468 78.845 -71.46 ;
      RECT 78.705 -71.865 78.845 -71.695 ;
      RECT 78.755 -70.66 78.845 -69.652 ;
      RECT 78.705 -70.425 78.845 -70.255 ;
      RECT 78.755 -69.238 78.845 -68.23 ;
      RECT 78.705 -68.635 78.845 -68.465 ;
      RECT 78.755 -67.43 78.845 -66.422 ;
      RECT 78.705 -67.195 78.845 -67.025 ;
      RECT 78.755 -66.008 78.845 -65 ;
      RECT 78.705 -65.405 78.845 -65.235 ;
      RECT 78.755 -64.2 78.845 -63.192 ;
      RECT 78.705 -63.965 78.845 -63.795 ;
      RECT 78.755 -62.778 78.845 -61.77 ;
      RECT 78.705 -62.175 78.845 -62.005 ;
      RECT 78.755 -60.97 78.845 -59.962 ;
      RECT 78.705 -60.735 78.845 -60.565 ;
      RECT 78.755 -59.548 78.845 -58.54 ;
      RECT 78.705 -58.945 78.845 -58.775 ;
      RECT 78.755 -57.74 78.845 -56.732 ;
      RECT 78.705 -57.505 78.845 -57.335 ;
      RECT 78.755 -56.318 78.845 -55.31 ;
      RECT 78.705 -55.715 78.845 -55.545 ;
      RECT 78.755 -54.51 78.845 -53.502 ;
      RECT 78.705 -54.275 78.845 -54.105 ;
      RECT 78.755 -53.088 78.845 -52.08 ;
      RECT 78.705 -52.485 78.845 -52.315 ;
      RECT 78.755 -51.28 78.845 -50.272 ;
      RECT 78.705 -51.045 78.845 -50.875 ;
      RECT 78.755 -49.858 78.845 -48.85 ;
      RECT 78.705 -49.255 78.845 -49.085 ;
      RECT 78.755 -48.05 78.845 -47.042 ;
      RECT 78.705 -47.815 78.845 -47.645 ;
      RECT 78.755 -46.628 78.845 -45.62 ;
      RECT 78.705 -46.025 78.845 -45.855 ;
      RECT 78.755 -44.82 78.845 -43.812 ;
      RECT 78.705 -44.585 78.845 -44.415 ;
      RECT 78.755 -43.398 78.845 -42.39 ;
      RECT 78.705 -42.795 78.845 -42.625 ;
      RECT 78.755 -41.59 78.845 -40.582 ;
      RECT 78.705 -41.355 78.845 -41.185 ;
      RECT 78.755 -40.168 78.845 -39.16 ;
      RECT 78.705 -39.565 78.845 -39.395 ;
      RECT 78.755 -38.36 78.845 -37.352 ;
      RECT 78.705 -38.125 78.845 -37.955 ;
      RECT 78.755 -36.938 78.845 -35.93 ;
      RECT 78.705 -36.335 78.845 -36.165 ;
      RECT 78.755 -35.13 78.845 -34.122 ;
      RECT 78.705 -34.895 78.845 -34.725 ;
      RECT 78.755 -33.708 78.845 -32.7 ;
      RECT 78.705 -33.105 78.845 -32.935 ;
      RECT 78.755 -31.9 78.845 -30.892 ;
      RECT 78.705 -31.665 78.845 -31.495 ;
      RECT 78.755 -30.478 78.845 -29.47 ;
      RECT 78.705 -29.875 78.845 -29.705 ;
      RECT 78.755 -28.67 78.845 -27.662 ;
      RECT 78.705 -28.435 78.845 -28.265 ;
      RECT 78.755 -27.248 78.845 -26.24 ;
      RECT 78.705 -26.645 78.845 -26.475 ;
      RECT 78.755 -25.44 78.845 -24.432 ;
      RECT 78.705 -25.205 78.845 -25.035 ;
      RECT 78.755 -24.018 78.845 -23.01 ;
      RECT 78.705 -23.415 78.845 -23.245 ;
      RECT 78.755 -22.21 78.845 -21.202 ;
      RECT 78.705 -21.975 78.845 -21.805 ;
      RECT 78.755 -20.788 78.845 -19.78 ;
      RECT 78.705 -20.185 78.845 -20.015 ;
      RECT 78.755 -18.98 78.845 -17.972 ;
      RECT 78.705 -18.745 78.845 -18.575 ;
      RECT 78.755 -17.558 78.845 -16.55 ;
      RECT 78.705 -16.955 78.845 -16.785 ;
      RECT 78.755 -15.75 78.845 -14.742 ;
      RECT 78.705 -15.515 78.845 -15.345 ;
      RECT 78.755 -14.328 78.845 -13.32 ;
      RECT 78.705 -13.725 78.845 -13.555 ;
      RECT 78.755 -12.52 78.845 -11.512 ;
      RECT 78.705 -12.285 78.845 -12.115 ;
      RECT 78.755 -11.098 78.845 -10.09 ;
      RECT 78.705 -10.495 78.845 -10.325 ;
      RECT 78.755 -9.29 78.845 -8.282 ;
      RECT 78.705 -9.055 78.845 -8.885 ;
      RECT 78.755 -7.868 78.845 -6.86 ;
      RECT 78.705 -7.265 78.845 -7.095 ;
      RECT 78.755 -6.06 78.845 -5.052 ;
      RECT 78.705 -5.825 78.845 -5.655 ;
      RECT 78.755 -4.638 78.845 -3.63 ;
      RECT 78.705 -4.035 78.845 -3.865 ;
      RECT 78.755 -2.83 78.845 -1.822 ;
      RECT 78.705 -2.595 78.845 -2.425 ;
      RECT 78.755 -1.408 78.845 -0.4 ;
      RECT 78.705 -0.805 78.845 -0.635 ;
      RECT 78.755 0.4 78.845 1.408 ;
      RECT 78.705 0.635 78.845 0.805 ;
      RECT 78.63 -114.685 78.805 -114.515 ;
      RECT 78.705 -114.895 78.805 -114.515 ;
      RECT 77.745 -113.555 77.845 -113.09 ;
      RECT 78.11 -113.555 78.21 -113.1 ;
      RECT 77.745 -113.555 78.59 -113.385 ;
      RECT 78.355 -101.538 78.445 -100.531 ;
      RECT 78.355 -101.225 78.495 -101.055 ;
      RECT 78.355 -99.729 78.445 -98.722 ;
      RECT 78.355 -99.205 78.495 -99.035 ;
      RECT 78.355 -98.308 78.445 -97.301 ;
      RECT 78.355 -97.995 78.495 -97.825 ;
      RECT 78.355 -96.499 78.445 -95.492 ;
      RECT 78.355 -95.975 78.495 -95.805 ;
      RECT 78.355 -95.078 78.445 -94.071 ;
      RECT 78.355 -94.765 78.495 -94.595 ;
      RECT 78.355 -93.269 78.445 -92.262 ;
      RECT 78.355 -92.745 78.495 -92.575 ;
      RECT 78.355 -91.848 78.445 -90.841 ;
      RECT 78.355 -91.535 78.495 -91.365 ;
      RECT 78.355 -90.039 78.445 -89.032 ;
      RECT 78.355 -89.515 78.495 -89.345 ;
      RECT 78.355 -88.618 78.445 -87.611 ;
      RECT 78.355 -88.305 78.495 -88.135 ;
      RECT 78.355 -86.809 78.445 -85.802 ;
      RECT 78.355 -86.285 78.495 -86.115 ;
      RECT 78.355 -85.388 78.445 -84.381 ;
      RECT 78.355 -85.075 78.495 -84.905 ;
      RECT 78.355 -83.579 78.445 -82.572 ;
      RECT 78.355 -83.055 78.495 -82.885 ;
      RECT 78.355 -82.158 78.445 -81.151 ;
      RECT 78.355 -81.845 78.495 -81.675 ;
      RECT 78.355 -80.349 78.445 -79.342 ;
      RECT 78.355 -79.825 78.495 -79.655 ;
      RECT 78.355 -78.928 78.445 -77.921 ;
      RECT 78.355 -78.615 78.495 -78.445 ;
      RECT 78.355 -77.119 78.445 -76.112 ;
      RECT 78.355 -76.595 78.495 -76.425 ;
      RECT 78.355 -75.698 78.445 -74.691 ;
      RECT 78.355 -75.385 78.495 -75.215 ;
      RECT 78.355 -73.889 78.445 -72.882 ;
      RECT 78.355 -73.365 78.495 -73.195 ;
      RECT 78.355 -72.468 78.445 -71.461 ;
      RECT 78.355 -72.155 78.495 -71.985 ;
      RECT 78.355 -70.659 78.445 -69.652 ;
      RECT 78.355 -70.135 78.495 -69.965 ;
      RECT 78.355 -69.238 78.445 -68.231 ;
      RECT 78.355 -68.925 78.495 -68.755 ;
      RECT 78.355 -67.429 78.445 -66.422 ;
      RECT 78.355 -66.905 78.495 -66.735 ;
      RECT 78.355 -66.008 78.445 -65.001 ;
      RECT 78.355 -65.695 78.495 -65.525 ;
      RECT 78.355 -64.199 78.445 -63.192 ;
      RECT 78.355 -63.675 78.495 -63.505 ;
      RECT 78.355 -62.778 78.445 -61.771 ;
      RECT 78.355 -62.465 78.495 -62.295 ;
      RECT 78.355 -60.969 78.445 -59.962 ;
      RECT 78.355 -60.445 78.495 -60.275 ;
      RECT 78.355 -59.548 78.445 -58.541 ;
      RECT 78.355 -59.235 78.495 -59.065 ;
      RECT 78.355 -57.739 78.445 -56.732 ;
      RECT 78.355 -57.215 78.495 -57.045 ;
      RECT 78.355 -56.318 78.445 -55.311 ;
      RECT 78.355 -56.005 78.495 -55.835 ;
      RECT 78.355 -54.509 78.445 -53.502 ;
      RECT 78.355 -53.985 78.495 -53.815 ;
      RECT 78.355 -53.088 78.445 -52.081 ;
      RECT 78.355 -52.775 78.495 -52.605 ;
      RECT 78.355 -51.279 78.445 -50.272 ;
      RECT 78.355 -50.755 78.495 -50.585 ;
      RECT 78.355 -49.858 78.445 -48.851 ;
      RECT 78.355 -49.545 78.495 -49.375 ;
      RECT 78.355 -48.049 78.445 -47.042 ;
      RECT 78.355 -47.525 78.495 -47.355 ;
      RECT 78.355 -46.628 78.445 -45.621 ;
      RECT 78.355 -46.315 78.495 -46.145 ;
      RECT 78.355 -44.819 78.445 -43.812 ;
      RECT 78.355 -44.295 78.495 -44.125 ;
      RECT 78.355 -43.398 78.445 -42.391 ;
      RECT 78.355 -43.085 78.495 -42.915 ;
      RECT 78.355 -41.589 78.445 -40.582 ;
      RECT 78.355 -41.065 78.495 -40.895 ;
      RECT 78.355 -40.168 78.445 -39.161 ;
      RECT 78.355 -39.855 78.495 -39.685 ;
      RECT 78.355 -38.359 78.445 -37.352 ;
      RECT 78.355 -37.835 78.495 -37.665 ;
      RECT 78.355 -36.938 78.445 -35.931 ;
      RECT 78.355 -36.625 78.495 -36.455 ;
      RECT 78.355 -35.129 78.445 -34.122 ;
      RECT 78.355 -34.605 78.495 -34.435 ;
      RECT 78.355 -33.708 78.445 -32.701 ;
      RECT 78.355 -33.395 78.495 -33.225 ;
      RECT 78.355 -31.899 78.445 -30.892 ;
      RECT 78.355 -31.375 78.495 -31.205 ;
      RECT 78.355 -30.478 78.445 -29.471 ;
      RECT 78.355 -30.165 78.495 -29.995 ;
      RECT 78.355 -28.669 78.445 -27.662 ;
      RECT 78.355 -28.145 78.495 -27.975 ;
      RECT 78.355 -27.248 78.445 -26.241 ;
      RECT 78.355 -26.935 78.495 -26.765 ;
      RECT 78.355 -25.439 78.445 -24.432 ;
      RECT 78.355 -24.915 78.495 -24.745 ;
      RECT 78.355 -24.018 78.445 -23.011 ;
      RECT 78.355 -23.705 78.495 -23.535 ;
      RECT 78.355 -22.209 78.445 -21.202 ;
      RECT 78.355 -21.685 78.495 -21.515 ;
      RECT 78.355 -20.788 78.445 -19.781 ;
      RECT 78.355 -20.475 78.495 -20.305 ;
      RECT 78.355 -18.979 78.445 -17.972 ;
      RECT 78.355 -18.455 78.495 -18.285 ;
      RECT 78.355 -17.558 78.445 -16.551 ;
      RECT 78.355 -17.245 78.495 -17.075 ;
      RECT 78.355 -15.749 78.445 -14.742 ;
      RECT 78.355 -15.225 78.495 -15.055 ;
      RECT 78.355 -14.328 78.445 -13.321 ;
      RECT 78.355 -14.015 78.495 -13.845 ;
      RECT 78.355 -12.519 78.445 -11.512 ;
      RECT 78.355 -11.995 78.495 -11.825 ;
      RECT 78.355 -11.098 78.445 -10.091 ;
      RECT 78.355 -10.785 78.495 -10.615 ;
      RECT 78.355 -9.289 78.445 -8.282 ;
      RECT 78.355 -8.765 78.495 -8.595 ;
      RECT 78.355 -7.868 78.445 -6.861 ;
      RECT 78.355 -7.555 78.495 -7.385 ;
      RECT 78.355 -6.059 78.445 -5.052 ;
      RECT 78.355 -5.535 78.495 -5.365 ;
      RECT 78.355 -4.638 78.445 -3.631 ;
      RECT 78.355 -4.325 78.495 -4.155 ;
      RECT 78.355 -2.829 78.445 -1.822 ;
      RECT 78.355 -2.305 78.495 -2.135 ;
      RECT 78.355 -1.408 78.445 -0.401 ;
      RECT 78.355 -1.095 78.495 -0.925 ;
      RECT 78.355 0.401 78.445 1.408 ;
      RECT 78.355 0.925 78.495 1.095 ;
      RECT 78.04 -114.685 78.21 -114.515 ;
      RECT 78.11 -114.895 78.21 -114.515 ;
      RECT 77.555 -101.538 77.645 -100.53 ;
      RECT 77.505 -100.935 77.645 -100.765 ;
      RECT 77.555 -99.73 77.645 -98.722 ;
      RECT 77.505 -99.495 77.645 -99.325 ;
      RECT 77.555 -98.308 77.645 -97.3 ;
      RECT 77.505 -97.705 77.645 -97.535 ;
      RECT 77.555 -96.5 77.645 -95.492 ;
      RECT 77.505 -96.265 77.645 -96.095 ;
      RECT 77.555 -95.078 77.645 -94.07 ;
      RECT 77.505 -94.475 77.645 -94.305 ;
      RECT 77.555 -93.27 77.645 -92.262 ;
      RECT 77.505 -93.035 77.645 -92.865 ;
      RECT 77.555 -91.848 77.645 -90.84 ;
      RECT 77.505 -91.245 77.645 -91.075 ;
      RECT 77.555 -90.04 77.645 -89.032 ;
      RECT 77.505 -89.805 77.645 -89.635 ;
      RECT 77.555 -88.618 77.645 -87.61 ;
      RECT 77.505 -88.015 77.645 -87.845 ;
      RECT 77.555 -86.81 77.645 -85.802 ;
      RECT 77.505 -86.575 77.645 -86.405 ;
      RECT 77.555 -85.388 77.645 -84.38 ;
      RECT 77.505 -84.785 77.645 -84.615 ;
      RECT 77.555 -83.58 77.645 -82.572 ;
      RECT 77.505 -83.345 77.645 -83.175 ;
      RECT 77.555 -82.158 77.645 -81.15 ;
      RECT 77.505 -81.555 77.645 -81.385 ;
      RECT 77.555 -80.35 77.645 -79.342 ;
      RECT 77.505 -80.115 77.645 -79.945 ;
      RECT 77.555 -78.928 77.645 -77.92 ;
      RECT 77.505 -78.325 77.645 -78.155 ;
      RECT 77.555 -77.12 77.645 -76.112 ;
      RECT 77.505 -76.885 77.645 -76.715 ;
      RECT 77.555 -75.698 77.645 -74.69 ;
      RECT 77.505 -75.095 77.645 -74.925 ;
      RECT 77.555 -73.89 77.645 -72.882 ;
      RECT 77.505 -73.655 77.645 -73.485 ;
      RECT 77.555 -72.468 77.645 -71.46 ;
      RECT 77.505 -71.865 77.645 -71.695 ;
      RECT 77.555 -70.66 77.645 -69.652 ;
      RECT 77.505 -70.425 77.645 -70.255 ;
      RECT 77.555 -69.238 77.645 -68.23 ;
      RECT 77.505 -68.635 77.645 -68.465 ;
      RECT 77.555 -67.43 77.645 -66.422 ;
      RECT 77.505 -67.195 77.645 -67.025 ;
      RECT 77.555 -66.008 77.645 -65 ;
      RECT 77.505 -65.405 77.645 -65.235 ;
      RECT 77.555 -64.2 77.645 -63.192 ;
      RECT 77.505 -63.965 77.645 -63.795 ;
      RECT 77.555 -62.778 77.645 -61.77 ;
      RECT 77.505 -62.175 77.645 -62.005 ;
      RECT 77.555 -60.97 77.645 -59.962 ;
      RECT 77.505 -60.735 77.645 -60.565 ;
      RECT 77.555 -59.548 77.645 -58.54 ;
      RECT 77.505 -58.945 77.645 -58.775 ;
      RECT 77.555 -57.74 77.645 -56.732 ;
      RECT 77.505 -57.505 77.645 -57.335 ;
      RECT 77.555 -56.318 77.645 -55.31 ;
      RECT 77.505 -55.715 77.645 -55.545 ;
      RECT 77.555 -54.51 77.645 -53.502 ;
      RECT 77.505 -54.275 77.645 -54.105 ;
      RECT 77.555 -53.088 77.645 -52.08 ;
      RECT 77.505 -52.485 77.645 -52.315 ;
      RECT 77.555 -51.28 77.645 -50.272 ;
      RECT 77.505 -51.045 77.645 -50.875 ;
      RECT 77.555 -49.858 77.645 -48.85 ;
      RECT 77.505 -49.255 77.645 -49.085 ;
      RECT 77.555 -48.05 77.645 -47.042 ;
      RECT 77.505 -47.815 77.645 -47.645 ;
      RECT 77.555 -46.628 77.645 -45.62 ;
      RECT 77.505 -46.025 77.645 -45.855 ;
      RECT 77.555 -44.82 77.645 -43.812 ;
      RECT 77.505 -44.585 77.645 -44.415 ;
      RECT 77.555 -43.398 77.645 -42.39 ;
      RECT 77.505 -42.795 77.645 -42.625 ;
      RECT 77.555 -41.59 77.645 -40.582 ;
      RECT 77.505 -41.355 77.645 -41.185 ;
      RECT 77.555 -40.168 77.645 -39.16 ;
      RECT 77.505 -39.565 77.645 -39.395 ;
      RECT 77.555 -38.36 77.645 -37.352 ;
      RECT 77.505 -38.125 77.645 -37.955 ;
      RECT 77.555 -36.938 77.645 -35.93 ;
      RECT 77.505 -36.335 77.645 -36.165 ;
      RECT 77.555 -35.13 77.645 -34.122 ;
      RECT 77.505 -34.895 77.645 -34.725 ;
      RECT 77.555 -33.708 77.645 -32.7 ;
      RECT 77.505 -33.105 77.645 -32.935 ;
      RECT 77.555 -31.9 77.645 -30.892 ;
      RECT 77.505 -31.665 77.645 -31.495 ;
      RECT 77.555 -30.478 77.645 -29.47 ;
      RECT 77.505 -29.875 77.645 -29.705 ;
      RECT 77.555 -28.67 77.645 -27.662 ;
      RECT 77.505 -28.435 77.645 -28.265 ;
      RECT 77.555 -27.248 77.645 -26.24 ;
      RECT 77.505 -26.645 77.645 -26.475 ;
      RECT 77.555 -25.44 77.645 -24.432 ;
      RECT 77.505 -25.205 77.645 -25.035 ;
      RECT 77.555 -24.018 77.645 -23.01 ;
      RECT 77.505 -23.415 77.645 -23.245 ;
      RECT 77.555 -22.21 77.645 -21.202 ;
      RECT 77.505 -21.975 77.645 -21.805 ;
      RECT 77.555 -20.788 77.645 -19.78 ;
      RECT 77.505 -20.185 77.645 -20.015 ;
      RECT 77.555 -18.98 77.645 -17.972 ;
      RECT 77.505 -18.745 77.645 -18.575 ;
      RECT 77.555 -17.558 77.645 -16.55 ;
      RECT 77.505 -16.955 77.645 -16.785 ;
      RECT 77.555 -15.75 77.645 -14.742 ;
      RECT 77.505 -15.515 77.645 -15.345 ;
      RECT 77.555 -14.328 77.645 -13.32 ;
      RECT 77.505 -13.725 77.645 -13.555 ;
      RECT 77.555 -12.52 77.645 -11.512 ;
      RECT 77.505 -12.285 77.645 -12.115 ;
      RECT 77.555 -11.098 77.645 -10.09 ;
      RECT 77.505 -10.495 77.645 -10.325 ;
      RECT 77.555 -9.29 77.645 -8.282 ;
      RECT 77.505 -9.055 77.645 -8.885 ;
      RECT 77.555 -7.868 77.645 -6.86 ;
      RECT 77.505 -7.265 77.645 -7.095 ;
      RECT 77.555 -6.06 77.645 -5.052 ;
      RECT 77.505 -5.825 77.645 -5.655 ;
      RECT 77.555 -4.638 77.645 -3.63 ;
      RECT 77.505 -4.035 77.645 -3.865 ;
      RECT 77.555 -2.83 77.645 -1.822 ;
      RECT 77.505 -2.595 77.645 -2.425 ;
      RECT 77.555 -1.408 77.645 -0.4 ;
      RECT 77.505 -0.805 77.645 -0.635 ;
      RECT 77.555 0.4 77.645 1.408 ;
      RECT 77.505 0.635 77.645 0.805 ;
      RECT 77.155 -101.538 77.245 -100.531 ;
      RECT 77.155 -101.225 77.295 -101.055 ;
      RECT 77.155 -99.729 77.245 -98.722 ;
      RECT 77.155 -99.205 77.295 -99.035 ;
      RECT 77.155 -98.308 77.245 -97.301 ;
      RECT 77.155 -97.995 77.295 -97.825 ;
      RECT 77.155 -96.499 77.245 -95.492 ;
      RECT 77.155 -95.975 77.295 -95.805 ;
      RECT 77.155 -95.078 77.245 -94.071 ;
      RECT 77.155 -94.765 77.295 -94.595 ;
      RECT 77.155 -93.269 77.245 -92.262 ;
      RECT 77.155 -92.745 77.295 -92.575 ;
      RECT 77.155 -91.848 77.245 -90.841 ;
      RECT 77.155 -91.535 77.295 -91.365 ;
      RECT 77.155 -90.039 77.245 -89.032 ;
      RECT 77.155 -89.515 77.295 -89.345 ;
      RECT 77.155 -88.618 77.245 -87.611 ;
      RECT 77.155 -88.305 77.295 -88.135 ;
      RECT 77.155 -86.809 77.245 -85.802 ;
      RECT 77.155 -86.285 77.295 -86.115 ;
      RECT 77.155 -85.388 77.245 -84.381 ;
      RECT 77.155 -85.075 77.295 -84.905 ;
      RECT 77.155 -83.579 77.245 -82.572 ;
      RECT 77.155 -83.055 77.295 -82.885 ;
      RECT 77.155 -82.158 77.245 -81.151 ;
      RECT 77.155 -81.845 77.295 -81.675 ;
      RECT 77.155 -80.349 77.245 -79.342 ;
      RECT 77.155 -79.825 77.295 -79.655 ;
      RECT 77.155 -78.928 77.245 -77.921 ;
      RECT 77.155 -78.615 77.295 -78.445 ;
      RECT 77.155 -77.119 77.245 -76.112 ;
      RECT 77.155 -76.595 77.295 -76.425 ;
      RECT 77.155 -75.698 77.245 -74.691 ;
      RECT 77.155 -75.385 77.295 -75.215 ;
      RECT 77.155 -73.889 77.245 -72.882 ;
      RECT 77.155 -73.365 77.295 -73.195 ;
      RECT 77.155 -72.468 77.245 -71.461 ;
      RECT 77.155 -72.155 77.295 -71.985 ;
      RECT 77.155 -70.659 77.245 -69.652 ;
      RECT 77.155 -70.135 77.295 -69.965 ;
      RECT 77.155 -69.238 77.245 -68.231 ;
      RECT 77.155 -68.925 77.295 -68.755 ;
      RECT 77.155 -67.429 77.245 -66.422 ;
      RECT 77.155 -66.905 77.295 -66.735 ;
      RECT 77.155 -66.008 77.245 -65.001 ;
      RECT 77.155 -65.695 77.295 -65.525 ;
      RECT 77.155 -64.199 77.245 -63.192 ;
      RECT 77.155 -63.675 77.295 -63.505 ;
      RECT 77.155 -62.778 77.245 -61.771 ;
      RECT 77.155 -62.465 77.295 -62.295 ;
      RECT 77.155 -60.969 77.245 -59.962 ;
      RECT 77.155 -60.445 77.295 -60.275 ;
      RECT 77.155 -59.548 77.245 -58.541 ;
      RECT 77.155 -59.235 77.295 -59.065 ;
      RECT 77.155 -57.739 77.245 -56.732 ;
      RECT 77.155 -57.215 77.295 -57.045 ;
      RECT 77.155 -56.318 77.245 -55.311 ;
      RECT 77.155 -56.005 77.295 -55.835 ;
      RECT 77.155 -54.509 77.245 -53.502 ;
      RECT 77.155 -53.985 77.295 -53.815 ;
      RECT 77.155 -53.088 77.245 -52.081 ;
      RECT 77.155 -52.775 77.295 -52.605 ;
      RECT 77.155 -51.279 77.245 -50.272 ;
      RECT 77.155 -50.755 77.295 -50.585 ;
      RECT 77.155 -49.858 77.245 -48.851 ;
      RECT 77.155 -49.545 77.295 -49.375 ;
      RECT 77.155 -48.049 77.245 -47.042 ;
      RECT 77.155 -47.525 77.295 -47.355 ;
      RECT 77.155 -46.628 77.245 -45.621 ;
      RECT 77.155 -46.315 77.295 -46.145 ;
      RECT 77.155 -44.819 77.245 -43.812 ;
      RECT 77.155 -44.295 77.295 -44.125 ;
      RECT 77.155 -43.398 77.245 -42.391 ;
      RECT 77.155 -43.085 77.295 -42.915 ;
      RECT 77.155 -41.589 77.245 -40.582 ;
      RECT 77.155 -41.065 77.295 -40.895 ;
      RECT 77.155 -40.168 77.245 -39.161 ;
      RECT 77.155 -39.855 77.295 -39.685 ;
      RECT 77.155 -38.359 77.245 -37.352 ;
      RECT 77.155 -37.835 77.295 -37.665 ;
      RECT 77.155 -36.938 77.245 -35.931 ;
      RECT 77.155 -36.625 77.295 -36.455 ;
      RECT 77.155 -35.129 77.245 -34.122 ;
      RECT 77.155 -34.605 77.295 -34.435 ;
      RECT 77.155 -33.708 77.245 -32.701 ;
      RECT 77.155 -33.395 77.295 -33.225 ;
      RECT 77.155 -31.899 77.245 -30.892 ;
      RECT 77.155 -31.375 77.295 -31.205 ;
      RECT 77.155 -30.478 77.245 -29.471 ;
      RECT 77.155 -30.165 77.295 -29.995 ;
      RECT 77.155 -28.669 77.245 -27.662 ;
      RECT 77.155 -28.145 77.295 -27.975 ;
      RECT 77.155 -27.248 77.245 -26.241 ;
      RECT 77.155 -26.935 77.295 -26.765 ;
      RECT 77.155 -25.439 77.245 -24.432 ;
      RECT 77.155 -24.915 77.295 -24.745 ;
      RECT 77.155 -24.018 77.245 -23.011 ;
      RECT 77.155 -23.705 77.295 -23.535 ;
      RECT 77.155 -22.209 77.245 -21.202 ;
      RECT 77.155 -21.685 77.295 -21.515 ;
      RECT 77.155 -20.788 77.245 -19.781 ;
      RECT 77.155 -20.475 77.295 -20.305 ;
      RECT 77.155 -18.979 77.245 -17.972 ;
      RECT 77.155 -18.455 77.295 -18.285 ;
      RECT 77.155 -17.558 77.245 -16.551 ;
      RECT 77.155 -17.245 77.295 -17.075 ;
      RECT 77.155 -15.749 77.245 -14.742 ;
      RECT 77.155 -15.225 77.295 -15.055 ;
      RECT 77.155 -14.328 77.245 -13.321 ;
      RECT 77.155 -14.015 77.295 -13.845 ;
      RECT 77.155 -12.519 77.245 -11.512 ;
      RECT 77.155 -11.995 77.295 -11.825 ;
      RECT 77.155 -11.098 77.245 -10.091 ;
      RECT 77.155 -10.785 77.295 -10.615 ;
      RECT 77.155 -9.289 77.245 -8.282 ;
      RECT 77.155 -8.765 77.295 -8.595 ;
      RECT 77.155 -7.868 77.245 -6.861 ;
      RECT 77.155 -7.555 77.295 -7.385 ;
      RECT 77.155 -6.059 77.245 -5.052 ;
      RECT 77.155 -5.535 77.295 -5.365 ;
      RECT 77.155 -4.638 77.245 -3.631 ;
      RECT 77.155 -4.325 77.295 -4.155 ;
      RECT 77.155 -2.829 77.245 -1.822 ;
      RECT 77.155 -2.305 77.295 -2.135 ;
      RECT 77.155 -1.408 77.245 -0.401 ;
      RECT 77.155 -1.095 77.295 -0.925 ;
      RECT 77.155 0.401 77.245 1.408 ;
      RECT 77.155 0.925 77.295 1.095 ;
      RECT 72.985 -108.935 76.765 -108.815 ;
      RECT 74.305 -109.475 74.405 -108.815 ;
      RECT 73.745 -109.475 73.845 -108.815 ;
      RECT 73.185 -109.475 73.285 -108.815 ;
      RECT 76.355 -101.538 76.445 -100.53 ;
      RECT 76.305 -100.935 76.445 -100.765 ;
      RECT 76.355 -99.73 76.445 -98.722 ;
      RECT 76.305 -99.495 76.445 -99.325 ;
      RECT 76.355 -98.308 76.445 -97.3 ;
      RECT 76.305 -97.705 76.445 -97.535 ;
      RECT 76.355 -96.5 76.445 -95.492 ;
      RECT 76.305 -96.265 76.445 -96.095 ;
      RECT 76.355 -95.078 76.445 -94.07 ;
      RECT 76.305 -94.475 76.445 -94.305 ;
      RECT 76.355 -93.27 76.445 -92.262 ;
      RECT 76.305 -93.035 76.445 -92.865 ;
      RECT 76.355 -91.848 76.445 -90.84 ;
      RECT 76.305 -91.245 76.445 -91.075 ;
      RECT 76.355 -90.04 76.445 -89.032 ;
      RECT 76.305 -89.805 76.445 -89.635 ;
      RECT 76.355 -88.618 76.445 -87.61 ;
      RECT 76.305 -88.015 76.445 -87.845 ;
      RECT 76.355 -86.81 76.445 -85.802 ;
      RECT 76.305 -86.575 76.445 -86.405 ;
      RECT 76.355 -85.388 76.445 -84.38 ;
      RECT 76.305 -84.785 76.445 -84.615 ;
      RECT 76.355 -83.58 76.445 -82.572 ;
      RECT 76.305 -83.345 76.445 -83.175 ;
      RECT 76.355 -82.158 76.445 -81.15 ;
      RECT 76.305 -81.555 76.445 -81.385 ;
      RECT 76.355 -80.35 76.445 -79.342 ;
      RECT 76.305 -80.115 76.445 -79.945 ;
      RECT 76.355 -78.928 76.445 -77.92 ;
      RECT 76.305 -78.325 76.445 -78.155 ;
      RECT 76.355 -77.12 76.445 -76.112 ;
      RECT 76.305 -76.885 76.445 -76.715 ;
      RECT 76.355 -75.698 76.445 -74.69 ;
      RECT 76.305 -75.095 76.445 -74.925 ;
      RECT 76.355 -73.89 76.445 -72.882 ;
      RECT 76.305 -73.655 76.445 -73.485 ;
      RECT 76.355 -72.468 76.445 -71.46 ;
      RECT 76.305 -71.865 76.445 -71.695 ;
      RECT 76.355 -70.66 76.445 -69.652 ;
      RECT 76.305 -70.425 76.445 -70.255 ;
      RECT 76.355 -69.238 76.445 -68.23 ;
      RECT 76.305 -68.635 76.445 -68.465 ;
      RECT 76.355 -67.43 76.445 -66.422 ;
      RECT 76.305 -67.195 76.445 -67.025 ;
      RECT 76.355 -66.008 76.445 -65 ;
      RECT 76.305 -65.405 76.445 -65.235 ;
      RECT 76.355 -64.2 76.445 -63.192 ;
      RECT 76.305 -63.965 76.445 -63.795 ;
      RECT 76.355 -62.778 76.445 -61.77 ;
      RECT 76.305 -62.175 76.445 -62.005 ;
      RECT 76.355 -60.97 76.445 -59.962 ;
      RECT 76.305 -60.735 76.445 -60.565 ;
      RECT 76.355 -59.548 76.445 -58.54 ;
      RECT 76.305 -58.945 76.445 -58.775 ;
      RECT 76.355 -57.74 76.445 -56.732 ;
      RECT 76.305 -57.505 76.445 -57.335 ;
      RECT 76.355 -56.318 76.445 -55.31 ;
      RECT 76.305 -55.715 76.445 -55.545 ;
      RECT 76.355 -54.51 76.445 -53.502 ;
      RECT 76.305 -54.275 76.445 -54.105 ;
      RECT 76.355 -53.088 76.445 -52.08 ;
      RECT 76.305 -52.485 76.445 -52.315 ;
      RECT 76.355 -51.28 76.445 -50.272 ;
      RECT 76.305 -51.045 76.445 -50.875 ;
      RECT 76.355 -49.858 76.445 -48.85 ;
      RECT 76.305 -49.255 76.445 -49.085 ;
      RECT 76.355 -48.05 76.445 -47.042 ;
      RECT 76.305 -47.815 76.445 -47.645 ;
      RECT 76.355 -46.628 76.445 -45.62 ;
      RECT 76.305 -46.025 76.445 -45.855 ;
      RECT 76.355 -44.82 76.445 -43.812 ;
      RECT 76.305 -44.585 76.445 -44.415 ;
      RECT 76.355 -43.398 76.445 -42.39 ;
      RECT 76.305 -42.795 76.445 -42.625 ;
      RECT 76.355 -41.59 76.445 -40.582 ;
      RECT 76.305 -41.355 76.445 -41.185 ;
      RECT 76.355 -40.168 76.445 -39.16 ;
      RECT 76.305 -39.565 76.445 -39.395 ;
      RECT 76.355 -38.36 76.445 -37.352 ;
      RECT 76.305 -38.125 76.445 -37.955 ;
      RECT 76.355 -36.938 76.445 -35.93 ;
      RECT 76.305 -36.335 76.445 -36.165 ;
      RECT 76.355 -35.13 76.445 -34.122 ;
      RECT 76.305 -34.895 76.445 -34.725 ;
      RECT 76.355 -33.708 76.445 -32.7 ;
      RECT 76.305 -33.105 76.445 -32.935 ;
      RECT 76.355 -31.9 76.445 -30.892 ;
      RECT 76.305 -31.665 76.445 -31.495 ;
      RECT 76.355 -30.478 76.445 -29.47 ;
      RECT 76.305 -29.875 76.445 -29.705 ;
      RECT 76.355 -28.67 76.445 -27.662 ;
      RECT 76.305 -28.435 76.445 -28.265 ;
      RECT 76.355 -27.248 76.445 -26.24 ;
      RECT 76.305 -26.645 76.445 -26.475 ;
      RECT 76.355 -25.44 76.445 -24.432 ;
      RECT 76.305 -25.205 76.445 -25.035 ;
      RECT 76.355 -24.018 76.445 -23.01 ;
      RECT 76.305 -23.415 76.445 -23.245 ;
      RECT 76.355 -22.21 76.445 -21.202 ;
      RECT 76.305 -21.975 76.445 -21.805 ;
      RECT 76.355 -20.788 76.445 -19.78 ;
      RECT 76.305 -20.185 76.445 -20.015 ;
      RECT 76.355 -18.98 76.445 -17.972 ;
      RECT 76.305 -18.745 76.445 -18.575 ;
      RECT 76.355 -17.558 76.445 -16.55 ;
      RECT 76.305 -16.955 76.445 -16.785 ;
      RECT 76.355 -15.75 76.445 -14.742 ;
      RECT 76.305 -15.515 76.445 -15.345 ;
      RECT 76.355 -14.328 76.445 -13.32 ;
      RECT 76.305 -13.725 76.445 -13.555 ;
      RECT 76.355 -12.52 76.445 -11.512 ;
      RECT 76.305 -12.285 76.445 -12.115 ;
      RECT 76.355 -11.098 76.445 -10.09 ;
      RECT 76.305 -10.495 76.445 -10.325 ;
      RECT 76.355 -9.29 76.445 -8.282 ;
      RECT 76.305 -9.055 76.445 -8.885 ;
      RECT 76.355 -7.868 76.445 -6.86 ;
      RECT 76.305 -7.265 76.445 -7.095 ;
      RECT 76.355 -6.06 76.445 -5.052 ;
      RECT 76.305 -5.825 76.445 -5.655 ;
      RECT 76.355 -4.638 76.445 -3.63 ;
      RECT 76.305 -4.035 76.445 -3.865 ;
      RECT 76.355 -2.83 76.445 -1.822 ;
      RECT 76.305 -2.595 76.445 -2.425 ;
      RECT 76.355 -1.408 76.445 -0.4 ;
      RECT 76.305 -0.805 76.445 -0.635 ;
      RECT 76.355 0.4 76.445 1.408 ;
      RECT 76.305 0.635 76.445 0.805 ;
      RECT 74.925 -111.685 76.405 -111.585 ;
      RECT 74.925 -112.195 75.025 -111.585 ;
      RECT 75.145 -109.15 76.405 -109.05 ;
      RECT 76.305 -109.475 76.405 -109.05 ;
      RECT 75.745 -109.475 75.845 -109.05 ;
      RECT 75.185 -109.475 75.285 -109.05 ;
      RECT 75.955 -101.538 76.045 -100.531 ;
      RECT 75.955 -101.225 76.095 -101.055 ;
      RECT 75.955 -99.729 76.045 -98.722 ;
      RECT 75.955 -99.205 76.095 -99.035 ;
      RECT 75.955 -98.308 76.045 -97.301 ;
      RECT 75.955 -97.995 76.095 -97.825 ;
      RECT 75.955 -96.499 76.045 -95.492 ;
      RECT 75.955 -95.975 76.095 -95.805 ;
      RECT 75.955 -95.078 76.045 -94.071 ;
      RECT 75.955 -94.765 76.095 -94.595 ;
      RECT 75.955 -93.269 76.045 -92.262 ;
      RECT 75.955 -92.745 76.095 -92.575 ;
      RECT 75.955 -91.848 76.045 -90.841 ;
      RECT 75.955 -91.535 76.095 -91.365 ;
      RECT 75.955 -90.039 76.045 -89.032 ;
      RECT 75.955 -89.515 76.095 -89.345 ;
      RECT 75.955 -88.618 76.045 -87.611 ;
      RECT 75.955 -88.305 76.095 -88.135 ;
      RECT 75.955 -86.809 76.045 -85.802 ;
      RECT 75.955 -86.285 76.095 -86.115 ;
      RECT 75.955 -85.388 76.045 -84.381 ;
      RECT 75.955 -85.075 76.095 -84.905 ;
      RECT 75.955 -83.579 76.045 -82.572 ;
      RECT 75.955 -83.055 76.095 -82.885 ;
      RECT 75.955 -82.158 76.045 -81.151 ;
      RECT 75.955 -81.845 76.095 -81.675 ;
      RECT 75.955 -80.349 76.045 -79.342 ;
      RECT 75.955 -79.825 76.095 -79.655 ;
      RECT 75.955 -78.928 76.045 -77.921 ;
      RECT 75.955 -78.615 76.095 -78.445 ;
      RECT 75.955 -77.119 76.045 -76.112 ;
      RECT 75.955 -76.595 76.095 -76.425 ;
      RECT 75.955 -75.698 76.045 -74.691 ;
      RECT 75.955 -75.385 76.095 -75.215 ;
      RECT 75.955 -73.889 76.045 -72.882 ;
      RECT 75.955 -73.365 76.095 -73.195 ;
      RECT 75.955 -72.468 76.045 -71.461 ;
      RECT 75.955 -72.155 76.095 -71.985 ;
      RECT 75.955 -70.659 76.045 -69.652 ;
      RECT 75.955 -70.135 76.095 -69.965 ;
      RECT 75.955 -69.238 76.045 -68.231 ;
      RECT 75.955 -68.925 76.095 -68.755 ;
      RECT 75.955 -67.429 76.045 -66.422 ;
      RECT 75.955 -66.905 76.095 -66.735 ;
      RECT 75.955 -66.008 76.045 -65.001 ;
      RECT 75.955 -65.695 76.095 -65.525 ;
      RECT 75.955 -64.199 76.045 -63.192 ;
      RECT 75.955 -63.675 76.095 -63.505 ;
      RECT 75.955 -62.778 76.045 -61.771 ;
      RECT 75.955 -62.465 76.095 -62.295 ;
      RECT 75.955 -60.969 76.045 -59.962 ;
      RECT 75.955 -60.445 76.095 -60.275 ;
      RECT 75.955 -59.548 76.045 -58.541 ;
      RECT 75.955 -59.235 76.095 -59.065 ;
      RECT 75.955 -57.739 76.045 -56.732 ;
      RECT 75.955 -57.215 76.095 -57.045 ;
      RECT 75.955 -56.318 76.045 -55.311 ;
      RECT 75.955 -56.005 76.095 -55.835 ;
      RECT 75.955 -54.509 76.045 -53.502 ;
      RECT 75.955 -53.985 76.095 -53.815 ;
      RECT 75.955 -53.088 76.045 -52.081 ;
      RECT 75.955 -52.775 76.095 -52.605 ;
      RECT 75.955 -51.279 76.045 -50.272 ;
      RECT 75.955 -50.755 76.095 -50.585 ;
      RECT 75.955 -49.858 76.045 -48.851 ;
      RECT 75.955 -49.545 76.095 -49.375 ;
      RECT 75.955 -48.049 76.045 -47.042 ;
      RECT 75.955 -47.525 76.095 -47.355 ;
      RECT 75.955 -46.628 76.045 -45.621 ;
      RECT 75.955 -46.315 76.095 -46.145 ;
      RECT 75.955 -44.819 76.045 -43.812 ;
      RECT 75.955 -44.295 76.095 -44.125 ;
      RECT 75.955 -43.398 76.045 -42.391 ;
      RECT 75.955 -43.085 76.095 -42.915 ;
      RECT 75.955 -41.589 76.045 -40.582 ;
      RECT 75.955 -41.065 76.095 -40.895 ;
      RECT 75.955 -40.168 76.045 -39.161 ;
      RECT 75.955 -39.855 76.095 -39.685 ;
      RECT 75.955 -38.359 76.045 -37.352 ;
      RECT 75.955 -37.835 76.095 -37.665 ;
      RECT 75.955 -36.938 76.045 -35.931 ;
      RECT 75.955 -36.625 76.095 -36.455 ;
      RECT 75.955 -35.129 76.045 -34.122 ;
      RECT 75.955 -34.605 76.095 -34.435 ;
      RECT 75.955 -33.708 76.045 -32.701 ;
      RECT 75.955 -33.395 76.095 -33.225 ;
      RECT 75.955 -31.899 76.045 -30.892 ;
      RECT 75.955 -31.375 76.095 -31.205 ;
      RECT 75.955 -30.478 76.045 -29.471 ;
      RECT 75.955 -30.165 76.095 -29.995 ;
      RECT 75.955 -28.669 76.045 -27.662 ;
      RECT 75.955 -28.145 76.095 -27.975 ;
      RECT 75.955 -27.248 76.045 -26.241 ;
      RECT 75.955 -26.935 76.095 -26.765 ;
      RECT 75.955 -25.439 76.045 -24.432 ;
      RECT 75.955 -24.915 76.095 -24.745 ;
      RECT 75.955 -24.018 76.045 -23.011 ;
      RECT 75.955 -23.705 76.095 -23.535 ;
      RECT 75.955 -22.209 76.045 -21.202 ;
      RECT 75.955 -21.685 76.095 -21.515 ;
      RECT 75.955 -20.788 76.045 -19.781 ;
      RECT 75.955 -20.475 76.095 -20.305 ;
      RECT 75.955 -18.979 76.045 -17.972 ;
      RECT 75.955 -18.455 76.095 -18.285 ;
      RECT 75.955 -17.558 76.045 -16.551 ;
      RECT 75.955 -17.245 76.095 -17.075 ;
      RECT 75.955 -15.749 76.045 -14.742 ;
      RECT 75.955 -15.225 76.095 -15.055 ;
      RECT 75.955 -14.328 76.045 -13.321 ;
      RECT 75.955 -14.015 76.095 -13.845 ;
      RECT 75.955 -12.519 76.045 -11.512 ;
      RECT 75.955 -11.995 76.095 -11.825 ;
      RECT 75.955 -11.098 76.045 -10.091 ;
      RECT 75.955 -10.785 76.095 -10.615 ;
      RECT 75.955 -9.289 76.045 -8.282 ;
      RECT 75.955 -8.765 76.095 -8.595 ;
      RECT 75.955 -7.868 76.045 -6.861 ;
      RECT 75.955 -7.555 76.095 -7.385 ;
      RECT 75.955 -6.059 76.045 -5.052 ;
      RECT 75.955 -5.535 76.095 -5.365 ;
      RECT 75.955 -4.638 76.045 -3.631 ;
      RECT 75.955 -4.325 76.095 -4.155 ;
      RECT 75.955 -2.829 76.045 -1.822 ;
      RECT 75.955 -2.305 76.095 -2.135 ;
      RECT 75.955 -1.408 76.045 -0.401 ;
      RECT 75.955 -1.095 76.095 -0.925 ;
      RECT 75.955 0.401 76.045 1.408 ;
      RECT 75.955 0.925 76.095 1.095 ;
      RECT 75.285 -111.495 75.455 -111.385 ;
      RECT 72.135 -111.495 75.455 -111.395 ;
      RECT 75.155 -101.538 75.245 -100.53 ;
      RECT 75.105 -100.935 75.245 -100.765 ;
      RECT 75.155 -99.73 75.245 -98.722 ;
      RECT 75.105 -99.495 75.245 -99.325 ;
      RECT 75.155 -98.308 75.245 -97.3 ;
      RECT 75.105 -97.705 75.245 -97.535 ;
      RECT 75.155 -96.5 75.245 -95.492 ;
      RECT 75.105 -96.265 75.245 -96.095 ;
      RECT 75.155 -95.078 75.245 -94.07 ;
      RECT 75.105 -94.475 75.245 -94.305 ;
      RECT 75.155 -93.27 75.245 -92.262 ;
      RECT 75.105 -93.035 75.245 -92.865 ;
      RECT 75.155 -91.848 75.245 -90.84 ;
      RECT 75.105 -91.245 75.245 -91.075 ;
      RECT 75.155 -90.04 75.245 -89.032 ;
      RECT 75.105 -89.805 75.245 -89.635 ;
      RECT 75.155 -88.618 75.245 -87.61 ;
      RECT 75.105 -88.015 75.245 -87.845 ;
      RECT 75.155 -86.81 75.245 -85.802 ;
      RECT 75.105 -86.575 75.245 -86.405 ;
      RECT 75.155 -85.388 75.245 -84.38 ;
      RECT 75.105 -84.785 75.245 -84.615 ;
      RECT 75.155 -83.58 75.245 -82.572 ;
      RECT 75.105 -83.345 75.245 -83.175 ;
      RECT 75.155 -82.158 75.245 -81.15 ;
      RECT 75.105 -81.555 75.245 -81.385 ;
      RECT 75.155 -80.35 75.245 -79.342 ;
      RECT 75.105 -80.115 75.245 -79.945 ;
      RECT 75.155 -78.928 75.245 -77.92 ;
      RECT 75.105 -78.325 75.245 -78.155 ;
      RECT 75.155 -77.12 75.245 -76.112 ;
      RECT 75.105 -76.885 75.245 -76.715 ;
      RECT 75.155 -75.698 75.245 -74.69 ;
      RECT 75.105 -75.095 75.245 -74.925 ;
      RECT 75.155 -73.89 75.245 -72.882 ;
      RECT 75.105 -73.655 75.245 -73.485 ;
      RECT 75.155 -72.468 75.245 -71.46 ;
      RECT 75.105 -71.865 75.245 -71.695 ;
      RECT 75.155 -70.66 75.245 -69.652 ;
      RECT 75.105 -70.425 75.245 -70.255 ;
      RECT 75.155 -69.238 75.245 -68.23 ;
      RECT 75.105 -68.635 75.245 -68.465 ;
      RECT 75.155 -67.43 75.245 -66.422 ;
      RECT 75.105 -67.195 75.245 -67.025 ;
      RECT 75.155 -66.008 75.245 -65 ;
      RECT 75.105 -65.405 75.245 -65.235 ;
      RECT 75.155 -64.2 75.245 -63.192 ;
      RECT 75.105 -63.965 75.245 -63.795 ;
      RECT 75.155 -62.778 75.245 -61.77 ;
      RECT 75.105 -62.175 75.245 -62.005 ;
      RECT 75.155 -60.97 75.245 -59.962 ;
      RECT 75.105 -60.735 75.245 -60.565 ;
      RECT 75.155 -59.548 75.245 -58.54 ;
      RECT 75.105 -58.945 75.245 -58.775 ;
      RECT 75.155 -57.74 75.245 -56.732 ;
      RECT 75.105 -57.505 75.245 -57.335 ;
      RECT 75.155 -56.318 75.245 -55.31 ;
      RECT 75.105 -55.715 75.245 -55.545 ;
      RECT 75.155 -54.51 75.245 -53.502 ;
      RECT 75.105 -54.275 75.245 -54.105 ;
      RECT 75.155 -53.088 75.245 -52.08 ;
      RECT 75.105 -52.485 75.245 -52.315 ;
      RECT 75.155 -51.28 75.245 -50.272 ;
      RECT 75.105 -51.045 75.245 -50.875 ;
      RECT 75.155 -49.858 75.245 -48.85 ;
      RECT 75.105 -49.255 75.245 -49.085 ;
      RECT 75.155 -48.05 75.245 -47.042 ;
      RECT 75.105 -47.815 75.245 -47.645 ;
      RECT 75.155 -46.628 75.245 -45.62 ;
      RECT 75.105 -46.025 75.245 -45.855 ;
      RECT 75.155 -44.82 75.245 -43.812 ;
      RECT 75.105 -44.585 75.245 -44.415 ;
      RECT 75.155 -43.398 75.245 -42.39 ;
      RECT 75.105 -42.795 75.245 -42.625 ;
      RECT 75.155 -41.59 75.245 -40.582 ;
      RECT 75.105 -41.355 75.245 -41.185 ;
      RECT 75.155 -40.168 75.245 -39.16 ;
      RECT 75.105 -39.565 75.245 -39.395 ;
      RECT 75.155 -38.36 75.245 -37.352 ;
      RECT 75.105 -38.125 75.245 -37.955 ;
      RECT 75.155 -36.938 75.245 -35.93 ;
      RECT 75.105 -36.335 75.245 -36.165 ;
      RECT 75.155 -35.13 75.245 -34.122 ;
      RECT 75.105 -34.895 75.245 -34.725 ;
      RECT 75.155 -33.708 75.245 -32.7 ;
      RECT 75.105 -33.105 75.245 -32.935 ;
      RECT 75.155 -31.9 75.245 -30.892 ;
      RECT 75.105 -31.665 75.245 -31.495 ;
      RECT 75.155 -30.478 75.245 -29.47 ;
      RECT 75.105 -29.875 75.245 -29.705 ;
      RECT 75.155 -28.67 75.245 -27.662 ;
      RECT 75.105 -28.435 75.245 -28.265 ;
      RECT 75.155 -27.248 75.245 -26.24 ;
      RECT 75.105 -26.645 75.245 -26.475 ;
      RECT 75.155 -25.44 75.245 -24.432 ;
      RECT 75.105 -25.205 75.245 -25.035 ;
      RECT 75.155 -24.018 75.245 -23.01 ;
      RECT 75.105 -23.415 75.245 -23.245 ;
      RECT 75.155 -22.21 75.245 -21.202 ;
      RECT 75.105 -21.975 75.245 -21.805 ;
      RECT 75.155 -20.788 75.245 -19.78 ;
      RECT 75.105 -20.185 75.245 -20.015 ;
      RECT 75.155 -18.98 75.245 -17.972 ;
      RECT 75.105 -18.745 75.245 -18.575 ;
      RECT 75.155 -17.558 75.245 -16.55 ;
      RECT 75.105 -16.955 75.245 -16.785 ;
      RECT 75.155 -15.75 75.245 -14.742 ;
      RECT 75.105 -15.515 75.245 -15.345 ;
      RECT 75.155 -14.328 75.245 -13.32 ;
      RECT 75.105 -13.725 75.245 -13.555 ;
      RECT 75.155 -12.52 75.245 -11.512 ;
      RECT 75.105 -12.285 75.245 -12.115 ;
      RECT 75.155 -11.098 75.245 -10.09 ;
      RECT 75.105 -10.495 75.245 -10.325 ;
      RECT 75.155 -9.29 75.245 -8.282 ;
      RECT 75.105 -9.055 75.245 -8.885 ;
      RECT 75.155 -7.868 75.245 -6.86 ;
      RECT 75.105 -7.265 75.245 -7.095 ;
      RECT 75.155 -6.06 75.245 -5.052 ;
      RECT 75.105 -5.825 75.245 -5.655 ;
      RECT 75.155 -4.638 75.245 -3.63 ;
      RECT 75.105 -4.035 75.245 -3.865 ;
      RECT 75.155 -2.83 75.245 -1.822 ;
      RECT 75.105 -2.595 75.245 -2.425 ;
      RECT 75.155 -1.408 75.245 -0.4 ;
      RECT 75.105 -0.805 75.245 -0.635 ;
      RECT 75.155 0.4 75.245 1.408 ;
      RECT 75.105 0.635 75.245 0.805 ;
      RECT 74.755 -101.538 74.845 -100.531 ;
      RECT 74.755 -101.225 74.895 -101.055 ;
      RECT 74.755 -99.729 74.845 -98.722 ;
      RECT 74.755 -99.205 74.895 -99.035 ;
      RECT 74.755 -98.308 74.845 -97.301 ;
      RECT 74.755 -97.995 74.895 -97.825 ;
      RECT 74.755 -96.499 74.845 -95.492 ;
      RECT 74.755 -95.975 74.895 -95.805 ;
      RECT 74.755 -95.078 74.845 -94.071 ;
      RECT 74.755 -94.765 74.895 -94.595 ;
      RECT 74.755 -93.269 74.845 -92.262 ;
      RECT 74.755 -92.745 74.895 -92.575 ;
      RECT 74.755 -91.848 74.845 -90.841 ;
      RECT 74.755 -91.535 74.895 -91.365 ;
      RECT 74.755 -90.039 74.845 -89.032 ;
      RECT 74.755 -89.515 74.895 -89.345 ;
      RECT 74.755 -88.618 74.845 -87.611 ;
      RECT 74.755 -88.305 74.895 -88.135 ;
      RECT 74.755 -86.809 74.845 -85.802 ;
      RECT 74.755 -86.285 74.895 -86.115 ;
      RECT 74.755 -85.388 74.845 -84.381 ;
      RECT 74.755 -85.075 74.895 -84.905 ;
      RECT 74.755 -83.579 74.845 -82.572 ;
      RECT 74.755 -83.055 74.895 -82.885 ;
      RECT 74.755 -82.158 74.845 -81.151 ;
      RECT 74.755 -81.845 74.895 -81.675 ;
      RECT 74.755 -80.349 74.845 -79.342 ;
      RECT 74.755 -79.825 74.895 -79.655 ;
      RECT 74.755 -78.928 74.845 -77.921 ;
      RECT 74.755 -78.615 74.895 -78.445 ;
      RECT 74.755 -77.119 74.845 -76.112 ;
      RECT 74.755 -76.595 74.895 -76.425 ;
      RECT 74.755 -75.698 74.845 -74.691 ;
      RECT 74.755 -75.385 74.895 -75.215 ;
      RECT 74.755 -73.889 74.845 -72.882 ;
      RECT 74.755 -73.365 74.895 -73.195 ;
      RECT 74.755 -72.468 74.845 -71.461 ;
      RECT 74.755 -72.155 74.895 -71.985 ;
      RECT 74.755 -70.659 74.845 -69.652 ;
      RECT 74.755 -70.135 74.895 -69.965 ;
      RECT 74.755 -69.238 74.845 -68.231 ;
      RECT 74.755 -68.925 74.895 -68.755 ;
      RECT 74.755 -67.429 74.845 -66.422 ;
      RECT 74.755 -66.905 74.895 -66.735 ;
      RECT 74.755 -66.008 74.845 -65.001 ;
      RECT 74.755 -65.695 74.895 -65.525 ;
      RECT 74.755 -64.199 74.845 -63.192 ;
      RECT 74.755 -63.675 74.895 -63.505 ;
      RECT 74.755 -62.778 74.845 -61.771 ;
      RECT 74.755 -62.465 74.895 -62.295 ;
      RECT 74.755 -60.969 74.845 -59.962 ;
      RECT 74.755 -60.445 74.895 -60.275 ;
      RECT 74.755 -59.548 74.845 -58.541 ;
      RECT 74.755 -59.235 74.895 -59.065 ;
      RECT 74.755 -57.739 74.845 -56.732 ;
      RECT 74.755 -57.215 74.895 -57.045 ;
      RECT 74.755 -56.318 74.845 -55.311 ;
      RECT 74.755 -56.005 74.895 -55.835 ;
      RECT 74.755 -54.509 74.845 -53.502 ;
      RECT 74.755 -53.985 74.895 -53.815 ;
      RECT 74.755 -53.088 74.845 -52.081 ;
      RECT 74.755 -52.775 74.895 -52.605 ;
      RECT 74.755 -51.279 74.845 -50.272 ;
      RECT 74.755 -50.755 74.895 -50.585 ;
      RECT 74.755 -49.858 74.845 -48.851 ;
      RECT 74.755 -49.545 74.895 -49.375 ;
      RECT 74.755 -48.049 74.845 -47.042 ;
      RECT 74.755 -47.525 74.895 -47.355 ;
      RECT 74.755 -46.628 74.845 -45.621 ;
      RECT 74.755 -46.315 74.895 -46.145 ;
      RECT 74.755 -44.819 74.845 -43.812 ;
      RECT 74.755 -44.295 74.895 -44.125 ;
      RECT 74.755 -43.398 74.845 -42.391 ;
      RECT 74.755 -43.085 74.895 -42.915 ;
      RECT 74.755 -41.589 74.845 -40.582 ;
      RECT 74.755 -41.065 74.895 -40.895 ;
      RECT 74.755 -40.168 74.845 -39.161 ;
      RECT 74.755 -39.855 74.895 -39.685 ;
      RECT 74.755 -38.359 74.845 -37.352 ;
      RECT 74.755 -37.835 74.895 -37.665 ;
      RECT 74.755 -36.938 74.845 -35.931 ;
      RECT 74.755 -36.625 74.895 -36.455 ;
      RECT 74.755 -35.129 74.845 -34.122 ;
      RECT 74.755 -34.605 74.895 -34.435 ;
      RECT 74.755 -33.708 74.845 -32.701 ;
      RECT 74.755 -33.395 74.895 -33.225 ;
      RECT 74.755 -31.899 74.845 -30.892 ;
      RECT 74.755 -31.375 74.895 -31.205 ;
      RECT 74.755 -30.478 74.845 -29.471 ;
      RECT 74.755 -30.165 74.895 -29.995 ;
      RECT 74.755 -28.669 74.845 -27.662 ;
      RECT 74.755 -28.145 74.895 -27.975 ;
      RECT 74.755 -27.248 74.845 -26.241 ;
      RECT 74.755 -26.935 74.895 -26.765 ;
      RECT 74.755 -25.439 74.845 -24.432 ;
      RECT 74.755 -24.915 74.895 -24.745 ;
      RECT 74.755 -24.018 74.845 -23.011 ;
      RECT 74.755 -23.705 74.895 -23.535 ;
      RECT 74.755 -22.209 74.845 -21.202 ;
      RECT 74.755 -21.685 74.895 -21.515 ;
      RECT 74.755 -20.788 74.845 -19.781 ;
      RECT 74.755 -20.475 74.895 -20.305 ;
      RECT 74.755 -18.979 74.845 -17.972 ;
      RECT 74.755 -18.455 74.895 -18.285 ;
      RECT 74.755 -17.558 74.845 -16.551 ;
      RECT 74.755 -17.245 74.895 -17.075 ;
      RECT 74.755 -15.749 74.845 -14.742 ;
      RECT 74.755 -15.225 74.895 -15.055 ;
      RECT 74.755 -14.328 74.845 -13.321 ;
      RECT 74.755 -14.015 74.895 -13.845 ;
      RECT 74.755 -12.519 74.845 -11.512 ;
      RECT 74.755 -11.995 74.895 -11.825 ;
      RECT 74.755 -11.098 74.845 -10.091 ;
      RECT 74.755 -10.785 74.895 -10.615 ;
      RECT 74.755 -9.289 74.845 -8.282 ;
      RECT 74.755 -8.765 74.895 -8.595 ;
      RECT 74.755 -7.868 74.845 -6.861 ;
      RECT 74.755 -7.555 74.895 -7.385 ;
      RECT 74.755 -6.059 74.845 -5.052 ;
      RECT 74.755 -5.535 74.895 -5.365 ;
      RECT 74.755 -4.638 74.845 -3.631 ;
      RECT 74.755 -4.325 74.895 -4.155 ;
      RECT 74.755 -2.829 74.845 -1.822 ;
      RECT 74.755 -2.305 74.895 -2.135 ;
      RECT 74.755 -1.408 74.845 -0.401 ;
      RECT 74.755 -1.095 74.895 -0.925 ;
      RECT 74.755 0.401 74.845 1.408 ;
      RECT 74.755 0.925 74.895 1.095 ;
      RECT 72.905 -111.685 74.385 -111.585 ;
      RECT 72.905 -112.055 73.005 -111.585 ;
      RECT 72.71 -114.395 74.285 -114.275 ;
      RECT 74.185 -114.895 74.285 -114.275 ;
      RECT 73.59 -114.895 73.69 -114.275 ;
      RECT 72.71 -114.85 72.81 -114.275 ;
      RECT 73.955 -101.538 74.045 -100.53 ;
      RECT 73.905 -100.935 74.045 -100.765 ;
      RECT 73.955 -99.73 74.045 -98.722 ;
      RECT 73.905 -99.495 74.045 -99.325 ;
      RECT 73.955 -98.308 74.045 -97.3 ;
      RECT 73.905 -97.705 74.045 -97.535 ;
      RECT 73.955 -96.5 74.045 -95.492 ;
      RECT 73.905 -96.265 74.045 -96.095 ;
      RECT 73.955 -95.078 74.045 -94.07 ;
      RECT 73.905 -94.475 74.045 -94.305 ;
      RECT 73.955 -93.27 74.045 -92.262 ;
      RECT 73.905 -93.035 74.045 -92.865 ;
      RECT 73.955 -91.848 74.045 -90.84 ;
      RECT 73.905 -91.245 74.045 -91.075 ;
      RECT 73.955 -90.04 74.045 -89.032 ;
      RECT 73.905 -89.805 74.045 -89.635 ;
      RECT 73.955 -88.618 74.045 -87.61 ;
      RECT 73.905 -88.015 74.045 -87.845 ;
      RECT 73.955 -86.81 74.045 -85.802 ;
      RECT 73.905 -86.575 74.045 -86.405 ;
      RECT 73.955 -85.388 74.045 -84.38 ;
      RECT 73.905 -84.785 74.045 -84.615 ;
      RECT 73.955 -83.58 74.045 -82.572 ;
      RECT 73.905 -83.345 74.045 -83.175 ;
      RECT 73.955 -82.158 74.045 -81.15 ;
      RECT 73.905 -81.555 74.045 -81.385 ;
      RECT 73.955 -80.35 74.045 -79.342 ;
      RECT 73.905 -80.115 74.045 -79.945 ;
      RECT 73.955 -78.928 74.045 -77.92 ;
      RECT 73.905 -78.325 74.045 -78.155 ;
      RECT 73.955 -77.12 74.045 -76.112 ;
      RECT 73.905 -76.885 74.045 -76.715 ;
      RECT 73.955 -75.698 74.045 -74.69 ;
      RECT 73.905 -75.095 74.045 -74.925 ;
      RECT 73.955 -73.89 74.045 -72.882 ;
      RECT 73.905 -73.655 74.045 -73.485 ;
      RECT 73.955 -72.468 74.045 -71.46 ;
      RECT 73.905 -71.865 74.045 -71.695 ;
      RECT 73.955 -70.66 74.045 -69.652 ;
      RECT 73.905 -70.425 74.045 -70.255 ;
      RECT 73.955 -69.238 74.045 -68.23 ;
      RECT 73.905 -68.635 74.045 -68.465 ;
      RECT 73.955 -67.43 74.045 -66.422 ;
      RECT 73.905 -67.195 74.045 -67.025 ;
      RECT 73.955 -66.008 74.045 -65 ;
      RECT 73.905 -65.405 74.045 -65.235 ;
      RECT 73.955 -64.2 74.045 -63.192 ;
      RECT 73.905 -63.965 74.045 -63.795 ;
      RECT 73.955 -62.778 74.045 -61.77 ;
      RECT 73.905 -62.175 74.045 -62.005 ;
      RECT 73.955 -60.97 74.045 -59.962 ;
      RECT 73.905 -60.735 74.045 -60.565 ;
      RECT 73.955 -59.548 74.045 -58.54 ;
      RECT 73.905 -58.945 74.045 -58.775 ;
      RECT 73.955 -57.74 74.045 -56.732 ;
      RECT 73.905 -57.505 74.045 -57.335 ;
      RECT 73.955 -56.318 74.045 -55.31 ;
      RECT 73.905 -55.715 74.045 -55.545 ;
      RECT 73.955 -54.51 74.045 -53.502 ;
      RECT 73.905 -54.275 74.045 -54.105 ;
      RECT 73.955 -53.088 74.045 -52.08 ;
      RECT 73.905 -52.485 74.045 -52.315 ;
      RECT 73.955 -51.28 74.045 -50.272 ;
      RECT 73.905 -51.045 74.045 -50.875 ;
      RECT 73.955 -49.858 74.045 -48.85 ;
      RECT 73.905 -49.255 74.045 -49.085 ;
      RECT 73.955 -48.05 74.045 -47.042 ;
      RECT 73.905 -47.815 74.045 -47.645 ;
      RECT 73.955 -46.628 74.045 -45.62 ;
      RECT 73.905 -46.025 74.045 -45.855 ;
      RECT 73.955 -44.82 74.045 -43.812 ;
      RECT 73.905 -44.585 74.045 -44.415 ;
      RECT 73.955 -43.398 74.045 -42.39 ;
      RECT 73.905 -42.795 74.045 -42.625 ;
      RECT 73.955 -41.59 74.045 -40.582 ;
      RECT 73.905 -41.355 74.045 -41.185 ;
      RECT 73.955 -40.168 74.045 -39.16 ;
      RECT 73.905 -39.565 74.045 -39.395 ;
      RECT 73.955 -38.36 74.045 -37.352 ;
      RECT 73.905 -38.125 74.045 -37.955 ;
      RECT 73.955 -36.938 74.045 -35.93 ;
      RECT 73.905 -36.335 74.045 -36.165 ;
      RECT 73.955 -35.13 74.045 -34.122 ;
      RECT 73.905 -34.895 74.045 -34.725 ;
      RECT 73.955 -33.708 74.045 -32.7 ;
      RECT 73.905 -33.105 74.045 -32.935 ;
      RECT 73.955 -31.9 74.045 -30.892 ;
      RECT 73.905 -31.665 74.045 -31.495 ;
      RECT 73.955 -30.478 74.045 -29.47 ;
      RECT 73.905 -29.875 74.045 -29.705 ;
      RECT 73.955 -28.67 74.045 -27.662 ;
      RECT 73.905 -28.435 74.045 -28.265 ;
      RECT 73.955 -27.248 74.045 -26.24 ;
      RECT 73.905 -26.645 74.045 -26.475 ;
      RECT 73.955 -25.44 74.045 -24.432 ;
      RECT 73.905 -25.205 74.045 -25.035 ;
      RECT 73.955 -24.018 74.045 -23.01 ;
      RECT 73.905 -23.415 74.045 -23.245 ;
      RECT 73.955 -22.21 74.045 -21.202 ;
      RECT 73.905 -21.975 74.045 -21.805 ;
      RECT 73.955 -20.788 74.045 -19.78 ;
      RECT 73.905 -20.185 74.045 -20.015 ;
      RECT 73.955 -18.98 74.045 -17.972 ;
      RECT 73.905 -18.745 74.045 -18.575 ;
      RECT 73.955 -17.558 74.045 -16.55 ;
      RECT 73.905 -16.955 74.045 -16.785 ;
      RECT 73.955 -15.75 74.045 -14.742 ;
      RECT 73.905 -15.515 74.045 -15.345 ;
      RECT 73.955 -14.328 74.045 -13.32 ;
      RECT 73.905 -13.725 74.045 -13.555 ;
      RECT 73.955 -12.52 74.045 -11.512 ;
      RECT 73.905 -12.285 74.045 -12.115 ;
      RECT 73.955 -11.098 74.045 -10.09 ;
      RECT 73.905 -10.495 74.045 -10.325 ;
      RECT 73.955 -9.29 74.045 -8.282 ;
      RECT 73.905 -9.055 74.045 -8.885 ;
      RECT 73.955 -7.868 74.045 -6.86 ;
      RECT 73.905 -7.265 74.045 -7.095 ;
      RECT 73.955 -6.06 74.045 -5.052 ;
      RECT 73.905 -5.825 74.045 -5.655 ;
      RECT 73.955 -4.638 74.045 -3.63 ;
      RECT 73.905 -4.035 74.045 -3.865 ;
      RECT 73.955 -2.83 74.045 -1.822 ;
      RECT 73.905 -2.595 74.045 -2.425 ;
      RECT 73.955 -1.408 74.045 -0.4 ;
      RECT 73.905 -0.805 74.045 -0.635 ;
      RECT 73.955 0.4 74.045 1.408 ;
      RECT 73.905 0.635 74.045 0.805 ;
      RECT 73.83 -114.685 74.005 -114.515 ;
      RECT 73.905 -114.895 74.005 -114.515 ;
      RECT 72.945 -113.555 73.045 -113.09 ;
      RECT 73.31 -113.555 73.41 -113.1 ;
      RECT 72.945 -113.555 73.79 -113.385 ;
      RECT 73.555 -101.538 73.645 -100.531 ;
      RECT 73.555 -101.225 73.695 -101.055 ;
      RECT 73.555 -99.729 73.645 -98.722 ;
      RECT 73.555 -99.205 73.695 -99.035 ;
      RECT 73.555 -98.308 73.645 -97.301 ;
      RECT 73.555 -97.995 73.695 -97.825 ;
      RECT 73.555 -96.499 73.645 -95.492 ;
      RECT 73.555 -95.975 73.695 -95.805 ;
      RECT 73.555 -95.078 73.645 -94.071 ;
      RECT 73.555 -94.765 73.695 -94.595 ;
      RECT 73.555 -93.269 73.645 -92.262 ;
      RECT 73.555 -92.745 73.695 -92.575 ;
      RECT 73.555 -91.848 73.645 -90.841 ;
      RECT 73.555 -91.535 73.695 -91.365 ;
      RECT 73.555 -90.039 73.645 -89.032 ;
      RECT 73.555 -89.515 73.695 -89.345 ;
      RECT 73.555 -88.618 73.645 -87.611 ;
      RECT 73.555 -88.305 73.695 -88.135 ;
      RECT 73.555 -86.809 73.645 -85.802 ;
      RECT 73.555 -86.285 73.695 -86.115 ;
      RECT 73.555 -85.388 73.645 -84.381 ;
      RECT 73.555 -85.075 73.695 -84.905 ;
      RECT 73.555 -83.579 73.645 -82.572 ;
      RECT 73.555 -83.055 73.695 -82.885 ;
      RECT 73.555 -82.158 73.645 -81.151 ;
      RECT 73.555 -81.845 73.695 -81.675 ;
      RECT 73.555 -80.349 73.645 -79.342 ;
      RECT 73.555 -79.825 73.695 -79.655 ;
      RECT 73.555 -78.928 73.645 -77.921 ;
      RECT 73.555 -78.615 73.695 -78.445 ;
      RECT 73.555 -77.119 73.645 -76.112 ;
      RECT 73.555 -76.595 73.695 -76.425 ;
      RECT 73.555 -75.698 73.645 -74.691 ;
      RECT 73.555 -75.385 73.695 -75.215 ;
      RECT 73.555 -73.889 73.645 -72.882 ;
      RECT 73.555 -73.365 73.695 -73.195 ;
      RECT 73.555 -72.468 73.645 -71.461 ;
      RECT 73.555 -72.155 73.695 -71.985 ;
      RECT 73.555 -70.659 73.645 -69.652 ;
      RECT 73.555 -70.135 73.695 -69.965 ;
      RECT 73.555 -69.238 73.645 -68.231 ;
      RECT 73.555 -68.925 73.695 -68.755 ;
      RECT 73.555 -67.429 73.645 -66.422 ;
      RECT 73.555 -66.905 73.695 -66.735 ;
      RECT 73.555 -66.008 73.645 -65.001 ;
      RECT 73.555 -65.695 73.695 -65.525 ;
      RECT 73.555 -64.199 73.645 -63.192 ;
      RECT 73.555 -63.675 73.695 -63.505 ;
      RECT 73.555 -62.778 73.645 -61.771 ;
      RECT 73.555 -62.465 73.695 -62.295 ;
      RECT 73.555 -60.969 73.645 -59.962 ;
      RECT 73.555 -60.445 73.695 -60.275 ;
      RECT 73.555 -59.548 73.645 -58.541 ;
      RECT 73.555 -59.235 73.695 -59.065 ;
      RECT 73.555 -57.739 73.645 -56.732 ;
      RECT 73.555 -57.215 73.695 -57.045 ;
      RECT 73.555 -56.318 73.645 -55.311 ;
      RECT 73.555 -56.005 73.695 -55.835 ;
      RECT 73.555 -54.509 73.645 -53.502 ;
      RECT 73.555 -53.985 73.695 -53.815 ;
      RECT 73.555 -53.088 73.645 -52.081 ;
      RECT 73.555 -52.775 73.695 -52.605 ;
      RECT 73.555 -51.279 73.645 -50.272 ;
      RECT 73.555 -50.755 73.695 -50.585 ;
      RECT 73.555 -49.858 73.645 -48.851 ;
      RECT 73.555 -49.545 73.695 -49.375 ;
      RECT 73.555 -48.049 73.645 -47.042 ;
      RECT 73.555 -47.525 73.695 -47.355 ;
      RECT 73.555 -46.628 73.645 -45.621 ;
      RECT 73.555 -46.315 73.695 -46.145 ;
      RECT 73.555 -44.819 73.645 -43.812 ;
      RECT 73.555 -44.295 73.695 -44.125 ;
      RECT 73.555 -43.398 73.645 -42.391 ;
      RECT 73.555 -43.085 73.695 -42.915 ;
      RECT 73.555 -41.589 73.645 -40.582 ;
      RECT 73.555 -41.065 73.695 -40.895 ;
      RECT 73.555 -40.168 73.645 -39.161 ;
      RECT 73.555 -39.855 73.695 -39.685 ;
      RECT 73.555 -38.359 73.645 -37.352 ;
      RECT 73.555 -37.835 73.695 -37.665 ;
      RECT 73.555 -36.938 73.645 -35.931 ;
      RECT 73.555 -36.625 73.695 -36.455 ;
      RECT 73.555 -35.129 73.645 -34.122 ;
      RECT 73.555 -34.605 73.695 -34.435 ;
      RECT 73.555 -33.708 73.645 -32.701 ;
      RECT 73.555 -33.395 73.695 -33.225 ;
      RECT 73.555 -31.899 73.645 -30.892 ;
      RECT 73.555 -31.375 73.695 -31.205 ;
      RECT 73.555 -30.478 73.645 -29.471 ;
      RECT 73.555 -30.165 73.695 -29.995 ;
      RECT 73.555 -28.669 73.645 -27.662 ;
      RECT 73.555 -28.145 73.695 -27.975 ;
      RECT 73.555 -27.248 73.645 -26.241 ;
      RECT 73.555 -26.935 73.695 -26.765 ;
      RECT 73.555 -25.439 73.645 -24.432 ;
      RECT 73.555 -24.915 73.695 -24.745 ;
      RECT 73.555 -24.018 73.645 -23.011 ;
      RECT 73.555 -23.705 73.695 -23.535 ;
      RECT 73.555 -22.209 73.645 -21.202 ;
      RECT 73.555 -21.685 73.695 -21.515 ;
      RECT 73.555 -20.788 73.645 -19.781 ;
      RECT 73.555 -20.475 73.695 -20.305 ;
      RECT 73.555 -18.979 73.645 -17.972 ;
      RECT 73.555 -18.455 73.695 -18.285 ;
      RECT 73.555 -17.558 73.645 -16.551 ;
      RECT 73.555 -17.245 73.695 -17.075 ;
      RECT 73.555 -15.749 73.645 -14.742 ;
      RECT 73.555 -15.225 73.695 -15.055 ;
      RECT 73.555 -14.328 73.645 -13.321 ;
      RECT 73.555 -14.015 73.695 -13.845 ;
      RECT 73.555 -12.519 73.645 -11.512 ;
      RECT 73.555 -11.995 73.695 -11.825 ;
      RECT 73.555 -11.098 73.645 -10.091 ;
      RECT 73.555 -10.785 73.695 -10.615 ;
      RECT 73.555 -9.289 73.645 -8.282 ;
      RECT 73.555 -8.765 73.695 -8.595 ;
      RECT 73.555 -7.868 73.645 -6.861 ;
      RECT 73.555 -7.555 73.695 -7.385 ;
      RECT 73.555 -6.059 73.645 -5.052 ;
      RECT 73.555 -5.535 73.695 -5.365 ;
      RECT 73.555 -4.638 73.645 -3.631 ;
      RECT 73.555 -4.325 73.695 -4.155 ;
      RECT 73.555 -2.829 73.645 -1.822 ;
      RECT 73.555 -2.305 73.695 -2.135 ;
      RECT 73.555 -1.408 73.645 -0.401 ;
      RECT 73.555 -1.095 73.695 -0.925 ;
      RECT 73.555 0.401 73.645 1.408 ;
      RECT 73.555 0.925 73.695 1.095 ;
      RECT 73.24 -114.685 73.41 -114.515 ;
      RECT 73.31 -114.895 73.41 -114.515 ;
      RECT 72.755 -101.538 72.845 -100.53 ;
      RECT 72.705 -100.935 72.845 -100.765 ;
      RECT 72.755 -99.73 72.845 -98.722 ;
      RECT 72.705 -99.495 72.845 -99.325 ;
      RECT 72.755 -98.308 72.845 -97.3 ;
      RECT 72.705 -97.705 72.845 -97.535 ;
      RECT 72.755 -96.5 72.845 -95.492 ;
      RECT 72.705 -96.265 72.845 -96.095 ;
      RECT 72.755 -95.078 72.845 -94.07 ;
      RECT 72.705 -94.475 72.845 -94.305 ;
      RECT 72.755 -93.27 72.845 -92.262 ;
      RECT 72.705 -93.035 72.845 -92.865 ;
      RECT 72.755 -91.848 72.845 -90.84 ;
      RECT 72.705 -91.245 72.845 -91.075 ;
      RECT 72.755 -90.04 72.845 -89.032 ;
      RECT 72.705 -89.805 72.845 -89.635 ;
      RECT 72.755 -88.618 72.845 -87.61 ;
      RECT 72.705 -88.015 72.845 -87.845 ;
      RECT 72.755 -86.81 72.845 -85.802 ;
      RECT 72.705 -86.575 72.845 -86.405 ;
      RECT 72.755 -85.388 72.845 -84.38 ;
      RECT 72.705 -84.785 72.845 -84.615 ;
      RECT 72.755 -83.58 72.845 -82.572 ;
      RECT 72.705 -83.345 72.845 -83.175 ;
      RECT 72.755 -82.158 72.845 -81.15 ;
      RECT 72.705 -81.555 72.845 -81.385 ;
      RECT 72.755 -80.35 72.845 -79.342 ;
      RECT 72.705 -80.115 72.845 -79.945 ;
      RECT 72.755 -78.928 72.845 -77.92 ;
      RECT 72.705 -78.325 72.845 -78.155 ;
      RECT 72.755 -77.12 72.845 -76.112 ;
      RECT 72.705 -76.885 72.845 -76.715 ;
      RECT 72.755 -75.698 72.845 -74.69 ;
      RECT 72.705 -75.095 72.845 -74.925 ;
      RECT 72.755 -73.89 72.845 -72.882 ;
      RECT 72.705 -73.655 72.845 -73.485 ;
      RECT 72.755 -72.468 72.845 -71.46 ;
      RECT 72.705 -71.865 72.845 -71.695 ;
      RECT 72.755 -70.66 72.845 -69.652 ;
      RECT 72.705 -70.425 72.845 -70.255 ;
      RECT 72.755 -69.238 72.845 -68.23 ;
      RECT 72.705 -68.635 72.845 -68.465 ;
      RECT 72.755 -67.43 72.845 -66.422 ;
      RECT 72.705 -67.195 72.845 -67.025 ;
      RECT 72.755 -66.008 72.845 -65 ;
      RECT 72.705 -65.405 72.845 -65.235 ;
      RECT 72.755 -64.2 72.845 -63.192 ;
      RECT 72.705 -63.965 72.845 -63.795 ;
      RECT 72.755 -62.778 72.845 -61.77 ;
      RECT 72.705 -62.175 72.845 -62.005 ;
      RECT 72.755 -60.97 72.845 -59.962 ;
      RECT 72.705 -60.735 72.845 -60.565 ;
      RECT 72.755 -59.548 72.845 -58.54 ;
      RECT 72.705 -58.945 72.845 -58.775 ;
      RECT 72.755 -57.74 72.845 -56.732 ;
      RECT 72.705 -57.505 72.845 -57.335 ;
      RECT 72.755 -56.318 72.845 -55.31 ;
      RECT 72.705 -55.715 72.845 -55.545 ;
      RECT 72.755 -54.51 72.845 -53.502 ;
      RECT 72.705 -54.275 72.845 -54.105 ;
      RECT 72.755 -53.088 72.845 -52.08 ;
      RECT 72.705 -52.485 72.845 -52.315 ;
      RECT 72.755 -51.28 72.845 -50.272 ;
      RECT 72.705 -51.045 72.845 -50.875 ;
      RECT 72.755 -49.858 72.845 -48.85 ;
      RECT 72.705 -49.255 72.845 -49.085 ;
      RECT 72.755 -48.05 72.845 -47.042 ;
      RECT 72.705 -47.815 72.845 -47.645 ;
      RECT 72.755 -46.628 72.845 -45.62 ;
      RECT 72.705 -46.025 72.845 -45.855 ;
      RECT 72.755 -44.82 72.845 -43.812 ;
      RECT 72.705 -44.585 72.845 -44.415 ;
      RECT 72.755 -43.398 72.845 -42.39 ;
      RECT 72.705 -42.795 72.845 -42.625 ;
      RECT 72.755 -41.59 72.845 -40.582 ;
      RECT 72.705 -41.355 72.845 -41.185 ;
      RECT 72.755 -40.168 72.845 -39.16 ;
      RECT 72.705 -39.565 72.845 -39.395 ;
      RECT 72.755 -38.36 72.845 -37.352 ;
      RECT 72.705 -38.125 72.845 -37.955 ;
      RECT 72.755 -36.938 72.845 -35.93 ;
      RECT 72.705 -36.335 72.845 -36.165 ;
      RECT 72.755 -35.13 72.845 -34.122 ;
      RECT 72.705 -34.895 72.845 -34.725 ;
      RECT 72.755 -33.708 72.845 -32.7 ;
      RECT 72.705 -33.105 72.845 -32.935 ;
      RECT 72.755 -31.9 72.845 -30.892 ;
      RECT 72.705 -31.665 72.845 -31.495 ;
      RECT 72.755 -30.478 72.845 -29.47 ;
      RECT 72.705 -29.875 72.845 -29.705 ;
      RECT 72.755 -28.67 72.845 -27.662 ;
      RECT 72.705 -28.435 72.845 -28.265 ;
      RECT 72.755 -27.248 72.845 -26.24 ;
      RECT 72.705 -26.645 72.845 -26.475 ;
      RECT 72.755 -25.44 72.845 -24.432 ;
      RECT 72.705 -25.205 72.845 -25.035 ;
      RECT 72.755 -24.018 72.845 -23.01 ;
      RECT 72.705 -23.415 72.845 -23.245 ;
      RECT 72.755 -22.21 72.845 -21.202 ;
      RECT 72.705 -21.975 72.845 -21.805 ;
      RECT 72.755 -20.788 72.845 -19.78 ;
      RECT 72.705 -20.185 72.845 -20.015 ;
      RECT 72.755 -18.98 72.845 -17.972 ;
      RECT 72.705 -18.745 72.845 -18.575 ;
      RECT 72.755 -17.558 72.845 -16.55 ;
      RECT 72.705 -16.955 72.845 -16.785 ;
      RECT 72.755 -15.75 72.845 -14.742 ;
      RECT 72.705 -15.515 72.845 -15.345 ;
      RECT 72.755 -14.328 72.845 -13.32 ;
      RECT 72.705 -13.725 72.845 -13.555 ;
      RECT 72.755 -12.52 72.845 -11.512 ;
      RECT 72.705 -12.285 72.845 -12.115 ;
      RECT 72.755 -11.098 72.845 -10.09 ;
      RECT 72.705 -10.495 72.845 -10.325 ;
      RECT 72.755 -9.29 72.845 -8.282 ;
      RECT 72.705 -9.055 72.845 -8.885 ;
      RECT 72.755 -7.868 72.845 -6.86 ;
      RECT 72.705 -7.265 72.845 -7.095 ;
      RECT 72.755 -6.06 72.845 -5.052 ;
      RECT 72.705 -5.825 72.845 -5.655 ;
      RECT 72.755 -4.638 72.845 -3.63 ;
      RECT 72.705 -4.035 72.845 -3.865 ;
      RECT 72.755 -2.83 72.845 -1.822 ;
      RECT 72.705 -2.595 72.845 -2.425 ;
      RECT 72.755 -1.408 72.845 -0.4 ;
      RECT 72.705 -0.805 72.845 -0.635 ;
      RECT 72.755 0.4 72.845 1.408 ;
      RECT 72.705 0.635 72.845 0.805 ;
      RECT 72.355 -101.538 72.445 -100.531 ;
      RECT 72.355 -101.225 72.495 -101.055 ;
      RECT 72.355 -99.729 72.445 -98.722 ;
      RECT 72.355 -99.205 72.495 -99.035 ;
      RECT 72.355 -98.308 72.445 -97.301 ;
      RECT 72.355 -97.995 72.495 -97.825 ;
      RECT 72.355 -96.499 72.445 -95.492 ;
      RECT 72.355 -95.975 72.495 -95.805 ;
      RECT 72.355 -95.078 72.445 -94.071 ;
      RECT 72.355 -94.765 72.495 -94.595 ;
      RECT 72.355 -93.269 72.445 -92.262 ;
      RECT 72.355 -92.745 72.495 -92.575 ;
      RECT 72.355 -91.848 72.445 -90.841 ;
      RECT 72.355 -91.535 72.495 -91.365 ;
      RECT 72.355 -90.039 72.445 -89.032 ;
      RECT 72.355 -89.515 72.495 -89.345 ;
      RECT 72.355 -88.618 72.445 -87.611 ;
      RECT 72.355 -88.305 72.495 -88.135 ;
      RECT 72.355 -86.809 72.445 -85.802 ;
      RECT 72.355 -86.285 72.495 -86.115 ;
      RECT 72.355 -85.388 72.445 -84.381 ;
      RECT 72.355 -85.075 72.495 -84.905 ;
      RECT 72.355 -83.579 72.445 -82.572 ;
      RECT 72.355 -83.055 72.495 -82.885 ;
      RECT 72.355 -82.158 72.445 -81.151 ;
      RECT 72.355 -81.845 72.495 -81.675 ;
      RECT 72.355 -80.349 72.445 -79.342 ;
      RECT 72.355 -79.825 72.495 -79.655 ;
      RECT 72.355 -78.928 72.445 -77.921 ;
      RECT 72.355 -78.615 72.495 -78.445 ;
      RECT 72.355 -77.119 72.445 -76.112 ;
      RECT 72.355 -76.595 72.495 -76.425 ;
      RECT 72.355 -75.698 72.445 -74.691 ;
      RECT 72.355 -75.385 72.495 -75.215 ;
      RECT 72.355 -73.889 72.445 -72.882 ;
      RECT 72.355 -73.365 72.495 -73.195 ;
      RECT 72.355 -72.468 72.445 -71.461 ;
      RECT 72.355 -72.155 72.495 -71.985 ;
      RECT 72.355 -70.659 72.445 -69.652 ;
      RECT 72.355 -70.135 72.495 -69.965 ;
      RECT 72.355 -69.238 72.445 -68.231 ;
      RECT 72.355 -68.925 72.495 -68.755 ;
      RECT 72.355 -67.429 72.445 -66.422 ;
      RECT 72.355 -66.905 72.495 -66.735 ;
      RECT 72.355 -66.008 72.445 -65.001 ;
      RECT 72.355 -65.695 72.495 -65.525 ;
      RECT 72.355 -64.199 72.445 -63.192 ;
      RECT 72.355 -63.675 72.495 -63.505 ;
      RECT 72.355 -62.778 72.445 -61.771 ;
      RECT 72.355 -62.465 72.495 -62.295 ;
      RECT 72.355 -60.969 72.445 -59.962 ;
      RECT 72.355 -60.445 72.495 -60.275 ;
      RECT 72.355 -59.548 72.445 -58.541 ;
      RECT 72.355 -59.235 72.495 -59.065 ;
      RECT 72.355 -57.739 72.445 -56.732 ;
      RECT 72.355 -57.215 72.495 -57.045 ;
      RECT 72.355 -56.318 72.445 -55.311 ;
      RECT 72.355 -56.005 72.495 -55.835 ;
      RECT 72.355 -54.509 72.445 -53.502 ;
      RECT 72.355 -53.985 72.495 -53.815 ;
      RECT 72.355 -53.088 72.445 -52.081 ;
      RECT 72.355 -52.775 72.495 -52.605 ;
      RECT 72.355 -51.279 72.445 -50.272 ;
      RECT 72.355 -50.755 72.495 -50.585 ;
      RECT 72.355 -49.858 72.445 -48.851 ;
      RECT 72.355 -49.545 72.495 -49.375 ;
      RECT 72.355 -48.049 72.445 -47.042 ;
      RECT 72.355 -47.525 72.495 -47.355 ;
      RECT 72.355 -46.628 72.445 -45.621 ;
      RECT 72.355 -46.315 72.495 -46.145 ;
      RECT 72.355 -44.819 72.445 -43.812 ;
      RECT 72.355 -44.295 72.495 -44.125 ;
      RECT 72.355 -43.398 72.445 -42.391 ;
      RECT 72.355 -43.085 72.495 -42.915 ;
      RECT 72.355 -41.589 72.445 -40.582 ;
      RECT 72.355 -41.065 72.495 -40.895 ;
      RECT 72.355 -40.168 72.445 -39.161 ;
      RECT 72.355 -39.855 72.495 -39.685 ;
      RECT 72.355 -38.359 72.445 -37.352 ;
      RECT 72.355 -37.835 72.495 -37.665 ;
      RECT 72.355 -36.938 72.445 -35.931 ;
      RECT 72.355 -36.625 72.495 -36.455 ;
      RECT 72.355 -35.129 72.445 -34.122 ;
      RECT 72.355 -34.605 72.495 -34.435 ;
      RECT 72.355 -33.708 72.445 -32.701 ;
      RECT 72.355 -33.395 72.495 -33.225 ;
      RECT 72.355 -31.899 72.445 -30.892 ;
      RECT 72.355 -31.375 72.495 -31.205 ;
      RECT 72.355 -30.478 72.445 -29.471 ;
      RECT 72.355 -30.165 72.495 -29.995 ;
      RECT 72.355 -28.669 72.445 -27.662 ;
      RECT 72.355 -28.145 72.495 -27.975 ;
      RECT 72.355 -27.248 72.445 -26.241 ;
      RECT 72.355 -26.935 72.495 -26.765 ;
      RECT 72.355 -25.439 72.445 -24.432 ;
      RECT 72.355 -24.915 72.495 -24.745 ;
      RECT 72.355 -24.018 72.445 -23.011 ;
      RECT 72.355 -23.705 72.495 -23.535 ;
      RECT 72.355 -22.209 72.445 -21.202 ;
      RECT 72.355 -21.685 72.495 -21.515 ;
      RECT 72.355 -20.788 72.445 -19.781 ;
      RECT 72.355 -20.475 72.495 -20.305 ;
      RECT 72.355 -18.979 72.445 -17.972 ;
      RECT 72.355 -18.455 72.495 -18.285 ;
      RECT 72.355 -17.558 72.445 -16.551 ;
      RECT 72.355 -17.245 72.495 -17.075 ;
      RECT 72.355 -15.749 72.445 -14.742 ;
      RECT 72.355 -15.225 72.495 -15.055 ;
      RECT 72.355 -14.328 72.445 -13.321 ;
      RECT 72.355 -14.015 72.495 -13.845 ;
      RECT 72.355 -12.519 72.445 -11.512 ;
      RECT 72.355 -11.995 72.495 -11.825 ;
      RECT 72.355 -11.098 72.445 -10.091 ;
      RECT 72.355 -10.785 72.495 -10.615 ;
      RECT 72.355 -9.289 72.445 -8.282 ;
      RECT 72.355 -8.765 72.495 -8.595 ;
      RECT 72.355 -7.868 72.445 -6.861 ;
      RECT 72.355 -7.555 72.495 -7.385 ;
      RECT 72.355 -6.059 72.445 -5.052 ;
      RECT 72.355 -5.535 72.495 -5.365 ;
      RECT 72.355 -4.638 72.445 -3.631 ;
      RECT 72.355 -4.325 72.495 -4.155 ;
      RECT 72.355 -2.829 72.445 -1.822 ;
      RECT 72.355 -2.305 72.495 -2.135 ;
      RECT 72.355 -1.408 72.445 -0.401 ;
      RECT 72.355 -1.095 72.495 -0.925 ;
      RECT 72.355 0.401 72.445 1.408 ;
      RECT 72.355 0.925 72.495 1.095 ;
      RECT 68.185 -108.935 71.965 -108.815 ;
      RECT 69.505 -109.475 69.605 -108.815 ;
      RECT 68.945 -109.475 69.045 -108.815 ;
      RECT 68.385 -109.475 68.485 -108.815 ;
      RECT 71.555 -101.538 71.645 -100.53 ;
      RECT 71.505 -100.935 71.645 -100.765 ;
      RECT 71.555 -99.73 71.645 -98.722 ;
      RECT 71.505 -99.495 71.645 -99.325 ;
      RECT 71.555 -98.308 71.645 -97.3 ;
      RECT 71.505 -97.705 71.645 -97.535 ;
      RECT 71.555 -96.5 71.645 -95.492 ;
      RECT 71.505 -96.265 71.645 -96.095 ;
      RECT 71.555 -95.078 71.645 -94.07 ;
      RECT 71.505 -94.475 71.645 -94.305 ;
      RECT 71.555 -93.27 71.645 -92.262 ;
      RECT 71.505 -93.035 71.645 -92.865 ;
      RECT 71.555 -91.848 71.645 -90.84 ;
      RECT 71.505 -91.245 71.645 -91.075 ;
      RECT 71.555 -90.04 71.645 -89.032 ;
      RECT 71.505 -89.805 71.645 -89.635 ;
      RECT 71.555 -88.618 71.645 -87.61 ;
      RECT 71.505 -88.015 71.645 -87.845 ;
      RECT 71.555 -86.81 71.645 -85.802 ;
      RECT 71.505 -86.575 71.645 -86.405 ;
      RECT 71.555 -85.388 71.645 -84.38 ;
      RECT 71.505 -84.785 71.645 -84.615 ;
      RECT 71.555 -83.58 71.645 -82.572 ;
      RECT 71.505 -83.345 71.645 -83.175 ;
      RECT 71.555 -82.158 71.645 -81.15 ;
      RECT 71.505 -81.555 71.645 -81.385 ;
      RECT 71.555 -80.35 71.645 -79.342 ;
      RECT 71.505 -80.115 71.645 -79.945 ;
      RECT 71.555 -78.928 71.645 -77.92 ;
      RECT 71.505 -78.325 71.645 -78.155 ;
      RECT 71.555 -77.12 71.645 -76.112 ;
      RECT 71.505 -76.885 71.645 -76.715 ;
      RECT 71.555 -75.698 71.645 -74.69 ;
      RECT 71.505 -75.095 71.645 -74.925 ;
      RECT 71.555 -73.89 71.645 -72.882 ;
      RECT 71.505 -73.655 71.645 -73.485 ;
      RECT 71.555 -72.468 71.645 -71.46 ;
      RECT 71.505 -71.865 71.645 -71.695 ;
      RECT 71.555 -70.66 71.645 -69.652 ;
      RECT 71.505 -70.425 71.645 -70.255 ;
      RECT 71.555 -69.238 71.645 -68.23 ;
      RECT 71.505 -68.635 71.645 -68.465 ;
      RECT 71.555 -67.43 71.645 -66.422 ;
      RECT 71.505 -67.195 71.645 -67.025 ;
      RECT 71.555 -66.008 71.645 -65 ;
      RECT 71.505 -65.405 71.645 -65.235 ;
      RECT 71.555 -64.2 71.645 -63.192 ;
      RECT 71.505 -63.965 71.645 -63.795 ;
      RECT 71.555 -62.778 71.645 -61.77 ;
      RECT 71.505 -62.175 71.645 -62.005 ;
      RECT 71.555 -60.97 71.645 -59.962 ;
      RECT 71.505 -60.735 71.645 -60.565 ;
      RECT 71.555 -59.548 71.645 -58.54 ;
      RECT 71.505 -58.945 71.645 -58.775 ;
      RECT 71.555 -57.74 71.645 -56.732 ;
      RECT 71.505 -57.505 71.645 -57.335 ;
      RECT 71.555 -56.318 71.645 -55.31 ;
      RECT 71.505 -55.715 71.645 -55.545 ;
      RECT 71.555 -54.51 71.645 -53.502 ;
      RECT 71.505 -54.275 71.645 -54.105 ;
      RECT 71.555 -53.088 71.645 -52.08 ;
      RECT 71.505 -52.485 71.645 -52.315 ;
      RECT 71.555 -51.28 71.645 -50.272 ;
      RECT 71.505 -51.045 71.645 -50.875 ;
      RECT 71.555 -49.858 71.645 -48.85 ;
      RECT 71.505 -49.255 71.645 -49.085 ;
      RECT 71.555 -48.05 71.645 -47.042 ;
      RECT 71.505 -47.815 71.645 -47.645 ;
      RECT 71.555 -46.628 71.645 -45.62 ;
      RECT 71.505 -46.025 71.645 -45.855 ;
      RECT 71.555 -44.82 71.645 -43.812 ;
      RECT 71.505 -44.585 71.645 -44.415 ;
      RECT 71.555 -43.398 71.645 -42.39 ;
      RECT 71.505 -42.795 71.645 -42.625 ;
      RECT 71.555 -41.59 71.645 -40.582 ;
      RECT 71.505 -41.355 71.645 -41.185 ;
      RECT 71.555 -40.168 71.645 -39.16 ;
      RECT 71.505 -39.565 71.645 -39.395 ;
      RECT 71.555 -38.36 71.645 -37.352 ;
      RECT 71.505 -38.125 71.645 -37.955 ;
      RECT 71.555 -36.938 71.645 -35.93 ;
      RECT 71.505 -36.335 71.645 -36.165 ;
      RECT 71.555 -35.13 71.645 -34.122 ;
      RECT 71.505 -34.895 71.645 -34.725 ;
      RECT 71.555 -33.708 71.645 -32.7 ;
      RECT 71.505 -33.105 71.645 -32.935 ;
      RECT 71.555 -31.9 71.645 -30.892 ;
      RECT 71.505 -31.665 71.645 -31.495 ;
      RECT 71.555 -30.478 71.645 -29.47 ;
      RECT 71.505 -29.875 71.645 -29.705 ;
      RECT 71.555 -28.67 71.645 -27.662 ;
      RECT 71.505 -28.435 71.645 -28.265 ;
      RECT 71.555 -27.248 71.645 -26.24 ;
      RECT 71.505 -26.645 71.645 -26.475 ;
      RECT 71.555 -25.44 71.645 -24.432 ;
      RECT 71.505 -25.205 71.645 -25.035 ;
      RECT 71.555 -24.018 71.645 -23.01 ;
      RECT 71.505 -23.415 71.645 -23.245 ;
      RECT 71.555 -22.21 71.645 -21.202 ;
      RECT 71.505 -21.975 71.645 -21.805 ;
      RECT 71.555 -20.788 71.645 -19.78 ;
      RECT 71.505 -20.185 71.645 -20.015 ;
      RECT 71.555 -18.98 71.645 -17.972 ;
      RECT 71.505 -18.745 71.645 -18.575 ;
      RECT 71.555 -17.558 71.645 -16.55 ;
      RECT 71.505 -16.955 71.645 -16.785 ;
      RECT 71.555 -15.75 71.645 -14.742 ;
      RECT 71.505 -15.515 71.645 -15.345 ;
      RECT 71.555 -14.328 71.645 -13.32 ;
      RECT 71.505 -13.725 71.645 -13.555 ;
      RECT 71.555 -12.52 71.645 -11.512 ;
      RECT 71.505 -12.285 71.645 -12.115 ;
      RECT 71.555 -11.098 71.645 -10.09 ;
      RECT 71.505 -10.495 71.645 -10.325 ;
      RECT 71.555 -9.29 71.645 -8.282 ;
      RECT 71.505 -9.055 71.645 -8.885 ;
      RECT 71.555 -7.868 71.645 -6.86 ;
      RECT 71.505 -7.265 71.645 -7.095 ;
      RECT 71.555 -6.06 71.645 -5.052 ;
      RECT 71.505 -5.825 71.645 -5.655 ;
      RECT 71.555 -4.638 71.645 -3.63 ;
      RECT 71.505 -4.035 71.645 -3.865 ;
      RECT 71.555 -2.83 71.645 -1.822 ;
      RECT 71.505 -2.595 71.645 -2.425 ;
      RECT 71.555 -1.408 71.645 -0.4 ;
      RECT 71.505 -0.805 71.645 -0.635 ;
      RECT 71.555 0.4 71.645 1.408 ;
      RECT 71.505 0.635 71.645 0.805 ;
      RECT 70.125 -111.685 71.605 -111.585 ;
      RECT 70.125 -112.195 70.225 -111.585 ;
      RECT 70.345 -109.15 71.605 -109.05 ;
      RECT 71.505 -109.475 71.605 -109.05 ;
      RECT 70.945 -109.475 71.045 -109.05 ;
      RECT 70.385 -109.475 70.485 -109.05 ;
      RECT 71.155 -101.538 71.245 -100.531 ;
      RECT 71.155 -101.225 71.295 -101.055 ;
      RECT 71.155 -99.729 71.245 -98.722 ;
      RECT 71.155 -99.205 71.295 -99.035 ;
      RECT 71.155 -98.308 71.245 -97.301 ;
      RECT 71.155 -97.995 71.295 -97.825 ;
      RECT 71.155 -96.499 71.245 -95.492 ;
      RECT 71.155 -95.975 71.295 -95.805 ;
      RECT 71.155 -95.078 71.245 -94.071 ;
      RECT 71.155 -94.765 71.295 -94.595 ;
      RECT 71.155 -93.269 71.245 -92.262 ;
      RECT 71.155 -92.745 71.295 -92.575 ;
      RECT 71.155 -91.848 71.245 -90.841 ;
      RECT 71.155 -91.535 71.295 -91.365 ;
      RECT 71.155 -90.039 71.245 -89.032 ;
      RECT 71.155 -89.515 71.295 -89.345 ;
      RECT 71.155 -88.618 71.245 -87.611 ;
      RECT 71.155 -88.305 71.295 -88.135 ;
      RECT 71.155 -86.809 71.245 -85.802 ;
      RECT 71.155 -86.285 71.295 -86.115 ;
      RECT 71.155 -85.388 71.245 -84.381 ;
      RECT 71.155 -85.075 71.295 -84.905 ;
      RECT 71.155 -83.579 71.245 -82.572 ;
      RECT 71.155 -83.055 71.295 -82.885 ;
      RECT 71.155 -82.158 71.245 -81.151 ;
      RECT 71.155 -81.845 71.295 -81.675 ;
      RECT 71.155 -80.349 71.245 -79.342 ;
      RECT 71.155 -79.825 71.295 -79.655 ;
      RECT 71.155 -78.928 71.245 -77.921 ;
      RECT 71.155 -78.615 71.295 -78.445 ;
      RECT 71.155 -77.119 71.245 -76.112 ;
      RECT 71.155 -76.595 71.295 -76.425 ;
      RECT 71.155 -75.698 71.245 -74.691 ;
      RECT 71.155 -75.385 71.295 -75.215 ;
      RECT 71.155 -73.889 71.245 -72.882 ;
      RECT 71.155 -73.365 71.295 -73.195 ;
      RECT 71.155 -72.468 71.245 -71.461 ;
      RECT 71.155 -72.155 71.295 -71.985 ;
      RECT 71.155 -70.659 71.245 -69.652 ;
      RECT 71.155 -70.135 71.295 -69.965 ;
      RECT 71.155 -69.238 71.245 -68.231 ;
      RECT 71.155 -68.925 71.295 -68.755 ;
      RECT 71.155 -67.429 71.245 -66.422 ;
      RECT 71.155 -66.905 71.295 -66.735 ;
      RECT 71.155 -66.008 71.245 -65.001 ;
      RECT 71.155 -65.695 71.295 -65.525 ;
      RECT 71.155 -64.199 71.245 -63.192 ;
      RECT 71.155 -63.675 71.295 -63.505 ;
      RECT 71.155 -62.778 71.245 -61.771 ;
      RECT 71.155 -62.465 71.295 -62.295 ;
      RECT 71.155 -60.969 71.245 -59.962 ;
      RECT 71.155 -60.445 71.295 -60.275 ;
      RECT 71.155 -59.548 71.245 -58.541 ;
      RECT 71.155 -59.235 71.295 -59.065 ;
      RECT 71.155 -57.739 71.245 -56.732 ;
      RECT 71.155 -57.215 71.295 -57.045 ;
      RECT 71.155 -56.318 71.245 -55.311 ;
      RECT 71.155 -56.005 71.295 -55.835 ;
      RECT 71.155 -54.509 71.245 -53.502 ;
      RECT 71.155 -53.985 71.295 -53.815 ;
      RECT 71.155 -53.088 71.245 -52.081 ;
      RECT 71.155 -52.775 71.295 -52.605 ;
      RECT 71.155 -51.279 71.245 -50.272 ;
      RECT 71.155 -50.755 71.295 -50.585 ;
      RECT 71.155 -49.858 71.245 -48.851 ;
      RECT 71.155 -49.545 71.295 -49.375 ;
      RECT 71.155 -48.049 71.245 -47.042 ;
      RECT 71.155 -47.525 71.295 -47.355 ;
      RECT 71.155 -46.628 71.245 -45.621 ;
      RECT 71.155 -46.315 71.295 -46.145 ;
      RECT 71.155 -44.819 71.245 -43.812 ;
      RECT 71.155 -44.295 71.295 -44.125 ;
      RECT 71.155 -43.398 71.245 -42.391 ;
      RECT 71.155 -43.085 71.295 -42.915 ;
      RECT 71.155 -41.589 71.245 -40.582 ;
      RECT 71.155 -41.065 71.295 -40.895 ;
      RECT 71.155 -40.168 71.245 -39.161 ;
      RECT 71.155 -39.855 71.295 -39.685 ;
      RECT 71.155 -38.359 71.245 -37.352 ;
      RECT 71.155 -37.835 71.295 -37.665 ;
      RECT 71.155 -36.938 71.245 -35.931 ;
      RECT 71.155 -36.625 71.295 -36.455 ;
      RECT 71.155 -35.129 71.245 -34.122 ;
      RECT 71.155 -34.605 71.295 -34.435 ;
      RECT 71.155 -33.708 71.245 -32.701 ;
      RECT 71.155 -33.395 71.295 -33.225 ;
      RECT 71.155 -31.899 71.245 -30.892 ;
      RECT 71.155 -31.375 71.295 -31.205 ;
      RECT 71.155 -30.478 71.245 -29.471 ;
      RECT 71.155 -30.165 71.295 -29.995 ;
      RECT 71.155 -28.669 71.245 -27.662 ;
      RECT 71.155 -28.145 71.295 -27.975 ;
      RECT 71.155 -27.248 71.245 -26.241 ;
      RECT 71.155 -26.935 71.295 -26.765 ;
      RECT 71.155 -25.439 71.245 -24.432 ;
      RECT 71.155 -24.915 71.295 -24.745 ;
      RECT 71.155 -24.018 71.245 -23.011 ;
      RECT 71.155 -23.705 71.295 -23.535 ;
      RECT 71.155 -22.209 71.245 -21.202 ;
      RECT 71.155 -21.685 71.295 -21.515 ;
      RECT 71.155 -20.788 71.245 -19.781 ;
      RECT 71.155 -20.475 71.295 -20.305 ;
      RECT 71.155 -18.979 71.245 -17.972 ;
      RECT 71.155 -18.455 71.295 -18.285 ;
      RECT 71.155 -17.558 71.245 -16.551 ;
      RECT 71.155 -17.245 71.295 -17.075 ;
      RECT 71.155 -15.749 71.245 -14.742 ;
      RECT 71.155 -15.225 71.295 -15.055 ;
      RECT 71.155 -14.328 71.245 -13.321 ;
      RECT 71.155 -14.015 71.295 -13.845 ;
      RECT 71.155 -12.519 71.245 -11.512 ;
      RECT 71.155 -11.995 71.295 -11.825 ;
      RECT 71.155 -11.098 71.245 -10.091 ;
      RECT 71.155 -10.785 71.295 -10.615 ;
      RECT 71.155 -9.289 71.245 -8.282 ;
      RECT 71.155 -8.765 71.295 -8.595 ;
      RECT 71.155 -7.868 71.245 -6.861 ;
      RECT 71.155 -7.555 71.295 -7.385 ;
      RECT 71.155 -6.059 71.245 -5.052 ;
      RECT 71.155 -5.535 71.295 -5.365 ;
      RECT 71.155 -4.638 71.245 -3.631 ;
      RECT 71.155 -4.325 71.295 -4.155 ;
      RECT 71.155 -2.829 71.245 -1.822 ;
      RECT 71.155 -2.305 71.295 -2.135 ;
      RECT 71.155 -1.408 71.245 -0.401 ;
      RECT 71.155 -1.095 71.295 -0.925 ;
      RECT 71.155 0.401 71.245 1.408 ;
      RECT 71.155 0.925 71.295 1.095 ;
      RECT 70.485 -111.495 70.655 -111.385 ;
      RECT 67.335 -111.495 70.655 -111.395 ;
      RECT 70.355 -101.538 70.445 -100.53 ;
      RECT 70.305 -100.935 70.445 -100.765 ;
      RECT 70.355 -99.73 70.445 -98.722 ;
      RECT 70.305 -99.495 70.445 -99.325 ;
      RECT 70.355 -98.308 70.445 -97.3 ;
      RECT 70.305 -97.705 70.445 -97.535 ;
      RECT 70.355 -96.5 70.445 -95.492 ;
      RECT 70.305 -96.265 70.445 -96.095 ;
      RECT 70.355 -95.078 70.445 -94.07 ;
      RECT 70.305 -94.475 70.445 -94.305 ;
      RECT 70.355 -93.27 70.445 -92.262 ;
      RECT 70.305 -93.035 70.445 -92.865 ;
      RECT 70.355 -91.848 70.445 -90.84 ;
      RECT 70.305 -91.245 70.445 -91.075 ;
      RECT 70.355 -90.04 70.445 -89.032 ;
      RECT 70.305 -89.805 70.445 -89.635 ;
      RECT 70.355 -88.618 70.445 -87.61 ;
      RECT 70.305 -88.015 70.445 -87.845 ;
      RECT 70.355 -86.81 70.445 -85.802 ;
      RECT 70.305 -86.575 70.445 -86.405 ;
      RECT 70.355 -85.388 70.445 -84.38 ;
      RECT 70.305 -84.785 70.445 -84.615 ;
      RECT 70.355 -83.58 70.445 -82.572 ;
      RECT 70.305 -83.345 70.445 -83.175 ;
      RECT 70.355 -82.158 70.445 -81.15 ;
      RECT 70.305 -81.555 70.445 -81.385 ;
      RECT 70.355 -80.35 70.445 -79.342 ;
      RECT 70.305 -80.115 70.445 -79.945 ;
      RECT 70.355 -78.928 70.445 -77.92 ;
      RECT 70.305 -78.325 70.445 -78.155 ;
      RECT 70.355 -77.12 70.445 -76.112 ;
      RECT 70.305 -76.885 70.445 -76.715 ;
      RECT 70.355 -75.698 70.445 -74.69 ;
      RECT 70.305 -75.095 70.445 -74.925 ;
      RECT 70.355 -73.89 70.445 -72.882 ;
      RECT 70.305 -73.655 70.445 -73.485 ;
      RECT 70.355 -72.468 70.445 -71.46 ;
      RECT 70.305 -71.865 70.445 -71.695 ;
      RECT 70.355 -70.66 70.445 -69.652 ;
      RECT 70.305 -70.425 70.445 -70.255 ;
      RECT 70.355 -69.238 70.445 -68.23 ;
      RECT 70.305 -68.635 70.445 -68.465 ;
      RECT 70.355 -67.43 70.445 -66.422 ;
      RECT 70.305 -67.195 70.445 -67.025 ;
      RECT 70.355 -66.008 70.445 -65 ;
      RECT 70.305 -65.405 70.445 -65.235 ;
      RECT 70.355 -64.2 70.445 -63.192 ;
      RECT 70.305 -63.965 70.445 -63.795 ;
      RECT 70.355 -62.778 70.445 -61.77 ;
      RECT 70.305 -62.175 70.445 -62.005 ;
      RECT 70.355 -60.97 70.445 -59.962 ;
      RECT 70.305 -60.735 70.445 -60.565 ;
      RECT 70.355 -59.548 70.445 -58.54 ;
      RECT 70.305 -58.945 70.445 -58.775 ;
      RECT 70.355 -57.74 70.445 -56.732 ;
      RECT 70.305 -57.505 70.445 -57.335 ;
      RECT 70.355 -56.318 70.445 -55.31 ;
      RECT 70.305 -55.715 70.445 -55.545 ;
      RECT 70.355 -54.51 70.445 -53.502 ;
      RECT 70.305 -54.275 70.445 -54.105 ;
      RECT 70.355 -53.088 70.445 -52.08 ;
      RECT 70.305 -52.485 70.445 -52.315 ;
      RECT 70.355 -51.28 70.445 -50.272 ;
      RECT 70.305 -51.045 70.445 -50.875 ;
      RECT 70.355 -49.858 70.445 -48.85 ;
      RECT 70.305 -49.255 70.445 -49.085 ;
      RECT 70.355 -48.05 70.445 -47.042 ;
      RECT 70.305 -47.815 70.445 -47.645 ;
      RECT 70.355 -46.628 70.445 -45.62 ;
      RECT 70.305 -46.025 70.445 -45.855 ;
      RECT 70.355 -44.82 70.445 -43.812 ;
      RECT 70.305 -44.585 70.445 -44.415 ;
      RECT 70.355 -43.398 70.445 -42.39 ;
      RECT 70.305 -42.795 70.445 -42.625 ;
      RECT 70.355 -41.59 70.445 -40.582 ;
      RECT 70.305 -41.355 70.445 -41.185 ;
      RECT 70.355 -40.168 70.445 -39.16 ;
      RECT 70.305 -39.565 70.445 -39.395 ;
      RECT 70.355 -38.36 70.445 -37.352 ;
      RECT 70.305 -38.125 70.445 -37.955 ;
      RECT 70.355 -36.938 70.445 -35.93 ;
      RECT 70.305 -36.335 70.445 -36.165 ;
      RECT 70.355 -35.13 70.445 -34.122 ;
      RECT 70.305 -34.895 70.445 -34.725 ;
      RECT 70.355 -33.708 70.445 -32.7 ;
      RECT 70.305 -33.105 70.445 -32.935 ;
      RECT 70.355 -31.9 70.445 -30.892 ;
      RECT 70.305 -31.665 70.445 -31.495 ;
      RECT 70.355 -30.478 70.445 -29.47 ;
      RECT 70.305 -29.875 70.445 -29.705 ;
      RECT 70.355 -28.67 70.445 -27.662 ;
      RECT 70.305 -28.435 70.445 -28.265 ;
      RECT 70.355 -27.248 70.445 -26.24 ;
      RECT 70.305 -26.645 70.445 -26.475 ;
      RECT 70.355 -25.44 70.445 -24.432 ;
      RECT 70.305 -25.205 70.445 -25.035 ;
      RECT 70.355 -24.018 70.445 -23.01 ;
      RECT 70.305 -23.415 70.445 -23.245 ;
      RECT 70.355 -22.21 70.445 -21.202 ;
      RECT 70.305 -21.975 70.445 -21.805 ;
      RECT 70.355 -20.788 70.445 -19.78 ;
      RECT 70.305 -20.185 70.445 -20.015 ;
      RECT 70.355 -18.98 70.445 -17.972 ;
      RECT 70.305 -18.745 70.445 -18.575 ;
      RECT 70.355 -17.558 70.445 -16.55 ;
      RECT 70.305 -16.955 70.445 -16.785 ;
      RECT 70.355 -15.75 70.445 -14.742 ;
      RECT 70.305 -15.515 70.445 -15.345 ;
      RECT 70.355 -14.328 70.445 -13.32 ;
      RECT 70.305 -13.725 70.445 -13.555 ;
      RECT 70.355 -12.52 70.445 -11.512 ;
      RECT 70.305 -12.285 70.445 -12.115 ;
      RECT 70.355 -11.098 70.445 -10.09 ;
      RECT 70.305 -10.495 70.445 -10.325 ;
      RECT 70.355 -9.29 70.445 -8.282 ;
      RECT 70.305 -9.055 70.445 -8.885 ;
      RECT 70.355 -7.868 70.445 -6.86 ;
      RECT 70.305 -7.265 70.445 -7.095 ;
      RECT 70.355 -6.06 70.445 -5.052 ;
      RECT 70.305 -5.825 70.445 -5.655 ;
      RECT 70.355 -4.638 70.445 -3.63 ;
      RECT 70.305 -4.035 70.445 -3.865 ;
      RECT 70.355 -2.83 70.445 -1.822 ;
      RECT 70.305 -2.595 70.445 -2.425 ;
      RECT 70.355 -1.408 70.445 -0.4 ;
      RECT 70.305 -0.805 70.445 -0.635 ;
      RECT 70.355 0.4 70.445 1.408 ;
      RECT 70.305 0.635 70.445 0.805 ;
      RECT 69.955 -101.538 70.045 -100.531 ;
      RECT 69.955 -101.225 70.095 -101.055 ;
      RECT 69.955 -99.729 70.045 -98.722 ;
      RECT 69.955 -99.205 70.095 -99.035 ;
      RECT 69.955 -98.308 70.045 -97.301 ;
      RECT 69.955 -97.995 70.095 -97.825 ;
      RECT 69.955 -96.499 70.045 -95.492 ;
      RECT 69.955 -95.975 70.095 -95.805 ;
      RECT 69.955 -95.078 70.045 -94.071 ;
      RECT 69.955 -94.765 70.095 -94.595 ;
      RECT 69.955 -93.269 70.045 -92.262 ;
      RECT 69.955 -92.745 70.095 -92.575 ;
      RECT 69.955 -91.848 70.045 -90.841 ;
      RECT 69.955 -91.535 70.095 -91.365 ;
      RECT 69.955 -90.039 70.045 -89.032 ;
      RECT 69.955 -89.515 70.095 -89.345 ;
      RECT 69.955 -88.618 70.045 -87.611 ;
      RECT 69.955 -88.305 70.095 -88.135 ;
      RECT 69.955 -86.809 70.045 -85.802 ;
      RECT 69.955 -86.285 70.095 -86.115 ;
      RECT 69.955 -85.388 70.045 -84.381 ;
      RECT 69.955 -85.075 70.095 -84.905 ;
      RECT 69.955 -83.579 70.045 -82.572 ;
      RECT 69.955 -83.055 70.095 -82.885 ;
      RECT 69.955 -82.158 70.045 -81.151 ;
      RECT 69.955 -81.845 70.095 -81.675 ;
      RECT 69.955 -80.349 70.045 -79.342 ;
      RECT 69.955 -79.825 70.095 -79.655 ;
      RECT 69.955 -78.928 70.045 -77.921 ;
      RECT 69.955 -78.615 70.095 -78.445 ;
      RECT 69.955 -77.119 70.045 -76.112 ;
      RECT 69.955 -76.595 70.095 -76.425 ;
      RECT 69.955 -75.698 70.045 -74.691 ;
      RECT 69.955 -75.385 70.095 -75.215 ;
      RECT 69.955 -73.889 70.045 -72.882 ;
      RECT 69.955 -73.365 70.095 -73.195 ;
      RECT 69.955 -72.468 70.045 -71.461 ;
      RECT 69.955 -72.155 70.095 -71.985 ;
      RECT 69.955 -70.659 70.045 -69.652 ;
      RECT 69.955 -70.135 70.095 -69.965 ;
      RECT 69.955 -69.238 70.045 -68.231 ;
      RECT 69.955 -68.925 70.095 -68.755 ;
      RECT 69.955 -67.429 70.045 -66.422 ;
      RECT 69.955 -66.905 70.095 -66.735 ;
      RECT 69.955 -66.008 70.045 -65.001 ;
      RECT 69.955 -65.695 70.095 -65.525 ;
      RECT 69.955 -64.199 70.045 -63.192 ;
      RECT 69.955 -63.675 70.095 -63.505 ;
      RECT 69.955 -62.778 70.045 -61.771 ;
      RECT 69.955 -62.465 70.095 -62.295 ;
      RECT 69.955 -60.969 70.045 -59.962 ;
      RECT 69.955 -60.445 70.095 -60.275 ;
      RECT 69.955 -59.548 70.045 -58.541 ;
      RECT 69.955 -59.235 70.095 -59.065 ;
      RECT 69.955 -57.739 70.045 -56.732 ;
      RECT 69.955 -57.215 70.095 -57.045 ;
      RECT 69.955 -56.318 70.045 -55.311 ;
      RECT 69.955 -56.005 70.095 -55.835 ;
      RECT 69.955 -54.509 70.045 -53.502 ;
      RECT 69.955 -53.985 70.095 -53.815 ;
      RECT 69.955 -53.088 70.045 -52.081 ;
      RECT 69.955 -52.775 70.095 -52.605 ;
      RECT 69.955 -51.279 70.045 -50.272 ;
      RECT 69.955 -50.755 70.095 -50.585 ;
      RECT 69.955 -49.858 70.045 -48.851 ;
      RECT 69.955 -49.545 70.095 -49.375 ;
      RECT 69.955 -48.049 70.045 -47.042 ;
      RECT 69.955 -47.525 70.095 -47.355 ;
      RECT 69.955 -46.628 70.045 -45.621 ;
      RECT 69.955 -46.315 70.095 -46.145 ;
      RECT 69.955 -44.819 70.045 -43.812 ;
      RECT 69.955 -44.295 70.095 -44.125 ;
      RECT 69.955 -43.398 70.045 -42.391 ;
      RECT 69.955 -43.085 70.095 -42.915 ;
      RECT 69.955 -41.589 70.045 -40.582 ;
      RECT 69.955 -41.065 70.095 -40.895 ;
      RECT 69.955 -40.168 70.045 -39.161 ;
      RECT 69.955 -39.855 70.095 -39.685 ;
      RECT 69.955 -38.359 70.045 -37.352 ;
      RECT 69.955 -37.835 70.095 -37.665 ;
      RECT 69.955 -36.938 70.045 -35.931 ;
      RECT 69.955 -36.625 70.095 -36.455 ;
      RECT 69.955 -35.129 70.045 -34.122 ;
      RECT 69.955 -34.605 70.095 -34.435 ;
      RECT 69.955 -33.708 70.045 -32.701 ;
      RECT 69.955 -33.395 70.095 -33.225 ;
      RECT 69.955 -31.899 70.045 -30.892 ;
      RECT 69.955 -31.375 70.095 -31.205 ;
      RECT 69.955 -30.478 70.045 -29.471 ;
      RECT 69.955 -30.165 70.095 -29.995 ;
      RECT 69.955 -28.669 70.045 -27.662 ;
      RECT 69.955 -28.145 70.095 -27.975 ;
      RECT 69.955 -27.248 70.045 -26.241 ;
      RECT 69.955 -26.935 70.095 -26.765 ;
      RECT 69.955 -25.439 70.045 -24.432 ;
      RECT 69.955 -24.915 70.095 -24.745 ;
      RECT 69.955 -24.018 70.045 -23.011 ;
      RECT 69.955 -23.705 70.095 -23.535 ;
      RECT 69.955 -22.209 70.045 -21.202 ;
      RECT 69.955 -21.685 70.095 -21.515 ;
      RECT 69.955 -20.788 70.045 -19.781 ;
      RECT 69.955 -20.475 70.095 -20.305 ;
      RECT 69.955 -18.979 70.045 -17.972 ;
      RECT 69.955 -18.455 70.095 -18.285 ;
      RECT 69.955 -17.558 70.045 -16.551 ;
      RECT 69.955 -17.245 70.095 -17.075 ;
      RECT 69.955 -15.749 70.045 -14.742 ;
      RECT 69.955 -15.225 70.095 -15.055 ;
      RECT 69.955 -14.328 70.045 -13.321 ;
      RECT 69.955 -14.015 70.095 -13.845 ;
      RECT 69.955 -12.519 70.045 -11.512 ;
      RECT 69.955 -11.995 70.095 -11.825 ;
      RECT 69.955 -11.098 70.045 -10.091 ;
      RECT 69.955 -10.785 70.095 -10.615 ;
      RECT 69.955 -9.289 70.045 -8.282 ;
      RECT 69.955 -8.765 70.095 -8.595 ;
      RECT 69.955 -7.868 70.045 -6.861 ;
      RECT 69.955 -7.555 70.095 -7.385 ;
      RECT 69.955 -6.059 70.045 -5.052 ;
      RECT 69.955 -5.535 70.095 -5.365 ;
      RECT 69.955 -4.638 70.045 -3.631 ;
      RECT 69.955 -4.325 70.095 -4.155 ;
      RECT 69.955 -2.829 70.045 -1.822 ;
      RECT 69.955 -2.305 70.095 -2.135 ;
      RECT 69.955 -1.408 70.045 -0.401 ;
      RECT 69.955 -1.095 70.095 -0.925 ;
      RECT 69.955 0.401 70.045 1.408 ;
      RECT 69.955 0.925 70.095 1.095 ;
      RECT 68.105 -111.685 69.585 -111.585 ;
      RECT 68.105 -112.055 68.205 -111.585 ;
      RECT 67.91 -114.395 69.485 -114.275 ;
      RECT 69.385 -114.895 69.485 -114.275 ;
      RECT 68.79 -114.895 68.89 -114.275 ;
      RECT 67.91 -114.85 68.01 -114.275 ;
      RECT 69.155 -101.538 69.245 -100.53 ;
      RECT 69.105 -100.935 69.245 -100.765 ;
      RECT 69.155 -99.73 69.245 -98.722 ;
      RECT 69.105 -99.495 69.245 -99.325 ;
      RECT 69.155 -98.308 69.245 -97.3 ;
      RECT 69.105 -97.705 69.245 -97.535 ;
      RECT 69.155 -96.5 69.245 -95.492 ;
      RECT 69.105 -96.265 69.245 -96.095 ;
      RECT 69.155 -95.078 69.245 -94.07 ;
      RECT 69.105 -94.475 69.245 -94.305 ;
      RECT 69.155 -93.27 69.245 -92.262 ;
      RECT 69.105 -93.035 69.245 -92.865 ;
      RECT 69.155 -91.848 69.245 -90.84 ;
      RECT 69.105 -91.245 69.245 -91.075 ;
      RECT 69.155 -90.04 69.245 -89.032 ;
      RECT 69.105 -89.805 69.245 -89.635 ;
      RECT 69.155 -88.618 69.245 -87.61 ;
      RECT 69.105 -88.015 69.245 -87.845 ;
      RECT 69.155 -86.81 69.245 -85.802 ;
      RECT 69.105 -86.575 69.245 -86.405 ;
      RECT 69.155 -85.388 69.245 -84.38 ;
      RECT 69.105 -84.785 69.245 -84.615 ;
      RECT 69.155 -83.58 69.245 -82.572 ;
      RECT 69.105 -83.345 69.245 -83.175 ;
      RECT 69.155 -82.158 69.245 -81.15 ;
      RECT 69.105 -81.555 69.245 -81.385 ;
      RECT 69.155 -80.35 69.245 -79.342 ;
      RECT 69.105 -80.115 69.245 -79.945 ;
      RECT 69.155 -78.928 69.245 -77.92 ;
      RECT 69.105 -78.325 69.245 -78.155 ;
      RECT 69.155 -77.12 69.245 -76.112 ;
      RECT 69.105 -76.885 69.245 -76.715 ;
      RECT 69.155 -75.698 69.245 -74.69 ;
      RECT 69.105 -75.095 69.245 -74.925 ;
      RECT 69.155 -73.89 69.245 -72.882 ;
      RECT 69.105 -73.655 69.245 -73.485 ;
      RECT 69.155 -72.468 69.245 -71.46 ;
      RECT 69.105 -71.865 69.245 -71.695 ;
      RECT 69.155 -70.66 69.245 -69.652 ;
      RECT 69.105 -70.425 69.245 -70.255 ;
      RECT 69.155 -69.238 69.245 -68.23 ;
      RECT 69.105 -68.635 69.245 -68.465 ;
      RECT 69.155 -67.43 69.245 -66.422 ;
      RECT 69.105 -67.195 69.245 -67.025 ;
      RECT 69.155 -66.008 69.245 -65 ;
      RECT 69.105 -65.405 69.245 -65.235 ;
      RECT 69.155 -64.2 69.245 -63.192 ;
      RECT 69.105 -63.965 69.245 -63.795 ;
      RECT 69.155 -62.778 69.245 -61.77 ;
      RECT 69.105 -62.175 69.245 -62.005 ;
      RECT 69.155 -60.97 69.245 -59.962 ;
      RECT 69.105 -60.735 69.245 -60.565 ;
      RECT 69.155 -59.548 69.245 -58.54 ;
      RECT 69.105 -58.945 69.245 -58.775 ;
      RECT 69.155 -57.74 69.245 -56.732 ;
      RECT 69.105 -57.505 69.245 -57.335 ;
      RECT 69.155 -56.318 69.245 -55.31 ;
      RECT 69.105 -55.715 69.245 -55.545 ;
      RECT 69.155 -54.51 69.245 -53.502 ;
      RECT 69.105 -54.275 69.245 -54.105 ;
      RECT 69.155 -53.088 69.245 -52.08 ;
      RECT 69.105 -52.485 69.245 -52.315 ;
      RECT 69.155 -51.28 69.245 -50.272 ;
      RECT 69.105 -51.045 69.245 -50.875 ;
      RECT 69.155 -49.858 69.245 -48.85 ;
      RECT 69.105 -49.255 69.245 -49.085 ;
      RECT 69.155 -48.05 69.245 -47.042 ;
      RECT 69.105 -47.815 69.245 -47.645 ;
      RECT 69.155 -46.628 69.245 -45.62 ;
      RECT 69.105 -46.025 69.245 -45.855 ;
      RECT 69.155 -44.82 69.245 -43.812 ;
      RECT 69.105 -44.585 69.245 -44.415 ;
      RECT 69.155 -43.398 69.245 -42.39 ;
      RECT 69.105 -42.795 69.245 -42.625 ;
      RECT 69.155 -41.59 69.245 -40.582 ;
      RECT 69.105 -41.355 69.245 -41.185 ;
      RECT 69.155 -40.168 69.245 -39.16 ;
      RECT 69.105 -39.565 69.245 -39.395 ;
      RECT 69.155 -38.36 69.245 -37.352 ;
      RECT 69.105 -38.125 69.245 -37.955 ;
      RECT 69.155 -36.938 69.245 -35.93 ;
      RECT 69.105 -36.335 69.245 -36.165 ;
      RECT 69.155 -35.13 69.245 -34.122 ;
      RECT 69.105 -34.895 69.245 -34.725 ;
      RECT 69.155 -33.708 69.245 -32.7 ;
      RECT 69.105 -33.105 69.245 -32.935 ;
      RECT 69.155 -31.9 69.245 -30.892 ;
      RECT 69.105 -31.665 69.245 -31.495 ;
      RECT 69.155 -30.478 69.245 -29.47 ;
      RECT 69.105 -29.875 69.245 -29.705 ;
      RECT 69.155 -28.67 69.245 -27.662 ;
      RECT 69.105 -28.435 69.245 -28.265 ;
      RECT 69.155 -27.248 69.245 -26.24 ;
      RECT 69.105 -26.645 69.245 -26.475 ;
      RECT 69.155 -25.44 69.245 -24.432 ;
      RECT 69.105 -25.205 69.245 -25.035 ;
      RECT 69.155 -24.018 69.245 -23.01 ;
      RECT 69.105 -23.415 69.245 -23.245 ;
      RECT 69.155 -22.21 69.245 -21.202 ;
      RECT 69.105 -21.975 69.245 -21.805 ;
      RECT 69.155 -20.788 69.245 -19.78 ;
      RECT 69.105 -20.185 69.245 -20.015 ;
      RECT 69.155 -18.98 69.245 -17.972 ;
      RECT 69.105 -18.745 69.245 -18.575 ;
      RECT 69.155 -17.558 69.245 -16.55 ;
      RECT 69.105 -16.955 69.245 -16.785 ;
      RECT 69.155 -15.75 69.245 -14.742 ;
      RECT 69.105 -15.515 69.245 -15.345 ;
      RECT 69.155 -14.328 69.245 -13.32 ;
      RECT 69.105 -13.725 69.245 -13.555 ;
      RECT 69.155 -12.52 69.245 -11.512 ;
      RECT 69.105 -12.285 69.245 -12.115 ;
      RECT 69.155 -11.098 69.245 -10.09 ;
      RECT 69.105 -10.495 69.245 -10.325 ;
      RECT 69.155 -9.29 69.245 -8.282 ;
      RECT 69.105 -9.055 69.245 -8.885 ;
      RECT 69.155 -7.868 69.245 -6.86 ;
      RECT 69.105 -7.265 69.245 -7.095 ;
      RECT 69.155 -6.06 69.245 -5.052 ;
      RECT 69.105 -5.825 69.245 -5.655 ;
      RECT 69.155 -4.638 69.245 -3.63 ;
      RECT 69.105 -4.035 69.245 -3.865 ;
      RECT 69.155 -2.83 69.245 -1.822 ;
      RECT 69.105 -2.595 69.245 -2.425 ;
      RECT 69.155 -1.408 69.245 -0.4 ;
      RECT 69.105 -0.805 69.245 -0.635 ;
      RECT 69.155 0.4 69.245 1.408 ;
      RECT 69.105 0.635 69.245 0.805 ;
      RECT 69.03 -114.685 69.205 -114.515 ;
      RECT 69.105 -114.895 69.205 -114.515 ;
      RECT 68.145 -113.555 68.245 -113.09 ;
      RECT 68.51 -113.555 68.61 -113.1 ;
      RECT 68.145 -113.555 68.99 -113.385 ;
      RECT 68.755 -101.538 68.845 -100.531 ;
      RECT 68.755 -101.225 68.895 -101.055 ;
      RECT 68.755 -99.729 68.845 -98.722 ;
      RECT 68.755 -99.205 68.895 -99.035 ;
      RECT 68.755 -98.308 68.845 -97.301 ;
      RECT 68.755 -97.995 68.895 -97.825 ;
      RECT 68.755 -96.499 68.845 -95.492 ;
      RECT 68.755 -95.975 68.895 -95.805 ;
      RECT 68.755 -95.078 68.845 -94.071 ;
      RECT 68.755 -94.765 68.895 -94.595 ;
      RECT 68.755 -93.269 68.845 -92.262 ;
      RECT 68.755 -92.745 68.895 -92.575 ;
      RECT 68.755 -91.848 68.845 -90.841 ;
      RECT 68.755 -91.535 68.895 -91.365 ;
      RECT 68.755 -90.039 68.845 -89.032 ;
      RECT 68.755 -89.515 68.895 -89.345 ;
      RECT 68.755 -88.618 68.845 -87.611 ;
      RECT 68.755 -88.305 68.895 -88.135 ;
      RECT 68.755 -86.809 68.845 -85.802 ;
      RECT 68.755 -86.285 68.895 -86.115 ;
      RECT 68.755 -85.388 68.845 -84.381 ;
      RECT 68.755 -85.075 68.895 -84.905 ;
      RECT 68.755 -83.579 68.845 -82.572 ;
      RECT 68.755 -83.055 68.895 -82.885 ;
      RECT 68.755 -82.158 68.845 -81.151 ;
      RECT 68.755 -81.845 68.895 -81.675 ;
      RECT 68.755 -80.349 68.845 -79.342 ;
      RECT 68.755 -79.825 68.895 -79.655 ;
      RECT 68.755 -78.928 68.845 -77.921 ;
      RECT 68.755 -78.615 68.895 -78.445 ;
      RECT 68.755 -77.119 68.845 -76.112 ;
      RECT 68.755 -76.595 68.895 -76.425 ;
      RECT 68.755 -75.698 68.845 -74.691 ;
      RECT 68.755 -75.385 68.895 -75.215 ;
      RECT 68.755 -73.889 68.845 -72.882 ;
      RECT 68.755 -73.365 68.895 -73.195 ;
      RECT 68.755 -72.468 68.845 -71.461 ;
      RECT 68.755 -72.155 68.895 -71.985 ;
      RECT 68.755 -70.659 68.845 -69.652 ;
      RECT 68.755 -70.135 68.895 -69.965 ;
      RECT 68.755 -69.238 68.845 -68.231 ;
      RECT 68.755 -68.925 68.895 -68.755 ;
      RECT 68.755 -67.429 68.845 -66.422 ;
      RECT 68.755 -66.905 68.895 -66.735 ;
      RECT 68.755 -66.008 68.845 -65.001 ;
      RECT 68.755 -65.695 68.895 -65.525 ;
      RECT 68.755 -64.199 68.845 -63.192 ;
      RECT 68.755 -63.675 68.895 -63.505 ;
      RECT 68.755 -62.778 68.845 -61.771 ;
      RECT 68.755 -62.465 68.895 -62.295 ;
      RECT 68.755 -60.969 68.845 -59.962 ;
      RECT 68.755 -60.445 68.895 -60.275 ;
      RECT 68.755 -59.548 68.845 -58.541 ;
      RECT 68.755 -59.235 68.895 -59.065 ;
      RECT 68.755 -57.739 68.845 -56.732 ;
      RECT 68.755 -57.215 68.895 -57.045 ;
      RECT 68.755 -56.318 68.845 -55.311 ;
      RECT 68.755 -56.005 68.895 -55.835 ;
      RECT 68.755 -54.509 68.845 -53.502 ;
      RECT 68.755 -53.985 68.895 -53.815 ;
      RECT 68.755 -53.088 68.845 -52.081 ;
      RECT 68.755 -52.775 68.895 -52.605 ;
      RECT 68.755 -51.279 68.845 -50.272 ;
      RECT 68.755 -50.755 68.895 -50.585 ;
      RECT 68.755 -49.858 68.845 -48.851 ;
      RECT 68.755 -49.545 68.895 -49.375 ;
      RECT 68.755 -48.049 68.845 -47.042 ;
      RECT 68.755 -47.525 68.895 -47.355 ;
      RECT 68.755 -46.628 68.845 -45.621 ;
      RECT 68.755 -46.315 68.895 -46.145 ;
      RECT 68.755 -44.819 68.845 -43.812 ;
      RECT 68.755 -44.295 68.895 -44.125 ;
      RECT 68.755 -43.398 68.845 -42.391 ;
      RECT 68.755 -43.085 68.895 -42.915 ;
      RECT 68.755 -41.589 68.845 -40.582 ;
      RECT 68.755 -41.065 68.895 -40.895 ;
      RECT 68.755 -40.168 68.845 -39.161 ;
      RECT 68.755 -39.855 68.895 -39.685 ;
      RECT 68.755 -38.359 68.845 -37.352 ;
      RECT 68.755 -37.835 68.895 -37.665 ;
      RECT 68.755 -36.938 68.845 -35.931 ;
      RECT 68.755 -36.625 68.895 -36.455 ;
      RECT 68.755 -35.129 68.845 -34.122 ;
      RECT 68.755 -34.605 68.895 -34.435 ;
      RECT 68.755 -33.708 68.845 -32.701 ;
      RECT 68.755 -33.395 68.895 -33.225 ;
      RECT 68.755 -31.899 68.845 -30.892 ;
      RECT 68.755 -31.375 68.895 -31.205 ;
      RECT 68.755 -30.478 68.845 -29.471 ;
      RECT 68.755 -30.165 68.895 -29.995 ;
      RECT 68.755 -28.669 68.845 -27.662 ;
      RECT 68.755 -28.145 68.895 -27.975 ;
      RECT 68.755 -27.248 68.845 -26.241 ;
      RECT 68.755 -26.935 68.895 -26.765 ;
      RECT 68.755 -25.439 68.845 -24.432 ;
      RECT 68.755 -24.915 68.895 -24.745 ;
      RECT 68.755 -24.018 68.845 -23.011 ;
      RECT 68.755 -23.705 68.895 -23.535 ;
      RECT 68.755 -22.209 68.845 -21.202 ;
      RECT 68.755 -21.685 68.895 -21.515 ;
      RECT 68.755 -20.788 68.845 -19.781 ;
      RECT 68.755 -20.475 68.895 -20.305 ;
      RECT 68.755 -18.979 68.845 -17.972 ;
      RECT 68.755 -18.455 68.895 -18.285 ;
      RECT 68.755 -17.558 68.845 -16.551 ;
      RECT 68.755 -17.245 68.895 -17.075 ;
      RECT 68.755 -15.749 68.845 -14.742 ;
      RECT 68.755 -15.225 68.895 -15.055 ;
      RECT 68.755 -14.328 68.845 -13.321 ;
      RECT 68.755 -14.015 68.895 -13.845 ;
      RECT 68.755 -12.519 68.845 -11.512 ;
      RECT 68.755 -11.995 68.895 -11.825 ;
      RECT 68.755 -11.098 68.845 -10.091 ;
      RECT 68.755 -10.785 68.895 -10.615 ;
      RECT 68.755 -9.289 68.845 -8.282 ;
      RECT 68.755 -8.765 68.895 -8.595 ;
      RECT 68.755 -7.868 68.845 -6.861 ;
      RECT 68.755 -7.555 68.895 -7.385 ;
      RECT 68.755 -6.059 68.845 -5.052 ;
      RECT 68.755 -5.535 68.895 -5.365 ;
      RECT 68.755 -4.638 68.845 -3.631 ;
      RECT 68.755 -4.325 68.895 -4.155 ;
      RECT 68.755 -2.829 68.845 -1.822 ;
      RECT 68.755 -2.305 68.895 -2.135 ;
      RECT 68.755 -1.408 68.845 -0.401 ;
      RECT 68.755 -1.095 68.895 -0.925 ;
      RECT 68.755 0.401 68.845 1.408 ;
      RECT 68.755 0.925 68.895 1.095 ;
      RECT 68.44 -114.685 68.61 -114.515 ;
      RECT 68.51 -114.895 68.61 -114.515 ;
      RECT 67.955 -101.538 68.045 -100.53 ;
      RECT 67.905 -100.935 68.045 -100.765 ;
      RECT 67.955 -99.73 68.045 -98.722 ;
      RECT 67.905 -99.495 68.045 -99.325 ;
      RECT 67.955 -98.308 68.045 -97.3 ;
      RECT 67.905 -97.705 68.045 -97.535 ;
      RECT 67.955 -96.5 68.045 -95.492 ;
      RECT 67.905 -96.265 68.045 -96.095 ;
      RECT 67.955 -95.078 68.045 -94.07 ;
      RECT 67.905 -94.475 68.045 -94.305 ;
      RECT 67.955 -93.27 68.045 -92.262 ;
      RECT 67.905 -93.035 68.045 -92.865 ;
      RECT 67.955 -91.848 68.045 -90.84 ;
      RECT 67.905 -91.245 68.045 -91.075 ;
      RECT 67.955 -90.04 68.045 -89.032 ;
      RECT 67.905 -89.805 68.045 -89.635 ;
      RECT 67.955 -88.618 68.045 -87.61 ;
      RECT 67.905 -88.015 68.045 -87.845 ;
      RECT 67.955 -86.81 68.045 -85.802 ;
      RECT 67.905 -86.575 68.045 -86.405 ;
      RECT 67.955 -85.388 68.045 -84.38 ;
      RECT 67.905 -84.785 68.045 -84.615 ;
      RECT 67.955 -83.58 68.045 -82.572 ;
      RECT 67.905 -83.345 68.045 -83.175 ;
      RECT 67.955 -82.158 68.045 -81.15 ;
      RECT 67.905 -81.555 68.045 -81.385 ;
      RECT 67.955 -80.35 68.045 -79.342 ;
      RECT 67.905 -80.115 68.045 -79.945 ;
      RECT 67.955 -78.928 68.045 -77.92 ;
      RECT 67.905 -78.325 68.045 -78.155 ;
      RECT 67.955 -77.12 68.045 -76.112 ;
      RECT 67.905 -76.885 68.045 -76.715 ;
      RECT 67.955 -75.698 68.045 -74.69 ;
      RECT 67.905 -75.095 68.045 -74.925 ;
      RECT 67.955 -73.89 68.045 -72.882 ;
      RECT 67.905 -73.655 68.045 -73.485 ;
      RECT 67.955 -72.468 68.045 -71.46 ;
      RECT 67.905 -71.865 68.045 -71.695 ;
      RECT 67.955 -70.66 68.045 -69.652 ;
      RECT 67.905 -70.425 68.045 -70.255 ;
      RECT 67.955 -69.238 68.045 -68.23 ;
      RECT 67.905 -68.635 68.045 -68.465 ;
      RECT 67.955 -67.43 68.045 -66.422 ;
      RECT 67.905 -67.195 68.045 -67.025 ;
      RECT 67.955 -66.008 68.045 -65 ;
      RECT 67.905 -65.405 68.045 -65.235 ;
      RECT 67.955 -64.2 68.045 -63.192 ;
      RECT 67.905 -63.965 68.045 -63.795 ;
      RECT 67.955 -62.778 68.045 -61.77 ;
      RECT 67.905 -62.175 68.045 -62.005 ;
      RECT 67.955 -60.97 68.045 -59.962 ;
      RECT 67.905 -60.735 68.045 -60.565 ;
      RECT 67.955 -59.548 68.045 -58.54 ;
      RECT 67.905 -58.945 68.045 -58.775 ;
      RECT 67.955 -57.74 68.045 -56.732 ;
      RECT 67.905 -57.505 68.045 -57.335 ;
      RECT 67.955 -56.318 68.045 -55.31 ;
      RECT 67.905 -55.715 68.045 -55.545 ;
      RECT 67.955 -54.51 68.045 -53.502 ;
      RECT 67.905 -54.275 68.045 -54.105 ;
      RECT 67.955 -53.088 68.045 -52.08 ;
      RECT 67.905 -52.485 68.045 -52.315 ;
      RECT 67.955 -51.28 68.045 -50.272 ;
      RECT 67.905 -51.045 68.045 -50.875 ;
      RECT 67.955 -49.858 68.045 -48.85 ;
      RECT 67.905 -49.255 68.045 -49.085 ;
      RECT 67.955 -48.05 68.045 -47.042 ;
      RECT 67.905 -47.815 68.045 -47.645 ;
      RECT 67.955 -46.628 68.045 -45.62 ;
      RECT 67.905 -46.025 68.045 -45.855 ;
      RECT 67.955 -44.82 68.045 -43.812 ;
      RECT 67.905 -44.585 68.045 -44.415 ;
      RECT 67.955 -43.398 68.045 -42.39 ;
      RECT 67.905 -42.795 68.045 -42.625 ;
      RECT 67.955 -41.59 68.045 -40.582 ;
      RECT 67.905 -41.355 68.045 -41.185 ;
      RECT 67.955 -40.168 68.045 -39.16 ;
      RECT 67.905 -39.565 68.045 -39.395 ;
      RECT 67.955 -38.36 68.045 -37.352 ;
      RECT 67.905 -38.125 68.045 -37.955 ;
      RECT 67.955 -36.938 68.045 -35.93 ;
      RECT 67.905 -36.335 68.045 -36.165 ;
      RECT 67.955 -35.13 68.045 -34.122 ;
      RECT 67.905 -34.895 68.045 -34.725 ;
      RECT 67.955 -33.708 68.045 -32.7 ;
      RECT 67.905 -33.105 68.045 -32.935 ;
      RECT 67.955 -31.9 68.045 -30.892 ;
      RECT 67.905 -31.665 68.045 -31.495 ;
      RECT 67.955 -30.478 68.045 -29.47 ;
      RECT 67.905 -29.875 68.045 -29.705 ;
      RECT 67.955 -28.67 68.045 -27.662 ;
      RECT 67.905 -28.435 68.045 -28.265 ;
      RECT 67.955 -27.248 68.045 -26.24 ;
      RECT 67.905 -26.645 68.045 -26.475 ;
      RECT 67.955 -25.44 68.045 -24.432 ;
      RECT 67.905 -25.205 68.045 -25.035 ;
      RECT 67.955 -24.018 68.045 -23.01 ;
      RECT 67.905 -23.415 68.045 -23.245 ;
      RECT 67.955 -22.21 68.045 -21.202 ;
      RECT 67.905 -21.975 68.045 -21.805 ;
      RECT 67.955 -20.788 68.045 -19.78 ;
      RECT 67.905 -20.185 68.045 -20.015 ;
      RECT 67.955 -18.98 68.045 -17.972 ;
      RECT 67.905 -18.745 68.045 -18.575 ;
      RECT 67.955 -17.558 68.045 -16.55 ;
      RECT 67.905 -16.955 68.045 -16.785 ;
      RECT 67.955 -15.75 68.045 -14.742 ;
      RECT 67.905 -15.515 68.045 -15.345 ;
      RECT 67.955 -14.328 68.045 -13.32 ;
      RECT 67.905 -13.725 68.045 -13.555 ;
      RECT 67.955 -12.52 68.045 -11.512 ;
      RECT 67.905 -12.285 68.045 -12.115 ;
      RECT 67.955 -11.098 68.045 -10.09 ;
      RECT 67.905 -10.495 68.045 -10.325 ;
      RECT 67.955 -9.29 68.045 -8.282 ;
      RECT 67.905 -9.055 68.045 -8.885 ;
      RECT 67.955 -7.868 68.045 -6.86 ;
      RECT 67.905 -7.265 68.045 -7.095 ;
      RECT 67.955 -6.06 68.045 -5.052 ;
      RECT 67.905 -5.825 68.045 -5.655 ;
      RECT 67.955 -4.638 68.045 -3.63 ;
      RECT 67.905 -4.035 68.045 -3.865 ;
      RECT 67.955 -2.83 68.045 -1.822 ;
      RECT 67.905 -2.595 68.045 -2.425 ;
      RECT 67.955 -1.408 68.045 -0.4 ;
      RECT 67.905 -0.805 68.045 -0.635 ;
      RECT 67.955 0.4 68.045 1.408 ;
      RECT 67.905 0.635 68.045 0.805 ;
      RECT 67.555 -101.538 67.645 -100.531 ;
      RECT 67.555 -101.225 67.695 -101.055 ;
      RECT 67.555 -99.729 67.645 -98.722 ;
      RECT 67.555 -99.205 67.695 -99.035 ;
      RECT 67.555 -98.308 67.645 -97.301 ;
      RECT 67.555 -97.995 67.695 -97.825 ;
      RECT 67.555 -96.499 67.645 -95.492 ;
      RECT 67.555 -95.975 67.695 -95.805 ;
      RECT 67.555 -95.078 67.645 -94.071 ;
      RECT 67.555 -94.765 67.695 -94.595 ;
      RECT 67.555 -93.269 67.645 -92.262 ;
      RECT 67.555 -92.745 67.695 -92.575 ;
      RECT 67.555 -91.848 67.645 -90.841 ;
      RECT 67.555 -91.535 67.695 -91.365 ;
      RECT 67.555 -90.039 67.645 -89.032 ;
      RECT 67.555 -89.515 67.695 -89.345 ;
      RECT 67.555 -88.618 67.645 -87.611 ;
      RECT 67.555 -88.305 67.695 -88.135 ;
      RECT 67.555 -86.809 67.645 -85.802 ;
      RECT 67.555 -86.285 67.695 -86.115 ;
      RECT 67.555 -85.388 67.645 -84.381 ;
      RECT 67.555 -85.075 67.695 -84.905 ;
      RECT 67.555 -83.579 67.645 -82.572 ;
      RECT 67.555 -83.055 67.695 -82.885 ;
      RECT 67.555 -82.158 67.645 -81.151 ;
      RECT 67.555 -81.845 67.695 -81.675 ;
      RECT 67.555 -80.349 67.645 -79.342 ;
      RECT 67.555 -79.825 67.695 -79.655 ;
      RECT 67.555 -78.928 67.645 -77.921 ;
      RECT 67.555 -78.615 67.695 -78.445 ;
      RECT 67.555 -77.119 67.645 -76.112 ;
      RECT 67.555 -76.595 67.695 -76.425 ;
      RECT 67.555 -75.698 67.645 -74.691 ;
      RECT 67.555 -75.385 67.695 -75.215 ;
      RECT 67.555 -73.889 67.645 -72.882 ;
      RECT 67.555 -73.365 67.695 -73.195 ;
      RECT 67.555 -72.468 67.645 -71.461 ;
      RECT 67.555 -72.155 67.695 -71.985 ;
      RECT 67.555 -70.659 67.645 -69.652 ;
      RECT 67.555 -70.135 67.695 -69.965 ;
      RECT 67.555 -69.238 67.645 -68.231 ;
      RECT 67.555 -68.925 67.695 -68.755 ;
      RECT 67.555 -67.429 67.645 -66.422 ;
      RECT 67.555 -66.905 67.695 -66.735 ;
      RECT 67.555 -66.008 67.645 -65.001 ;
      RECT 67.555 -65.695 67.695 -65.525 ;
      RECT 67.555 -64.199 67.645 -63.192 ;
      RECT 67.555 -63.675 67.695 -63.505 ;
      RECT 67.555 -62.778 67.645 -61.771 ;
      RECT 67.555 -62.465 67.695 -62.295 ;
      RECT 67.555 -60.969 67.645 -59.962 ;
      RECT 67.555 -60.445 67.695 -60.275 ;
      RECT 67.555 -59.548 67.645 -58.541 ;
      RECT 67.555 -59.235 67.695 -59.065 ;
      RECT 67.555 -57.739 67.645 -56.732 ;
      RECT 67.555 -57.215 67.695 -57.045 ;
      RECT 67.555 -56.318 67.645 -55.311 ;
      RECT 67.555 -56.005 67.695 -55.835 ;
      RECT 67.555 -54.509 67.645 -53.502 ;
      RECT 67.555 -53.985 67.695 -53.815 ;
      RECT 67.555 -53.088 67.645 -52.081 ;
      RECT 67.555 -52.775 67.695 -52.605 ;
      RECT 67.555 -51.279 67.645 -50.272 ;
      RECT 67.555 -50.755 67.695 -50.585 ;
      RECT 67.555 -49.858 67.645 -48.851 ;
      RECT 67.555 -49.545 67.695 -49.375 ;
      RECT 67.555 -48.049 67.645 -47.042 ;
      RECT 67.555 -47.525 67.695 -47.355 ;
      RECT 67.555 -46.628 67.645 -45.621 ;
      RECT 67.555 -46.315 67.695 -46.145 ;
      RECT 67.555 -44.819 67.645 -43.812 ;
      RECT 67.555 -44.295 67.695 -44.125 ;
      RECT 67.555 -43.398 67.645 -42.391 ;
      RECT 67.555 -43.085 67.695 -42.915 ;
      RECT 67.555 -41.589 67.645 -40.582 ;
      RECT 67.555 -41.065 67.695 -40.895 ;
      RECT 67.555 -40.168 67.645 -39.161 ;
      RECT 67.555 -39.855 67.695 -39.685 ;
      RECT 67.555 -38.359 67.645 -37.352 ;
      RECT 67.555 -37.835 67.695 -37.665 ;
      RECT 67.555 -36.938 67.645 -35.931 ;
      RECT 67.555 -36.625 67.695 -36.455 ;
      RECT 67.555 -35.129 67.645 -34.122 ;
      RECT 67.555 -34.605 67.695 -34.435 ;
      RECT 67.555 -33.708 67.645 -32.701 ;
      RECT 67.555 -33.395 67.695 -33.225 ;
      RECT 67.555 -31.899 67.645 -30.892 ;
      RECT 67.555 -31.375 67.695 -31.205 ;
      RECT 67.555 -30.478 67.645 -29.471 ;
      RECT 67.555 -30.165 67.695 -29.995 ;
      RECT 67.555 -28.669 67.645 -27.662 ;
      RECT 67.555 -28.145 67.695 -27.975 ;
      RECT 67.555 -27.248 67.645 -26.241 ;
      RECT 67.555 -26.935 67.695 -26.765 ;
      RECT 67.555 -25.439 67.645 -24.432 ;
      RECT 67.555 -24.915 67.695 -24.745 ;
      RECT 67.555 -24.018 67.645 -23.011 ;
      RECT 67.555 -23.705 67.695 -23.535 ;
      RECT 67.555 -22.209 67.645 -21.202 ;
      RECT 67.555 -21.685 67.695 -21.515 ;
      RECT 67.555 -20.788 67.645 -19.781 ;
      RECT 67.555 -20.475 67.695 -20.305 ;
      RECT 67.555 -18.979 67.645 -17.972 ;
      RECT 67.555 -18.455 67.695 -18.285 ;
      RECT 67.555 -17.558 67.645 -16.551 ;
      RECT 67.555 -17.245 67.695 -17.075 ;
      RECT 67.555 -15.749 67.645 -14.742 ;
      RECT 67.555 -15.225 67.695 -15.055 ;
      RECT 67.555 -14.328 67.645 -13.321 ;
      RECT 67.555 -14.015 67.695 -13.845 ;
      RECT 67.555 -12.519 67.645 -11.512 ;
      RECT 67.555 -11.995 67.695 -11.825 ;
      RECT 67.555 -11.098 67.645 -10.091 ;
      RECT 67.555 -10.785 67.695 -10.615 ;
      RECT 67.555 -9.289 67.645 -8.282 ;
      RECT 67.555 -8.765 67.695 -8.595 ;
      RECT 67.555 -7.868 67.645 -6.861 ;
      RECT 67.555 -7.555 67.695 -7.385 ;
      RECT 67.555 -6.059 67.645 -5.052 ;
      RECT 67.555 -5.535 67.695 -5.365 ;
      RECT 67.555 -4.638 67.645 -3.631 ;
      RECT 67.555 -4.325 67.695 -4.155 ;
      RECT 67.555 -2.829 67.645 -1.822 ;
      RECT 67.555 -2.305 67.695 -2.135 ;
      RECT 67.555 -1.408 67.645 -0.401 ;
      RECT 67.555 -1.095 67.695 -0.925 ;
      RECT 67.555 0.401 67.645 1.408 ;
      RECT 67.555 0.925 67.695 1.095 ;
      RECT 63.385 -108.935 67.165 -108.815 ;
      RECT 64.705 -109.475 64.805 -108.815 ;
      RECT 64.145 -109.475 64.245 -108.815 ;
      RECT 63.585 -109.475 63.685 -108.815 ;
      RECT 66.755 -101.538 66.845 -100.53 ;
      RECT 66.705 -100.935 66.845 -100.765 ;
      RECT 66.755 -99.73 66.845 -98.722 ;
      RECT 66.705 -99.495 66.845 -99.325 ;
      RECT 66.755 -98.308 66.845 -97.3 ;
      RECT 66.705 -97.705 66.845 -97.535 ;
      RECT 66.755 -96.5 66.845 -95.492 ;
      RECT 66.705 -96.265 66.845 -96.095 ;
      RECT 66.755 -95.078 66.845 -94.07 ;
      RECT 66.705 -94.475 66.845 -94.305 ;
      RECT 66.755 -93.27 66.845 -92.262 ;
      RECT 66.705 -93.035 66.845 -92.865 ;
      RECT 66.755 -91.848 66.845 -90.84 ;
      RECT 66.705 -91.245 66.845 -91.075 ;
      RECT 66.755 -90.04 66.845 -89.032 ;
      RECT 66.705 -89.805 66.845 -89.635 ;
      RECT 66.755 -88.618 66.845 -87.61 ;
      RECT 66.705 -88.015 66.845 -87.845 ;
      RECT 66.755 -86.81 66.845 -85.802 ;
      RECT 66.705 -86.575 66.845 -86.405 ;
      RECT 66.755 -85.388 66.845 -84.38 ;
      RECT 66.705 -84.785 66.845 -84.615 ;
      RECT 66.755 -83.58 66.845 -82.572 ;
      RECT 66.705 -83.345 66.845 -83.175 ;
      RECT 66.755 -82.158 66.845 -81.15 ;
      RECT 66.705 -81.555 66.845 -81.385 ;
      RECT 66.755 -80.35 66.845 -79.342 ;
      RECT 66.705 -80.115 66.845 -79.945 ;
      RECT 66.755 -78.928 66.845 -77.92 ;
      RECT 66.705 -78.325 66.845 -78.155 ;
      RECT 66.755 -77.12 66.845 -76.112 ;
      RECT 66.705 -76.885 66.845 -76.715 ;
      RECT 66.755 -75.698 66.845 -74.69 ;
      RECT 66.705 -75.095 66.845 -74.925 ;
      RECT 66.755 -73.89 66.845 -72.882 ;
      RECT 66.705 -73.655 66.845 -73.485 ;
      RECT 66.755 -72.468 66.845 -71.46 ;
      RECT 66.705 -71.865 66.845 -71.695 ;
      RECT 66.755 -70.66 66.845 -69.652 ;
      RECT 66.705 -70.425 66.845 -70.255 ;
      RECT 66.755 -69.238 66.845 -68.23 ;
      RECT 66.705 -68.635 66.845 -68.465 ;
      RECT 66.755 -67.43 66.845 -66.422 ;
      RECT 66.705 -67.195 66.845 -67.025 ;
      RECT 66.755 -66.008 66.845 -65 ;
      RECT 66.705 -65.405 66.845 -65.235 ;
      RECT 66.755 -64.2 66.845 -63.192 ;
      RECT 66.705 -63.965 66.845 -63.795 ;
      RECT 66.755 -62.778 66.845 -61.77 ;
      RECT 66.705 -62.175 66.845 -62.005 ;
      RECT 66.755 -60.97 66.845 -59.962 ;
      RECT 66.705 -60.735 66.845 -60.565 ;
      RECT 66.755 -59.548 66.845 -58.54 ;
      RECT 66.705 -58.945 66.845 -58.775 ;
      RECT 66.755 -57.74 66.845 -56.732 ;
      RECT 66.705 -57.505 66.845 -57.335 ;
      RECT 66.755 -56.318 66.845 -55.31 ;
      RECT 66.705 -55.715 66.845 -55.545 ;
      RECT 66.755 -54.51 66.845 -53.502 ;
      RECT 66.705 -54.275 66.845 -54.105 ;
      RECT 66.755 -53.088 66.845 -52.08 ;
      RECT 66.705 -52.485 66.845 -52.315 ;
      RECT 66.755 -51.28 66.845 -50.272 ;
      RECT 66.705 -51.045 66.845 -50.875 ;
      RECT 66.755 -49.858 66.845 -48.85 ;
      RECT 66.705 -49.255 66.845 -49.085 ;
      RECT 66.755 -48.05 66.845 -47.042 ;
      RECT 66.705 -47.815 66.845 -47.645 ;
      RECT 66.755 -46.628 66.845 -45.62 ;
      RECT 66.705 -46.025 66.845 -45.855 ;
      RECT 66.755 -44.82 66.845 -43.812 ;
      RECT 66.705 -44.585 66.845 -44.415 ;
      RECT 66.755 -43.398 66.845 -42.39 ;
      RECT 66.705 -42.795 66.845 -42.625 ;
      RECT 66.755 -41.59 66.845 -40.582 ;
      RECT 66.705 -41.355 66.845 -41.185 ;
      RECT 66.755 -40.168 66.845 -39.16 ;
      RECT 66.705 -39.565 66.845 -39.395 ;
      RECT 66.755 -38.36 66.845 -37.352 ;
      RECT 66.705 -38.125 66.845 -37.955 ;
      RECT 66.755 -36.938 66.845 -35.93 ;
      RECT 66.705 -36.335 66.845 -36.165 ;
      RECT 66.755 -35.13 66.845 -34.122 ;
      RECT 66.705 -34.895 66.845 -34.725 ;
      RECT 66.755 -33.708 66.845 -32.7 ;
      RECT 66.705 -33.105 66.845 -32.935 ;
      RECT 66.755 -31.9 66.845 -30.892 ;
      RECT 66.705 -31.665 66.845 -31.495 ;
      RECT 66.755 -30.478 66.845 -29.47 ;
      RECT 66.705 -29.875 66.845 -29.705 ;
      RECT 66.755 -28.67 66.845 -27.662 ;
      RECT 66.705 -28.435 66.845 -28.265 ;
      RECT 66.755 -27.248 66.845 -26.24 ;
      RECT 66.705 -26.645 66.845 -26.475 ;
      RECT 66.755 -25.44 66.845 -24.432 ;
      RECT 66.705 -25.205 66.845 -25.035 ;
      RECT 66.755 -24.018 66.845 -23.01 ;
      RECT 66.705 -23.415 66.845 -23.245 ;
      RECT 66.755 -22.21 66.845 -21.202 ;
      RECT 66.705 -21.975 66.845 -21.805 ;
      RECT 66.755 -20.788 66.845 -19.78 ;
      RECT 66.705 -20.185 66.845 -20.015 ;
      RECT 66.755 -18.98 66.845 -17.972 ;
      RECT 66.705 -18.745 66.845 -18.575 ;
      RECT 66.755 -17.558 66.845 -16.55 ;
      RECT 66.705 -16.955 66.845 -16.785 ;
      RECT 66.755 -15.75 66.845 -14.742 ;
      RECT 66.705 -15.515 66.845 -15.345 ;
      RECT 66.755 -14.328 66.845 -13.32 ;
      RECT 66.705 -13.725 66.845 -13.555 ;
      RECT 66.755 -12.52 66.845 -11.512 ;
      RECT 66.705 -12.285 66.845 -12.115 ;
      RECT 66.755 -11.098 66.845 -10.09 ;
      RECT 66.705 -10.495 66.845 -10.325 ;
      RECT 66.755 -9.29 66.845 -8.282 ;
      RECT 66.705 -9.055 66.845 -8.885 ;
      RECT 66.755 -7.868 66.845 -6.86 ;
      RECT 66.705 -7.265 66.845 -7.095 ;
      RECT 66.755 -6.06 66.845 -5.052 ;
      RECT 66.705 -5.825 66.845 -5.655 ;
      RECT 66.755 -4.638 66.845 -3.63 ;
      RECT 66.705 -4.035 66.845 -3.865 ;
      RECT 66.755 -2.83 66.845 -1.822 ;
      RECT 66.705 -2.595 66.845 -2.425 ;
      RECT 66.755 -1.408 66.845 -0.4 ;
      RECT 66.705 -0.805 66.845 -0.635 ;
      RECT 66.755 0.4 66.845 1.408 ;
      RECT 66.705 0.635 66.845 0.805 ;
      RECT 65.325 -111.685 66.805 -111.585 ;
      RECT 65.325 -112.195 65.425 -111.585 ;
      RECT 65.545 -109.15 66.805 -109.05 ;
      RECT 66.705 -109.475 66.805 -109.05 ;
      RECT 66.145 -109.475 66.245 -109.05 ;
      RECT 65.585 -109.475 65.685 -109.05 ;
      RECT 66.355 -101.538 66.445 -100.531 ;
      RECT 66.355 -101.225 66.495 -101.055 ;
      RECT 66.355 -99.729 66.445 -98.722 ;
      RECT 66.355 -99.205 66.495 -99.035 ;
      RECT 66.355 -98.308 66.445 -97.301 ;
      RECT 66.355 -97.995 66.495 -97.825 ;
      RECT 66.355 -96.499 66.445 -95.492 ;
      RECT 66.355 -95.975 66.495 -95.805 ;
      RECT 66.355 -95.078 66.445 -94.071 ;
      RECT 66.355 -94.765 66.495 -94.595 ;
      RECT 66.355 -93.269 66.445 -92.262 ;
      RECT 66.355 -92.745 66.495 -92.575 ;
      RECT 66.355 -91.848 66.445 -90.841 ;
      RECT 66.355 -91.535 66.495 -91.365 ;
      RECT 66.355 -90.039 66.445 -89.032 ;
      RECT 66.355 -89.515 66.495 -89.345 ;
      RECT 66.355 -88.618 66.445 -87.611 ;
      RECT 66.355 -88.305 66.495 -88.135 ;
      RECT 66.355 -86.809 66.445 -85.802 ;
      RECT 66.355 -86.285 66.495 -86.115 ;
      RECT 66.355 -85.388 66.445 -84.381 ;
      RECT 66.355 -85.075 66.495 -84.905 ;
      RECT 66.355 -83.579 66.445 -82.572 ;
      RECT 66.355 -83.055 66.495 -82.885 ;
      RECT 66.355 -82.158 66.445 -81.151 ;
      RECT 66.355 -81.845 66.495 -81.675 ;
      RECT 66.355 -80.349 66.445 -79.342 ;
      RECT 66.355 -79.825 66.495 -79.655 ;
      RECT 66.355 -78.928 66.445 -77.921 ;
      RECT 66.355 -78.615 66.495 -78.445 ;
      RECT 66.355 -77.119 66.445 -76.112 ;
      RECT 66.355 -76.595 66.495 -76.425 ;
      RECT 66.355 -75.698 66.445 -74.691 ;
      RECT 66.355 -75.385 66.495 -75.215 ;
      RECT 66.355 -73.889 66.445 -72.882 ;
      RECT 66.355 -73.365 66.495 -73.195 ;
      RECT 66.355 -72.468 66.445 -71.461 ;
      RECT 66.355 -72.155 66.495 -71.985 ;
      RECT 66.355 -70.659 66.445 -69.652 ;
      RECT 66.355 -70.135 66.495 -69.965 ;
      RECT 66.355 -69.238 66.445 -68.231 ;
      RECT 66.355 -68.925 66.495 -68.755 ;
      RECT 66.355 -67.429 66.445 -66.422 ;
      RECT 66.355 -66.905 66.495 -66.735 ;
      RECT 66.355 -66.008 66.445 -65.001 ;
      RECT 66.355 -65.695 66.495 -65.525 ;
      RECT 66.355 -64.199 66.445 -63.192 ;
      RECT 66.355 -63.675 66.495 -63.505 ;
      RECT 66.355 -62.778 66.445 -61.771 ;
      RECT 66.355 -62.465 66.495 -62.295 ;
      RECT 66.355 -60.969 66.445 -59.962 ;
      RECT 66.355 -60.445 66.495 -60.275 ;
      RECT 66.355 -59.548 66.445 -58.541 ;
      RECT 66.355 -59.235 66.495 -59.065 ;
      RECT 66.355 -57.739 66.445 -56.732 ;
      RECT 66.355 -57.215 66.495 -57.045 ;
      RECT 66.355 -56.318 66.445 -55.311 ;
      RECT 66.355 -56.005 66.495 -55.835 ;
      RECT 66.355 -54.509 66.445 -53.502 ;
      RECT 66.355 -53.985 66.495 -53.815 ;
      RECT 66.355 -53.088 66.445 -52.081 ;
      RECT 66.355 -52.775 66.495 -52.605 ;
      RECT 66.355 -51.279 66.445 -50.272 ;
      RECT 66.355 -50.755 66.495 -50.585 ;
      RECT 66.355 -49.858 66.445 -48.851 ;
      RECT 66.355 -49.545 66.495 -49.375 ;
      RECT 66.355 -48.049 66.445 -47.042 ;
      RECT 66.355 -47.525 66.495 -47.355 ;
      RECT 66.355 -46.628 66.445 -45.621 ;
      RECT 66.355 -46.315 66.495 -46.145 ;
      RECT 66.355 -44.819 66.445 -43.812 ;
      RECT 66.355 -44.295 66.495 -44.125 ;
      RECT 66.355 -43.398 66.445 -42.391 ;
      RECT 66.355 -43.085 66.495 -42.915 ;
      RECT 66.355 -41.589 66.445 -40.582 ;
      RECT 66.355 -41.065 66.495 -40.895 ;
      RECT 66.355 -40.168 66.445 -39.161 ;
      RECT 66.355 -39.855 66.495 -39.685 ;
      RECT 66.355 -38.359 66.445 -37.352 ;
      RECT 66.355 -37.835 66.495 -37.665 ;
      RECT 66.355 -36.938 66.445 -35.931 ;
      RECT 66.355 -36.625 66.495 -36.455 ;
      RECT 66.355 -35.129 66.445 -34.122 ;
      RECT 66.355 -34.605 66.495 -34.435 ;
      RECT 66.355 -33.708 66.445 -32.701 ;
      RECT 66.355 -33.395 66.495 -33.225 ;
      RECT 66.355 -31.899 66.445 -30.892 ;
      RECT 66.355 -31.375 66.495 -31.205 ;
      RECT 66.355 -30.478 66.445 -29.471 ;
      RECT 66.355 -30.165 66.495 -29.995 ;
      RECT 66.355 -28.669 66.445 -27.662 ;
      RECT 66.355 -28.145 66.495 -27.975 ;
      RECT 66.355 -27.248 66.445 -26.241 ;
      RECT 66.355 -26.935 66.495 -26.765 ;
      RECT 66.355 -25.439 66.445 -24.432 ;
      RECT 66.355 -24.915 66.495 -24.745 ;
      RECT 66.355 -24.018 66.445 -23.011 ;
      RECT 66.355 -23.705 66.495 -23.535 ;
      RECT 66.355 -22.209 66.445 -21.202 ;
      RECT 66.355 -21.685 66.495 -21.515 ;
      RECT 66.355 -20.788 66.445 -19.781 ;
      RECT 66.355 -20.475 66.495 -20.305 ;
      RECT 66.355 -18.979 66.445 -17.972 ;
      RECT 66.355 -18.455 66.495 -18.285 ;
      RECT 66.355 -17.558 66.445 -16.551 ;
      RECT 66.355 -17.245 66.495 -17.075 ;
      RECT 66.355 -15.749 66.445 -14.742 ;
      RECT 66.355 -15.225 66.495 -15.055 ;
      RECT 66.355 -14.328 66.445 -13.321 ;
      RECT 66.355 -14.015 66.495 -13.845 ;
      RECT 66.355 -12.519 66.445 -11.512 ;
      RECT 66.355 -11.995 66.495 -11.825 ;
      RECT 66.355 -11.098 66.445 -10.091 ;
      RECT 66.355 -10.785 66.495 -10.615 ;
      RECT 66.355 -9.289 66.445 -8.282 ;
      RECT 66.355 -8.765 66.495 -8.595 ;
      RECT 66.355 -7.868 66.445 -6.861 ;
      RECT 66.355 -7.555 66.495 -7.385 ;
      RECT 66.355 -6.059 66.445 -5.052 ;
      RECT 66.355 -5.535 66.495 -5.365 ;
      RECT 66.355 -4.638 66.445 -3.631 ;
      RECT 66.355 -4.325 66.495 -4.155 ;
      RECT 66.355 -2.829 66.445 -1.822 ;
      RECT 66.355 -2.305 66.495 -2.135 ;
      RECT 66.355 -1.408 66.445 -0.401 ;
      RECT 66.355 -1.095 66.495 -0.925 ;
      RECT 66.355 0.401 66.445 1.408 ;
      RECT 66.355 0.925 66.495 1.095 ;
      RECT 65.685 -111.495 65.855 -111.385 ;
      RECT 62.535 -111.495 65.855 -111.395 ;
      RECT 65.555 -101.538 65.645 -100.53 ;
      RECT 65.505 -100.935 65.645 -100.765 ;
      RECT 65.555 -99.73 65.645 -98.722 ;
      RECT 65.505 -99.495 65.645 -99.325 ;
      RECT 65.555 -98.308 65.645 -97.3 ;
      RECT 65.505 -97.705 65.645 -97.535 ;
      RECT 65.555 -96.5 65.645 -95.492 ;
      RECT 65.505 -96.265 65.645 -96.095 ;
      RECT 65.555 -95.078 65.645 -94.07 ;
      RECT 65.505 -94.475 65.645 -94.305 ;
      RECT 65.555 -93.27 65.645 -92.262 ;
      RECT 65.505 -93.035 65.645 -92.865 ;
      RECT 65.555 -91.848 65.645 -90.84 ;
      RECT 65.505 -91.245 65.645 -91.075 ;
      RECT 65.555 -90.04 65.645 -89.032 ;
      RECT 65.505 -89.805 65.645 -89.635 ;
      RECT 65.555 -88.618 65.645 -87.61 ;
      RECT 65.505 -88.015 65.645 -87.845 ;
      RECT 65.555 -86.81 65.645 -85.802 ;
      RECT 65.505 -86.575 65.645 -86.405 ;
      RECT 65.555 -85.388 65.645 -84.38 ;
      RECT 65.505 -84.785 65.645 -84.615 ;
      RECT 65.555 -83.58 65.645 -82.572 ;
      RECT 65.505 -83.345 65.645 -83.175 ;
      RECT 65.555 -82.158 65.645 -81.15 ;
      RECT 65.505 -81.555 65.645 -81.385 ;
      RECT 65.555 -80.35 65.645 -79.342 ;
      RECT 65.505 -80.115 65.645 -79.945 ;
      RECT 65.555 -78.928 65.645 -77.92 ;
      RECT 65.505 -78.325 65.645 -78.155 ;
      RECT 65.555 -77.12 65.645 -76.112 ;
      RECT 65.505 -76.885 65.645 -76.715 ;
      RECT 65.555 -75.698 65.645 -74.69 ;
      RECT 65.505 -75.095 65.645 -74.925 ;
      RECT 65.555 -73.89 65.645 -72.882 ;
      RECT 65.505 -73.655 65.645 -73.485 ;
      RECT 65.555 -72.468 65.645 -71.46 ;
      RECT 65.505 -71.865 65.645 -71.695 ;
      RECT 65.555 -70.66 65.645 -69.652 ;
      RECT 65.505 -70.425 65.645 -70.255 ;
      RECT 65.555 -69.238 65.645 -68.23 ;
      RECT 65.505 -68.635 65.645 -68.465 ;
      RECT 65.555 -67.43 65.645 -66.422 ;
      RECT 65.505 -67.195 65.645 -67.025 ;
      RECT 65.555 -66.008 65.645 -65 ;
      RECT 65.505 -65.405 65.645 -65.235 ;
      RECT 65.555 -64.2 65.645 -63.192 ;
      RECT 65.505 -63.965 65.645 -63.795 ;
      RECT 65.555 -62.778 65.645 -61.77 ;
      RECT 65.505 -62.175 65.645 -62.005 ;
      RECT 65.555 -60.97 65.645 -59.962 ;
      RECT 65.505 -60.735 65.645 -60.565 ;
      RECT 65.555 -59.548 65.645 -58.54 ;
      RECT 65.505 -58.945 65.645 -58.775 ;
      RECT 65.555 -57.74 65.645 -56.732 ;
      RECT 65.505 -57.505 65.645 -57.335 ;
      RECT 65.555 -56.318 65.645 -55.31 ;
      RECT 65.505 -55.715 65.645 -55.545 ;
      RECT 65.555 -54.51 65.645 -53.502 ;
      RECT 65.505 -54.275 65.645 -54.105 ;
      RECT 65.555 -53.088 65.645 -52.08 ;
      RECT 65.505 -52.485 65.645 -52.315 ;
      RECT 65.555 -51.28 65.645 -50.272 ;
      RECT 65.505 -51.045 65.645 -50.875 ;
      RECT 65.555 -49.858 65.645 -48.85 ;
      RECT 65.505 -49.255 65.645 -49.085 ;
      RECT 65.555 -48.05 65.645 -47.042 ;
      RECT 65.505 -47.815 65.645 -47.645 ;
      RECT 65.555 -46.628 65.645 -45.62 ;
      RECT 65.505 -46.025 65.645 -45.855 ;
      RECT 65.555 -44.82 65.645 -43.812 ;
      RECT 65.505 -44.585 65.645 -44.415 ;
      RECT 65.555 -43.398 65.645 -42.39 ;
      RECT 65.505 -42.795 65.645 -42.625 ;
      RECT 65.555 -41.59 65.645 -40.582 ;
      RECT 65.505 -41.355 65.645 -41.185 ;
      RECT 65.555 -40.168 65.645 -39.16 ;
      RECT 65.505 -39.565 65.645 -39.395 ;
      RECT 65.555 -38.36 65.645 -37.352 ;
      RECT 65.505 -38.125 65.645 -37.955 ;
      RECT 65.555 -36.938 65.645 -35.93 ;
      RECT 65.505 -36.335 65.645 -36.165 ;
      RECT 65.555 -35.13 65.645 -34.122 ;
      RECT 65.505 -34.895 65.645 -34.725 ;
      RECT 65.555 -33.708 65.645 -32.7 ;
      RECT 65.505 -33.105 65.645 -32.935 ;
      RECT 65.555 -31.9 65.645 -30.892 ;
      RECT 65.505 -31.665 65.645 -31.495 ;
      RECT 65.555 -30.478 65.645 -29.47 ;
      RECT 65.505 -29.875 65.645 -29.705 ;
      RECT 65.555 -28.67 65.645 -27.662 ;
      RECT 65.505 -28.435 65.645 -28.265 ;
      RECT 65.555 -27.248 65.645 -26.24 ;
      RECT 65.505 -26.645 65.645 -26.475 ;
      RECT 65.555 -25.44 65.645 -24.432 ;
      RECT 65.505 -25.205 65.645 -25.035 ;
      RECT 65.555 -24.018 65.645 -23.01 ;
      RECT 65.505 -23.415 65.645 -23.245 ;
      RECT 65.555 -22.21 65.645 -21.202 ;
      RECT 65.505 -21.975 65.645 -21.805 ;
      RECT 65.555 -20.788 65.645 -19.78 ;
      RECT 65.505 -20.185 65.645 -20.015 ;
      RECT 65.555 -18.98 65.645 -17.972 ;
      RECT 65.505 -18.745 65.645 -18.575 ;
      RECT 65.555 -17.558 65.645 -16.55 ;
      RECT 65.505 -16.955 65.645 -16.785 ;
      RECT 65.555 -15.75 65.645 -14.742 ;
      RECT 65.505 -15.515 65.645 -15.345 ;
      RECT 65.555 -14.328 65.645 -13.32 ;
      RECT 65.505 -13.725 65.645 -13.555 ;
      RECT 65.555 -12.52 65.645 -11.512 ;
      RECT 65.505 -12.285 65.645 -12.115 ;
      RECT 65.555 -11.098 65.645 -10.09 ;
      RECT 65.505 -10.495 65.645 -10.325 ;
      RECT 65.555 -9.29 65.645 -8.282 ;
      RECT 65.505 -9.055 65.645 -8.885 ;
      RECT 65.555 -7.868 65.645 -6.86 ;
      RECT 65.505 -7.265 65.645 -7.095 ;
      RECT 65.555 -6.06 65.645 -5.052 ;
      RECT 65.505 -5.825 65.645 -5.655 ;
      RECT 65.555 -4.638 65.645 -3.63 ;
      RECT 65.505 -4.035 65.645 -3.865 ;
      RECT 65.555 -2.83 65.645 -1.822 ;
      RECT 65.505 -2.595 65.645 -2.425 ;
      RECT 65.555 -1.408 65.645 -0.4 ;
      RECT 65.505 -0.805 65.645 -0.635 ;
      RECT 65.555 0.4 65.645 1.408 ;
      RECT 65.505 0.635 65.645 0.805 ;
      RECT 65.155 -101.538 65.245 -100.531 ;
      RECT 65.155 -101.225 65.295 -101.055 ;
      RECT 65.155 -99.729 65.245 -98.722 ;
      RECT 65.155 -99.205 65.295 -99.035 ;
      RECT 65.155 -98.308 65.245 -97.301 ;
      RECT 65.155 -97.995 65.295 -97.825 ;
      RECT 65.155 -96.499 65.245 -95.492 ;
      RECT 65.155 -95.975 65.295 -95.805 ;
      RECT 65.155 -95.078 65.245 -94.071 ;
      RECT 65.155 -94.765 65.295 -94.595 ;
      RECT 65.155 -93.269 65.245 -92.262 ;
      RECT 65.155 -92.745 65.295 -92.575 ;
      RECT 65.155 -91.848 65.245 -90.841 ;
      RECT 65.155 -91.535 65.295 -91.365 ;
      RECT 65.155 -90.039 65.245 -89.032 ;
      RECT 65.155 -89.515 65.295 -89.345 ;
      RECT 65.155 -88.618 65.245 -87.611 ;
      RECT 65.155 -88.305 65.295 -88.135 ;
      RECT 65.155 -86.809 65.245 -85.802 ;
      RECT 65.155 -86.285 65.295 -86.115 ;
      RECT 65.155 -85.388 65.245 -84.381 ;
      RECT 65.155 -85.075 65.295 -84.905 ;
      RECT 65.155 -83.579 65.245 -82.572 ;
      RECT 65.155 -83.055 65.295 -82.885 ;
      RECT 65.155 -82.158 65.245 -81.151 ;
      RECT 65.155 -81.845 65.295 -81.675 ;
      RECT 65.155 -80.349 65.245 -79.342 ;
      RECT 65.155 -79.825 65.295 -79.655 ;
      RECT 65.155 -78.928 65.245 -77.921 ;
      RECT 65.155 -78.615 65.295 -78.445 ;
      RECT 65.155 -77.119 65.245 -76.112 ;
      RECT 65.155 -76.595 65.295 -76.425 ;
      RECT 65.155 -75.698 65.245 -74.691 ;
      RECT 65.155 -75.385 65.295 -75.215 ;
      RECT 65.155 -73.889 65.245 -72.882 ;
      RECT 65.155 -73.365 65.295 -73.195 ;
      RECT 65.155 -72.468 65.245 -71.461 ;
      RECT 65.155 -72.155 65.295 -71.985 ;
      RECT 65.155 -70.659 65.245 -69.652 ;
      RECT 65.155 -70.135 65.295 -69.965 ;
      RECT 65.155 -69.238 65.245 -68.231 ;
      RECT 65.155 -68.925 65.295 -68.755 ;
      RECT 65.155 -67.429 65.245 -66.422 ;
      RECT 65.155 -66.905 65.295 -66.735 ;
      RECT 65.155 -66.008 65.245 -65.001 ;
      RECT 65.155 -65.695 65.295 -65.525 ;
      RECT 65.155 -64.199 65.245 -63.192 ;
      RECT 65.155 -63.675 65.295 -63.505 ;
      RECT 65.155 -62.778 65.245 -61.771 ;
      RECT 65.155 -62.465 65.295 -62.295 ;
      RECT 65.155 -60.969 65.245 -59.962 ;
      RECT 65.155 -60.445 65.295 -60.275 ;
      RECT 65.155 -59.548 65.245 -58.541 ;
      RECT 65.155 -59.235 65.295 -59.065 ;
      RECT 65.155 -57.739 65.245 -56.732 ;
      RECT 65.155 -57.215 65.295 -57.045 ;
      RECT 65.155 -56.318 65.245 -55.311 ;
      RECT 65.155 -56.005 65.295 -55.835 ;
      RECT 65.155 -54.509 65.245 -53.502 ;
      RECT 65.155 -53.985 65.295 -53.815 ;
      RECT 65.155 -53.088 65.245 -52.081 ;
      RECT 65.155 -52.775 65.295 -52.605 ;
      RECT 65.155 -51.279 65.245 -50.272 ;
      RECT 65.155 -50.755 65.295 -50.585 ;
      RECT 65.155 -49.858 65.245 -48.851 ;
      RECT 65.155 -49.545 65.295 -49.375 ;
      RECT 65.155 -48.049 65.245 -47.042 ;
      RECT 65.155 -47.525 65.295 -47.355 ;
      RECT 65.155 -46.628 65.245 -45.621 ;
      RECT 65.155 -46.315 65.295 -46.145 ;
      RECT 65.155 -44.819 65.245 -43.812 ;
      RECT 65.155 -44.295 65.295 -44.125 ;
      RECT 65.155 -43.398 65.245 -42.391 ;
      RECT 65.155 -43.085 65.295 -42.915 ;
      RECT 65.155 -41.589 65.245 -40.582 ;
      RECT 65.155 -41.065 65.295 -40.895 ;
      RECT 65.155 -40.168 65.245 -39.161 ;
      RECT 65.155 -39.855 65.295 -39.685 ;
      RECT 65.155 -38.359 65.245 -37.352 ;
      RECT 65.155 -37.835 65.295 -37.665 ;
      RECT 65.155 -36.938 65.245 -35.931 ;
      RECT 65.155 -36.625 65.295 -36.455 ;
      RECT 65.155 -35.129 65.245 -34.122 ;
      RECT 65.155 -34.605 65.295 -34.435 ;
      RECT 65.155 -33.708 65.245 -32.701 ;
      RECT 65.155 -33.395 65.295 -33.225 ;
      RECT 65.155 -31.899 65.245 -30.892 ;
      RECT 65.155 -31.375 65.295 -31.205 ;
      RECT 65.155 -30.478 65.245 -29.471 ;
      RECT 65.155 -30.165 65.295 -29.995 ;
      RECT 65.155 -28.669 65.245 -27.662 ;
      RECT 65.155 -28.145 65.295 -27.975 ;
      RECT 65.155 -27.248 65.245 -26.241 ;
      RECT 65.155 -26.935 65.295 -26.765 ;
      RECT 65.155 -25.439 65.245 -24.432 ;
      RECT 65.155 -24.915 65.295 -24.745 ;
      RECT 65.155 -24.018 65.245 -23.011 ;
      RECT 65.155 -23.705 65.295 -23.535 ;
      RECT 65.155 -22.209 65.245 -21.202 ;
      RECT 65.155 -21.685 65.295 -21.515 ;
      RECT 65.155 -20.788 65.245 -19.781 ;
      RECT 65.155 -20.475 65.295 -20.305 ;
      RECT 65.155 -18.979 65.245 -17.972 ;
      RECT 65.155 -18.455 65.295 -18.285 ;
      RECT 65.155 -17.558 65.245 -16.551 ;
      RECT 65.155 -17.245 65.295 -17.075 ;
      RECT 65.155 -15.749 65.245 -14.742 ;
      RECT 65.155 -15.225 65.295 -15.055 ;
      RECT 65.155 -14.328 65.245 -13.321 ;
      RECT 65.155 -14.015 65.295 -13.845 ;
      RECT 65.155 -12.519 65.245 -11.512 ;
      RECT 65.155 -11.995 65.295 -11.825 ;
      RECT 65.155 -11.098 65.245 -10.091 ;
      RECT 65.155 -10.785 65.295 -10.615 ;
      RECT 65.155 -9.289 65.245 -8.282 ;
      RECT 65.155 -8.765 65.295 -8.595 ;
      RECT 65.155 -7.868 65.245 -6.861 ;
      RECT 65.155 -7.555 65.295 -7.385 ;
      RECT 65.155 -6.059 65.245 -5.052 ;
      RECT 65.155 -5.535 65.295 -5.365 ;
      RECT 65.155 -4.638 65.245 -3.631 ;
      RECT 65.155 -4.325 65.295 -4.155 ;
      RECT 65.155 -2.829 65.245 -1.822 ;
      RECT 65.155 -2.305 65.295 -2.135 ;
      RECT 65.155 -1.408 65.245 -0.401 ;
      RECT 65.155 -1.095 65.295 -0.925 ;
      RECT 65.155 0.401 65.245 1.408 ;
      RECT 65.155 0.925 65.295 1.095 ;
      RECT 63.305 -111.685 64.785 -111.585 ;
      RECT 63.305 -112.055 63.405 -111.585 ;
      RECT 63.11 -114.395 64.685 -114.275 ;
      RECT 64.585 -114.895 64.685 -114.275 ;
      RECT 63.99 -114.895 64.09 -114.275 ;
      RECT 63.11 -114.85 63.21 -114.275 ;
      RECT 64.355 -101.538 64.445 -100.53 ;
      RECT 64.305 -100.935 64.445 -100.765 ;
      RECT 64.355 -99.73 64.445 -98.722 ;
      RECT 64.305 -99.495 64.445 -99.325 ;
      RECT 64.355 -98.308 64.445 -97.3 ;
      RECT 64.305 -97.705 64.445 -97.535 ;
      RECT 64.355 -96.5 64.445 -95.492 ;
      RECT 64.305 -96.265 64.445 -96.095 ;
      RECT 64.355 -95.078 64.445 -94.07 ;
      RECT 64.305 -94.475 64.445 -94.305 ;
      RECT 64.355 -93.27 64.445 -92.262 ;
      RECT 64.305 -93.035 64.445 -92.865 ;
      RECT 64.355 -91.848 64.445 -90.84 ;
      RECT 64.305 -91.245 64.445 -91.075 ;
      RECT 64.355 -90.04 64.445 -89.032 ;
      RECT 64.305 -89.805 64.445 -89.635 ;
      RECT 64.355 -88.618 64.445 -87.61 ;
      RECT 64.305 -88.015 64.445 -87.845 ;
      RECT 64.355 -86.81 64.445 -85.802 ;
      RECT 64.305 -86.575 64.445 -86.405 ;
      RECT 64.355 -85.388 64.445 -84.38 ;
      RECT 64.305 -84.785 64.445 -84.615 ;
      RECT 64.355 -83.58 64.445 -82.572 ;
      RECT 64.305 -83.345 64.445 -83.175 ;
      RECT 64.355 -82.158 64.445 -81.15 ;
      RECT 64.305 -81.555 64.445 -81.385 ;
      RECT 64.355 -80.35 64.445 -79.342 ;
      RECT 64.305 -80.115 64.445 -79.945 ;
      RECT 64.355 -78.928 64.445 -77.92 ;
      RECT 64.305 -78.325 64.445 -78.155 ;
      RECT 64.355 -77.12 64.445 -76.112 ;
      RECT 64.305 -76.885 64.445 -76.715 ;
      RECT 64.355 -75.698 64.445 -74.69 ;
      RECT 64.305 -75.095 64.445 -74.925 ;
      RECT 64.355 -73.89 64.445 -72.882 ;
      RECT 64.305 -73.655 64.445 -73.485 ;
      RECT 64.355 -72.468 64.445 -71.46 ;
      RECT 64.305 -71.865 64.445 -71.695 ;
      RECT 64.355 -70.66 64.445 -69.652 ;
      RECT 64.305 -70.425 64.445 -70.255 ;
      RECT 64.355 -69.238 64.445 -68.23 ;
      RECT 64.305 -68.635 64.445 -68.465 ;
      RECT 64.355 -67.43 64.445 -66.422 ;
      RECT 64.305 -67.195 64.445 -67.025 ;
      RECT 64.355 -66.008 64.445 -65 ;
      RECT 64.305 -65.405 64.445 -65.235 ;
      RECT 64.355 -64.2 64.445 -63.192 ;
      RECT 64.305 -63.965 64.445 -63.795 ;
      RECT 64.355 -62.778 64.445 -61.77 ;
      RECT 64.305 -62.175 64.445 -62.005 ;
      RECT 64.355 -60.97 64.445 -59.962 ;
      RECT 64.305 -60.735 64.445 -60.565 ;
      RECT 64.355 -59.548 64.445 -58.54 ;
      RECT 64.305 -58.945 64.445 -58.775 ;
      RECT 64.355 -57.74 64.445 -56.732 ;
      RECT 64.305 -57.505 64.445 -57.335 ;
      RECT 64.355 -56.318 64.445 -55.31 ;
      RECT 64.305 -55.715 64.445 -55.545 ;
      RECT 64.355 -54.51 64.445 -53.502 ;
      RECT 64.305 -54.275 64.445 -54.105 ;
      RECT 64.355 -53.088 64.445 -52.08 ;
      RECT 64.305 -52.485 64.445 -52.315 ;
      RECT 64.355 -51.28 64.445 -50.272 ;
      RECT 64.305 -51.045 64.445 -50.875 ;
      RECT 64.355 -49.858 64.445 -48.85 ;
      RECT 64.305 -49.255 64.445 -49.085 ;
      RECT 64.355 -48.05 64.445 -47.042 ;
      RECT 64.305 -47.815 64.445 -47.645 ;
      RECT 64.355 -46.628 64.445 -45.62 ;
      RECT 64.305 -46.025 64.445 -45.855 ;
      RECT 64.355 -44.82 64.445 -43.812 ;
      RECT 64.305 -44.585 64.445 -44.415 ;
      RECT 64.355 -43.398 64.445 -42.39 ;
      RECT 64.305 -42.795 64.445 -42.625 ;
      RECT 64.355 -41.59 64.445 -40.582 ;
      RECT 64.305 -41.355 64.445 -41.185 ;
      RECT 64.355 -40.168 64.445 -39.16 ;
      RECT 64.305 -39.565 64.445 -39.395 ;
      RECT 64.355 -38.36 64.445 -37.352 ;
      RECT 64.305 -38.125 64.445 -37.955 ;
      RECT 64.355 -36.938 64.445 -35.93 ;
      RECT 64.305 -36.335 64.445 -36.165 ;
      RECT 64.355 -35.13 64.445 -34.122 ;
      RECT 64.305 -34.895 64.445 -34.725 ;
      RECT 64.355 -33.708 64.445 -32.7 ;
      RECT 64.305 -33.105 64.445 -32.935 ;
      RECT 64.355 -31.9 64.445 -30.892 ;
      RECT 64.305 -31.665 64.445 -31.495 ;
      RECT 64.355 -30.478 64.445 -29.47 ;
      RECT 64.305 -29.875 64.445 -29.705 ;
      RECT 64.355 -28.67 64.445 -27.662 ;
      RECT 64.305 -28.435 64.445 -28.265 ;
      RECT 64.355 -27.248 64.445 -26.24 ;
      RECT 64.305 -26.645 64.445 -26.475 ;
      RECT 64.355 -25.44 64.445 -24.432 ;
      RECT 64.305 -25.205 64.445 -25.035 ;
      RECT 64.355 -24.018 64.445 -23.01 ;
      RECT 64.305 -23.415 64.445 -23.245 ;
      RECT 64.355 -22.21 64.445 -21.202 ;
      RECT 64.305 -21.975 64.445 -21.805 ;
      RECT 64.355 -20.788 64.445 -19.78 ;
      RECT 64.305 -20.185 64.445 -20.015 ;
      RECT 64.355 -18.98 64.445 -17.972 ;
      RECT 64.305 -18.745 64.445 -18.575 ;
      RECT 64.355 -17.558 64.445 -16.55 ;
      RECT 64.305 -16.955 64.445 -16.785 ;
      RECT 64.355 -15.75 64.445 -14.742 ;
      RECT 64.305 -15.515 64.445 -15.345 ;
      RECT 64.355 -14.328 64.445 -13.32 ;
      RECT 64.305 -13.725 64.445 -13.555 ;
      RECT 64.355 -12.52 64.445 -11.512 ;
      RECT 64.305 -12.285 64.445 -12.115 ;
      RECT 64.355 -11.098 64.445 -10.09 ;
      RECT 64.305 -10.495 64.445 -10.325 ;
      RECT 64.355 -9.29 64.445 -8.282 ;
      RECT 64.305 -9.055 64.445 -8.885 ;
      RECT 64.355 -7.868 64.445 -6.86 ;
      RECT 64.305 -7.265 64.445 -7.095 ;
      RECT 64.355 -6.06 64.445 -5.052 ;
      RECT 64.305 -5.825 64.445 -5.655 ;
      RECT 64.355 -4.638 64.445 -3.63 ;
      RECT 64.305 -4.035 64.445 -3.865 ;
      RECT 64.355 -2.83 64.445 -1.822 ;
      RECT 64.305 -2.595 64.445 -2.425 ;
      RECT 64.355 -1.408 64.445 -0.4 ;
      RECT 64.305 -0.805 64.445 -0.635 ;
      RECT 64.355 0.4 64.445 1.408 ;
      RECT 64.305 0.635 64.445 0.805 ;
      RECT 64.23 -114.685 64.405 -114.515 ;
      RECT 64.305 -114.895 64.405 -114.515 ;
      RECT 63.345 -113.555 63.445 -113.09 ;
      RECT 63.71 -113.555 63.81 -113.1 ;
      RECT 63.345 -113.555 64.19 -113.385 ;
      RECT 63.955 -101.538 64.045 -100.531 ;
      RECT 63.955 -101.225 64.095 -101.055 ;
      RECT 63.955 -99.729 64.045 -98.722 ;
      RECT 63.955 -99.205 64.095 -99.035 ;
      RECT 63.955 -98.308 64.045 -97.301 ;
      RECT 63.955 -97.995 64.095 -97.825 ;
      RECT 63.955 -96.499 64.045 -95.492 ;
      RECT 63.955 -95.975 64.095 -95.805 ;
      RECT 63.955 -95.078 64.045 -94.071 ;
      RECT 63.955 -94.765 64.095 -94.595 ;
      RECT 63.955 -93.269 64.045 -92.262 ;
      RECT 63.955 -92.745 64.095 -92.575 ;
      RECT 63.955 -91.848 64.045 -90.841 ;
      RECT 63.955 -91.535 64.095 -91.365 ;
      RECT 63.955 -90.039 64.045 -89.032 ;
      RECT 63.955 -89.515 64.095 -89.345 ;
      RECT 63.955 -88.618 64.045 -87.611 ;
      RECT 63.955 -88.305 64.095 -88.135 ;
      RECT 63.955 -86.809 64.045 -85.802 ;
      RECT 63.955 -86.285 64.095 -86.115 ;
      RECT 63.955 -85.388 64.045 -84.381 ;
      RECT 63.955 -85.075 64.095 -84.905 ;
      RECT 63.955 -83.579 64.045 -82.572 ;
      RECT 63.955 -83.055 64.095 -82.885 ;
      RECT 63.955 -82.158 64.045 -81.151 ;
      RECT 63.955 -81.845 64.095 -81.675 ;
      RECT 63.955 -80.349 64.045 -79.342 ;
      RECT 63.955 -79.825 64.095 -79.655 ;
      RECT 63.955 -78.928 64.045 -77.921 ;
      RECT 63.955 -78.615 64.095 -78.445 ;
      RECT 63.955 -77.119 64.045 -76.112 ;
      RECT 63.955 -76.595 64.095 -76.425 ;
      RECT 63.955 -75.698 64.045 -74.691 ;
      RECT 63.955 -75.385 64.095 -75.215 ;
      RECT 63.955 -73.889 64.045 -72.882 ;
      RECT 63.955 -73.365 64.095 -73.195 ;
      RECT 63.955 -72.468 64.045 -71.461 ;
      RECT 63.955 -72.155 64.095 -71.985 ;
      RECT 63.955 -70.659 64.045 -69.652 ;
      RECT 63.955 -70.135 64.095 -69.965 ;
      RECT 63.955 -69.238 64.045 -68.231 ;
      RECT 63.955 -68.925 64.095 -68.755 ;
      RECT 63.955 -67.429 64.045 -66.422 ;
      RECT 63.955 -66.905 64.095 -66.735 ;
      RECT 63.955 -66.008 64.045 -65.001 ;
      RECT 63.955 -65.695 64.095 -65.525 ;
      RECT 63.955 -64.199 64.045 -63.192 ;
      RECT 63.955 -63.675 64.095 -63.505 ;
      RECT 63.955 -62.778 64.045 -61.771 ;
      RECT 63.955 -62.465 64.095 -62.295 ;
      RECT 63.955 -60.969 64.045 -59.962 ;
      RECT 63.955 -60.445 64.095 -60.275 ;
      RECT 63.955 -59.548 64.045 -58.541 ;
      RECT 63.955 -59.235 64.095 -59.065 ;
      RECT 63.955 -57.739 64.045 -56.732 ;
      RECT 63.955 -57.215 64.095 -57.045 ;
      RECT 63.955 -56.318 64.045 -55.311 ;
      RECT 63.955 -56.005 64.095 -55.835 ;
      RECT 63.955 -54.509 64.045 -53.502 ;
      RECT 63.955 -53.985 64.095 -53.815 ;
      RECT 63.955 -53.088 64.045 -52.081 ;
      RECT 63.955 -52.775 64.095 -52.605 ;
      RECT 63.955 -51.279 64.045 -50.272 ;
      RECT 63.955 -50.755 64.095 -50.585 ;
      RECT 63.955 -49.858 64.045 -48.851 ;
      RECT 63.955 -49.545 64.095 -49.375 ;
      RECT 63.955 -48.049 64.045 -47.042 ;
      RECT 63.955 -47.525 64.095 -47.355 ;
      RECT 63.955 -46.628 64.045 -45.621 ;
      RECT 63.955 -46.315 64.095 -46.145 ;
      RECT 63.955 -44.819 64.045 -43.812 ;
      RECT 63.955 -44.295 64.095 -44.125 ;
      RECT 63.955 -43.398 64.045 -42.391 ;
      RECT 63.955 -43.085 64.095 -42.915 ;
      RECT 63.955 -41.589 64.045 -40.582 ;
      RECT 63.955 -41.065 64.095 -40.895 ;
      RECT 63.955 -40.168 64.045 -39.161 ;
      RECT 63.955 -39.855 64.095 -39.685 ;
      RECT 63.955 -38.359 64.045 -37.352 ;
      RECT 63.955 -37.835 64.095 -37.665 ;
      RECT 63.955 -36.938 64.045 -35.931 ;
      RECT 63.955 -36.625 64.095 -36.455 ;
      RECT 63.955 -35.129 64.045 -34.122 ;
      RECT 63.955 -34.605 64.095 -34.435 ;
      RECT 63.955 -33.708 64.045 -32.701 ;
      RECT 63.955 -33.395 64.095 -33.225 ;
      RECT 63.955 -31.899 64.045 -30.892 ;
      RECT 63.955 -31.375 64.095 -31.205 ;
      RECT 63.955 -30.478 64.045 -29.471 ;
      RECT 63.955 -30.165 64.095 -29.995 ;
      RECT 63.955 -28.669 64.045 -27.662 ;
      RECT 63.955 -28.145 64.095 -27.975 ;
      RECT 63.955 -27.248 64.045 -26.241 ;
      RECT 63.955 -26.935 64.095 -26.765 ;
      RECT 63.955 -25.439 64.045 -24.432 ;
      RECT 63.955 -24.915 64.095 -24.745 ;
      RECT 63.955 -24.018 64.045 -23.011 ;
      RECT 63.955 -23.705 64.095 -23.535 ;
      RECT 63.955 -22.209 64.045 -21.202 ;
      RECT 63.955 -21.685 64.095 -21.515 ;
      RECT 63.955 -20.788 64.045 -19.781 ;
      RECT 63.955 -20.475 64.095 -20.305 ;
      RECT 63.955 -18.979 64.045 -17.972 ;
      RECT 63.955 -18.455 64.095 -18.285 ;
      RECT 63.955 -17.558 64.045 -16.551 ;
      RECT 63.955 -17.245 64.095 -17.075 ;
      RECT 63.955 -15.749 64.045 -14.742 ;
      RECT 63.955 -15.225 64.095 -15.055 ;
      RECT 63.955 -14.328 64.045 -13.321 ;
      RECT 63.955 -14.015 64.095 -13.845 ;
      RECT 63.955 -12.519 64.045 -11.512 ;
      RECT 63.955 -11.995 64.095 -11.825 ;
      RECT 63.955 -11.098 64.045 -10.091 ;
      RECT 63.955 -10.785 64.095 -10.615 ;
      RECT 63.955 -9.289 64.045 -8.282 ;
      RECT 63.955 -8.765 64.095 -8.595 ;
      RECT 63.955 -7.868 64.045 -6.861 ;
      RECT 63.955 -7.555 64.095 -7.385 ;
      RECT 63.955 -6.059 64.045 -5.052 ;
      RECT 63.955 -5.535 64.095 -5.365 ;
      RECT 63.955 -4.638 64.045 -3.631 ;
      RECT 63.955 -4.325 64.095 -4.155 ;
      RECT 63.955 -2.829 64.045 -1.822 ;
      RECT 63.955 -2.305 64.095 -2.135 ;
      RECT 63.955 -1.408 64.045 -0.401 ;
      RECT 63.955 -1.095 64.095 -0.925 ;
      RECT 63.955 0.401 64.045 1.408 ;
      RECT 63.955 0.925 64.095 1.095 ;
      RECT 63.64 -114.685 63.81 -114.515 ;
      RECT 63.71 -114.895 63.81 -114.515 ;
      RECT 63.155 -101.538 63.245 -100.53 ;
      RECT 63.105 -100.935 63.245 -100.765 ;
      RECT 63.155 -99.73 63.245 -98.722 ;
      RECT 63.105 -99.495 63.245 -99.325 ;
      RECT 63.155 -98.308 63.245 -97.3 ;
      RECT 63.105 -97.705 63.245 -97.535 ;
      RECT 63.155 -96.5 63.245 -95.492 ;
      RECT 63.105 -96.265 63.245 -96.095 ;
      RECT 63.155 -95.078 63.245 -94.07 ;
      RECT 63.105 -94.475 63.245 -94.305 ;
      RECT 63.155 -93.27 63.245 -92.262 ;
      RECT 63.105 -93.035 63.245 -92.865 ;
      RECT 63.155 -91.848 63.245 -90.84 ;
      RECT 63.105 -91.245 63.245 -91.075 ;
      RECT 63.155 -90.04 63.245 -89.032 ;
      RECT 63.105 -89.805 63.245 -89.635 ;
      RECT 63.155 -88.618 63.245 -87.61 ;
      RECT 63.105 -88.015 63.245 -87.845 ;
      RECT 63.155 -86.81 63.245 -85.802 ;
      RECT 63.105 -86.575 63.245 -86.405 ;
      RECT 63.155 -85.388 63.245 -84.38 ;
      RECT 63.105 -84.785 63.245 -84.615 ;
      RECT 63.155 -83.58 63.245 -82.572 ;
      RECT 63.105 -83.345 63.245 -83.175 ;
      RECT 63.155 -82.158 63.245 -81.15 ;
      RECT 63.105 -81.555 63.245 -81.385 ;
      RECT 63.155 -80.35 63.245 -79.342 ;
      RECT 63.105 -80.115 63.245 -79.945 ;
      RECT 63.155 -78.928 63.245 -77.92 ;
      RECT 63.105 -78.325 63.245 -78.155 ;
      RECT 63.155 -77.12 63.245 -76.112 ;
      RECT 63.105 -76.885 63.245 -76.715 ;
      RECT 63.155 -75.698 63.245 -74.69 ;
      RECT 63.105 -75.095 63.245 -74.925 ;
      RECT 63.155 -73.89 63.245 -72.882 ;
      RECT 63.105 -73.655 63.245 -73.485 ;
      RECT 63.155 -72.468 63.245 -71.46 ;
      RECT 63.105 -71.865 63.245 -71.695 ;
      RECT 63.155 -70.66 63.245 -69.652 ;
      RECT 63.105 -70.425 63.245 -70.255 ;
      RECT 63.155 -69.238 63.245 -68.23 ;
      RECT 63.105 -68.635 63.245 -68.465 ;
      RECT 63.155 -67.43 63.245 -66.422 ;
      RECT 63.105 -67.195 63.245 -67.025 ;
      RECT 63.155 -66.008 63.245 -65 ;
      RECT 63.105 -65.405 63.245 -65.235 ;
      RECT 63.155 -64.2 63.245 -63.192 ;
      RECT 63.105 -63.965 63.245 -63.795 ;
      RECT 63.155 -62.778 63.245 -61.77 ;
      RECT 63.105 -62.175 63.245 -62.005 ;
      RECT 63.155 -60.97 63.245 -59.962 ;
      RECT 63.105 -60.735 63.245 -60.565 ;
      RECT 63.155 -59.548 63.245 -58.54 ;
      RECT 63.105 -58.945 63.245 -58.775 ;
      RECT 63.155 -57.74 63.245 -56.732 ;
      RECT 63.105 -57.505 63.245 -57.335 ;
      RECT 63.155 -56.318 63.245 -55.31 ;
      RECT 63.105 -55.715 63.245 -55.545 ;
      RECT 63.155 -54.51 63.245 -53.502 ;
      RECT 63.105 -54.275 63.245 -54.105 ;
      RECT 63.155 -53.088 63.245 -52.08 ;
      RECT 63.105 -52.485 63.245 -52.315 ;
      RECT 63.155 -51.28 63.245 -50.272 ;
      RECT 63.105 -51.045 63.245 -50.875 ;
      RECT 63.155 -49.858 63.245 -48.85 ;
      RECT 63.105 -49.255 63.245 -49.085 ;
      RECT 63.155 -48.05 63.245 -47.042 ;
      RECT 63.105 -47.815 63.245 -47.645 ;
      RECT 63.155 -46.628 63.245 -45.62 ;
      RECT 63.105 -46.025 63.245 -45.855 ;
      RECT 63.155 -44.82 63.245 -43.812 ;
      RECT 63.105 -44.585 63.245 -44.415 ;
      RECT 63.155 -43.398 63.245 -42.39 ;
      RECT 63.105 -42.795 63.245 -42.625 ;
      RECT 63.155 -41.59 63.245 -40.582 ;
      RECT 63.105 -41.355 63.245 -41.185 ;
      RECT 63.155 -40.168 63.245 -39.16 ;
      RECT 63.105 -39.565 63.245 -39.395 ;
      RECT 63.155 -38.36 63.245 -37.352 ;
      RECT 63.105 -38.125 63.245 -37.955 ;
      RECT 63.155 -36.938 63.245 -35.93 ;
      RECT 63.105 -36.335 63.245 -36.165 ;
      RECT 63.155 -35.13 63.245 -34.122 ;
      RECT 63.105 -34.895 63.245 -34.725 ;
      RECT 63.155 -33.708 63.245 -32.7 ;
      RECT 63.105 -33.105 63.245 -32.935 ;
      RECT 63.155 -31.9 63.245 -30.892 ;
      RECT 63.105 -31.665 63.245 -31.495 ;
      RECT 63.155 -30.478 63.245 -29.47 ;
      RECT 63.105 -29.875 63.245 -29.705 ;
      RECT 63.155 -28.67 63.245 -27.662 ;
      RECT 63.105 -28.435 63.245 -28.265 ;
      RECT 63.155 -27.248 63.245 -26.24 ;
      RECT 63.105 -26.645 63.245 -26.475 ;
      RECT 63.155 -25.44 63.245 -24.432 ;
      RECT 63.105 -25.205 63.245 -25.035 ;
      RECT 63.155 -24.018 63.245 -23.01 ;
      RECT 63.105 -23.415 63.245 -23.245 ;
      RECT 63.155 -22.21 63.245 -21.202 ;
      RECT 63.105 -21.975 63.245 -21.805 ;
      RECT 63.155 -20.788 63.245 -19.78 ;
      RECT 63.105 -20.185 63.245 -20.015 ;
      RECT 63.155 -18.98 63.245 -17.972 ;
      RECT 63.105 -18.745 63.245 -18.575 ;
      RECT 63.155 -17.558 63.245 -16.55 ;
      RECT 63.105 -16.955 63.245 -16.785 ;
      RECT 63.155 -15.75 63.245 -14.742 ;
      RECT 63.105 -15.515 63.245 -15.345 ;
      RECT 63.155 -14.328 63.245 -13.32 ;
      RECT 63.105 -13.725 63.245 -13.555 ;
      RECT 63.155 -12.52 63.245 -11.512 ;
      RECT 63.105 -12.285 63.245 -12.115 ;
      RECT 63.155 -11.098 63.245 -10.09 ;
      RECT 63.105 -10.495 63.245 -10.325 ;
      RECT 63.155 -9.29 63.245 -8.282 ;
      RECT 63.105 -9.055 63.245 -8.885 ;
      RECT 63.155 -7.868 63.245 -6.86 ;
      RECT 63.105 -7.265 63.245 -7.095 ;
      RECT 63.155 -6.06 63.245 -5.052 ;
      RECT 63.105 -5.825 63.245 -5.655 ;
      RECT 63.155 -4.638 63.245 -3.63 ;
      RECT 63.105 -4.035 63.245 -3.865 ;
      RECT 63.155 -2.83 63.245 -1.822 ;
      RECT 63.105 -2.595 63.245 -2.425 ;
      RECT 63.155 -1.408 63.245 -0.4 ;
      RECT 63.105 -0.805 63.245 -0.635 ;
      RECT 63.155 0.4 63.245 1.408 ;
      RECT 63.105 0.635 63.245 0.805 ;
      RECT 62.755 -101.538 62.845 -100.531 ;
      RECT 62.755 -101.225 62.895 -101.055 ;
      RECT 62.755 -99.729 62.845 -98.722 ;
      RECT 62.755 -99.205 62.895 -99.035 ;
      RECT 62.755 -98.308 62.845 -97.301 ;
      RECT 62.755 -97.995 62.895 -97.825 ;
      RECT 62.755 -96.499 62.845 -95.492 ;
      RECT 62.755 -95.975 62.895 -95.805 ;
      RECT 62.755 -95.078 62.845 -94.071 ;
      RECT 62.755 -94.765 62.895 -94.595 ;
      RECT 62.755 -93.269 62.845 -92.262 ;
      RECT 62.755 -92.745 62.895 -92.575 ;
      RECT 62.755 -91.848 62.845 -90.841 ;
      RECT 62.755 -91.535 62.895 -91.365 ;
      RECT 62.755 -90.039 62.845 -89.032 ;
      RECT 62.755 -89.515 62.895 -89.345 ;
      RECT 62.755 -88.618 62.845 -87.611 ;
      RECT 62.755 -88.305 62.895 -88.135 ;
      RECT 62.755 -86.809 62.845 -85.802 ;
      RECT 62.755 -86.285 62.895 -86.115 ;
      RECT 62.755 -85.388 62.845 -84.381 ;
      RECT 62.755 -85.075 62.895 -84.905 ;
      RECT 62.755 -83.579 62.845 -82.572 ;
      RECT 62.755 -83.055 62.895 -82.885 ;
      RECT 62.755 -82.158 62.845 -81.151 ;
      RECT 62.755 -81.845 62.895 -81.675 ;
      RECT 62.755 -80.349 62.845 -79.342 ;
      RECT 62.755 -79.825 62.895 -79.655 ;
      RECT 62.755 -78.928 62.845 -77.921 ;
      RECT 62.755 -78.615 62.895 -78.445 ;
      RECT 62.755 -77.119 62.845 -76.112 ;
      RECT 62.755 -76.595 62.895 -76.425 ;
      RECT 62.755 -75.698 62.845 -74.691 ;
      RECT 62.755 -75.385 62.895 -75.215 ;
      RECT 62.755 -73.889 62.845 -72.882 ;
      RECT 62.755 -73.365 62.895 -73.195 ;
      RECT 62.755 -72.468 62.845 -71.461 ;
      RECT 62.755 -72.155 62.895 -71.985 ;
      RECT 62.755 -70.659 62.845 -69.652 ;
      RECT 62.755 -70.135 62.895 -69.965 ;
      RECT 62.755 -69.238 62.845 -68.231 ;
      RECT 62.755 -68.925 62.895 -68.755 ;
      RECT 62.755 -67.429 62.845 -66.422 ;
      RECT 62.755 -66.905 62.895 -66.735 ;
      RECT 62.755 -66.008 62.845 -65.001 ;
      RECT 62.755 -65.695 62.895 -65.525 ;
      RECT 62.755 -64.199 62.845 -63.192 ;
      RECT 62.755 -63.675 62.895 -63.505 ;
      RECT 62.755 -62.778 62.845 -61.771 ;
      RECT 62.755 -62.465 62.895 -62.295 ;
      RECT 62.755 -60.969 62.845 -59.962 ;
      RECT 62.755 -60.445 62.895 -60.275 ;
      RECT 62.755 -59.548 62.845 -58.541 ;
      RECT 62.755 -59.235 62.895 -59.065 ;
      RECT 62.755 -57.739 62.845 -56.732 ;
      RECT 62.755 -57.215 62.895 -57.045 ;
      RECT 62.755 -56.318 62.845 -55.311 ;
      RECT 62.755 -56.005 62.895 -55.835 ;
      RECT 62.755 -54.509 62.845 -53.502 ;
      RECT 62.755 -53.985 62.895 -53.815 ;
      RECT 62.755 -53.088 62.845 -52.081 ;
      RECT 62.755 -52.775 62.895 -52.605 ;
      RECT 62.755 -51.279 62.845 -50.272 ;
      RECT 62.755 -50.755 62.895 -50.585 ;
      RECT 62.755 -49.858 62.845 -48.851 ;
      RECT 62.755 -49.545 62.895 -49.375 ;
      RECT 62.755 -48.049 62.845 -47.042 ;
      RECT 62.755 -47.525 62.895 -47.355 ;
      RECT 62.755 -46.628 62.845 -45.621 ;
      RECT 62.755 -46.315 62.895 -46.145 ;
      RECT 62.755 -44.819 62.845 -43.812 ;
      RECT 62.755 -44.295 62.895 -44.125 ;
      RECT 62.755 -43.398 62.845 -42.391 ;
      RECT 62.755 -43.085 62.895 -42.915 ;
      RECT 62.755 -41.589 62.845 -40.582 ;
      RECT 62.755 -41.065 62.895 -40.895 ;
      RECT 62.755 -40.168 62.845 -39.161 ;
      RECT 62.755 -39.855 62.895 -39.685 ;
      RECT 62.755 -38.359 62.845 -37.352 ;
      RECT 62.755 -37.835 62.895 -37.665 ;
      RECT 62.755 -36.938 62.845 -35.931 ;
      RECT 62.755 -36.625 62.895 -36.455 ;
      RECT 62.755 -35.129 62.845 -34.122 ;
      RECT 62.755 -34.605 62.895 -34.435 ;
      RECT 62.755 -33.708 62.845 -32.701 ;
      RECT 62.755 -33.395 62.895 -33.225 ;
      RECT 62.755 -31.899 62.845 -30.892 ;
      RECT 62.755 -31.375 62.895 -31.205 ;
      RECT 62.755 -30.478 62.845 -29.471 ;
      RECT 62.755 -30.165 62.895 -29.995 ;
      RECT 62.755 -28.669 62.845 -27.662 ;
      RECT 62.755 -28.145 62.895 -27.975 ;
      RECT 62.755 -27.248 62.845 -26.241 ;
      RECT 62.755 -26.935 62.895 -26.765 ;
      RECT 62.755 -25.439 62.845 -24.432 ;
      RECT 62.755 -24.915 62.895 -24.745 ;
      RECT 62.755 -24.018 62.845 -23.011 ;
      RECT 62.755 -23.705 62.895 -23.535 ;
      RECT 62.755 -22.209 62.845 -21.202 ;
      RECT 62.755 -21.685 62.895 -21.515 ;
      RECT 62.755 -20.788 62.845 -19.781 ;
      RECT 62.755 -20.475 62.895 -20.305 ;
      RECT 62.755 -18.979 62.845 -17.972 ;
      RECT 62.755 -18.455 62.895 -18.285 ;
      RECT 62.755 -17.558 62.845 -16.551 ;
      RECT 62.755 -17.245 62.895 -17.075 ;
      RECT 62.755 -15.749 62.845 -14.742 ;
      RECT 62.755 -15.225 62.895 -15.055 ;
      RECT 62.755 -14.328 62.845 -13.321 ;
      RECT 62.755 -14.015 62.895 -13.845 ;
      RECT 62.755 -12.519 62.845 -11.512 ;
      RECT 62.755 -11.995 62.895 -11.825 ;
      RECT 62.755 -11.098 62.845 -10.091 ;
      RECT 62.755 -10.785 62.895 -10.615 ;
      RECT 62.755 -9.289 62.845 -8.282 ;
      RECT 62.755 -8.765 62.895 -8.595 ;
      RECT 62.755 -7.868 62.845 -6.861 ;
      RECT 62.755 -7.555 62.895 -7.385 ;
      RECT 62.755 -6.059 62.845 -5.052 ;
      RECT 62.755 -5.535 62.895 -5.365 ;
      RECT 62.755 -4.638 62.845 -3.631 ;
      RECT 62.755 -4.325 62.895 -4.155 ;
      RECT 62.755 -2.829 62.845 -1.822 ;
      RECT 62.755 -2.305 62.895 -2.135 ;
      RECT 62.755 -1.408 62.845 -0.401 ;
      RECT 62.755 -1.095 62.895 -0.925 ;
      RECT 62.755 0.401 62.845 1.408 ;
      RECT 62.755 0.925 62.895 1.095 ;
      RECT 58.585 -108.935 62.365 -108.815 ;
      RECT 59.905 -109.475 60.005 -108.815 ;
      RECT 59.345 -109.475 59.445 -108.815 ;
      RECT 58.785 -109.475 58.885 -108.815 ;
      RECT 61.955 -101.538 62.045 -100.53 ;
      RECT 61.905 -100.935 62.045 -100.765 ;
      RECT 61.955 -99.73 62.045 -98.722 ;
      RECT 61.905 -99.495 62.045 -99.325 ;
      RECT 61.955 -98.308 62.045 -97.3 ;
      RECT 61.905 -97.705 62.045 -97.535 ;
      RECT 61.955 -96.5 62.045 -95.492 ;
      RECT 61.905 -96.265 62.045 -96.095 ;
      RECT 61.955 -95.078 62.045 -94.07 ;
      RECT 61.905 -94.475 62.045 -94.305 ;
      RECT 61.955 -93.27 62.045 -92.262 ;
      RECT 61.905 -93.035 62.045 -92.865 ;
      RECT 61.955 -91.848 62.045 -90.84 ;
      RECT 61.905 -91.245 62.045 -91.075 ;
      RECT 61.955 -90.04 62.045 -89.032 ;
      RECT 61.905 -89.805 62.045 -89.635 ;
      RECT 61.955 -88.618 62.045 -87.61 ;
      RECT 61.905 -88.015 62.045 -87.845 ;
      RECT 61.955 -86.81 62.045 -85.802 ;
      RECT 61.905 -86.575 62.045 -86.405 ;
      RECT 61.955 -85.388 62.045 -84.38 ;
      RECT 61.905 -84.785 62.045 -84.615 ;
      RECT 61.955 -83.58 62.045 -82.572 ;
      RECT 61.905 -83.345 62.045 -83.175 ;
      RECT 61.955 -82.158 62.045 -81.15 ;
      RECT 61.905 -81.555 62.045 -81.385 ;
      RECT 61.955 -80.35 62.045 -79.342 ;
      RECT 61.905 -80.115 62.045 -79.945 ;
      RECT 61.955 -78.928 62.045 -77.92 ;
      RECT 61.905 -78.325 62.045 -78.155 ;
      RECT 61.955 -77.12 62.045 -76.112 ;
      RECT 61.905 -76.885 62.045 -76.715 ;
      RECT 61.955 -75.698 62.045 -74.69 ;
      RECT 61.905 -75.095 62.045 -74.925 ;
      RECT 61.955 -73.89 62.045 -72.882 ;
      RECT 61.905 -73.655 62.045 -73.485 ;
      RECT 61.955 -72.468 62.045 -71.46 ;
      RECT 61.905 -71.865 62.045 -71.695 ;
      RECT 61.955 -70.66 62.045 -69.652 ;
      RECT 61.905 -70.425 62.045 -70.255 ;
      RECT 61.955 -69.238 62.045 -68.23 ;
      RECT 61.905 -68.635 62.045 -68.465 ;
      RECT 61.955 -67.43 62.045 -66.422 ;
      RECT 61.905 -67.195 62.045 -67.025 ;
      RECT 61.955 -66.008 62.045 -65 ;
      RECT 61.905 -65.405 62.045 -65.235 ;
      RECT 61.955 -64.2 62.045 -63.192 ;
      RECT 61.905 -63.965 62.045 -63.795 ;
      RECT 61.955 -62.778 62.045 -61.77 ;
      RECT 61.905 -62.175 62.045 -62.005 ;
      RECT 61.955 -60.97 62.045 -59.962 ;
      RECT 61.905 -60.735 62.045 -60.565 ;
      RECT 61.955 -59.548 62.045 -58.54 ;
      RECT 61.905 -58.945 62.045 -58.775 ;
      RECT 61.955 -57.74 62.045 -56.732 ;
      RECT 61.905 -57.505 62.045 -57.335 ;
      RECT 61.955 -56.318 62.045 -55.31 ;
      RECT 61.905 -55.715 62.045 -55.545 ;
      RECT 61.955 -54.51 62.045 -53.502 ;
      RECT 61.905 -54.275 62.045 -54.105 ;
      RECT 61.955 -53.088 62.045 -52.08 ;
      RECT 61.905 -52.485 62.045 -52.315 ;
      RECT 61.955 -51.28 62.045 -50.272 ;
      RECT 61.905 -51.045 62.045 -50.875 ;
      RECT 61.955 -49.858 62.045 -48.85 ;
      RECT 61.905 -49.255 62.045 -49.085 ;
      RECT 61.955 -48.05 62.045 -47.042 ;
      RECT 61.905 -47.815 62.045 -47.645 ;
      RECT 61.955 -46.628 62.045 -45.62 ;
      RECT 61.905 -46.025 62.045 -45.855 ;
      RECT 61.955 -44.82 62.045 -43.812 ;
      RECT 61.905 -44.585 62.045 -44.415 ;
      RECT 61.955 -43.398 62.045 -42.39 ;
      RECT 61.905 -42.795 62.045 -42.625 ;
      RECT 61.955 -41.59 62.045 -40.582 ;
      RECT 61.905 -41.355 62.045 -41.185 ;
      RECT 61.955 -40.168 62.045 -39.16 ;
      RECT 61.905 -39.565 62.045 -39.395 ;
      RECT 61.955 -38.36 62.045 -37.352 ;
      RECT 61.905 -38.125 62.045 -37.955 ;
      RECT 61.955 -36.938 62.045 -35.93 ;
      RECT 61.905 -36.335 62.045 -36.165 ;
      RECT 61.955 -35.13 62.045 -34.122 ;
      RECT 61.905 -34.895 62.045 -34.725 ;
      RECT 61.955 -33.708 62.045 -32.7 ;
      RECT 61.905 -33.105 62.045 -32.935 ;
      RECT 61.955 -31.9 62.045 -30.892 ;
      RECT 61.905 -31.665 62.045 -31.495 ;
      RECT 61.955 -30.478 62.045 -29.47 ;
      RECT 61.905 -29.875 62.045 -29.705 ;
      RECT 61.955 -28.67 62.045 -27.662 ;
      RECT 61.905 -28.435 62.045 -28.265 ;
      RECT 61.955 -27.248 62.045 -26.24 ;
      RECT 61.905 -26.645 62.045 -26.475 ;
      RECT 61.955 -25.44 62.045 -24.432 ;
      RECT 61.905 -25.205 62.045 -25.035 ;
      RECT 61.955 -24.018 62.045 -23.01 ;
      RECT 61.905 -23.415 62.045 -23.245 ;
      RECT 61.955 -22.21 62.045 -21.202 ;
      RECT 61.905 -21.975 62.045 -21.805 ;
      RECT 61.955 -20.788 62.045 -19.78 ;
      RECT 61.905 -20.185 62.045 -20.015 ;
      RECT 61.955 -18.98 62.045 -17.972 ;
      RECT 61.905 -18.745 62.045 -18.575 ;
      RECT 61.955 -17.558 62.045 -16.55 ;
      RECT 61.905 -16.955 62.045 -16.785 ;
      RECT 61.955 -15.75 62.045 -14.742 ;
      RECT 61.905 -15.515 62.045 -15.345 ;
      RECT 61.955 -14.328 62.045 -13.32 ;
      RECT 61.905 -13.725 62.045 -13.555 ;
      RECT 61.955 -12.52 62.045 -11.512 ;
      RECT 61.905 -12.285 62.045 -12.115 ;
      RECT 61.955 -11.098 62.045 -10.09 ;
      RECT 61.905 -10.495 62.045 -10.325 ;
      RECT 61.955 -9.29 62.045 -8.282 ;
      RECT 61.905 -9.055 62.045 -8.885 ;
      RECT 61.955 -7.868 62.045 -6.86 ;
      RECT 61.905 -7.265 62.045 -7.095 ;
      RECT 61.955 -6.06 62.045 -5.052 ;
      RECT 61.905 -5.825 62.045 -5.655 ;
      RECT 61.955 -4.638 62.045 -3.63 ;
      RECT 61.905 -4.035 62.045 -3.865 ;
      RECT 61.955 -2.83 62.045 -1.822 ;
      RECT 61.905 -2.595 62.045 -2.425 ;
      RECT 61.955 -1.408 62.045 -0.4 ;
      RECT 61.905 -0.805 62.045 -0.635 ;
      RECT 61.955 0.4 62.045 1.408 ;
      RECT 61.905 0.635 62.045 0.805 ;
      RECT 60.525 -111.685 62.005 -111.585 ;
      RECT 60.525 -112.195 60.625 -111.585 ;
      RECT 60.745 -109.15 62.005 -109.05 ;
      RECT 61.905 -109.475 62.005 -109.05 ;
      RECT 61.345 -109.475 61.445 -109.05 ;
      RECT 60.785 -109.475 60.885 -109.05 ;
      RECT 61.555 -101.538 61.645 -100.531 ;
      RECT 61.555 -101.225 61.695 -101.055 ;
      RECT 61.555 -99.729 61.645 -98.722 ;
      RECT 61.555 -99.205 61.695 -99.035 ;
      RECT 61.555 -98.308 61.645 -97.301 ;
      RECT 61.555 -97.995 61.695 -97.825 ;
      RECT 61.555 -96.499 61.645 -95.492 ;
      RECT 61.555 -95.975 61.695 -95.805 ;
      RECT 61.555 -95.078 61.645 -94.071 ;
      RECT 61.555 -94.765 61.695 -94.595 ;
      RECT 61.555 -93.269 61.645 -92.262 ;
      RECT 61.555 -92.745 61.695 -92.575 ;
      RECT 61.555 -91.848 61.645 -90.841 ;
      RECT 61.555 -91.535 61.695 -91.365 ;
      RECT 61.555 -90.039 61.645 -89.032 ;
      RECT 61.555 -89.515 61.695 -89.345 ;
      RECT 61.555 -88.618 61.645 -87.611 ;
      RECT 61.555 -88.305 61.695 -88.135 ;
      RECT 61.555 -86.809 61.645 -85.802 ;
      RECT 61.555 -86.285 61.695 -86.115 ;
      RECT 61.555 -85.388 61.645 -84.381 ;
      RECT 61.555 -85.075 61.695 -84.905 ;
      RECT 61.555 -83.579 61.645 -82.572 ;
      RECT 61.555 -83.055 61.695 -82.885 ;
      RECT 61.555 -82.158 61.645 -81.151 ;
      RECT 61.555 -81.845 61.695 -81.675 ;
      RECT 61.555 -80.349 61.645 -79.342 ;
      RECT 61.555 -79.825 61.695 -79.655 ;
      RECT 61.555 -78.928 61.645 -77.921 ;
      RECT 61.555 -78.615 61.695 -78.445 ;
      RECT 61.555 -77.119 61.645 -76.112 ;
      RECT 61.555 -76.595 61.695 -76.425 ;
      RECT 61.555 -75.698 61.645 -74.691 ;
      RECT 61.555 -75.385 61.695 -75.215 ;
      RECT 61.555 -73.889 61.645 -72.882 ;
      RECT 61.555 -73.365 61.695 -73.195 ;
      RECT 61.555 -72.468 61.645 -71.461 ;
      RECT 61.555 -72.155 61.695 -71.985 ;
      RECT 61.555 -70.659 61.645 -69.652 ;
      RECT 61.555 -70.135 61.695 -69.965 ;
      RECT 61.555 -69.238 61.645 -68.231 ;
      RECT 61.555 -68.925 61.695 -68.755 ;
      RECT 61.555 -67.429 61.645 -66.422 ;
      RECT 61.555 -66.905 61.695 -66.735 ;
      RECT 61.555 -66.008 61.645 -65.001 ;
      RECT 61.555 -65.695 61.695 -65.525 ;
      RECT 61.555 -64.199 61.645 -63.192 ;
      RECT 61.555 -63.675 61.695 -63.505 ;
      RECT 61.555 -62.778 61.645 -61.771 ;
      RECT 61.555 -62.465 61.695 -62.295 ;
      RECT 61.555 -60.969 61.645 -59.962 ;
      RECT 61.555 -60.445 61.695 -60.275 ;
      RECT 61.555 -59.548 61.645 -58.541 ;
      RECT 61.555 -59.235 61.695 -59.065 ;
      RECT 61.555 -57.739 61.645 -56.732 ;
      RECT 61.555 -57.215 61.695 -57.045 ;
      RECT 61.555 -56.318 61.645 -55.311 ;
      RECT 61.555 -56.005 61.695 -55.835 ;
      RECT 61.555 -54.509 61.645 -53.502 ;
      RECT 61.555 -53.985 61.695 -53.815 ;
      RECT 61.555 -53.088 61.645 -52.081 ;
      RECT 61.555 -52.775 61.695 -52.605 ;
      RECT 61.555 -51.279 61.645 -50.272 ;
      RECT 61.555 -50.755 61.695 -50.585 ;
      RECT 61.555 -49.858 61.645 -48.851 ;
      RECT 61.555 -49.545 61.695 -49.375 ;
      RECT 61.555 -48.049 61.645 -47.042 ;
      RECT 61.555 -47.525 61.695 -47.355 ;
      RECT 61.555 -46.628 61.645 -45.621 ;
      RECT 61.555 -46.315 61.695 -46.145 ;
      RECT 61.555 -44.819 61.645 -43.812 ;
      RECT 61.555 -44.295 61.695 -44.125 ;
      RECT 61.555 -43.398 61.645 -42.391 ;
      RECT 61.555 -43.085 61.695 -42.915 ;
      RECT 61.555 -41.589 61.645 -40.582 ;
      RECT 61.555 -41.065 61.695 -40.895 ;
      RECT 61.555 -40.168 61.645 -39.161 ;
      RECT 61.555 -39.855 61.695 -39.685 ;
      RECT 61.555 -38.359 61.645 -37.352 ;
      RECT 61.555 -37.835 61.695 -37.665 ;
      RECT 61.555 -36.938 61.645 -35.931 ;
      RECT 61.555 -36.625 61.695 -36.455 ;
      RECT 61.555 -35.129 61.645 -34.122 ;
      RECT 61.555 -34.605 61.695 -34.435 ;
      RECT 61.555 -33.708 61.645 -32.701 ;
      RECT 61.555 -33.395 61.695 -33.225 ;
      RECT 61.555 -31.899 61.645 -30.892 ;
      RECT 61.555 -31.375 61.695 -31.205 ;
      RECT 61.555 -30.478 61.645 -29.471 ;
      RECT 61.555 -30.165 61.695 -29.995 ;
      RECT 61.555 -28.669 61.645 -27.662 ;
      RECT 61.555 -28.145 61.695 -27.975 ;
      RECT 61.555 -27.248 61.645 -26.241 ;
      RECT 61.555 -26.935 61.695 -26.765 ;
      RECT 61.555 -25.439 61.645 -24.432 ;
      RECT 61.555 -24.915 61.695 -24.745 ;
      RECT 61.555 -24.018 61.645 -23.011 ;
      RECT 61.555 -23.705 61.695 -23.535 ;
      RECT 61.555 -22.209 61.645 -21.202 ;
      RECT 61.555 -21.685 61.695 -21.515 ;
      RECT 61.555 -20.788 61.645 -19.781 ;
      RECT 61.555 -20.475 61.695 -20.305 ;
      RECT 61.555 -18.979 61.645 -17.972 ;
      RECT 61.555 -18.455 61.695 -18.285 ;
      RECT 61.555 -17.558 61.645 -16.551 ;
      RECT 61.555 -17.245 61.695 -17.075 ;
      RECT 61.555 -15.749 61.645 -14.742 ;
      RECT 61.555 -15.225 61.695 -15.055 ;
      RECT 61.555 -14.328 61.645 -13.321 ;
      RECT 61.555 -14.015 61.695 -13.845 ;
      RECT 61.555 -12.519 61.645 -11.512 ;
      RECT 61.555 -11.995 61.695 -11.825 ;
      RECT 61.555 -11.098 61.645 -10.091 ;
      RECT 61.555 -10.785 61.695 -10.615 ;
      RECT 61.555 -9.289 61.645 -8.282 ;
      RECT 61.555 -8.765 61.695 -8.595 ;
      RECT 61.555 -7.868 61.645 -6.861 ;
      RECT 61.555 -7.555 61.695 -7.385 ;
      RECT 61.555 -6.059 61.645 -5.052 ;
      RECT 61.555 -5.535 61.695 -5.365 ;
      RECT 61.555 -4.638 61.645 -3.631 ;
      RECT 61.555 -4.325 61.695 -4.155 ;
      RECT 61.555 -2.829 61.645 -1.822 ;
      RECT 61.555 -2.305 61.695 -2.135 ;
      RECT 61.555 -1.408 61.645 -0.401 ;
      RECT 61.555 -1.095 61.695 -0.925 ;
      RECT 61.555 0.401 61.645 1.408 ;
      RECT 61.555 0.925 61.695 1.095 ;
      RECT 60.885 -111.495 61.055 -111.385 ;
      RECT 57.735 -111.495 61.055 -111.395 ;
      RECT 60.755 -101.538 60.845 -100.53 ;
      RECT 60.705 -100.935 60.845 -100.765 ;
      RECT 60.755 -99.73 60.845 -98.722 ;
      RECT 60.705 -99.495 60.845 -99.325 ;
      RECT 60.755 -98.308 60.845 -97.3 ;
      RECT 60.705 -97.705 60.845 -97.535 ;
      RECT 60.755 -96.5 60.845 -95.492 ;
      RECT 60.705 -96.265 60.845 -96.095 ;
      RECT 60.755 -95.078 60.845 -94.07 ;
      RECT 60.705 -94.475 60.845 -94.305 ;
      RECT 60.755 -93.27 60.845 -92.262 ;
      RECT 60.705 -93.035 60.845 -92.865 ;
      RECT 60.755 -91.848 60.845 -90.84 ;
      RECT 60.705 -91.245 60.845 -91.075 ;
      RECT 60.755 -90.04 60.845 -89.032 ;
      RECT 60.705 -89.805 60.845 -89.635 ;
      RECT 60.755 -88.618 60.845 -87.61 ;
      RECT 60.705 -88.015 60.845 -87.845 ;
      RECT 60.755 -86.81 60.845 -85.802 ;
      RECT 60.705 -86.575 60.845 -86.405 ;
      RECT 60.755 -85.388 60.845 -84.38 ;
      RECT 60.705 -84.785 60.845 -84.615 ;
      RECT 60.755 -83.58 60.845 -82.572 ;
      RECT 60.705 -83.345 60.845 -83.175 ;
      RECT 60.755 -82.158 60.845 -81.15 ;
      RECT 60.705 -81.555 60.845 -81.385 ;
      RECT 60.755 -80.35 60.845 -79.342 ;
      RECT 60.705 -80.115 60.845 -79.945 ;
      RECT 60.755 -78.928 60.845 -77.92 ;
      RECT 60.705 -78.325 60.845 -78.155 ;
      RECT 60.755 -77.12 60.845 -76.112 ;
      RECT 60.705 -76.885 60.845 -76.715 ;
      RECT 60.755 -75.698 60.845 -74.69 ;
      RECT 60.705 -75.095 60.845 -74.925 ;
      RECT 60.755 -73.89 60.845 -72.882 ;
      RECT 60.705 -73.655 60.845 -73.485 ;
      RECT 60.755 -72.468 60.845 -71.46 ;
      RECT 60.705 -71.865 60.845 -71.695 ;
      RECT 60.755 -70.66 60.845 -69.652 ;
      RECT 60.705 -70.425 60.845 -70.255 ;
      RECT 60.755 -69.238 60.845 -68.23 ;
      RECT 60.705 -68.635 60.845 -68.465 ;
      RECT 60.755 -67.43 60.845 -66.422 ;
      RECT 60.705 -67.195 60.845 -67.025 ;
      RECT 60.755 -66.008 60.845 -65 ;
      RECT 60.705 -65.405 60.845 -65.235 ;
      RECT 60.755 -64.2 60.845 -63.192 ;
      RECT 60.705 -63.965 60.845 -63.795 ;
      RECT 60.755 -62.778 60.845 -61.77 ;
      RECT 60.705 -62.175 60.845 -62.005 ;
      RECT 60.755 -60.97 60.845 -59.962 ;
      RECT 60.705 -60.735 60.845 -60.565 ;
      RECT 60.755 -59.548 60.845 -58.54 ;
      RECT 60.705 -58.945 60.845 -58.775 ;
      RECT 60.755 -57.74 60.845 -56.732 ;
      RECT 60.705 -57.505 60.845 -57.335 ;
      RECT 60.755 -56.318 60.845 -55.31 ;
      RECT 60.705 -55.715 60.845 -55.545 ;
      RECT 60.755 -54.51 60.845 -53.502 ;
      RECT 60.705 -54.275 60.845 -54.105 ;
      RECT 60.755 -53.088 60.845 -52.08 ;
      RECT 60.705 -52.485 60.845 -52.315 ;
      RECT 60.755 -51.28 60.845 -50.272 ;
      RECT 60.705 -51.045 60.845 -50.875 ;
      RECT 60.755 -49.858 60.845 -48.85 ;
      RECT 60.705 -49.255 60.845 -49.085 ;
      RECT 60.755 -48.05 60.845 -47.042 ;
      RECT 60.705 -47.815 60.845 -47.645 ;
      RECT 60.755 -46.628 60.845 -45.62 ;
      RECT 60.705 -46.025 60.845 -45.855 ;
      RECT 60.755 -44.82 60.845 -43.812 ;
      RECT 60.705 -44.585 60.845 -44.415 ;
      RECT 60.755 -43.398 60.845 -42.39 ;
      RECT 60.705 -42.795 60.845 -42.625 ;
      RECT 60.755 -41.59 60.845 -40.582 ;
      RECT 60.705 -41.355 60.845 -41.185 ;
      RECT 60.755 -40.168 60.845 -39.16 ;
      RECT 60.705 -39.565 60.845 -39.395 ;
      RECT 60.755 -38.36 60.845 -37.352 ;
      RECT 60.705 -38.125 60.845 -37.955 ;
      RECT 60.755 -36.938 60.845 -35.93 ;
      RECT 60.705 -36.335 60.845 -36.165 ;
      RECT 60.755 -35.13 60.845 -34.122 ;
      RECT 60.705 -34.895 60.845 -34.725 ;
      RECT 60.755 -33.708 60.845 -32.7 ;
      RECT 60.705 -33.105 60.845 -32.935 ;
      RECT 60.755 -31.9 60.845 -30.892 ;
      RECT 60.705 -31.665 60.845 -31.495 ;
      RECT 60.755 -30.478 60.845 -29.47 ;
      RECT 60.705 -29.875 60.845 -29.705 ;
      RECT 60.755 -28.67 60.845 -27.662 ;
      RECT 60.705 -28.435 60.845 -28.265 ;
      RECT 60.755 -27.248 60.845 -26.24 ;
      RECT 60.705 -26.645 60.845 -26.475 ;
      RECT 60.755 -25.44 60.845 -24.432 ;
      RECT 60.705 -25.205 60.845 -25.035 ;
      RECT 60.755 -24.018 60.845 -23.01 ;
      RECT 60.705 -23.415 60.845 -23.245 ;
      RECT 60.755 -22.21 60.845 -21.202 ;
      RECT 60.705 -21.975 60.845 -21.805 ;
      RECT 60.755 -20.788 60.845 -19.78 ;
      RECT 60.705 -20.185 60.845 -20.015 ;
      RECT 60.755 -18.98 60.845 -17.972 ;
      RECT 60.705 -18.745 60.845 -18.575 ;
      RECT 60.755 -17.558 60.845 -16.55 ;
      RECT 60.705 -16.955 60.845 -16.785 ;
      RECT 60.755 -15.75 60.845 -14.742 ;
      RECT 60.705 -15.515 60.845 -15.345 ;
      RECT 60.755 -14.328 60.845 -13.32 ;
      RECT 60.705 -13.725 60.845 -13.555 ;
      RECT 60.755 -12.52 60.845 -11.512 ;
      RECT 60.705 -12.285 60.845 -12.115 ;
      RECT 60.755 -11.098 60.845 -10.09 ;
      RECT 60.705 -10.495 60.845 -10.325 ;
      RECT 60.755 -9.29 60.845 -8.282 ;
      RECT 60.705 -9.055 60.845 -8.885 ;
      RECT 60.755 -7.868 60.845 -6.86 ;
      RECT 60.705 -7.265 60.845 -7.095 ;
      RECT 60.755 -6.06 60.845 -5.052 ;
      RECT 60.705 -5.825 60.845 -5.655 ;
      RECT 60.755 -4.638 60.845 -3.63 ;
      RECT 60.705 -4.035 60.845 -3.865 ;
      RECT 60.755 -2.83 60.845 -1.822 ;
      RECT 60.705 -2.595 60.845 -2.425 ;
      RECT 60.755 -1.408 60.845 -0.4 ;
      RECT 60.705 -0.805 60.845 -0.635 ;
      RECT 60.755 0.4 60.845 1.408 ;
      RECT 60.705 0.635 60.845 0.805 ;
      RECT 60.355 -101.538 60.445 -100.531 ;
      RECT 60.355 -101.225 60.495 -101.055 ;
      RECT 60.355 -99.729 60.445 -98.722 ;
      RECT 60.355 -99.205 60.495 -99.035 ;
      RECT 60.355 -98.308 60.445 -97.301 ;
      RECT 60.355 -97.995 60.495 -97.825 ;
      RECT 60.355 -96.499 60.445 -95.492 ;
      RECT 60.355 -95.975 60.495 -95.805 ;
      RECT 60.355 -95.078 60.445 -94.071 ;
      RECT 60.355 -94.765 60.495 -94.595 ;
      RECT 60.355 -93.269 60.445 -92.262 ;
      RECT 60.355 -92.745 60.495 -92.575 ;
      RECT 60.355 -91.848 60.445 -90.841 ;
      RECT 60.355 -91.535 60.495 -91.365 ;
      RECT 60.355 -90.039 60.445 -89.032 ;
      RECT 60.355 -89.515 60.495 -89.345 ;
      RECT 60.355 -88.618 60.445 -87.611 ;
      RECT 60.355 -88.305 60.495 -88.135 ;
      RECT 60.355 -86.809 60.445 -85.802 ;
      RECT 60.355 -86.285 60.495 -86.115 ;
      RECT 60.355 -85.388 60.445 -84.381 ;
      RECT 60.355 -85.075 60.495 -84.905 ;
      RECT 60.355 -83.579 60.445 -82.572 ;
      RECT 60.355 -83.055 60.495 -82.885 ;
      RECT 60.355 -82.158 60.445 -81.151 ;
      RECT 60.355 -81.845 60.495 -81.675 ;
      RECT 60.355 -80.349 60.445 -79.342 ;
      RECT 60.355 -79.825 60.495 -79.655 ;
      RECT 60.355 -78.928 60.445 -77.921 ;
      RECT 60.355 -78.615 60.495 -78.445 ;
      RECT 60.355 -77.119 60.445 -76.112 ;
      RECT 60.355 -76.595 60.495 -76.425 ;
      RECT 60.355 -75.698 60.445 -74.691 ;
      RECT 60.355 -75.385 60.495 -75.215 ;
      RECT 60.355 -73.889 60.445 -72.882 ;
      RECT 60.355 -73.365 60.495 -73.195 ;
      RECT 60.355 -72.468 60.445 -71.461 ;
      RECT 60.355 -72.155 60.495 -71.985 ;
      RECT 60.355 -70.659 60.445 -69.652 ;
      RECT 60.355 -70.135 60.495 -69.965 ;
      RECT 60.355 -69.238 60.445 -68.231 ;
      RECT 60.355 -68.925 60.495 -68.755 ;
      RECT 60.355 -67.429 60.445 -66.422 ;
      RECT 60.355 -66.905 60.495 -66.735 ;
      RECT 60.355 -66.008 60.445 -65.001 ;
      RECT 60.355 -65.695 60.495 -65.525 ;
      RECT 60.355 -64.199 60.445 -63.192 ;
      RECT 60.355 -63.675 60.495 -63.505 ;
      RECT 60.355 -62.778 60.445 -61.771 ;
      RECT 60.355 -62.465 60.495 -62.295 ;
      RECT 60.355 -60.969 60.445 -59.962 ;
      RECT 60.355 -60.445 60.495 -60.275 ;
      RECT 60.355 -59.548 60.445 -58.541 ;
      RECT 60.355 -59.235 60.495 -59.065 ;
      RECT 60.355 -57.739 60.445 -56.732 ;
      RECT 60.355 -57.215 60.495 -57.045 ;
      RECT 60.355 -56.318 60.445 -55.311 ;
      RECT 60.355 -56.005 60.495 -55.835 ;
      RECT 60.355 -54.509 60.445 -53.502 ;
      RECT 60.355 -53.985 60.495 -53.815 ;
      RECT 60.355 -53.088 60.445 -52.081 ;
      RECT 60.355 -52.775 60.495 -52.605 ;
      RECT 60.355 -51.279 60.445 -50.272 ;
      RECT 60.355 -50.755 60.495 -50.585 ;
      RECT 60.355 -49.858 60.445 -48.851 ;
      RECT 60.355 -49.545 60.495 -49.375 ;
      RECT 60.355 -48.049 60.445 -47.042 ;
      RECT 60.355 -47.525 60.495 -47.355 ;
      RECT 60.355 -46.628 60.445 -45.621 ;
      RECT 60.355 -46.315 60.495 -46.145 ;
      RECT 60.355 -44.819 60.445 -43.812 ;
      RECT 60.355 -44.295 60.495 -44.125 ;
      RECT 60.355 -43.398 60.445 -42.391 ;
      RECT 60.355 -43.085 60.495 -42.915 ;
      RECT 60.355 -41.589 60.445 -40.582 ;
      RECT 60.355 -41.065 60.495 -40.895 ;
      RECT 60.355 -40.168 60.445 -39.161 ;
      RECT 60.355 -39.855 60.495 -39.685 ;
      RECT 60.355 -38.359 60.445 -37.352 ;
      RECT 60.355 -37.835 60.495 -37.665 ;
      RECT 60.355 -36.938 60.445 -35.931 ;
      RECT 60.355 -36.625 60.495 -36.455 ;
      RECT 60.355 -35.129 60.445 -34.122 ;
      RECT 60.355 -34.605 60.495 -34.435 ;
      RECT 60.355 -33.708 60.445 -32.701 ;
      RECT 60.355 -33.395 60.495 -33.225 ;
      RECT 60.355 -31.899 60.445 -30.892 ;
      RECT 60.355 -31.375 60.495 -31.205 ;
      RECT 60.355 -30.478 60.445 -29.471 ;
      RECT 60.355 -30.165 60.495 -29.995 ;
      RECT 60.355 -28.669 60.445 -27.662 ;
      RECT 60.355 -28.145 60.495 -27.975 ;
      RECT 60.355 -27.248 60.445 -26.241 ;
      RECT 60.355 -26.935 60.495 -26.765 ;
      RECT 60.355 -25.439 60.445 -24.432 ;
      RECT 60.355 -24.915 60.495 -24.745 ;
      RECT 60.355 -24.018 60.445 -23.011 ;
      RECT 60.355 -23.705 60.495 -23.535 ;
      RECT 60.355 -22.209 60.445 -21.202 ;
      RECT 60.355 -21.685 60.495 -21.515 ;
      RECT 60.355 -20.788 60.445 -19.781 ;
      RECT 60.355 -20.475 60.495 -20.305 ;
      RECT 60.355 -18.979 60.445 -17.972 ;
      RECT 60.355 -18.455 60.495 -18.285 ;
      RECT 60.355 -17.558 60.445 -16.551 ;
      RECT 60.355 -17.245 60.495 -17.075 ;
      RECT 60.355 -15.749 60.445 -14.742 ;
      RECT 60.355 -15.225 60.495 -15.055 ;
      RECT 60.355 -14.328 60.445 -13.321 ;
      RECT 60.355 -14.015 60.495 -13.845 ;
      RECT 60.355 -12.519 60.445 -11.512 ;
      RECT 60.355 -11.995 60.495 -11.825 ;
      RECT 60.355 -11.098 60.445 -10.091 ;
      RECT 60.355 -10.785 60.495 -10.615 ;
      RECT 60.355 -9.289 60.445 -8.282 ;
      RECT 60.355 -8.765 60.495 -8.595 ;
      RECT 60.355 -7.868 60.445 -6.861 ;
      RECT 60.355 -7.555 60.495 -7.385 ;
      RECT 60.355 -6.059 60.445 -5.052 ;
      RECT 60.355 -5.535 60.495 -5.365 ;
      RECT 60.355 -4.638 60.445 -3.631 ;
      RECT 60.355 -4.325 60.495 -4.155 ;
      RECT 60.355 -2.829 60.445 -1.822 ;
      RECT 60.355 -2.305 60.495 -2.135 ;
      RECT 60.355 -1.408 60.445 -0.401 ;
      RECT 60.355 -1.095 60.495 -0.925 ;
      RECT 60.355 0.401 60.445 1.408 ;
      RECT 60.355 0.925 60.495 1.095 ;
      RECT 58.505 -111.685 59.985 -111.585 ;
      RECT 58.505 -112.055 58.605 -111.585 ;
      RECT 58.31 -114.395 59.885 -114.275 ;
      RECT 59.785 -114.895 59.885 -114.275 ;
      RECT 59.19 -114.895 59.29 -114.275 ;
      RECT 58.31 -114.85 58.41 -114.275 ;
      RECT 59.555 -101.538 59.645 -100.53 ;
      RECT 59.505 -100.935 59.645 -100.765 ;
      RECT 59.555 -99.73 59.645 -98.722 ;
      RECT 59.505 -99.495 59.645 -99.325 ;
      RECT 59.555 -98.308 59.645 -97.3 ;
      RECT 59.505 -97.705 59.645 -97.535 ;
      RECT 59.555 -96.5 59.645 -95.492 ;
      RECT 59.505 -96.265 59.645 -96.095 ;
      RECT 59.555 -95.078 59.645 -94.07 ;
      RECT 59.505 -94.475 59.645 -94.305 ;
      RECT 59.555 -93.27 59.645 -92.262 ;
      RECT 59.505 -93.035 59.645 -92.865 ;
      RECT 59.555 -91.848 59.645 -90.84 ;
      RECT 59.505 -91.245 59.645 -91.075 ;
      RECT 59.555 -90.04 59.645 -89.032 ;
      RECT 59.505 -89.805 59.645 -89.635 ;
      RECT 59.555 -88.618 59.645 -87.61 ;
      RECT 59.505 -88.015 59.645 -87.845 ;
      RECT 59.555 -86.81 59.645 -85.802 ;
      RECT 59.505 -86.575 59.645 -86.405 ;
      RECT 59.555 -85.388 59.645 -84.38 ;
      RECT 59.505 -84.785 59.645 -84.615 ;
      RECT 59.555 -83.58 59.645 -82.572 ;
      RECT 59.505 -83.345 59.645 -83.175 ;
      RECT 59.555 -82.158 59.645 -81.15 ;
      RECT 59.505 -81.555 59.645 -81.385 ;
      RECT 59.555 -80.35 59.645 -79.342 ;
      RECT 59.505 -80.115 59.645 -79.945 ;
      RECT 59.555 -78.928 59.645 -77.92 ;
      RECT 59.505 -78.325 59.645 -78.155 ;
      RECT 59.555 -77.12 59.645 -76.112 ;
      RECT 59.505 -76.885 59.645 -76.715 ;
      RECT 59.555 -75.698 59.645 -74.69 ;
      RECT 59.505 -75.095 59.645 -74.925 ;
      RECT 59.555 -73.89 59.645 -72.882 ;
      RECT 59.505 -73.655 59.645 -73.485 ;
      RECT 59.555 -72.468 59.645 -71.46 ;
      RECT 59.505 -71.865 59.645 -71.695 ;
      RECT 59.555 -70.66 59.645 -69.652 ;
      RECT 59.505 -70.425 59.645 -70.255 ;
      RECT 59.555 -69.238 59.645 -68.23 ;
      RECT 59.505 -68.635 59.645 -68.465 ;
      RECT 59.555 -67.43 59.645 -66.422 ;
      RECT 59.505 -67.195 59.645 -67.025 ;
      RECT 59.555 -66.008 59.645 -65 ;
      RECT 59.505 -65.405 59.645 -65.235 ;
      RECT 59.555 -64.2 59.645 -63.192 ;
      RECT 59.505 -63.965 59.645 -63.795 ;
      RECT 59.555 -62.778 59.645 -61.77 ;
      RECT 59.505 -62.175 59.645 -62.005 ;
      RECT 59.555 -60.97 59.645 -59.962 ;
      RECT 59.505 -60.735 59.645 -60.565 ;
      RECT 59.555 -59.548 59.645 -58.54 ;
      RECT 59.505 -58.945 59.645 -58.775 ;
      RECT 59.555 -57.74 59.645 -56.732 ;
      RECT 59.505 -57.505 59.645 -57.335 ;
      RECT 59.555 -56.318 59.645 -55.31 ;
      RECT 59.505 -55.715 59.645 -55.545 ;
      RECT 59.555 -54.51 59.645 -53.502 ;
      RECT 59.505 -54.275 59.645 -54.105 ;
      RECT 59.555 -53.088 59.645 -52.08 ;
      RECT 59.505 -52.485 59.645 -52.315 ;
      RECT 59.555 -51.28 59.645 -50.272 ;
      RECT 59.505 -51.045 59.645 -50.875 ;
      RECT 59.555 -49.858 59.645 -48.85 ;
      RECT 59.505 -49.255 59.645 -49.085 ;
      RECT 59.555 -48.05 59.645 -47.042 ;
      RECT 59.505 -47.815 59.645 -47.645 ;
      RECT 59.555 -46.628 59.645 -45.62 ;
      RECT 59.505 -46.025 59.645 -45.855 ;
      RECT 59.555 -44.82 59.645 -43.812 ;
      RECT 59.505 -44.585 59.645 -44.415 ;
      RECT 59.555 -43.398 59.645 -42.39 ;
      RECT 59.505 -42.795 59.645 -42.625 ;
      RECT 59.555 -41.59 59.645 -40.582 ;
      RECT 59.505 -41.355 59.645 -41.185 ;
      RECT 59.555 -40.168 59.645 -39.16 ;
      RECT 59.505 -39.565 59.645 -39.395 ;
      RECT 59.555 -38.36 59.645 -37.352 ;
      RECT 59.505 -38.125 59.645 -37.955 ;
      RECT 59.555 -36.938 59.645 -35.93 ;
      RECT 59.505 -36.335 59.645 -36.165 ;
      RECT 59.555 -35.13 59.645 -34.122 ;
      RECT 59.505 -34.895 59.645 -34.725 ;
      RECT 59.555 -33.708 59.645 -32.7 ;
      RECT 59.505 -33.105 59.645 -32.935 ;
      RECT 59.555 -31.9 59.645 -30.892 ;
      RECT 59.505 -31.665 59.645 -31.495 ;
      RECT 59.555 -30.478 59.645 -29.47 ;
      RECT 59.505 -29.875 59.645 -29.705 ;
      RECT 59.555 -28.67 59.645 -27.662 ;
      RECT 59.505 -28.435 59.645 -28.265 ;
      RECT 59.555 -27.248 59.645 -26.24 ;
      RECT 59.505 -26.645 59.645 -26.475 ;
      RECT 59.555 -25.44 59.645 -24.432 ;
      RECT 59.505 -25.205 59.645 -25.035 ;
      RECT 59.555 -24.018 59.645 -23.01 ;
      RECT 59.505 -23.415 59.645 -23.245 ;
      RECT 59.555 -22.21 59.645 -21.202 ;
      RECT 59.505 -21.975 59.645 -21.805 ;
      RECT 59.555 -20.788 59.645 -19.78 ;
      RECT 59.505 -20.185 59.645 -20.015 ;
      RECT 59.555 -18.98 59.645 -17.972 ;
      RECT 59.505 -18.745 59.645 -18.575 ;
      RECT 59.555 -17.558 59.645 -16.55 ;
      RECT 59.505 -16.955 59.645 -16.785 ;
      RECT 59.555 -15.75 59.645 -14.742 ;
      RECT 59.505 -15.515 59.645 -15.345 ;
      RECT 59.555 -14.328 59.645 -13.32 ;
      RECT 59.505 -13.725 59.645 -13.555 ;
      RECT 59.555 -12.52 59.645 -11.512 ;
      RECT 59.505 -12.285 59.645 -12.115 ;
      RECT 59.555 -11.098 59.645 -10.09 ;
      RECT 59.505 -10.495 59.645 -10.325 ;
      RECT 59.555 -9.29 59.645 -8.282 ;
      RECT 59.505 -9.055 59.645 -8.885 ;
      RECT 59.555 -7.868 59.645 -6.86 ;
      RECT 59.505 -7.265 59.645 -7.095 ;
      RECT 59.555 -6.06 59.645 -5.052 ;
      RECT 59.505 -5.825 59.645 -5.655 ;
      RECT 59.555 -4.638 59.645 -3.63 ;
      RECT 59.505 -4.035 59.645 -3.865 ;
      RECT 59.555 -2.83 59.645 -1.822 ;
      RECT 59.505 -2.595 59.645 -2.425 ;
      RECT 59.555 -1.408 59.645 -0.4 ;
      RECT 59.505 -0.805 59.645 -0.635 ;
      RECT 59.555 0.4 59.645 1.408 ;
      RECT 59.505 0.635 59.645 0.805 ;
      RECT 59.43 -114.685 59.605 -114.515 ;
      RECT 59.505 -114.895 59.605 -114.515 ;
      RECT 58.545 -113.555 58.645 -113.09 ;
      RECT 58.91 -113.555 59.01 -113.1 ;
      RECT 58.545 -113.555 59.39 -113.385 ;
      RECT 59.155 -101.538 59.245 -100.531 ;
      RECT 59.155 -101.225 59.295 -101.055 ;
      RECT 59.155 -99.729 59.245 -98.722 ;
      RECT 59.155 -99.205 59.295 -99.035 ;
      RECT 59.155 -98.308 59.245 -97.301 ;
      RECT 59.155 -97.995 59.295 -97.825 ;
      RECT 59.155 -96.499 59.245 -95.492 ;
      RECT 59.155 -95.975 59.295 -95.805 ;
      RECT 59.155 -95.078 59.245 -94.071 ;
      RECT 59.155 -94.765 59.295 -94.595 ;
      RECT 59.155 -93.269 59.245 -92.262 ;
      RECT 59.155 -92.745 59.295 -92.575 ;
      RECT 59.155 -91.848 59.245 -90.841 ;
      RECT 59.155 -91.535 59.295 -91.365 ;
      RECT 59.155 -90.039 59.245 -89.032 ;
      RECT 59.155 -89.515 59.295 -89.345 ;
      RECT 59.155 -88.618 59.245 -87.611 ;
      RECT 59.155 -88.305 59.295 -88.135 ;
      RECT 59.155 -86.809 59.245 -85.802 ;
      RECT 59.155 -86.285 59.295 -86.115 ;
      RECT 59.155 -85.388 59.245 -84.381 ;
      RECT 59.155 -85.075 59.295 -84.905 ;
      RECT 59.155 -83.579 59.245 -82.572 ;
      RECT 59.155 -83.055 59.295 -82.885 ;
      RECT 59.155 -82.158 59.245 -81.151 ;
      RECT 59.155 -81.845 59.295 -81.675 ;
      RECT 59.155 -80.349 59.245 -79.342 ;
      RECT 59.155 -79.825 59.295 -79.655 ;
      RECT 59.155 -78.928 59.245 -77.921 ;
      RECT 59.155 -78.615 59.295 -78.445 ;
      RECT 59.155 -77.119 59.245 -76.112 ;
      RECT 59.155 -76.595 59.295 -76.425 ;
      RECT 59.155 -75.698 59.245 -74.691 ;
      RECT 59.155 -75.385 59.295 -75.215 ;
      RECT 59.155 -73.889 59.245 -72.882 ;
      RECT 59.155 -73.365 59.295 -73.195 ;
      RECT 59.155 -72.468 59.245 -71.461 ;
      RECT 59.155 -72.155 59.295 -71.985 ;
      RECT 59.155 -70.659 59.245 -69.652 ;
      RECT 59.155 -70.135 59.295 -69.965 ;
      RECT 59.155 -69.238 59.245 -68.231 ;
      RECT 59.155 -68.925 59.295 -68.755 ;
      RECT 59.155 -67.429 59.245 -66.422 ;
      RECT 59.155 -66.905 59.295 -66.735 ;
      RECT 59.155 -66.008 59.245 -65.001 ;
      RECT 59.155 -65.695 59.295 -65.525 ;
      RECT 59.155 -64.199 59.245 -63.192 ;
      RECT 59.155 -63.675 59.295 -63.505 ;
      RECT 59.155 -62.778 59.245 -61.771 ;
      RECT 59.155 -62.465 59.295 -62.295 ;
      RECT 59.155 -60.969 59.245 -59.962 ;
      RECT 59.155 -60.445 59.295 -60.275 ;
      RECT 59.155 -59.548 59.245 -58.541 ;
      RECT 59.155 -59.235 59.295 -59.065 ;
      RECT 59.155 -57.739 59.245 -56.732 ;
      RECT 59.155 -57.215 59.295 -57.045 ;
      RECT 59.155 -56.318 59.245 -55.311 ;
      RECT 59.155 -56.005 59.295 -55.835 ;
      RECT 59.155 -54.509 59.245 -53.502 ;
      RECT 59.155 -53.985 59.295 -53.815 ;
      RECT 59.155 -53.088 59.245 -52.081 ;
      RECT 59.155 -52.775 59.295 -52.605 ;
      RECT 59.155 -51.279 59.245 -50.272 ;
      RECT 59.155 -50.755 59.295 -50.585 ;
      RECT 59.155 -49.858 59.245 -48.851 ;
      RECT 59.155 -49.545 59.295 -49.375 ;
      RECT 59.155 -48.049 59.245 -47.042 ;
      RECT 59.155 -47.525 59.295 -47.355 ;
      RECT 59.155 -46.628 59.245 -45.621 ;
      RECT 59.155 -46.315 59.295 -46.145 ;
      RECT 59.155 -44.819 59.245 -43.812 ;
      RECT 59.155 -44.295 59.295 -44.125 ;
      RECT 59.155 -43.398 59.245 -42.391 ;
      RECT 59.155 -43.085 59.295 -42.915 ;
      RECT 59.155 -41.589 59.245 -40.582 ;
      RECT 59.155 -41.065 59.295 -40.895 ;
      RECT 59.155 -40.168 59.245 -39.161 ;
      RECT 59.155 -39.855 59.295 -39.685 ;
      RECT 59.155 -38.359 59.245 -37.352 ;
      RECT 59.155 -37.835 59.295 -37.665 ;
      RECT 59.155 -36.938 59.245 -35.931 ;
      RECT 59.155 -36.625 59.295 -36.455 ;
      RECT 59.155 -35.129 59.245 -34.122 ;
      RECT 59.155 -34.605 59.295 -34.435 ;
      RECT 59.155 -33.708 59.245 -32.701 ;
      RECT 59.155 -33.395 59.295 -33.225 ;
      RECT 59.155 -31.899 59.245 -30.892 ;
      RECT 59.155 -31.375 59.295 -31.205 ;
      RECT 59.155 -30.478 59.245 -29.471 ;
      RECT 59.155 -30.165 59.295 -29.995 ;
      RECT 59.155 -28.669 59.245 -27.662 ;
      RECT 59.155 -28.145 59.295 -27.975 ;
      RECT 59.155 -27.248 59.245 -26.241 ;
      RECT 59.155 -26.935 59.295 -26.765 ;
      RECT 59.155 -25.439 59.245 -24.432 ;
      RECT 59.155 -24.915 59.295 -24.745 ;
      RECT 59.155 -24.018 59.245 -23.011 ;
      RECT 59.155 -23.705 59.295 -23.535 ;
      RECT 59.155 -22.209 59.245 -21.202 ;
      RECT 59.155 -21.685 59.295 -21.515 ;
      RECT 59.155 -20.788 59.245 -19.781 ;
      RECT 59.155 -20.475 59.295 -20.305 ;
      RECT 59.155 -18.979 59.245 -17.972 ;
      RECT 59.155 -18.455 59.295 -18.285 ;
      RECT 59.155 -17.558 59.245 -16.551 ;
      RECT 59.155 -17.245 59.295 -17.075 ;
      RECT 59.155 -15.749 59.245 -14.742 ;
      RECT 59.155 -15.225 59.295 -15.055 ;
      RECT 59.155 -14.328 59.245 -13.321 ;
      RECT 59.155 -14.015 59.295 -13.845 ;
      RECT 59.155 -12.519 59.245 -11.512 ;
      RECT 59.155 -11.995 59.295 -11.825 ;
      RECT 59.155 -11.098 59.245 -10.091 ;
      RECT 59.155 -10.785 59.295 -10.615 ;
      RECT 59.155 -9.289 59.245 -8.282 ;
      RECT 59.155 -8.765 59.295 -8.595 ;
      RECT 59.155 -7.868 59.245 -6.861 ;
      RECT 59.155 -7.555 59.295 -7.385 ;
      RECT 59.155 -6.059 59.245 -5.052 ;
      RECT 59.155 -5.535 59.295 -5.365 ;
      RECT 59.155 -4.638 59.245 -3.631 ;
      RECT 59.155 -4.325 59.295 -4.155 ;
      RECT 59.155 -2.829 59.245 -1.822 ;
      RECT 59.155 -2.305 59.295 -2.135 ;
      RECT 59.155 -1.408 59.245 -0.401 ;
      RECT 59.155 -1.095 59.295 -0.925 ;
      RECT 59.155 0.401 59.245 1.408 ;
      RECT 59.155 0.925 59.295 1.095 ;
      RECT 58.84 -114.685 59.01 -114.515 ;
      RECT 58.91 -114.895 59.01 -114.515 ;
      RECT 58.355 -101.538 58.445 -100.53 ;
      RECT 58.305 -100.935 58.445 -100.765 ;
      RECT 58.355 -99.73 58.445 -98.722 ;
      RECT 58.305 -99.495 58.445 -99.325 ;
      RECT 58.355 -98.308 58.445 -97.3 ;
      RECT 58.305 -97.705 58.445 -97.535 ;
      RECT 58.355 -96.5 58.445 -95.492 ;
      RECT 58.305 -96.265 58.445 -96.095 ;
      RECT 58.355 -95.078 58.445 -94.07 ;
      RECT 58.305 -94.475 58.445 -94.305 ;
      RECT 58.355 -93.27 58.445 -92.262 ;
      RECT 58.305 -93.035 58.445 -92.865 ;
      RECT 58.355 -91.848 58.445 -90.84 ;
      RECT 58.305 -91.245 58.445 -91.075 ;
      RECT 58.355 -90.04 58.445 -89.032 ;
      RECT 58.305 -89.805 58.445 -89.635 ;
      RECT 58.355 -88.618 58.445 -87.61 ;
      RECT 58.305 -88.015 58.445 -87.845 ;
      RECT 58.355 -86.81 58.445 -85.802 ;
      RECT 58.305 -86.575 58.445 -86.405 ;
      RECT 58.355 -85.388 58.445 -84.38 ;
      RECT 58.305 -84.785 58.445 -84.615 ;
      RECT 58.355 -83.58 58.445 -82.572 ;
      RECT 58.305 -83.345 58.445 -83.175 ;
      RECT 58.355 -82.158 58.445 -81.15 ;
      RECT 58.305 -81.555 58.445 -81.385 ;
      RECT 58.355 -80.35 58.445 -79.342 ;
      RECT 58.305 -80.115 58.445 -79.945 ;
      RECT 58.355 -78.928 58.445 -77.92 ;
      RECT 58.305 -78.325 58.445 -78.155 ;
      RECT 58.355 -77.12 58.445 -76.112 ;
      RECT 58.305 -76.885 58.445 -76.715 ;
      RECT 58.355 -75.698 58.445 -74.69 ;
      RECT 58.305 -75.095 58.445 -74.925 ;
      RECT 58.355 -73.89 58.445 -72.882 ;
      RECT 58.305 -73.655 58.445 -73.485 ;
      RECT 58.355 -72.468 58.445 -71.46 ;
      RECT 58.305 -71.865 58.445 -71.695 ;
      RECT 58.355 -70.66 58.445 -69.652 ;
      RECT 58.305 -70.425 58.445 -70.255 ;
      RECT 58.355 -69.238 58.445 -68.23 ;
      RECT 58.305 -68.635 58.445 -68.465 ;
      RECT 58.355 -67.43 58.445 -66.422 ;
      RECT 58.305 -67.195 58.445 -67.025 ;
      RECT 58.355 -66.008 58.445 -65 ;
      RECT 58.305 -65.405 58.445 -65.235 ;
      RECT 58.355 -64.2 58.445 -63.192 ;
      RECT 58.305 -63.965 58.445 -63.795 ;
      RECT 58.355 -62.778 58.445 -61.77 ;
      RECT 58.305 -62.175 58.445 -62.005 ;
      RECT 58.355 -60.97 58.445 -59.962 ;
      RECT 58.305 -60.735 58.445 -60.565 ;
      RECT 58.355 -59.548 58.445 -58.54 ;
      RECT 58.305 -58.945 58.445 -58.775 ;
      RECT 58.355 -57.74 58.445 -56.732 ;
      RECT 58.305 -57.505 58.445 -57.335 ;
      RECT 58.355 -56.318 58.445 -55.31 ;
      RECT 58.305 -55.715 58.445 -55.545 ;
      RECT 58.355 -54.51 58.445 -53.502 ;
      RECT 58.305 -54.275 58.445 -54.105 ;
      RECT 58.355 -53.088 58.445 -52.08 ;
      RECT 58.305 -52.485 58.445 -52.315 ;
      RECT 58.355 -51.28 58.445 -50.272 ;
      RECT 58.305 -51.045 58.445 -50.875 ;
      RECT 58.355 -49.858 58.445 -48.85 ;
      RECT 58.305 -49.255 58.445 -49.085 ;
      RECT 58.355 -48.05 58.445 -47.042 ;
      RECT 58.305 -47.815 58.445 -47.645 ;
      RECT 58.355 -46.628 58.445 -45.62 ;
      RECT 58.305 -46.025 58.445 -45.855 ;
      RECT 58.355 -44.82 58.445 -43.812 ;
      RECT 58.305 -44.585 58.445 -44.415 ;
      RECT 58.355 -43.398 58.445 -42.39 ;
      RECT 58.305 -42.795 58.445 -42.625 ;
      RECT 58.355 -41.59 58.445 -40.582 ;
      RECT 58.305 -41.355 58.445 -41.185 ;
      RECT 58.355 -40.168 58.445 -39.16 ;
      RECT 58.305 -39.565 58.445 -39.395 ;
      RECT 58.355 -38.36 58.445 -37.352 ;
      RECT 58.305 -38.125 58.445 -37.955 ;
      RECT 58.355 -36.938 58.445 -35.93 ;
      RECT 58.305 -36.335 58.445 -36.165 ;
      RECT 58.355 -35.13 58.445 -34.122 ;
      RECT 58.305 -34.895 58.445 -34.725 ;
      RECT 58.355 -33.708 58.445 -32.7 ;
      RECT 58.305 -33.105 58.445 -32.935 ;
      RECT 58.355 -31.9 58.445 -30.892 ;
      RECT 58.305 -31.665 58.445 -31.495 ;
      RECT 58.355 -30.478 58.445 -29.47 ;
      RECT 58.305 -29.875 58.445 -29.705 ;
      RECT 58.355 -28.67 58.445 -27.662 ;
      RECT 58.305 -28.435 58.445 -28.265 ;
      RECT 58.355 -27.248 58.445 -26.24 ;
      RECT 58.305 -26.645 58.445 -26.475 ;
      RECT 58.355 -25.44 58.445 -24.432 ;
      RECT 58.305 -25.205 58.445 -25.035 ;
      RECT 58.355 -24.018 58.445 -23.01 ;
      RECT 58.305 -23.415 58.445 -23.245 ;
      RECT 58.355 -22.21 58.445 -21.202 ;
      RECT 58.305 -21.975 58.445 -21.805 ;
      RECT 58.355 -20.788 58.445 -19.78 ;
      RECT 58.305 -20.185 58.445 -20.015 ;
      RECT 58.355 -18.98 58.445 -17.972 ;
      RECT 58.305 -18.745 58.445 -18.575 ;
      RECT 58.355 -17.558 58.445 -16.55 ;
      RECT 58.305 -16.955 58.445 -16.785 ;
      RECT 58.355 -15.75 58.445 -14.742 ;
      RECT 58.305 -15.515 58.445 -15.345 ;
      RECT 58.355 -14.328 58.445 -13.32 ;
      RECT 58.305 -13.725 58.445 -13.555 ;
      RECT 58.355 -12.52 58.445 -11.512 ;
      RECT 58.305 -12.285 58.445 -12.115 ;
      RECT 58.355 -11.098 58.445 -10.09 ;
      RECT 58.305 -10.495 58.445 -10.325 ;
      RECT 58.355 -9.29 58.445 -8.282 ;
      RECT 58.305 -9.055 58.445 -8.885 ;
      RECT 58.355 -7.868 58.445 -6.86 ;
      RECT 58.305 -7.265 58.445 -7.095 ;
      RECT 58.355 -6.06 58.445 -5.052 ;
      RECT 58.305 -5.825 58.445 -5.655 ;
      RECT 58.355 -4.638 58.445 -3.63 ;
      RECT 58.305 -4.035 58.445 -3.865 ;
      RECT 58.355 -2.83 58.445 -1.822 ;
      RECT 58.305 -2.595 58.445 -2.425 ;
      RECT 58.355 -1.408 58.445 -0.4 ;
      RECT 58.305 -0.805 58.445 -0.635 ;
      RECT 58.355 0.4 58.445 1.408 ;
      RECT 58.305 0.635 58.445 0.805 ;
      RECT 57.955 -101.538 58.045 -100.531 ;
      RECT 57.955 -101.225 58.095 -101.055 ;
      RECT 57.955 -99.729 58.045 -98.722 ;
      RECT 57.955 -99.205 58.095 -99.035 ;
      RECT 57.955 -98.308 58.045 -97.301 ;
      RECT 57.955 -97.995 58.095 -97.825 ;
      RECT 57.955 -96.499 58.045 -95.492 ;
      RECT 57.955 -95.975 58.095 -95.805 ;
      RECT 57.955 -95.078 58.045 -94.071 ;
      RECT 57.955 -94.765 58.095 -94.595 ;
      RECT 57.955 -93.269 58.045 -92.262 ;
      RECT 57.955 -92.745 58.095 -92.575 ;
      RECT 57.955 -91.848 58.045 -90.841 ;
      RECT 57.955 -91.535 58.095 -91.365 ;
      RECT 57.955 -90.039 58.045 -89.032 ;
      RECT 57.955 -89.515 58.095 -89.345 ;
      RECT 57.955 -88.618 58.045 -87.611 ;
      RECT 57.955 -88.305 58.095 -88.135 ;
      RECT 57.955 -86.809 58.045 -85.802 ;
      RECT 57.955 -86.285 58.095 -86.115 ;
      RECT 57.955 -85.388 58.045 -84.381 ;
      RECT 57.955 -85.075 58.095 -84.905 ;
      RECT 57.955 -83.579 58.045 -82.572 ;
      RECT 57.955 -83.055 58.095 -82.885 ;
      RECT 57.955 -82.158 58.045 -81.151 ;
      RECT 57.955 -81.845 58.095 -81.675 ;
      RECT 57.955 -80.349 58.045 -79.342 ;
      RECT 57.955 -79.825 58.095 -79.655 ;
      RECT 57.955 -78.928 58.045 -77.921 ;
      RECT 57.955 -78.615 58.095 -78.445 ;
      RECT 57.955 -77.119 58.045 -76.112 ;
      RECT 57.955 -76.595 58.095 -76.425 ;
      RECT 57.955 -75.698 58.045 -74.691 ;
      RECT 57.955 -75.385 58.095 -75.215 ;
      RECT 57.955 -73.889 58.045 -72.882 ;
      RECT 57.955 -73.365 58.095 -73.195 ;
      RECT 57.955 -72.468 58.045 -71.461 ;
      RECT 57.955 -72.155 58.095 -71.985 ;
      RECT 57.955 -70.659 58.045 -69.652 ;
      RECT 57.955 -70.135 58.095 -69.965 ;
      RECT 57.955 -69.238 58.045 -68.231 ;
      RECT 57.955 -68.925 58.095 -68.755 ;
      RECT 57.955 -67.429 58.045 -66.422 ;
      RECT 57.955 -66.905 58.095 -66.735 ;
      RECT 57.955 -66.008 58.045 -65.001 ;
      RECT 57.955 -65.695 58.095 -65.525 ;
      RECT 57.955 -64.199 58.045 -63.192 ;
      RECT 57.955 -63.675 58.095 -63.505 ;
      RECT 57.955 -62.778 58.045 -61.771 ;
      RECT 57.955 -62.465 58.095 -62.295 ;
      RECT 57.955 -60.969 58.045 -59.962 ;
      RECT 57.955 -60.445 58.095 -60.275 ;
      RECT 57.955 -59.548 58.045 -58.541 ;
      RECT 57.955 -59.235 58.095 -59.065 ;
      RECT 57.955 -57.739 58.045 -56.732 ;
      RECT 57.955 -57.215 58.095 -57.045 ;
      RECT 57.955 -56.318 58.045 -55.311 ;
      RECT 57.955 -56.005 58.095 -55.835 ;
      RECT 57.955 -54.509 58.045 -53.502 ;
      RECT 57.955 -53.985 58.095 -53.815 ;
      RECT 57.955 -53.088 58.045 -52.081 ;
      RECT 57.955 -52.775 58.095 -52.605 ;
      RECT 57.955 -51.279 58.045 -50.272 ;
      RECT 57.955 -50.755 58.095 -50.585 ;
      RECT 57.955 -49.858 58.045 -48.851 ;
      RECT 57.955 -49.545 58.095 -49.375 ;
      RECT 57.955 -48.049 58.045 -47.042 ;
      RECT 57.955 -47.525 58.095 -47.355 ;
      RECT 57.955 -46.628 58.045 -45.621 ;
      RECT 57.955 -46.315 58.095 -46.145 ;
      RECT 57.955 -44.819 58.045 -43.812 ;
      RECT 57.955 -44.295 58.095 -44.125 ;
      RECT 57.955 -43.398 58.045 -42.391 ;
      RECT 57.955 -43.085 58.095 -42.915 ;
      RECT 57.955 -41.589 58.045 -40.582 ;
      RECT 57.955 -41.065 58.095 -40.895 ;
      RECT 57.955 -40.168 58.045 -39.161 ;
      RECT 57.955 -39.855 58.095 -39.685 ;
      RECT 57.955 -38.359 58.045 -37.352 ;
      RECT 57.955 -37.835 58.095 -37.665 ;
      RECT 57.955 -36.938 58.045 -35.931 ;
      RECT 57.955 -36.625 58.095 -36.455 ;
      RECT 57.955 -35.129 58.045 -34.122 ;
      RECT 57.955 -34.605 58.095 -34.435 ;
      RECT 57.955 -33.708 58.045 -32.701 ;
      RECT 57.955 -33.395 58.095 -33.225 ;
      RECT 57.955 -31.899 58.045 -30.892 ;
      RECT 57.955 -31.375 58.095 -31.205 ;
      RECT 57.955 -30.478 58.045 -29.471 ;
      RECT 57.955 -30.165 58.095 -29.995 ;
      RECT 57.955 -28.669 58.045 -27.662 ;
      RECT 57.955 -28.145 58.095 -27.975 ;
      RECT 57.955 -27.248 58.045 -26.241 ;
      RECT 57.955 -26.935 58.095 -26.765 ;
      RECT 57.955 -25.439 58.045 -24.432 ;
      RECT 57.955 -24.915 58.095 -24.745 ;
      RECT 57.955 -24.018 58.045 -23.011 ;
      RECT 57.955 -23.705 58.095 -23.535 ;
      RECT 57.955 -22.209 58.045 -21.202 ;
      RECT 57.955 -21.685 58.095 -21.515 ;
      RECT 57.955 -20.788 58.045 -19.781 ;
      RECT 57.955 -20.475 58.095 -20.305 ;
      RECT 57.955 -18.979 58.045 -17.972 ;
      RECT 57.955 -18.455 58.095 -18.285 ;
      RECT 57.955 -17.558 58.045 -16.551 ;
      RECT 57.955 -17.245 58.095 -17.075 ;
      RECT 57.955 -15.749 58.045 -14.742 ;
      RECT 57.955 -15.225 58.095 -15.055 ;
      RECT 57.955 -14.328 58.045 -13.321 ;
      RECT 57.955 -14.015 58.095 -13.845 ;
      RECT 57.955 -12.519 58.045 -11.512 ;
      RECT 57.955 -11.995 58.095 -11.825 ;
      RECT 57.955 -11.098 58.045 -10.091 ;
      RECT 57.955 -10.785 58.095 -10.615 ;
      RECT 57.955 -9.289 58.045 -8.282 ;
      RECT 57.955 -8.765 58.095 -8.595 ;
      RECT 57.955 -7.868 58.045 -6.861 ;
      RECT 57.955 -7.555 58.095 -7.385 ;
      RECT 57.955 -6.059 58.045 -5.052 ;
      RECT 57.955 -5.535 58.095 -5.365 ;
      RECT 57.955 -4.638 58.045 -3.631 ;
      RECT 57.955 -4.325 58.095 -4.155 ;
      RECT 57.955 -2.829 58.045 -1.822 ;
      RECT 57.955 -2.305 58.095 -2.135 ;
      RECT 57.955 -1.408 58.045 -0.401 ;
      RECT 57.955 -1.095 58.095 -0.925 ;
      RECT 57.955 0.401 58.045 1.408 ;
      RECT 57.955 0.925 58.095 1.095 ;
      RECT 53.785 -108.935 57.565 -108.815 ;
      RECT 55.105 -109.475 55.205 -108.815 ;
      RECT 54.545 -109.475 54.645 -108.815 ;
      RECT 53.985 -109.475 54.085 -108.815 ;
      RECT 57.155 -101.538 57.245 -100.53 ;
      RECT 57.105 -100.935 57.245 -100.765 ;
      RECT 57.155 -99.73 57.245 -98.722 ;
      RECT 57.105 -99.495 57.245 -99.325 ;
      RECT 57.155 -98.308 57.245 -97.3 ;
      RECT 57.105 -97.705 57.245 -97.535 ;
      RECT 57.155 -96.5 57.245 -95.492 ;
      RECT 57.105 -96.265 57.245 -96.095 ;
      RECT 57.155 -95.078 57.245 -94.07 ;
      RECT 57.105 -94.475 57.245 -94.305 ;
      RECT 57.155 -93.27 57.245 -92.262 ;
      RECT 57.105 -93.035 57.245 -92.865 ;
      RECT 57.155 -91.848 57.245 -90.84 ;
      RECT 57.105 -91.245 57.245 -91.075 ;
      RECT 57.155 -90.04 57.245 -89.032 ;
      RECT 57.105 -89.805 57.245 -89.635 ;
      RECT 57.155 -88.618 57.245 -87.61 ;
      RECT 57.105 -88.015 57.245 -87.845 ;
      RECT 57.155 -86.81 57.245 -85.802 ;
      RECT 57.105 -86.575 57.245 -86.405 ;
      RECT 57.155 -85.388 57.245 -84.38 ;
      RECT 57.105 -84.785 57.245 -84.615 ;
      RECT 57.155 -83.58 57.245 -82.572 ;
      RECT 57.105 -83.345 57.245 -83.175 ;
      RECT 57.155 -82.158 57.245 -81.15 ;
      RECT 57.105 -81.555 57.245 -81.385 ;
      RECT 57.155 -80.35 57.245 -79.342 ;
      RECT 57.105 -80.115 57.245 -79.945 ;
      RECT 57.155 -78.928 57.245 -77.92 ;
      RECT 57.105 -78.325 57.245 -78.155 ;
      RECT 57.155 -77.12 57.245 -76.112 ;
      RECT 57.105 -76.885 57.245 -76.715 ;
      RECT 57.155 -75.698 57.245 -74.69 ;
      RECT 57.105 -75.095 57.245 -74.925 ;
      RECT 57.155 -73.89 57.245 -72.882 ;
      RECT 57.105 -73.655 57.245 -73.485 ;
      RECT 57.155 -72.468 57.245 -71.46 ;
      RECT 57.105 -71.865 57.245 -71.695 ;
      RECT 57.155 -70.66 57.245 -69.652 ;
      RECT 57.105 -70.425 57.245 -70.255 ;
      RECT 57.155 -69.238 57.245 -68.23 ;
      RECT 57.105 -68.635 57.245 -68.465 ;
      RECT 57.155 -67.43 57.245 -66.422 ;
      RECT 57.105 -67.195 57.245 -67.025 ;
      RECT 57.155 -66.008 57.245 -65 ;
      RECT 57.105 -65.405 57.245 -65.235 ;
      RECT 57.155 -64.2 57.245 -63.192 ;
      RECT 57.105 -63.965 57.245 -63.795 ;
      RECT 57.155 -62.778 57.245 -61.77 ;
      RECT 57.105 -62.175 57.245 -62.005 ;
      RECT 57.155 -60.97 57.245 -59.962 ;
      RECT 57.105 -60.735 57.245 -60.565 ;
      RECT 57.155 -59.548 57.245 -58.54 ;
      RECT 57.105 -58.945 57.245 -58.775 ;
      RECT 57.155 -57.74 57.245 -56.732 ;
      RECT 57.105 -57.505 57.245 -57.335 ;
      RECT 57.155 -56.318 57.245 -55.31 ;
      RECT 57.105 -55.715 57.245 -55.545 ;
      RECT 57.155 -54.51 57.245 -53.502 ;
      RECT 57.105 -54.275 57.245 -54.105 ;
      RECT 57.155 -53.088 57.245 -52.08 ;
      RECT 57.105 -52.485 57.245 -52.315 ;
      RECT 57.155 -51.28 57.245 -50.272 ;
      RECT 57.105 -51.045 57.245 -50.875 ;
      RECT 57.155 -49.858 57.245 -48.85 ;
      RECT 57.105 -49.255 57.245 -49.085 ;
      RECT 57.155 -48.05 57.245 -47.042 ;
      RECT 57.105 -47.815 57.245 -47.645 ;
      RECT 57.155 -46.628 57.245 -45.62 ;
      RECT 57.105 -46.025 57.245 -45.855 ;
      RECT 57.155 -44.82 57.245 -43.812 ;
      RECT 57.105 -44.585 57.245 -44.415 ;
      RECT 57.155 -43.398 57.245 -42.39 ;
      RECT 57.105 -42.795 57.245 -42.625 ;
      RECT 57.155 -41.59 57.245 -40.582 ;
      RECT 57.105 -41.355 57.245 -41.185 ;
      RECT 57.155 -40.168 57.245 -39.16 ;
      RECT 57.105 -39.565 57.245 -39.395 ;
      RECT 57.155 -38.36 57.245 -37.352 ;
      RECT 57.105 -38.125 57.245 -37.955 ;
      RECT 57.155 -36.938 57.245 -35.93 ;
      RECT 57.105 -36.335 57.245 -36.165 ;
      RECT 57.155 -35.13 57.245 -34.122 ;
      RECT 57.105 -34.895 57.245 -34.725 ;
      RECT 57.155 -33.708 57.245 -32.7 ;
      RECT 57.105 -33.105 57.245 -32.935 ;
      RECT 57.155 -31.9 57.245 -30.892 ;
      RECT 57.105 -31.665 57.245 -31.495 ;
      RECT 57.155 -30.478 57.245 -29.47 ;
      RECT 57.105 -29.875 57.245 -29.705 ;
      RECT 57.155 -28.67 57.245 -27.662 ;
      RECT 57.105 -28.435 57.245 -28.265 ;
      RECT 57.155 -27.248 57.245 -26.24 ;
      RECT 57.105 -26.645 57.245 -26.475 ;
      RECT 57.155 -25.44 57.245 -24.432 ;
      RECT 57.105 -25.205 57.245 -25.035 ;
      RECT 57.155 -24.018 57.245 -23.01 ;
      RECT 57.105 -23.415 57.245 -23.245 ;
      RECT 57.155 -22.21 57.245 -21.202 ;
      RECT 57.105 -21.975 57.245 -21.805 ;
      RECT 57.155 -20.788 57.245 -19.78 ;
      RECT 57.105 -20.185 57.245 -20.015 ;
      RECT 57.155 -18.98 57.245 -17.972 ;
      RECT 57.105 -18.745 57.245 -18.575 ;
      RECT 57.155 -17.558 57.245 -16.55 ;
      RECT 57.105 -16.955 57.245 -16.785 ;
      RECT 57.155 -15.75 57.245 -14.742 ;
      RECT 57.105 -15.515 57.245 -15.345 ;
      RECT 57.155 -14.328 57.245 -13.32 ;
      RECT 57.105 -13.725 57.245 -13.555 ;
      RECT 57.155 -12.52 57.245 -11.512 ;
      RECT 57.105 -12.285 57.245 -12.115 ;
      RECT 57.155 -11.098 57.245 -10.09 ;
      RECT 57.105 -10.495 57.245 -10.325 ;
      RECT 57.155 -9.29 57.245 -8.282 ;
      RECT 57.105 -9.055 57.245 -8.885 ;
      RECT 57.155 -7.868 57.245 -6.86 ;
      RECT 57.105 -7.265 57.245 -7.095 ;
      RECT 57.155 -6.06 57.245 -5.052 ;
      RECT 57.105 -5.825 57.245 -5.655 ;
      RECT 57.155 -4.638 57.245 -3.63 ;
      RECT 57.105 -4.035 57.245 -3.865 ;
      RECT 57.155 -2.83 57.245 -1.822 ;
      RECT 57.105 -2.595 57.245 -2.425 ;
      RECT 57.155 -1.408 57.245 -0.4 ;
      RECT 57.105 -0.805 57.245 -0.635 ;
      RECT 57.155 0.4 57.245 1.408 ;
      RECT 57.105 0.635 57.245 0.805 ;
      RECT 55.725 -111.685 57.205 -111.585 ;
      RECT 55.725 -112.195 55.825 -111.585 ;
      RECT 55.945 -109.15 57.205 -109.05 ;
      RECT 57.105 -109.475 57.205 -109.05 ;
      RECT 56.545 -109.475 56.645 -109.05 ;
      RECT 55.985 -109.475 56.085 -109.05 ;
      RECT 56.755 -101.538 56.845 -100.531 ;
      RECT 56.755 -101.225 56.895 -101.055 ;
      RECT 56.755 -99.729 56.845 -98.722 ;
      RECT 56.755 -99.205 56.895 -99.035 ;
      RECT 56.755 -98.308 56.845 -97.301 ;
      RECT 56.755 -97.995 56.895 -97.825 ;
      RECT 56.755 -96.499 56.845 -95.492 ;
      RECT 56.755 -95.975 56.895 -95.805 ;
      RECT 56.755 -95.078 56.845 -94.071 ;
      RECT 56.755 -94.765 56.895 -94.595 ;
      RECT 56.755 -93.269 56.845 -92.262 ;
      RECT 56.755 -92.745 56.895 -92.575 ;
      RECT 56.755 -91.848 56.845 -90.841 ;
      RECT 56.755 -91.535 56.895 -91.365 ;
      RECT 56.755 -90.039 56.845 -89.032 ;
      RECT 56.755 -89.515 56.895 -89.345 ;
      RECT 56.755 -88.618 56.845 -87.611 ;
      RECT 56.755 -88.305 56.895 -88.135 ;
      RECT 56.755 -86.809 56.845 -85.802 ;
      RECT 56.755 -86.285 56.895 -86.115 ;
      RECT 56.755 -85.388 56.845 -84.381 ;
      RECT 56.755 -85.075 56.895 -84.905 ;
      RECT 56.755 -83.579 56.845 -82.572 ;
      RECT 56.755 -83.055 56.895 -82.885 ;
      RECT 56.755 -82.158 56.845 -81.151 ;
      RECT 56.755 -81.845 56.895 -81.675 ;
      RECT 56.755 -80.349 56.845 -79.342 ;
      RECT 56.755 -79.825 56.895 -79.655 ;
      RECT 56.755 -78.928 56.845 -77.921 ;
      RECT 56.755 -78.615 56.895 -78.445 ;
      RECT 56.755 -77.119 56.845 -76.112 ;
      RECT 56.755 -76.595 56.895 -76.425 ;
      RECT 56.755 -75.698 56.845 -74.691 ;
      RECT 56.755 -75.385 56.895 -75.215 ;
      RECT 56.755 -73.889 56.845 -72.882 ;
      RECT 56.755 -73.365 56.895 -73.195 ;
      RECT 56.755 -72.468 56.845 -71.461 ;
      RECT 56.755 -72.155 56.895 -71.985 ;
      RECT 56.755 -70.659 56.845 -69.652 ;
      RECT 56.755 -70.135 56.895 -69.965 ;
      RECT 56.755 -69.238 56.845 -68.231 ;
      RECT 56.755 -68.925 56.895 -68.755 ;
      RECT 56.755 -67.429 56.845 -66.422 ;
      RECT 56.755 -66.905 56.895 -66.735 ;
      RECT 56.755 -66.008 56.845 -65.001 ;
      RECT 56.755 -65.695 56.895 -65.525 ;
      RECT 56.755 -64.199 56.845 -63.192 ;
      RECT 56.755 -63.675 56.895 -63.505 ;
      RECT 56.755 -62.778 56.845 -61.771 ;
      RECT 56.755 -62.465 56.895 -62.295 ;
      RECT 56.755 -60.969 56.845 -59.962 ;
      RECT 56.755 -60.445 56.895 -60.275 ;
      RECT 56.755 -59.548 56.845 -58.541 ;
      RECT 56.755 -59.235 56.895 -59.065 ;
      RECT 56.755 -57.739 56.845 -56.732 ;
      RECT 56.755 -57.215 56.895 -57.045 ;
      RECT 56.755 -56.318 56.845 -55.311 ;
      RECT 56.755 -56.005 56.895 -55.835 ;
      RECT 56.755 -54.509 56.845 -53.502 ;
      RECT 56.755 -53.985 56.895 -53.815 ;
      RECT 56.755 -53.088 56.845 -52.081 ;
      RECT 56.755 -52.775 56.895 -52.605 ;
      RECT 56.755 -51.279 56.845 -50.272 ;
      RECT 56.755 -50.755 56.895 -50.585 ;
      RECT 56.755 -49.858 56.845 -48.851 ;
      RECT 56.755 -49.545 56.895 -49.375 ;
      RECT 56.755 -48.049 56.845 -47.042 ;
      RECT 56.755 -47.525 56.895 -47.355 ;
      RECT 56.755 -46.628 56.845 -45.621 ;
      RECT 56.755 -46.315 56.895 -46.145 ;
      RECT 56.755 -44.819 56.845 -43.812 ;
      RECT 56.755 -44.295 56.895 -44.125 ;
      RECT 56.755 -43.398 56.845 -42.391 ;
      RECT 56.755 -43.085 56.895 -42.915 ;
      RECT 56.755 -41.589 56.845 -40.582 ;
      RECT 56.755 -41.065 56.895 -40.895 ;
      RECT 56.755 -40.168 56.845 -39.161 ;
      RECT 56.755 -39.855 56.895 -39.685 ;
      RECT 56.755 -38.359 56.845 -37.352 ;
      RECT 56.755 -37.835 56.895 -37.665 ;
      RECT 56.755 -36.938 56.845 -35.931 ;
      RECT 56.755 -36.625 56.895 -36.455 ;
      RECT 56.755 -35.129 56.845 -34.122 ;
      RECT 56.755 -34.605 56.895 -34.435 ;
      RECT 56.755 -33.708 56.845 -32.701 ;
      RECT 56.755 -33.395 56.895 -33.225 ;
      RECT 56.755 -31.899 56.845 -30.892 ;
      RECT 56.755 -31.375 56.895 -31.205 ;
      RECT 56.755 -30.478 56.845 -29.471 ;
      RECT 56.755 -30.165 56.895 -29.995 ;
      RECT 56.755 -28.669 56.845 -27.662 ;
      RECT 56.755 -28.145 56.895 -27.975 ;
      RECT 56.755 -27.248 56.845 -26.241 ;
      RECT 56.755 -26.935 56.895 -26.765 ;
      RECT 56.755 -25.439 56.845 -24.432 ;
      RECT 56.755 -24.915 56.895 -24.745 ;
      RECT 56.755 -24.018 56.845 -23.011 ;
      RECT 56.755 -23.705 56.895 -23.535 ;
      RECT 56.755 -22.209 56.845 -21.202 ;
      RECT 56.755 -21.685 56.895 -21.515 ;
      RECT 56.755 -20.788 56.845 -19.781 ;
      RECT 56.755 -20.475 56.895 -20.305 ;
      RECT 56.755 -18.979 56.845 -17.972 ;
      RECT 56.755 -18.455 56.895 -18.285 ;
      RECT 56.755 -17.558 56.845 -16.551 ;
      RECT 56.755 -17.245 56.895 -17.075 ;
      RECT 56.755 -15.749 56.845 -14.742 ;
      RECT 56.755 -15.225 56.895 -15.055 ;
      RECT 56.755 -14.328 56.845 -13.321 ;
      RECT 56.755 -14.015 56.895 -13.845 ;
      RECT 56.755 -12.519 56.845 -11.512 ;
      RECT 56.755 -11.995 56.895 -11.825 ;
      RECT 56.755 -11.098 56.845 -10.091 ;
      RECT 56.755 -10.785 56.895 -10.615 ;
      RECT 56.755 -9.289 56.845 -8.282 ;
      RECT 56.755 -8.765 56.895 -8.595 ;
      RECT 56.755 -7.868 56.845 -6.861 ;
      RECT 56.755 -7.555 56.895 -7.385 ;
      RECT 56.755 -6.059 56.845 -5.052 ;
      RECT 56.755 -5.535 56.895 -5.365 ;
      RECT 56.755 -4.638 56.845 -3.631 ;
      RECT 56.755 -4.325 56.895 -4.155 ;
      RECT 56.755 -2.829 56.845 -1.822 ;
      RECT 56.755 -2.305 56.895 -2.135 ;
      RECT 56.755 -1.408 56.845 -0.401 ;
      RECT 56.755 -1.095 56.895 -0.925 ;
      RECT 56.755 0.401 56.845 1.408 ;
      RECT 56.755 0.925 56.895 1.095 ;
      RECT 56.085 -111.495 56.255 -111.385 ;
      RECT 52.935 -111.495 56.255 -111.395 ;
      RECT 55.955 -101.538 56.045 -100.53 ;
      RECT 55.905 -100.935 56.045 -100.765 ;
      RECT 55.955 -99.73 56.045 -98.722 ;
      RECT 55.905 -99.495 56.045 -99.325 ;
      RECT 55.955 -98.308 56.045 -97.3 ;
      RECT 55.905 -97.705 56.045 -97.535 ;
      RECT 55.955 -96.5 56.045 -95.492 ;
      RECT 55.905 -96.265 56.045 -96.095 ;
      RECT 55.955 -95.078 56.045 -94.07 ;
      RECT 55.905 -94.475 56.045 -94.305 ;
      RECT 55.955 -93.27 56.045 -92.262 ;
      RECT 55.905 -93.035 56.045 -92.865 ;
      RECT 55.955 -91.848 56.045 -90.84 ;
      RECT 55.905 -91.245 56.045 -91.075 ;
      RECT 55.955 -90.04 56.045 -89.032 ;
      RECT 55.905 -89.805 56.045 -89.635 ;
      RECT 55.955 -88.618 56.045 -87.61 ;
      RECT 55.905 -88.015 56.045 -87.845 ;
      RECT 55.955 -86.81 56.045 -85.802 ;
      RECT 55.905 -86.575 56.045 -86.405 ;
      RECT 55.955 -85.388 56.045 -84.38 ;
      RECT 55.905 -84.785 56.045 -84.615 ;
      RECT 55.955 -83.58 56.045 -82.572 ;
      RECT 55.905 -83.345 56.045 -83.175 ;
      RECT 55.955 -82.158 56.045 -81.15 ;
      RECT 55.905 -81.555 56.045 -81.385 ;
      RECT 55.955 -80.35 56.045 -79.342 ;
      RECT 55.905 -80.115 56.045 -79.945 ;
      RECT 55.955 -78.928 56.045 -77.92 ;
      RECT 55.905 -78.325 56.045 -78.155 ;
      RECT 55.955 -77.12 56.045 -76.112 ;
      RECT 55.905 -76.885 56.045 -76.715 ;
      RECT 55.955 -75.698 56.045 -74.69 ;
      RECT 55.905 -75.095 56.045 -74.925 ;
      RECT 55.955 -73.89 56.045 -72.882 ;
      RECT 55.905 -73.655 56.045 -73.485 ;
      RECT 55.955 -72.468 56.045 -71.46 ;
      RECT 55.905 -71.865 56.045 -71.695 ;
      RECT 55.955 -70.66 56.045 -69.652 ;
      RECT 55.905 -70.425 56.045 -70.255 ;
      RECT 55.955 -69.238 56.045 -68.23 ;
      RECT 55.905 -68.635 56.045 -68.465 ;
      RECT 55.955 -67.43 56.045 -66.422 ;
      RECT 55.905 -67.195 56.045 -67.025 ;
      RECT 55.955 -66.008 56.045 -65 ;
      RECT 55.905 -65.405 56.045 -65.235 ;
      RECT 55.955 -64.2 56.045 -63.192 ;
      RECT 55.905 -63.965 56.045 -63.795 ;
      RECT 55.955 -62.778 56.045 -61.77 ;
      RECT 55.905 -62.175 56.045 -62.005 ;
      RECT 55.955 -60.97 56.045 -59.962 ;
      RECT 55.905 -60.735 56.045 -60.565 ;
      RECT 55.955 -59.548 56.045 -58.54 ;
      RECT 55.905 -58.945 56.045 -58.775 ;
      RECT 55.955 -57.74 56.045 -56.732 ;
      RECT 55.905 -57.505 56.045 -57.335 ;
      RECT 55.955 -56.318 56.045 -55.31 ;
      RECT 55.905 -55.715 56.045 -55.545 ;
      RECT 55.955 -54.51 56.045 -53.502 ;
      RECT 55.905 -54.275 56.045 -54.105 ;
      RECT 55.955 -53.088 56.045 -52.08 ;
      RECT 55.905 -52.485 56.045 -52.315 ;
      RECT 55.955 -51.28 56.045 -50.272 ;
      RECT 55.905 -51.045 56.045 -50.875 ;
      RECT 55.955 -49.858 56.045 -48.85 ;
      RECT 55.905 -49.255 56.045 -49.085 ;
      RECT 55.955 -48.05 56.045 -47.042 ;
      RECT 55.905 -47.815 56.045 -47.645 ;
      RECT 55.955 -46.628 56.045 -45.62 ;
      RECT 55.905 -46.025 56.045 -45.855 ;
      RECT 55.955 -44.82 56.045 -43.812 ;
      RECT 55.905 -44.585 56.045 -44.415 ;
      RECT 55.955 -43.398 56.045 -42.39 ;
      RECT 55.905 -42.795 56.045 -42.625 ;
      RECT 55.955 -41.59 56.045 -40.582 ;
      RECT 55.905 -41.355 56.045 -41.185 ;
      RECT 55.955 -40.168 56.045 -39.16 ;
      RECT 55.905 -39.565 56.045 -39.395 ;
      RECT 55.955 -38.36 56.045 -37.352 ;
      RECT 55.905 -38.125 56.045 -37.955 ;
      RECT 55.955 -36.938 56.045 -35.93 ;
      RECT 55.905 -36.335 56.045 -36.165 ;
      RECT 55.955 -35.13 56.045 -34.122 ;
      RECT 55.905 -34.895 56.045 -34.725 ;
      RECT 55.955 -33.708 56.045 -32.7 ;
      RECT 55.905 -33.105 56.045 -32.935 ;
      RECT 55.955 -31.9 56.045 -30.892 ;
      RECT 55.905 -31.665 56.045 -31.495 ;
      RECT 55.955 -30.478 56.045 -29.47 ;
      RECT 55.905 -29.875 56.045 -29.705 ;
      RECT 55.955 -28.67 56.045 -27.662 ;
      RECT 55.905 -28.435 56.045 -28.265 ;
      RECT 55.955 -27.248 56.045 -26.24 ;
      RECT 55.905 -26.645 56.045 -26.475 ;
      RECT 55.955 -25.44 56.045 -24.432 ;
      RECT 55.905 -25.205 56.045 -25.035 ;
      RECT 55.955 -24.018 56.045 -23.01 ;
      RECT 55.905 -23.415 56.045 -23.245 ;
      RECT 55.955 -22.21 56.045 -21.202 ;
      RECT 55.905 -21.975 56.045 -21.805 ;
      RECT 55.955 -20.788 56.045 -19.78 ;
      RECT 55.905 -20.185 56.045 -20.015 ;
      RECT 55.955 -18.98 56.045 -17.972 ;
      RECT 55.905 -18.745 56.045 -18.575 ;
      RECT 55.955 -17.558 56.045 -16.55 ;
      RECT 55.905 -16.955 56.045 -16.785 ;
      RECT 55.955 -15.75 56.045 -14.742 ;
      RECT 55.905 -15.515 56.045 -15.345 ;
      RECT 55.955 -14.328 56.045 -13.32 ;
      RECT 55.905 -13.725 56.045 -13.555 ;
      RECT 55.955 -12.52 56.045 -11.512 ;
      RECT 55.905 -12.285 56.045 -12.115 ;
      RECT 55.955 -11.098 56.045 -10.09 ;
      RECT 55.905 -10.495 56.045 -10.325 ;
      RECT 55.955 -9.29 56.045 -8.282 ;
      RECT 55.905 -9.055 56.045 -8.885 ;
      RECT 55.955 -7.868 56.045 -6.86 ;
      RECT 55.905 -7.265 56.045 -7.095 ;
      RECT 55.955 -6.06 56.045 -5.052 ;
      RECT 55.905 -5.825 56.045 -5.655 ;
      RECT 55.955 -4.638 56.045 -3.63 ;
      RECT 55.905 -4.035 56.045 -3.865 ;
      RECT 55.955 -2.83 56.045 -1.822 ;
      RECT 55.905 -2.595 56.045 -2.425 ;
      RECT 55.955 -1.408 56.045 -0.4 ;
      RECT 55.905 -0.805 56.045 -0.635 ;
      RECT 55.955 0.4 56.045 1.408 ;
      RECT 55.905 0.635 56.045 0.805 ;
      RECT 55.555 -101.538 55.645 -100.531 ;
      RECT 55.555 -101.225 55.695 -101.055 ;
      RECT 55.555 -99.729 55.645 -98.722 ;
      RECT 55.555 -99.205 55.695 -99.035 ;
      RECT 55.555 -98.308 55.645 -97.301 ;
      RECT 55.555 -97.995 55.695 -97.825 ;
      RECT 55.555 -96.499 55.645 -95.492 ;
      RECT 55.555 -95.975 55.695 -95.805 ;
      RECT 55.555 -95.078 55.645 -94.071 ;
      RECT 55.555 -94.765 55.695 -94.595 ;
      RECT 55.555 -93.269 55.645 -92.262 ;
      RECT 55.555 -92.745 55.695 -92.575 ;
      RECT 55.555 -91.848 55.645 -90.841 ;
      RECT 55.555 -91.535 55.695 -91.365 ;
      RECT 55.555 -90.039 55.645 -89.032 ;
      RECT 55.555 -89.515 55.695 -89.345 ;
      RECT 55.555 -88.618 55.645 -87.611 ;
      RECT 55.555 -88.305 55.695 -88.135 ;
      RECT 55.555 -86.809 55.645 -85.802 ;
      RECT 55.555 -86.285 55.695 -86.115 ;
      RECT 55.555 -85.388 55.645 -84.381 ;
      RECT 55.555 -85.075 55.695 -84.905 ;
      RECT 55.555 -83.579 55.645 -82.572 ;
      RECT 55.555 -83.055 55.695 -82.885 ;
      RECT 55.555 -82.158 55.645 -81.151 ;
      RECT 55.555 -81.845 55.695 -81.675 ;
      RECT 55.555 -80.349 55.645 -79.342 ;
      RECT 55.555 -79.825 55.695 -79.655 ;
      RECT 55.555 -78.928 55.645 -77.921 ;
      RECT 55.555 -78.615 55.695 -78.445 ;
      RECT 55.555 -77.119 55.645 -76.112 ;
      RECT 55.555 -76.595 55.695 -76.425 ;
      RECT 55.555 -75.698 55.645 -74.691 ;
      RECT 55.555 -75.385 55.695 -75.215 ;
      RECT 55.555 -73.889 55.645 -72.882 ;
      RECT 55.555 -73.365 55.695 -73.195 ;
      RECT 55.555 -72.468 55.645 -71.461 ;
      RECT 55.555 -72.155 55.695 -71.985 ;
      RECT 55.555 -70.659 55.645 -69.652 ;
      RECT 55.555 -70.135 55.695 -69.965 ;
      RECT 55.555 -69.238 55.645 -68.231 ;
      RECT 55.555 -68.925 55.695 -68.755 ;
      RECT 55.555 -67.429 55.645 -66.422 ;
      RECT 55.555 -66.905 55.695 -66.735 ;
      RECT 55.555 -66.008 55.645 -65.001 ;
      RECT 55.555 -65.695 55.695 -65.525 ;
      RECT 55.555 -64.199 55.645 -63.192 ;
      RECT 55.555 -63.675 55.695 -63.505 ;
      RECT 55.555 -62.778 55.645 -61.771 ;
      RECT 55.555 -62.465 55.695 -62.295 ;
      RECT 55.555 -60.969 55.645 -59.962 ;
      RECT 55.555 -60.445 55.695 -60.275 ;
      RECT 55.555 -59.548 55.645 -58.541 ;
      RECT 55.555 -59.235 55.695 -59.065 ;
      RECT 55.555 -57.739 55.645 -56.732 ;
      RECT 55.555 -57.215 55.695 -57.045 ;
      RECT 55.555 -56.318 55.645 -55.311 ;
      RECT 55.555 -56.005 55.695 -55.835 ;
      RECT 55.555 -54.509 55.645 -53.502 ;
      RECT 55.555 -53.985 55.695 -53.815 ;
      RECT 55.555 -53.088 55.645 -52.081 ;
      RECT 55.555 -52.775 55.695 -52.605 ;
      RECT 55.555 -51.279 55.645 -50.272 ;
      RECT 55.555 -50.755 55.695 -50.585 ;
      RECT 55.555 -49.858 55.645 -48.851 ;
      RECT 55.555 -49.545 55.695 -49.375 ;
      RECT 55.555 -48.049 55.645 -47.042 ;
      RECT 55.555 -47.525 55.695 -47.355 ;
      RECT 55.555 -46.628 55.645 -45.621 ;
      RECT 55.555 -46.315 55.695 -46.145 ;
      RECT 55.555 -44.819 55.645 -43.812 ;
      RECT 55.555 -44.295 55.695 -44.125 ;
      RECT 55.555 -43.398 55.645 -42.391 ;
      RECT 55.555 -43.085 55.695 -42.915 ;
      RECT 55.555 -41.589 55.645 -40.582 ;
      RECT 55.555 -41.065 55.695 -40.895 ;
      RECT 55.555 -40.168 55.645 -39.161 ;
      RECT 55.555 -39.855 55.695 -39.685 ;
      RECT 55.555 -38.359 55.645 -37.352 ;
      RECT 55.555 -37.835 55.695 -37.665 ;
      RECT 55.555 -36.938 55.645 -35.931 ;
      RECT 55.555 -36.625 55.695 -36.455 ;
      RECT 55.555 -35.129 55.645 -34.122 ;
      RECT 55.555 -34.605 55.695 -34.435 ;
      RECT 55.555 -33.708 55.645 -32.701 ;
      RECT 55.555 -33.395 55.695 -33.225 ;
      RECT 55.555 -31.899 55.645 -30.892 ;
      RECT 55.555 -31.375 55.695 -31.205 ;
      RECT 55.555 -30.478 55.645 -29.471 ;
      RECT 55.555 -30.165 55.695 -29.995 ;
      RECT 55.555 -28.669 55.645 -27.662 ;
      RECT 55.555 -28.145 55.695 -27.975 ;
      RECT 55.555 -27.248 55.645 -26.241 ;
      RECT 55.555 -26.935 55.695 -26.765 ;
      RECT 55.555 -25.439 55.645 -24.432 ;
      RECT 55.555 -24.915 55.695 -24.745 ;
      RECT 55.555 -24.018 55.645 -23.011 ;
      RECT 55.555 -23.705 55.695 -23.535 ;
      RECT 55.555 -22.209 55.645 -21.202 ;
      RECT 55.555 -21.685 55.695 -21.515 ;
      RECT 55.555 -20.788 55.645 -19.781 ;
      RECT 55.555 -20.475 55.695 -20.305 ;
      RECT 55.555 -18.979 55.645 -17.972 ;
      RECT 55.555 -18.455 55.695 -18.285 ;
      RECT 55.555 -17.558 55.645 -16.551 ;
      RECT 55.555 -17.245 55.695 -17.075 ;
      RECT 55.555 -15.749 55.645 -14.742 ;
      RECT 55.555 -15.225 55.695 -15.055 ;
      RECT 55.555 -14.328 55.645 -13.321 ;
      RECT 55.555 -14.015 55.695 -13.845 ;
      RECT 55.555 -12.519 55.645 -11.512 ;
      RECT 55.555 -11.995 55.695 -11.825 ;
      RECT 55.555 -11.098 55.645 -10.091 ;
      RECT 55.555 -10.785 55.695 -10.615 ;
      RECT 55.555 -9.289 55.645 -8.282 ;
      RECT 55.555 -8.765 55.695 -8.595 ;
      RECT 55.555 -7.868 55.645 -6.861 ;
      RECT 55.555 -7.555 55.695 -7.385 ;
      RECT 55.555 -6.059 55.645 -5.052 ;
      RECT 55.555 -5.535 55.695 -5.365 ;
      RECT 55.555 -4.638 55.645 -3.631 ;
      RECT 55.555 -4.325 55.695 -4.155 ;
      RECT 55.555 -2.829 55.645 -1.822 ;
      RECT 55.555 -2.305 55.695 -2.135 ;
      RECT 55.555 -1.408 55.645 -0.401 ;
      RECT 55.555 -1.095 55.695 -0.925 ;
      RECT 55.555 0.401 55.645 1.408 ;
      RECT 55.555 0.925 55.695 1.095 ;
      RECT 53.705 -111.685 55.185 -111.585 ;
      RECT 53.705 -112.055 53.805 -111.585 ;
      RECT 53.51 -114.395 55.085 -114.275 ;
      RECT 54.985 -114.895 55.085 -114.275 ;
      RECT 54.39 -114.895 54.49 -114.275 ;
      RECT 53.51 -114.85 53.61 -114.275 ;
      RECT 54.755 -101.538 54.845 -100.53 ;
      RECT 54.705 -100.935 54.845 -100.765 ;
      RECT 54.755 -99.73 54.845 -98.722 ;
      RECT 54.705 -99.495 54.845 -99.325 ;
      RECT 54.755 -98.308 54.845 -97.3 ;
      RECT 54.705 -97.705 54.845 -97.535 ;
      RECT 54.755 -96.5 54.845 -95.492 ;
      RECT 54.705 -96.265 54.845 -96.095 ;
      RECT 54.755 -95.078 54.845 -94.07 ;
      RECT 54.705 -94.475 54.845 -94.305 ;
      RECT 54.755 -93.27 54.845 -92.262 ;
      RECT 54.705 -93.035 54.845 -92.865 ;
      RECT 54.755 -91.848 54.845 -90.84 ;
      RECT 54.705 -91.245 54.845 -91.075 ;
      RECT 54.755 -90.04 54.845 -89.032 ;
      RECT 54.705 -89.805 54.845 -89.635 ;
      RECT 54.755 -88.618 54.845 -87.61 ;
      RECT 54.705 -88.015 54.845 -87.845 ;
      RECT 54.755 -86.81 54.845 -85.802 ;
      RECT 54.705 -86.575 54.845 -86.405 ;
      RECT 54.755 -85.388 54.845 -84.38 ;
      RECT 54.705 -84.785 54.845 -84.615 ;
      RECT 54.755 -83.58 54.845 -82.572 ;
      RECT 54.705 -83.345 54.845 -83.175 ;
      RECT 54.755 -82.158 54.845 -81.15 ;
      RECT 54.705 -81.555 54.845 -81.385 ;
      RECT 54.755 -80.35 54.845 -79.342 ;
      RECT 54.705 -80.115 54.845 -79.945 ;
      RECT 54.755 -78.928 54.845 -77.92 ;
      RECT 54.705 -78.325 54.845 -78.155 ;
      RECT 54.755 -77.12 54.845 -76.112 ;
      RECT 54.705 -76.885 54.845 -76.715 ;
      RECT 54.755 -75.698 54.845 -74.69 ;
      RECT 54.705 -75.095 54.845 -74.925 ;
      RECT 54.755 -73.89 54.845 -72.882 ;
      RECT 54.705 -73.655 54.845 -73.485 ;
      RECT 54.755 -72.468 54.845 -71.46 ;
      RECT 54.705 -71.865 54.845 -71.695 ;
      RECT 54.755 -70.66 54.845 -69.652 ;
      RECT 54.705 -70.425 54.845 -70.255 ;
      RECT 54.755 -69.238 54.845 -68.23 ;
      RECT 54.705 -68.635 54.845 -68.465 ;
      RECT 54.755 -67.43 54.845 -66.422 ;
      RECT 54.705 -67.195 54.845 -67.025 ;
      RECT 54.755 -66.008 54.845 -65 ;
      RECT 54.705 -65.405 54.845 -65.235 ;
      RECT 54.755 -64.2 54.845 -63.192 ;
      RECT 54.705 -63.965 54.845 -63.795 ;
      RECT 54.755 -62.778 54.845 -61.77 ;
      RECT 54.705 -62.175 54.845 -62.005 ;
      RECT 54.755 -60.97 54.845 -59.962 ;
      RECT 54.705 -60.735 54.845 -60.565 ;
      RECT 54.755 -59.548 54.845 -58.54 ;
      RECT 54.705 -58.945 54.845 -58.775 ;
      RECT 54.755 -57.74 54.845 -56.732 ;
      RECT 54.705 -57.505 54.845 -57.335 ;
      RECT 54.755 -56.318 54.845 -55.31 ;
      RECT 54.705 -55.715 54.845 -55.545 ;
      RECT 54.755 -54.51 54.845 -53.502 ;
      RECT 54.705 -54.275 54.845 -54.105 ;
      RECT 54.755 -53.088 54.845 -52.08 ;
      RECT 54.705 -52.485 54.845 -52.315 ;
      RECT 54.755 -51.28 54.845 -50.272 ;
      RECT 54.705 -51.045 54.845 -50.875 ;
      RECT 54.755 -49.858 54.845 -48.85 ;
      RECT 54.705 -49.255 54.845 -49.085 ;
      RECT 54.755 -48.05 54.845 -47.042 ;
      RECT 54.705 -47.815 54.845 -47.645 ;
      RECT 54.755 -46.628 54.845 -45.62 ;
      RECT 54.705 -46.025 54.845 -45.855 ;
      RECT 54.755 -44.82 54.845 -43.812 ;
      RECT 54.705 -44.585 54.845 -44.415 ;
      RECT 54.755 -43.398 54.845 -42.39 ;
      RECT 54.705 -42.795 54.845 -42.625 ;
      RECT 54.755 -41.59 54.845 -40.582 ;
      RECT 54.705 -41.355 54.845 -41.185 ;
      RECT 54.755 -40.168 54.845 -39.16 ;
      RECT 54.705 -39.565 54.845 -39.395 ;
      RECT 54.755 -38.36 54.845 -37.352 ;
      RECT 54.705 -38.125 54.845 -37.955 ;
      RECT 54.755 -36.938 54.845 -35.93 ;
      RECT 54.705 -36.335 54.845 -36.165 ;
      RECT 54.755 -35.13 54.845 -34.122 ;
      RECT 54.705 -34.895 54.845 -34.725 ;
      RECT 54.755 -33.708 54.845 -32.7 ;
      RECT 54.705 -33.105 54.845 -32.935 ;
      RECT 54.755 -31.9 54.845 -30.892 ;
      RECT 54.705 -31.665 54.845 -31.495 ;
      RECT 54.755 -30.478 54.845 -29.47 ;
      RECT 54.705 -29.875 54.845 -29.705 ;
      RECT 54.755 -28.67 54.845 -27.662 ;
      RECT 54.705 -28.435 54.845 -28.265 ;
      RECT 54.755 -27.248 54.845 -26.24 ;
      RECT 54.705 -26.645 54.845 -26.475 ;
      RECT 54.755 -25.44 54.845 -24.432 ;
      RECT 54.705 -25.205 54.845 -25.035 ;
      RECT 54.755 -24.018 54.845 -23.01 ;
      RECT 54.705 -23.415 54.845 -23.245 ;
      RECT 54.755 -22.21 54.845 -21.202 ;
      RECT 54.705 -21.975 54.845 -21.805 ;
      RECT 54.755 -20.788 54.845 -19.78 ;
      RECT 54.705 -20.185 54.845 -20.015 ;
      RECT 54.755 -18.98 54.845 -17.972 ;
      RECT 54.705 -18.745 54.845 -18.575 ;
      RECT 54.755 -17.558 54.845 -16.55 ;
      RECT 54.705 -16.955 54.845 -16.785 ;
      RECT 54.755 -15.75 54.845 -14.742 ;
      RECT 54.705 -15.515 54.845 -15.345 ;
      RECT 54.755 -14.328 54.845 -13.32 ;
      RECT 54.705 -13.725 54.845 -13.555 ;
      RECT 54.755 -12.52 54.845 -11.512 ;
      RECT 54.705 -12.285 54.845 -12.115 ;
      RECT 54.755 -11.098 54.845 -10.09 ;
      RECT 54.705 -10.495 54.845 -10.325 ;
      RECT 54.755 -9.29 54.845 -8.282 ;
      RECT 54.705 -9.055 54.845 -8.885 ;
      RECT 54.755 -7.868 54.845 -6.86 ;
      RECT 54.705 -7.265 54.845 -7.095 ;
      RECT 54.755 -6.06 54.845 -5.052 ;
      RECT 54.705 -5.825 54.845 -5.655 ;
      RECT 54.755 -4.638 54.845 -3.63 ;
      RECT 54.705 -4.035 54.845 -3.865 ;
      RECT 54.755 -2.83 54.845 -1.822 ;
      RECT 54.705 -2.595 54.845 -2.425 ;
      RECT 54.755 -1.408 54.845 -0.4 ;
      RECT 54.705 -0.805 54.845 -0.635 ;
      RECT 54.755 0.4 54.845 1.408 ;
      RECT 54.705 0.635 54.845 0.805 ;
      RECT 54.63 -114.685 54.805 -114.515 ;
      RECT 54.705 -114.895 54.805 -114.515 ;
      RECT 53.745 -113.555 53.845 -113.09 ;
      RECT 54.11 -113.555 54.21 -113.1 ;
      RECT 53.745 -113.555 54.59 -113.385 ;
      RECT 54.355 -101.538 54.445 -100.531 ;
      RECT 54.355 -101.225 54.495 -101.055 ;
      RECT 54.355 -99.729 54.445 -98.722 ;
      RECT 54.355 -99.205 54.495 -99.035 ;
      RECT 54.355 -98.308 54.445 -97.301 ;
      RECT 54.355 -97.995 54.495 -97.825 ;
      RECT 54.355 -96.499 54.445 -95.492 ;
      RECT 54.355 -95.975 54.495 -95.805 ;
      RECT 54.355 -95.078 54.445 -94.071 ;
      RECT 54.355 -94.765 54.495 -94.595 ;
      RECT 54.355 -93.269 54.445 -92.262 ;
      RECT 54.355 -92.745 54.495 -92.575 ;
      RECT 54.355 -91.848 54.445 -90.841 ;
      RECT 54.355 -91.535 54.495 -91.365 ;
      RECT 54.355 -90.039 54.445 -89.032 ;
      RECT 54.355 -89.515 54.495 -89.345 ;
      RECT 54.355 -88.618 54.445 -87.611 ;
      RECT 54.355 -88.305 54.495 -88.135 ;
      RECT 54.355 -86.809 54.445 -85.802 ;
      RECT 54.355 -86.285 54.495 -86.115 ;
      RECT 54.355 -85.388 54.445 -84.381 ;
      RECT 54.355 -85.075 54.495 -84.905 ;
      RECT 54.355 -83.579 54.445 -82.572 ;
      RECT 54.355 -83.055 54.495 -82.885 ;
      RECT 54.355 -82.158 54.445 -81.151 ;
      RECT 54.355 -81.845 54.495 -81.675 ;
      RECT 54.355 -80.349 54.445 -79.342 ;
      RECT 54.355 -79.825 54.495 -79.655 ;
      RECT 54.355 -78.928 54.445 -77.921 ;
      RECT 54.355 -78.615 54.495 -78.445 ;
      RECT 54.355 -77.119 54.445 -76.112 ;
      RECT 54.355 -76.595 54.495 -76.425 ;
      RECT 54.355 -75.698 54.445 -74.691 ;
      RECT 54.355 -75.385 54.495 -75.215 ;
      RECT 54.355 -73.889 54.445 -72.882 ;
      RECT 54.355 -73.365 54.495 -73.195 ;
      RECT 54.355 -72.468 54.445 -71.461 ;
      RECT 54.355 -72.155 54.495 -71.985 ;
      RECT 54.355 -70.659 54.445 -69.652 ;
      RECT 54.355 -70.135 54.495 -69.965 ;
      RECT 54.355 -69.238 54.445 -68.231 ;
      RECT 54.355 -68.925 54.495 -68.755 ;
      RECT 54.355 -67.429 54.445 -66.422 ;
      RECT 54.355 -66.905 54.495 -66.735 ;
      RECT 54.355 -66.008 54.445 -65.001 ;
      RECT 54.355 -65.695 54.495 -65.525 ;
      RECT 54.355 -64.199 54.445 -63.192 ;
      RECT 54.355 -63.675 54.495 -63.505 ;
      RECT 54.355 -62.778 54.445 -61.771 ;
      RECT 54.355 -62.465 54.495 -62.295 ;
      RECT 54.355 -60.969 54.445 -59.962 ;
      RECT 54.355 -60.445 54.495 -60.275 ;
      RECT 54.355 -59.548 54.445 -58.541 ;
      RECT 54.355 -59.235 54.495 -59.065 ;
      RECT 54.355 -57.739 54.445 -56.732 ;
      RECT 54.355 -57.215 54.495 -57.045 ;
      RECT 54.355 -56.318 54.445 -55.311 ;
      RECT 54.355 -56.005 54.495 -55.835 ;
      RECT 54.355 -54.509 54.445 -53.502 ;
      RECT 54.355 -53.985 54.495 -53.815 ;
      RECT 54.355 -53.088 54.445 -52.081 ;
      RECT 54.355 -52.775 54.495 -52.605 ;
      RECT 54.355 -51.279 54.445 -50.272 ;
      RECT 54.355 -50.755 54.495 -50.585 ;
      RECT 54.355 -49.858 54.445 -48.851 ;
      RECT 54.355 -49.545 54.495 -49.375 ;
      RECT 54.355 -48.049 54.445 -47.042 ;
      RECT 54.355 -47.525 54.495 -47.355 ;
      RECT 54.355 -46.628 54.445 -45.621 ;
      RECT 54.355 -46.315 54.495 -46.145 ;
      RECT 54.355 -44.819 54.445 -43.812 ;
      RECT 54.355 -44.295 54.495 -44.125 ;
      RECT 54.355 -43.398 54.445 -42.391 ;
      RECT 54.355 -43.085 54.495 -42.915 ;
      RECT 54.355 -41.589 54.445 -40.582 ;
      RECT 54.355 -41.065 54.495 -40.895 ;
      RECT 54.355 -40.168 54.445 -39.161 ;
      RECT 54.355 -39.855 54.495 -39.685 ;
      RECT 54.355 -38.359 54.445 -37.352 ;
      RECT 54.355 -37.835 54.495 -37.665 ;
      RECT 54.355 -36.938 54.445 -35.931 ;
      RECT 54.355 -36.625 54.495 -36.455 ;
      RECT 54.355 -35.129 54.445 -34.122 ;
      RECT 54.355 -34.605 54.495 -34.435 ;
      RECT 54.355 -33.708 54.445 -32.701 ;
      RECT 54.355 -33.395 54.495 -33.225 ;
      RECT 54.355 -31.899 54.445 -30.892 ;
      RECT 54.355 -31.375 54.495 -31.205 ;
      RECT 54.355 -30.478 54.445 -29.471 ;
      RECT 54.355 -30.165 54.495 -29.995 ;
      RECT 54.355 -28.669 54.445 -27.662 ;
      RECT 54.355 -28.145 54.495 -27.975 ;
      RECT 54.355 -27.248 54.445 -26.241 ;
      RECT 54.355 -26.935 54.495 -26.765 ;
      RECT 54.355 -25.439 54.445 -24.432 ;
      RECT 54.355 -24.915 54.495 -24.745 ;
      RECT 54.355 -24.018 54.445 -23.011 ;
      RECT 54.355 -23.705 54.495 -23.535 ;
      RECT 54.355 -22.209 54.445 -21.202 ;
      RECT 54.355 -21.685 54.495 -21.515 ;
      RECT 54.355 -20.788 54.445 -19.781 ;
      RECT 54.355 -20.475 54.495 -20.305 ;
      RECT 54.355 -18.979 54.445 -17.972 ;
      RECT 54.355 -18.455 54.495 -18.285 ;
      RECT 54.355 -17.558 54.445 -16.551 ;
      RECT 54.355 -17.245 54.495 -17.075 ;
      RECT 54.355 -15.749 54.445 -14.742 ;
      RECT 54.355 -15.225 54.495 -15.055 ;
      RECT 54.355 -14.328 54.445 -13.321 ;
      RECT 54.355 -14.015 54.495 -13.845 ;
      RECT 54.355 -12.519 54.445 -11.512 ;
      RECT 54.355 -11.995 54.495 -11.825 ;
      RECT 54.355 -11.098 54.445 -10.091 ;
      RECT 54.355 -10.785 54.495 -10.615 ;
      RECT 54.355 -9.289 54.445 -8.282 ;
      RECT 54.355 -8.765 54.495 -8.595 ;
      RECT 54.355 -7.868 54.445 -6.861 ;
      RECT 54.355 -7.555 54.495 -7.385 ;
      RECT 54.355 -6.059 54.445 -5.052 ;
      RECT 54.355 -5.535 54.495 -5.365 ;
      RECT 54.355 -4.638 54.445 -3.631 ;
      RECT 54.355 -4.325 54.495 -4.155 ;
      RECT 54.355 -2.829 54.445 -1.822 ;
      RECT 54.355 -2.305 54.495 -2.135 ;
      RECT 54.355 -1.408 54.445 -0.401 ;
      RECT 54.355 -1.095 54.495 -0.925 ;
      RECT 54.355 0.401 54.445 1.408 ;
      RECT 54.355 0.925 54.495 1.095 ;
      RECT 54.04 -114.685 54.21 -114.515 ;
      RECT 54.11 -114.895 54.21 -114.515 ;
      RECT 53.555 -101.538 53.645 -100.53 ;
      RECT 53.505 -100.935 53.645 -100.765 ;
      RECT 53.555 -99.73 53.645 -98.722 ;
      RECT 53.505 -99.495 53.645 -99.325 ;
      RECT 53.555 -98.308 53.645 -97.3 ;
      RECT 53.505 -97.705 53.645 -97.535 ;
      RECT 53.555 -96.5 53.645 -95.492 ;
      RECT 53.505 -96.265 53.645 -96.095 ;
      RECT 53.555 -95.078 53.645 -94.07 ;
      RECT 53.505 -94.475 53.645 -94.305 ;
      RECT 53.555 -93.27 53.645 -92.262 ;
      RECT 53.505 -93.035 53.645 -92.865 ;
      RECT 53.555 -91.848 53.645 -90.84 ;
      RECT 53.505 -91.245 53.645 -91.075 ;
      RECT 53.555 -90.04 53.645 -89.032 ;
      RECT 53.505 -89.805 53.645 -89.635 ;
      RECT 53.555 -88.618 53.645 -87.61 ;
      RECT 53.505 -88.015 53.645 -87.845 ;
      RECT 53.555 -86.81 53.645 -85.802 ;
      RECT 53.505 -86.575 53.645 -86.405 ;
      RECT 53.555 -85.388 53.645 -84.38 ;
      RECT 53.505 -84.785 53.645 -84.615 ;
      RECT 53.555 -83.58 53.645 -82.572 ;
      RECT 53.505 -83.345 53.645 -83.175 ;
      RECT 53.555 -82.158 53.645 -81.15 ;
      RECT 53.505 -81.555 53.645 -81.385 ;
      RECT 53.555 -80.35 53.645 -79.342 ;
      RECT 53.505 -80.115 53.645 -79.945 ;
      RECT 53.555 -78.928 53.645 -77.92 ;
      RECT 53.505 -78.325 53.645 -78.155 ;
      RECT 53.555 -77.12 53.645 -76.112 ;
      RECT 53.505 -76.885 53.645 -76.715 ;
      RECT 53.555 -75.698 53.645 -74.69 ;
      RECT 53.505 -75.095 53.645 -74.925 ;
      RECT 53.555 -73.89 53.645 -72.882 ;
      RECT 53.505 -73.655 53.645 -73.485 ;
      RECT 53.555 -72.468 53.645 -71.46 ;
      RECT 53.505 -71.865 53.645 -71.695 ;
      RECT 53.555 -70.66 53.645 -69.652 ;
      RECT 53.505 -70.425 53.645 -70.255 ;
      RECT 53.555 -69.238 53.645 -68.23 ;
      RECT 53.505 -68.635 53.645 -68.465 ;
      RECT 53.555 -67.43 53.645 -66.422 ;
      RECT 53.505 -67.195 53.645 -67.025 ;
      RECT 53.555 -66.008 53.645 -65 ;
      RECT 53.505 -65.405 53.645 -65.235 ;
      RECT 53.555 -64.2 53.645 -63.192 ;
      RECT 53.505 -63.965 53.645 -63.795 ;
      RECT 53.555 -62.778 53.645 -61.77 ;
      RECT 53.505 -62.175 53.645 -62.005 ;
      RECT 53.555 -60.97 53.645 -59.962 ;
      RECT 53.505 -60.735 53.645 -60.565 ;
      RECT 53.555 -59.548 53.645 -58.54 ;
      RECT 53.505 -58.945 53.645 -58.775 ;
      RECT 53.555 -57.74 53.645 -56.732 ;
      RECT 53.505 -57.505 53.645 -57.335 ;
      RECT 53.555 -56.318 53.645 -55.31 ;
      RECT 53.505 -55.715 53.645 -55.545 ;
      RECT 53.555 -54.51 53.645 -53.502 ;
      RECT 53.505 -54.275 53.645 -54.105 ;
      RECT 53.555 -53.088 53.645 -52.08 ;
      RECT 53.505 -52.485 53.645 -52.315 ;
      RECT 53.555 -51.28 53.645 -50.272 ;
      RECT 53.505 -51.045 53.645 -50.875 ;
      RECT 53.555 -49.858 53.645 -48.85 ;
      RECT 53.505 -49.255 53.645 -49.085 ;
      RECT 53.555 -48.05 53.645 -47.042 ;
      RECT 53.505 -47.815 53.645 -47.645 ;
      RECT 53.555 -46.628 53.645 -45.62 ;
      RECT 53.505 -46.025 53.645 -45.855 ;
      RECT 53.555 -44.82 53.645 -43.812 ;
      RECT 53.505 -44.585 53.645 -44.415 ;
      RECT 53.555 -43.398 53.645 -42.39 ;
      RECT 53.505 -42.795 53.645 -42.625 ;
      RECT 53.555 -41.59 53.645 -40.582 ;
      RECT 53.505 -41.355 53.645 -41.185 ;
      RECT 53.555 -40.168 53.645 -39.16 ;
      RECT 53.505 -39.565 53.645 -39.395 ;
      RECT 53.555 -38.36 53.645 -37.352 ;
      RECT 53.505 -38.125 53.645 -37.955 ;
      RECT 53.555 -36.938 53.645 -35.93 ;
      RECT 53.505 -36.335 53.645 -36.165 ;
      RECT 53.555 -35.13 53.645 -34.122 ;
      RECT 53.505 -34.895 53.645 -34.725 ;
      RECT 53.555 -33.708 53.645 -32.7 ;
      RECT 53.505 -33.105 53.645 -32.935 ;
      RECT 53.555 -31.9 53.645 -30.892 ;
      RECT 53.505 -31.665 53.645 -31.495 ;
      RECT 53.555 -30.478 53.645 -29.47 ;
      RECT 53.505 -29.875 53.645 -29.705 ;
      RECT 53.555 -28.67 53.645 -27.662 ;
      RECT 53.505 -28.435 53.645 -28.265 ;
      RECT 53.555 -27.248 53.645 -26.24 ;
      RECT 53.505 -26.645 53.645 -26.475 ;
      RECT 53.555 -25.44 53.645 -24.432 ;
      RECT 53.505 -25.205 53.645 -25.035 ;
      RECT 53.555 -24.018 53.645 -23.01 ;
      RECT 53.505 -23.415 53.645 -23.245 ;
      RECT 53.555 -22.21 53.645 -21.202 ;
      RECT 53.505 -21.975 53.645 -21.805 ;
      RECT 53.555 -20.788 53.645 -19.78 ;
      RECT 53.505 -20.185 53.645 -20.015 ;
      RECT 53.555 -18.98 53.645 -17.972 ;
      RECT 53.505 -18.745 53.645 -18.575 ;
      RECT 53.555 -17.558 53.645 -16.55 ;
      RECT 53.505 -16.955 53.645 -16.785 ;
      RECT 53.555 -15.75 53.645 -14.742 ;
      RECT 53.505 -15.515 53.645 -15.345 ;
      RECT 53.555 -14.328 53.645 -13.32 ;
      RECT 53.505 -13.725 53.645 -13.555 ;
      RECT 53.555 -12.52 53.645 -11.512 ;
      RECT 53.505 -12.285 53.645 -12.115 ;
      RECT 53.555 -11.098 53.645 -10.09 ;
      RECT 53.505 -10.495 53.645 -10.325 ;
      RECT 53.555 -9.29 53.645 -8.282 ;
      RECT 53.505 -9.055 53.645 -8.885 ;
      RECT 53.555 -7.868 53.645 -6.86 ;
      RECT 53.505 -7.265 53.645 -7.095 ;
      RECT 53.555 -6.06 53.645 -5.052 ;
      RECT 53.505 -5.825 53.645 -5.655 ;
      RECT 53.555 -4.638 53.645 -3.63 ;
      RECT 53.505 -4.035 53.645 -3.865 ;
      RECT 53.555 -2.83 53.645 -1.822 ;
      RECT 53.505 -2.595 53.645 -2.425 ;
      RECT 53.555 -1.408 53.645 -0.4 ;
      RECT 53.505 -0.805 53.645 -0.635 ;
      RECT 53.555 0.4 53.645 1.408 ;
      RECT 53.505 0.635 53.645 0.805 ;
      RECT 53.155 -101.538 53.245 -100.531 ;
      RECT 53.155 -101.225 53.295 -101.055 ;
      RECT 53.155 -99.729 53.245 -98.722 ;
      RECT 53.155 -99.205 53.295 -99.035 ;
      RECT 53.155 -98.308 53.245 -97.301 ;
      RECT 53.155 -97.995 53.295 -97.825 ;
      RECT 53.155 -96.499 53.245 -95.492 ;
      RECT 53.155 -95.975 53.295 -95.805 ;
      RECT 53.155 -95.078 53.245 -94.071 ;
      RECT 53.155 -94.765 53.295 -94.595 ;
      RECT 53.155 -93.269 53.245 -92.262 ;
      RECT 53.155 -92.745 53.295 -92.575 ;
      RECT 53.155 -91.848 53.245 -90.841 ;
      RECT 53.155 -91.535 53.295 -91.365 ;
      RECT 53.155 -90.039 53.245 -89.032 ;
      RECT 53.155 -89.515 53.295 -89.345 ;
      RECT 53.155 -88.618 53.245 -87.611 ;
      RECT 53.155 -88.305 53.295 -88.135 ;
      RECT 53.155 -86.809 53.245 -85.802 ;
      RECT 53.155 -86.285 53.295 -86.115 ;
      RECT 53.155 -85.388 53.245 -84.381 ;
      RECT 53.155 -85.075 53.295 -84.905 ;
      RECT 53.155 -83.579 53.245 -82.572 ;
      RECT 53.155 -83.055 53.295 -82.885 ;
      RECT 53.155 -82.158 53.245 -81.151 ;
      RECT 53.155 -81.845 53.295 -81.675 ;
      RECT 53.155 -80.349 53.245 -79.342 ;
      RECT 53.155 -79.825 53.295 -79.655 ;
      RECT 53.155 -78.928 53.245 -77.921 ;
      RECT 53.155 -78.615 53.295 -78.445 ;
      RECT 53.155 -77.119 53.245 -76.112 ;
      RECT 53.155 -76.595 53.295 -76.425 ;
      RECT 53.155 -75.698 53.245 -74.691 ;
      RECT 53.155 -75.385 53.295 -75.215 ;
      RECT 53.155 -73.889 53.245 -72.882 ;
      RECT 53.155 -73.365 53.295 -73.195 ;
      RECT 53.155 -72.468 53.245 -71.461 ;
      RECT 53.155 -72.155 53.295 -71.985 ;
      RECT 53.155 -70.659 53.245 -69.652 ;
      RECT 53.155 -70.135 53.295 -69.965 ;
      RECT 53.155 -69.238 53.245 -68.231 ;
      RECT 53.155 -68.925 53.295 -68.755 ;
      RECT 53.155 -67.429 53.245 -66.422 ;
      RECT 53.155 -66.905 53.295 -66.735 ;
      RECT 53.155 -66.008 53.245 -65.001 ;
      RECT 53.155 -65.695 53.295 -65.525 ;
      RECT 53.155 -64.199 53.245 -63.192 ;
      RECT 53.155 -63.675 53.295 -63.505 ;
      RECT 53.155 -62.778 53.245 -61.771 ;
      RECT 53.155 -62.465 53.295 -62.295 ;
      RECT 53.155 -60.969 53.245 -59.962 ;
      RECT 53.155 -60.445 53.295 -60.275 ;
      RECT 53.155 -59.548 53.245 -58.541 ;
      RECT 53.155 -59.235 53.295 -59.065 ;
      RECT 53.155 -57.739 53.245 -56.732 ;
      RECT 53.155 -57.215 53.295 -57.045 ;
      RECT 53.155 -56.318 53.245 -55.311 ;
      RECT 53.155 -56.005 53.295 -55.835 ;
      RECT 53.155 -54.509 53.245 -53.502 ;
      RECT 53.155 -53.985 53.295 -53.815 ;
      RECT 53.155 -53.088 53.245 -52.081 ;
      RECT 53.155 -52.775 53.295 -52.605 ;
      RECT 53.155 -51.279 53.245 -50.272 ;
      RECT 53.155 -50.755 53.295 -50.585 ;
      RECT 53.155 -49.858 53.245 -48.851 ;
      RECT 53.155 -49.545 53.295 -49.375 ;
      RECT 53.155 -48.049 53.245 -47.042 ;
      RECT 53.155 -47.525 53.295 -47.355 ;
      RECT 53.155 -46.628 53.245 -45.621 ;
      RECT 53.155 -46.315 53.295 -46.145 ;
      RECT 53.155 -44.819 53.245 -43.812 ;
      RECT 53.155 -44.295 53.295 -44.125 ;
      RECT 53.155 -43.398 53.245 -42.391 ;
      RECT 53.155 -43.085 53.295 -42.915 ;
      RECT 53.155 -41.589 53.245 -40.582 ;
      RECT 53.155 -41.065 53.295 -40.895 ;
      RECT 53.155 -40.168 53.245 -39.161 ;
      RECT 53.155 -39.855 53.295 -39.685 ;
      RECT 53.155 -38.359 53.245 -37.352 ;
      RECT 53.155 -37.835 53.295 -37.665 ;
      RECT 53.155 -36.938 53.245 -35.931 ;
      RECT 53.155 -36.625 53.295 -36.455 ;
      RECT 53.155 -35.129 53.245 -34.122 ;
      RECT 53.155 -34.605 53.295 -34.435 ;
      RECT 53.155 -33.708 53.245 -32.701 ;
      RECT 53.155 -33.395 53.295 -33.225 ;
      RECT 53.155 -31.899 53.245 -30.892 ;
      RECT 53.155 -31.375 53.295 -31.205 ;
      RECT 53.155 -30.478 53.245 -29.471 ;
      RECT 53.155 -30.165 53.295 -29.995 ;
      RECT 53.155 -28.669 53.245 -27.662 ;
      RECT 53.155 -28.145 53.295 -27.975 ;
      RECT 53.155 -27.248 53.245 -26.241 ;
      RECT 53.155 -26.935 53.295 -26.765 ;
      RECT 53.155 -25.439 53.245 -24.432 ;
      RECT 53.155 -24.915 53.295 -24.745 ;
      RECT 53.155 -24.018 53.245 -23.011 ;
      RECT 53.155 -23.705 53.295 -23.535 ;
      RECT 53.155 -22.209 53.245 -21.202 ;
      RECT 53.155 -21.685 53.295 -21.515 ;
      RECT 53.155 -20.788 53.245 -19.781 ;
      RECT 53.155 -20.475 53.295 -20.305 ;
      RECT 53.155 -18.979 53.245 -17.972 ;
      RECT 53.155 -18.455 53.295 -18.285 ;
      RECT 53.155 -17.558 53.245 -16.551 ;
      RECT 53.155 -17.245 53.295 -17.075 ;
      RECT 53.155 -15.749 53.245 -14.742 ;
      RECT 53.155 -15.225 53.295 -15.055 ;
      RECT 53.155 -14.328 53.245 -13.321 ;
      RECT 53.155 -14.015 53.295 -13.845 ;
      RECT 53.155 -12.519 53.245 -11.512 ;
      RECT 53.155 -11.995 53.295 -11.825 ;
      RECT 53.155 -11.098 53.245 -10.091 ;
      RECT 53.155 -10.785 53.295 -10.615 ;
      RECT 53.155 -9.289 53.245 -8.282 ;
      RECT 53.155 -8.765 53.295 -8.595 ;
      RECT 53.155 -7.868 53.245 -6.861 ;
      RECT 53.155 -7.555 53.295 -7.385 ;
      RECT 53.155 -6.059 53.245 -5.052 ;
      RECT 53.155 -5.535 53.295 -5.365 ;
      RECT 53.155 -4.638 53.245 -3.631 ;
      RECT 53.155 -4.325 53.295 -4.155 ;
      RECT 53.155 -2.829 53.245 -1.822 ;
      RECT 53.155 -2.305 53.295 -2.135 ;
      RECT 53.155 -1.408 53.245 -0.401 ;
      RECT 53.155 -1.095 53.295 -0.925 ;
      RECT 53.155 0.401 53.245 1.408 ;
      RECT 53.155 0.925 53.295 1.095 ;
      RECT 48.985 -108.935 52.765 -108.815 ;
      RECT 50.305 -109.475 50.405 -108.815 ;
      RECT 49.745 -109.475 49.845 -108.815 ;
      RECT 49.185 -109.475 49.285 -108.815 ;
      RECT 52.355 -101.538 52.445 -100.53 ;
      RECT 52.305 -100.935 52.445 -100.765 ;
      RECT 52.355 -99.73 52.445 -98.722 ;
      RECT 52.305 -99.495 52.445 -99.325 ;
      RECT 52.355 -98.308 52.445 -97.3 ;
      RECT 52.305 -97.705 52.445 -97.535 ;
      RECT 52.355 -96.5 52.445 -95.492 ;
      RECT 52.305 -96.265 52.445 -96.095 ;
      RECT 52.355 -95.078 52.445 -94.07 ;
      RECT 52.305 -94.475 52.445 -94.305 ;
      RECT 52.355 -93.27 52.445 -92.262 ;
      RECT 52.305 -93.035 52.445 -92.865 ;
      RECT 52.355 -91.848 52.445 -90.84 ;
      RECT 52.305 -91.245 52.445 -91.075 ;
      RECT 52.355 -90.04 52.445 -89.032 ;
      RECT 52.305 -89.805 52.445 -89.635 ;
      RECT 52.355 -88.618 52.445 -87.61 ;
      RECT 52.305 -88.015 52.445 -87.845 ;
      RECT 52.355 -86.81 52.445 -85.802 ;
      RECT 52.305 -86.575 52.445 -86.405 ;
      RECT 52.355 -85.388 52.445 -84.38 ;
      RECT 52.305 -84.785 52.445 -84.615 ;
      RECT 52.355 -83.58 52.445 -82.572 ;
      RECT 52.305 -83.345 52.445 -83.175 ;
      RECT 52.355 -82.158 52.445 -81.15 ;
      RECT 52.305 -81.555 52.445 -81.385 ;
      RECT 52.355 -80.35 52.445 -79.342 ;
      RECT 52.305 -80.115 52.445 -79.945 ;
      RECT 52.355 -78.928 52.445 -77.92 ;
      RECT 52.305 -78.325 52.445 -78.155 ;
      RECT 52.355 -77.12 52.445 -76.112 ;
      RECT 52.305 -76.885 52.445 -76.715 ;
      RECT 52.355 -75.698 52.445 -74.69 ;
      RECT 52.305 -75.095 52.445 -74.925 ;
      RECT 52.355 -73.89 52.445 -72.882 ;
      RECT 52.305 -73.655 52.445 -73.485 ;
      RECT 52.355 -72.468 52.445 -71.46 ;
      RECT 52.305 -71.865 52.445 -71.695 ;
      RECT 52.355 -70.66 52.445 -69.652 ;
      RECT 52.305 -70.425 52.445 -70.255 ;
      RECT 52.355 -69.238 52.445 -68.23 ;
      RECT 52.305 -68.635 52.445 -68.465 ;
      RECT 52.355 -67.43 52.445 -66.422 ;
      RECT 52.305 -67.195 52.445 -67.025 ;
      RECT 52.355 -66.008 52.445 -65 ;
      RECT 52.305 -65.405 52.445 -65.235 ;
      RECT 52.355 -64.2 52.445 -63.192 ;
      RECT 52.305 -63.965 52.445 -63.795 ;
      RECT 52.355 -62.778 52.445 -61.77 ;
      RECT 52.305 -62.175 52.445 -62.005 ;
      RECT 52.355 -60.97 52.445 -59.962 ;
      RECT 52.305 -60.735 52.445 -60.565 ;
      RECT 52.355 -59.548 52.445 -58.54 ;
      RECT 52.305 -58.945 52.445 -58.775 ;
      RECT 52.355 -57.74 52.445 -56.732 ;
      RECT 52.305 -57.505 52.445 -57.335 ;
      RECT 52.355 -56.318 52.445 -55.31 ;
      RECT 52.305 -55.715 52.445 -55.545 ;
      RECT 52.355 -54.51 52.445 -53.502 ;
      RECT 52.305 -54.275 52.445 -54.105 ;
      RECT 52.355 -53.088 52.445 -52.08 ;
      RECT 52.305 -52.485 52.445 -52.315 ;
      RECT 52.355 -51.28 52.445 -50.272 ;
      RECT 52.305 -51.045 52.445 -50.875 ;
      RECT 52.355 -49.858 52.445 -48.85 ;
      RECT 52.305 -49.255 52.445 -49.085 ;
      RECT 52.355 -48.05 52.445 -47.042 ;
      RECT 52.305 -47.815 52.445 -47.645 ;
      RECT 52.355 -46.628 52.445 -45.62 ;
      RECT 52.305 -46.025 52.445 -45.855 ;
      RECT 52.355 -44.82 52.445 -43.812 ;
      RECT 52.305 -44.585 52.445 -44.415 ;
      RECT 52.355 -43.398 52.445 -42.39 ;
      RECT 52.305 -42.795 52.445 -42.625 ;
      RECT 52.355 -41.59 52.445 -40.582 ;
      RECT 52.305 -41.355 52.445 -41.185 ;
      RECT 52.355 -40.168 52.445 -39.16 ;
      RECT 52.305 -39.565 52.445 -39.395 ;
      RECT 52.355 -38.36 52.445 -37.352 ;
      RECT 52.305 -38.125 52.445 -37.955 ;
      RECT 52.355 -36.938 52.445 -35.93 ;
      RECT 52.305 -36.335 52.445 -36.165 ;
      RECT 52.355 -35.13 52.445 -34.122 ;
      RECT 52.305 -34.895 52.445 -34.725 ;
      RECT 52.355 -33.708 52.445 -32.7 ;
      RECT 52.305 -33.105 52.445 -32.935 ;
      RECT 52.355 -31.9 52.445 -30.892 ;
      RECT 52.305 -31.665 52.445 -31.495 ;
      RECT 52.355 -30.478 52.445 -29.47 ;
      RECT 52.305 -29.875 52.445 -29.705 ;
      RECT 52.355 -28.67 52.445 -27.662 ;
      RECT 52.305 -28.435 52.445 -28.265 ;
      RECT 52.355 -27.248 52.445 -26.24 ;
      RECT 52.305 -26.645 52.445 -26.475 ;
      RECT 52.355 -25.44 52.445 -24.432 ;
      RECT 52.305 -25.205 52.445 -25.035 ;
      RECT 52.355 -24.018 52.445 -23.01 ;
      RECT 52.305 -23.415 52.445 -23.245 ;
      RECT 52.355 -22.21 52.445 -21.202 ;
      RECT 52.305 -21.975 52.445 -21.805 ;
      RECT 52.355 -20.788 52.445 -19.78 ;
      RECT 52.305 -20.185 52.445 -20.015 ;
      RECT 52.355 -18.98 52.445 -17.972 ;
      RECT 52.305 -18.745 52.445 -18.575 ;
      RECT 52.355 -17.558 52.445 -16.55 ;
      RECT 52.305 -16.955 52.445 -16.785 ;
      RECT 52.355 -15.75 52.445 -14.742 ;
      RECT 52.305 -15.515 52.445 -15.345 ;
      RECT 52.355 -14.328 52.445 -13.32 ;
      RECT 52.305 -13.725 52.445 -13.555 ;
      RECT 52.355 -12.52 52.445 -11.512 ;
      RECT 52.305 -12.285 52.445 -12.115 ;
      RECT 52.355 -11.098 52.445 -10.09 ;
      RECT 52.305 -10.495 52.445 -10.325 ;
      RECT 52.355 -9.29 52.445 -8.282 ;
      RECT 52.305 -9.055 52.445 -8.885 ;
      RECT 52.355 -7.868 52.445 -6.86 ;
      RECT 52.305 -7.265 52.445 -7.095 ;
      RECT 52.355 -6.06 52.445 -5.052 ;
      RECT 52.305 -5.825 52.445 -5.655 ;
      RECT 52.355 -4.638 52.445 -3.63 ;
      RECT 52.305 -4.035 52.445 -3.865 ;
      RECT 52.355 -2.83 52.445 -1.822 ;
      RECT 52.305 -2.595 52.445 -2.425 ;
      RECT 52.355 -1.408 52.445 -0.4 ;
      RECT 52.305 -0.805 52.445 -0.635 ;
      RECT 52.355 0.4 52.445 1.408 ;
      RECT 52.305 0.635 52.445 0.805 ;
      RECT 50.925 -111.685 52.405 -111.585 ;
      RECT 50.925 -112.195 51.025 -111.585 ;
      RECT 51.145 -109.15 52.405 -109.05 ;
      RECT 52.305 -109.475 52.405 -109.05 ;
      RECT 51.745 -109.475 51.845 -109.05 ;
      RECT 51.185 -109.475 51.285 -109.05 ;
      RECT 51.955 -101.538 52.045 -100.531 ;
      RECT 51.955 -101.225 52.095 -101.055 ;
      RECT 51.955 -99.729 52.045 -98.722 ;
      RECT 51.955 -99.205 52.095 -99.035 ;
      RECT 51.955 -98.308 52.045 -97.301 ;
      RECT 51.955 -97.995 52.095 -97.825 ;
      RECT 51.955 -96.499 52.045 -95.492 ;
      RECT 51.955 -95.975 52.095 -95.805 ;
      RECT 51.955 -95.078 52.045 -94.071 ;
      RECT 51.955 -94.765 52.095 -94.595 ;
      RECT 51.955 -93.269 52.045 -92.262 ;
      RECT 51.955 -92.745 52.095 -92.575 ;
      RECT 51.955 -91.848 52.045 -90.841 ;
      RECT 51.955 -91.535 52.095 -91.365 ;
      RECT 51.955 -90.039 52.045 -89.032 ;
      RECT 51.955 -89.515 52.095 -89.345 ;
      RECT 51.955 -88.618 52.045 -87.611 ;
      RECT 51.955 -88.305 52.095 -88.135 ;
      RECT 51.955 -86.809 52.045 -85.802 ;
      RECT 51.955 -86.285 52.095 -86.115 ;
      RECT 51.955 -85.388 52.045 -84.381 ;
      RECT 51.955 -85.075 52.095 -84.905 ;
      RECT 51.955 -83.579 52.045 -82.572 ;
      RECT 51.955 -83.055 52.095 -82.885 ;
      RECT 51.955 -82.158 52.045 -81.151 ;
      RECT 51.955 -81.845 52.095 -81.675 ;
      RECT 51.955 -80.349 52.045 -79.342 ;
      RECT 51.955 -79.825 52.095 -79.655 ;
      RECT 51.955 -78.928 52.045 -77.921 ;
      RECT 51.955 -78.615 52.095 -78.445 ;
      RECT 51.955 -77.119 52.045 -76.112 ;
      RECT 51.955 -76.595 52.095 -76.425 ;
      RECT 51.955 -75.698 52.045 -74.691 ;
      RECT 51.955 -75.385 52.095 -75.215 ;
      RECT 51.955 -73.889 52.045 -72.882 ;
      RECT 51.955 -73.365 52.095 -73.195 ;
      RECT 51.955 -72.468 52.045 -71.461 ;
      RECT 51.955 -72.155 52.095 -71.985 ;
      RECT 51.955 -70.659 52.045 -69.652 ;
      RECT 51.955 -70.135 52.095 -69.965 ;
      RECT 51.955 -69.238 52.045 -68.231 ;
      RECT 51.955 -68.925 52.095 -68.755 ;
      RECT 51.955 -67.429 52.045 -66.422 ;
      RECT 51.955 -66.905 52.095 -66.735 ;
      RECT 51.955 -66.008 52.045 -65.001 ;
      RECT 51.955 -65.695 52.095 -65.525 ;
      RECT 51.955 -64.199 52.045 -63.192 ;
      RECT 51.955 -63.675 52.095 -63.505 ;
      RECT 51.955 -62.778 52.045 -61.771 ;
      RECT 51.955 -62.465 52.095 -62.295 ;
      RECT 51.955 -60.969 52.045 -59.962 ;
      RECT 51.955 -60.445 52.095 -60.275 ;
      RECT 51.955 -59.548 52.045 -58.541 ;
      RECT 51.955 -59.235 52.095 -59.065 ;
      RECT 51.955 -57.739 52.045 -56.732 ;
      RECT 51.955 -57.215 52.095 -57.045 ;
      RECT 51.955 -56.318 52.045 -55.311 ;
      RECT 51.955 -56.005 52.095 -55.835 ;
      RECT 51.955 -54.509 52.045 -53.502 ;
      RECT 51.955 -53.985 52.095 -53.815 ;
      RECT 51.955 -53.088 52.045 -52.081 ;
      RECT 51.955 -52.775 52.095 -52.605 ;
      RECT 51.955 -51.279 52.045 -50.272 ;
      RECT 51.955 -50.755 52.095 -50.585 ;
      RECT 51.955 -49.858 52.045 -48.851 ;
      RECT 51.955 -49.545 52.095 -49.375 ;
      RECT 51.955 -48.049 52.045 -47.042 ;
      RECT 51.955 -47.525 52.095 -47.355 ;
      RECT 51.955 -46.628 52.045 -45.621 ;
      RECT 51.955 -46.315 52.095 -46.145 ;
      RECT 51.955 -44.819 52.045 -43.812 ;
      RECT 51.955 -44.295 52.095 -44.125 ;
      RECT 51.955 -43.398 52.045 -42.391 ;
      RECT 51.955 -43.085 52.095 -42.915 ;
      RECT 51.955 -41.589 52.045 -40.582 ;
      RECT 51.955 -41.065 52.095 -40.895 ;
      RECT 51.955 -40.168 52.045 -39.161 ;
      RECT 51.955 -39.855 52.095 -39.685 ;
      RECT 51.955 -38.359 52.045 -37.352 ;
      RECT 51.955 -37.835 52.095 -37.665 ;
      RECT 51.955 -36.938 52.045 -35.931 ;
      RECT 51.955 -36.625 52.095 -36.455 ;
      RECT 51.955 -35.129 52.045 -34.122 ;
      RECT 51.955 -34.605 52.095 -34.435 ;
      RECT 51.955 -33.708 52.045 -32.701 ;
      RECT 51.955 -33.395 52.095 -33.225 ;
      RECT 51.955 -31.899 52.045 -30.892 ;
      RECT 51.955 -31.375 52.095 -31.205 ;
      RECT 51.955 -30.478 52.045 -29.471 ;
      RECT 51.955 -30.165 52.095 -29.995 ;
      RECT 51.955 -28.669 52.045 -27.662 ;
      RECT 51.955 -28.145 52.095 -27.975 ;
      RECT 51.955 -27.248 52.045 -26.241 ;
      RECT 51.955 -26.935 52.095 -26.765 ;
      RECT 51.955 -25.439 52.045 -24.432 ;
      RECT 51.955 -24.915 52.095 -24.745 ;
      RECT 51.955 -24.018 52.045 -23.011 ;
      RECT 51.955 -23.705 52.095 -23.535 ;
      RECT 51.955 -22.209 52.045 -21.202 ;
      RECT 51.955 -21.685 52.095 -21.515 ;
      RECT 51.955 -20.788 52.045 -19.781 ;
      RECT 51.955 -20.475 52.095 -20.305 ;
      RECT 51.955 -18.979 52.045 -17.972 ;
      RECT 51.955 -18.455 52.095 -18.285 ;
      RECT 51.955 -17.558 52.045 -16.551 ;
      RECT 51.955 -17.245 52.095 -17.075 ;
      RECT 51.955 -15.749 52.045 -14.742 ;
      RECT 51.955 -15.225 52.095 -15.055 ;
      RECT 51.955 -14.328 52.045 -13.321 ;
      RECT 51.955 -14.015 52.095 -13.845 ;
      RECT 51.955 -12.519 52.045 -11.512 ;
      RECT 51.955 -11.995 52.095 -11.825 ;
      RECT 51.955 -11.098 52.045 -10.091 ;
      RECT 51.955 -10.785 52.095 -10.615 ;
      RECT 51.955 -9.289 52.045 -8.282 ;
      RECT 51.955 -8.765 52.095 -8.595 ;
      RECT 51.955 -7.868 52.045 -6.861 ;
      RECT 51.955 -7.555 52.095 -7.385 ;
      RECT 51.955 -6.059 52.045 -5.052 ;
      RECT 51.955 -5.535 52.095 -5.365 ;
      RECT 51.955 -4.638 52.045 -3.631 ;
      RECT 51.955 -4.325 52.095 -4.155 ;
      RECT 51.955 -2.829 52.045 -1.822 ;
      RECT 51.955 -2.305 52.095 -2.135 ;
      RECT 51.955 -1.408 52.045 -0.401 ;
      RECT 51.955 -1.095 52.095 -0.925 ;
      RECT 51.955 0.401 52.045 1.408 ;
      RECT 51.955 0.925 52.095 1.095 ;
      RECT 51.285 -111.495 51.455 -111.385 ;
      RECT 48.135 -111.495 51.455 -111.395 ;
      RECT 51.155 -101.538 51.245 -100.53 ;
      RECT 51.105 -100.935 51.245 -100.765 ;
      RECT 51.155 -99.73 51.245 -98.722 ;
      RECT 51.105 -99.495 51.245 -99.325 ;
      RECT 51.155 -98.308 51.245 -97.3 ;
      RECT 51.105 -97.705 51.245 -97.535 ;
      RECT 51.155 -96.5 51.245 -95.492 ;
      RECT 51.105 -96.265 51.245 -96.095 ;
      RECT 51.155 -95.078 51.245 -94.07 ;
      RECT 51.105 -94.475 51.245 -94.305 ;
      RECT 51.155 -93.27 51.245 -92.262 ;
      RECT 51.105 -93.035 51.245 -92.865 ;
      RECT 51.155 -91.848 51.245 -90.84 ;
      RECT 51.105 -91.245 51.245 -91.075 ;
      RECT 51.155 -90.04 51.245 -89.032 ;
      RECT 51.105 -89.805 51.245 -89.635 ;
      RECT 51.155 -88.618 51.245 -87.61 ;
      RECT 51.105 -88.015 51.245 -87.845 ;
      RECT 51.155 -86.81 51.245 -85.802 ;
      RECT 51.105 -86.575 51.245 -86.405 ;
      RECT 51.155 -85.388 51.245 -84.38 ;
      RECT 51.105 -84.785 51.245 -84.615 ;
      RECT 51.155 -83.58 51.245 -82.572 ;
      RECT 51.105 -83.345 51.245 -83.175 ;
      RECT 51.155 -82.158 51.245 -81.15 ;
      RECT 51.105 -81.555 51.245 -81.385 ;
      RECT 51.155 -80.35 51.245 -79.342 ;
      RECT 51.105 -80.115 51.245 -79.945 ;
      RECT 51.155 -78.928 51.245 -77.92 ;
      RECT 51.105 -78.325 51.245 -78.155 ;
      RECT 51.155 -77.12 51.245 -76.112 ;
      RECT 51.105 -76.885 51.245 -76.715 ;
      RECT 51.155 -75.698 51.245 -74.69 ;
      RECT 51.105 -75.095 51.245 -74.925 ;
      RECT 51.155 -73.89 51.245 -72.882 ;
      RECT 51.105 -73.655 51.245 -73.485 ;
      RECT 51.155 -72.468 51.245 -71.46 ;
      RECT 51.105 -71.865 51.245 -71.695 ;
      RECT 51.155 -70.66 51.245 -69.652 ;
      RECT 51.105 -70.425 51.245 -70.255 ;
      RECT 51.155 -69.238 51.245 -68.23 ;
      RECT 51.105 -68.635 51.245 -68.465 ;
      RECT 51.155 -67.43 51.245 -66.422 ;
      RECT 51.105 -67.195 51.245 -67.025 ;
      RECT 51.155 -66.008 51.245 -65 ;
      RECT 51.105 -65.405 51.245 -65.235 ;
      RECT 51.155 -64.2 51.245 -63.192 ;
      RECT 51.105 -63.965 51.245 -63.795 ;
      RECT 51.155 -62.778 51.245 -61.77 ;
      RECT 51.105 -62.175 51.245 -62.005 ;
      RECT 51.155 -60.97 51.245 -59.962 ;
      RECT 51.105 -60.735 51.245 -60.565 ;
      RECT 51.155 -59.548 51.245 -58.54 ;
      RECT 51.105 -58.945 51.245 -58.775 ;
      RECT 51.155 -57.74 51.245 -56.732 ;
      RECT 51.105 -57.505 51.245 -57.335 ;
      RECT 51.155 -56.318 51.245 -55.31 ;
      RECT 51.105 -55.715 51.245 -55.545 ;
      RECT 51.155 -54.51 51.245 -53.502 ;
      RECT 51.105 -54.275 51.245 -54.105 ;
      RECT 51.155 -53.088 51.245 -52.08 ;
      RECT 51.105 -52.485 51.245 -52.315 ;
      RECT 51.155 -51.28 51.245 -50.272 ;
      RECT 51.105 -51.045 51.245 -50.875 ;
      RECT 51.155 -49.858 51.245 -48.85 ;
      RECT 51.105 -49.255 51.245 -49.085 ;
      RECT 51.155 -48.05 51.245 -47.042 ;
      RECT 51.105 -47.815 51.245 -47.645 ;
      RECT 51.155 -46.628 51.245 -45.62 ;
      RECT 51.105 -46.025 51.245 -45.855 ;
      RECT 51.155 -44.82 51.245 -43.812 ;
      RECT 51.105 -44.585 51.245 -44.415 ;
      RECT 51.155 -43.398 51.245 -42.39 ;
      RECT 51.105 -42.795 51.245 -42.625 ;
      RECT 51.155 -41.59 51.245 -40.582 ;
      RECT 51.105 -41.355 51.245 -41.185 ;
      RECT 51.155 -40.168 51.245 -39.16 ;
      RECT 51.105 -39.565 51.245 -39.395 ;
      RECT 51.155 -38.36 51.245 -37.352 ;
      RECT 51.105 -38.125 51.245 -37.955 ;
      RECT 51.155 -36.938 51.245 -35.93 ;
      RECT 51.105 -36.335 51.245 -36.165 ;
      RECT 51.155 -35.13 51.245 -34.122 ;
      RECT 51.105 -34.895 51.245 -34.725 ;
      RECT 51.155 -33.708 51.245 -32.7 ;
      RECT 51.105 -33.105 51.245 -32.935 ;
      RECT 51.155 -31.9 51.245 -30.892 ;
      RECT 51.105 -31.665 51.245 -31.495 ;
      RECT 51.155 -30.478 51.245 -29.47 ;
      RECT 51.105 -29.875 51.245 -29.705 ;
      RECT 51.155 -28.67 51.245 -27.662 ;
      RECT 51.105 -28.435 51.245 -28.265 ;
      RECT 51.155 -27.248 51.245 -26.24 ;
      RECT 51.105 -26.645 51.245 -26.475 ;
      RECT 51.155 -25.44 51.245 -24.432 ;
      RECT 51.105 -25.205 51.245 -25.035 ;
      RECT 51.155 -24.018 51.245 -23.01 ;
      RECT 51.105 -23.415 51.245 -23.245 ;
      RECT 51.155 -22.21 51.245 -21.202 ;
      RECT 51.105 -21.975 51.245 -21.805 ;
      RECT 51.155 -20.788 51.245 -19.78 ;
      RECT 51.105 -20.185 51.245 -20.015 ;
      RECT 51.155 -18.98 51.245 -17.972 ;
      RECT 51.105 -18.745 51.245 -18.575 ;
      RECT 51.155 -17.558 51.245 -16.55 ;
      RECT 51.105 -16.955 51.245 -16.785 ;
      RECT 51.155 -15.75 51.245 -14.742 ;
      RECT 51.105 -15.515 51.245 -15.345 ;
      RECT 51.155 -14.328 51.245 -13.32 ;
      RECT 51.105 -13.725 51.245 -13.555 ;
      RECT 51.155 -12.52 51.245 -11.512 ;
      RECT 51.105 -12.285 51.245 -12.115 ;
      RECT 51.155 -11.098 51.245 -10.09 ;
      RECT 51.105 -10.495 51.245 -10.325 ;
      RECT 51.155 -9.29 51.245 -8.282 ;
      RECT 51.105 -9.055 51.245 -8.885 ;
      RECT 51.155 -7.868 51.245 -6.86 ;
      RECT 51.105 -7.265 51.245 -7.095 ;
      RECT 51.155 -6.06 51.245 -5.052 ;
      RECT 51.105 -5.825 51.245 -5.655 ;
      RECT 51.155 -4.638 51.245 -3.63 ;
      RECT 51.105 -4.035 51.245 -3.865 ;
      RECT 51.155 -2.83 51.245 -1.822 ;
      RECT 51.105 -2.595 51.245 -2.425 ;
      RECT 51.155 -1.408 51.245 -0.4 ;
      RECT 51.105 -0.805 51.245 -0.635 ;
      RECT 51.155 0.4 51.245 1.408 ;
      RECT 51.105 0.635 51.245 0.805 ;
      RECT 50.755 -101.538 50.845 -100.531 ;
      RECT 50.755 -101.225 50.895 -101.055 ;
      RECT 50.755 -99.729 50.845 -98.722 ;
      RECT 50.755 -99.205 50.895 -99.035 ;
      RECT 50.755 -98.308 50.845 -97.301 ;
      RECT 50.755 -97.995 50.895 -97.825 ;
      RECT 50.755 -96.499 50.845 -95.492 ;
      RECT 50.755 -95.975 50.895 -95.805 ;
      RECT 50.755 -95.078 50.845 -94.071 ;
      RECT 50.755 -94.765 50.895 -94.595 ;
      RECT 50.755 -93.269 50.845 -92.262 ;
      RECT 50.755 -92.745 50.895 -92.575 ;
      RECT 50.755 -91.848 50.845 -90.841 ;
      RECT 50.755 -91.535 50.895 -91.365 ;
      RECT 50.755 -90.039 50.845 -89.032 ;
      RECT 50.755 -89.515 50.895 -89.345 ;
      RECT 50.755 -88.618 50.845 -87.611 ;
      RECT 50.755 -88.305 50.895 -88.135 ;
      RECT 50.755 -86.809 50.845 -85.802 ;
      RECT 50.755 -86.285 50.895 -86.115 ;
      RECT 50.755 -85.388 50.845 -84.381 ;
      RECT 50.755 -85.075 50.895 -84.905 ;
      RECT 50.755 -83.579 50.845 -82.572 ;
      RECT 50.755 -83.055 50.895 -82.885 ;
      RECT 50.755 -82.158 50.845 -81.151 ;
      RECT 50.755 -81.845 50.895 -81.675 ;
      RECT 50.755 -80.349 50.845 -79.342 ;
      RECT 50.755 -79.825 50.895 -79.655 ;
      RECT 50.755 -78.928 50.845 -77.921 ;
      RECT 50.755 -78.615 50.895 -78.445 ;
      RECT 50.755 -77.119 50.845 -76.112 ;
      RECT 50.755 -76.595 50.895 -76.425 ;
      RECT 50.755 -75.698 50.845 -74.691 ;
      RECT 50.755 -75.385 50.895 -75.215 ;
      RECT 50.755 -73.889 50.845 -72.882 ;
      RECT 50.755 -73.365 50.895 -73.195 ;
      RECT 50.755 -72.468 50.845 -71.461 ;
      RECT 50.755 -72.155 50.895 -71.985 ;
      RECT 50.755 -70.659 50.845 -69.652 ;
      RECT 50.755 -70.135 50.895 -69.965 ;
      RECT 50.755 -69.238 50.845 -68.231 ;
      RECT 50.755 -68.925 50.895 -68.755 ;
      RECT 50.755 -67.429 50.845 -66.422 ;
      RECT 50.755 -66.905 50.895 -66.735 ;
      RECT 50.755 -66.008 50.845 -65.001 ;
      RECT 50.755 -65.695 50.895 -65.525 ;
      RECT 50.755 -64.199 50.845 -63.192 ;
      RECT 50.755 -63.675 50.895 -63.505 ;
      RECT 50.755 -62.778 50.845 -61.771 ;
      RECT 50.755 -62.465 50.895 -62.295 ;
      RECT 50.755 -60.969 50.845 -59.962 ;
      RECT 50.755 -60.445 50.895 -60.275 ;
      RECT 50.755 -59.548 50.845 -58.541 ;
      RECT 50.755 -59.235 50.895 -59.065 ;
      RECT 50.755 -57.739 50.845 -56.732 ;
      RECT 50.755 -57.215 50.895 -57.045 ;
      RECT 50.755 -56.318 50.845 -55.311 ;
      RECT 50.755 -56.005 50.895 -55.835 ;
      RECT 50.755 -54.509 50.845 -53.502 ;
      RECT 50.755 -53.985 50.895 -53.815 ;
      RECT 50.755 -53.088 50.845 -52.081 ;
      RECT 50.755 -52.775 50.895 -52.605 ;
      RECT 50.755 -51.279 50.845 -50.272 ;
      RECT 50.755 -50.755 50.895 -50.585 ;
      RECT 50.755 -49.858 50.845 -48.851 ;
      RECT 50.755 -49.545 50.895 -49.375 ;
      RECT 50.755 -48.049 50.845 -47.042 ;
      RECT 50.755 -47.525 50.895 -47.355 ;
      RECT 50.755 -46.628 50.845 -45.621 ;
      RECT 50.755 -46.315 50.895 -46.145 ;
      RECT 50.755 -44.819 50.845 -43.812 ;
      RECT 50.755 -44.295 50.895 -44.125 ;
      RECT 50.755 -43.398 50.845 -42.391 ;
      RECT 50.755 -43.085 50.895 -42.915 ;
      RECT 50.755 -41.589 50.845 -40.582 ;
      RECT 50.755 -41.065 50.895 -40.895 ;
      RECT 50.755 -40.168 50.845 -39.161 ;
      RECT 50.755 -39.855 50.895 -39.685 ;
      RECT 50.755 -38.359 50.845 -37.352 ;
      RECT 50.755 -37.835 50.895 -37.665 ;
      RECT 50.755 -36.938 50.845 -35.931 ;
      RECT 50.755 -36.625 50.895 -36.455 ;
      RECT 50.755 -35.129 50.845 -34.122 ;
      RECT 50.755 -34.605 50.895 -34.435 ;
      RECT 50.755 -33.708 50.845 -32.701 ;
      RECT 50.755 -33.395 50.895 -33.225 ;
      RECT 50.755 -31.899 50.845 -30.892 ;
      RECT 50.755 -31.375 50.895 -31.205 ;
      RECT 50.755 -30.478 50.845 -29.471 ;
      RECT 50.755 -30.165 50.895 -29.995 ;
      RECT 50.755 -28.669 50.845 -27.662 ;
      RECT 50.755 -28.145 50.895 -27.975 ;
      RECT 50.755 -27.248 50.845 -26.241 ;
      RECT 50.755 -26.935 50.895 -26.765 ;
      RECT 50.755 -25.439 50.845 -24.432 ;
      RECT 50.755 -24.915 50.895 -24.745 ;
      RECT 50.755 -24.018 50.845 -23.011 ;
      RECT 50.755 -23.705 50.895 -23.535 ;
      RECT 50.755 -22.209 50.845 -21.202 ;
      RECT 50.755 -21.685 50.895 -21.515 ;
      RECT 50.755 -20.788 50.845 -19.781 ;
      RECT 50.755 -20.475 50.895 -20.305 ;
      RECT 50.755 -18.979 50.845 -17.972 ;
      RECT 50.755 -18.455 50.895 -18.285 ;
      RECT 50.755 -17.558 50.845 -16.551 ;
      RECT 50.755 -17.245 50.895 -17.075 ;
      RECT 50.755 -15.749 50.845 -14.742 ;
      RECT 50.755 -15.225 50.895 -15.055 ;
      RECT 50.755 -14.328 50.845 -13.321 ;
      RECT 50.755 -14.015 50.895 -13.845 ;
      RECT 50.755 -12.519 50.845 -11.512 ;
      RECT 50.755 -11.995 50.895 -11.825 ;
      RECT 50.755 -11.098 50.845 -10.091 ;
      RECT 50.755 -10.785 50.895 -10.615 ;
      RECT 50.755 -9.289 50.845 -8.282 ;
      RECT 50.755 -8.765 50.895 -8.595 ;
      RECT 50.755 -7.868 50.845 -6.861 ;
      RECT 50.755 -7.555 50.895 -7.385 ;
      RECT 50.755 -6.059 50.845 -5.052 ;
      RECT 50.755 -5.535 50.895 -5.365 ;
      RECT 50.755 -4.638 50.845 -3.631 ;
      RECT 50.755 -4.325 50.895 -4.155 ;
      RECT 50.755 -2.829 50.845 -1.822 ;
      RECT 50.755 -2.305 50.895 -2.135 ;
      RECT 50.755 -1.408 50.845 -0.401 ;
      RECT 50.755 -1.095 50.895 -0.925 ;
      RECT 50.755 0.401 50.845 1.408 ;
      RECT 50.755 0.925 50.895 1.095 ;
      RECT 48.905 -111.685 50.385 -111.585 ;
      RECT 48.905 -112.055 49.005 -111.585 ;
      RECT 48.71 -114.395 50.285 -114.275 ;
      RECT 50.185 -114.895 50.285 -114.275 ;
      RECT 49.59 -114.895 49.69 -114.275 ;
      RECT 48.71 -114.85 48.81 -114.275 ;
      RECT 49.955 -101.538 50.045 -100.53 ;
      RECT 49.905 -100.935 50.045 -100.765 ;
      RECT 49.955 -99.73 50.045 -98.722 ;
      RECT 49.905 -99.495 50.045 -99.325 ;
      RECT 49.955 -98.308 50.045 -97.3 ;
      RECT 49.905 -97.705 50.045 -97.535 ;
      RECT 49.955 -96.5 50.045 -95.492 ;
      RECT 49.905 -96.265 50.045 -96.095 ;
      RECT 49.955 -95.078 50.045 -94.07 ;
      RECT 49.905 -94.475 50.045 -94.305 ;
      RECT 49.955 -93.27 50.045 -92.262 ;
      RECT 49.905 -93.035 50.045 -92.865 ;
      RECT 49.955 -91.848 50.045 -90.84 ;
      RECT 49.905 -91.245 50.045 -91.075 ;
      RECT 49.955 -90.04 50.045 -89.032 ;
      RECT 49.905 -89.805 50.045 -89.635 ;
      RECT 49.955 -88.618 50.045 -87.61 ;
      RECT 49.905 -88.015 50.045 -87.845 ;
      RECT 49.955 -86.81 50.045 -85.802 ;
      RECT 49.905 -86.575 50.045 -86.405 ;
      RECT 49.955 -85.388 50.045 -84.38 ;
      RECT 49.905 -84.785 50.045 -84.615 ;
      RECT 49.955 -83.58 50.045 -82.572 ;
      RECT 49.905 -83.345 50.045 -83.175 ;
      RECT 49.955 -82.158 50.045 -81.15 ;
      RECT 49.905 -81.555 50.045 -81.385 ;
      RECT 49.955 -80.35 50.045 -79.342 ;
      RECT 49.905 -80.115 50.045 -79.945 ;
      RECT 49.955 -78.928 50.045 -77.92 ;
      RECT 49.905 -78.325 50.045 -78.155 ;
      RECT 49.955 -77.12 50.045 -76.112 ;
      RECT 49.905 -76.885 50.045 -76.715 ;
      RECT 49.955 -75.698 50.045 -74.69 ;
      RECT 49.905 -75.095 50.045 -74.925 ;
      RECT 49.955 -73.89 50.045 -72.882 ;
      RECT 49.905 -73.655 50.045 -73.485 ;
      RECT 49.955 -72.468 50.045 -71.46 ;
      RECT 49.905 -71.865 50.045 -71.695 ;
      RECT 49.955 -70.66 50.045 -69.652 ;
      RECT 49.905 -70.425 50.045 -70.255 ;
      RECT 49.955 -69.238 50.045 -68.23 ;
      RECT 49.905 -68.635 50.045 -68.465 ;
      RECT 49.955 -67.43 50.045 -66.422 ;
      RECT 49.905 -67.195 50.045 -67.025 ;
      RECT 49.955 -66.008 50.045 -65 ;
      RECT 49.905 -65.405 50.045 -65.235 ;
      RECT 49.955 -64.2 50.045 -63.192 ;
      RECT 49.905 -63.965 50.045 -63.795 ;
      RECT 49.955 -62.778 50.045 -61.77 ;
      RECT 49.905 -62.175 50.045 -62.005 ;
      RECT 49.955 -60.97 50.045 -59.962 ;
      RECT 49.905 -60.735 50.045 -60.565 ;
      RECT 49.955 -59.548 50.045 -58.54 ;
      RECT 49.905 -58.945 50.045 -58.775 ;
      RECT 49.955 -57.74 50.045 -56.732 ;
      RECT 49.905 -57.505 50.045 -57.335 ;
      RECT 49.955 -56.318 50.045 -55.31 ;
      RECT 49.905 -55.715 50.045 -55.545 ;
      RECT 49.955 -54.51 50.045 -53.502 ;
      RECT 49.905 -54.275 50.045 -54.105 ;
      RECT 49.955 -53.088 50.045 -52.08 ;
      RECT 49.905 -52.485 50.045 -52.315 ;
      RECT 49.955 -51.28 50.045 -50.272 ;
      RECT 49.905 -51.045 50.045 -50.875 ;
      RECT 49.955 -49.858 50.045 -48.85 ;
      RECT 49.905 -49.255 50.045 -49.085 ;
      RECT 49.955 -48.05 50.045 -47.042 ;
      RECT 49.905 -47.815 50.045 -47.645 ;
      RECT 49.955 -46.628 50.045 -45.62 ;
      RECT 49.905 -46.025 50.045 -45.855 ;
      RECT 49.955 -44.82 50.045 -43.812 ;
      RECT 49.905 -44.585 50.045 -44.415 ;
      RECT 49.955 -43.398 50.045 -42.39 ;
      RECT 49.905 -42.795 50.045 -42.625 ;
      RECT 49.955 -41.59 50.045 -40.582 ;
      RECT 49.905 -41.355 50.045 -41.185 ;
      RECT 49.955 -40.168 50.045 -39.16 ;
      RECT 49.905 -39.565 50.045 -39.395 ;
      RECT 49.955 -38.36 50.045 -37.352 ;
      RECT 49.905 -38.125 50.045 -37.955 ;
      RECT 49.955 -36.938 50.045 -35.93 ;
      RECT 49.905 -36.335 50.045 -36.165 ;
      RECT 49.955 -35.13 50.045 -34.122 ;
      RECT 49.905 -34.895 50.045 -34.725 ;
      RECT 49.955 -33.708 50.045 -32.7 ;
      RECT 49.905 -33.105 50.045 -32.935 ;
      RECT 49.955 -31.9 50.045 -30.892 ;
      RECT 49.905 -31.665 50.045 -31.495 ;
      RECT 49.955 -30.478 50.045 -29.47 ;
      RECT 49.905 -29.875 50.045 -29.705 ;
      RECT 49.955 -28.67 50.045 -27.662 ;
      RECT 49.905 -28.435 50.045 -28.265 ;
      RECT 49.955 -27.248 50.045 -26.24 ;
      RECT 49.905 -26.645 50.045 -26.475 ;
      RECT 49.955 -25.44 50.045 -24.432 ;
      RECT 49.905 -25.205 50.045 -25.035 ;
      RECT 49.955 -24.018 50.045 -23.01 ;
      RECT 49.905 -23.415 50.045 -23.245 ;
      RECT 49.955 -22.21 50.045 -21.202 ;
      RECT 49.905 -21.975 50.045 -21.805 ;
      RECT 49.955 -20.788 50.045 -19.78 ;
      RECT 49.905 -20.185 50.045 -20.015 ;
      RECT 49.955 -18.98 50.045 -17.972 ;
      RECT 49.905 -18.745 50.045 -18.575 ;
      RECT 49.955 -17.558 50.045 -16.55 ;
      RECT 49.905 -16.955 50.045 -16.785 ;
      RECT 49.955 -15.75 50.045 -14.742 ;
      RECT 49.905 -15.515 50.045 -15.345 ;
      RECT 49.955 -14.328 50.045 -13.32 ;
      RECT 49.905 -13.725 50.045 -13.555 ;
      RECT 49.955 -12.52 50.045 -11.512 ;
      RECT 49.905 -12.285 50.045 -12.115 ;
      RECT 49.955 -11.098 50.045 -10.09 ;
      RECT 49.905 -10.495 50.045 -10.325 ;
      RECT 49.955 -9.29 50.045 -8.282 ;
      RECT 49.905 -9.055 50.045 -8.885 ;
      RECT 49.955 -7.868 50.045 -6.86 ;
      RECT 49.905 -7.265 50.045 -7.095 ;
      RECT 49.955 -6.06 50.045 -5.052 ;
      RECT 49.905 -5.825 50.045 -5.655 ;
      RECT 49.955 -4.638 50.045 -3.63 ;
      RECT 49.905 -4.035 50.045 -3.865 ;
      RECT 49.955 -2.83 50.045 -1.822 ;
      RECT 49.905 -2.595 50.045 -2.425 ;
      RECT 49.955 -1.408 50.045 -0.4 ;
      RECT 49.905 -0.805 50.045 -0.635 ;
      RECT 49.955 0.4 50.045 1.408 ;
      RECT 49.905 0.635 50.045 0.805 ;
      RECT 49.83 -114.685 50.005 -114.515 ;
      RECT 49.905 -114.895 50.005 -114.515 ;
      RECT 48.945 -113.555 49.045 -113.09 ;
      RECT 49.31 -113.555 49.41 -113.1 ;
      RECT 48.945 -113.555 49.79 -113.385 ;
      RECT 49.555 -101.538 49.645 -100.531 ;
      RECT 49.555 -101.225 49.695 -101.055 ;
      RECT 49.555 -99.729 49.645 -98.722 ;
      RECT 49.555 -99.205 49.695 -99.035 ;
      RECT 49.555 -98.308 49.645 -97.301 ;
      RECT 49.555 -97.995 49.695 -97.825 ;
      RECT 49.555 -96.499 49.645 -95.492 ;
      RECT 49.555 -95.975 49.695 -95.805 ;
      RECT 49.555 -95.078 49.645 -94.071 ;
      RECT 49.555 -94.765 49.695 -94.595 ;
      RECT 49.555 -93.269 49.645 -92.262 ;
      RECT 49.555 -92.745 49.695 -92.575 ;
      RECT 49.555 -91.848 49.645 -90.841 ;
      RECT 49.555 -91.535 49.695 -91.365 ;
      RECT 49.555 -90.039 49.645 -89.032 ;
      RECT 49.555 -89.515 49.695 -89.345 ;
      RECT 49.555 -88.618 49.645 -87.611 ;
      RECT 49.555 -88.305 49.695 -88.135 ;
      RECT 49.555 -86.809 49.645 -85.802 ;
      RECT 49.555 -86.285 49.695 -86.115 ;
      RECT 49.555 -85.388 49.645 -84.381 ;
      RECT 49.555 -85.075 49.695 -84.905 ;
      RECT 49.555 -83.579 49.645 -82.572 ;
      RECT 49.555 -83.055 49.695 -82.885 ;
      RECT 49.555 -82.158 49.645 -81.151 ;
      RECT 49.555 -81.845 49.695 -81.675 ;
      RECT 49.555 -80.349 49.645 -79.342 ;
      RECT 49.555 -79.825 49.695 -79.655 ;
      RECT 49.555 -78.928 49.645 -77.921 ;
      RECT 49.555 -78.615 49.695 -78.445 ;
      RECT 49.555 -77.119 49.645 -76.112 ;
      RECT 49.555 -76.595 49.695 -76.425 ;
      RECT 49.555 -75.698 49.645 -74.691 ;
      RECT 49.555 -75.385 49.695 -75.215 ;
      RECT 49.555 -73.889 49.645 -72.882 ;
      RECT 49.555 -73.365 49.695 -73.195 ;
      RECT 49.555 -72.468 49.645 -71.461 ;
      RECT 49.555 -72.155 49.695 -71.985 ;
      RECT 49.555 -70.659 49.645 -69.652 ;
      RECT 49.555 -70.135 49.695 -69.965 ;
      RECT 49.555 -69.238 49.645 -68.231 ;
      RECT 49.555 -68.925 49.695 -68.755 ;
      RECT 49.555 -67.429 49.645 -66.422 ;
      RECT 49.555 -66.905 49.695 -66.735 ;
      RECT 49.555 -66.008 49.645 -65.001 ;
      RECT 49.555 -65.695 49.695 -65.525 ;
      RECT 49.555 -64.199 49.645 -63.192 ;
      RECT 49.555 -63.675 49.695 -63.505 ;
      RECT 49.555 -62.778 49.645 -61.771 ;
      RECT 49.555 -62.465 49.695 -62.295 ;
      RECT 49.555 -60.969 49.645 -59.962 ;
      RECT 49.555 -60.445 49.695 -60.275 ;
      RECT 49.555 -59.548 49.645 -58.541 ;
      RECT 49.555 -59.235 49.695 -59.065 ;
      RECT 49.555 -57.739 49.645 -56.732 ;
      RECT 49.555 -57.215 49.695 -57.045 ;
      RECT 49.555 -56.318 49.645 -55.311 ;
      RECT 49.555 -56.005 49.695 -55.835 ;
      RECT 49.555 -54.509 49.645 -53.502 ;
      RECT 49.555 -53.985 49.695 -53.815 ;
      RECT 49.555 -53.088 49.645 -52.081 ;
      RECT 49.555 -52.775 49.695 -52.605 ;
      RECT 49.555 -51.279 49.645 -50.272 ;
      RECT 49.555 -50.755 49.695 -50.585 ;
      RECT 49.555 -49.858 49.645 -48.851 ;
      RECT 49.555 -49.545 49.695 -49.375 ;
      RECT 49.555 -48.049 49.645 -47.042 ;
      RECT 49.555 -47.525 49.695 -47.355 ;
      RECT 49.555 -46.628 49.645 -45.621 ;
      RECT 49.555 -46.315 49.695 -46.145 ;
      RECT 49.555 -44.819 49.645 -43.812 ;
      RECT 49.555 -44.295 49.695 -44.125 ;
      RECT 49.555 -43.398 49.645 -42.391 ;
      RECT 49.555 -43.085 49.695 -42.915 ;
      RECT 49.555 -41.589 49.645 -40.582 ;
      RECT 49.555 -41.065 49.695 -40.895 ;
      RECT 49.555 -40.168 49.645 -39.161 ;
      RECT 49.555 -39.855 49.695 -39.685 ;
      RECT 49.555 -38.359 49.645 -37.352 ;
      RECT 49.555 -37.835 49.695 -37.665 ;
      RECT 49.555 -36.938 49.645 -35.931 ;
      RECT 49.555 -36.625 49.695 -36.455 ;
      RECT 49.555 -35.129 49.645 -34.122 ;
      RECT 49.555 -34.605 49.695 -34.435 ;
      RECT 49.555 -33.708 49.645 -32.701 ;
      RECT 49.555 -33.395 49.695 -33.225 ;
      RECT 49.555 -31.899 49.645 -30.892 ;
      RECT 49.555 -31.375 49.695 -31.205 ;
      RECT 49.555 -30.478 49.645 -29.471 ;
      RECT 49.555 -30.165 49.695 -29.995 ;
      RECT 49.555 -28.669 49.645 -27.662 ;
      RECT 49.555 -28.145 49.695 -27.975 ;
      RECT 49.555 -27.248 49.645 -26.241 ;
      RECT 49.555 -26.935 49.695 -26.765 ;
      RECT 49.555 -25.439 49.645 -24.432 ;
      RECT 49.555 -24.915 49.695 -24.745 ;
      RECT 49.555 -24.018 49.645 -23.011 ;
      RECT 49.555 -23.705 49.695 -23.535 ;
      RECT 49.555 -22.209 49.645 -21.202 ;
      RECT 49.555 -21.685 49.695 -21.515 ;
      RECT 49.555 -20.788 49.645 -19.781 ;
      RECT 49.555 -20.475 49.695 -20.305 ;
      RECT 49.555 -18.979 49.645 -17.972 ;
      RECT 49.555 -18.455 49.695 -18.285 ;
      RECT 49.555 -17.558 49.645 -16.551 ;
      RECT 49.555 -17.245 49.695 -17.075 ;
      RECT 49.555 -15.749 49.645 -14.742 ;
      RECT 49.555 -15.225 49.695 -15.055 ;
      RECT 49.555 -14.328 49.645 -13.321 ;
      RECT 49.555 -14.015 49.695 -13.845 ;
      RECT 49.555 -12.519 49.645 -11.512 ;
      RECT 49.555 -11.995 49.695 -11.825 ;
      RECT 49.555 -11.098 49.645 -10.091 ;
      RECT 49.555 -10.785 49.695 -10.615 ;
      RECT 49.555 -9.289 49.645 -8.282 ;
      RECT 49.555 -8.765 49.695 -8.595 ;
      RECT 49.555 -7.868 49.645 -6.861 ;
      RECT 49.555 -7.555 49.695 -7.385 ;
      RECT 49.555 -6.059 49.645 -5.052 ;
      RECT 49.555 -5.535 49.695 -5.365 ;
      RECT 49.555 -4.638 49.645 -3.631 ;
      RECT 49.555 -4.325 49.695 -4.155 ;
      RECT 49.555 -2.829 49.645 -1.822 ;
      RECT 49.555 -2.305 49.695 -2.135 ;
      RECT 49.555 -1.408 49.645 -0.401 ;
      RECT 49.555 -1.095 49.695 -0.925 ;
      RECT 49.555 0.401 49.645 1.408 ;
      RECT 49.555 0.925 49.695 1.095 ;
      RECT 49.24 -114.685 49.41 -114.515 ;
      RECT 49.31 -114.895 49.41 -114.515 ;
      RECT 48.755 -101.538 48.845 -100.53 ;
      RECT 48.705 -100.935 48.845 -100.765 ;
      RECT 48.755 -99.73 48.845 -98.722 ;
      RECT 48.705 -99.495 48.845 -99.325 ;
      RECT 48.755 -98.308 48.845 -97.3 ;
      RECT 48.705 -97.705 48.845 -97.535 ;
      RECT 48.755 -96.5 48.845 -95.492 ;
      RECT 48.705 -96.265 48.845 -96.095 ;
      RECT 48.755 -95.078 48.845 -94.07 ;
      RECT 48.705 -94.475 48.845 -94.305 ;
      RECT 48.755 -93.27 48.845 -92.262 ;
      RECT 48.705 -93.035 48.845 -92.865 ;
      RECT 48.755 -91.848 48.845 -90.84 ;
      RECT 48.705 -91.245 48.845 -91.075 ;
      RECT 48.755 -90.04 48.845 -89.032 ;
      RECT 48.705 -89.805 48.845 -89.635 ;
      RECT 48.755 -88.618 48.845 -87.61 ;
      RECT 48.705 -88.015 48.845 -87.845 ;
      RECT 48.755 -86.81 48.845 -85.802 ;
      RECT 48.705 -86.575 48.845 -86.405 ;
      RECT 48.755 -85.388 48.845 -84.38 ;
      RECT 48.705 -84.785 48.845 -84.615 ;
      RECT 48.755 -83.58 48.845 -82.572 ;
      RECT 48.705 -83.345 48.845 -83.175 ;
      RECT 48.755 -82.158 48.845 -81.15 ;
      RECT 48.705 -81.555 48.845 -81.385 ;
      RECT 48.755 -80.35 48.845 -79.342 ;
      RECT 48.705 -80.115 48.845 -79.945 ;
      RECT 48.755 -78.928 48.845 -77.92 ;
      RECT 48.705 -78.325 48.845 -78.155 ;
      RECT 48.755 -77.12 48.845 -76.112 ;
      RECT 48.705 -76.885 48.845 -76.715 ;
      RECT 48.755 -75.698 48.845 -74.69 ;
      RECT 48.705 -75.095 48.845 -74.925 ;
      RECT 48.755 -73.89 48.845 -72.882 ;
      RECT 48.705 -73.655 48.845 -73.485 ;
      RECT 48.755 -72.468 48.845 -71.46 ;
      RECT 48.705 -71.865 48.845 -71.695 ;
      RECT 48.755 -70.66 48.845 -69.652 ;
      RECT 48.705 -70.425 48.845 -70.255 ;
      RECT 48.755 -69.238 48.845 -68.23 ;
      RECT 48.705 -68.635 48.845 -68.465 ;
      RECT 48.755 -67.43 48.845 -66.422 ;
      RECT 48.705 -67.195 48.845 -67.025 ;
      RECT 48.755 -66.008 48.845 -65 ;
      RECT 48.705 -65.405 48.845 -65.235 ;
      RECT 48.755 -64.2 48.845 -63.192 ;
      RECT 48.705 -63.965 48.845 -63.795 ;
      RECT 48.755 -62.778 48.845 -61.77 ;
      RECT 48.705 -62.175 48.845 -62.005 ;
      RECT 48.755 -60.97 48.845 -59.962 ;
      RECT 48.705 -60.735 48.845 -60.565 ;
      RECT 48.755 -59.548 48.845 -58.54 ;
      RECT 48.705 -58.945 48.845 -58.775 ;
      RECT 48.755 -57.74 48.845 -56.732 ;
      RECT 48.705 -57.505 48.845 -57.335 ;
      RECT 48.755 -56.318 48.845 -55.31 ;
      RECT 48.705 -55.715 48.845 -55.545 ;
      RECT 48.755 -54.51 48.845 -53.502 ;
      RECT 48.705 -54.275 48.845 -54.105 ;
      RECT 48.755 -53.088 48.845 -52.08 ;
      RECT 48.705 -52.485 48.845 -52.315 ;
      RECT 48.755 -51.28 48.845 -50.272 ;
      RECT 48.705 -51.045 48.845 -50.875 ;
      RECT 48.755 -49.858 48.845 -48.85 ;
      RECT 48.705 -49.255 48.845 -49.085 ;
      RECT 48.755 -48.05 48.845 -47.042 ;
      RECT 48.705 -47.815 48.845 -47.645 ;
      RECT 48.755 -46.628 48.845 -45.62 ;
      RECT 48.705 -46.025 48.845 -45.855 ;
      RECT 48.755 -44.82 48.845 -43.812 ;
      RECT 48.705 -44.585 48.845 -44.415 ;
      RECT 48.755 -43.398 48.845 -42.39 ;
      RECT 48.705 -42.795 48.845 -42.625 ;
      RECT 48.755 -41.59 48.845 -40.582 ;
      RECT 48.705 -41.355 48.845 -41.185 ;
      RECT 48.755 -40.168 48.845 -39.16 ;
      RECT 48.705 -39.565 48.845 -39.395 ;
      RECT 48.755 -38.36 48.845 -37.352 ;
      RECT 48.705 -38.125 48.845 -37.955 ;
      RECT 48.755 -36.938 48.845 -35.93 ;
      RECT 48.705 -36.335 48.845 -36.165 ;
      RECT 48.755 -35.13 48.845 -34.122 ;
      RECT 48.705 -34.895 48.845 -34.725 ;
      RECT 48.755 -33.708 48.845 -32.7 ;
      RECT 48.705 -33.105 48.845 -32.935 ;
      RECT 48.755 -31.9 48.845 -30.892 ;
      RECT 48.705 -31.665 48.845 -31.495 ;
      RECT 48.755 -30.478 48.845 -29.47 ;
      RECT 48.705 -29.875 48.845 -29.705 ;
      RECT 48.755 -28.67 48.845 -27.662 ;
      RECT 48.705 -28.435 48.845 -28.265 ;
      RECT 48.755 -27.248 48.845 -26.24 ;
      RECT 48.705 -26.645 48.845 -26.475 ;
      RECT 48.755 -25.44 48.845 -24.432 ;
      RECT 48.705 -25.205 48.845 -25.035 ;
      RECT 48.755 -24.018 48.845 -23.01 ;
      RECT 48.705 -23.415 48.845 -23.245 ;
      RECT 48.755 -22.21 48.845 -21.202 ;
      RECT 48.705 -21.975 48.845 -21.805 ;
      RECT 48.755 -20.788 48.845 -19.78 ;
      RECT 48.705 -20.185 48.845 -20.015 ;
      RECT 48.755 -18.98 48.845 -17.972 ;
      RECT 48.705 -18.745 48.845 -18.575 ;
      RECT 48.755 -17.558 48.845 -16.55 ;
      RECT 48.705 -16.955 48.845 -16.785 ;
      RECT 48.755 -15.75 48.845 -14.742 ;
      RECT 48.705 -15.515 48.845 -15.345 ;
      RECT 48.755 -14.328 48.845 -13.32 ;
      RECT 48.705 -13.725 48.845 -13.555 ;
      RECT 48.755 -12.52 48.845 -11.512 ;
      RECT 48.705 -12.285 48.845 -12.115 ;
      RECT 48.755 -11.098 48.845 -10.09 ;
      RECT 48.705 -10.495 48.845 -10.325 ;
      RECT 48.755 -9.29 48.845 -8.282 ;
      RECT 48.705 -9.055 48.845 -8.885 ;
      RECT 48.755 -7.868 48.845 -6.86 ;
      RECT 48.705 -7.265 48.845 -7.095 ;
      RECT 48.755 -6.06 48.845 -5.052 ;
      RECT 48.705 -5.825 48.845 -5.655 ;
      RECT 48.755 -4.638 48.845 -3.63 ;
      RECT 48.705 -4.035 48.845 -3.865 ;
      RECT 48.755 -2.83 48.845 -1.822 ;
      RECT 48.705 -2.595 48.845 -2.425 ;
      RECT 48.755 -1.408 48.845 -0.4 ;
      RECT 48.705 -0.805 48.845 -0.635 ;
      RECT 48.755 0.4 48.845 1.408 ;
      RECT 48.705 0.635 48.845 0.805 ;
      RECT 48.355 -101.538 48.445 -100.531 ;
      RECT 48.355 -101.225 48.495 -101.055 ;
      RECT 48.355 -99.729 48.445 -98.722 ;
      RECT 48.355 -99.205 48.495 -99.035 ;
      RECT 48.355 -98.308 48.445 -97.301 ;
      RECT 48.355 -97.995 48.495 -97.825 ;
      RECT 48.355 -96.499 48.445 -95.492 ;
      RECT 48.355 -95.975 48.495 -95.805 ;
      RECT 48.355 -95.078 48.445 -94.071 ;
      RECT 48.355 -94.765 48.495 -94.595 ;
      RECT 48.355 -93.269 48.445 -92.262 ;
      RECT 48.355 -92.745 48.495 -92.575 ;
      RECT 48.355 -91.848 48.445 -90.841 ;
      RECT 48.355 -91.535 48.495 -91.365 ;
      RECT 48.355 -90.039 48.445 -89.032 ;
      RECT 48.355 -89.515 48.495 -89.345 ;
      RECT 48.355 -88.618 48.445 -87.611 ;
      RECT 48.355 -88.305 48.495 -88.135 ;
      RECT 48.355 -86.809 48.445 -85.802 ;
      RECT 48.355 -86.285 48.495 -86.115 ;
      RECT 48.355 -85.388 48.445 -84.381 ;
      RECT 48.355 -85.075 48.495 -84.905 ;
      RECT 48.355 -83.579 48.445 -82.572 ;
      RECT 48.355 -83.055 48.495 -82.885 ;
      RECT 48.355 -82.158 48.445 -81.151 ;
      RECT 48.355 -81.845 48.495 -81.675 ;
      RECT 48.355 -80.349 48.445 -79.342 ;
      RECT 48.355 -79.825 48.495 -79.655 ;
      RECT 48.355 -78.928 48.445 -77.921 ;
      RECT 48.355 -78.615 48.495 -78.445 ;
      RECT 48.355 -77.119 48.445 -76.112 ;
      RECT 48.355 -76.595 48.495 -76.425 ;
      RECT 48.355 -75.698 48.445 -74.691 ;
      RECT 48.355 -75.385 48.495 -75.215 ;
      RECT 48.355 -73.889 48.445 -72.882 ;
      RECT 48.355 -73.365 48.495 -73.195 ;
      RECT 48.355 -72.468 48.445 -71.461 ;
      RECT 48.355 -72.155 48.495 -71.985 ;
      RECT 48.355 -70.659 48.445 -69.652 ;
      RECT 48.355 -70.135 48.495 -69.965 ;
      RECT 48.355 -69.238 48.445 -68.231 ;
      RECT 48.355 -68.925 48.495 -68.755 ;
      RECT 48.355 -67.429 48.445 -66.422 ;
      RECT 48.355 -66.905 48.495 -66.735 ;
      RECT 48.355 -66.008 48.445 -65.001 ;
      RECT 48.355 -65.695 48.495 -65.525 ;
      RECT 48.355 -64.199 48.445 -63.192 ;
      RECT 48.355 -63.675 48.495 -63.505 ;
      RECT 48.355 -62.778 48.445 -61.771 ;
      RECT 48.355 -62.465 48.495 -62.295 ;
      RECT 48.355 -60.969 48.445 -59.962 ;
      RECT 48.355 -60.445 48.495 -60.275 ;
      RECT 48.355 -59.548 48.445 -58.541 ;
      RECT 48.355 -59.235 48.495 -59.065 ;
      RECT 48.355 -57.739 48.445 -56.732 ;
      RECT 48.355 -57.215 48.495 -57.045 ;
      RECT 48.355 -56.318 48.445 -55.311 ;
      RECT 48.355 -56.005 48.495 -55.835 ;
      RECT 48.355 -54.509 48.445 -53.502 ;
      RECT 48.355 -53.985 48.495 -53.815 ;
      RECT 48.355 -53.088 48.445 -52.081 ;
      RECT 48.355 -52.775 48.495 -52.605 ;
      RECT 48.355 -51.279 48.445 -50.272 ;
      RECT 48.355 -50.755 48.495 -50.585 ;
      RECT 48.355 -49.858 48.445 -48.851 ;
      RECT 48.355 -49.545 48.495 -49.375 ;
      RECT 48.355 -48.049 48.445 -47.042 ;
      RECT 48.355 -47.525 48.495 -47.355 ;
      RECT 48.355 -46.628 48.445 -45.621 ;
      RECT 48.355 -46.315 48.495 -46.145 ;
      RECT 48.355 -44.819 48.445 -43.812 ;
      RECT 48.355 -44.295 48.495 -44.125 ;
      RECT 48.355 -43.398 48.445 -42.391 ;
      RECT 48.355 -43.085 48.495 -42.915 ;
      RECT 48.355 -41.589 48.445 -40.582 ;
      RECT 48.355 -41.065 48.495 -40.895 ;
      RECT 48.355 -40.168 48.445 -39.161 ;
      RECT 48.355 -39.855 48.495 -39.685 ;
      RECT 48.355 -38.359 48.445 -37.352 ;
      RECT 48.355 -37.835 48.495 -37.665 ;
      RECT 48.355 -36.938 48.445 -35.931 ;
      RECT 48.355 -36.625 48.495 -36.455 ;
      RECT 48.355 -35.129 48.445 -34.122 ;
      RECT 48.355 -34.605 48.495 -34.435 ;
      RECT 48.355 -33.708 48.445 -32.701 ;
      RECT 48.355 -33.395 48.495 -33.225 ;
      RECT 48.355 -31.899 48.445 -30.892 ;
      RECT 48.355 -31.375 48.495 -31.205 ;
      RECT 48.355 -30.478 48.445 -29.471 ;
      RECT 48.355 -30.165 48.495 -29.995 ;
      RECT 48.355 -28.669 48.445 -27.662 ;
      RECT 48.355 -28.145 48.495 -27.975 ;
      RECT 48.355 -27.248 48.445 -26.241 ;
      RECT 48.355 -26.935 48.495 -26.765 ;
      RECT 48.355 -25.439 48.445 -24.432 ;
      RECT 48.355 -24.915 48.495 -24.745 ;
      RECT 48.355 -24.018 48.445 -23.011 ;
      RECT 48.355 -23.705 48.495 -23.535 ;
      RECT 48.355 -22.209 48.445 -21.202 ;
      RECT 48.355 -21.685 48.495 -21.515 ;
      RECT 48.355 -20.788 48.445 -19.781 ;
      RECT 48.355 -20.475 48.495 -20.305 ;
      RECT 48.355 -18.979 48.445 -17.972 ;
      RECT 48.355 -18.455 48.495 -18.285 ;
      RECT 48.355 -17.558 48.445 -16.551 ;
      RECT 48.355 -17.245 48.495 -17.075 ;
      RECT 48.355 -15.749 48.445 -14.742 ;
      RECT 48.355 -15.225 48.495 -15.055 ;
      RECT 48.355 -14.328 48.445 -13.321 ;
      RECT 48.355 -14.015 48.495 -13.845 ;
      RECT 48.355 -12.519 48.445 -11.512 ;
      RECT 48.355 -11.995 48.495 -11.825 ;
      RECT 48.355 -11.098 48.445 -10.091 ;
      RECT 48.355 -10.785 48.495 -10.615 ;
      RECT 48.355 -9.289 48.445 -8.282 ;
      RECT 48.355 -8.765 48.495 -8.595 ;
      RECT 48.355 -7.868 48.445 -6.861 ;
      RECT 48.355 -7.555 48.495 -7.385 ;
      RECT 48.355 -6.059 48.445 -5.052 ;
      RECT 48.355 -5.535 48.495 -5.365 ;
      RECT 48.355 -4.638 48.445 -3.631 ;
      RECT 48.355 -4.325 48.495 -4.155 ;
      RECT 48.355 -2.829 48.445 -1.822 ;
      RECT 48.355 -2.305 48.495 -2.135 ;
      RECT 48.355 -1.408 48.445 -0.401 ;
      RECT 48.355 -1.095 48.495 -0.925 ;
      RECT 48.355 0.401 48.445 1.408 ;
      RECT 48.355 0.925 48.495 1.095 ;
      RECT 44.185 -108.935 47.965 -108.815 ;
      RECT 45.505 -109.475 45.605 -108.815 ;
      RECT 44.945 -109.475 45.045 -108.815 ;
      RECT 44.385 -109.475 44.485 -108.815 ;
      RECT 47.555 -101.538 47.645 -100.53 ;
      RECT 47.505 -100.935 47.645 -100.765 ;
      RECT 47.555 -99.73 47.645 -98.722 ;
      RECT 47.505 -99.495 47.645 -99.325 ;
      RECT 47.555 -98.308 47.645 -97.3 ;
      RECT 47.505 -97.705 47.645 -97.535 ;
      RECT 47.555 -96.5 47.645 -95.492 ;
      RECT 47.505 -96.265 47.645 -96.095 ;
      RECT 47.555 -95.078 47.645 -94.07 ;
      RECT 47.505 -94.475 47.645 -94.305 ;
      RECT 47.555 -93.27 47.645 -92.262 ;
      RECT 47.505 -93.035 47.645 -92.865 ;
      RECT 47.555 -91.848 47.645 -90.84 ;
      RECT 47.505 -91.245 47.645 -91.075 ;
      RECT 47.555 -90.04 47.645 -89.032 ;
      RECT 47.505 -89.805 47.645 -89.635 ;
      RECT 47.555 -88.618 47.645 -87.61 ;
      RECT 47.505 -88.015 47.645 -87.845 ;
      RECT 47.555 -86.81 47.645 -85.802 ;
      RECT 47.505 -86.575 47.645 -86.405 ;
      RECT 47.555 -85.388 47.645 -84.38 ;
      RECT 47.505 -84.785 47.645 -84.615 ;
      RECT 47.555 -83.58 47.645 -82.572 ;
      RECT 47.505 -83.345 47.645 -83.175 ;
      RECT 47.555 -82.158 47.645 -81.15 ;
      RECT 47.505 -81.555 47.645 -81.385 ;
      RECT 47.555 -80.35 47.645 -79.342 ;
      RECT 47.505 -80.115 47.645 -79.945 ;
      RECT 47.555 -78.928 47.645 -77.92 ;
      RECT 47.505 -78.325 47.645 -78.155 ;
      RECT 47.555 -77.12 47.645 -76.112 ;
      RECT 47.505 -76.885 47.645 -76.715 ;
      RECT 47.555 -75.698 47.645 -74.69 ;
      RECT 47.505 -75.095 47.645 -74.925 ;
      RECT 47.555 -73.89 47.645 -72.882 ;
      RECT 47.505 -73.655 47.645 -73.485 ;
      RECT 47.555 -72.468 47.645 -71.46 ;
      RECT 47.505 -71.865 47.645 -71.695 ;
      RECT 47.555 -70.66 47.645 -69.652 ;
      RECT 47.505 -70.425 47.645 -70.255 ;
      RECT 47.555 -69.238 47.645 -68.23 ;
      RECT 47.505 -68.635 47.645 -68.465 ;
      RECT 47.555 -67.43 47.645 -66.422 ;
      RECT 47.505 -67.195 47.645 -67.025 ;
      RECT 47.555 -66.008 47.645 -65 ;
      RECT 47.505 -65.405 47.645 -65.235 ;
      RECT 47.555 -64.2 47.645 -63.192 ;
      RECT 47.505 -63.965 47.645 -63.795 ;
      RECT 47.555 -62.778 47.645 -61.77 ;
      RECT 47.505 -62.175 47.645 -62.005 ;
      RECT 47.555 -60.97 47.645 -59.962 ;
      RECT 47.505 -60.735 47.645 -60.565 ;
      RECT 47.555 -59.548 47.645 -58.54 ;
      RECT 47.505 -58.945 47.645 -58.775 ;
      RECT 47.555 -57.74 47.645 -56.732 ;
      RECT 47.505 -57.505 47.645 -57.335 ;
      RECT 47.555 -56.318 47.645 -55.31 ;
      RECT 47.505 -55.715 47.645 -55.545 ;
      RECT 47.555 -54.51 47.645 -53.502 ;
      RECT 47.505 -54.275 47.645 -54.105 ;
      RECT 47.555 -53.088 47.645 -52.08 ;
      RECT 47.505 -52.485 47.645 -52.315 ;
      RECT 47.555 -51.28 47.645 -50.272 ;
      RECT 47.505 -51.045 47.645 -50.875 ;
      RECT 47.555 -49.858 47.645 -48.85 ;
      RECT 47.505 -49.255 47.645 -49.085 ;
      RECT 47.555 -48.05 47.645 -47.042 ;
      RECT 47.505 -47.815 47.645 -47.645 ;
      RECT 47.555 -46.628 47.645 -45.62 ;
      RECT 47.505 -46.025 47.645 -45.855 ;
      RECT 47.555 -44.82 47.645 -43.812 ;
      RECT 47.505 -44.585 47.645 -44.415 ;
      RECT 47.555 -43.398 47.645 -42.39 ;
      RECT 47.505 -42.795 47.645 -42.625 ;
      RECT 47.555 -41.59 47.645 -40.582 ;
      RECT 47.505 -41.355 47.645 -41.185 ;
      RECT 47.555 -40.168 47.645 -39.16 ;
      RECT 47.505 -39.565 47.645 -39.395 ;
      RECT 47.555 -38.36 47.645 -37.352 ;
      RECT 47.505 -38.125 47.645 -37.955 ;
      RECT 47.555 -36.938 47.645 -35.93 ;
      RECT 47.505 -36.335 47.645 -36.165 ;
      RECT 47.555 -35.13 47.645 -34.122 ;
      RECT 47.505 -34.895 47.645 -34.725 ;
      RECT 47.555 -33.708 47.645 -32.7 ;
      RECT 47.505 -33.105 47.645 -32.935 ;
      RECT 47.555 -31.9 47.645 -30.892 ;
      RECT 47.505 -31.665 47.645 -31.495 ;
      RECT 47.555 -30.478 47.645 -29.47 ;
      RECT 47.505 -29.875 47.645 -29.705 ;
      RECT 47.555 -28.67 47.645 -27.662 ;
      RECT 47.505 -28.435 47.645 -28.265 ;
      RECT 47.555 -27.248 47.645 -26.24 ;
      RECT 47.505 -26.645 47.645 -26.475 ;
      RECT 47.555 -25.44 47.645 -24.432 ;
      RECT 47.505 -25.205 47.645 -25.035 ;
      RECT 47.555 -24.018 47.645 -23.01 ;
      RECT 47.505 -23.415 47.645 -23.245 ;
      RECT 47.555 -22.21 47.645 -21.202 ;
      RECT 47.505 -21.975 47.645 -21.805 ;
      RECT 47.555 -20.788 47.645 -19.78 ;
      RECT 47.505 -20.185 47.645 -20.015 ;
      RECT 47.555 -18.98 47.645 -17.972 ;
      RECT 47.505 -18.745 47.645 -18.575 ;
      RECT 47.555 -17.558 47.645 -16.55 ;
      RECT 47.505 -16.955 47.645 -16.785 ;
      RECT 47.555 -15.75 47.645 -14.742 ;
      RECT 47.505 -15.515 47.645 -15.345 ;
      RECT 47.555 -14.328 47.645 -13.32 ;
      RECT 47.505 -13.725 47.645 -13.555 ;
      RECT 47.555 -12.52 47.645 -11.512 ;
      RECT 47.505 -12.285 47.645 -12.115 ;
      RECT 47.555 -11.098 47.645 -10.09 ;
      RECT 47.505 -10.495 47.645 -10.325 ;
      RECT 47.555 -9.29 47.645 -8.282 ;
      RECT 47.505 -9.055 47.645 -8.885 ;
      RECT 47.555 -7.868 47.645 -6.86 ;
      RECT 47.505 -7.265 47.645 -7.095 ;
      RECT 47.555 -6.06 47.645 -5.052 ;
      RECT 47.505 -5.825 47.645 -5.655 ;
      RECT 47.555 -4.638 47.645 -3.63 ;
      RECT 47.505 -4.035 47.645 -3.865 ;
      RECT 47.555 -2.83 47.645 -1.822 ;
      RECT 47.505 -2.595 47.645 -2.425 ;
      RECT 47.555 -1.408 47.645 -0.4 ;
      RECT 47.505 -0.805 47.645 -0.635 ;
      RECT 47.555 0.4 47.645 1.408 ;
      RECT 47.505 0.635 47.645 0.805 ;
      RECT 46.125 -111.685 47.605 -111.585 ;
      RECT 46.125 -112.195 46.225 -111.585 ;
      RECT 46.345 -109.15 47.605 -109.05 ;
      RECT 47.505 -109.475 47.605 -109.05 ;
      RECT 46.945 -109.475 47.045 -109.05 ;
      RECT 46.385 -109.475 46.485 -109.05 ;
      RECT 47.155 -101.538 47.245 -100.531 ;
      RECT 47.155 -101.225 47.295 -101.055 ;
      RECT 47.155 -99.729 47.245 -98.722 ;
      RECT 47.155 -99.205 47.295 -99.035 ;
      RECT 47.155 -98.308 47.245 -97.301 ;
      RECT 47.155 -97.995 47.295 -97.825 ;
      RECT 47.155 -96.499 47.245 -95.492 ;
      RECT 47.155 -95.975 47.295 -95.805 ;
      RECT 47.155 -95.078 47.245 -94.071 ;
      RECT 47.155 -94.765 47.295 -94.595 ;
      RECT 47.155 -93.269 47.245 -92.262 ;
      RECT 47.155 -92.745 47.295 -92.575 ;
      RECT 47.155 -91.848 47.245 -90.841 ;
      RECT 47.155 -91.535 47.295 -91.365 ;
      RECT 47.155 -90.039 47.245 -89.032 ;
      RECT 47.155 -89.515 47.295 -89.345 ;
      RECT 47.155 -88.618 47.245 -87.611 ;
      RECT 47.155 -88.305 47.295 -88.135 ;
      RECT 47.155 -86.809 47.245 -85.802 ;
      RECT 47.155 -86.285 47.295 -86.115 ;
      RECT 47.155 -85.388 47.245 -84.381 ;
      RECT 47.155 -85.075 47.295 -84.905 ;
      RECT 47.155 -83.579 47.245 -82.572 ;
      RECT 47.155 -83.055 47.295 -82.885 ;
      RECT 47.155 -82.158 47.245 -81.151 ;
      RECT 47.155 -81.845 47.295 -81.675 ;
      RECT 47.155 -80.349 47.245 -79.342 ;
      RECT 47.155 -79.825 47.295 -79.655 ;
      RECT 47.155 -78.928 47.245 -77.921 ;
      RECT 47.155 -78.615 47.295 -78.445 ;
      RECT 47.155 -77.119 47.245 -76.112 ;
      RECT 47.155 -76.595 47.295 -76.425 ;
      RECT 47.155 -75.698 47.245 -74.691 ;
      RECT 47.155 -75.385 47.295 -75.215 ;
      RECT 47.155 -73.889 47.245 -72.882 ;
      RECT 47.155 -73.365 47.295 -73.195 ;
      RECT 47.155 -72.468 47.245 -71.461 ;
      RECT 47.155 -72.155 47.295 -71.985 ;
      RECT 47.155 -70.659 47.245 -69.652 ;
      RECT 47.155 -70.135 47.295 -69.965 ;
      RECT 47.155 -69.238 47.245 -68.231 ;
      RECT 47.155 -68.925 47.295 -68.755 ;
      RECT 47.155 -67.429 47.245 -66.422 ;
      RECT 47.155 -66.905 47.295 -66.735 ;
      RECT 47.155 -66.008 47.245 -65.001 ;
      RECT 47.155 -65.695 47.295 -65.525 ;
      RECT 47.155 -64.199 47.245 -63.192 ;
      RECT 47.155 -63.675 47.295 -63.505 ;
      RECT 47.155 -62.778 47.245 -61.771 ;
      RECT 47.155 -62.465 47.295 -62.295 ;
      RECT 47.155 -60.969 47.245 -59.962 ;
      RECT 47.155 -60.445 47.295 -60.275 ;
      RECT 47.155 -59.548 47.245 -58.541 ;
      RECT 47.155 -59.235 47.295 -59.065 ;
      RECT 47.155 -57.739 47.245 -56.732 ;
      RECT 47.155 -57.215 47.295 -57.045 ;
      RECT 47.155 -56.318 47.245 -55.311 ;
      RECT 47.155 -56.005 47.295 -55.835 ;
      RECT 47.155 -54.509 47.245 -53.502 ;
      RECT 47.155 -53.985 47.295 -53.815 ;
      RECT 47.155 -53.088 47.245 -52.081 ;
      RECT 47.155 -52.775 47.295 -52.605 ;
      RECT 47.155 -51.279 47.245 -50.272 ;
      RECT 47.155 -50.755 47.295 -50.585 ;
      RECT 47.155 -49.858 47.245 -48.851 ;
      RECT 47.155 -49.545 47.295 -49.375 ;
      RECT 47.155 -48.049 47.245 -47.042 ;
      RECT 47.155 -47.525 47.295 -47.355 ;
      RECT 47.155 -46.628 47.245 -45.621 ;
      RECT 47.155 -46.315 47.295 -46.145 ;
      RECT 47.155 -44.819 47.245 -43.812 ;
      RECT 47.155 -44.295 47.295 -44.125 ;
      RECT 47.155 -43.398 47.245 -42.391 ;
      RECT 47.155 -43.085 47.295 -42.915 ;
      RECT 47.155 -41.589 47.245 -40.582 ;
      RECT 47.155 -41.065 47.295 -40.895 ;
      RECT 47.155 -40.168 47.245 -39.161 ;
      RECT 47.155 -39.855 47.295 -39.685 ;
      RECT 47.155 -38.359 47.245 -37.352 ;
      RECT 47.155 -37.835 47.295 -37.665 ;
      RECT 47.155 -36.938 47.245 -35.931 ;
      RECT 47.155 -36.625 47.295 -36.455 ;
      RECT 47.155 -35.129 47.245 -34.122 ;
      RECT 47.155 -34.605 47.295 -34.435 ;
      RECT 47.155 -33.708 47.245 -32.701 ;
      RECT 47.155 -33.395 47.295 -33.225 ;
      RECT 47.155 -31.899 47.245 -30.892 ;
      RECT 47.155 -31.375 47.295 -31.205 ;
      RECT 47.155 -30.478 47.245 -29.471 ;
      RECT 47.155 -30.165 47.295 -29.995 ;
      RECT 47.155 -28.669 47.245 -27.662 ;
      RECT 47.155 -28.145 47.295 -27.975 ;
      RECT 47.155 -27.248 47.245 -26.241 ;
      RECT 47.155 -26.935 47.295 -26.765 ;
      RECT 47.155 -25.439 47.245 -24.432 ;
      RECT 47.155 -24.915 47.295 -24.745 ;
      RECT 47.155 -24.018 47.245 -23.011 ;
      RECT 47.155 -23.705 47.295 -23.535 ;
      RECT 47.155 -22.209 47.245 -21.202 ;
      RECT 47.155 -21.685 47.295 -21.515 ;
      RECT 47.155 -20.788 47.245 -19.781 ;
      RECT 47.155 -20.475 47.295 -20.305 ;
      RECT 47.155 -18.979 47.245 -17.972 ;
      RECT 47.155 -18.455 47.295 -18.285 ;
      RECT 47.155 -17.558 47.245 -16.551 ;
      RECT 47.155 -17.245 47.295 -17.075 ;
      RECT 47.155 -15.749 47.245 -14.742 ;
      RECT 47.155 -15.225 47.295 -15.055 ;
      RECT 47.155 -14.328 47.245 -13.321 ;
      RECT 47.155 -14.015 47.295 -13.845 ;
      RECT 47.155 -12.519 47.245 -11.512 ;
      RECT 47.155 -11.995 47.295 -11.825 ;
      RECT 47.155 -11.098 47.245 -10.091 ;
      RECT 47.155 -10.785 47.295 -10.615 ;
      RECT 47.155 -9.289 47.245 -8.282 ;
      RECT 47.155 -8.765 47.295 -8.595 ;
      RECT 47.155 -7.868 47.245 -6.861 ;
      RECT 47.155 -7.555 47.295 -7.385 ;
      RECT 47.155 -6.059 47.245 -5.052 ;
      RECT 47.155 -5.535 47.295 -5.365 ;
      RECT 47.155 -4.638 47.245 -3.631 ;
      RECT 47.155 -4.325 47.295 -4.155 ;
      RECT 47.155 -2.829 47.245 -1.822 ;
      RECT 47.155 -2.305 47.295 -2.135 ;
      RECT 47.155 -1.408 47.245 -0.401 ;
      RECT 47.155 -1.095 47.295 -0.925 ;
      RECT 47.155 0.401 47.245 1.408 ;
      RECT 47.155 0.925 47.295 1.095 ;
      RECT 46.485 -111.495 46.655 -111.385 ;
      RECT 43.335 -111.495 46.655 -111.395 ;
      RECT 46.355 -101.538 46.445 -100.53 ;
      RECT 46.305 -100.935 46.445 -100.765 ;
      RECT 46.355 -99.73 46.445 -98.722 ;
      RECT 46.305 -99.495 46.445 -99.325 ;
      RECT 46.355 -98.308 46.445 -97.3 ;
      RECT 46.305 -97.705 46.445 -97.535 ;
      RECT 46.355 -96.5 46.445 -95.492 ;
      RECT 46.305 -96.265 46.445 -96.095 ;
      RECT 46.355 -95.078 46.445 -94.07 ;
      RECT 46.305 -94.475 46.445 -94.305 ;
      RECT 46.355 -93.27 46.445 -92.262 ;
      RECT 46.305 -93.035 46.445 -92.865 ;
      RECT 46.355 -91.848 46.445 -90.84 ;
      RECT 46.305 -91.245 46.445 -91.075 ;
      RECT 46.355 -90.04 46.445 -89.032 ;
      RECT 46.305 -89.805 46.445 -89.635 ;
      RECT 46.355 -88.618 46.445 -87.61 ;
      RECT 46.305 -88.015 46.445 -87.845 ;
      RECT 46.355 -86.81 46.445 -85.802 ;
      RECT 46.305 -86.575 46.445 -86.405 ;
      RECT 46.355 -85.388 46.445 -84.38 ;
      RECT 46.305 -84.785 46.445 -84.615 ;
      RECT 46.355 -83.58 46.445 -82.572 ;
      RECT 46.305 -83.345 46.445 -83.175 ;
      RECT 46.355 -82.158 46.445 -81.15 ;
      RECT 46.305 -81.555 46.445 -81.385 ;
      RECT 46.355 -80.35 46.445 -79.342 ;
      RECT 46.305 -80.115 46.445 -79.945 ;
      RECT 46.355 -78.928 46.445 -77.92 ;
      RECT 46.305 -78.325 46.445 -78.155 ;
      RECT 46.355 -77.12 46.445 -76.112 ;
      RECT 46.305 -76.885 46.445 -76.715 ;
      RECT 46.355 -75.698 46.445 -74.69 ;
      RECT 46.305 -75.095 46.445 -74.925 ;
      RECT 46.355 -73.89 46.445 -72.882 ;
      RECT 46.305 -73.655 46.445 -73.485 ;
      RECT 46.355 -72.468 46.445 -71.46 ;
      RECT 46.305 -71.865 46.445 -71.695 ;
      RECT 46.355 -70.66 46.445 -69.652 ;
      RECT 46.305 -70.425 46.445 -70.255 ;
      RECT 46.355 -69.238 46.445 -68.23 ;
      RECT 46.305 -68.635 46.445 -68.465 ;
      RECT 46.355 -67.43 46.445 -66.422 ;
      RECT 46.305 -67.195 46.445 -67.025 ;
      RECT 46.355 -66.008 46.445 -65 ;
      RECT 46.305 -65.405 46.445 -65.235 ;
      RECT 46.355 -64.2 46.445 -63.192 ;
      RECT 46.305 -63.965 46.445 -63.795 ;
      RECT 46.355 -62.778 46.445 -61.77 ;
      RECT 46.305 -62.175 46.445 -62.005 ;
      RECT 46.355 -60.97 46.445 -59.962 ;
      RECT 46.305 -60.735 46.445 -60.565 ;
      RECT 46.355 -59.548 46.445 -58.54 ;
      RECT 46.305 -58.945 46.445 -58.775 ;
      RECT 46.355 -57.74 46.445 -56.732 ;
      RECT 46.305 -57.505 46.445 -57.335 ;
      RECT 46.355 -56.318 46.445 -55.31 ;
      RECT 46.305 -55.715 46.445 -55.545 ;
      RECT 46.355 -54.51 46.445 -53.502 ;
      RECT 46.305 -54.275 46.445 -54.105 ;
      RECT 46.355 -53.088 46.445 -52.08 ;
      RECT 46.305 -52.485 46.445 -52.315 ;
      RECT 46.355 -51.28 46.445 -50.272 ;
      RECT 46.305 -51.045 46.445 -50.875 ;
      RECT 46.355 -49.858 46.445 -48.85 ;
      RECT 46.305 -49.255 46.445 -49.085 ;
      RECT 46.355 -48.05 46.445 -47.042 ;
      RECT 46.305 -47.815 46.445 -47.645 ;
      RECT 46.355 -46.628 46.445 -45.62 ;
      RECT 46.305 -46.025 46.445 -45.855 ;
      RECT 46.355 -44.82 46.445 -43.812 ;
      RECT 46.305 -44.585 46.445 -44.415 ;
      RECT 46.355 -43.398 46.445 -42.39 ;
      RECT 46.305 -42.795 46.445 -42.625 ;
      RECT 46.355 -41.59 46.445 -40.582 ;
      RECT 46.305 -41.355 46.445 -41.185 ;
      RECT 46.355 -40.168 46.445 -39.16 ;
      RECT 46.305 -39.565 46.445 -39.395 ;
      RECT 46.355 -38.36 46.445 -37.352 ;
      RECT 46.305 -38.125 46.445 -37.955 ;
      RECT 46.355 -36.938 46.445 -35.93 ;
      RECT 46.305 -36.335 46.445 -36.165 ;
      RECT 46.355 -35.13 46.445 -34.122 ;
      RECT 46.305 -34.895 46.445 -34.725 ;
      RECT 46.355 -33.708 46.445 -32.7 ;
      RECT 46.305 -33.105 46.445 -32.935 ;
      RECT 46.355 -31.9 46.445 -30.892 ;
      RECT 46.305 -31.665 46.445 -31.495 ;
      RECT 46.355 -30.478 46.445 -29.47 ;
      RECT 46.305 -29.875 46.445 -29.705 ;
      RECT 46.355 -28.67 46.445 -27.662 ;
      RECT 46.305 -28.435 46.445 -28.265 ;
      RECT 46.355 -27.248 46.445 -26.24 ;
      RECT 46.305 -26.645 46.445 -26.475 ;
      RECT 46.355 -25.44 46.445 -24.432 ;
      RECT 46.305 -25.205 46.445 -25.035 ;
      RECT 46.355 -24.018 46.445 -23.01 ;
      RECT 46.305 -23.415 46.445 -23.245 ;
      RECT 46.355 -22.21 46.445 -21.202 ;
      RECT 46.305 -21.975 46.445 -21.805 ;
      RECT 46.355 -20.788 46.445 -19.78 ;
      RECT 46.305 -20.185 46.445 -20.015 ;
      RECT 46.355 -18.98 46.445 -17.972 ;
      RECT 46.305 -18.745 46.445 -18.575 ;
      RECT 46.355 -17.558 46.445 -16.55 ;
      RECT 46.305 -16.955 46.445 -16.785 ;
      RECT 46.355 -15.75 46.445 -14.742 ;
      RECT 46.305 -15.515 46.445 -15.345 ;
      RECT 46.355 -14.328 46.445 -13.32 ;
      RECT 46.305 -13.725 46.445 -13.555 ;
      RECT 46.355 -12.52 46.445 -11.512 ;
      RECT 46.305 -12.285 46.445 -12.115 ;
      RECT 46.355 -11.098 46.445 -10.09 ;
      RECT 46.305 -10.495 46.445 -10.325 ;
      RECT 46.355 -9.29 46.445 -8.282 ;
      RECT 46.305 -9.055 46.445 -8.885 ;
      RECT 46.355 -7.868 46.445 -6.86 ;
      RECT 46.305 -7.265 46.445 -7.095 ;
      RECT 46.355 -6.06 46.445 -5.052 ;
      RECT 46.305 -5.825 46.445 -5.655 ;
      RECT 46.355 -4.638 46.445 -3.63 ;
      RECT 46.305 -4.035 46.445 -3.865 ;
      RECT 46.355 -2.83 46.445 -1.822 ;
      RECT 46.305 -2.595 46.445 -2.425 ;
      RECT 46.355 -1.408 46.445 -0.4 ;
      RECT 46.305 -0.805 46.445 -0.635 ;
      RECT 46.355 0.4 46.445 1.408 ;
      RECT 46.305 0.635 46.445 0.805 ;
      RECT 45.955 -101.538 46.045 -100.531 ;
      RECT 45.955 -101.225 46.095 -101.055 ;
      RECT 45.955 -99.729 46.045 -98.722 ;
      RECT 45.955 -99.205 46.095 -99.035 ;
      RECT 45.955 -98.308 46.045 -97.301 ;
      RECT 45.955 -97.995 46.095 -97.825 ;
      RECT 45.955 -96.499 46.045 -95.492 ;
      RECT 45.955 -95.975 46.095 -95.805 ;
      RECT 45.955 -95.078 46.045 -94.071 ;
      RECT 45.955 -94.765 46.095 -94.595 ;
      RECT 45.955 -93.269 46.045 -92.262 ;
      RECT 45.955 -92.745 46.095 -92.575 ;
      RECT 45.955 -91.848 46.045 -90.841 ;
      RECT 45.955 -91.535 46.095 -91.365 ;
      RECT 45.955 -90.039 46.045 -89.032 ;
      RECT 45.955 -89.515 46.095 -89.345 ;
      RECT 45.955 -88.618 46.045 -87.611 ;
      RECT 45.955 -88.305 46.095 -88.135 ;
      RECT 45.955 -86.809 46.045 -85.802 ;
      RECT 45.955 -86.285 46.095 -86.115 ;
      RECT 45.955 -85.388 46.045 -84.381 ;
      RECT 45.955 -85.075 46.095 -84.905 ;
      RECT 45.955 -83.579 46.045 -82.572 ;
      RECT 45.955 -83.055 46.095 -82.885 ;
      RECT 45.955 -82.158 46.045 -81.151 ;
      RECT 45.955 -81.845 46.095 -81.675 ;
      RECT 45.955 -80.349 46.045 -79.342 ;
      RECT 45.955 -79.825 46.095 -79.655 ;
      RECT 45.955 -78.928 46.045 -77.921 ;
      RECT 45.955 -78.615 46.095 -78.445 ;
      RECT 45.955 -77.119 46.045 -76.112 ;
      RECT 45.955 -76.595 46.095 -76.425 ;
      RECT 45.955 -75.698 46.045 -74.691 ;
      RECT 45.955 -75.385 46.095 -75.215 ;
      RECT 45.955 -73.889 46.045 -72.882 ;
      RECT 45.955 -73.365 46.095 -73.195 ;
      RECT 45.955 -72.468 46.045 -71.461 ;
      RECT 45.955 -72.155 46.095 -71.985 ;
      RECT 45.955 -70.659 46.045 -69.652 ;
      RECT 45.955 -70.135 46.095 -69.965 ;
      RECT 45.955 -69.238 46.045 -68.231 ;
      RECT 45.955 -68.925 46.095 -68.755 ;
      RECT 45.955 -67.429 46.045 -66.422 ;
      RECT 45.955 -66.905 46.095 -66.735 ;
      RECT 45.955 -66.008 46.045 -65.001 ;
      RECT 45.955 -65.695 46.095 -65.525 ;
      RECT 45.955 -64.199 46.045 -63.192 ;
      RECT 45.955 -63.675 46.095 -63.505 ;
      RECT 45.955 -62.778 46.045 -61.771 ;
      RECT 45.955 -62.465 46.095 -62.295 ;
      RECT 45.955 -60.969 46.045 -59.962 ;
      RECT 45.955 -60.445 46.095 -60.275 ;
      RECT 45.955 -59.548 46.045 -58.541 ;
      RECT 45.955 -59.235 46.095 -59.065 ;
      RECT 45.955 -57.739 46.045 -56.732 ;
      RECT 45.955 -57.215 46.095 -57.045 ;
      RECT 45.955 -56.318 46.045 -55.311 ;
      RECT 45.955 -56.005 46.095 -55.835 ;
      RECT 45.955 -54.509 46.045 -53.502 ;
      RECT 45.955 -53.985 46.095 -53.815 ;
      RECT 45.955 -53.088 46.045 -52.081 ;
      RECT 45.955 -52.775 46.095 -52.605 ;
      RECT 45.955 -51.279 46.045 -50.272 ;
      RECT 45.955 -50.755 46.095 -50.585 ;
      RECT 45.955 -49.858 46.045 -48.851 ;
      RECT 45.955 -49.545 46.095 -49.375 ;
      RECT 45.955 -48.049 46.045 -47.042 ;
      RECT 45.955 -47.525 46.095 -47.355 ;
      RECT 45.955 -46.628 46.045 -45.621 ;
      RECT 45.955 -46.315 46.095 -46.145 ;
      RECT 45.955 -44.819 46.045 -43.812 ;
      RECT 45.955 -44.295 46.095 -44.125 ;
      RECT 45.955 -43.398 46.045 -42.391 ;
      RECT 45.955 -43.085 46.095 -42.915 ;
      RECT 45.955 -41.589 46.045 -40.582 ;
      RECT 45.955 -41.065 46.095 -40.895 ;
      RECT 45.955 -40.168 46.045 -39.161 ;
      RECT 45.955 -39.855 46.095 -39.685 ;
      RECT 45.955 -38.359 46.045 -37.352 ;
      RECT 45.955 -37.835 46.095 -37.665 ;
      RECT 45.955 -36.938 46.045 -35.931 ;
      RECT 45.955 -36.625 46.095 -36.455 ;
      RECT 45.955 -35.129 46.045 -34.122 ;
      RECT 45.955 -34.605 46.095 -34.435 ;
      RECT 45.955 -33.708 46.045 -32.701 ;
      RECT 45.955 -33.395 46.095 -33.225 ;
      RECT 45.955 -31.899 46.045 -30.892 ;
      RECT 45.955 -31.375 46.095 -31.205 ;
      RECT 45.955 -30.478 46.045 -29.471 ;
      RECT 45.955 -30.165 46.095 -29.995 ;
      RECT 45.955 -28.669 46.045 -27.662 ;
      RECT 45.955 -28.145 46.095 -27.975 ;
      RECT 45.955 -27.248 46.045 -26.241 ;
      RECT 45.955 -26.935 46.095 -26.765 ;
      RECT 45.955 -25.439 46.045 -24.432 ;
      RECT 45.955 -24.915 46.095 -24.745 ;
      RECT 45.955 -24.018 46.045 -23.011 ;
      RECT 45.955 -23.705 46.095 -23.535 ;
      RECT 45.955 -22.209 46.045 -21.202 ;
      RECT 45.955 -21.685 46.095 -21.515 ;
      RECT 45.955 -20.788 46.045 -19.781 ;
      RECT 45.955 -20.475 46.095 -20.305 ;
      RECT 45.955 -18.979 46.045 -17.972 ;
      RECT 45.955 -18.455 46.095 -18.285 ;
      RECT 45.955 -17.558 46.045 -16.551 ;
      RECT 45.955 -17.245 46.095 -17.075 ;
      RECT 45.955 -15.749 46.045 -14.742 ;
      RECT 45.955 -15.225 46.095 -15.055 ;
      RECT 45.955 -14.328 46.045 -13.321 ;
      RECT 45.955 -14.015 46.095 -13.845 ;
      RECT 45.955 -12.519 46.045 -11.512 ;
      RECT 45.955 -11.995 46.095 -11.825 ;
      RECT 45.955 -11.098 46.045 -10.091 ;
      RECT 45.955 -10.785 46.095 -10.615 ;
      RECT 45.955 -9.289 46.045 -8.282 ;
      RECT 45.955 -8.765 46.095 -8.595 ;
      RECT 45.955 -7.868 46.045 -6.861 ;
      RECT 45.955 -7.555 46.095 -7.385 ;
      RECT 45.955 -6.059 46.045 -5.052 ;
      RECT 45.955 -5.535 46.095 -5.365 ;
      RECT 45.955 -4.638 46.045 -3.631 ;
      RECT 45.955 -4.325 46.095 -4.155 ;
      RECT 45.955 -2.829 46.045 -1.822 ;
      RECT 45.955 -2.305 46.095 -2.135 ;
      RECT 45.955 -1.408 46.045 -0.401 ;
      RECT 45.955 -1.095 46.095 -0.925 ;
      RECT 45.955 0.401 46.045 1.408 ;
      RECT 45.955 0.925 46.095 1.095 ;
      RECT 44.105 -111.685 45.585 -111.585 ;
      RECT 44.105 -112.055 44.205 -111.585 ;
      RECT 43.91 -114.395 45.485 -114.275 ;
      RECT 45.385 -114.895 45.485 -114.275 ;
      RECT 44.79 -114.895 44.89 -114.275 ;
      RECT 43.91 -114.85 44.01 -114.275 ;
      RECT 45.155 -101.538 45.245 -100.53 ;
      RECT 45.105 -100.935 45.245 -100.765 ;
      RECT 45.155 -99.73 45.245 -98.722 ;
      RECT 45.105 -99.495 45.245 -99.325 ;
      RECT 45.155 -98.308 45.245 -97.3 ;
      RECT 45.105 -97.705 45.245 -97.535 ;
      RECT 45.155 -96.5 45.245 -95.492 ;
      RECT 45.105 -96.265 45.245 -96.095 ;
      RECT 45.155 -95.078 45.245 -94.07 ;
      RECT 45.105 -94.475 45.245 -94.305 ;
      RECT 45.155 -93.27 45.245 -92.262 ;
      RECT 45.105 -93.035 45.245 -92.865 ;
      RECT 45.155 -91.848 45.245 -90.84 ;
      RECT 45.105 -91.245 45.245 -91.075 ;
      RECT 45.155 -90.04 45.245 -89.032 ;
      RECT 45.105 -89.805 45.245 -89.635 ;
      RECT 45.155 -88.618 45.245 -87.61 ;
      RECT 45.105 -88.015 45.245 -87.845 ;
      RECT 45.155 -86.81 45.245 -85.802 ;
      RECT 45.105 -86.575 45.245 -86.405 ;
      RECT 45.155 -85.388 45.245 -84.38 ;
      RECT 45.105 -84.785 45.245 -84.615 ;
      RECT 45.155 -83.58 45.245 -82.572 ;
      RECT 45.105 -83.345 45.245 -83.175 ;
      RECT 45.155 -82.158 45.245 -81.15 ;
      RECT 45.105 -81.555 45.245 -81.385 ;
      RECT 45.155 -80.35 45.245 -79.342 ;
      RECT 45.105 -80.115 45.245 -79.945 ;
      RECT 45.155 -78.928 45.245 -77.92 ;
      RECT 45.105 -78.325 45.245 -78.155 ;
      RECT 45.155 -77.12 45.245 -76.112 ;
      RECT 45.105 -76.885 45.245 -76.715 ;
      RECT 45.155 -75.698 45.245 -74.69 ;
      RECT 45.105 -75.095 45.245 -74.925 ;
      RECT 45.155 -73.89 45.245 -72.882 ;
      RECT 45.105 -73.655 45.245 -73.485 ;
      RECT 45.155 -72.468 45.245 -71.46 ;
      RECT 45.105 -71.865 45.245 -71.695 ;
      RECT 45.155 -70.66 45.245 -69.652 ;
      RECT 45.105 -70.425 45.245 -70.255 ;
      RECT 45.155 -69.238 45.245 -68.23 ;
      RECT 45.105 -68.635 45.245 -68.465 ;
      RECT 45.155 -67.43 45.245 -66.422 ;
      RECT 45.105 -67.195 45.245 -67.025 ;
      RECT 45.155 -66.008 45.245 -65 ;
      RECT 45.105 -65.405 45.245 -65.235 ;
      RECT 45.155 -64.2 45.245 -63.192 ;
      RECT 45.105 -63.965 45.245 -63.795 ;
      RECT 45.155 -62.778 45.245 -61.77 ;
      RECT 45.105 -62.175 45.245 -62.005 ;
      RECT 45.155 -60.97 45.245 -59.962 ;
      RECT 45.105 -60.735 45.245 -60.565 ;
      RECT 45.155 -59.548 45.245 -58.54 ;
      RECT 45.105 -58.945 45.245 -58.775 ;
      RECT 45.155 -57.74 45.245 -56.732 ;
      RECT 45.105 -57.505 45.245 -57.335 ;
      RECT 45.155 -56.318 45.245 -55.31 ;
      RECT 45.105 -55.715 45.245 -55.545 ;
      RECT 45.155 -54.51 45.245 -53.502 ;
      RECT 45.105 -54.275 45.245 -54.105 ;
      RECT 45.155 -53.088 45.245 -52.08 ;
      RECT 45.105 -52.485 45.245 -52.315 ;
      RECT 45.155 -51.28 45.245 -50.272 ;
      RECT 45.105 -51.045 45.245 -50.875 ;
      RECT 45.155 -49.858 45.245 -48.85 ;
      RECT 45.105 -49.255 45.245 -49.085 ;
      RECT 45.155 -48.05 45.245 -47.042 ;
      RECT 45.105 -47.815 45.245 -47.645 ;
      RECT 45.155 -46.628 45.245 -45.62 ;
      RECT 45.105 -46.025 45.245 -45.855 ;
      RECT 45.155 -44.82 45.245 -43.812 ;
      RECT 45.105 -44.585 45.245 -44.415 ;
      RECT 45.155 -43.398 45.245 -42.39 ;
      RECT 45.105 -42.795 45.245 -42.625 ;
      RECT 45.155 -41.59 45.245 -40.582 ;
      RECT 45.105 -41.355 45.245 -41.185 ;
      RECT 45.155 -40.168 45.245 -39.16 ;
      RECT 45.105 -39.565 45.245 -39.395 ;
      RECT 45.155 -38.36 45.245 -37.352 ;
      RECT 45.105 -38.125 45.245 -37.955 ;
      RECT 45.155 -36.938 45.245 -35.93 ;
      RECT 45.105 -36.335 45.245 -36.165 ;
      RECT 45.155 -35.13 45.245 -34.122 ;
      RECT 45.105 -34.895 45.245 -34.725 ;
      RECT 45.155 -33.708 45.245 -32.7 ;
      RECT 45.105 -33.105 45.245 -32.935 ;
      RECT 45.155 -31.9 45.245 -30.892 ;
      RECT 45.105 -31.665 45.245 -31.495 ;
      RECT 45.155 -30.478 45.245 -29.47 ;
      RECT 45.105 -29.875 45.245 -29.705 ;
      RECT 45.155 -28.67 45.245 -27.662 ;
      RECT 45.105 -28.435 45.245 -28.265 ;
      RECT 45.155 -27.248 45.245 -26.24 ;
      RECT 45.105 -26.645 45.245 -26.475 ;
      RECT 45.155 -25.44 45.245 -24.432 ;
      RECT 45.105 -25.205 45.245 -25.035 ;
      RECT 45.155 -24.018 45.245 -23.01 ;
      RECT 45.105 -23.415 45.245 -23.245 ;
      RECT 45.155 -22.21 45.245 -21.202 ;
      RECT 45.105 -21.975 45.245 -21.805 ;
      RECT 45.155 -20.788 45.245 -19.78 ;
      RECT 45.105 -20.185 45.245 -20.015 ;
      RECT 45.155 -18.98 45.245 -17.972 ;
      RECT 45.105 -18.745 45.245 -18.575 ;
      RECT 45.155 -17.558 45.245 -16.55 ;
      RECT 45.105 -16.955 45.245 -16.785 ;
      RECT 45.155 -15.75 45.245 -14.742 ;
      RECT 45.105 -15.515 45.245 -15.345 ;
      RECT 45.155 -14.328 45.245 -13.32 ;
      RECT 45.105 -13.725 45.245 -13.555 ;
      RECT 45.155 -12.52 45.245 -11.512 ;
      RECT 45.105 -12.285 45.245 -12.115 ;
      RECT 45.155 -11.098 45.245 -10.09 ;
      RECT 45.105 -10.495 45.245 -10.325 ;
      RECT 45.155 -9.29 45.245 -8.282 ;
      RECT 45.105 -9.055 45.245 -8.885 ;
      RECT 45.155 -7.868 45.245 -6.86 ;
      RECT 45.105 -7.265 45.245 -7.095 ;
      RECT 45.155 -6.06 45.245 -5.052 ;
      RECT 45.105 -5.825 45.245 -5.655 ;
      RECT 45.155 -4.638 45.245 -3.63 ;
      RECT 45.105 -4.035 45.245 -3.865 ;
      RECT 45.155 -2.83 45.245 -1.822 ;
      RECT 45.105 -2.595 45.245 -2.425 ;
      RECT 45.155 -1.408 45.245 -0.4 ;
      RECT 45.105 -0.805 45.245 -0.635 ;
      RECT 45.155 0.4 45.245 1.408 ;
      RECT 45.105 0.635 45.245 0.805 ;
      RECT 45.03 -114.685 45.205 -114.515 ;
      RECT 45.105 -114.895 45.205 -114.515 ;
      RECT 44.145 -113.555 44.245 -113.09 ;
      RECT 44.51 -113.555 44.61 -113.1 ;
      RECT 44.145 -113.555 44.99 -113.385 ;
      RECT 44.755 -101.538 44.845 -100.531 ;
      RECT 44.755 -101.225 44.895 -101.055 ;
      RECT 44.755 -99.729 44.845 -98.722 ;
      RECT 44.755 -99.205 44.895 -99.035 ;
      RECT 44.755 -98.308 44.845 -97.301 ;
      RECT 44.755 -97.995 44.895 -97.825 ;
      RECT 44.755 -96.499 44.845 -95.492 ;
      RECT 44.755 -95.975 44.895 -95.805 ;
      RECT 44.755 -95.078 44.845 -94.071 ;
      RECT 44.755 -94.765 44.895 -94.595 ;
      RECT 44.755 -93.269 44.845 -92.262 ;
      RECT 44.755 -92.745 44.895 -92.575 ;
      RECT 44.755 -91.848 44.845 -90.841 ;
      RECT 44.755 -91.535 44.895 -91.365 ;
      RECT 44.755 -90.039 44.845 -89.032 ;
      RECT 44.755 -89.515 44.895 -89.345 ;
      RECT 44.755 -88.618 44.845 -87.611 ;
      RECT 44.755 -88.305 44.895 -88.135 ;
      RECT 44.755 -86.809 44.845 -85.802 ;
      RECT 44.755 -86.285 44.895 -86.115 ;
      RECT 44.755 -85.388 44.845 -84.381 ;
      RECT 44.755 -85.075 44.895 -84.905 ;
      RECT 44.755 -83.579 44.845 -82.572 ;
      RECT 44.755 -83.055 44.895 -82.885 ;
      RECT 44.755 -82.158 44.845 -81.151 ;
      RECT 44.755 -81.845 44.895 -81.675 ;
      RECT 44.755 -80.349 44.845 -79.342 ;
      RECT 44.755 -79.825 44.895 -79.655 ;
      RECT 44.755 -78.928 44.845 -77.921 ;
      RECT 44.755 -78.615 44.895 -78.445 ;
      RECT 44.755 -77.119 44.845 -76.112 ;
      RECT 44.755 -76.595 44.895 -76.425 ;
      RECT 44.755 -75.698 44.845 -74.691 ;
      RECT 44.755 -75.385 44.895 -75.215 ;
      RECT 44.755 -73.889 44.845 -72.882 ;
      RECT 44.755 -73.365 44.895 -73.195 ;
      RECT 44.755 -72.468 44.845 -71.461 ;
      RECT 44.755 -72.155 44.895 -71.985 ;
      RECT 44.755 -70.659 44.845 -69.652 ;
      RECT 44.755 -70.135 44.895 -69.965 ;
      RECT 44.755 -69.238 44.845 -68.231 ;
      RECT 44.755 -68.925 44.895 -68.755 ;
      RECT 44.755 -67.429 44.845 -66.422 ;
      RECT 44.755 -66.905 44.895 -66.735 ;
      RECT 44.755 -66.008 44.845 -65.001 ;
      RECT 44.755 -65.695 44.895 -65.525 ;
      RECT 44.755 -64.199 44.845 -63.192 ;
      RECT 44.755 -63.675 44.895 -63.505 ;
      RECT 44.755 -62.778 44.845 -61.771 ;
      RECT 44.755 -62.465 44.895 -62.295 ;
      RECT 44.755 -60.969 44.845 -59.962 ;
      RECT 44.755 -60.445 44.895 -60.275 ;
      RECT 44.755 -59.548 44.845 -58.541 ;
      RECT 44.755 -59.235 44.895 -59.065 ;
      RECT 44.755 -57.739 44.845 -56.732 ;
      RECT 44.755 -57.215 44.895 -57.045 ;
      RECT 44.755 -56.318 44.845 -55.311 ;
      RECT 44.755 -56.005 44.895 -55.835 ;
      RECT 44.755 -54.509 44.845 -53.502 ;
      RECT 44.755 -53.985 44.895 -53.815 ;
      RECT 44.755 -53.088 44.845 -52.081 ;
      RECT 44.755 -52.775 44.895 -52.605 ;
      RECT 44.755 -51.279 44.845 -50.272 ;
      RECT 44.755 -50.755 44.895 -50.585 ;
      RECT 44.755 -49.858 44.845 -48.851 ;
      RECT 44.755 -49.545 44.895 -49.375 ;
      RECT 44.755 -48.049 44.845 -47.042 ;
      RECT 44.755 -47.525 44.895 -47.355 ;
      RECT 44.755 -46.628 44.845 -45.621 ;
      RECT 44.755 -46.315 44.895 -46.145 ;
      RECT 44.755 -44.819 44.845 -43.812 ;
      RECT 44.755 -44.295 44.895 -44.125 ;
      RECT 44.755 -43.398 44.845 -42.391 ;
      RECT 44.755 -43.085 44.895 -42.915 ;
      RECT 44.755 -41.589 44.845 -40.582 ;
      RECT 44.755 -41.065 44.895 -40.895 ;
      RECT 44.755 -40.168 44.845 -39.161 ;
      RECT 44.755 -39.855 44.895 -39.685 ;
      RECT 44.755 -38.359 44.845 -37.352 ;
      RECT 44.755 -37.835 44.895 -37.665 ;
      RECT 44.755 -36.938 44.845 -35.931 ;
      RECT 44.755 -36.625 44.895 -36.455 ;
      RECT 44.755 -35.129 44.845 -34.122 ;
      RECT 44.755 -34.605 44.895 -34.435 ;
      RECT 44.755 -33.708 44.845 -32.701 ;
      RECT 44.755 -33.395 44.895 -33.225 ;
      RECT 44.755 -31.899 44.845 -30.892 ;
      RECT 44.755 -31.375 44.895 -31.205 ;
      RECT 44.755 -30.478 44.845 -29.471 ;
      RECT 44.755 -30.165 44.895 -29.995 ;
      RECT 44.755 -28.669 44.845 -27.662 ;
      RECT 44.755 -28.145 44.895 -27.975 ;
      RECT 44.755 -27.248 44.845 -26.241 ;
      RECT 44.755 -26.935 44.895 -26.765 ;
      RECT 44.755 -25.439 44.845 -24.432 ;
      RECT 44.755 -24.915 44.895 -24.745 ;
      RECT 44.755 -24.018 44.845 -23.011 ;
      RECT 44.755 -23.705 44.895 -23.535 ;
      RECT 44.755 -22.209 44.845 -21.202 ;
      RECT 44.755 -21.685 44.895 -21.515 ;
      RECT 44.755 -20.788 44.845 -19.781 ;
      RECT 44.755 -20.475 44.895 -20.305 ;
      RECT 44.755 -18.979 44.845 -17.972 ;
      RECT 44.755 -18.455 44.895 -18.285 ;
      RECT 44.755 -17.558 44.845 -16.551 ;
      RECT 44.755 -17.245 44.895 -17.075 ;
      RECT 44.755 -15.749 44.845 -14.742 ;
      RECT 44.755 -15.225 44.895 -15.055 ;
      RECT 44.755 -14.328 44.845 -13.321 ;
      RECT 44.755 -14.015 44.895 -13.845 ;
      RECT 44.755 -12.519 44.845 -11.512 ;
      RECT 44.755 -11.995 44.895 -11.825 ;
      RECT 44.755 -11.098 44.845 -10.091 ;
      RECT 44.755 -10.785 44.895 -10.615 ;
      RECT 44.755 -9.289 44.845 -8.282 ;
      RECT 44.755 -8.765 44.895 -8.595 ;
      RECT 44.755 -7.868 44.845 -6.861 ;
      RECT 44.755 -7.555 44.895 -7.385 ;
      RECT 44.755 -6.059 44.845 -5.052 ;
      RECT 44.755 -5.535 44.895 -5.365 ;
      RECT 44.755 -4.638 44.845 -3.631 ;
      RECT 44.755 -4.325 44.895 -4.155 ;
      RECT 44.755 -2.829 44.845 -1.822 ;
      RECT 44.755 -2.305 44.895 -2.135 ;
      RECT 44.755 -1.408 44.845 -0.401 ;
      RECT 44.755 -1.095 44.895 -0.925 ;
      RECT 44.755 0.401 44.845 1.408 ;
      RECT 44.755 0.925 44.895 1.095 ;
      RECT 44.44 -114.685 44.61 -114.515 ;
      RECT 44.51 -114.895 44.61 -114.515 ;
      RECT 43.955 -101.538 44.045 -100.53 ;
      RECT 43.905 -100.935 44.045 -100.765 ;
      RECT 43.955 -99.73 44.045 -98.722 ;
      RECT 43.905 -99.495 44.045 -99.325 ;
      RECT 43.955 -98.308 44.045 -97.3 ;
      RECT 43.905 -97.705 44.045 -97.535 ;
      RECT 43.955 -96.5 44.045 -95.492 ;
      RECT 43.905 -96.265 44.045 -96.095 ;
      RECT 43.955 -95.078 44.045 -94.07 ;
      RECT 43.905 -94.475 44.045 -94.305 ;
      RECT 43.955 -93.27 44.045 -92.262 ;
      RECT 43.905 -93.035 44.045 -92.865 ;
      RECT 43.955 -91.848 44.045 -90.84 ;
      RECT 43.905 -91.245 44.045 -91.075 ;
      RECT 43.955 -90.04 44.045 -89.032 ;
      RECT 43.905 -89.805 44.045 -89.635 ;
      RECT 43.955 -88.618 44.045 -87.61 ;
      RECT 43.905 -88.015 44.045 -87.845 ;
      RECT 43.955 -86.81 44.045 -85.802 ;
      RECT 43.905 -86.575 44.045 -86.405 ;
      RECT 43.955 -85.388 44.045 -84.38 ;
      RECT 43.905 -84.785 44.045 -84.615 ;
      RECT 43.955 -83.58 44.045 -82.572 ;
      RECT 43.905 -83.345 44.045 -83.175 ;
      RECT 43.955 -82.158 44.045 -81.15 ;
      RECT 43.905 -81.555 44.045 -81.385 ;
      RECT 43.955 -80.35 44.045 -79.342 ;
      RECT 43.905 -80.115 44.045 -79.945 ;
      RECT 43.955 -78.928 44.045 -77.92 ;
      RECT 43.905 -78.325 44.045 -78.155 ;
      RECT 43.955 -77.12 44.045 -76.112 ;
      RECT 43.905 -76.885 44.045 -76.715 ;
      RECT 43.955 -75.698 44.045 -74.69 ;
      RECT 43.905 -75.095 44.045 -74.925 ;
      RECT 43.955 -73.89 44.045 -72.882 ;
      RECT 43.905 -73.655 44.045 -73.485 ;
      RECT 43.955 -72.468 44.045 -71.46 ;
      RECT 43.905 -71.865 44.045 -71.695 ;
      RECT 43.955 -70.66 44.045 -69.652 ;
      RECT 43.905 -70.425 44.045 -70.255 ;
      RECT 43.955 -69.238 44.045 -68.23 ;
      RECT 43.905 -68.635 44.045 -68.465 ;
      RECT 43.955 -67.43 44.045 -66.422 ;
      RECT 43.905 -67.195 44.045 -67.025 ;
      RECT 43.955 -66.008 44.045 -65 ;
      RECT 43.905 -65.405 44.045 -65.235 ;
      RECT 43.955 -64.2 44.045 -63.192 ;
      RECT 43.905 -63.965 44.045 -63.795 ;
      RECT 43.955 -62.778 44.045 -61.77 ;
      RECT 43.905 -62.175 44.045 -62.005 ;
      RECT 43.955 -60.97 44.045 -59.962 ;
      RECT 43.905 -60.735 44.045 -60.565 ;
      RECT 43.955 -59.548 44.045 -58.54 ;
      RECT 43.905 -58.945 44.045 -58.775 ;
      RECT 43.955 -57.74 44.045 -56.732 ;
      RECT 43.905 -57.505 44.045 -57.335 ;
      RECT 43.955 -56.318 44.045 -55.31 ;
      RECT 43.905 -55.715 44.045 -55.545 ;
      RECT 43.955 -54.51 44.045 -53.502 ;
      RECT 43.905 -54.275 44.045 -54.105 ;
      RECT 43.955 -53.088 44.045 -52.08 ;
      RECT 43.905 -52.485 44.045 -52.315 ;
      RECT 43.955 -51.28 44.045 -50.272 ;
      RECT 43.905 -51.045 44.045 -50.875 ;
      RECT 43.955 -49.858 44.045 -48.85 ;
      RECT 43.905 -49.255 44.045 -49.085 ;
      RECT 43.955 -48.05 44.045 -47.042 ;
      RECT 43.905 -47.815 44.045 -47.645 ;
      RECT 43.955 -46.628 44.045 -45.62 ;
      RECT 43.905 -46.025 44.045 -45.855 ;
      RECT 43.955 -44.82 44.045 -43.812 ;
      RECT 43.905 -44.585 44.045 -44.415 ;
      RECT 43.955 -43.398 44.045 -42.39 ;
      RECT 43.905 -42.795 44.045 -42.625 ;
      RECT 43.955 -41.59 44.045 -40.582 ;
      RECT 43.905 -41.355 44.045 -41.185 ;
      RECT 43.955 -40.168 44.045 -39.16 ;
      RECT 43.905 -39.565 44.045 -39.395 ;
      RECT 43.955 -38.36 44.045 -37.352 ;
      RECT 43.905 -38.125 44.045 -37.955 ;
      RECT 43.955 -36.938 44.045 -35.93 ;
      RECT 43.905 -36.335 44.045 -36.165 ;
      RECT 43.955 -35.13 44.045 -34.122 ;
      RECT 43.905 -34.895 44.045 -34.725 ;
      RECT 43.955 -33.708 44.045 -32.7 ;
      RECT 43.905 -33.105 44.045 -32.935 ;
      RECT 43.955 -31.9 44.045 -30.892 ;
      RECT 43.905 -31.665 44.045 -31.495 ;
      RECT 43.955 -30.478 44.045 -29.47 ;
      RECT 43.905 -29.875 44.045 -29.705 ;
      RECT 43.955 -28.67 44.045 -27.662 ;
      RECT 43.905 -28.435 44.045 -28.265 ;
      RECT 43.955 -27.248 44.045 -26.24 ;
      RECT 43.905 -26.645 44.045 -26.475 ;
      RECT 43.955 -25.44 44.045 -24.432 ;
      RECT 43.905 -25.205 44.045 -25.035 ;
      RECT 43.955 -24.018 44.045 -23.01 ;
      RECT 43.905 -23.415 44.045 -23.245 ;
      RECT 43.955 -22.21 44.045 -21.202 ;
      RECT 43.905 -21.975 44.045 -21.805 ;
      RECT 43.955 -20.788 44.045 -19.78 ;
      RECT 43.905 -20.185 44.045 -20.015 ;
      RECT 43.955 -18.98 44.045 -17.972 ;
      RECT 43.905 -18.745 44.045 -18.575 ;
      RECT 43.955 -17.558 44.045 -16.55 ;
      RECT 43.905 -16.955 44.045 -16.785 ;
      RECT 43.955 -15.75 44.045 -14.742 ;
      RECT 43.905 -15.515 44.045 -15.345 ;
      RECT 43.955 -14.328 44.045 -13.32 ;
      RECT 43.905 -13.725 44.045 -13.555 ;
      RECT 43.955 -12.52 44.045 -11.512 ;
      RECT 43.905 -12.285 44.045 -12.115 ;
      RECT 43.955 -11.098 44.045 -10.09 ;
      RECT 43.905 -10.495 44.045 -10.325 ;
      RECT 43.955 -9.29 44.045 -8.282 ;
      RECT 43.905 -9.055 44.045 -8.885 ;
      RECT 43.955 -7.868 44.045 -6.86 ;
      RECT 43.905 -7.265 44.045 -7.095 ;
      RECT 43.955 -6.06 44.045 -5.052 ;
      RECT 43.905 -5.825 44.045 -5.655 ;
      RECT 43.955 -4.638 44.045 -3.63 ;
      RECT 43.905 -4.035 44.045 -3.865 ;
      RECT 43.955 -2.83 44.045 -1.822 ;
      RECT 43.905 -2.595 44.045 -2.425 ;
      RECT 43.955 -1.408 44.045 -0.4 ;
      RECT 43.905 -0.805 44.045 -0.635 ;
      RECT 43.955 0.4 44.045 1.408 ;
      RECT 43.905 0.635 44.045 0.805 ;
      RECT 43.555 -101.538 43.645 -100.531 ;
      RECT 43.555 -101.225 43.695 -101.055 ;
      RECT 43.555 -99.729 43.645 -98.722 ;
      RECT 43.555 -99.205 43.695 -99.035 ;
      RECT 43.555 -98.308 43.645 -97.301 ;
      RECT 43.555 -97.995 43.695 -97.825 ;
      RECT 43.555 -96.499 43.645 -95.492 ;
      RECT 43.555 -95.975 43.695 -95.805 ;
      RECT 43.555 -95.078 43.645 -94.071 ;
      RECT 43.555 -94.765 43.695 -94.595 ;
      RECT 43.555 -93.269 43.645 -92.262 ;
      RECT 43.555 -92.745 43.695 -92.575 ;
      RECT 43.555 -91.848 43.645 -90.841 ;
      RECT 43.555 -91.535 43.695 -91.365 ;
      RECT 43.555 -90.039 43.645 -89.032 ;
      RECT 43.555 -89.515 43.695 -89.345 ;
      RECT 43.555 -88.618 43.645 -87.611 ;
      RECT 43.555 -88.305 43.695 -88.135 ;
      RECT 43.555 -86.809 43.645 -85.802 ;
      RECT 43.555 -86.285 43.695 -86.115 ;
      RECT 43.555 -85.388 43.645 -84.381 ;
      RECT 43.555 -85.075 43.695 -84.905 ;
      RECT 43.555 -83.579 43.645 -82.572 ;
      RECT 43.555 -83.055 43.695 -82.885 ;
      RECT 43.555 -82.158 43.645 -81.151 ;
      RECT 43.555 -81.845 43.695 -81.675 ;
      RECT 43.555 -80.349 43.645 -79.342 ;
      RECT 43.555 -79.825 43.695 -79.655 ;
      RECT 43.555 -78.928 43.645 -77.921 ;
      RECT 43.555 -78.615 43.695 -78.445 ;
      RECT 43.555 -77.119 43.645 -76.112 ;
      RECT 43.555 -76.595 43.695 -76.425 ;
      RECT 43.555 -75.698 43.645 -74.691 ;
      RECT 43.555 -75.385 43.695 -75.215 ;
      RECT 43.555 -73.889 43.645 -72.882 ;
      RECT 43.555 -73.365 43.695 -73.195 ;
      RECT 43.555 -72.468 43.645 -71.461 ;
      RECT 43.555 -72.155 43.695 -71.985 ;
      RECT 43.555 -70.659 43.645 -69.652 ;
      RECT 43.555 -70.135 43.695 -69.965 ;
      RECT 43.555 -69.238 43.645 -68.231 ;
      RECT 43.555 -68.925 43.695 -68.755 ;
      RECT 43.555 -67.429 43.645 -66.422 ;
      RECT 43.555 -66.905 43.695 -66.735 ;
      RECT 43.555 -66.008 43.645 -65.001 ;
      RECT 43.555 -65.695 43.695 -65.525 ;
      RECT 43.555 -64.199 43.645 -63.192 ;
      RECT 43.555 -63.675 43.695 -63.505 ;
      RECT 43.555 -62.778 43.645 -61.771 ;
      RECT 43.555 -62.465 43.695 -62.295 ;
      RECT 43.555 -60.969 43.645 -59.962 ;
      RECT 43.555 -60.445 43.695 -60.275 ;
      RECT 43.555 -59.548 43.645 -58.541 ;
      RECT 43.555 -59.235 43.695 -59.065 ;
      RECT 43.555 -57.739 43.645 -56.732 ;
      RECT 43.555 -57.215 43.695 -57.045 ;
      RECT 43.555 -56.318 43.645 -55.311 ;
      RECT 43.555 -56.005 43.695 -55.835 ;
      RECT 43.555 -54.509 43.645 -53.502 ;
      RECT 43.555 -53.985 43.695 -53.815 ;
      RECT 43.555 -53.088 43.645 -52.081 ;
      RECT 43.555 -52.775 43.695 -52.605 ;
      RECT 43.555 -51.279 43.645 -50.272 ;
      RECT 43.555 -50.755 43.695 -50.585 ;
      RECT 43.555 -49.858 43.645 -48.851 ;
      RECT 43.555 -49.545 43.695 -49.375 ;
      RECT 43.555 -48.049 43.645 -47.042 ;
      RECT 43.555 -47.525 43.695 -47.355 ;
      RECT 43.555 -46.628 43.645 -45.621 ;
      RECT 43.555 -46.315 43.695 -46.145 ;
      RECT 43.555 -44.819 43.645 -43.812 ;
      RECT 43.555 -44.295 43.695 -44.125 ;
      RECT 43.555 -43.398 43.645 -42.391 ;
      RECT 43.555 -43.085 43.695 -42.915 ;
      RECT 43.555 -41.589 43.645 -40.582 ;
      RECT 43.555 -41.065 43.695 -40.895 ;
      RECT 43.555 -40.168 43.645 -39.161 ;
      RECT 43.555 -39.855 43.695 -39.685 ;
      RECT 43.555 -38.359 43.645 -37.352 ;
      RECT 43.555 -37.835 43.695 -37.665 ;
      RECT 43.555 -36.938 43.645 -35.931 ;
      RECT 43.555 -36.625 43.695 -36.455 ;
      RECT 43.555 -35.129 43.645 -34.122 ;
      RECT 43.555 -34.605 43.695 -34.435 ;
      RECT 43.555 -33.708 43.645 -32.701 ;
      RECT 43.555 -33.395 43.695 -33.225 ;
      RECT 43.555 -31.899 43.645 -30.892 ;
      RECT 43.555 -31.375 43.695 -31.205 ;
      RECT 43.555 -30.478 43.645 -29.471 ;
      RECT 43.555 -30.165 43.695 -29.995 ;
      RECT 43.555 -28.669 43.645 -27.662 ;
      RECT 43.555 -28.145 43.695 -27.975 ;
      RECT 43.555 -27.248 43.645 -26.241 ;
      RECT 43.555 -26.935 43.695 -26.765 ;
      RECT 43.555 -25.439 43.645 -24.432 ;
      RECT 43.555 -24.915 43.695 -24.745 ;
      RECT 43.555 -24.018 43.645 -23.011 ;
      RECT 43.555 -23.705 43.695 -23.535 ;
      RECT 43.555 -22.209 43.645 -21.202 ;
      RECT 43.555 -21.685 43.695 -21.515 ;
      RECT 43.555 -20.788 43.645 -19.781 ;
      RECT 43.555 -20.475 43.695 -20.305 ;
      RECT 43.555 -18.979 43.645 -17.972 ;
      RECT 43.555 -18.455 43.695 -18.285 ;
      RECT 43.555 -17.558 43.645 -16.551 ;
      RECT 43.555 -17.245 43.695 -17.075 ;
      RECT 43.555 -15.749 43.645 -14.742 ;
      RECT 43.555 -15.225 43.695 -15.055 ;
      RECT 43.555 -14.328 43.645 -13.321 ;
      RECT 43.555 -14.015 43.695 -13.845 ;
      RECT 43.555 -12.519 43.645 -11.512 ;
      RECT 43.555 -11.995 43.695 -11.825 ;
      RECT 43.555 -11.098 43.645 -10.091 ;
      RECT 43.555 -10.785 43.695 -10.615 ;
      RECT 43.555 -9.289 43.645 -8.282 ;
      RECT 43.555 -8.765 43.695 -8.595 ;
      RECT 43.555 -7.868 43.645 -6.861 ;
      RECT 43.555 -7.555 43.695 -7.385 ;
      RECT 43.555 -6.059 43.645 -5.052 ;
      RECT 43.555 -5.535 43.695 -5.365 ;
      RECT 43.555 -4.638 43.645 -3.631 ;
      RECT 43.555 -4.325 43.695 -4.155 ;
      RECT 43.555 -2.829 43.645 -1.822 ;
      RECT 43.555 -2.305 43.695 -2.135 ;
      RECT 43.555 -1.408 43.645 -0.401 ;
      RECT 43.555 -1.095 43.695 -0.925 ;
      RECT 43.555 0.401 43.645 1.408 ;
      RECT 43.555 0.925 43.695 1.095 ;
      RECT 39.385 -108.935 43.165 -108.815 ;
      RECT 40.705 -109.475 40.805 -108.815 ;
      RECT 40.145 -109.475 40.245 -108.815 ;
      RECT 39.585 -109.475 39.685 -108.815 ;
      RECT 42.755 -101.538 42.845 -100.53 ;
      RECT 42.705 -100.935 42.845 -100.765 ;
      RECT 42.755 -99.73 42.845 -98.722 ;
      RECT 42.705 -99.495 42.845 -99.325 ;
      RECT 42.755 -98.308 42.845 -97.3 ;
      RECT 42.705 -97.705 42.845 -97.535 ;
      RECT 42.755 -96.5 42.845 -95.492 ;
      RECT 42.705 -96.265 42.845 -96.095 ;
      RECT 42.755 -95.078 42.845 -94.07 ;
      RECT 42.705 -94.475 42.845 -94.305 ;
      RECT 42.755 -93.27 42.845 -92.262 ;
      RECT 42.705 -93.035 42.845 -92.865 ;
      RECT 42.755 -91.848 42.845 -90.84 ;
      RECT 42.705 -91.245 42.845 -91.075 ;
      RECT 42.755 -90.04 42.845 -89.032 ;
      RECT 42.705 -89.805 42.845 -89.635 ;
      RECT 42.755 -88.618 42.845 -87.61 ;
      RECT 42.705 -88.015 42.845 -87.845 ;
      RECT 42.755 -86.81 42.845 -85.802 ;
      RECT 42.705 -86.575 42.845 -86.405 ;
      RECT 42.755 -85.388 42.845 -84.38 ;
      RECT 42.705 -84.785 42.845 -84.615 ;
      RECT 42.755 -83.58 42.845 -82.572 ;
      RECT 42.705 -83.345 42.845 -83.175 ;
      RECT 42.755 -82.158 42.845 -81.15 ;
      RECT 42.705 -81.555 42.845 -81.385 ;
      RECT 42.755 -80.35 42.845 -79.342 ;
      RECT 42.705 -80.115 42.845 -79.945 ;
      RECT 42.755 -78.928 42.845 -77.92 ;
      RECT 42.705 -78.325 42.845 -78.155 ;
      RECT 42.755 -77.12 42.845 -76.112 ;
      RECT 42.705 -76.885 42.845 -76.715 ;
      RECT 42.755 -75.698 42.845 -74.69 ;
      RECT 42.705 -75.095 42.845 -74.925 ;
      RECT 42.755 -73.89 42.845 -72.882 ;
      RECT 42.705 -73.655 42.845 -73.485 ;
      RECT 42.755 -72.468 42.845 -71.46 ;
      RECT 42.705 -71.865 42.845 -71.695 ;
      RECT 42.755 -70.66 42.845 -69.652 ;
      RECT 42.705 -70.425 42.845 -70.255 ;
      RECT 42.755 -69.238 42.845 -68.23 ;
      RECT 42.705 -68.635 42.845 -68.465 ;
      RECT 42.755 -67.43 42.845 -66.422 ;
      RECT 42.705 -67.195 42.845 -67.025 ;
      RECT 42.755 -66.008 42.845 -65 ;
      RECT 42.705 -65.405 42.845 -65.235 ;
      RECT 42.755 -64.2 42.845 -63.192 ;
      RECT 42.705 -63.965 42.845 -63.795 ;
      RECT 42.755 -62.778 42.845 -61.77 ;
      RECT 42.705 -62.175 42.845 -62.005 ;
      RECT 42.755 -60.97 42.845 -59.962 ;
      RECT 42.705 -60.735 42.845 -60.565 ;
      RECT 42.755 -59.548 42.845 -58.54 ;
      RECT 42.705 -58.945 42.845 -58.775 ;
      RECT 42.755 -57.74 42.845 -56.732 ;
      RECT 42.705 -57.505 42.845 -57.335 ;
      RECT 42.755 -56.318 42.845 -55.31 ;
      RECT 42.705 -55.715 42.845 -55.545 ;
      RECT 42.755 -54.51 42.845 -53.502 ;
      RECT 42.705 -54.275 42.845 -54.105 ;
      RECT 42.755 -53.088 42.845 -52.08 ;
      RECT 42.705 -52.485 42.845 -52.315 ;
      RECT 42.755 -51.28 42.845 -50.272 ;
      RECT 42.705 -51.045 42.845 -50.875 ;
      RECT 42.755 -49.858 42.845 -48.85 ;
      RECT 42.705 -49.255 42.845 -49.085 ;
      RECT 42.755 -48.05 42.845 -47.042 ;
      RECT 42.705 -47.815 42.845 -47.645 ;
      RECT 42.755 -46.628 42.845 -45.62 ;
      RECT 42.705 -46.025 42.845 -45.855 ;
      RECT 42.755 -44.82 42.845 -43.812 ;
      RECT 42.705 -44.585 42.845 -44.415 ;
      RECT 42.755 -43.398 42.845 -42.39 ;
      RECT 42.705 -42.795 42.845 -42.625 ;
      RECT 42.755 -41.59 42.845 -40.582 ;
      RECT 42.705 -41.355 42.845 -41.185 ;
      RECT 42.755 -40.168 42.845 -39.16 ;
      RECT 42.705 -39.565 42.845 -39.395 ;
      RECT 42.755 -38.36 42.845 -37.352 ;
      RECT 42.705 -38.125 42.845 -37.955 ;
      RECT 42.755 -36.938 42.845 -35.93 ;
      RECT 42.705 -36.335 42.845 -36.165 ;
      RECT 42.755 -35.13 42.845 -34.122 ;
      RECT 42.705 -34.895 42.845 -34.725 ;
      RECT 42.755 -33.708 42.845 -32.7 ;
      RECT 42.705 -33.105 42.845 -32.935 ;
      RECT 42.755 -31.9 42.845 -30.892 ;
      RECT 42.705 -31.665 42.845 -31.495 ;
      RECT 42.755 -30.478 42.845 -29.47 ;
      RECT 42.705 -29.875 42.845 -29.705 ;
      RECT 42.755 -28.67 42.845 -27.662 ;
      RECT 42.705 -28.435 42.845 -28.265 ;
      RECT 42.755 -27.248 42.845 -26.24 ;
      RECT 42.705 -26.645 42.845 -26.475 ;
      RECT 42.755 -25.44 42.845 -24.432 ;
      RECT 42.705 -25.205 42.845 -25.035 ;
      RECT 42.755 -24.018 42.845 -23.01 ;
      RECT 42.705 -23.415 42.845 -23.245 ;
      RECT 42.755 -22.21 42.845 -21.202 ;
      RECT 42.705 -21.975 42.845 -21.805 ;
      RECT 42.755 -20.788 42.845 -19.78 ;
      RECT 42.705 -20.185 42.845 -20.015 ;
      RECT 42.755 -18.98 42.845 -17.972 ;
      RECT 42.705 -18.745 42.845 -18.575 ;
      RECT 42.755 -17.558 42.845 -16.55 ;
      RECT 42.705 -16.955 42.845 -16.785 ;
      RECT 42.755 -15.75 42.845 -14.742 ;
      RECT 42.705 -15.515 42.845 -15.345 ;
      RECT 42.755 -14.328 42.845 -13.32 ;
      RECT 42.705 -13.725 42.845 -13.555 ;
      RECT 42.755 -12.52 42.845 -11.512 ;
      RECT 42.705 -12.285 42.845 -12.115 ;
      RECT 42.755 -11.098 42.845 -10.09 ;
      RECT 42.705 -10.495 42.845 -10.325 ;
      RECT 42.755 -9.29 42.845 -8.282 ;
      RECT 42.705 -9.055 42.845 -8.885 ;
      RECT 42.755 -7.868 42.845 -6.86 ;
      RECT 42.705 -7.265 42.845 -7.095 ;
      RECT 42.755 -6.06 42.845 -5.052 ;
      RECT 42.705 -5.825 42.845 -5.655 ;
      RECT 42.755 -4.638 42.845 -3.63 ;
      RECT 42.705 -4.035 42.845 -3.865 ;
      RECT 42.755 -2.83 42.845 -1.822 ;
      RECT 42.705 -2.595 42.845 -2.425 ;
      RECT 42.755 -1.408 42.845 -0.4 ;
      RECT 42.705 -0.805 42.845 -0.635 ;
      RECT 42.755 0.4 42.845 1.408 ;
      RECT 42.705 0.635 42.845 0.805 ;
      RECT 41.325 -111.685 42.805 -111.585 ;
      RECT 41.325 -112.195 41.425 -111.585 ;
      RECT 41.545 -109.15 42.805 -109.05 ;
      RECT 42.705 -109.475 42.805 -109.05 ;
      RECT 42.145 -109.475 42.245 -109.05 ;
      RECT 41.585 -109.475 41.685 -109.05 ;
      RECT 42.355 -101.538 42.445 -100.531 ;
      RECT 42.355 -101.225 42.495 -101.055 ;
      RECT 42.355 -99.729 42.445 -98.722 ;
      RECT 42.355 -99.205 42.495 -99.035 ;
      RECT 42.355 -98.308 42.445 -97.301 ;
      RECT 42.355 -97.995 42.495 -97.825 ;
      RECT 42.355 -96.499 42.445 -95.492 ;
      RECT 42.355 -95.975 42.495 -95.805 ;
      RECT 42.355 -95.078 42.445 -94.071 ;
      RECT 42.355 -94.765 42.495 -94.595 ;
      RECT 42.355 -93.269 42.445 -92.262 ;
      RECT 42.355 -92.745 42.495 -92.575 ;
      RECT 42.355 -91.848 42.445 -90.841 ;
      RECT 42.355 -91.535 42.495 -91.365 ;
      RECT 42.355 -90.039 42.445 -89.032 ;
      RECT 42.355 -89.515 42.495 -89.345 ;
      RECT 42.355 -88.618 42.445 -87.611 ;
      RECT 42.355 -88.305 42.495 -88.135 ;
      RECT 42.355 -86.809 42.445 -85.802 ;
      RECT 42.355 -86.285 42.495 -86.115 ;
      RECT 42.355 -85.388 42.445 -84.381 ;
      RECT 42.355 -85.075 42.495 -84.905 ;
      RECT 42.355 -83.579 42.445 -82.572 ;
      RECT 42.355 -83.055 42.495 -82.885 ;
      RECT 42.355 -82.158 42.445 -81.151 ;
      RECT 42.355 -81.845 42.495 -81.675 ;
      RECT 42.355 -80.349 42.445 -79.342 ;
      RECT 42.355 -79.825 42.495 -79.655 ;
      RECT 42.355 -78.928 42.445 -77.921 ;
      RECT 42.355 -78.615 42.495 -78.445 ;
      RECT 42.355 -77.119 42.445 -76.112 ;
      RECT 42.355 -76.595 42.495 -76.425 ;
      RECT 42.355 -75.698 42.445 -74.691 ;
      RECT 42.355 -75.385 42.495 -75.215 ;
      RECT 42.355 -73.889 42.445 -72.882 ;
      RECT 42.355 -73.365 42.495 -73.195 ;
      RECT 42.355 -72.468 42.445 -71.461 ;
      RECT 42.355 -72.155 42.495 -71.985 ;
      RECT 42.355 -70.659 42.445 -69.652 ;
      RECT 42.355 -70.135 42.495 -69.965 ;
      RECT 42.355 -69.238 42.445 -68.231 ;
      RECT 42.355 -68.925 42.495 -68.755 ;
      RECT 42.355 -67.429 42.445 -66.422 ;
      RECT 42.355 -66.905 42.495 -66.735 ;
      RECT 42.355 -66.008 42.445 -65.001 ;
      RECT 42.355 -65.695 42.495 -65.525 ;
      RECT 42.355 -64.199 42.445 -63.192 ;
      RECT 42.355 -63.675 42.495 -63.505 ;
      RECT 42.355 -62.778 42.445 -61.771 ;
      RECT 42.355 -62.465 42.495 -62.295 ;
      RECT 42.355 -60.969 42.445 -59.962 ;
      RECT 42.355 -60.445 42.495 -60.275 ;
      RECT 42.355 -59.548 42.445 -58.541 ;
      RECT 42.355 -59.235 42.495 -59.065 ;
      RECT 42.355 -57.739 42.445 -56.732 ;
      RECT 42.355 -57.215 42.495 -57.045 ;
      RECT 42.355 -56.318 42.445 -55.311 ;
      RECT 42.355 -56.005 42.495 -55.835 ;
      RECT 42.355 -54.509 42.445 -53.502 ;
      RECT 42.355 -53.985 42.495 -53.815 ;
      RECT 42.355 -53.088 42.445 -52.081 ;
      RECT 42.355 -52.775 42.495 -52.605 ;
      RECT 42.355 -51.279 42.445 -50.272 ;
      RECT 42.355 -50.755 42.495 -50.585 ;
      RECT 42.355 -49.858 42.445 -48.851 ;
      RECT 42.355 -49.545 42.495 -49.375 ;
      RECT 42.355 -48.049 42.445 -47.042 ;
      RECT 42.355 -47.525 42.495 -47.355 ;
      RECT 42.355 -46.628 42.445 -45.621 ;
      RECT 42.355 -46.315 42.495 -46.145 ;
      RECT 42.355 -44.819 42.445 -43.812 ;
      RECT 42.355 -44.295 42.495 -44.125 ;
      RECT 42.355 -43.398 42.445 -42.391 ;
      RECT 42.355 -43.085 42.495 -42.915 ;
      RECT 42.355 -41.589 42.445 -40.582 ;
      RECT 42.355 -41.065 42.495 -40.895 ;
      RECT 42.355 -40.168 42.445 -39.161 ;
      RECT 42.355 -39.855 42.495 -39.685 ;
      RECT 42.355 -38.359 42.445 -37.352 ;
      RECT 42.355 -37.835 42.495 -37.665 ;
      RECT 42.355 -36.938 42.445 -35.931 ;
      RECT 42.355 -36.625 42.495 -36.455 ;
      RECT 42.355 -35.129 42.445 -34.122 ;
      RECT 42.355 -34.605 42.495 -34.435 ;
      RECT 42.355 -33.708 42.445 -32.701 ;
      RECT 42.355 -33.395 42.495 -33.225 ;
      RECT 42.355 -31.899 42.445 -30.892 ;
      RECT 42.355 -31.375 42.495 -31.205 ;
      RECT 42.355 -30.478 42.445 -29.471 ;
      RECT 42.355 -30.165 42.495 -29.995 ;
      RECT 42.355 -28.669 42.445 -27.662 ;
      RECT 42.355 -28.145 42.495 -27.975 ;
      RECT 42.355 -27.248 42.445 -26.241 ;
      RECT 42.355 -26.935 42.495 -26.765 ;
      RECT 42.355 -25.439 42.445 -24.432 ;
      RECT 42.355 -24.915 42.495 -24.745 ;
      RECT 42.355 -24.018 42.445 -23.011 ;
      RECT 42.355 -23.705 42.495 -23.535 ;
      RECT 42.355 -22.209 42.445 -21.202 ;
      RECT 42.355 -21.685 42.495 -21.515 ;
      RECT 42.355 -20.788 42.445 -19.781 ;
      RECT 42.355 -20.475 42.495 -20.305 ;
      RECT 42.355 -18.979 42.445 -17.972 ;
      RECT 42.355 -18.455 42.495 -18.285 ;
      RECT 42.355 -17.558 42.445 -16.551 ;
      RECT 42.355 -17.245 42.495 -17.075 ;
      RECT 42.355 -15.749 42.445 -14.742 ;
      RECT 42.355 -15.225 42.495 -15.055 ;
      RECT 42.355 -14.328 42.445 -13.321 ;
      RECT 42.355 -14.015 42.495 -13.845 ;
      RECT 42.355 -12.519 42.445 -11.512 ;
      RECT 42.355 -11.995 42.495 -11.825 ;
      RECT 42.355 -11.098 42.445 -10.091 ;
      RECT 42.355 -10.785 42.495 -10.615 ;
      RECT 42.355 -9.289 42.445 -8.282 ;
      RECT 42.355 -8.765 42.495 -8.595 ;
      RECT 42.355 -7.868 42.445 -6.861 ;
      RECT 42.355 -7.555 42.495 -7.385 ;
      RECT 42.355 -6.059 42.445 -5.052 ;
      RECT 42.355 -5.535 42.495 -5.365 ;
      RECT 42.355 -4.638 42.445 -3.631 ;
      RECT 42.355 -4.325 42.495 -4.155 ;
      RECT 42.355 -2.829 42.445 -1.822 ;
      RECT 42.355 -2.305 42.495 -2.135 ;
      RECT 42.355 -1.408 42.445 -0.401 ;
      RECT 42.355 -1.095 42.495 -0.925 ;
      RECT 42.355 0.401 42.445 1.408 ;
      RECT 42.355 0.925 42.495 1.095 ;
      RECT 41.685 -111.495 41.855 -111.385 ;
      RECT 38.535 -111.495 41.855 -111.395 ;
      RECT 41.555 -101.538 41.645 -100.53 ;
      RECT 41.505 -100.935 41.645 -100.765 ;
      RECT 41.555 -99.73 41.645 -98.722 ;
      RECT 41.505 -99.495 41.645 -99.325 ;
      RECT 41.555 -98.308 41.645 -97.3 ;
      RECT 41.505 -97.705 41.645 -97.535 ;
      RECT 41.555 -96.5 41.645 -95.492 ;
      RECT 41.505 -96.265 41.645 -96.095 ;
      RECT 41.555 -95.078 41.645 -94.07 ;
      RECT 41.505 -94.475 41.645 -94.305 ;
      RECT 41.555 -93.27 41.645 -92.262 ;
      RECT 41.505 -93.035 41.645 -92.865 ;
      RECT 41.555 -91.848 41.645 -90.84 ;
      RECT 41.505 -91.245 41.645 -91.075 ;
      RECT 41.555 -90.04 41.645 -89.032 ;
      RECT 41.505 -89.805 41.645 -89.635 ;
      RECT 41.555 -88.618 41.645 -87.61 ;
      RECT 41.505 -88.015 41.645 -87.845 ;
      RECT 41.555 -86.81 41.645 -85.802 ;
      RECT 41.505 -86.575 41.645 -86.405 ;
      RECT 41.555 -85.388 41.645 -84.38 ;
      RECT 41.505 -84.785 41.645 -84.615 ;
      RECT 41.555 -83.58 41.645 -82.572 ;
      RECT 41.505 -83.345 41.645 -83.175 ;
      RECT 41.555 -82.158 41.645 -81.15 ;
      RECT 41.505 -81.555 41.645 -81.385 ;
      RECT 41.555 -80.35 41.645 -79.342 ;
      RECT 41.505 -80.115 41.645 -79.945 ;
      RECT 41.555 -78.928 41.645 -77.92 ;
      RECT 41.505 -78.325 41.645 -78.155 ;
      RECT 41.555 -77.12 41.645 -76.112 ;
      RECT 41.505 -76.885 41.645 -76.715 ;
      RECT 41.555 -75.698 41.645 -74.69 ;
      RECT 41.505 -75.095 41.645 -74.925 ;
      RECT 41.555 -73.89 41.645 -72.882 ;
      RECT 41.505 -73.655 41.645 -73.485 ;
      RECT 41.555 -72.468 41.645 -71.46 ;
      RECT 41.505 -71.865 41.645 -71.695 ;
      RECT 41.555 -70.66 41.645 -69.652 ;
      RECT 41.505 -70.425 41.645 -70.255 ;
      RECT 41.555 -69.238 41.645 -68.23 ;
      RECT 41.505 -68.635 41.645 -68.465 ;
      RECT 41.555 -67.43 41.645 -66.422 ;
      RECT 41.505 -67.195 41.645 -67.025 ;
      RECT 41.555 -66.008 41.645 -65 ;
      RECT 41.505 -65.405 41.645 -65.235 ;
      RECT 41.555 -64.2 41.645 -63.192 ;
      RECT 41.505 -63.965 41.645 -63.795 ;
      RECT 41.555 -62.778 41.645 -61.77 ;
      RECT 41.505 -62.175 41.645 -62.005 ;
      RECT 41.555 -60.97 41.645 -59.962 ;
      RECT 41.505 -60.735 41.645 -60.565 ;
      RECT 41.555 -59.548 41.645 -58.54 ;
      RECT 41.505 -58.945 41.645 -58.775 ;
      RECT 41.555 -57.74 41.645 -56.732 ;
      RECT 41.505 -57.505 41.645 -57.335 ;
      RECT 41.555 -56.318 41.645 -55.31 ;
      RECT 41.505 -55.715 41.645 -55.545 ;
      RECT 41.555 -54.51 41.645 -53.502 ;
      RECT 41.505 -54.275 41.645 -54.105 ;
      RECT 41.555 -53.088 41.645 -52.08 ;
      RECT 41.505 -52.485 41.645 -52.315 ;
      RECT 41.555 -51.28 41.645 -50.272 ;
      RECT 41.505 -51.045 41.645 -50.875 ;
      RECT 41.555 -49.858 41.645 -48.85 ;
      RECT 41.505 -49.255 41.645 -49.085 ;
      RECT 41.555 -48.05 41.645 -47.042 ;
      RECT 41.505 -47.815 41.645 -47.645 ;
      RECT 41.555 -46.628 41.645 -45.62 ;
      RECT 41.505 -46.025 41.645 -45.855 ;
      RECT 41.555 -44.82 41.645 -43.812 ;
      RECT 41.505 -44.585 41.645 -44.415 ;
      RECT 41.555 -43.398 41.645 -42.39 ;
      RECT 41.505 -42.795 41.645 -42.625 ;
      RECT 41.555 -41.59 41.645 -40.582 ;
      RECT 41.505 -41.355 41.645 -41.185 ;
      RECT 41.555 -40.168 41.645 -39.16 ;
      RECT 41.505 -39.565 41.645 -39.395 ;
      RECT 41.555 -38.36 41.645 -37.352 ;
      RECT 41.505 -38.125 41.645 -37.955 ;
      RECT 41.555 -36.938 41.645 -35.93 ;
      RECT 41.505 -36.335 41.645 -36.165 ;
      RECT 41.555 -35.13 41.645 -34.122 ;
      RECT 41.505 -34.895 41.645 -34.725 ;
      RECT 41.555 -33.708 41.645 -32.7 ;
      RECT 41.505 -33.105 41.645 -32.935 ;
      RECT 41.555 -31.9 41.645 -30.892 ;
      RECT 41.505 -31.665 41.645 -31.495 ;
      RECT 41.555 -30.478 41.645 -29.47 ;
      RECT 41.505 -29.875 41.645 -29.705 ;
      RECT 41.555 -28.67 41.645 -27.662 ;
      RECT 41.505 -28.435 41.645 -28.265 ;
      RECT 41.555 -27.248 41.645 -26.24 ;
      RECT 41.505 -26.645 41.645 -26.475 ;
      RECT 41.555 -25.44 41.645 -24.432 ;
      RECT 41.505 -25.205 41.645 -25.035 ;
      RECT 41.555 -24.018 41.645 -23.01 ;
      RECT 41.505 -23.415 41.645 -23.245 ;
      RECT 41.555 -22.21 41.645 -21.202 ;
      RECT 41.505 -21.975 41.645 -21.805 ;
      RECT 41.555 -20.788 41.645 -19.78 ;
      RECT 41.505 -20.185 41.645 -20.015 ;
      RECT 41.555 -18.98 41.645 -17.972 ;
      RECT 41.505 -18.745 41.645 -18.575 ;
      RECT 41.555 -17.558 41.645 -16.55 ;
      RECT 41.505 -16.955 41.645 -16.785 ;
      RECT 41.555 -15.75 41.645 -14.742 ;
      RECT 41.505 -15.515 41.645 -15.345 ;
      RECT 41.555 -14.328 41.645 -13.32 ;
      RECT 41.505 -13.725 41.645 -13.555 ;
      RECT 41.555 -12.52 41.645 -11.512 ;
      RECT 41.505 -12.285 41.645 -12.115 ;
      RECT 41.555 -11.098 41.645 -10.09 ;
      RECT 41.505 -10.495 41.645 -10.325 ;
      RECT 41.555 -9.29 41.645 -8.282 ;
      RECT 41.505 -9.055 41.645 -8.885 ;
      RECT 41.555 -7.868 41.645 -6.86 ;
      RECT 41.505 -7.265 41.645 -7.095 ;
      RECT 41.555 -6.06 41.645 -5.052 ;
      RECT 41.505 -5.825 41.645 -5.655 ;
      RECT 41.555 -4.638 41.645 -3.63 ;
      RECT 41.505 -4.035 41.645 -3.865 ;
      RECT 41.555 -2.83 41.645 -1.822 ;
      RECT 41.505 -2.595 41.645 -2.425 ;
      RECT 41.555 -1.408 41.645 -0.4 ;
      RECT 41.505 -0.805 41.645 -0.635 ;
      RECT 41.555 0.4 41.645 1.408 ;
      RECT 41.505 0.635 41.645 0.805 ;
      RECT 41.155 -101.538 41.245 -100.531 ;
      RECT 41.155 -101.225 41.295 -101.055 ;
      RECT 41.155 -99.729 41.245 -98.722 ;
      RECT 41.155 -99.205 41.295 -99.035 ;
      RECT 41.155 -98.308 41.245 -97.301 ;
      RECT 41.155 -97.995 41.295 -97.825 ;
      RECT 41.155 -96.499 41.245 -95.492 ;
      RECT 41.155 -95.975 41.295 -95.805 ;
      RECT 41.155 -95.078 41.245 -94.071 ;
      RECT 41.155 -94.765 41.295 -94.595 ;
      RECT 41.155 -93.269 41.245 -92.262 ;
      RECT 41.155 -92.745 41.295 -92.575 ;
      RECT 41.155 -91.848 41.245 -90.841 ;
      RECT 41.155 -91.535 41.295 -91.365 ;
      RECT 41.155 -90.039 41.245 -89.032 ;
      RECT 41.155 -89.515 41.295 -89.345 ;
      RECT 41.155 -88.618 41.245 -87.611 ;
      RECT 41.155 -88.305 41.295 -88.135 ;
      RECT 41.155 -86.809 41.245 -85.802 ;
      RECT 41.155 -86.285 41.295 -86.115 ;
      RECT 41.155 -85.388 41.245 -84.381 ;
      RECT 41.155 -85.075 41.295 -84.905 ;
      RECT 41.155 -83.579 41.245 -82.572 ;
      RECT 41.155 -83.055 41.295 -82.885 ;
      RECT 41.155 -82.158 41.245 -81.151 ;
      RECT 41.155 -81.845 41.295 -81.675 ;
      RECT 41.155 -80.349 41.245 -79.342 ;
      RECT 41.155 -79.825 41.295 -79.655 ;
      RECT 41.155 -78.928 41.245 -77.921 ;
      RECT 41.155 -78.615 41.295 -78.445 ;
      RECT 41.155 -77.119 41.245 -76.112 ;
      RECT 41.155 -76.595 41.295 -76.425 ;
      RECT 41.155 -75.698 41.245 -74.691 ;
      RECT 41.155 -75.385 41.295 -75.215 ;
      RECT 41.155 -73.889 41.245 -72.882 ;
      RECT 41.155 -73.365 41.295 -73.195 ;
      RECT 41.155 -72.468 41.245 -71.461 ;
      RECT 41.155 -72.155 41.295 -71.985 ;
      RECT 41.155 -70.659 41.245 -69.652 ;
      RECT 41.155 -70.135 41.295 -69.965 ;
      RECT 41.155 -69.238 41.245 -68.231 ;
      RECT 41.155 -68.925 41.295 -68.755 ;
      RECT 41.155 -67.429 41.245 -66.422 ;
      RECT 41.155 -66.905 41.295 -66.735 ;
      RECT 41.155 -66.008 41.245 -65.001 ;
      RECT 41.155 -65.695 41.295 -65.525 ;
      RECT 41.155 -64.199 41.245 -63.192 ;
      RECT 41.155 -63.675 41.295 -63.505 ;
      RECT 41.155 -62.778 41.245 -61.771 ;
      RECT 41.155 -62.465 41.295 -62.295 ;
      RECT 41.155 -60.969 41.245 -59.962 ;
      RECT 41.155 -60.445 41.295 -60.275 ;
      RECT 41.155 -59.548 41.245 -58.541 ;
      RECT 41.155 -59.235 41.295 -59.065 ;
      RECT 41.155 -57.739 41.245 -56.732 ;
      RECT 41.155 -57.215 41.295 -57.045 ;
      RECT 41.155 -56.318 41.245 -55.311 ;
      RECT 41.155 -56.005 41.295 -55.835 ;
      RECT 41.155 -54.509 41.245 -53.502 ;
      RECT 41.155 -53.985 41.295 -53.815 ;
      RECT 41.155 -53.088 41.245 -52.081 ;
      RECT 41.155 -52.775 41.295 -52.605 ;
      RECT 41.155 -51.279 41.245 -50.272 ;
      RECT 41.155 -50.755 41.295 -50.585 ;
      RECT 41.155 -49.858 41.245 -48.851 ;
      RECT 41.155 -49.545 41.295 -49.375 ;
      RECT 41.155 -48.049 41.245 -47.042 ;
      RECT 41.155 -47.525 41.295 -47.355 ;
      RECT 41.155 -46.628 41.245 -45.621 ;
      RECT 41.155 -46.315 41.295 -46.145 ;
      RECT 41.155 -44.819 41.245 -43.812 ;
      RECT 41.155 -44.295 41.295 -44.125 ;
      RECT 41.155 -43.398 41.245 -42.391 ;
      RECT 41.155 -43.085 41.295 -42.915 ;
      RECT 41.155 -41.589 41.245 -40.582 ;
      RECT 41.155 -41.065 41.295 -40.895 ;
      RECT 41.155 -40.168 41.245 -39.161 ;
      RECT 41.155 -39.855 41.295 -39.685 ;
      RECT 41.155 -38.359 41.245 -37.352 ;
      RECT 41.155 -37.835 41.295 -37.665 ;
      RECT 41.155 -36.938 41.245 -35.931 ;
      RECT 41.155 -36.625 41.295 -36.455 ;
      RECT 41.155 -35.129 41.245 -34.122 ;
      RECT 41.155 -34.605 41.295 -34.435 ;
      RECT 41.155 -33.708 41.245 -32.701 ;
      RECT 41.155 -33.395 41.295 -33.225 ;
      RECT 41.155 -31.899 41.245 -30.892 ;
      RECT 41.155 -31.375 41.295 -31.205 ;
      RECT 41.155 -30.478 41.245 -29.471 ;
      RECT 41.155 -30.165 41.295 -29.995 ;
      RECT 41.155 -28.669 41.245 -27.662 ;
      RECT 41.155 -28.145 41.295 -27.975 ;
      RECT 41.155 -27.248 41.245 -26.241 ;
      RECT 41.155 -26.935 41.295 -26.765 ;
      RECT 41.155 -25.439 41.245 -24.432 ;
      RECT 41.155 -24.915 41.295 -24.745 ;
      RECT 41.155 -24.018 41.245 -23.011 ;
      RECT 41.155 -23.705 41.295 -23.535 ;
      RECT 41.155 -22.209 41.245 -21.202 ;
      RECT 41.155 -21.685 41.295 -21.515 ;
      RECT 41.155 -20.788 41.245 -19.781 ;
      RECT 41.155 -20.475 41.295 -20.305 ;
      RECT 41.155 -18.979 41.245 -17.972 ;
      RECT 41.155 -18.455 41.295 -18.285 ;
      RECT 41.155 -17.558 41.245 -16.551 ;
      RECT 41.155 -17.245 41.295 -17.075 ;
      RECT 41.155 -15.749 41.245 -14.742 ;
      RECT 41.155 -15.225 41.295 -15.055 ;
      RECT 41.155 -14.328 41.245 -13.321 ;
      RECT 41.155 -14.015 41.295 -13.845 ;
      RECT 41.155 -12.519 41.245 -11.512 ;
      RECT 41.155 -11.995 41.295 -11.825 ;
      RECT 41.155 -11.098 41.245 -10.091 ;
      RECT 41.155 -10.785 41.295 -10.615 ;
      RECT 41.155 -9.289 41.245 -8.282 ;
      RECT 41.155 -8.765 41.295 -8.595 ;
      RECT 41.155 -7.868 41.245 -6.861 ;
      RECT 41.155 -7.555 41.295 -7.385 ;
      RECT 41.155 -6.059 41.245 -5.052 ;
      RECT 41.155 -5.535 41.295 -5.365 ;
      RECT 41.155 -4.638 41.245 -3.631 ;
      RECT 41.155 -4.325 41.295 -4.155 ;
      RECT 41.155 -2.829 41.245 -1.822 ;
      RECT 41.155 -2.305 41.295 -2.135 ;
      RECT 41.155 -1.408 41.245 -0.401 ;
      RECT 41.155 -1.095 41.295 -0.925 ;
      RECT 41.155 0.401 41.245 1.408 ;
      RECT 41.155 0.925 41.295 1.095 ;
      RECT 39.305 -111.685 40.785 -111.585 ;
      RECT 39.305 -112.055 39.405 -111.585 ;
      RECT 39.11 -114.395 40.685 -114.275 ;
      RECT 40.585 -114.895 40.685 -114.275 ;
      RECT 39.99 -114.895 40.09 -114.275 ;
      RECT 39.11 -114.85 39.21 -114.275 ;
      RECT 40.355 -101.538 40.445 -100.53 ;
      RECT 40.305 -100.935 40.445 -100.765 ;
      RECT 40.355 -99.73 40.445 -98.722 ;
      RECT 40.305 -99.495 40.445 -99.325 ;
      RECT 40.355 -98.308 40.445 -97.3 ;
      RECT 40.305 -97.705 40.445 -97.535 ;
      RECT 40.355 -96.5 40.445 -95.492 ;
      RECT 40.305 -96.265 40.445 -96.095 ;
      RECT 40.355 -95.078 40.445 -94.07 ;
      RECT 40.305 -94.475 40.445 -94.305 ;
      RECT 40.355 -93.27 40.445 -92.262 ;
      RECT 40.305 -93.035 40.445 -92.865 ;
      RECT 40.355 -91.848 40.445 -90.84 ;
      RECT 40.305 -91.245 40.445 -91.075 ;
      RECT 40.355 -90.04 40.445 -89.032 ;
      RECT 40.305 -89.805 40.445 -89.635 ;
      RECT 40.355 -88.618 40.445 -87.61 ;
      RECT 40.305 -88.015 40.445 -87.845 ;
      RECT 40.355 -86.81 40.445 -85.802 ;
      RECT 40.305 -86.575 40.445 -86.405 ;
      RECT 40.355 -85.388 40.445 -84.38 ;
      RECT 40.305 -84.785 40.445 -84.615 ;
      RECT 40.355 -83.58 40.445 -82.572 ;
      RECT 40.305 -83.345 40.445 -83.175 ;
      RECT 40.355 -82.158 40.445 -81.15 ;
      RECT 40.305 -81.555 40.445 -81.385 ;
      RECT 40.355 -80.35 40.445 -79.342 ;
      RECT 40.305 -80.115 40.445 -79.945 ;
      RECT 40.355 -78.928 40.445 -77.92 ;
      RECT 40.305 -78.325 40.445 -78.155 ;
      RECT 40.355 -77.12 40.445 -76.112 ;
      RECT 40.305 -76.885 40.445 -76.715 ;
      RECT 40.355 -75.698 40.445 -74.69 ;
      RECT 40.305 -75.095 40.445 -74.925 ;
      RECT 40.355 -73.89 40.445 -72.882 ;
      RECT 40.305 -73.655 40.445 -73.485 ;
      RECT 40.355 -72.468 40.445 -71.46 ;
      RECT 40.305 -71.865 40.445 -71.695 ;
      RECT 40.355 -70.66 40.445 -69.652 ;
      RECT 40.305 -70.425 40.445 -70.255 ;
      RECT 40.355 -69.238 40.445 -68.23 ;
      RECT 40.305 -68.635 40.445 -68.465 ;
      RECT 40.355 -67.43 40.445 -66.422 ;
      RECT 40.305 -67.195 40.445 -67.025 ;
      RECT 40.355 -66.008 40.445 -65 ;
      RECT 40.305 -65.405 40.445 -65.235 ;
      RECT 40.355 -64.2 40.445 -63.192 ;
      RECT 40.305 -63.965 40.445 -63.795 ;
      RECT 40.355 -62.778 40.445 -61.77 ;
      RECT 40.305 -62.175 40.445 -62.005 ;
      RECT 40.355 -60.97 40.445 -59.962 ;
      RECT 40.305 -60.735 40.445 -60.565 ;
      RECT 40.355 -59.548 40.445 -58.54 ;
      RECT 40.305 -58.945 40.445 -58.775 ;
      RECT 40.355 -57.74 40.445 -56.732 ;
      RECT 40.305 -57.505 40.445 -57.335 ;
      RECT 40.355 -56.318 40.445 -55.31 ;
      RECT 40.305 -55.715 40.445 -55.545 ;
      RECT 40.355 -54.51 40.445 -53.502 ;
      RECT 40.305 -54.275 40.445 -54.105 ;
      RECT 40.355 -53.088 40.445 -52.08 ;
      RECT 40.305 -52.485 40.445 -52.315 ;
      RECT 40.355 -51.28 40.445 -50.272 ;
      RECT 40.305 -51.045 40.445 -50.875 ;
      RECT 40.355 -49.858 40.445 -48.85 ;
      RECT 40.305 -49.255 40.445 -49.085 ;
      RECT 40.355 -48.05 40.445 -47.042 ;
      RECT 40.305 -47.815 40.445 -47.645 ;
      RECT 40.355 -46.628 40.445 -45.62 ;
      RECT 40.305 -46.025 40.445 -45.855 ;
      RECT 40.355 -44.82 40.445 -43.812 ;
      RECT 40.305 -44.585 40.445 -44.415 ;
      RECT 40.355 -43.398 40.445 -42.39 ;
      RECT 40.305 -42.795 40.445 -42.625 ;
      RECT 40.355 -41.59 40.445 -40.582 ;
      RECT 40.305 -41.355 40.445 -41.185 ;
      RECT 40.355 -40.168 40.445 -39.16 ;
      RECT 40.305 -39.565 40.445 -39.395 ;
      RECT 40.355 -38.36 40.445 -37.352 ;
      RECT 40.305 -38.125 40.445 -37.955 ;
      RECT 40.355 -36.938 40.445 -35.93 ;
      RECT 40.305 -36.335 40.445 -36.165 ;
      RECT 40.355 -35.13 40.445 -34.122 ;
      RECT 40.305 -34.895 40.445 -34.725 ;
      RECT 40.355 -33.708 40.445 -32.7 ;
      RECT 40.305 -33.105 40.445 -32.935 ;
      RECT 40.355 -31.9 40.445 -30.892 ;
      RECT 40.305 -31.665 40.445 -31.495 ;
      RECT 40.355 -30.478 40.445 -29.47 ;
      RECT 40.305 -29.875 40.445 -29.705 ;
      RECT 40.355 -28.67 40.445 -27.662 ;
      RECT 40.305 -28.435 40.445 -28.265 ;
      RECT 40.355 -27.248 40.445 -26.24 ;
      RECT 40.305 -26.645 40.445 -26.475 ;
      RECT 40.355 -25.44 40.445 -24.432 ;
      RECT 40.305 -25.205 40.445 -25.035 ;
      RECT 40.355 -24.018 40.445 -23.01 ;
      RECT 40.305 -23.415 40.445 -23.245 ;
      RECT 40.355 -22.21 40.445 -21.202 ;
      RECT 40.305 -21.975 40.445 -21.805 ;
      RECT 40.355 -20.788 40.445 -19.78 ;
      RECT 40.305 -20.185 40.445 -20.015 ;
      RECT 40.355 -18.98 40.445 -17.972 ;
      RECT 40.305 -18.745 40.445 -18.575 ;
      RECT 40.355 -17.558 40.445 -16.55 ;
      RECT 40.305 -16.955 40.445 -16.785 ;
      RECT 40.355 -15.75 40.445 -14.742 ;
      RECT 40.305 -15.515 40.445 -15.345 ;
      RECT 40.355 -14.328 40.445 -13.32 ;
      RECT 40.305 -13.725 40.445 -13.555 ;
      RECT 40.355 -12.52 40.445 -11.512 ;
      RECT 40.305 -12.285 40.445 -12.115 ;
      RECT 40.355 -11.098 40.445 -10.09 ;
      RECT 40.305 -10.495 40.445 -10.325 ;
      RECT 40.355 -9.29 40.445 -8.282 ;
      RECT 40.305 -9.055 40.445 -8.885 ;
      RECT 40.355 -7.868 40.445 -6.86 ;
      RECT 40.305 -7.265 40.445 -7.095 ;
      RECT 40.355 -6.06 40.445 -5.052 ;
      RECT 40.305 -5.825 40.445 -5.655 ;
      RECT 40.355 -4.638 40.445 -3.63 ;
      RECT 40.305 -4.035 40.445 -3.865 ;
      RECT 40.355 -2.83 40.445 -1.822 ;
      RECT 40.305 -2.595 40.445 -2.425 ;
      RECT 40.355 -1.408 40.445 -0.4 ;
      RECT 40.305 -0.805 40.445 -0.635 ;
      RECT 40.355 0.4 40.445 1.408 ;
      RECT 40.305 0.635 40.445 0.805 ;
      RECT 40.23 -114.685 40.405 -114.515 ;
      RECT 40.305 -114.895 40.405 -114.515 ;
      RECT 39.345 -113.555 39.445 -113.09 ;
      RECT 39.71 -113.555 39.81 -113.1 ;
      RECT 39.345 -113.555 40.19 -113.385 ;
      RECT 39.955 -101.538 40.045 -100.531 ;
      RECT 39.955 -101.225 40.095 -101.055 ;
      RECT 39.955 -99.729 40.045 -98.722 ;
      RECT 39.955 -99.205 40.095 -99.035 ;
      RECT 39.955 -98.308 40.045 -97.301 ;
      RECT 39.955 -97.995 40.095 -97.825 ;
      RECT 39.955 -96.499 40.045 -95.492 ;
      RECT 39.955 -95.975 40.095 -95.805 ;
      RECT 39.955 -95.078 40.045 -94.071 ;
      RECT 39.955 -94.765 40.095 -94.595 ;
      RECT 39.955 -93.269 40.045 -92.262 ;
      RECT 39.955 -92.745 40.095 -92.575 ;
      RECT 39.955 -91.848 40.045 -90.841 ;
      RECT 39.955 -91.535 40.095 -91.365 ;
      RECT 39.955 -90.039 40.045 -89.032 ;
      RECT 39.955 -89.515 40.095 -89.345 ;
      RECT 39.955 -88.618 40.045 -87.611 ;
      RECT 39.955 -88.305 40.095 -88.135 ;
      RECT 39.955 -86.809 40.045 -85.802 ;
      RECT 39.955 -86.285 40.095 -86.115 ;
      RECT 39.955 -85.388 40.045 -84.381 ;
      RECT 39.955 -85.075 40.095 -84.905 ;
      RECT 39.955 -83.579 40.045 -82.572 ;
      RECT 39.955 -83.055 40.095 -82.885 ;
      RECT 39.955 -82.158 40.045 -81.151 ;
      RECT 39.955 -81.845 40.095 -81.675 ;
      RECT 39.955 -80.349 40.045 -79.342 ;
      RECT 39.955 -79.825 40.095 -79.655 ;
      RECT 39.955 -78.928 40.045 -77.921 ;
      RECT 39.955 -78.615 40.095 -78.445 ;
      RECT 39.955 -77.119 40.045 -76.112 ;
      RECT 39.955 -76.595 40.095 -76.425 ;
      RECT 39.955 -75.698 40.045 -74.691 ;
      RECT 39.955 -75.385 40.095 -75.215 ;
      RECT 39.955 -73.889 40.045 -72.882 ;
      RECT 39.955 -73.365 40.095 -73.195 ;
      RECT 39.955 -72.468 40.045 -71.461 ;
      RECT 39.955 -72.155 40.095 -71.985 ;
      RECT 39.955 -70.659 40.045 -69.652 ;
      RECT 39.955 -70.135 40.095 -69.965 ;
      RECT 39.955 -69.238 40.045 -68.231 ;
      RECT 39.955 -68.925 40.095 -68.755 ;
      RECT 39.955 -67.429 40.045 -66.422 ;
      RECT 39.955 -66.905 40.095 -66.735 ;
      RECT 39.955 -66.008 40.045 -65.001 ;
      RECT 39.955 -65.695 40.095 -65.525 ;
      RECT 39.955 -64.199 40.045 -63.192 ;
      RECT 39.955 -63.675 40.095 -63.505 ;
      RECT 39.955 -62.778 40.045 -61.771 ;
      RECT 39.955 -62.465 40.095 -62.295 ;
      RECT 39.955 -60.969 40.045 -59.962 ;
      RECT 39.955 -60.445 40.095 -60.275 ;
      RECT 39.955 -59.548 40.045 -58.541 ;
      RECT 39.955 -59.235 40.095 -59.065 ;
      RECT 39.955 -57.739 40.045 -56.732 ;
      RECT 39.955 -57.215 40.095 -57.045 ;
      RECT 39.955 -56.318 40.045 -55.311 ;
      RECT 39.955 -56.005 40.095 -55.835 ;
      RECT 39.955 -54.509 40.045 -53.502 ;
      RECT 39.955 -53.985 40.095 -53.815 ;
      RECT 39.955 -53.088 40.045 -52.081 ;
      RECT 39.955 -52.775 40.095 -52.605 ;
      RECT 39.955 -51.279 40.045 -50.272 ;
      RECT 39.955 -50.755 40.095 -50.585 ;
      RECT 39.955 -49.858 40.045 -48.851 ;
      RECT 39.955 -49.545 40.095 -49.375 ;
      RECT 39.955 -48.049 40.045 -47.042 ;
      RECT 39.955 -47.525 40.095 -47.355 ;
      RECT 39.955 -46.628 40.045 -45.621 ;
      RECT 39.955 -46.315 40.095 -46.145 ;
      RECT 39.955 -44.819 40.045 -43.812 ;
      RECT 39.955 -44.295 40.095 -44.125 ;
      RECT 39.955 -43.398 40.045 -42.391 ;
      RECT 39.955 -43.085 40.095 -42.915 ;
      RECT 39.955 -41.589 40.045 -40.582 ;
      RECT 39.955 -41.065 40.095 -40.895 ;
      RECT 39.955 -40.168 40.045 -39.161 ;
      RECT 39.955 -39.855 40.095 -39.685 ;
      RECT 39.955 -38.359 40.045 -37.352 ;
      RECT 39.955 -37.835 40.095 -37.665 ;
      RECT 39.955 -36.938 40.045 -35.931 ;
      RECT 39.955 -36.625 40.095 -36.455 ;
      RECT 39.955 -35.129 40.045 -34.122 ;
      RECT 39.955 -34.605 40.095 -34.435 ;
      RECT 39.955 -33.708 40.045 -32.701 ;
      RECT 39.955 -33.395 40.095 -33.225 ;
      RECT 39.955 -31.899 40.045 -30.892 ;
      RECT 39.955 -31.375 40.095 -31.205 ;
      RECT 39.955 -30.478 40.045 -29.471 ;
      RECT 39.955 -30.165 40.095 -29.995 ;
      RECT 39.955 -28.669 40.045 -27.662 ;
      RECT 39.955 -28.145 40.095 -27.975 ;
      RECT 39.955 -27.248 40.045 -26.241 ;
      RECT 39.955 -26.935 40.095 -26.765 ;
      RECT 39.955 -25.439 40.045 -24.432 ;
      RECT 39.955 -24.915 40.095 -24.745 ;
      RECT 39.955 -24.018 40.045 -23.011 ;
      RECT 39.955 -23.705 40.095 -23.535 ;
      RECT 39.955 -22.209 40.045 -21.202 ;
      RECT 39.955 -21.685 40.095 -21.515 ;
      RECT 39.955 -20.788 40.045 -19.781 ;
      RECT 39.955 -20.475 40.095 -20.305 ;
      RECT 39.955 -18.979 40.045 -17.972 ;
      RECT 39.955 -18.455 40.095 -18.285 ;
      RECT 39.955 -17.558 40.045 -16.551 ;
      RECT 39.955 -17.245 40.095 -17.075 ;
      RECT 39.955 -15.749 40.045 -14.742 ;
      RECT 39.955 -15.225 40.095 -15.055 ;
      RECT 39.955 -14.328 40.045 -13.321 ;
      RECT 39.955 -14.015 40.095 -13.845 ;
      RECT 39.955 -12.519 40.045 -11.512 ;
      RECT 39.955 -11.995 40.095 -11.825 ;
      RECT 39.955 -11.098 40.045 -10.091 ;
      RECT 39.955 -10.785 40.095 -10.615 ;
      RECT 39.955 -9.289 40.045 -8.282 ;
      RECT 39.955 -8.765 40.095 -8.595 ;
      RECT 39.955 -7.868 40.045 -6.861 ;
      RECT 39.955 -7.555 40.095 -7.385 ;
      RECT 39.955 -6.059 40.045 -5.052 ;
      RECT 39.955 -5.535 40.095 -5.365 ;
      RECT 39.955 -4.638 40.045 -3.631 ;
      RECT 39.955 -4.325 40.095 -4.155 ;
      RECT 39.955 -2.829 40.045 -1.822 ;
      RECT 39.955 -2.305 40.095 -2.135 ;
      RECT 39.955 -1.408 40.045 -0.401 ;
      RECT 39.955 -1.095 40.095 -0.925 ;
      RECT 39.955 0.401 40.045 1.408 ;
      RECT 39.955 0.925 40.095 1.095 ;
      RECT 39.64 -114.685 39.81 -114.515 ;
      RECT 39.71 -114.895 39.81 -114.515 ;
      RECT 39.155 -101.538 39.245 -100.53 ;
      RECT 39.105 -100.935 39.245 -100.765 ;
      RECT 39.155 -99.73 39.245 -98.722 ;
      RECT 39.105 -99.495 39.245 -99.325 ;
      RECT 39.155 -98.308 39.245 -97.3 ;
      RECT 39.105 -97.705 39.245 -97.535 ;
      RECT 39.155 -96.5 39.245 -95.492 ;
      RECT 39.105 -96.265 39.245 -96.095 ;
      RECT 39.155 -95.078 39.245 -94.07 ;
      RECT 39.105 -94.475 39.245 -94.305 ;
      RECT 39.155 -93.27 39.245 -92.262 ;
      RECT 39.105 -93.035 39.245 -92.865 ;
      RECT 39.155 -91.848 39.245 -90.84 ;
      RECT 39.105 -91.245 39.245 -91.075 ;
      RECT 39.155 -90.04 39.245 -89.032 ;
      RECT 39.105 -89.805 39.245 -89.635 ;
      RECT 39.155 -88.618 39.245 -87.61 ;
      RECT 39.105 -88.015 39.245 -87.845 ;
      RECT 39.155 -86.81 39.245 -85.802 ;
      RECT 39.105 -86.575 39.245 -86.405 ;
      RECT 39.155 -85.388 39.245 -84.38 ;
      RECT 39.105 -84.785 39.245 -84.615 ;
      RECT 39.155 -83.58 39.245 -82.572 ;
      RECT 39.105 -83.345 39.245 -83.175 ;
      RECT 39.155 -82.158 39.245 -81.15 ;
      RECT 39.105 -81.555 39.245 -81.385 ;
      RECT 39.155 -80.35 39.245 -79.342 ;
      RECT 39.105 -80.115 39.245 -79.945 ;
      RECT 39.155 -78.928 39.245 -77.92 ;
      RECT 39.105 -78.325 39.245 -78.155 ;
      RECT 39.155 -77.12 39.245 -76.112 ;
      RECT 39.105 -76.885 39.245 -76.715 ;
      RECT 39.155 -75.698 39.245 -74.69 ;
      RECT 39.105 -75.095 39.245 -74.925 ;
      RECT 39.155 -73.89 39.245 -72.882 ;
      RECT 39.105 -73.655 39.245 -73.485 ;
      RECT 39.155 -72.468 39.245 -71.46 ;
      RECT 39.105 -71.865 39.245 -71.695 ;
      RECT 39.155 -70.66 39.245 -69.652 ;
      RECT 39.105 -70.425 39.245 -70.255 ;
      RECT 39.155 -69.238 39.245 -68.23 ;
      RECT 39.105 -68.635 39.245 -68.465 ;
      RECT 39.155 -67.43 39.245 -66.422 ;
      RECT 39.105 -67.195 39.245 -67.025 ;
      RECT 39.155 -66.008 39.245 -65 ;
      RECT 39.105 -65.405 39.245 -65.235 ;
      RECT 39.155 -64.2 39.245 -63.192 ;
      RECT 39.105 -63.965 39.245 -63.795 ;
      RECT 39.155 -62.778 39.245 -61.77 ;
      RECT 39.105 -62.175 39.245 -62.005 ;
      RECT 39.155 -60.97 39.245 -59.962 ;
      RECT 39.105 -60.735 39.245 -60.565 ;
      RECT 39.155 -59.548 39.245 -58.54 ;
      RECT 39.105 -58.945 39.245 -58.775 ;
      RECT 39.155 -57.74 39.245 -56.732 ;
      RECT 39.105 -57.505 39.245 -57.335 ;
      RECT 39.155 -56.318 39.245 -55.31 ;
      RECT 39.105 -55.715 39.245 -55.545 ;
      RECT 39.155 -54.51 39.245 -53.502 ;
      RECT 39.105 -54.275 39.245 -54.105 ;
      RECT 39.155 -53.088 39.245 -52.08 ;
      RECT 39.105 -52.485 39.245 -52.315 ;
      RECT 39.155 -51.28 39.245 -50.272 ;
      RECT 39.105 -51.045 39.245 -50.875 ;
      RECT 39.155 -49.858 39.245 -48.85 ;
      RECT 39.105 -49.255 39.245 -49.085 ;
      RECT 39.155 -48.05 39.245 -47.042 ;
      RECT 39.105 -47.815 39.245 -47.645 ;
      RECT 39.155 -46.628 39.245 -45.62 ;
      RECT 39.105 -46.025 39.245 -45.855 ;
      RECT 39.155 -44.82 39.245 -43.812 ;
      RECT 39.105 -44.585 39.245 -44.415 ;
      RECT 39.155 -43.398 39.245 -42.39 ;
      RECT 39.105 -42.795 39.245 -42.625 ;
      RECT 39.155 -41.59 39.245 -40.582 ;
      RECT 39.105 -41.355 39.245 -41.185 ;
      RECT 39.155 -40.168 39.245 -39.16 ;
      RECT 39.105 -39.565 39.245 -39.395 ;
      RECT 39.155 -38.36 39.245 -37.352 ;
      RECT 39.105 -38.125 39.245 -37.955 ;
      RECT 39.155 -36.938 39.245 -35.93 ;
      RECT 39.105 -36.335 39.245 -36.165 ;
      RECT 39.155 -35.13 39.245 -34.122 ;
      RECT 39.105 -34.895 39.245 -34.725 ;
      RECT 39.155 -33.708 39.245 -32.7 ;
      RECT 39.105 -33.105 39.245 -32.935 ;
      RECT 39.155 -31.9 39.245 -30.892 ;
      RECT 39.105 -31.665 39.245 -31.495 ;
      RECT 39.155 -30.478 39.245 -29.47 ;
      RECT 39.105 -29.875 39.245 -29.705 ;
      RECT 39.155 -28.67 39.245 -27.662 ;
      RECT 39.105 -28.435 39.245 -28.265 ;
      RECT 39.155 -27.248 39.245 -26.24 ;
      RECT 39.105 -26.645 39.245 -26.475 ;
      RECT 39.155 -25.44 39.245 -24.432 ;
      RECT 39.105 -25.205 39.245 -25.035 ;
      RECT 39.155 -24.018 39.245 -23.01 ;
      RECT 39.105 -23.415 39.245 -23.245 ;
      RECT 39.155 -22.21 39.245 -21.202 ;
      RECT 39.105 -21.975 39.245 -21.805 ;
      RECT 39.155 -20.788 39.245 -19.78 ;
      RECT 39.105 -20.185 39.245 -20.015 ;
      RECT 39.155 -18.98 39.245 -17.972 ;
      RECT 39.105 -18.745 39.245 -18.575 ;
      RECT 39.155 -17.558 39.245 -16.55 ;
      RECT 39.105 -16.955 39.245 -16.785 ;
      RECT 39.155 -15.75 39.245 -14.742 ;
      RECT 39.105 -15.515 39.245 -15.345 ;
      RECT 39.155 -14.328 39.245 -13.32 ;
      RECT 39.105 -13.725 39.245 -13.555 ;
      RECT 39.155 -12.52 39.245 -11.512 ;
      RECT 39.105 -12.285 39.245 -12.115 ;
      RECT 39.155 -11.098 39.245 -10.09 ;
      RECT 39.105 -10.495 39.245 -10.325 ;
      RECT 39.155 -9.29 39.245 -8.282 ;
      RECT 39.105 -9.055 39.245 -8.885 ;
      RECT 39.155 -7.868 39.245 -6.86 ;
      RECT 39.105 -7.265 39.245 -7.095 ;
      RECT 39.155 -6.06 39.245 -5.052 ;
      RECT 39.105 -5.825 39.245 -5.655 ;
      RECT 39.155 -4.638 39.245 -3.63 ;
      RECT 39.105 -4.035 39.245 -3.865 ;
      RECT 39.155 -2.83 39.245 -1.822 ;
      RECT 39.105 -2.595 39.245 -2.425 ;
      RECT 39.155 -1.408 39.245 -0.4 ;
      RECT 39.105 -0.805 39.245 -0.635 ;
      RECT 39.155 0.4 39.245 1.408 ;
      RECT 39.105 0.635 39.245 0.805 ;
      RECT 38.755 -101.538 38.845 -100.531 ;
      RECT 38.755 -101.225 38.895 -101.055 ;
      RECT 38.755 -99.729 38.845 -98.722 ;
      RECT 38.755 -99.205 38.895 -99.035 ;
      RECT 38.755 -98.308 38.845 -97.301 ;
      RECT 38.755 -97.995 38.895 -97.825 ;
      RECT 38.755 -96.499 38.845 -95.492 ;
      RECT 38.755 -95.975 38.895 -95.805 ;
      RECT 38.755 -95.078 38.845 -94.071 ;
      RECT 38.755 -94.765 38.895 -94.595 ;
      RECT 38.755 -93.269 38.845 -92.262 ;
      RECT 38.755 -92.745 38.895 -92.575 ;
      RECT 38.755 -91.848 38.845 -90.841 ;
      RECT 38.755 -91.535 38.895 -91.365 ;
      RECT 38.755 -90.039 38.845 -89.032 ;
      RECT 38.755 -89.515 38.895 -89.345 ;
      RECT 38.755 -88.618 38.845 -87.611 ;
      RECT 38.755 -88.305 38.895 -88.135 ;
      RECT 38.755 -86.809 38.845 -85.802 ;
      RECT 38.755 -86.285 38.895 -86.115 ;
      RECT 38.755 -85.388 38.845 -84.381 ;
      RECT 38.755 -85.075 38.895 -84.905 ;
      RECT 38.755 -83.579 38.845 -82.572 ;
      RECT 38.755 -83.055 38.895 -82.885 ;
      RECT 38.755 -82.158 38.845 -81.151 ;
      RECT 38.755 -81.845 38.895 -81.675 ;
      RECT 38.755 -80.349 38.845 -79.342 ;
      RECT 38.755 -79.825 38.895 -79.655 ;
      RECT 38.755 -78.928 38.845 -77.921 ;
      RECT 38.755 -78.615 38.895 -78.445 ;
      RECT 38.755 -77.119 38.845 -76.112 ;
      RECT 38.755 -76.595 38.895 -76.425 ;
      RECT 38.755 -75.698 38.845 -74.691 ;
      RECT 38.755 -75.385 38.895 -75.215 ;
      RECT 38.755 -73.889 38.845 -72.882 ;
      RECT 38.755 -73.365 38.895 -73.195 ;
      RECT 38.755 -72.468 38.845 -71.461 ;
      RECT 38.755 -72.155 38.895 -71.985 ;
      RECT 38.755 -70.659 38.845 -69.652 ;
      RECT 38.755 -70.135 38.895 -69.965 ;
      RECT 38.755 -69.238 38.845 -68.231 ;
      RECT 38.755 -68.925 38.895 -68.755 ;
      RECT 38.755 -67.429 38.845 -66.422 ;
      RECT 38.755 -66.905 38.895 -66.735 ;
      RECT 38.755 -66.008 38.845 -65.001 ;
      RECT 38.755 -65.695 38.895 -65.525 ;
      RECT 38.755 -64.199 38.845 -63.192 ;
      RECT 38.755 -63.675 38.895 -63.505 ;
      RECT 38.755 -62.778 38.845 -61.771 ;
      RECT 38.755 -62.465 38.895 -62.295 ;
      RECT 38.755 -60.969 38.845 -59.962 ;
      RECT 38.755 -60.445 38.895 -60.275 ;
      RECT 38.755 -59.548 38.845 -58.541 ;
      RECT 38.755 -59.235 38.895 -59.065 ;
      RECT 38.755 -57.739 38.845 -56.732 ;
      RECT 38.755 -57.215 38.895 -57.045 ;
      RECT 38.755 -56.318 38.845 -55.311 ;
      RECT 38.755 -56.005 38.895 -55.835 ;
      RECT 38.755 -54.509 38.845 -53.502 ;
      RECT 38.755 -53.985 38.895 -53.815 ;
      RECT 38.755 -53.088 38.845 -52.081 ;
      RECT 38.755 -52.775 38.895 -52.605 ;
      RECT 38.755 -51.279 38.845 -50.272 ;
      RECT 38.755 -50.755 38.895 -50.585 ;
      RECT 38.755 -49.858 38.845 -48.851 ;
      RECT 38.755 -49.545 38.895 -49.375 ;
      RECT 38.755 -48.049 38.845 -47.042 ;
      RECT 38.755 -47.525 38.895 -47.355 ;
      RECT 38.755 -46.628 38.845 -45.621 ;
      RECT 38.755 -46.315 38.895 -46.145 ;
      RECT 38.755 -44.819 38.845 -43.812 ;
      RECT 38.755 -44.295 38.895 -44.125 ;
      RECT 38.755 -43.398 38.845 -42.391 ;
      RECT 38.755 -43.085 38.895 -42.915 ;
      RECT 38.755 -41.589 38.845 -40.582 ;
      RECT 38.755 -41.065 38.895 -40.895 ;
      RECT 38.755 -40.168 38.845 -39.161 ;
      RECT 38.755 -39.855 38.895 -39.685 ;
      RECT 38.755 -38.359 38.845 -37.352 ;
      RECT 38.755 -37.835 38.895 -37.665 ;
      RECT 38.755 -36.938 38.845 -35.931 ;
      RECT 38.755 -36.625 38.895 -36.455 ;
      RECT 38.755 -35.129 38.845 -34.122 ;
      RECT 38.755 -34.605 38.895 -34.435 ;
      RECT 38.755 -33.708 38.845 -32.701 ;
      RECT 38.755 -33.395 38.895 -33.225 ;
      RECT 38.755 -31.899 38.845 -30.892 ;
      RECT 38.755 -31.375 38.895 -31.205 ;
      RECT 38.755 -30.478 38.845 -29.471 ;
      RECT 38.755 -30.165 38.895 -29.995 ;
      RECT 38.755 -28.669 38.845 -27.662 ;
      RECT 38.755 -28.145 38.895 -27.975 ;
      RECT 38.755 -27.248 38.845 -26.241 ;
      RECT 38.755 -26.935 38.895 -26.765 ;
      RECT 38.755 -25.439 38.845 -24.432 ;
      RECT 38.755 -24.915 38.895 -24.745 ;
      RECT 38.755 -24.018 38.845 -23.011 ;
      RECT 38.755 -23.705 38.895 -23.535 ;
      RECT 38.755 -22.209 38.845 -21.202 ;
      RECT 38.755 -21.685 38.895 -21.515 ;
      RECT 38.755 -20.788 38.845 -19.781 ;
      RECT 38.755 -20.475 38.895 -20.305 ;
      RECT 38.755 -18.979 38.845 -17.972 ;
      RECT 38.755 -18.455 38.895 -18.285 ;
      RECT 38.755 -17.558 38.845 -16.551 ;
      RECT 38.755 -17.245 38.895 -17.075 ;
      RECT 38.755 -15.749 38.845 -14.742 ;
      RECT 38.755 -15.225 38.895 -15.055 ;
      RECT 38.755 -14.328 38.845 -13.321 ;
      RECT 38.755 -14.015 38.895 -13.845 ;
      RECT 38.755 -12.519 38.845 -11.512 ;
      RECT 38.755 -11.995 38.895 -11.825 ;
      RECT 38.755 -11.098 38.845 -10.091 ;
      RECT 38.755 -10.785 38.895 -10.615 ;
      RECT 38.755 -9.289 38.845 -8.282 ;
      RECT 38.755 -8.765 38.895 -8.595 ;
      RECT 38.755 -7.868 38.845 -6.861 ;
      RECT 38.755 -7.555 38.895 -7.385 ;
      RECT 38.755 -6.059 38.845 -5.052 ;
      RECT 38.755 -5.535 38.895 -5.365 ;
      RECT 38.755 -4.638 38.845 -3.631 ;
      RECT 38.755 -4.325 38.895 -4.155 ;
      RECT 38.755 -2.829 38.845 -1.822 ;
      RECT 38.755 -2.305 38.895 -2.135 ;
      RECT 38.755 -1.408 38.845 -0.401 ;
      RECT 38.755 -1.095 38.895 -0.925 ;
      RECT 38.755 0.401 38.845 1.408 ;
      RECT 38.755 0.925 38.895 1.095 ;
      RECT 34.585 -108.935 38.365 -108.815 ;
      RECT 35.905 -109.475 36.005 -108.815 ;
      RECT 35.345 -109.475 35.445 -108.815 ;
      RECT 34.785 -109.475 34.885 -108.815 ;
      RECT 37.955 -101.538 38.045 -100.53 ;
      RECT 37.905 -100.935 38.045 -100.765 ;
      RECT 37.955 -99.73 38.045 -98.722 ;
      RECT 37.905 -99.495 38.045 -99.325 ;
      RECT 37.955 -98.308 38.045 -97.3 ;
      RECT 37.905 -97.705 38.045 -97.535 ;
      RECT 37.955 -96.5 38.045 -95.492 ;
      RECT 37.905 -96.265 38.045 -96.095 ;
      RECT 37.955 -95.078 38.045 -94.07 ;
      RECT 37.905 -94.475 38.045 -94.305 ;
      RECT 37.955 -93.27 38.045 -92.262 ;
      RECT 37.905 -93.035 38.045 -92.865 ;
      RECT 37.955 -91.848 38.045 -90.84 ;
      RECT 37.905 -91.245 38.045 -91.075 ;
      RECT 37.955 -90.04 38.045 -89.032 ;
      RECT 37.905 -89.805 38.045 -89.635 ;
      RECT 37.955 -88.618 38.045 -87.61 ;
      RECT 37.905 -88.015 38.045 -87.845 ;
      RECT 37.955 -86.81 38.045 -85.802 ;
      RECT 37.905 -86.575 38.045 -86.405 ;
      RECT 37.955 -85.388 38.045 -84.38 ;
      RECT 37.905 -84.785 38.045 -84.615 ;
      RECT 37.955 -83.58 38.045 -82.572 ;
      RECT 37.905 -83.345 38.045 -83.175 ;
      RECT 37.955 -82.158 38.045 -81.15 ;
      RECT 37.905 -81.555 38.045 -81.385 ;
      RECT 37.955 -80.35 38.045 -79.342 ;
      RECT 37.905 -80.115 38.045 -79.945 ;
      RECT 37.955 -78.928 38.045 -77.92 ;
      RECT 37.905 -78.325 38.045 -78.155 ;
      RECT 37.955 -77.12 38.045 -76.112 ;
      RECT 37.905 -76.885 38.045 -76.715 ;
      RECT 37.955 -75.698 38.045 -74.69 ;
      RECT 37.905 -75.095 38.045 -74.925 ;
      RECT 37.955 -73.89 38.045 -72.882 ;
      RECT 37.905 -73.655 38.045 -73.485 ;
      RECT 37.955 -72.468 38.045 -71.46 ;
      RECT 37.905 -71.865 38.045 -71.695 ;
      RECT 37.955 -70.66 38.045 -69.652 ;
      RECT 37.905 -70.425 38.045 -70.255 ;
      RECT 37.955 -69.238 38.045 -68.23 ;
      RECT 37.905 -68.635 38.045 -68.465 ;
      RECT 37.955 -67.43 38.045 -66.422 ;
      RECT 37.905 -67.195 38.045 -67.025 ;
      RECT 37.955 -66.008 38.045 -65 ;
      RECT 37.905 -65.405 38.045 -65.235 ;
      RECT 37.955 -64.2 38.045 -63.192 ;
      RECT 37.905 -63.965 38.045 -63.795 ;
      RECT 37.955 -62.778 38.045 -61.77 ;
      RECT 37.905 -62.175 38.045 -62.005 ;
      RECT 37.955 -60.97 38.045 -59.962 ;
      RECT 37.905 -60.735 38.045 -60.565 ;
      RECT 37.955 -59.548 38.045 -58.54 ;
      RECT 37.905 -58.945 38.045 -58.775 ;
      RECT 37.955 -57.74 38.045 -56.732 ;
      RECT 37.905 -57.505 38.045 -57.335 ;
      RECT 37.955 -56.318 38.045 -55.31 ;
      RECT 37.905 -55.715 38.045 -55.545 ;
      RECT 37.955 -54.51 38.045 -53.502 ;
      RECT 37.905 -54.275 38.045 -54.105 ;
      RECT 37.955 -53.088 38.045 -52.08 ;
      RECT 37.905 -52.485 38.045 -52.315 ;
      RECT 37.955 -51.28 38.045 -50.272 ;
      RECT 37.905 -51.045 38.045 -50.875 ;
      RECT 37.955 -49.858 38.045 -48.85 ;
      RECT 37.905 -49.255 38.045 -49.085 ;
      RECT 37.955 -48.05 38.045 -47.042 ;
      RECT 37.905 -47.815 38.045 -47.645 ;
      RECT 37.955 -46.628 38.045 -45.62 ;
      RECT 37.905 -46.025 38.045 -45.855 ;
      RECT 37.955 -44.82 38.045 -43.812 ;
      RECT 37.905 -44.585 38.045 -44.415 ;
      RECT 37.955 -43.398 38.045 -42.39 ;
      RECT 37.905 -42.795 38.045 -42.625 ;
      RECT 37.955 -41.59 38.045 -40.582 ;
      RECT 37.905 -41.355 38.045 -41.185 ;
      RECT 37.955 -40.168 38.045 -39.16 ;
      RECT 37.905 -39.565 38.045 -39.395 ;
      RECT 37.955 -38.36 38.045 -37.352 ;
      RECT 37.905 -38.125 38.045 -37.955 ;
      RECT 37.955 -36.938 38.045 -35.93 ;
      RECT 37.905 -36.335 38.045 -36.165 ;
      RECT 37.955 -35.13 38.045 -34.122 ;
      RECT 37.905 -34.895 38.045 -34.725 ;
      RECT 37.955 -33.708 38.045 -32.7 ;
      RECT 37.905 -33.105 38.045 -32.935 ;
      RECT 37.955 -31.9 38.045 -30.892 ;
      RECT 37.905 -31.665 38.045 -31.495 ;
      RECT 37.955 -30.478 38.045 -29.47 ;
      RECT 37.905 -29.875 38.045 -29.705 ;
      RECT 37.955 -28.67 38.045 -27.662 ;
      RECT 37.905 -28.435 38.045 -28.265 ;
      RECT 37.955 -27.248 38.045 -26.24 ;
      RECT 37.905 -26.645 38.045 -26.475 ;
      RECT 37.955 -25.44 38.045 -24.432 ;
      RECT 37.905 -25.205 38.045 -25.035 ;
      RECT 37.955 -24.018 38.045 -23.01 ;
      RECT 37.905 -23.415 38.045 -23.245 ;
      RECT 37.955 -22.21 38.045 -21.202 ;
      RECT 37.905 -21.975 38.045 -21.805 ;
      RECT 37.955 -20.788 38.045 -19.78 ;
      RECT 37.905 -20.185 38.045 -20.015 ;
      RECT 37.955 -18.98 38.045 -17.972 ;
      RECT 37.905 -18.745 38.045 -18.575 ;
      RECT 37.955 -17.558 38.045 -16.55 ;
      RECT 37.905 -16.955 38.045 -16.785 ;
      RECT 37.955 -15.75 38.045 -14.742 ;
      RECT 37.905 -15.515 38.045 -15.345 ;
      RECT 37.955 -14.328 38.045 -13.32 ;
      RECT 37.905 -13.725 38.045 -13.555 ;
      RECT 37.955 -12.52 38.045 -11.512 ;
      RECT 37.905 -12.285 38.045 -12.115 ;
      RECT 37.955 -11.098 38.045 -10.09 ;
      RECT 37.905 -10.495 38.045 -10.325 ;
      RECT 37.955 -9.29 38.045 -8.282 ;
      RECT 37.905 -9.055 38.045 -8.885 ;
      RECT 37.955 -7.868 38.045 -6.86 ;
      RECT 37.905 -7.265 38.045 -7.095 ;
      RECT 37.955 -6.06 38.045 -5.052 ;
      RECT 37.905 -5.825 38.045 -5.655 ;
      RECT 37.955 -4.638 38.045 -3.63 ;
      RECT 37.905 -4.035 38.045 -3.865 ;
      RECT 37.955 -2.83 38.045 -1.822 ;
      RECT 37.905 -2.595 38.045 -2.425 ;
      RECT 37.955 -1.408 38.045 -0.4 ;
      RECT 37.905 -0.805 38.045 -0.635 ;
      RECT 37.955 0.4 38.045 1.408 ;
      RECT 37.905 0.635 38.045 0.805 ;
      RECT 36.525 -111.685 38.005 -111.585 ;
      RECT 36.525 -112.195 36.625 -111.585 ;
      RECT 36.745 -109.15 38.005 -109.05 ;
      RECT 37.905 -109.475 38.005 -109.05 ;
      RECT 37.345 -109.475 37.445 -109.05 ;
      RECT 36.785 -109.475 36.885 -109.05 ;
      RECT 37.555 -101.538 37.645 -100.531 ;
      RECT 37.555 -101.225 37.695 -101.055 ;
      RECT 37.555 -99.729 37.645 -98.722 ;
      RECT 37.555 -99.205 37.695 -99.035 ;
      RECT 37.555 -98.308 37.645 -97.301 ;
      RECT 37.555 -97.995 37.695 -97.825 ;
      RECT 37.555 -96.499 37.645 -95.492 ;
      RECT 37.555 -95.975 37.695 -95.805 ;
      RECT 37.555 -95.078 37.645 -94.071 ;
      RECT 37.555 -94.765 37.695 -94.595 ;
      RECT 37.555 -93.269 37.645 -92.262 ;
      RECT 37.555 -92.745 37.695 -92.575 ;
      RECT 37.555 -91.848 37.645 -90.841 ;
      RECT 37.555 -91.535 37.695 -91.365 ;
      RECT 37.555 -90.039 37.645 -89.032 ;
      RECT 37.555 -89.515 37.695 -89.345 ;
      RECT 37.555 -88.618 37.645 -87.611 ;
      RECT 37.555 -88.305 37.695 -88.135 ;
      RECT 37.555 -86.809 37.645 -85.802 ;
      RECT 37.555 -86.285 37.695 -86.115 ;
      RECT 37.555 -85.388 37.645 -84.381 ;
      RECT 37.555 -85.075 37.695 -84.905 ;
      RECT 37.555 -83.579 37.645 -82.572 ;
      RECT 37.555 -83.055 37.695 -82.885 ;
      RECT 37.555 -82.158 37.645 -81.151 ;
      RECT 37.555 -81.845 37.695 -81.675 ;
      RECT 37.555 -80.349 37.645 -79.342 ;
      RECT 37.555 -79.825 37.695 -79.655 ;
      RECT 37.555 -78.928 37.645 -77.921 ;
      RECT 37.555 -78.615 37.695 -78.445 ;
      RECT 37.555 -77.119 37.645 -76.112 ;
      RECT 37.555 -76.595 37.695 -76.425 ;
      RECT 37.555 -75.698 37.645 -74.691 ;
      RECT 37.555 -75.385 37.695 -75.215 ;
      RECT 37.555 -73.889 37.645 -72.882 ;
      RECT 37.555 -73.365 37.695 -73.195 ;
      RECT 37.555 -72.468 37.645 -71.461 ;
      RECT 37.555 -72.155 37.695 -71.985 ;
      RECT 37.555 -70.659 37.645 -69.652 ;
      RECT 37.555 -70.135 37.695 -69.965 ;
      RECT 37.555 -69.238 37.645 -68.231 ;
      RECT 37.555 -68.925 37.695 -68.755 ;
      RECT 37.555 -67.429 37.645 -66.422 ;
      RECT 37.555 -66.905 37.695 -66.735 ;
      RECT 37.555 -66.008 37.645 -65.001 ;
      RECT 37.555 -65.695 37.695 -65.525 ;
      RECT 37.555 -64.199 37.645 -63.192 ;
      RECT 37.555 -63.675 37.695 -63.505 ;
      RECT 37.555 -62.778 37.645 -61.771 ;
      RECT 37.555 -62.465 37.695 -62.295 ;
      RECT 37.555 -60.969 37.645 -59.962 ;
      RECT 37.555 -60.445 37.695 -60.275 ;
      RECT 37.555 -59.548 37.645 -58.541 ;
      RECT 37.555 -59.235 37.695 -59.065 ;
      RECT 37.555 -57.739 37.645 -56.732 ;
      RECT 37.555 -57.215 37.695 -57.045 ;
      RECT 37.555 -56.318 37.645 -55.311 ;
      RECT 37.555 -56.005 37.695 -55.835 ;
      RECT 37.555 -54.509 37.645 -53.502 ;
      RECT 37.555 -53.985 37.695 -53.815 ;
      RECT 37.555 -53.088 37.645 -52.081 ;
      RECT 37.555 -52.775 37.695 -52.605 ;
      RECT 37.555 -51.279 37.645 -50.272 ;
      RECT 37.555 -50.755 37.695 -50.585 ;
      RECT 37.555 -49.858 37.645 -48.851 ;
      RECT 37.555 -49.545 37.695 -49.375 ;
      RECT 37.555 -48.049 37.645 -47.042 ;
      RECT 37.555 -47.525 37.695 -47.355 ;
      RECT 37.555 -46.628 37.645 -45.621 ;
      RECT 37.555 -46.315 37.695 -46.145 ;
      RECT 37.555 -44.819 37.645 -43.812 ;
      RECT 37.555 -44.295 37.695 -44.125 ;
      RECT 37.555 -43.398 37.645 -42.391 ;
      RECT 37.555 -43.085 37.695 -42.915 ;
      RECT 37.555 -41.589 37.645 -40.582 ;
      RECT 37.555 -41.065 37.695 -40.895 ;
      RECT 37.555 -40.168 37.645 -39.161 ;
      RECT 37.555 -39.855 37.695 -39.685 ;
      RECT 37.555 -38.359 37.645 -37.352 ;
      RECT 37.555 -37.835 37.695 -37.665 ;
      RECT 37.555 -36.938 37.645 -35.931 ;
      RECT 37.555 -36.625 37.695 -36.455 ;
      RECT 37.555 -35.129 37.645 -34.122 ;
      RECT 37.555 -34.605 37.695 -34.435 ;
      RECT 37.555 -33.708 37.645 -32.701 ;
      RECT 37.555 -33.395 37.695 -33.225 ;
      RECT 37.555 -31.899 37.645 -30.892 ;
      RECT 37.555 -31.375 37.695 -31.205 ;
      RECT 37.555 -30.478 37.645 -29.471 ;
      RECT 37.555 -30.165 37.695 -29.995 ;
      RECT 37.555 -28.669 37.645 -27.662 ;
      RECT 37.555 -28.145 37.695 -27.975 ;
      RECT 37.555 -27.248 37.645 -26.241 ;
      RECT 37.555 -26.935 37.695 -26.765 ;
      RECT 37.555 -25.439 37.645 -24.432 ;
      RECT 37.555 -24.915 37.695 -24.745 ;
      RECT 37.555 -24.018 37.645 -23.011 ;
      RECT 37.555 -23.705 37.695 -23.535 ;
      RECT 37.555 -22.209 37.645 -21.202 ;
      RECT 37.555 -21.685 37.695 -21.515 ;
      RECT 37.555 -20.788 37.645 -19.781 ;
      RECT 37.555 -20.475 37.695 -20.305 ;
      RECT 37.555 -18.979 37.645 -17.972 ;
      RECT 37.555 -18.455 37.695 -18.285 ;
      RECT 37.555 -17.558 37.645 -16.551 ;
      RECT 37.555 -17.245 37.695 -17.075 ;
      RECT 37.555 -15.749 37.645 -14.742 ;
      RECT 37.555 -15.225 37.695 -15.055 ;
      RECT 37.555 -14.328 37.645 -13.321 ;
      RECT 37.555 -14.015 37.695 -13.845 ;
      RECT 37.555 -12.519 37.645 -11.512 ;
      RECT 37.555 -11.995 37.695 -11.825 ;
      RECT 37.555 -11.098 37.645 -10.091 ;
      RECT 37.555 -10.785 37.695 -10.615 ;
      RECT 37.555 -9.289 37.645 -8.282 ;
      RECT 37.555 -8.765 37.695 -8.595 ;
      RECT 37.555 -7.868 37.645 -6.861 ;
      RECT 37.555 -7.555 37.695 -7.385 ;
      RECT 37.555 -6.059 37.645 -5.052 ;
      RECT 37.555 -5.535 37.695 -5.365 ;
      RECT 37.555 -4.638 37.645 -3.631 ;
      RECT 37.555 -4.325 37.695 -4.155 ;
      RECT 37.555 -2.829 37.645 -1.822 ;
      RECT 37.555 -2.305 37.695 -2.135 ;
      RECT 37.555 -1.408 37.645 -0.401 ;
      RECT 37.555 -1.095 37.695 -0.925 ;
      RECT 37.555 0.401 37.645 1.408 ;
      RECT 37.555 0.925 37.695 1.095 ;
      RECT 36.885 -111.495 37.055 -111.385 ;
      RECT 33.735 -111.495 37.055 -111.395 ;
      RECT 36.755 -101.538 36.845 -100.53 ;
      RECT 36.705 -100.935 36.845 -100.765 ;
      RECT 36.755 -99.73 36.845 -98.722 ;
      RECT 36.705 -99.495 36.845 -99.325 ;
      RECT 36.755 -98.308 36.845 -97.3 ;
      RECT 36.705 -97.705 36.845 -97.535 ;
      RECT 36.755 -96.5 36.845 -95.492 ;
      RECT 36.705 -96.265 36.845 -96.095 ;
      RECT 36.755 -95.078 36.845 -94.07 ;
      RECT 36.705 -94.475 36.845 -94.305 ;
      RECT 36.755 -93.27 36.845 -92.262 ;
      RECT 36.705 -93.035 36.845 -92.865 ;
      RECT 36.755 -91.848 36.845 -90.84 ;
      RECT 36.705 -91.245 36.845 -91.075 ;
      RECT 36.755 -90.04 36.845 -89.032 ;
      RECT 36.705 -89.805 36.845 -89.635 ;
      RECT 36.755 -88.618 36.845 -87.61 ;
      RECT 36.705 -88.015 36.845 -87.845 ;
      RECT 36.755 -86.81 36.845 -85.802 ;
      RECT 36.705 -86.575 36.845 -86.405 ;
      RECT 36.755 -85.388 36.845 -84.38 ;
      RECT 36.705 -84.785 36.845 -84.615 ;
      RECT 36.755 -83.58 36.845 -82.572 ;
      RECT 36.705 -83.345 36.845 -83.175 ;
      RECT 36.755 -82.158 36.845 -81.15 ;
      RECT 36.705 -81.555 36.845 -81.385 ;
      RECT 36.755 -80.35 36.845 -79.342 ;
      RECT 36.705 -80.115 36.845 -79.945 ;
      RECT 36.755 -78.928 36.845 -77.92 ;
      RECT 36.705 -78.325 36.845 -78.155 ;
      RECT 36.755 -77.12 36.845 -76.112 ;
      RECT 36.705 -76.885 36.845 -76.715 ;
      RECT 36.755 -75.698 36.845 -74.69 ;
      RECT 36.705 -75.095 36.845 -74.925 ;
      RECT 36.755 -73.89 36.845 -72.882 ;
      RECT 36.705 -73.655 36.845 -73.485 ;
      RECT 36.755 -72.468 36.845 -71.46 ;
      RECT 36.705 -71.865 36.845 -71.695 ;
      RECT 36.755 -70.66 36.845 -69.652 ;
      RECT 36.705 -70.425 36.845 -70.255 ;
      RECT 36.755 -69.238 36.845 -68.23 ;
      RECT 36.705 -68.635 36.845 -68.465 ;
      RECT 36.755 -67.43 36.845 -66.422 ;
      RECT 36.705 -67.195 36.845 -67.025 ;
      RECT 36.755 -66.008 36.845 -65 ;
      RECT 36.705 -65.405 36.845 -65.235 ;
      RECT 36.755 -64.2 36.845 -63.192 ;
      RECT 36.705 -63.965 36.845 -63.795 ;
      RECT 36.755 -62.778 36.845 -61.77 ;
      RECT 36.705 -62.175 36.845 -62.005 ;
      RECT 36.755 -60.97 36.845 -59.962 ;
      RECT 36.705 -60.735 36.845 -60.565 ;
      RECT 36.755 -59.548 36.845 -58.54 ;
      RECT 36.705 -58.945 36.845 -58.775 ;
      RECT 36.755 -57.74 36.845 -56.732 ;
      RECT 36.705 -57.505 36.845 -57.335 ;
      RECT 36.755 -56.318 36.845 -55.31 ;
      RECT 36.705 -55.715 36.845 -55.545 ;
      RECT 36.755 -54.51 36.845 -53.502 ;
      RECT 36.705 -54.275 36.845 -54.105 ;
      RECT 36.755 -53.088 36.845 -52.08 ;
      RECT 36.705 -52.485 36.845 -52.315 ;
      RECT 36.755 -51.28 36.845 -50.272 ;
      RECT 36.705 -51.045 36.845 -50.875 ;
      RECT 36.755 -49.858 36.845 -48.85 ;
      RECT 36.705 -49.255 36.845 -49.085 ;
      RECT 36.755 -48.05 36.845 -47.042 ;
      RECT 36.705 -47.815 36.845 -47.645 ;
      RECT 36.755 -46.628 36.845 -45.62 ;
      RECT 36.705 -46.025 36.845 -45.855 ;
      RECT 36.755 -44.82 36.845 -43.812 ;
      RECT 36.705 -44.585 36.845 -44.415 ;
      RECT 36.755 -43.398 36.845 -42.39 ;
      RECT 36.705 -42.795 36.845 -42.625 ;
      RECT 36.755 -41.59 36.845 -40.582 ;
      RECT 36.705 -41.355 36.845 -41.185 ;
      RECT 36.755 -40.168 36.845 -39.16 ;
      RECT 36.705 -39.565 36.845 -39.395 ;
      RECT 36.755 -38.36 36.845 -37.352 ;
      RECT 36.705 -38.125 36.845 -37.955 ;
      RECT 36.755 -36.938 36.845 -35.93 ;
      RECT 36.705 -36.335 36.845 -36.165 ;
      RECT 36.755 -35.13 36.845 -34.122 ;
      RECT 36.705 -34.895 36.845 -34.725 ;
      RECT 36.755 -33.708 36.845 -32.7 ;
      RECT 36.705 -33.105 36.845 -32.935 ;
      RECT 36.755 -31.9 36.845 -30.892 ;
      RECT 36.705 -31.665 36.845 -31.495 ;
      RECT 36.755 -30.478 36.845 -29.47 ;
      RECT 36.705 -29.875 36.845 -29.705 ;
      RECT 36.755 -28.67 36.845 -27.662 ;
      RECT 36.705 -28.435 36.845 -28.265 ;
      RECT 36.755 -27.248 36.845 -26.24 ;
      RECT 36.705 -26.645 36.845 -26.475 ;
      RECT 36.755 -25.44 36.845 -24.432 ;
      RECT 36.705 -25.205 36.845 -25.035 ;
      RECT 36.755 -24.018 36.845 -23.01 ;
      RECT 36.705 -23.415 36.845 -23.245 ;
      RECT 36.755 -22.21 36.845 -21.202 ;
      RECT 36.705 -21.975 36.845 -21.805 ;
      RECT 36.755 -20.788 36.845 -19.78 ;
      RECT 36.705 -20.185 36.845 -20.015 ;
      RECT 36.755 -18.98 36.845 -17.972 ;
      RECT 36.705 -18.745 36.845 -18.575 ;
      RECT 36.755 -17.558 36.845 -16.55 ;
      RECT 36.705 -16.955 36.845 -16.785 ;
      RECT 36.755 -15.75 36.845 -14.742 ;
      RECT 36.705 -15.515 36.845 -15.345 ;
      RECT 36.755 -14.328 36.845 -13.32 ;
      RECT 36.705 -13.725 36.845 -13.555 ;
      RECT 36.755 -12.52 36.845 -11.512 ;
      RECT 36.705 -12.285 36.845 -12.115 ;
      RECT 36.755 -11.098 36.845 -10.09 ;
      RECT 36.705 -10.495 36.845 -10.325 ;
      RECT 36.755 -9.29 36.845 -8.282 ;
      RECT 36.705 -9.055 36.845 -8.885 ;
      RECT 36.755 -7.868 36.845 -6.86 ;
      RECT 36.705 -7.265 36.845 -7.095 ;
      RECT 36.755 -6.06 36.845 -5.052 ;
      RECT 36.705 -5.825 36.845 -5.655 ;
      RECT 36.755 -4.638 36.845 -3.63 ;
      RECT 36.705 -4.035 36.845 -3.865 ;
      RECT 36.755 -2.83 36.845 -1.822 ;
      RECT 36.705 -2.595 36.845 -2.425 ;
      RECT 36.755 -1.408 36.845 -0.4 ;
      RECT 36.705 -0.805 36.845 -0.635 ;
      RECT 36.755 0.4 36.845 1.408 ;
      RECT 36.705 0.635 36.845 0.805 ;
      RECT 36.355 -101.538 36.445 -100.531 ;
      RECT 36.355 -101.225 36.495 -101.055 ;
      RECT 36.355 -99.729 36.445 -98.722 ;
      RECT 36.355 -99.205 36.495 -99.035 ;
      RECT 36.355 -98.308 36.445 -97.301 ;
      RECT 36.355 -97.995 36.495 -97.825 ;
      RECT 36.355 -96.499 36.445 -95.492 ;
      RECT 36.355 -95.975 36.495 -95.805 ;
      RECT 36.355 -95.078 36.445 -94.071 ;
      RECT 36.355 -94.765 36.495 -94.595 ;
      RECT 36.355 -93.269 36.445 -92.262 ;
      RECT 36.355 -92.745 36.495 -92.575 ;
      RECT 36.355 -91.848 36.445 -90.841 ;
      RECT 36.355 -91.535 36.495 -91.365 ;
      RECT 36.355 -90.039 36.445 -89.032 ;
      RECT 36.355 -89.515 36.495 -89.345 ;
      RECT 36.355 -88.618 36.445 -87.611 ;
      RECT 36.355 -88.305 36.495 -88.135 ;
      RECT 36.355 -86.809 36.445 -85.802 ;
      RECT 36.355 -86.285 36.495 -86.115 ;
      RECT 36.355 -85.388 36.445 -84.381 ;
      RECT 36.355 -85.075 36.495 -84.905 ;
      RECT 36.355 -83.579 36.445 -82.572 ;
      RECT 36.355 -83.055 36.495 -82.885 ;
      RECT 36.355 -82.158 36.445 -81.151 ;
      RECT 36.355 -81.845 36.495 -81.675 ;
      RECT 36.355 -80.349 36.445 -79.342 ;
      RECT 36.355 -79.825 36.495 -79.655 ;
      RECT 36.355 -78.928 36.445 -77.921 ;
      RECT 36.355 -78.615 36.495 -78.445 ;
      RECT 36.355 -77.119 36.445 -76.112 ;
      RECT 36.355 -76.595 36.495 -76.425 ;
      RECT 36.355 -75.698 36.445 -74.691 ;
      RECT 36.355 -75.385 36.495 -75.215 ;
      RECT 36.355 -73.889 36.445 -72.882 ;
      RECT 36.355 -73.365 36.495 -73.195 ;
      RECT 36.355 -72.468 36.445 -71.461 ;
      RECT 36.355 -72.155 36.495 -71.985 ;
      RECT 36.355 -70.659 36.445 -69.652 ;
      RECT 36.355 -70.135 36.495 -69.965 ;
      RECT 36.355 -69.238 36.445 -68.231 ;
      RECT 36.355 -68.925 36.495 -68.755 ;
      RECT 36.355 -67.429 36.445 -66.422 ;
      RECT 36.355 -66.905 36.495 -66.735 ;
      RECT 36.355 -66.008 36.445 -65.001 ;
      RECT 36.355 -65.695 36.495 -65.525 ;
      RECT 36.355 -64.199 36.445 -63.192 ;
      RECT 36.355 -63.675 36.495 -63.505 ;
      RECT 36.355 -62.778 36.445 -61.771 ;
      RECT 36.355 -62.465 36.495 -62.295 ;
      RECT 36.355 -60.969 36.445 -59.962 ;
      RECT 36.355 -60.445 36.495 -60.275 ;
      RECT 36.355 -59.548 36.445 -58.541 ;
      RECT 36.355 -59.235 36.495 -59.065 ;
      RECT 36.355 -57.739 36.445 -56.732 ;
      RECT 36.355 -57.215 36.495 -57.045 ;
      RECT 36.355 -56.318 36.445 -55.311 ;
      RECT 36.355 -56.005 36.495 -55.835 ;
      RECT 36.355 -54.509 36.445 -53.502 ;
      RECT 36.355 -53.985 36.495 -53.815 ;
      RECT 36.355 -53.088 36.445 -52.081 ;
      RECT 36.355 -52.775 36.495 -52.605 ;
      RECT 36.355 -51.279 36.445 -50.272 ;
      RECT 36.355 -50.755 36.495 -50.585 ;
      RECT 36.355 -49.858 36.445 -48.851 ;
      RECT 36.355 -49.545 36.495 -49.375 ;
      RECT 36.355 -48.049 36.445 -47.042 ;
      RECT 36.355 -47.525 36.495 -47.355 ;
      RECT 36.355 -46.628 36.445 -45.621 ;
      RECT 36.355 -46.315 36.495 -46.145 ;
      RECT 36.355 -44.819 36.445 -43.812 ;
      RECT 36.355 -44.295 36.495 -44.125 ;
      RECT 36.355 -43.398 36.445 -42.391 ;
      RECT 36.355 -43.085 36.495 -42.915 ;
      RECT 36.355 -41.589 36.445 -40.582 ;
      RECT 36.355 -41.065 36.495 -40.895 ;
      RECT 36.355 -40.168 36.445 -39.161 ;
      RECT 36.355 -39.855 36.495 -39.685 ;
      RECT 36.355 -38.359 36.445 -37.352 ;
      RECT 36.355 -37.835 36.495 -37.665 ;
      RECT 36.355 -36.938 36.445 -35.931 ;
      RECT 36.355 -36.625 36.495 -36.455 ;
      RECT 36.355 -35.129 36.445 -34.122 ;
      RECT 36.355 -34.605 36.495 -34.435 ;
      RECT 36.355 -33.708 36.445 -32.701 ;
      RECT 36.355 -33.395 36.495 -33.225 ;
      RECT 36.355 -31.899 36.445 -30.892 ;
      RECT 36.355 -31.375 36.495 -31.205 ;
      RECT 36.355 -30.478 36.445 -29.471 ;
      RECT 36.355 -30.165 36.495 -29.995 ;
      RECT 36.355 -28.669 36.445 -27.662 ;
      RECT 36.355 -28.145 36.495 -27.975 ;
      RECT 36.355 -27.248 36.445 -26.241 ;
      RECT 36.355 -26.935 36.495 -26.765 ;
      RECT 36.355 -25.439 36.445 -24.432 ;
      RECT 36.355 -24.915 36.495 -24.745 ;
      RECT 36.355 -24.018 36.445 -23.011 ;
      RECT 36.355 -23.705 36.495 -23.535 ;
      RECT 36.355 -22.209 36.445 -21.202 ;
      RECT 36.355 -21.685 36.495 -21.515 ;
      RECT 36.355 -20.788 36.445 -19.781 ;
      RECT 36.355 -20.475 36.495 -20.305 ;
      RECT 36.355 -18.979 36.445 -17.972 ;
      RECT 36.355 -18.455 36.495 -18.285 ;
      RECT 36.355 -17.558 36.445 -16.551 ;
      RECT 36.355 -17.245 36.495 -17.075 ;
      RECT 36.355 -15.749 36.445 -14.742 ;
      RECT 36.355 -15.225 36.495 -15.055 ;
      RECT 36.355 -14.328 36.445 -13.321 ;
      RECT 36.355 -14.015 36.495 -13.845 ;
      RECT 36.355 -12.519 36.445 -11.512 ;
      RECT 36.355 -11.995 36.495 -11.825 ;
      RECT 36.355 -11.098 36.445 -10.091 ;
      RECT 36.355 -10.785 36.495 -10.615 ;
      RECT 36.355 -9.289 36.445 -8.282 ;
      RECT 36.355 -8.765 36.495 -8.595 ;
      RECT 36.355 -7.868 36.445 -6.861 ;
      RECT 36.355 -7.555 36.495 -7.385 ;
      RECT 36.355 -6.059 36.445 -5.052 ;
      RECT 36.355 -5.535 36.495 -5.365 ;
      RECT 36.355 -4.638 36.445 -3.631 ;
      RECT 36.355 -4.325 36.495 -4.155 ;
      RECT 36.355 -2.829 36.445 -1.822 ;
      RECT 36.355 -2.305 36.495 -2.135 ;
      RECT 36.355 -1.408 36.445 -0.401 ;
      RECT 36.355 -1.095 36.495 -0.925 ;
      RECT 36.355 0.401 36.445 1.408 ;
      RECT 36.355 0.925 36.495 1.095 ;
      RECT 34.505 -111.685 35.985 -111.585 ;
      RECT 34.505 -112.055 34.605 -111.585 ;
      RECT 34.31 -114.395 35.885 -114.275 ;
      RECT 35.785 -114.895 35.885 -114.275 ;
      RECT 35.19 -114.895 35.29 -114.275 ;
      RECT 34.31 -114.85 34.41 -114.275 ;
      RECT 35.555 -101.538 35.645 -100.53 ;
      RECT 35.505 -100.935 35.645 -100.765 ;
      RECT 35.555 -99.73 35.645 -98.722 ;
      RECT 35.505 -99.495 35.645 -99.325 ;
      RECT 35.555 -98.308 35.645 -97.3 ;
      RECT 35.505 -97.705 35.645 -97.535 ;
      RECT 35.555 -96.5 35.645 -95.492 ;
      RECT 35.505 -96.265 35.645 -96.095 ;
      RECT 35.555 -95.078 35.645 -94.07 ;
      RECT 35.505 -94.475 35.645 -94.305 ;
      RECT 35.555 -93.27 35.645 -92.262 ;
      RECT 35.505 -93.035 35.645 -92.865 ;
      RECT 35.555 -91.848 35.645 -90.84 ;
      RECT 35.505 -91.245 35.645 -91.075 ;
      RECT 35.555 -90.04 35.645 -89.032 ;
      RECT 35.505 -89.805 35.645 -89.635 ;
      RECT 35.555 -88.618 35.645 -87.61 ;
      RECT 35.505 -88.015 35.645 -87.845 ;
      RECT 35.555 -86.81 35.645 -85.802 ;
      RECT 35.505 -86.575 35.645 -86.405 ;
      RECT 35.555 -85.388 35.645 -84.38 ;
      RECT 35.505 -84.785 35.645 -84.615 ;
      RECT 35.555 -83.58 35.645 -82.572 ;
      RECT 35.505 -83.345 35.645 -83.175 ;
      RECT 35.555 -82.158 35.645 -81.15 ;
      RECT 35.505 -81.555 35.645 -81.385 ;
      RECT 35.555 -80.35 35.645 -79.342 ;
      RECT 35.505 -80.115 35.645 -79.945 ;
      RECT 35.555 -78.928 35.645 -77.92 ;
      RECT 35.505 -78.325 35.645 -78.155 ;
      RECT 35.555 -77.12 35.645 -76.112 ;
      RECT 35.505 -76.885 35.645 -76.715 ;
      RECT 35.555 -75.698 35.645 -74.69 ;
      RECT 35.505 -75.095 35.645 -74.925 ;
      RECT 35.555 -73.89 35.645 -72.882 ;
      RECT 35.505 -73.655 35.645 -73.485 ;
      RECT 35.555 -72.468 35.645 -71.46 ;
      RECT 35.505 -71.865 35.645 -71.695 ;
      RECT 35.555 -70.66 35.645 -69.652 ;
      RECT 35.505 -70.425 35.645 -70.255 ;
      RECT 35.555 -69.238 35.645 -68.23 ;
      RECT 35.505 -68.635 35.645 -68.465 ;
      RECT 35.555 -67.43 35.645 -66.422 ;
      RECT 35.505 -67.195 35.645 -67.025 ;
      RECT 35.555 -66.008 35.645 -65 ;
      RECT 35.505 -65.405 35.645 -65.235 ;
      RECT 35.555 -64.2 35.645 -63.192 ;
      RECT 35.505 -63.965 35.645 -63.795 ;
      RECT 35.555 -62.778 35.645 -61.77 ;
      RECT 35.505 -62.175 35.645 -62.005 ;
      RECT 35.555 -60.97 35.645 -59.962 ;
      RECT 35.505 -60.735 35.645 -60.565 ;
      RECT 35.555 -59.548 35.645 -58.54 ;
      RECT 35.505 -58.945 35.645 -58.775 ;
      RECT 35.555 -57.74 35.645 -56.732 ;
      RECT 35.505 -57.505 35.645 -57.335 ;
      RECT 35.555 -56.318 35.645 -55.31 ;
      RECT 35.505 -55.715 35.645 -55.545 ;
      RECT 35.555 -54.51 35.645 -53.502 ;
      RECT 35.505 -54.275 35.645 -54.105 ;
      RECT 35.555 -53.088 35.645 -52.08 ;
      RECT 35.505 -52.485 35.645 -52.315 ;
      RECT 35.555 -51.28 35.645 -50.272 ;
      RECT 35.505 -51.045 35.645 -50.875 ;
      RECT 35.555 -49.858 35.645 -48.85 ;
      RECT 35.505 -49.255 35.645 -49.085 ;
      RECT 35.555 -48.05 35.645 -47.042 ;
      RECT 35.505 -47.815 35.645 -47.645 ;
      RECT 35.555 -46.628 35.645 -45.62 ;
      RECT 35.505 -46.025 35.645 -45.855 ;
      RECT 35.555 -44.82 35.645 -43.812 ;
      RECT 35.505 -44.585 35.645 -44.415 ;
      RECT 35.555 -43.398 35.645 -42.39 ;
      RECT 35.505 -42.795 35.645 -42.625 ;
      RECT 35.555 -41.59 35.645 -40.582 ;
      RECT 35.505 -41.355 35.645 -41.185 ;
      RECT 35.555 -40.168 35.645 -39.16 ;
      RECT 35.505 -39.565 35.645 -39.395 ;
      RECT 35.555 -38.36 35.645 -37.352 ;
      RECT 35.505 -38.125 35.645 -37.955 ;
      RECT 35.555 -36.938 35.645 -35.93 ;
      RECT 35.505 -36.335 35.645 -36.165 ;
      RECT 35.555 -35.13 35.645 -34.122 ;
      RECT 35.505 -34.895 35.645 -34.725 ;
      RECT 35.555 -33.708 35.645 -32.7 ;
      RECT 35.505 -33.105 35.645 -32.935 ;
      RECT 35.555 -31.9 35.645 -30.892 ;
      RECT 35.505 -31.665 35.645 -31.495 ;
      RECT 35.555 -30.478 35.645 -29.47 ;
      RECT 35.505 -29.875 35.645 -29.705 ;
      RECT 35.555 -28.67 35.645 -27.662 ;
      RECT 35.505 -28.435 35.645 -28.265 ;
      RECT 35.555 -27.248 35.645 -26.24 ;
      RECT 35.505 -26.645 35.645 -26.475 ;
      RECT 35.555 -25.44 35.645 -24.432 ;
      RECT 35.505 -25.205 35.645 -25.035 ;
      RECT 35.555 -24.018 35.645 -23.01 ;
      RECT 35.505 -23.415 35.645 -23.245 ;
      RECT 35.555 -22.21 35.645 -21.202 ;
      RECT 35.505 -21.975 35.645 -21.805 ;
      RECT 35.555 -20.788 35.645 -19.78 ;
      RECT 35.505 -20.185 35.645 -20.015 ;
      RECT 35.555 -18.98 35.645 -17.972 ;
      RECT 35.505 -18.745 35.645 -18.575 ;
      RECT 35.555 -17.558 35.645 -16.55 ;
      RECT 35.505 -16.955 35.645 -16.785 ;
      RECT 35.555 -15.75 35.645 -14.742 ;
      RECT 35.505 -15.515 35.645 -15.345 ;
      RECT 35.555 -14.328 35.645 -13.32 ;
      RECT 35.505 -13.725 35.645 -13.555 ;
      RECT 35.555 -12.52 35.645 -11.512 ;
      RECT 35.505 -12.285 35.645 -12.115 ;
      RECT 35.555 -11.098 35.645 -10.09 ;
      RECT 35.505 -10.495 35.645 -10.325 ;
      RECT 35.555 -9.29 35.645 -8.282 ;
      RECT 35.505 -9.055 35.645 -8.885 ;
      RECT 35.555 -7.868 35.645 -6.86 ;
      RECT 35.505 -7.265 35.645 -7.095 ;
      RECT 35.555 -6.06 35.645 -5.052 ;
      RECT 35.505 -5.825 35.645 -5.655 ;
      RECT 35.555 -4.638 35.645 -3.63 ;
      RECT 35.505 -4.035 35.645 -3.865 ;
      RECT 35.555 -2.83 35.645 -1.822 ;
      RECT 35.505 -2.595 35.645 -2.425 ;
      RECT 35.555 -1.408 35.645 -0.4 ;
      RECT 35.505 -0.805 35.645 -0.635 ;
      RECT 35.555 0.4 35.645 1.408 ;
      RECT 35.505 0.635 35.645 0.805 ;
      RECT 35.43 -114.685 35.605 -114.515 ;
      RECT 35.505 -114.895 35.605 -114.515 ;
      RECT 34.545 -113.555 34.645 -113.09 ;
      RECT 34.91 -113.555 35.01 -113.1 ;
      RECT 34.545 -113.555 35.39 -113.385 ;
      RECT 35.155 -101.538 35.245 -100.531 ;
      RECT 35.155 -101.225 35.295 -101.055 ;
      RECT 35.155 -99.729 35.245 -98.722 ;
      RECT 35.155 -99.205 35.295 -99.035 ;
      RECT 35.155 -98.308 35.245 -97.301 ;
      RECT 35.155 -97.995 35.295 -97.825 ;
      RECT 35.155 -96.499 35.245 -95.492 ;
      RECT 35.155 -95.975 35.295 -95.805 ;
      RECT 35.155 -95.078 35.245 -94.071 ;
      RECT 35.155 -94.765 35.295 -94.595 ;
      RECT 35.155 -93.269 35.245 -92.262 ;
      RECT 35.155 -92.745 35.295 -92.575 ;
      RECT 35.155 -91.848 35.245 -90.841 ;
      RECT 35.155 -91.535 35.295 -91.365 ;
      RECT 35.155 -90.039 35.245 -89.032 ;
      RECT 35.155 -89.515 35.295 -89.345 ;
      RECT 35.155 -88.618 35.245 -87.611 ;
      RECT 35.155 -88.305 35.295 -88.135 ;
      RECT 35.155 -86.809 35.245 -85.802 ;
      RECT 35.155 -86.285 35.295 -86.115 ;
      RECT 35.155 -85.388 35.245 -84.381 ;
      RECT 35.155 -85.075 35.295 -84.905 ;
      RECT 35.155 -83.579 35.245 -82.572 ;
      RECT 35.155 -83.055 35.295 -82.885 ;
      RECT 35.155 -82.158 35.245 -81.151 ;
      RECT 35.155 -81.845 35.295 -81.675 ;
      RECT 35.155 -80.349 35.245 -79.342 ;
      RECT 35.155 -79.825 35.295 -79.655 ;
      RECT 35.155 -78.928 35.245 -77.921 ;
      RECT 35.155 -78.615 35.295 -78.445 ;
      RECT 35.155 -77.119 35.245 -76.112 ;
      RECT 35.155 -76.595 35.295 -76.425 ;
      RECT 35.155 -75.698 35.245 -74.691 ;
      RECT 35.155 -75.385 35.295 -75.215 ;
      RECT 35.155 -73.889 35.245 -72.882 ;
      RECT 35.155 -73.365 35.295 -73.195 ;
      RECT 35.155 -72.468 35.245 -71.461 ;
      RECT 35.155 -72.155 35.295 -71.985 ;
      RECT 35.155 -70.659 35.245 -69.652 ;
      RECT 35.155 -70.135 35.295 -69.965 ;
      RECT 35.155 -69.238 35.245 -68.231 ;
      RECT 35.155 -68.925 35.295 -68.755 ;
      RECT 35.155 -67.429 35.245 -66.422 ;
      RECT 35.155 -66.905 35.295 -66.735 ;
      RECT 35.155 -66.008 35.245 -65.001 ;
      RECT 35.155 -65.695 35.295 -65.525 ;
      RECT 35.155 -64.199 35.245 -63.192 ;
      RECT 35.155 -63.675 35.295 -63.505 ;
      RECT 35.155 -62.778 35.245 -61.771 ;
      RECT 35.155 -62.465 35.295 -62.295 ;
      RECT 35.155 -60.969 35.245 -59.962 ;
      RECT 35.155 -60.445 35.295 -60.275 ;
      RECT 35.155 -59.548 35.245 -58.541 ;
      RECT 35.155 -59.235 35.295 -59.065 ;
      RECT 35.155 -57.739 35.245 -56.732 ;
      RECT 35.155 -57.215 35.295 -57.045 ;
      RECT 35.155 -56.318 35.245 -55.311 ;
      RECT 35.155 -56.005 35.295 -55.835 ;
      RECT 35.155 -54.509 35.245 -53.502 ;
      RECT 35.155 -53.985 35.295 -53.815 ;
      RECT 35.155 -53.088 35.245 -52.081 ;
      RECT 35.155 -52.775 35.295 -52.605 ;
      RECT 35.155 -51.279 35.245 -50.272 ;
      RECT 35.155 -50.755 35.295 -50.585 ;
      RECT 35.155 -49.858 35.245 -48.851 ;
      RECT 35.155 -49.545 35.295 -49.375 ;
      RECT 35.155 -48.049 35.245 -47.042 ;
      RECT 35.155 -47.525 35.295 -47.355 ;
      RECT 35.155 -46.628 35.245 -45.621 ;
      RECT 35.155 -46.315 35.295 -46.145 ;
      RECT 35.155 -44.819 35.245 -43.812 ;
      RECT 35.155 -44.295 35.295 -44.125 ;
      RECT 35.155 -43.398 35.245 -42.391 ;
      RECT 35.155 -43.085 35.295 -42.915 ;
      RECT 35.155 -41.589 35.245 -40.582 ;
      RECT 35.155 -41.065 35.295 -40.895 ;
      RECT 35.155 -40.168 35.245 -39.161 ;
      RECT 35.155 -39.855 35.295 -39.685 ;
      RECT 35.155 -38.359 35.245 -37.352 ;
      RECT 35.155 -37.835 35.295 -37.665 ;
      RECT 35.155 -36.938 35.245 -35.931 ;
      RECT 35.155 -36.625 35.295 -36.455 ;
      RECT 35.155 -35.129 35.245 -34.122 ;
      RECT 35.155 -34.605 35.295 -34.435 ;
      RECT 35.155 -33.708 35.245 -32.701 ;
      RECT 35.155 -33.395 35.295 -33.225 ;
      RECT 35.155 -31.899 35.245 -30.892 ;
      RECT 35.155 -31.375 35.295 -31.205 ;
      RECT 35.155 -30.478 35.245 -29.471 ;
      RECT 35.155 -30.165 35.295 -29.995 ;
      RECT 35.155 -28.669 35.245 -27.662 ;
      RECT 35.155 -28.145 35.295 -27.975 ;
      RECT 35.155 -27.248 35.245 -26.241 ;
      RECT 35.155 -26.935 35.295 -26.765 ;
      RECT 35.155 -25.439 35.245 -24.432 ;
      RECT 35.155 -24.915 35.295 -24.745 ;
      RECT 35.155 -24.018 35.245 -23.011 ;
      RECT 35.155 -23.705 35.295 -23.535 ;
      RECT 35.155 -22.209 35.245 -21.202 ;
      RECT 35.155 -21.685 35.295 -21.515 ;
      RECT 35.155 -20.788 35.245 -19.781 ;
      RECT 35.155 -20.475 35.295 -20.305 ;
      RECT 35.155 -18.979 35.245 -17.972 ;
      RECT 35.155 -18.455 35.295 -18.285 ;
      RECT 35.155 -17.558 35.245 -16.551 ;
      RECT 35.155 -17.245 35.295 -17.075 ;
      RECT 35.155 -15.749 35.245 -14.742 ;
      RECT 35.155 -15.225 35.295 -15.055 ;
      RECT 35.155 -14.328 35.245 -13.321 ;
      RECT 35.155 -14.015 35.295 -13.845 ;
      RECT 35.155 -12.519 35.245 -11.512 ;
      RECT 35.155 -11.995 35.295 -11.825 ;
      RECT 35.155 -11.098 35.245 -10.091 ;
      RECT 35.155 -10.785 35.295 -10.615 ;
      RECT 35.155 -9.289 35.245 -8.282 ;
      RECT 35.155 -8.765 35.295 -8.595 ;
      RECT 35.155 -7.868 35.245 -6.861 ;
      RECT 35.155 -7.555 35.295 -7.385 ;
      RECT 35.155 -6.059 35.245 -5.052 ;
      RECT 35.155 -5.535 35.295 -5.365 ;
      RECT 35.155 -4.638 35.245 -3.631 ;
      RECT 35.155 -4.325 35.295 -4.155 ;
      RECT 35.155 -2.829 35.245 -1.822 ;
      RECT 35.155 -2.305 35.295 -2.135 ;
      RECT 35.155 -1.408 35.245 -0.401 ;
      RECT 35.155 -1.095 35.295 -0.925 ;
      RECT 35.155 0.401 35.245 1.408 ;
      RECT 35.155 0.925 35.295 1.095 ;
      RECT 34.84 -114.685 35.01 -114.515 ;
      RECT 34.91 -114.895 35.01 -114.515 ;
      RECT 34.355 -101.538 34.445 -100.53 ;
      RECT 34.305 -100.935 34.445 -100.765 ;
      RECT 34.355 -99.73 34.445 -98.722 ;
      RECT 34.305 -99.495 34.445 -99.325 ;
      RECT 34.355 -98.308 34.445 -97.3 ;
      RECT 34.305 -97.705 34.445 -97.535 ;
      RECT 34.355 -96.5 34.445 -95.492 ;
      RECT 34.305 -96.265 34.445 -96.095 ;
      RECT 34.355 -95.078 34.445 -94.07 ;
      RECT 34.305 -94.475 34.445 -94.305 ;
      RECT 34.355 -93.27 34.445 -92.262 ;
      RECT 34.305 -93.035 34.445 -92.865 ;
      RECT 34.355 -91.848 34.445 -90.84 ;
      RECT 34.305 -91.245 34.445 -91.075 ;
      RECT 34.355 -90.04 34.445 -89.032 ;
      RECT 34.305 -89.805 34.445 -89.635 ;
      RECT 34.355 -88.618 34.445 -87.61 ;
      RECT 34.305 -88.015 34.445 -87.845 ;
      RECT 34.355 -86.81 34.445 -85.802 ;
      RECT 34.305 -86.575 34.445 -86.405 ;
      RECT 34.355 -85.388 34.445 -84.38 ;
      RECT 34.305 -84.785 34.445 -84.615 ;
      RECT 34.355 -83.58 34.445 -82.572 ;
      RECT 34.305 -83.345 34.445 -83.175 ;
      RECT 34.355 -82.158 34.445 -81.15 ;
      RECT 34.305 -81.555 34.445 -81.385 ;
      RECT 34.355 -80.35 34.445 -79.342 ;
      RECT 34.305 -80.115 34.445 -79.945 ;
      RECT 34.355 -78.928 34.445 -77.92 ;
      RECT 34.305 -78.325 34.445 -78.155 ;
      RECT 34.355 -77.12 34.445 -76.112 ;
      RECT 34.305 -76.885 34.445 -76.715 ;
      RECT 34.355 -75.698 34.445 -74.69 ;
      RECT 34.305 -75.095 34.445 -74.925 ;
      RECT 34.355 -73.89 34.445 -72.882 ;
      RECT 34.305 -73.655 34.445 -73.485 ;
      RECT 34.355 -72.468 34.445 -71.46 ;
      RECT 34.305 -71.865 34.445 -71.695 ;
      RECT 34.355 -70.66 34.445 -69.652 ;
      RECT 34.305 -70.425 34.445 -70.255 ;
      RECT 34.355 -69.238 34.445 -68.23 ;
      RECT 34.305 -68.635 34.445 -68.465 ;
      RECT 34.355 -67.43 34.445 -66.422 ;
      RECT 34.305 -67.195 34.445 -67.025 ;
      RECT 34.355 -66.008 34.445 -65 ;
      RECT 34.305 -65.405 34.445 -65.235 ;
      RECT 34.355 -64.2 34.445 -63.192 ;
      RECT 34.305 -63.965 34.445 -63.795 ;
      RECT 34.355 -62.778 34.445 -61.77 ;
      RECT 34.305 -62.175 34.445 -62.005 ;
      RECT 34.355 -60.97 34.445 -59.962 ;
      RECT 34.305 -60.735 34.445 -60.565 ;
      RECT 34.355 -59.548 34.445 -58.54 ;
      RECT 34.305 -58.945 34.445 -58.775 ;
      RECT 34.355 -57.74 34.445 -56.732 ;
      RECT 34.305 -57.505 34.445 -57.335 ;
      RECT 34.355 -56.318 34.445 -55.31 ;
      RECT 34.305 -55.715 34.445 -55.545 ;
      RECT 34.355 -54.51 34.445 -53.502 ;
      RECT 34.305 -54.275 34.445 -54.105 ;
      RECT 34.355 -53.088 34.445 -52.08 ;
      RECT 34.305 -52.485 34.445 -52.315 ;
      RECT 34.355 -51.28 34.445 -50.272 ;
      RECT 34.305 -51.045 34.445 -50.875 ;
      RECT 34.355 -49.858 34.445 -48.85 ;
      RECT 34.305 -49.255 34.445 -49.085 ;
      RECT 34.355 -48.05 34.445 -47.042 ;
      RECT 34.305 -47.815 34.445 -47.645 ;
      RECT 34.355 -46.628 34.445 -45.62 ;
      RECT 34.305 -46.025 34.445 -45.855 ;
      RECT 34.355 -44.82 34.445 -43.812 ;
      RECT 34.305 -44.585 34.445 -44.415 ;
      RECT 34.355 -43.398 34.445 -42.39 ;
      RECT 34.305 -42.795 34.445 -42.625 ;
      RECT 34.355 -41.59 34.445 -40.582 ;
      RECT 34.305 -41.355 34.445 -41.185 ;
      RECT 34.355 -40.168 34.445 -39.16 ;
      RECT 34.305 -39.565 34.445 -39.395 ;
      RECT 34.355 -38.36 34.445 -37.352 ;
      RECT 34.305 -38.125 34.445 -37.955 ;
      RECT 34.355 -36.938 34.445 -35.93 ;
      RECT 34.305 -36.335 34.445 -36.165 ;
      RECT 34.355 -35.13 34.445 -34.122 ;
      RECT 34.305 -34.895 34.445 -34.725 ;
      RECT 34.355 -33.708 34.445 -32.7 ;
      RECT 34.305 -33.105 34.445 -32.935 ;
      RECT 34.355 -31.9 34.445 -30.892 ;
      RECT 34.305 -31.665 34.445 -31.495 ;
      RECT 34.355 -30.478 34.445 -29.47 ;
      RECT 34.305 -29.875 34.445 -29.705 ;
      RECT 34.355 -28.67 34.445 -27.662 ;
      RECT 34.305 -28.435 34.445 -28.265 ;
      RECT 34.355 -27.248 34.445 -26.24 ;
      RECT 34.305 -26.645 34.445 -26.475 ;
      RECT 34.355 -25.44 34.445 -24.432 ;
      RECT 34.305 -25.205 34.445 -25.035 ;
      RECT 34.355 -24.018 34.445 -23.01 ;
      RECT 34.305 -23.415 34.445 -23.245 ;
      RECT 34.355 -22.21 34.445 -21.202 ;
      RECT 34.305 -21.975 34.445 -21.805 ;
      RECT 34.355 -20.788 34.445 -19.78 ;
      RECT 34.305 -20.185 34.445 -20.015 ;
      RECT 34.355 -18.98 34.445 -17.972 ;
      RECT 34.305 -18.745 34.445 -18.575 ;
      RECT 34.355 -17.558 34.445 -16.55 ;
      RECT 34.305 -16.955 34.445 -16.785 ;
      RECT 34.355 -15.75 34.445 -14.742 ;
      RECT 34.305 -15.515 34.445 -15.345 ;
      RECT 34.355 -14.328 34.445 -13.32 ;
      RECT 34.305 -13.725 34.445 -13.555 ;
      RECT 34.355 -12.52 34.445 -11.512 ;
      RECT 34.305 -12.285 34.445 -12.115 ;
      RECT 34.355 -11.098 34.445 -10.09 ;
      RECT 34.305 -10.495 34.445 -10.325 ;
      RECT 34.355 -9.29 34.445 -8.282 ;
      RECT 34.305 -9.055 34.445 -8.885 ;
      RECT 34.355 -7.868 34.445 -6.86 ;
      RECT 34.305 -7.265 34.445 -7.095 ;
      RECT 34.355 -6.06 34.445 -5.052 ;
      RECT 34.305 -5.825 34.445 -5.655 ;
      RECT 34.355 -4.638 34.445 -3.63 ;
      RECT 34.305 -4.035 34.445 -3.865 ;
      RECT 34.355 -2.83 34.445 -1.822 ;
      RECT 34.305 -2.595 34.445 -2.425 ;
      RECT 34.355 -1.408 34.445 -0.4 ;
      RECT 34.305 -0.805 34.445 -0.635 ;
      RECT 34.355 0.4 34.445 1.408 ;
      RECT 34.305 0.635 34.445 0.805 ;
      RECT 33.955 -101.538 34.045 -100.531 ;
      RECT 33.955 -101.225 34.095 -101.055 ;
      RECT 33.955 -99.729 34.045 -98.722 ;
      RECT 33.955 -99.205 34.095 -99.035 ;
      RECT 33.955 -98.308 34.045 -97.301 ;
      RECT 33.955 -97.995 34.095 -97.825 ;
      RECT 33.955 -96.499 34.045 -95.492 ;
      RECT 33.955 -95.975 34.095 -95.805 ;
      RECT 33.955 -95.078 34.045 -94.071 ;
      RECT 33.955 -94.765 34.095 -94.595 ;
      RECT 33.955 -93.269 34.045 -92.262 ;
      RECT 33.955 -92.745 34.095 -92.575 ;
      RECT 33.955 -91.848 34.045 -90.841 ;
      RECT 33.955 -91.535 34.095 -91.365 ;
      RECT 33.955 -90.039 34.045 -89.032 ;
      RECT 33.955 -89.515 34.095 -89.345 ;
      RECT 33.955 -88.618 34.045 -87.611 ;
      RECT 33.955 -88.305 34.095 -88.135 ;
      RECT 33.955 -86.809 34.045 -85.802 ;
      RECT 33.955 -86.285 34.095 -86.115 ;
      RECT 33.955 -85.388 34.045 -84.381 ;
      RECT 33.955 -85.075 34.095 -84.905 ;
      RECT 33.955 -83.579 34.045 -82.572 ;
      RECT 33.955 -83.055 34.095 -82.885 ;
      RECT 33.955 -82.158 34.045 -81.151 ;
      RECT 33.955 -81.845 34.095 -81.675 ;
      RECT 33.955 -80.349 34.045 -79.342 ;
      RECT 33.955 -79.825 34.095 -79.655 ;
      RECT 33.955 -78.928 34.045 -77.921 ;
      RECT 33.955 -78.615 34.095 -78.445 ;
      RECT 33.955 -77.119 34.045 -76.112 ;
      RECT 33.955 -76.595 34.095 -76.425 ;
      RECT 33.955 -75.698 34.045 -74.691 ;
      RECT 33.955 -75.385 34.095 -75.215 ;
      RECT 33.955 -73.889 34.045 -72.882 ;
      RECT 33.955 -73.365 34.095 -73.195 ;
      RECT 33.955 -72.468 34.045 -71.461 ;
      RECT 33.955 -72.155 34.095 -71.985 ;
      RECT 33.955 -70.659 34.045 -69.652 ;
      RECT 33.955 -70.135 34.095 -69.965 ;
      RECT 33.955 -69.238 34.045 -68.231 ;
      RECT 33.955 -68.925 34.095 -68.755 ;
      RECT 33.955 -67.429 34.045 -66.422 ;
      RECT 33.955 -66.905 34.095 -66.735 ;
      RECT 33.955 -66.008 34.045 -65.001 ;
      RECT 33.955 -65.695 34.095 -65.525 ;
      RECT 33.955 -64.199 34.045 -63.192 ;
      RECT 33.955 -63.675 34.095 -63.505 ;
      RECT 33.955 -62.778 34.045 -61.771 ;
      RECT 33.955 -62.465 34.095 -62.295 ;
      RECT 33.955 -60.969 34.045 -59.962 ;
      RECT 33.955 -60.445 34.095 -60.275 ;
      RECT 33.955 -59.548 34.045 -58.541 ;
      RECT 33.955 -59.235 34.095 -59.065 ;
      RECT 33.955 -57.739 34.045 -56.732 ;
      RECT 33.955 -57.215 34.095 -57.045 ;
      RECT 33.955 -56.318 34.045 -55.311 ;
      RECT 33.955 -56.005 34.095 -55.835 ;
      RECT 33.955 -54.509 34.045 -53.502 ;
      RECT 33.955 -53.985 34.095 -53.815 ;
      RECT 33.955 -53.088 34.045 -52.081 ;
      RECT 33.955 -52.775 34.095 -52.605 ;
      RECT 33.955 -51.279 34.045 -50.272 ;
      RECT 33.955 -50.755 34.095 -50.585 ;
      RECT 33.955 -49.858 34.045 -48.851 ;
      RECT 33.955 -49.545 34.095 -49.375 ;
      RECT 33.955 -48.049 34.045 -47.042 ;
      RECT 33.955 -47.525 34.095 -47.355 ;
      RECT 33.955 -46.628 34.045 -45.621 ;
      RECT 33.955 -46.315 34.095 -46.145 ;
      RECT 33.955 -44.819 34.045 -43.812 ;
      RECT 33.955 -44.295 34.095 -44.125 ;
      RECT 33.955 -43.398 34.045 -42.391 ;
      RECT 33.955 -43.085 34.095 -42.915 ;
      RECT 33.955 -41.589 34.045 -40.582 ;
      RECT 33.955 -41.065 34.095 -40.895 ;
      RECT 33.955 -40.168 34.045 -39.161 ;
      RECT 33.955 -39.855 34.095 -39.685 ;
      RECT 33.955 -38.359 34.045 -37.352 ;
      RECT 33.955 -37.835 34.095 -37.665 ;
      RECT 33.955 -36.938 34.045 -35.931 ;
      RECT 33.955 -36.625 34.095 -36.455 ;
      RECT 33.955 -35.129 34.045 -34.122 ;
      RECT 33.955 -34.605 34.095 -34.435 ;
      RECT 33.955 -33.708 34.045 -32.701 ;
      RECT 33.955 -33.395 34.095 -33.225 ;
      RECT 33.955 -31.899 34.045 -30.892 ;
      RECT 33.955 -31.375 34.095 -31.205 ;
      RECT 33.955 -30.478 34.045 -29.471 ;
      RECT 33.955 -30.165 34.095 -29.995 ;
      RECT 33.955 -28.669 34.045 -27.662 ;
      RECT 33.955 -28.145 34.095 -27.975 ;
      RECT 33.955 -27.248 34.045 -26.241 ;
      RECT 33.955 -26.935 34.095 -26.765 ;
      RECT 33.955 -25.439 34.045 -24.432 ;
      RECT 33.955 -24.915 34.095 -24.745 ;
      RECT 33.955 -24.018 34.045 -23.011 ;
      RECT 33.955 -23.705 34.095 -23.535 ;
      RECT 33.955 -22.209 34.045 -21.202 ;
      RECT 33.955 -21.685 34.095 -21.515 ;
      RECT 33.955 -20.788 34.045 -19.781 ;
      RECT 33.955 -20.475 34.095 -20.305 ;
      RECT 33.955 -18.979 34.045 -17.972 ;
      RECT 33.955 -18.455 34.095 -18.285 ;
      RECT 33.955 -17.558 34.045 -16.551 ;
      RECT 33.955 -17.245 34.095 -17.075 ;
      RECT 33.955 -15.749 34.045 -14.742 ;
      RECT 33.955 -15.225 34.095 -15.055 ;
      RECT 33.955 -14.328 34.045 -13.321 ;
      RECT 33.955 -14.015 34.095 -13.845 ;
      RECT 33.955 -12.519 34.045 -11.512 ;
      RECT 33.955 -11.995 34.095 -11.825 ;
      RECT 33.955 -11.098 34.045 -10.091 ;
      RECT 33.955 -10.785 34.095 -10.615 ;
      RECT 33.955 -9.289 34.045 -8.282 ;
      RECT 33.955 -8.765 34.095 -8.595 ;
      RECT 33.955 -7.868 34.045 -6.861 ;
      RECT 33.955 -7.555 34.095 -7.385 ;
      RECT 33.955 -6.059 34.045 -5.052 ;
      RECT 33.955 -5.535 34.095 -5.365 ;
      RECT 33.955 -4.638 34.045 -3.631 ;
      RECT 33.955 -4.325 34.095 -4.155 ;
      RECT 33.955 -2.829 34.045 -1.822 ;
      RECT 33.955 -2.305 34.095 -2.135 ;
      RECT 33.955 -1.408 34.045 -0.401 ;
      RECT 33.955 -1.095 34.095 -0.925 ;
      RECT 33.955 0.401 34.045 1.408 ;
      RECT 33.955 0.925 34.095 1.095 ;
      RECT 29.785 -108.935 33.565 -108.815 ;
      RECT 31.105 -109.475 31.205 -108.815 ;
      RECT 30.545 -109.475 30.645 -108.815 ;
      RECT 29.985 -109.475 30.085 -108.815 ;
      RECT 33.155 -101.538 33.245 -100.53 ;
      RECT 33.105 -100.935 33.245 -100.765 ;
      RECT 33.155 -99.73 33.245 -98.722 ;
      RECT 33.105 -99.495 33.245 -99.325 ;
      RECT 33.155 -98.308 33.245 -97.3 ;
      RECT 33.105 -97.705 33.245 -97.535 ;
      RECT 33.155 -96.5 33.245 -95.492 ;
      RECT 33.105 -96.265 33.245 -96.095 ;
      RECT 33.155 -95.078 33.245 -94.07 ;
      RECT 33.105 -94.475 33.245 -94.305 ;
      RECT 33.155 -93.27 33.245 -92.262 ;
      RECT 33.105 -93.035 33.245 -92.865 ;
      RECT 33.155 -91.848 33.245 -90.84 ;
      RECT 33.105 -91.245 33.245 -91.075 ;
      RECT 33.155 -90.04 33.245 -89.032 ;
      RECT 33.105 -89.805 33.245 -89.635 ;
      RECT 33.155 -88.618 33.245 -87.61 ;
      RECT 33.105 -88.015 33.245 -87.845 ;
      RECT 33.155 -86.81 33.245 -85.802 ;
      RECT 33.105 -86.575 33.245 -86.405 ;
      RECT 33.155 -85.388 33.245 -84.38 ;
      RECT 33.105 -84.785 33.245 -84.615 ;
      RECT 33.155 -83.58 33.245 -82.572 ;
      RECT 33.105 -83.345 33.245 -83.175 ;
      RECT 33.155 -82.158 33.245 -81.15 ;
      RECT 33.105 -81.555 33.245 -81.385 ;
      RECT 33.155 -80.35 33.245 -79.342 ;
      RECT 33.105 -80.115 33.245 -79.945 ;
      RECT 33.155 -78.928 33.245 -77.92 ;
      RECT 33.105 -78.325 33.245 -78.155 ;
      RECT 33.155 -77.12 33.245 -76.112 ;
      RECT 33.105 -76.885 33.245 -76.715 ;
      RECT 33.155 -75.698 33.245 -74.69 ;
      RECT 33.105 -75.095 33.245 -74.925 ;
      RECT 33.155 -73.89 33.245 -72.882 ;
      RECT 33.105 -73.655 33.245 -73.485 ;
      RECT 33.155 -72.468 33.245 -71.46 ;
      RECT 33.105 -71.865 33.245 -71.695 ;
      RECT 33.155 -70.66 33.245 -69.652 ;
      RECT 33.105 -70.425 33.245 -70.255 ;
      RECT 33.155 -69.238 33.245 -68.23 ;
      RECT 33.105 -68.635 33.245 -68.465 ;
      RECT 33.155 -67.43 33.245 -66.422 ;
      RECT 33.105 -67.195 33.245 -67.025 ;
      RECT 33.155 -66.008 33.245 -65 ;
      RECT 33.105 -65.405 33.245 -65.235 ;
      RECT 33.155 -64.2 33.245 -63.192 ;
      RECT 33.105 -63.965 33.245 -63.795 ;
      RECT 33.155 -62.778 33.245 -61.77 ;
      RECT 33.105 -62.175 33.245 -62.005 ;
      RECT 33.155 -60.97 33.245 -59.962 ;
      RECT 33.105 -60.735 33.245 -60.565 ;
      RECT 33.155 -59.548 33.245 -58.54 ;
      RECT 33.105 -58.945 33.245 -58.775 ;
      RECT 33.155 -57.74 33.245 -56.732 ;
      RECT 33.105 -57.505 33.245 -57.335 ;
      RECT 33.155 -56.318 33.245 -55.31 ;
      RECT 33.105 -55.715 33.245 -55.545 ;
      RECT 33.155 -54.51 33.245 -53.502 ;
      RECT 33.105 -54.275 33.245 -54.105 ;
      RECT 33.155 -53.088 33.245 -52.08 ;
      RECT 33.105 -52.485 33.245 -52.315 ;
      RECT 33.155 -51.28 33.245 -50.272 ;
      RECT 33.105 -51.045 33.245 -50.875 ;
      RECT 33.155 -49.858 33.245 -48.85 ;
      RECT 33.105 -49.255 33.245 -49.085 ;
      RECT 33.155 -48.05 33.245 -47.042 ;
      RECT 33.105 -47.815 33.245 -47.645 ;
      RECT 33.155 -46.628 33.245 -45.62 ;
      RECT 33.105 -46.025 33.245 -45.855 ;
      RECT 33.155 -44.82 33.245 -43.812 ;
      RECT 33.105 -44.585 33.245 -44.415 ;
      RECT 33.155 -43.398 33.245 -42.39 ;
      RECT 33.105 -42.795 33.245 -42.625 ;
      RECT 33.155 -41.59 33.245 -40.582 ;
      RECT 33.105 -41.355 33.245 -41.185 ;
      RECT 33.155 -40.168 33.245 -39.16 ;
      RECT 33.105 -39.565 33.245 -39.395 ;
      RECT 33.155 -38.36 33.245 -37.352 ;
      RECT 33.105 -38.125 33.245 -37.955 ;
      RECT 33.155 -36.938 33.245 -35.93 ;
      RECT 33.105 -36.335 33.245 -36.165 ;
      RECT 33.155 -35.13 33.245 -34.122 ;
      RECT 33.105 -34.895 33.245 -34.725 ;
      RECT 33.155 -33.708 33.245 -32.7 ;
      RECT 33.105 -33.105 33.245 -32.935 ;
      RECT 33.155 -31.9 33.245 -30.892 ;
      RECT 33.105 -31.665 33.245 -31.495 ;
      RECT 33.155 -30.478 33.245 -29.47 ;
      RECT 33.105 -29.875 33.245 -29.705 ;
      RECT 33.155 -28.67 33.245 -27.662 ;
      RECT 33.105 -28.435 33.245 -28.265 ;
      RECT 33.155 -27.248 33.245 -26.24 ;
      RECT 33.105 -26.645 33.245 -26.475 ;
      RECT 33.155 -25.44 33.245 -24.432 ;
      RECT 33.105 -25.205 33.245 -25.035 ;
      RECT 33.155 -24.018 33.245 -23.01 ;
      RECT 33.105 -23.415 33.245 -23.245 ;
      RECT 33.155 -22.21 33.245 -21.202 ;
      RECT 33.105 -21.975 33.245 -21.805 ;
      RECT 33.155 -20.788 33.245 -19.78 ;
      RECT 33.105 -20.185 33.245 -20.015 ;
      RECT 33.155 -18.98 33.245 -17.972 ;
      RECT 33.105 -18.745 33.245 -18.575 ;
      RECT 33.155 -17.558 33.245 -16.55 ;
      RECT 33.105 -16.955 33.245 -16.785 ;
      RECT 33.155 -15.75 33.245 -14.742 ;
      RECT 33.105 -15.515 33.245 -15.345 ;
      RECT 33.155 -14.328 33.245 -13.32 ;
      RECT 33.105 -13.725 33.245 -13.555 ;
      RECT 33.155 -12.52 33.245 -11.512 ;
      RECT 33.105 -12.285 33.245 -12.115 ;
      RECT 33.155 -11.098 33.245 -10.09 ;
      RECT 33.105 -10.495 33.245 -10.325 ;
      RECT 33.155 -9.29 33.245 -8.282 ;
      RECT 33.105 -9.055 33.245 -8.885 ;
      RECT 33.155 -7.868 33.245 -6.86 ;
      RECT 33.105 -7.265 33.245 -7.095 ;
      RECT 33.155 -6.06 33.245 -5.052 ;
      RECT 33.105 -5.825 33.245 -5.655 ;
      RECT 33.155 -4.638 33.245 -3.63 ;
      RECT 33.105 -4.035 33.245 -3.865 ;
      RECT 33.155 -2.83 33.245 -1.822 ;
      RECT 33.105 -2.595 33.245 -2.425 ;
      RECT 33.155 -1.408 33.245 -0.4 ;
      RECT 33.105 -0.805 33.245 -0.635 ;
      RECT 33.155 0.4 33.245 1.408 ;
      RECT 33.105 0.635 33.245 0.805 ;
      RECT 31.725 -111.685 33.205 -111.585 ;
      RECT 31.725 -112.195 31.825 -111.585 ;
      RECT 31.945 -109.15 33.205 -109.05 ;
      RECT 33.105 -109.475 33.205 -109.05 ;
      RECT 32.545 -109.475 32.645 -109.05 ;
      RECT 31.985 -109.475 32.085 -109.05 ;
      RECT 32.755 -101.538 32.845 -100.531 ;
      RECT 32.755 -101.225 32.895 -101.055 ;
      RECT 32.755 -99.729 32.845 -98.722 ;
      RECT 32.755 -99.205 32.895 -99.035 ;
      RECT 32.755 -98.308 32.845 -97.301 ;
      RECT 32.755 -97.995 32.895 -97.825 ;
      RECT 32.755 -96.499 32.845 -95.492 ;
      RECT 32.755 -95.975 32.895 -95.805 ;
      RECT 32.755 -95.078 32.845 -94.071 ;
      RECT 32.755 -94.765 32.895 -94.595 ;
      RECT 32.755 -93.269 32.845 -92.262 ;
      RECT 32.755 -92.745 32.895 -92.575 ;
      RECT 32.755 -91.848 32.845 -90.841 ;
      RECT 32.755 -91.535 32.895 -91.365 ;
      RECT 32.755 -90.039 32.845 -89.032 ;
      RECT 32.755 -89.515 32.895 -89.345 ;
      RECT 32.755 -88.618 32.845 -87.611 ;
      RECT 32.755 -88.305 32.895 -88.135 ;
      RECT 32.755 -86.809 32.845 -85.802 ;
      RECT 32.755 -86.285 32.895 -86.115 ;
      RECT 32.755 -85.388 32.845 -84.381 ;
      RECT 32.755 -85.075 32.895 -84.905 ;
      RECT 32.755 -83.579 32.845 -82.572 ;
      RECT 32.755 -83.055 32.895 -82.885 ;
      RECT 32.755 -82.158 32.845 -81.151 ;
      RECT 32.755 -81.845 32.895 -81.675 ;
      RECT 32.755 -80.349 32.845 -79.342 ;
      RECT 32.755 -79.825 32.895 -79.655 ;
      RECT 32.755 -78.928 32.845 -77.921 ;
      RECT 32.755 -78.615 32.895 -78.445 ;
      RECT 32.755 -77.119 32.845 -76.112 ;
      RECT 32.755 -76.595 32.895 -76.425 ;
      RECT 32.755 -75.698 32.845 -74.691 ;
      RECT 32.755 -75.385 32.895 -75.215 ;
      RECT 32.755 -73.889 32.845 -72.882 ;
      RECT 32.755 -73.365 32.895 -73.195 ;
      RECT 32.755 -72.468 32.845 -71.461 ;
      RECT 32.755 -72.155 32.895 -71.985 ;
      RECT 32.755 -70.659 32.845 -69.652 ;
      RECT 32.755 -70.135 32.895 -69.965 ;
      RECT 32.755 -69.238 32.845 -68.231 ;
      RECT 32.755 -68.925 32.895 -68.755 ;
      RECT 32.755 -67.429 32.845 -66.422 ;
      RECT 32.755 -66.905 32.895 -66.735 ;
      RECT 32.755 -66.008 32.845 -65.001 ;
      RECT 32.755 -65.695 32.895 -65.525 ;
      RECT 32.755 -64.199 32.845 -63.192 ;
      RECT 32.755 -63.675 32.895 -63.505 ;
      RECT 32.755 -62.778 32.845 -61.771 ;
      RECT 32.755 -62.465 32.895 -62.295 ;
      RECT 32.755 -60.969 32.845 -59.962 ;
      RECT 32.755 -60.445 32.895 -60.275 ;
      RECT 32.755 -59.548 32.845 -58.541 ;
      RECT 32.755 -59.235 32.895 -59.065 ;
      RECT 32.755 -57.739 32.845 -56.732 ;
      RECT 32.755 -57.215 32.895 -57.045 ;
      RECT 32.755 -56.318 32.845 -55.311 ;
      RECT 32.755 -56.005 32.895 -55.835 ;
      RECT 32.755 -54.509 32.845 -53.502 ;
      RECT 32.755 -53.985 32.895 -53.815 ;
      RECT 32.755 -53.088 32.845 -52.081 ;
      RECT 32.755 -52.775 32.895 -52.605 ;
      RECT 32.755 -51.279 32.845 -50.272 ;
      RECT 32.755 -50.755 32.895 -50.585 ;
      RECT 32.755 -49.858 32.845 -48.851 ;
      RECT 32.755 -49.545 32.895 -49.375 ;
      RECT 32.755 -48.049 32.845 -47.042 ;
      RECT 32.755 -47.525 32.895 -47.355 ;
      RECT 32.755 -46.628 32.845 -45.621 ;
      RECT 32.755 -46.315 32.895 -46.145 ;
      RECT 32.755 -44.819 32.845 -43.812 ;
      RECT 32.755 -44.295 32.895 -44.125 ;
      RECT 32.755 -43.398 32.845 -42.391 ;
      RECT 32.755 -43.085 32.895 -42.915 ;
      RECT 32.755 -41.589 32.845 -40.582 ;
      RECT 32.755 -41.065 32.895 -40.895 ;
      RECT 32.755 -40.168 32.845 -39.161 ;
      RECT 32.755 -39.855 32.895 -39.685 ;
      RECT 32.755 -38.359 32.845 -37.352 ;
      RECT 32.755 -37.835 32.895 -37.665 ;
      RECT 32.755 -36.938 32.845 -35.931 ;
      RECT 32.755 -36.625 32.895 -36.455 ;
      RECT 32.755 -35.129 32.845 -34.122 ;
      RECT 32.755 -34.605 32.895 -34.435 ;
      RECT 32.755 -33.708 32.845 -32.701 ;
      RECT 32.755 -33.395 32.895 -33.225 ;
      RECT 32.755 -31.899 32.845 -30.892 ;
      RECT 32.755 -31.375 32.895 -31.205 ;
      RECT 32.755 -30.478 32.845 -29.471 ;
      RECT 32.755 -30.165 32.895 -29.995 ;
      RECT 32.755 -28.669 32.845 -27.662 ;
      RECT 32.755 -28.145 32.895 -27.975 ;
      RECT 32.755 -27.248 32.845 -26.241 ;
      RECT 32.755 -26.935 32.895 -26.765 ;
      RECT 32.755 -25.439 32.845 -24.432 ;
      RECT 32.755 -24.915 32.895 -24.745 ;
      RECT 32.755 -24.018 32.845 -23.011 ;
      RECT 32.755 -23.705 32.895 -23.535 ;
      RECT 32.755 -22.209 32.845 -21.202 ;
      RECT 32.755 -21.685 32.895 -21.515 ;
      RECT 32.755 -20.788 32.845 -19.781 ;
      RECT 32.755 -20.475 32.895 -20.305 ;
      RECT 32.755 -18.979 32.845 -17.972 ;
      RECT 32.755 -18.455 32.895 -18.285 ;
      RECT 32.755 -17.558 32.845 -16.551 ;
      RECT 32.755 -17.245 32.895 -17.075 ;
      RECT 32.755 -15.749 32.845 -14.742 ;
      RECT 32.755 -15.225 32.895 -15.055 ;
      RECT 32.755 -14.328 32.845 -13.321 ;
      RECT 32.755 -14.015 32.895 -13.845 ;
      RECT 32.755 -12.519 32.845 -11.512 ;
      RECT 32.755 -11.995 32.895 -11.825 ;
      RECT 32.755 -11.098 32.845 -10.091 ;
      RECT 32.755 -10.785 32.895 -10.615 ;
      RECT 32.755 -9.289 32.845 -8.282 ;
      RECT 32.755 -8.765 32.895 -8.595 ;
      RECT 32.755 -7.868 32.845 -6.861 ;
      RECT 32.755 -7.555 32.895 -7.385 ;
      RECT 32.755 -6.059 32.845 -5.052 ;
      RECT 32.755 -5.535 32.895 -5.365 ;
      RECT 32.755 -4.638 32.845 -3.631 ;
      RECT 32.755 -4.325 32.895 -4.155 ;
      RECT 32.755 -2.829 32.845 -1.822 ;
      RECT 32.755 -2.305 32.895 -2.135 ;
      RECT 32.755 -1.408 32.845 -0.401 ;
      RECT 32.755 -1.095 32.895 -0.925 ;
      RECT 32.755 0.401 32.845 1.408 ;
      RECT 32.755 0.925 32.895 1.095 ;
      RECT 32.085 -111.495 32.255 -111.385 ;
      RECT 28.935 -111.495 32.255 -111.395 ;
      RECT 31.955 -101.538 32.045 -100.53 ;
      RECT 31.905 -100.935 32.045 -100.765 ;
      RECT 31.955 -99.73 32.045 -98.722 ;
      RECT 31.905 -99.495 32.045 -99.325 ;
      RECT 31.955 -98.308 32.045 -97.3 ;
      RECT 31.905 -97.705 32.045 -97.535 ;
      RECT 31.955 -96.5 32.045 -95.492 ;
      RECT 31.905 -96.265 32.045 -96.095 ;
      RECT 31.955 -95.078 32.045 -94.07 ;
      RECT 31.905 -94.475 32.045 -94.305 ;
      RECT 31.955 -93.27 32.045 -92.262 ;
      RECT 31.905 -93.035 32.045 -92.865 ;
      RECT 31.955 -91.848 32.045 -90.84 ;
      RECT 31.905 -91.245 32.045 -91.075 ;
      RECT 31.955 -90.04 32.045 -89.032 ;
      RECT 31.905 -89.805 32.045 -89.635 ;
      RECT 31.955 -88.618 32.045 -87.61 ;
      RECT 31.905 -88.015 32.045 -87.845 ;
      RECT 31.955 -86.81 32.045 -85.802 ;
      RECT 31.905 -86.575 32.045 -86.405 ;
      RECT 31.955 -85.388 32.045 -84.38 ;
      RECT 31.905 -84.785 32.045 -84.615 ;
      RECT 31.955 -83.58 32.045 -82.572 ;
      RECT 31.905 -83.345 32.045 -83.175 ;
      RECT 31.955 -82.158 32.045 -81.15 ;
      RECT 31.905 -81.555 32.045 -81.385 ;
      RECT 31.955 -80.35 32.045 -79.342 ;
      RECT 31.905 -80.115 32.045 -79.945 ;
      RECT 31.955 -78.928 32.045 -77.92 ;
      RECT 31.905 -78.325 32.045 -78.155 ;
      RECT 31.955 -77.12 32.045 -76.112 ;
      RECT 31.905 -76.885 32.045 -76.715 ;
      RECT 31.955 -75.698 32.045 -74.69 ;
      RECT 31.905 -75.095 32.045 -74.925 ;
      RECT 31.955 -73.89 32.045 -72.882 ;
      RECT 31.905 -73.655 32.045 -73.485 ;
      RECT 31.955 -72.468 32.045 -71.46 ;
      RECT 31.905 -71.865 32.045 -71.695 ;
      RECT 31.955 -70.66 32.045 -69.652 ;
      RECT 31.905 -70.425 32.045 -70.255 ;
      RECT 31.955 -69.238 32.045 -68.23 ;
      RECT 31.905 -68.635 32.045 -68.465 ;
      RECT 31.955 -67.43 32.045 -66.422 ;
      RECT 31.905 -67.195 32.045 -67.025 ;
      RECT 31.955 -66.008 32.045 -65 ;
      RECT 31.905 -65.405 32.045 -65.235 ;
      RECT 31.955 -64.2 32.045 -63.192 ;
      RECT 31.905 -63.965 32.045 -63.795 ;
      RECT 31.955 -62.778 32.045 -61.77 ;
      RECT 31.905 -62.175 32.045 -62.005 ;
      RECT 31.955 -60.97 32.045 -59.962 ;
      RECT 31.905 -60.735 32.045 -60.565 ;
      RECT 31.955 -59.548 32.045 -58.54 ;
      RECT 31.905 -58.945 32.045 -58.775 ;
      RECT 31.955 -57.74 32.045 -56.732 ;
      RECT 31.905 -57.505 32.045 -57.335 ;
      RECT 31.955 -56.318 32.045 -55.31 ;
      RECT 31.905 -55.715 32.045 -55.545 ;
      RECT 31.955 -54.51 32.045 -53.502 ;
      RECT 31.905 -54.275 32.045 -54.105 ;
      RECT 31.955 -53.088 32.045 -52.08 ;
      RECT 31.905 -52.485 32.045 -52.315 ;
      RECT 31.955 -51.28 32.045 -50.272 ;
      RECT 31.905 -51.045 32.045 -50.875 ;
      RECT 31.955 -49.858 32.045 -48.85 ;
      RECT 31.905 -49.255 32.045 -49.085 ;
      RECT 31.955 -48.05 32.045 -47.042 ;
      RECT 31.905 -47.815 32.045 -47.645 ;
      RECT 31.955 -46.628 32.045 -45.62 ;
      RECT 31.905 -46.025 32.045 -45.855 ;
      RECT 31.955 -44.82 32.045 -43.812 ;
      RECT 31.905 -44.585 32.045 -44.415 ;
      RECT 31.955 -43.398 32.045 -42.39 ;
      RECT 31.905 -42.795 32.045 -42.625 ;
      RECT 31.955 -41.59 32.045 -40.582 ;
      RECT 31.905 -41.355 32.045 -41.185 ;
      RECT 31.955 -40.168 32.045 -39.16 ;
      RECT 31.905 -39.565 32.045 -39.395 ;
      RECT 31.955 -38.36 32.045 -37.352 ;
      RECT 31.905 -38.125 32.045 -37.955 ;
      RECT 31.955 -36.938 32.045 -35.93 ;
      RECT 31.905 -36.335 32.045 -36.165 ;
      RECT 31.955 -35.13 32.045 -34.122 ;
      RECT 31.905 -34.895 32.045 -34.725 ;
      RECT 31.955 -33.708 32.045 -32.7 ;
      RECT 31.905 -33.105 32.045 -32.935 ;
      RECT 31.955 -31.9 32.045 -30.892 ;
      RECT 31.905 -31.665 32.045 -31.495 ;
      RECT 31.955 -30.478 32.045 -29.47 ;
      RECT 31.905 -29.875 32.045 -29.705 ;
      RECT 31.955 -28.67 32.045 -27.662 ;
      RECT 31.905 -28.435 32.045 -28.265 ;
      RECT 31.955 -27.248 32.045 -26.24 ;
      RECT 31.905 -26.645 32.045 -26.475 ;
      RECT 31.955 -25.44 32.045 -24.432 ;
      RECT 31.905 -25.205 32.045 -25.035 ;
      RECT 31.955 -24.018 32.045 -23.01 ;
      RECT 31.905 -23.415 32.045 -23.245 ;
      RECT 31.955 -22.21 32.045 -21.202 ;
      RECT 31.905 -21.975 32.045 -21.805 ;
      RECT 31.955 -20.788 32.045 -19.78 ;
      RECT 31.905 -20.185 32.045 -20.015 ;
      RECT 31.955 -18.98 32.045 -17.972 ;
      RECT 31.905 -18.745 32.045 -18.575 ;
      RECT 31.955 -17.558 32.045 -16.55 ;
      RECT 31.905 -16.955 32.045 -16.785 ;
      RECT 31.955 -15.75 32.045 -14.742 ;
      RECT 31.905 -15.515 32.045 -15.345 ;
      RECT 31.955 -14.328 32.045 -13.32 ;
      RECT 31.905 -13.725 32.045 -13.555 ;
      RECT 31.955 -12.52 32.045 -11.512 ;
      RECT 31.905 -12.285 32.045 -12.115 ;
      RECT 31.955 -11.098 32.045 -10.09 ;
      RECT 31.905 -10.495 32.045 -10.325 ;
      RECT 31.955 -9.29 32.045 -8.282 ;
      RECT 31.905 -9.055 32.045 -8.885 ;
      RECT 31.955 -7.868 32.045 -6.86 ;
      RECT 31.905 -7.265 32.045 -7.095 ;
      RECT 31.955 -6.06 32.045 -5.052 ;
      RECT 31.905 -5.825 32.045 -5.655 ;
      RECT 31.955 -4.638 32.045 -3.63 ;
      RECT 31.905 -4.035 32.045 -3.865 ;
      RECT 31.955 -2.83 32.045 -1.822 ;
      RECT 31.905 -2.595 32.045 -2.425 ;
      RECT 31.955 -1.408 32.045 -0.4 ;
      RECT 31.905 -0.805 32.045 -0.635 ;
      RECT 31.955 0.4 32.045 1.408 ;
      RECT 31.905 0.635 32.045 0.805 ;
      RECT 31.555 -101.538 31.645 -100.531 ;
      RECT 31.555 -101.225 31.695 -101.055 ;
      RECT 31.555 -99.729 31.645 -98.722 ;
      RECT 31.555 -99.205 31.695 -99.035 ;
      RECT 31.555 -98.308 31.645 -97.301 ;
      RECT 31.555 -97.995 31.695 -97.825 ;
      RECT 31.555 -96.499 31.645 -95.492 ;
      RECT 31.555 -95.975 31.695 -95.805 ;
      RECT 31.555 -95.078 31.645 -94.071 ;
      RECT 31.555 -94.765 31.695 -94.595 ;
      RECT 31.555 -93.269 31.645 -92.262 ;
      RECT 31.555 -92.745 31.695 -92.575 ;
      RECT 31.555 -91.848 31.645 -90.841 ;
      RECT 31.555 -91.535 31.695 -91.365 ;
      RECT 31.555 -90.039 31.645 -89.032 ;
      RECT 31.555 -89.515 31.695 -89.345 ;
      RECT 31.555 -88.618 31.645 -87.611 ;
      RECT 31.555 -88.305 31.695 -88.135 ;
      RECT 31.555 -86.809 31.645 -85.802 ;
      RECT 31.555 -86.285 31.695 -86.115 ;
      RECT 31.555 -85.388 31.645 -84.381 ;
      RECT 31.555 -85.075 31.695 -84.905 ;
      RECT 31.555 -83.579 31.645 -82.572 ;
      RECT 31.555 -83.055 31.695 -82.885 ;
      RECT 31.555 -82.158 31.645 -81.151 ;
      RECT 31.555 -81.845 31.695 -81.675 ;
      RECT 31.555 -80.349 31.645 -79.342 ;
      RECT 31.555 -79.825 31.695 -79.655 ;
      RECT 31.555 -78.928 31.645 -77.921 ;
      RECT 31.555 -78.615 31.695 -78.445 ;
      RECT 31.555 -77.119 31.645 -76.112 ;
      RECT 31.555 -76.595 31.695 -76.425 ;
      RECT 31.555 -75.698 31.645 -74.691 ;
      RECT 31.555 -75.385 31.695 -75.215 ;
      RECT 31.555 -73.889 31.645 -72.882 ;
      RECT 31.555 -73.365 31.695 -73.195 ;
      RECT 31.555 -72.468 31.645 -71.461 ;
      RECT 31.555 -72.155 31.695 -71.985 ;
      RECT 31.555 -70.659 31.645 -69.652 ;
      RECT 31.555 -70.135 31.695 -69.965 ;
      RECT 31.555 -69.238 31.645 -68.231 ;
      RECT 31.555 -68.925 31.695 -68.755 ;
      RECT 31.555 -67.429 31.645 -66.422 ;
      RECT 31.555 -66.905 31.695 -66.735 ;
      RECT 31.555 -66.008 31.645 -65.001 ;
      RECT 31.555 -65.695 31.695 -65.525 ;
      RECT 31.555 -64.199 31.645 -63.192 ;
      RECT 31.555 -63.675 31.695 -63.505 ;
      RECT 31.555 -62.778 31.645 -61.771 ;
      RECT 31.555 -62.465 31.695 -62.295 ;
      RECT 31.555 -60.969 31.645 -59.962 ;
      RECT 31.555 -60.445 31.695 -60.275 ;
      RECT 31.555 -59.548 31.645 -58.541 ;
      RECT 31.555 -59.235 31.695 -59.065 ;
      RECT 31.555 -57.739 31.645 -56.732 ;
      RECT 31.555 -57.215 31.695 -57.045 ;
      RECT 31.555 -56.318 31.645 -55.311 ;
      RECT 31.555 -56.005 31.695 -55.835 ;
      RECT 31.555 -54.509 31.645 -53.502 ;
      RECT 31.555 -53.985 31.695 -53.815 ;
      RECT 31.555 -53.088 31.645 -52.081 ;
      RECT 31.555 -52.775 31.695 -52.605 ;
      RECT 31.555 -51.279 31.645 -50.272 ;
      RECT 31.555 -50.755 31.695 -50.585 ;
      RECT 31.555 -49.858 31.645 -48.851 ;
      RECT 31.555 -49.545 31.695 -49.375 ;
      RECT 31.555 -48.049 31.645 -47.042 ;
      RECT 31.555 -47.525 31.695 -47.355 ;
      RECT 31.555 -46.628 31.645 -45.621 ;
      RECT 31.555 -46.315 31.695 -46.145 ;
      RECT 31.555 -44.819 31.645 -43.812 ;
      RECT 31.555 -44.295 31.695 -44.125 ;
      RECT 31.555 -43.398 31.645 -42.391 ;
      RECT 31.555 -43.085 31.695 -42.915 ;
      RECT 31.555 -41.589 31.645 -40.582 ;
      RECT 31.555 -41.065 31.695 -40.895 ;
      RECT 31.555 -40.168 31.645 -39.161 ;
      RECT 31.555 -39.855 31.695 -39.685 ;
      RECT 31.555 -38.359 31.645 -37.352 ;
      RECT 31.555 -37.835 31.695 -37.665 ;
      RECT 31.555 -36.938 31.645 -35.931 ;
      RECT 31.555 -36.625 31.695 -36.455 ;
      RECT 31.555 -35.129 31.645 -34.122 ;
      RECT 31.555 -34.605 31.695 -34.435 ;
      RECT 31.555 -33.708 31.645 -32.701 ;
      RECT 31.555 -33.395 31.695 -33.225 ;
      RECT 31.555 -31.899 31.645 -30.892 ;
      RECT 31.555 -31.375 31.695 -31.205 ;
      RECT 31.555 -30.478 31.645 -29.471 ;
      RECT 31.555 -30.165 31.695 -29.995 ;
      RECT 31.555 -28.669 31.645 -27.662 ;
      RECT 31.555 -28.145 31.695 -27.975 ;
      RECT 31.555 -27.248 31.645 -26.241 ;
      RECT 31.555 -26.935 31.695 -26.765 ;
      RECT 31.555 -25.439 31.645 -24.432 ;
      RECT 31.555 -24.915 31.695 -24.745 ;
      RECT 31.555 -24.018 31.645 -23.011 ;
      RECT 31.555 -23.705 31.695 -23.535 ;
      RECT 31.555 -22.209 31.645 -21.202 ;
      RECT 31.555 -21.685 31.695 -21.515 ;
      RECT 31.555 -20.788 31.645 -19.781 ;
      RECT 31.555 -20.475 31.695 -20.305 ;
      RECT 31.555 -18.979 31.645 -17.972 ;
      RECT 31.555 -18.455 31.695 -18.285 ;
      RECT 31.555 -17.558 31.645 -16.551 ;
      RECT 31.555 -17.245 31.695 -17.075 ;
      RECT 31.555 -15.749 31.645 -14.742 ;
      RECT 31.555 -15.225 31.695 -15.055 ;
      RECT 31.555 -14.328 31.645 -13.321 ;
      RECT 31.555 -14.015 31.695 -13.845 ;
      RECT 31.555 -12.519 31.645 -11.512 ;
      RECT 31.555 -11.995 31.695 -11.825 ;
      RECT 31.555 -11.098 31.645 -10.091 ;
      RECT 31.555 -10.785 31.695 -10.615 ;
      RECT 31.555 -9.289 31.645 -8.282 ;
      RECT 31.555 -8.765 31.695 -8.595 ;
      RECT 31.555 -7.868 31.645 -6.861 ;
      RECT 31.555 -7.555 31.695 -7.385 ;
      RECT 31.555 -6.059 31.645 -5.052 ;
      RECT 31.555 -5.535 31.695 -5.365 ;
      RECT 31.555 -4.638 31.645 -3.631 ;
      RECT 31.555 -4.325 31.695 -4.155 ;
      RECT 31.555 -2.829 31.645 -1.822 ;
      RECT 31.555 -2.305 31.695 -2.135 ;
      RECT 31.555 -1.408 31.645 -0.401 ;
      RECT 31.555 -1.095 31.695 -0.925 ;
      RECT 31.555 0.401 31.645 1.408 ;
      RECT 31.555 0.925 31.695 1.095 ;
      RECT 29.705 -111.685 31.185 -111.585 ;
      RECT 29.705 -112.055 29.805 -111.585 ;
      RECT 29.51 -114.395 31.085 -114.275 ;
      RECT 30.985 -114.895 31.085 -114.275 ;
      RECT 30.39 -114.895 30.49 -114.275 ;
      RECT 29.51 -114.85 29.61 -114.275 ;
      RECT 30.755 -101.538 30.845 -100.53 ;
      RECT 30.705 -100.935 30.845 -100.765 ;
      RECT 30.755 -99.73 30.845 -98.722 ;
      RECT 30.705 -99.495 30.845 -99.325 ;
      RECT 30.755 -98.308 30.845 -97.3 ;
      RECT 30.705 -97.705 30.845 -97.535 ;
      RECT 30.755 -96.5 30.845 -95.492 ;
      RECT 30.705 -96.265 30.845 -96.095 ;
      RECT 30.755 -95.078 30.845 -94.07 ;
      RECT 30.705 -94.475 30.845 -94.305 ;
      RECT 30.755 -93.27 30.845 -92.262 ;
      RECT 30.705 -93.035 30.845 -92.865 ;
      RECT 30.755 -91.848 30.845 -90.84 ;
      RECT 30.705 -91.245 30.845 -91.075 ;
      RECT 30.755 -90.04 30.845 -89.032 ;
      RECT 30.705 -89.805 30.845 -89.635 ;
      RECT 30.755 -88.618 30.845 -87.61 ;
      RECT 30.705 -88.015 30.845 -87.845 ;
      RECT 30.755 -86.81 30.845 -85.802 ;
      RECT 30.705 -86.575 30.845 -86.405 ;
      RECT 30.755 -85.388 30.845 -84.38 ;
      RECT 30.705 -84.785 30.845 -84.615 ;
      RECT 30.755 -83.58 30.845 -82.572 ;
      RECT 30.705 -83.345 30.845 -83.175 ;
      RECT 30.755 -82.158 30.845 -81.15 ;
      RECT 30.705 -81.555 30.845 -81.385 ;
      RECT 30.755 -80.35 30.845 -79.342 ;
      RECT 30.705 -80.115 30.845 -79.945 ;
      RECT 30.755 -78.928 30.845 -77.92 ;
      RECT 30.705 -78.325 30.845 -78.155 ;
      RECT 30.755 -77.12 30.845 -76.112 ;
      RECT 30.705 -76.885 30.845 -76.715 ;
      RECT 30.755 -75.698 30.845 -74.69 ;
      RECT 30.705 -75.095 30.845 -74.925 ;
      RECT 30.755 -73.89 30.845 -72.882 ;
      RECT 30.705 -73.655 30.845 -73.485 ;
      RECT 30.755 -72.468 30.845 -71.46 ;
      RECT 30.705 -71.865 30.845 -71.695 ;
      RECT 30.755 -70.66 30.845 -69.652 ;
      RECT 30.705 -70.425 30.845 -70.255 ;
      RECT 30.755 -69.238 30.845 -68.23 ;
      RECT 30.705 -68.635 30.845 -68.465 ;
      RECT 30.755 -67.43 30.845 -66.422 ;
      RECT 30.705 -67.195 30.845 -67.025 ;
      RECT 30.755 -66.008 30.845 -65 ;
      RECT 30.705 -65.405 30.845 -65.235 ;
      RECT 30.755 -64.2 30.845 -63.192 ;
      RECT 30.705 -63.965 30.845 -63.795 ;
      RECT 30.755 -62.778 30.845 -61.77 ;
      RECT 30.705 -62.175 30.845 -62.005 ;
      RECT 30.755 -60.97 30.845 -59.962 ;
      RECT 30.705 -60.735 30.845 -60.565 ;
      RECT 30.755 -59.548 30.845 -58.54 ;
      RECT 30.705 -58.945 30.845 -58.775 ;
      RECT 30.755 -57.74 30.845 -56.732 ;
      RECT 30.705 -57.505 30.845 -57.335 ;
      RECT 30.755 -56.318 30.845 -55.31 ;
      RECT 30.705 -55.715 30.845 -55.545 ;
      RECT 30.755 -54.51 30.845 -53.502 ;
      RECT 30.705 -54.275 30.845 -54.105 ;
      RECT 30.755 -53.088 30.845 -52.08 ;
      RECT 30.705 -52.485 30.845 -52.315 ;
      RECT 30.755 -51.28 30.845 -50.272 ;
      RECT 30.705 -51.045 30.845 -50.875 ;
      RECT 30.755 -49.858 30.845 -48.85 ;
      RECT 30.705 -49.255 30.845 -49.085 ;
      RECT 30.755 -48.05 30.845 -47.042 ;
      RECT 30.705 -47.815 30.845 -47.645 ;
      RECT 30.755 -46.628 30.845 -45.62 ;
      RECT 30.705 -46.025 30.845 -45.855 ;
      RECT 30.755 -44.82 30.845 -43.812 ;
      RECT 30.705 -44.585 30.845 -44.415 ;
      RECT 30.755 -43.398 30.845 -42.39 ;
      RECT 30.705 -42.795 30.845 -42.625 ;
      RECT 30.755 -41.59 30.845 -40.582 ;
      RECT 30.705 -41.355 30.845 -41.185 ;
      RECT 30.755 -40.168 30.845 -39.16 ;
      RECT 30.705 -39.565 30.845 -39.395 ;
      RECT 30.755 -38.36 30.845 -37.352 ;
      RECT 30.705 -38.125 30.845 -37.955 ;
      RECT 30.755 -36.938 30.845 -35.93 ;
      RECT 30.705 -36.335 30.845 -36.165 ;
      RECT 30.755 -35.13 30.845 -34.122 ;
      RECT 30.705 -34.895 30.845 -34.725 ;
      RECT 30.755 -33.708 30.845 -32.7 ;
      RECT 30.705 -33.105 30.845 -32.935 ;
      RECT 30.755 -31.9 30.845 -30.892 ;
      RECT 30.705 -31.665 30.845 -31.495 ;
      RECT 30.755 -30.478 30.845 -29.47 ;
      RECT 30.705 -29.875 30.845 -29.705 ;
      RECT 30.755 -28.67 30.845 -27.662 ;
      RECT 30.705 -28.435 30.845 -28.265 ;
      RECT 30.755 -27.248 30.845 -26.24 ;
      RECT 30.705 -26.645 30.845 -26.475 ;
      RECT 30.755 -25.44 30.845 -24.432 ;
      RECT 30.705 -25.205 30.845 -25.035 ;
      RECT 30.755 -24.018 30.845 -23.01 ;
      RECT 30.705 -23.415 30.845 -23.245 ;
      RECT 30.755 -22.21 30.845 -21.202 ;
      RECT 30.705 -21.975 30.845 -21.805 ;
      RECT 30.755 -20.788 30.845 -19.78 ;
      RECT 30.705 -20.185 30.845 -20.015 ;
      RECT 30.755 -18.98 30.845 -17.972 ;
      RECT 30.705 -18.745 30.845 -18.575 ;
      RECT 30.755 -17.558 30.845 -16.55 ;
      RECT 30.705 -16.955 30.845 -16.785 ;
      RECT 30.755 -15.75 30.845 -14.742 ;
      RECT 30.705 -15.515 30.845 -15.345 ;
      RECT 30.755 -14.328 30.845 -13.32 ;
      RECT 30.705 -13.725 30.845 -13.555 ;
      RECT 30.755 -12.52 30.845 -11.512 ;
      RECT 30.705 -12.285 30.845 -12.115 ;
      RECT 30.755 -11.098 30.845 -10.09 ;
      RECT 30.705 -10.495 30.845 -10.325 ;
      RECT 30.755 -9.29 30.845 -8.282 ;
      RECT 30.705 -9.055 30.845 -8.885 ;
      RECT 30.755 -7.868 30.845 -6.86 ;
      RECT 30.705 -7.265 30.845 -7.095 ;
      RECT 30.755 -6.06 30.845 -5.052 ;
      RECT 30.705 -5.825 30.845 -5.655 ;
      RECT 30.755 -4.638 30.845 -3.63 ;
      RECT 30.705 -4.035 30.845 -3.865 ;
      RECT 30.755 -2.83 30.845 -1.822 ;
      RECT 30.705 -2.595 30.845 -2.425 ;
      RECT 30.755 -1.408 30.845 -0.4 ;
      RECT 30.705 -0.805 30.845 -0.635 ;
      RECT 30.755 0.4 30.845 1.408 ;
      RECT 30.705 0.635 30.845 0.805 ;
      RECT 30.63 -114.685 30.805 -114.515 ;
      RECT 30.705 -114.895 30.805 -114.515 ;
      RECT 29.745 -113.555 29.845 -113.09 ;
      RECT 30.11 -113.555 30.21 -113.1 ;
      RECT 29.745 -113.555 30.59 -113.385 ;
      RECT 30.355 -101.538 30.445 -100.531 ;
      RECT 30.355 -101.225 30.495 -101.055 ;
      RECT 30.355 -99.729 30.445 -98.722 ;
      RECT 30.355 -99.205 30.495 -99.035 ;
      RECT 30.355 -98.308 30.445 -97.301 ;
      RECT 30.355 -97.995 30.495 -97.825 ;
      RECT 30.355 -96.499 30.445 -95.492 ;
      RECT 30.355 -95.975 30.495 -95.805 ;
      RECT 30.355 -95.078 30.445 -94.071 ;
      RECT 30.355 -94.765 30.495 -94.595 ;
      RECT 30.355 -93.269 30.445 -92.262 ;
      RECT 30.355 -92.745 30.495 -92.575 ;
      RECT 30.355 -91.848 30.445 -90.841 ;
      RECT 30.355 -91.535 30.495 -91.365 ;
      RECT 30.355 -90.039 30.445 -89.032 ;
      RECT 30.355 -89.515 30.495 -89.345 ;
      RECT 30.355 -88.618 30.445 -87.611 ;
      RECT 30.355 -88.305 30.495 -88.135 ;
      RECT 30.355 -86.809 30.445 -85.802 ;
      RECT 30.355 -86.285 30.495 -86.115 ;
      RECT 30.355 -85.388 30.445 -84.381 ;
      RECT 30.355 -85.075 30.495 -84.905 ;
      RECT 30.355 -83.579 30.445 -82.572 ;
      RECT 30.355 -83.055 30.495 -82.885 ;
      RECT 30.355 -82.158 30.445 -81.151 ;
      RECT 30.355 -81.845 30.495 -81.675 ;
      RECT 30.355 -80.349 30.445 -79.342 ;
      RECT 30.355 -79.825 30.495 -79.655 ;
      RECT 30.355 -78.928 30.445 -77.921 ;
      RECT 30.355 -78.615 30.495 -78.445 ;
      RECT 30.355 -77.119 30.445 -76.112 ;
      RECT 30.355 -76.595 30.495 -76.425 ;
      RECT 30.355 -75.698 30.445 -74.691 ;
      RECT 30.355 -75.385 30.495 -75.215 ;
      RECT 30.355 -73.889 30.445 -72.882 ;
      RECT 30.355 -73.365 30.495 -73.195 ;
      RECT 30.355 -72.468 30.445 -71.461 ;
      RECT 30.355 -72.155 30.495 -71.985 ;
      RECT 30.355 -70.659 30.445 -69.652 ;
      RECT 30.355 -70.135 30.495 -69.965 ;
      RECT 30.355 -69.238 30.445 -68.231 ;
      RECT 30.355 -68.925 30.495 -68.755 ;
      RECT 30.355 -67.429 30.445 -66.422 ;
      RECT 30.355 -66.905 30.495 -66.735 ;
      RECT 30.355 -66.008 30.445 -65.001 ;
      RECT 30.355 -65.695 30.495 -65.525 ;
      RECT 30.355 -64.199 30.445 -63.192 ;
      RECT 30.355 -63.675 30.495 -63.505 ;
      RECT 30.355 -62.778 30.445 -61.771 ;
      RECT 30.355 -62.465 30.495 -62.295 ;
      RECT 30.355 -60.969 30.445 -59.962 ;
      RECT 30.355 -60.445 30.495 -60.275 ;
      RECT 30.355 -59.548 30.445 -58.541 ;
      RECT 30.355 -59.235 30.495 -59.065 ;
      RECT 30.355 -57.739 30.445 -56.732 ;
      RECT 30.355 -57.215 30.495 -57.045 ;
      RECT 30.355 -56.318 30.445 -55.311 ;
      RECT 30.355 -56.005 30.495 -55.835 ;
      RECT 30.355 -54.509 30.445 -53.502 ;
      RECT 30.355 -53.985 30.495 -53.815 ;
      RECT 30.355 -53.088 30.445 -52.081 ;
      RECT 30.355 -52.775 30.495 -52.605 ;
      RECT 30.355 -51.279 30.445 -50.272 ;
      RECT 30.355 -50.755 30.495 -50.585 ;
      RECT 30.355 -49.858 30.445 -48.851 ;
      RECT 30.355 -49.545 30.495 -49.375 ;
      RECT 30.355 -48.049 30.445 -47.042 ;
      RECT 30.355 -47.525 30.495 -47.355 ;
      RECT 30.355 -46.628 30.445 -45.621 ;
      RECT 30.355 -46.315 30.495 -46.145 ;
      RECT 30.355 -44.819 30.445 -43.812 ;
      RECT 30.355 -44.295 30.495 -44.125 ;
      RECT 30.355 -43.398 30.445 -42.391 ;
      RECT 30.355 -43.085 30.495 -42.915 ;
      RECT 30.355 -41.589 30.445 -40.582 ;
      RECT 30.355 -41.065 30.495 -40.895 ;
      RECT 30.355 -40.168 30.445 -39.161 ;
      RECT 30.355 -39.855 30.495 -39.685 ;
      RECT 30.355 -38.359 30.445 -37.352 ;
      RECT 30.355 -37.835 30.495 -37.665 ;
      RECT 30.355 -36.938 30.445 -35.931 ;
      RECT 30.355 -36.625 30.495 -36.455 ;
      RECT 30.355 -35.129 30.445 -34.122 ;
      RECT 30.355 -34.605 30.495 -34.435 ;
      RECT 30.355 -33.708 30.445 -32.701 ;
      RECT 30.355 -33.395 30.495 -33.225 ;
      RECT 30.355 -31.899 30.445 -30.892 ;
      RECT 30.355 -31.375 30.495 -31.205 ;
      RECT 30.355 -30.478 30.445 -29.471 ;
      RECT 30.355 -30.165 30.495 -29.995 ;
      RECT 30.355 -28.669 30.445 -27.662 ;
      RECT 30.355 -28.145 30.495 -27.975 ;
      RECT 30.355 -27.248 30.445 -26.241 ;
      RECT 30.355 -26.935 30.495 -26.765 ;
      RECT 30.355 -25.439 30.445 -24.432 ;
      RECT 30.355 -24.915 30.495 -24.745 ;
      RECT 30.355 -24.018 30.445 -23.011 ;
      RECT 30.355 -23.705 30.495 -23.535 ;
      RECT 30.355 -22.209 30.445 -21.202 ;
      RECT 30.355 -21.685 30.495 -21.515 ;
      RECT 30.355 -20.788 30.445 -19.781 ;
      RECT 30.355 -20.475 30.495 -20.305 ;
      RECT 30.355 -18.979 30.445 -17.972 ;
      RECT 30.355 -18.455 30.495 -18.285 ;
      RECT 30.355 -17.558 30.445 -16.551 ;
      RECT 30.355 -17.245 30.495 -17.075 ;
      RECT 30.355 -15.749 30.445 -14.742 ;
      RECT 30.355 -15.225 30.495 -15.055 ;
      RECT 30.355 -14.328 30.445 -13.321 ;
      RECT 30.355 -14.015 30.495 -13.845 ;
      RECT 30.355 -12.519 30.445 -11.512 ;
      RECT 30.355 -11.995 30.495 -11.825 ;
      RECT 30.355 -11.098 30.445 -10.091 ;
      RECT 30.355 -10.785 30.495 -10.615 ;
      RECT 30.355 -9.289 30.445 -8.282 ;
      RECT 30.355 -8.765 30.495 -8.595 ;
      RECT 30.355 -7.868 30.445 -6.861 ;
      RECT 30.355 -7.555 30.495 -7.385 ;
      RECT 30.355 -6.059 30.445 -5.052 ;
      RECT 30.355 -5.535 30.495 -5.365 ;
      RECT 30.355 -4.638 30.445 -3.631 ;
      RECT 30.355 -4.325 30.495 -4.155 ;
      RECT 30.355 -2.829 30.445 -1.822 ;
      RECT 30.355 -2.305 30.495 -2.135 ;
      RECT 30.355 -1.408 30.445 -0.401 ;
      RECT 30.355 -1.095 30.495 -0.925 ;
      RECT 30.355 0.401 30.445 1.408 ;
      RECT 30.355 0.925 30.495 1.095 ;
      RECT 30.04 -114.685 30.21 -114.515 ;
      RECT 30.11 -114.895 30.21 -114.515 ;
      RECT 29.555 -101.538 29.645 -100.53 ;
      RECT 29.505 -100.935 29.645 -100.765 ;
      RECT 29.555 -99.73 29.645 -98.722 ;
      RECT 29.505 -99.495 29.645 -99.325 ;
      RECT 29.555 -98.308 29.645 -97.3 ;
      RECT 29.505 -97.705 29.645 -97.535 ;
      RECT 29.555 -96.5 29.645 -95.492 ;
      RECT 29.505 -96.265 29.645 -96.095 ;
      RECT 29.555 -95.078 29.645 -94.07 ;
      RECT 29.505 -94.475 29.645 -94.305 ;
      RECT 29.555 -93.27 29.645 -92.262 ;
      RECT 29.505 -93.035 29.645 -92.865 ;
      RECT 29.555 -91.848 29.645 -90.84 ;
      RECT 29.505 -91.245 29.645 -91.075 ;
      RECT 29.555 -90.04 29.645 -89.032 ;
      RECT 29.505 -89.805 29.645 -89.635 ;
      RECT 29.555 -88.618 29.645 -87.61 ;
      RECT 29.505 -88.015 29.645 -87.845 ;
      RECT 29.555 -86.81 29.645 -85.802 ;
      RECT 29.505 -86.575 29.645 -86.405 ;
      RECT 29.555 -85.388 29.645 -84.38 ;
      RECT 29.505 -84.785 29.645 -84.615 ;
      RECT 29.555 -83.58 29.645 -82.572 ;
      RECT 29.505 -83.345 29.645 -83.175 ;
      RECT 29.555 -82.158 29.645 -81.15 ;
      RECT 29.505 -81.555 29.645 -81.385 ;
      RECT 29.555 -80.35 29.645 -79.342 ;
      RECT 29.505 -80.115 29.645 -79.945 ;
      RECT 29.555 -78.928 29.645 -77.92 ;
      RECT 29.505 -78.325 29.645 -78.155 ;
      RECT 29.555 -77.12 29.645 -76.112 ;
      RECT 29.505 -76.885 29.645 -76.715 ;
      RECT 29.555 -75.698 29.645 -74.69 ;
      RECT 29.505 -75.095 29.645 -74.925 ;
      RECT 29.555 -73.89 29.645 -72.882 ;
      RECT 29.505 -73.655 29.645 -73.485 ;
      RECT 29.555 -72.468 29.645 -71.46 ;
      RECT 29.505 -71.865 29.645 -71.695 ;
      RECT 29.555 -70.66 29.645 -69.652 ;
      RECT 29.505 -70.425 29.645 -70.255 ;
      RECT 29.555 -69.238 29.645 -68.23 ;
      RECT 29.505 -68.635 29.645 -68.465 ;
      RECT 29.555 -67.43 29.645 -66.422 ;
      RECT 29.505 -67.195 29.645 -67.025 ;
      RECT 29.555 -66.008 29.645 -65 ;
      RECT 29.505 -65.405 29.645 -65.235 ;
      RECT 29.555 -64.2 29.645 -63.192 ;
      RECT 29.505 -63.965 29.645 -63.795 ;
      RECT 29.555 -62.778 29.645 -61.77 ;
      RECT 29.505 -62.175 29.645 -62.005 ;
      RECT 29.555 -60.97 29.645 -59.962 ;
      RECT 29.505 -60.735 29.645 -60.565 ;
      RECT 29.555 -59.548 29.645 -58.54 ;
      RECT 29.505 -58.945 29.645 -58.775 ;
      RECT 29.555 -57.74 29.645 -56.732 ;
      RECT 29.505 -57.505 29.645 -57.335 ;
      RECT 29.555 -56.318 29.645 -55.31 ;
      RECT 29.505 -55.715 29.645 -55.545 ;
      RECT 29.555 -54.51 29.645 -53.502 ;
      RECT 29.505 -54.275 29.645 -54.105 ;
      RECT 29.555 -53.088 29.645 -52.08 ;
      RECT 29.505 -52.485 29.645 -52.315 ;
      RECT 29.555 -51.28 29.645 -50.272 ;
      RECT 29.505 -51.045 29.645 -50.875 ;
      RECT 29.555 -49.858 29.645 -48.85 ;
      RECT 29.505 -49.255 29.645 -49.085 ;
      RECT 29.555 -48.05 29.645 -47.042 ;
      RECT 29.505 -47.815 29.645 -47.645 ;
      RECT 29.555 -46.628 29.645 -45.62 ;
      RECT 29.505 -46.025 29.645 -45.855 ;
      RECT 29.555 -44.82 29.645 -43.812 ;
      RECT 29.505 -44.585 29.645 -44.415 ;
      RECT 29.555 -43.398 29.645 -42.39 ;
      RECT 29.505 -42.795 29.645 -42.625 ;
      RECT 29.555 -41.59 29.645 -40.582 ;
      RECT 29.505 -41.355 29.645 -41.185 ;
      RECT 29.555 -40.168 29.645 -39.16 ;
      RECT 29.505 -39.565 29.645 -39.395 ;
      RECT 29.555 -38.36 29.645 -37.352 ;
      RECT 29.505 -38.125 29.645 -37.955 ;
      RECT 29.555 -36.938 29.645 -35.93 ;
      RECT 29.505 -36.335 29.645 -36.165 ;
      RECT 29.555 -35.13 29.645 -34.122 ;
      RECT 29.505 -34.895 29.645 -34.725 ;
      RECT 29.555 -33.708 29.645 -32.7 ;
      RECT 29.505 -33.105 29.645 -32.935 ;
      RECT 29.555 -31.9 29.645 -30.892 ;
      RECT 29.505 -31.665 29.645 -31.495 ;
      RECT 29.555 -30.478 29.645 -29.47 ;
      RECT 29.505 -29.875 29.645 -29.705 ;
      RECT 29.555 -28.67 29.645 -27.662 ;
      RECT 29.505 -28.435 29.645 -28.265 ;
      RECT 29.555 -27.248 29.645 -26.24 ;
      RECT 29.505 -26.645 29.645 -26.475 ;
      RECT 29.555 -25.44 29.645 -24.432 ;
      RECT 29.505 -25.205 29.645 -25.035 ;
      RECT 29.555 -24.018 29.645 -23.01 ;
      RECT 29.505 -23.415 29.645 -23.245 ;
      RECT 29.555 -22.21 29.645 -21.202 ;
      RECT 29.505 -21.975 29.645 -21.805 ;
      RECT 29.555 -20.788 29.645 -19.78 ;
      RECT 29.505 -20.185 29.645 -20.015 ;
      RECT 29.555 -18.98 29.645 -17.972 ;
      RECT 29.505 -18.745 29.645 -18.575 ;
      RECT 29.555 -17.558 29.645 -16.55 ;
      RECT 29.505 -16.955 29.645 -16.785 ;
      RECT 29.555 -15.75 29.645 -14.742 ;
      RECT 29.505 -15.515 29.645 -15.345 ;
      RECT 29.555 -14.328 29.645 -13.32 ;
      RECT 29.505 -13.725 29.645 -13.555 ;
      RECT 29.555 -12.52 29.645 -11.512 ;
      RECT 29.505 -12.285 29.645 -12.115 ;
      RECT 29.555 -11.098 29.645 -10.09 ;
      RECT 29.505 -10.495 29.645 -10.325 ;
      RECT 29.555 -9.29 29.645 -8.282 ;
      RECT 29.505 -9.055 29.645 -8.885 ;
      RECT 29.555 -7.868 29.645 -6.86 ;
      RECT 29.505 -7.265 29.645 -7.095 ;
      RECT 29.555 -6.06 29.645 -5.052 ;
      RECT 29.505 -5.825 29.645 -5.655 ;
      RECT 29.555 -4.638 29.645 -3.63 ;
      RECT 29.505 -4.035 29.645 -3.865 ;
      RECT 29.555 -2.83 29.645 -1.822 ;
      RECT 29.505 -2.595 29.645 -2.425 ;
      RECT 29.555 -1.408 29.645 -0.4 ;
      RECT 29.505 -0.805 29.645 -0.635 ;
      RECT 29.555 0.4 29.645 1.408 ;
      RECT 29.505 0.635 29.645 0.805 ;
      RECT 29.155 -101.538 29.245 -100.531 ;
      RECT 29.155 -101.225 29.295 -101.055 ;
      RECT 29.155 -99.729 29.245 -98.722 ;
      RECT 29.155 -99.205 29.295 -99.035 ;
      RECT 29.155 -98.308 29.245 -97.301 ;
      RECT 29.155 -97.995 29.295 -97.825 ;
      RECT 29.155 -96.499 29.245 -95.492 ;
      RECT 29.155 -95.975 29.295 -95.805 ;
      RECT 29.155 -95.078 29.245 -94.071 ;
      RECT 29.155 -94.765 29.295 -94.595 ;
      RECT 29.155 -93.269 29.245 -92.262 ;
      RECT 29.155 -92.745 29.295 -92.575 ;
      RECT 29.155 -91.848 29.245 -90.841 ;
      RECT 29.155 -91.535 29.295 -91.365 ;
      RECT 29.155 -90.039 29.245 -89.032 ;
      RECT 29.155 -89.515 29.295 -89.345 ;
      RECT 29.155 -88.618 29.245 -87.611 ;
      RECT 29.155 -88.305 29.295 -88.135 ;
      RECT 29.155 -86.809 29.245 -85.802 ;
      RECT 29.155 -86.285 29.295 -86.115 ;
      RECT 29.155 -85.388 29.245 -84.381 ;
      RECT 29.155 -85.075 29.295 -84.905 ;
      RECT 29.155 -83.579 29.245 -82.572 ;
      RECT 29.155 -83.055 29.295 -82.885 ;
      RECT 29.155 -82.158 29.245 -81.151 ;
      RECT 29.155 -81.845 29.295 -81.675 ;
      RECT 29.155 -80.349 29.245 -79.342 ;
      RECT 29.155 -79.825 29.295 -79.655 ;
      RECT 29.155 -78.928 29.245 -77.921 ;
      RECT 29.155 -78.615 29.295 -78.445 ;
      RECT 29.155 -77.119 29.245 -76.112 ;
      RECT 29.155 -76.595 29.295 -76.425 ;
      RECT 29.155 -75.698 29.245 -74.691 ;
      RECT 29.155 -75.385 29.295 -75.215 ;
      RECT 29.155 -73.889 29.245 -72.882 ;
      RECT 29.155 -73.365 29.295 -73.195 ;
      RECT 29.155 -72.468 29.245 -71.461 ;
      RECT 29.155 -72.155 29.295 -71.985 ;
      RECT 29.155 -70.659 29.245 -69.652 ;
      RECT 29.155 -70.135 29.295 -69.965 ;
      RECT 29.155 -69.238 29.245 -68.231 ;
      RECT 29.155 -68.925 29.295 -68.755 ;
      RECT 29.155 -67.429 29.245 -66.422 ;
      RECT 29.155 -66.905 29.295 -66.735 ;
      RECT 29.155 -66.008 29.245 -65.001 ;
      RECT 29.155 -65.695 29.295 -65.525 ;
      RECT 29.155 -64.199 29.245 -63.192 ;
      RECT 29.155 -63.675 29.295 -63.505 ;
      RECT 29.155 -62.778 29.245 -61.771 ;
      RECT 29.155 -62.465 29.295 -62.295 ;
      RECT 29.155 -60.969 29.245 -59.962 ;
      RECT 29.155 -60.445 29.295 -60.275 ;
      RECT 29.155 -59.548 29.245 -58.541 ;
      RECT 29.155 -59.235 29.295 -59.065 ;
      RECT 29.155 -57.739 29.245 -56.732 ;
      RECT 29.155 -57.215 29.295 -57.045 ;
      RECT 29.155 -56.318 29.245 -55.311 ;
      RECT 29.155 -56.005 29.295 -55.835 ;
      RECT 29.155 -54.509 29.245 -53.502 ;
      RECT 29.155 -53.985 29.295 -53.815 ;
      RECT 29.155 -53.088 29.245 -52.081 ;
      RECT 29.155 -52.775 29.295 -52.605 ;
      RECT 29.155 -51.279 29.245 -50.272 ;
      RECT 29.155 -50.755 29.295 -50.585 ;
      RECT 29.155 -49.858 29.245 -48.851 ;
      RECT 29.155 -49.545 29.295 -49.375 ;
      RECT 29.155 -48.049 29.245 -47.042 ;
      RECT 29.155 -47.525 29.295 -47.355 ;
      RECT 29.155 -46.628 29.245 -45.621 ;
      RECT 29.155 -46.315 29.295 -46.145 ;
      RECT 29.155 -44.819 29.245 -43.812 ;
      RECT 29.155 -44.295 29.295 -44.125 ;
      RECT 29.155 -43.398 29.245 -42.391 ;
      RECT 29.155 -43.085 29.295 -42.915 ;
      RECT 29.155 -41.589 29.245 -40.582 ;
      RECT 29.155 -41.065 29.295 -40.895 ;
      RECT 29.155 -40.168 29.245 -39.161 ;
      RECT 29.155 -39.855 29.295 -39.685 ;
      RECT 29.155 -38.359 29.245 -37.352 ;
      RECT 29.155 -37.835 29.295 -37.665 ;
      RECT 29.155 -36.938 29.245 -35.931 ;
      RECT 29.155 -36.625 29.295 -36.455 ;
      RECT 29.155 -35.129 29.245 -34.122 ;
      RECT 29.155 -34.605 29.295 -34.435 ;
      RECT 29.155 -33.708 29.245 -32.701 ;
      RECT 29.155 -33.395 29.295 -33.225 ;
      RECT 29.155 -31.899 29.245 -30.892 ;
      RECT 29.155 -31.375 29.295 -31.205 ;
      RECT 29.155 -30.478 29.245 -29.471 ;
      RECT 29.155 -30.165 29.295 -29.995 ;
      RECT 29.155 -28.669 29.245 -27.662 ;
      RECT 29.155 -28.145 29.295 -27.975 ;
      RECT 29.155 -27.248 29.245 -26.241 ;
      RECT 29.155 -26.935 29.295 -26.765 ;
      RECT 29.155 -25.439 29.245 -24.432 ;
      RECT 29.155 -24.915 29.295 -24.745 ;
      RECT 29.155 -24.018 29.245 -23.011 ;
      RECT 29.155 -23.705 29.295 -23.535 ;
      RECT 29.155 -22.209 29.245 -21.202 ;
      RECT 29.155 -21.685 29.295 -21.515 ;
      RECT 29.155 -20.788 29.245 -19.781 ;
      RECT 29.155 -20.475 29.295 -20.305 ;
      RECT 29.155 -18.979 29.245 -17.972 ;
      RECT 29.155 -18.455 29.295 -18.285 ;
      RECT 29.155 -17.558 29.245 -16.551 ;
      RECT 29.155 -17.245 29.295 -17.075 ;
      RECT 29.155 -15.749 29.245 -14.742 ;
      RECT 29.155 -15.225 29.295 -15.055 ;
      RECT 29.155 -14.328 29.245 -13.321 ;
      RECT 29.155 -14.015 29.295 -13.845 ;
      RECT 29.155 -12.519 29.245 -11.512 ;
      RECT 29.155 -11.995 29.295 -11.825 ;
      RECT 29.155 -11.098 29.245 -10.091 ;
      RECT 29.155 -10.785 29.295 -10.615 ;
      RECT 29.155 -9.289 29.245 -8.282 ;
      RECT 29.155 -8.765 29.295 -8.595 ;
      RECT 29.155 -7.868 29.245 -6.861 ;
      RECT 29.155 -7.555 29.295 -7.385 ;
      RECT 29.155 -6.059 29.245 -5.052 ;
      RECT 29.155 -5.535 29.295 -5.365 ;
      RECT 29.155 -4.638 29.245 -3.631 ;
      RECT 29.155 -4.325 29.295 -4.155 ;
      RECT 29.155 -2.829 29.245 -1.822 ;
      RECT 29.155 -2.305 29.295 -2.135 ;
      RECT 29.155 -1.408 29.245 -0.401 ;
      RECT 29.155 -1.095 29.295 -0.925 ;
      RECT 29.155 0.401 29.245 1.408 ;
      RECT 29.155 0.925 29.295 1.095 ;
      RECT 24.985 -108.935 28.765 -108.815 ;
      RECT 26.305 -109.475 26.405 -108.815 ;
      RECT 25.745 -109.475 25.845 -108.815 ;
      RECT 25.185 -109.475 25.285 -108.815 ;
      RECT 28.355 -101.538 28.445 -100.53 ;
      RECT 28.305 -100.935 28.445 -100.765 ;
      RECT 28.355 -99.73 28.445 -98.722 ;
      RECT 28.305 -99.495 28.445 -99.325 ;
      RECT 28.355 -98.308 28.445 -97.3 ;
      RECT 28.305 -97.705 28.445 -97.535 ;
      RECT 28.355 -96.5 28.445 -95.492 ;
      RECT 28.305 -96.265 28.445 -96.095 ;
      RECT 28.355 -95.078 28.445 -94.07 ;
      RECT 28.305 -94.475 28.445 -94.305 ;
      RECT 28.355 -93.27 28.445 -92.262 ;
      RECT 28.305 -93.035 28.445 -92.865 ;
      RECT 28.355 -91.848 28.445 -90.84 ;
      RECT 28.305 -91.245 28.445 -91.075 ;
      RECT 28.355 -90.04 28.445 -89.032 ;
      RECT 28.305 -89.805 28.445 -89.635 ;
      RECT 28.355 -88.618 28.445 -87.61 ;
      RECT 28.305 -88.015 28.445 -87.845 ;
      RECT 28.355 -86.81 28.445 -85.802 ;
      RECT 28.305 -86.575 28.445 -86.405 ;
      RECT 28.355 -85.388 28.445 -84.38 ;
      RECT 28.305 -84.785 28.445 -84.615 ;
      RECT 28.355 -83.58 28.445 -82.572 ;
      RECT 28.305 -83.345 28.445 -83.175 ;
      RECT 28.355 -82.158 28.445 -81.15 ;
      RECT 28.305 -81.555 28.445 -81.385 ;
      RECT 28.355 -80.35 28.445 -79.342 ;
      RECT 28.305 -80.115 28.445 -79.945 ;
      RECT 28.355 -78.928 28.445 -77.92 ;
      RECT 28.305 -78.325 28.445 -78.155 ;
      RECT 28.355 -77.12 28.445 -76.112 ;
      RECT 28.305 -76.885 28.445 -76.715 ;
      RECT 28.355 -75.698 28.445 -74.69 ;
      RECT 28.305 -75.095 28.445 -74.925 ;
      RECT 28.355 -73.89 28.445 -72.882 ;
      RECT 28.305 -73.655 28.445 -73.485 ;
      RECT 28.355 -72.468 28.445 -71.46 ;
      RECT 28.305 -71.865 28.445 -71.695 ;
      RECT 28.355 -70.66 28.445 -69.652 ;
      RECT 28.305 -70.425 28.445 -70.255 ;
      RECT 28.355 -69.238 28.445 -68.23 ;
      RECT 28.305 -68.635 28.445 -68.465 ;
      RECT 28.355 -67.43 28.445 -66.422 ;
      RECT 28.305 -67.195 28.445 -67.025 ;
      RECT 28.355 -66.008 28.445 -65 ;
      RECT 28.305 -65.405 28.445 -65.235 ;
      RECT 28.355 -64.2 28.445 -63.192 ;
      RECT 28.305 -63.965 28.445 -63.795 ;
      RECT 28.355 -62.778 28.445 -61.77 ;
      RECT 28.305 -62.175 28.445 -62.005 ;
      RECT 28.355 -60.97 28.445 -59.962 ;
      RECT 28.305 -60.735 28.445 -60.565 ;
      RECT 28.355 -59.548 28.445 -58.54 ;
      RECT 28.305 -58.945 28.445 -58.775 ;
      RECT 28.355 -57.74 28.445 -56.732 ;
      RECT 28.305 -57.505 28.445 -57.335 ;
      RECT 28.355 -56.318 28.445 -55.31 ;
      RECT 28.305 -55.715 28.445 -55.545 ;
      RECT 28.355 -54.51 28.445 -53.502 ;
      RECT 28.305 -54.275 28.445 -54.105 ;
      RECT 28.355 -53.088 28.445 -52.08 ;
      RECT 28.305 -52.485 28.445 -52.315 ;
      RECT 28.355 -51.28 28.445 -50.272 ;
      RECT 28.305 -51.045 28.445 -50.875 ;
      RECT 28.355 -49.858 28.445 -48.85 ;
      RECT 28.305 -49.255 28.445 -49.085 ;
      RECT 28.355 -48.05 28.445 -47.042 ;
      RECT 28.305 -47.815 28.445 -47.645 ;
      RECT 28.355 -46.628 28.445 -45.62 ;
      RECT 28.305 -46.025 28.445 -45.855 ;
      RECT 28.355 -44.82 28.445 -43.812 ;
      RECT 28.305 -44.585 28.445 -44.415 ;
      RECT 28.355 -43.398 28.445 -42.39 ;
      RECT 28.305 -42.795 28.445 -42.625 ;
      RECT 28.355 -41.59 28.445 -40.582 ;
      RECT 28.305 -41.355 28.445 -41.185 ;
      RECT 28.355 -40.168 28.445 -39.16 ;
      RECT 28.305 -39.565 28.445 -39.395 ;
      RECT 28.355 -38.36 28.445 -37.352 ;
      RECT 28.305 -38.125 28.445 -37.955 ;
      RECT 28.355 -36.938 28.445 -35.93 ;
      RECT 28.305 -36.335 28.445 -36.165 ;
      RECT 28.355 -35.13 28.445 -34.122 ;
      RECT 28.305 -34.895 28.445 -34.725 ;
      RECT 28.355 -33.708 28.445 -32.7 ;
      RECT 28.305 -33.105 28.445 -32.935 ;
      RECT 28.355 -31.9 28.445 -30.892 ;
      RECT 28.305 -31.665 28.445 -31.495 ;
      RECT 28.355 -30.478 28.445 -29.47 ;
      RECT 28.305 -29.875 28.445 -29.705 ;
      RECT 28.355 -28.67 28.445 -27.662 ;
      RECT 28.305 -28.435 28.445 -28.265 ;
      RECT 28.355 -27.248 28.445 -26.24 ;
      RECT 28.305 -26.645 28.445 -26.475 ;
      RECT 28.355 -25.44 28.445 -24.432 ;
      RECT 28.305 -25.205 28.445 -25.035 ;
      RECT 28.355 -24.018 28.445 -23.01 ;
      RECT 28.305 -23.415 28.445 -23.245 ;
      RECT 28.355 -22.21 28.445 -21.202 ;
      RECT 28.305 -21.975 28.445 -21.805 ;
      RECT 28.355 -20.788 28.445 -19.78 ;
      RECT 28.305 -20.185 28.445 -20.015 ;
      RECT 28.355 -18.98 28.445 -17.972 ;
      RECT 28.305 -18.745 28.445 -18.575 ;
      RECT 28.355 -17.558 28.445 -16.55 ;
      RECT 28.305 -16.955 28.445 -16.785 ;
      RECT 28.355 -15.75 28.445 -14.742 ;
      RECT 28.305 -15.515 28.445 -15.345 ;
      RECT 28.355 -14.328 28.445 -13.32 ;
      RECT 28.305 -13.725 28.445 -13.555 ;
      RECT 28.355 -12.52 28.445 -11.512 ;
      RECT 28.305 -12.285 28.445 -12.115 ;
      RECT 28.355 -11.098 28.445 -10.09 ;
      RECT 28.305 -10.495 28.445 -10.325 ;
      RECT 28.355 -9.29 28.445 -8.282 ;
      RECT 28.305 -9.055 28.445 -8.885 ;
      RECT 28.355 -7.868 28.445 -6.86 ;
      RECT 28.305 -7.265 28.445 -7.095 ;
      RECT 28.355 -6.06 28.445 -5.052 ;
      RECT 28.305 -5.825 28.445 -5.655 ;
      RECT 28.355 -4.638 28.445 -3.63 ;
      RECT 28.305 -4.035 28.445 -3.865 ;
      RECT 28.355 -2.83 28.445 -1.822 ;
      RECT 28.305 -2.595 28.445 -2.425 ;
      RECT 28.355 -1.408 28.445 -0.4 ;
      RECT 28.305 -0.805 28.445 -0.635 ;
      RECT 28.355 0.4 28.445 1.408 ;
      RECT 28.305 0.635 28.445 0.805 ;
      RECT 26.925 -111.685 28.405 -111.585 ;
      RECT 26.925 -112.195 27.025 -111.585 ;
      RECT 27.145 -109.15 28.405 -109.05 ;
      RECT 28.305 -109.475 28.405 -109.05 ;
      RECT 27.745 -109.475 27.845 -109.05 ;
      RECT 27.185 -109.475 27.285 -109.05 ;
      RECT 27.955 -101.538 28.045 -100.531 ;
      RECT 27.955 -101.225 28.095 -101.055 ;
      RECT 27.955 -99.729 28.045 -98.722 ;
      RECT 27.955 -99.205 28.095 -99.035 ;
      RECT 27.955 -98.308 28.045 -97.301 ;
      RECT 27.955 -97.995 28.095 -97.825 ;
      RECT 27.955 -96.499 28.045 -95.492 ;
      RECT 27.955 -95.975 28.095 -95.805 ;
      RECT 27.955 -95.078 28.045 -94.071 ;
      RECT 27.955 -94.765 28.095 -94.595 ;
      RECT 27.955 -93.269 28.045 -92.262 ;
      RECT 27.955 -92.745 28.095 -92.575 ;
      RECT 27.955 -91.848 28.045 -90.841 ;
      RECT 27.955 -91.535 28.095 -91.365 ;
      RECT 27.955 -90.039 28.045 -89.032 ;
      RECT 27.955 -89.515 28.095 -89.345 ;
      RECT 27.955 -88.618 28.045 -87.611 ;
      RECT 27.955 -88.305 28.095 -88.135 ;
      RECT 27.955 -86.809 28.045 -85.802 ;
      RECT 27.955 -86.285 28.095 -86.115 ;
      RECT 27.955 -85.388 28.045 -84.381 ;
      RECT 27.955 -85.075 28.095 -84.905 ;
      RECT 27.955 -83.579 28.045 -82.572 ;
      RECT 27.955 -83.055 28.095 -82.885 ;
      RECT 27.955 -82.158 28.045 -81.151 ;
      RECT 27.955 -81.845 28.095 -81.675 ;
      RECT 27.955 -80.349 28.045 -79.342 ;
      RECT 27.955 -79.825 28.095 -79.655 ;
      RECT 27.955 -78.928 28.045 -77.921 ;
      RECT 27.955 -78.615 28.095 -78.445 ;
      RECT 27.955 -77.119 28.045 -76.112 ;
      RECT 27.955 -76.595 28.095 -76.425 ;
      RECT 27.955 -75.698 28.045 -74.691 ;
      RECT 27.955 -75.385 28.095 -75.215 ;
      RECT 27.955 -73.889 28.045 -72.882 ;
      RECT 27.955 -73.365 28.095 -73.195 ;
      RECT 27.955 -72.468 28.045 -71.461 ;
      RECT 27.955 -72.155 28.095 -71.985 ;
      RECT 27.955 -70.659 28.045 -69.652 ;
      RECT 27.955 -70.135 28.095 -69.965 ;
      RECT 27.955 -69.238 28.045 -68.231 ;
      RECT 27.955 -68.925 28.095 -68.755 ;
      RECT 27.955 -67.429 28.045 -66.422 ;
      RECT 27.955 -66.905 28.095 -66.735 ;
      RECT 27.955 -66.008 28.045 -65.001 ;
      RECT 27.955 -65.695 28.095 -65.525 ;
      RECT 27.955 -64.199 28.045 -63.192 ;
      RECT 27.955 -63.675 28.095 -63.505 ;
      RECT 27.955 -62.778 28.045 -61.771 ;
      RECT 27.955 -62.465 28.095 -62.295 ;
      RECT 27.955 -60.969 28.045 -59.962 ;
      RECT 27.955 -60.445 28.095 -60.275 ;
      RECT 27.955 -59.548 28.045 -58.541 ;
      RECT 27.955 -59.235 28.095 -59.065 ;
      RECT 27.955 -57.739 28.045 -56.732 ;
      RECT 27.955 -57.215 28.095 -57.045 ;
      RECT 27.955 -56.318 28.045 -55.311 ;
      RECT 27.955 -56.005 28.095 -55.835 ;
      RECT 27.955 -54.509 28.045 -53.502 ;
      RECT 27.955 -53.985 28.095 -53.815 ;
      RECT 27.955 -53.088 28.045 -52.081 ;
      RECT 27.955 -52.775 28.095 -52.605 ;
      RECT 27.955 -51.279 28.045 -50.272 ;
      RECT 27.955 -50.755 28.095 -50.585 ;
      RECT 27.955 -49.858 28.045 -48.851 ;
      RECT 27.955 -49.545 28.095 -49.375 ;
      RECT 27.955 -48.049 28.045 -47.042 ;
      RECT 27.955 -47.525 28.095 -47.355 ;
      RECT 27.955 -46.628 28.045 -45.621 ;
      RECT 27.955 -46.315 28.095 -46.145 ;
      RECT 27.955 -44.819 28.045 -43.812 ;
      RECT 27.955 -44.295 28.095 -44.125 ;
      RECT 27.955 -43.398 28.045 -42.391 ;
      RECT 27.955 -43.085 28.095 -42.915 ;
      RECT 27.955 -41.589 28.045 -40.582 ;
      RECT 27.955 -41.065 28.095 -40.895 ;
      RECT 27.955 -40.168 28.045 -39.161 ;
      RECT 27.955 -39.855 28.095 -39.685 ;
      RECT 27.955 -38.359 28.045 -37.352 ;
      RECT 27.955 -37.835 28.095 -37.665 ;
      RECT 27.955 -36.938 28.045 -35.931 ;
      RECT 27.955 -36.625 28.095 -36.455 ;
      RECT 27.955 -35.129 28.045 -34.122 ;
      RECT 27.955 -34.605 28.095 -34.435 ;
      RECT 27.955 -33.708 28.045 -32.701 ;
      RECT 27.955 -33.395 28.095 -33.225 ;
      RECT 27.955 -31.899 28.045 -30.892 ;
      RECT 27.955 -31.375 28.095 -31.205 ;
      RECT 27.955 -30.478 28.045 -29.471 ;
      RECT 27.955 -30.165 28.095 -29.995 ;
      RECT 27.955 -28.669 28.045 -27.662 ;
      RECT 27.955 -28.145 28.095 -27.975 ;
      RECT 27.955 -27.248 28.045 -26.241 ;
      RECT 27.955 -26.935 28.095 -26.765 ;
      RECT 27.955 -25.439 28.045 -24.432 ;
      RECT 27.955 -24.915 28.095 -24.745 ;
      RECT 27.955 -24.018 28.045 -23.011 ;
      RECT 27.955 -23.705 28.095 -23.535 ;
      RECT 27.955 -22.209 28.045 -21.202 ;
      RECT 27.955 -21.685 28.095 -21.515 ;
      RECT 27.955 -20.788 28.045 -19.781 ;
      RECT 27.955 -20.475 28.095 -20.305 ;
      RECT 27.955 -18.979 28.045 -17.972 ;
      RECT 27.955 -18.455 28.095 -18.285 ;
      RECT 27.955 -17.558 28.045 -16.551 ;
      RECT 27.955 -17.245 28.095 -17.075 ;
      RECT 27.955 -15.749 28.045 -14.742 ;
      RECT 27.955 -15.225 28.095 -15.055 ;
      RECT 27.955 -14.328 28.045 -13.321 ;
      RECT 27.955 -14.015 28.095 -13.845 ;
      RECT 27.955 -12.519 28.045 -11.512 ;
      RECT 27.955 -11.995 28.095 -11.825 ;
      RECT 27.955 -11.098 28.045 -10.091 ;
      RECT 27.955 -10.785 28.095 -10.615 ;
      RECT 27.955 -9.289 28.045 -8.282 ;
      RECT 27.955 -8.765 28.095 -8.595 ;
      RECT 27.955 -7.868 28.045 -6.861 ;
      RECT 27.955 -7.555 28.095 -7.385 ;
      RECT 27.955 -6.059 28.045 -5.052 ;
      RECT 27.955 -5.535 28.095 -5.365 ;
      RECT 27.955 -4.638 28.045 -3.631 ;
      RECT 27.955 -4.325 28.095 -4.155 ;
      RECT 27.955 -2.829 28.045 -1.822 ;
      RECT 27.955 -2.305 28.095 -2.135 ;
      RECT 27.955 -1.408 28.045 -0.401 ;
      RECT 27.955 -1.095 28.095 -0.925 ;
      RECT 27.955 0.401 28.045 1.408 ;
      RECT 27.955 0.925 28.095 1.095 ;
      RECT 27.285 -111.495 27.455 -111.385 ;
      RECT 24.135 -111.495 27.455 -111.395 ;
      RECT 27.155 -101.538 27.245 -100.53 ;
      RECT 27.105 -100.935 27.245 -100.765 ;
      RECT 27.155 -99.73 27.245 -98.722 ;
      RECT 27.105 -99.495 27.245 -99.325 ;
      RECT 27.155 -98.308 27.245 -97.3 ;
      RECT 27.105 -97.705 27.245 -97.535 ;
      RECT 27.155 -96.5 27.245 -95.492 ;
      RECT 27.105 -96.265 27.245 -96.095 ;
      RECT 27.155 -95.078 27.245 -94.07 ;
      RECT 27.105 -94.475 27.245 -94.305 ;
      RECT 27.155 -93.27 27.245 -92.262 ;
      RECT 27.105 -93.035 27.245 -92.865 ;
      RECT 27.155 -91.848 27.245 -90.84 ;
      RECT 27.105 -91.245 27.245 -91.075 ;
      RECT 27.155 -90.04 27.245 -89.032 ;
      RECT 27.105 -89.805 27.245 -89.635 ;
      RECT 27.155 -88.618 27.245 -87.61 ;
      RECT 27.105 -88.015 27.245 -87.845 ;
      RECT 27.155 -86.81 27.245 -85.802 ;
      RECT 27.105 -86.575 27.245 -86.405 ;
      RECT 27.155 -85.388 27.245 -84.38 ;
      RECT 27.105 -84.785 27.245 -84.615 ;
      RECT 27.155 -83.58 27.245 -82.572 ;
      RECT 27.105 -83.345 27.245 -83.175 ;
      RECT 27.155 -82.158 27.245 -81.15 ;
      RECT 27.105 -81.555 27.245 -81.385 ;
      RECT 27.155 -80.35 27.245 -79.342 ;
      RECT 27.105 -80.115 27.245 -79.945 ;
      RECT 27.155 -78.928 27.245 -77.92 ;
      RECT 27.105 -78.325 27.245 -78.155 ;
      RECT 27.155 -77.12 27.245 -76.112 ;
      RECT 27.105 -76.885 27.245 -76.715 ;
      RECT 27.155 -75.698 27.245 -74.69 ;
      RECT 27.105 -75.095 27.245 -74.925 ;
      RECT 27.155 -73.89 27.245 -72.882 ;
      RECT 27.105 -73.655 27.245 -73.485 ;
      RECT 27.155 -72.468 27.245 -71.46 ;
      RECT 27.105 -71.865 27.245 -71.695 ;
      RECT 27.155 -70.66 27.245 -69.652 ;
      RECT 27.105 -70.425 27.245 -70.255 ;
      RECT 27.155 -69.238 27.245 -68.23 ;
      RECT 27.105 -68.635 27.245 -68.465 ;
      RECT 27.155 -67.43 27.245 -66.422 ;
      RECT 27.105 -67.195 27.245 -67.025 ;
      RECT 27.155 -66.008 27.245 -65 ;
      RECT 27.105 -65.405 27.245 -65.235 ;
      RECT 27.155 -64.2 27.245 -63.192 ;
      RECT 27.105 -63.965 27.245 -63.795 ;
      RECT 27.155 -62.778 27.245 -61.77 ;
      RECT 27.105 -62.175 27.245 -62.005 ;
      RECT 27.155 -60.97 27.245 -59.962 ;
      RECT 27.105 -60.735 27.245 -60.565 ;
      RECT 27.155 -59.548 27.245 -58.54 ;
      RECT 27.105 -58.945 27.245 -58.775 ;
      RECT 27.155 -57.74 27.245 -56.732 ;
      RECT 27.105 -57.505 27.245 -57.335 ;
      RECT 27.155 -56.318 27.245 -55.31 ;
      RECT 27.105 -55.715 27.245 -55.545 ;
      RECT 27.155 -54.51 27.245 -53.502 ;
      RECT 27.105 -54.275 27.245 -54.105 ;
      RECT 27.155 -53.088 27.245 -52.08 ;
      RECT 27.105 -52.485 27.245 -52.315 ;
      RECT 27.155 -51.28 27.245 -50.272 ;
      RECT 27.105 -51.045 27.245 -50.875 ;
      RECT 27.155 -49.858 27.245 -48.85 ;
      RECT 27.105 -49.255 27.245 -49.085 ;
      RECT 27.155 -48.05 27.245 -47.042 ;
      RECT 27.105 -47.815 27.245 -47.645 ;
      RECT 27.155 -46.628 27.245 -45.62 ;
      RECT 27.105 -46.025 27.245 -45.855 ;
      RECT 27.155 -44.82 27.245 -43.812 ;
      RECT 27.105 -44.585 27.245 -44.415 ;
      RECT 27.155 -43.398 27.245 -42.39 ;
      RECT 27.105 -42.795 27.245 -42.625 ;
      RECT 27.155 -41.59 27.245 -40.582 ;
      RECT 27.105 -41.355 27.245 -41.185 ;
      RECT 27.155 -40.168 27.245 -39.16 ;
      RECT 27.105 -39.565 27.245 -39.395 ;
      RECT 27.155 -38.36 27.245 -37.352 ;
      RECT 27.105 -38.125 27.245 -37.955 ;
      RECT 27.155 -36.938 27.245 -35.93 ;
      RECT 27.105 -36.335 27.245 -36.165 ;
      RECT 27.155 -35.13 27.245 -34.122 ;
      RECT 27.105 -34.895 27.245 -34.725 ;
      RECT 27.155 -33.708 27.245 -32.7 ;
      RECT 27.105 -33.105 27.245 -32.935 ;
      RECT 27.155 -31.9 27.245 -30.892 ;
      RECT 27.105 -31.665 27.245 -31.495 ;
      RECT 27.155 -30.478 27.245 -29.47 ;
      RECT 27.105 -29.875 27.245 -29.705 ;
      RECT 27.155 -28.67 27.245 -27.662 ;
      RECT 27.105 -28.435 27.245 -28.265 ;
      RECT 27.155 -27.248 27.245 -26.24 ;
      RECT 27.105 -26.645 27.245 -26.475 ;
      RECT 27.155 -25.44 27.245 -24.432 ;
      RECT 27.105 -25.205 27.245 -25.035 ;
      RECT 27.155 -24.018 27.245 -23.01 ;
      RECT 27.105 -23.415 27.245 -23.245 ;
      RECT 27.155 -22.21 27.245 -21.202 ;
      RECT 27.105 -21.975 27.245 -21.805 ;
      RECT 27.155 -20.788 27.245 -19.78 ;
      RECT 27.105 -20.185 27.245 -20.015 ;
      RECT 27.155 -18.98 27.245 -17.972 ;
      RECT 27.105 -18.745 27.245 -18.575 ;
      RECT 27.155 -17.558 27.245 -16.55 ;
      RECT 27.105 -16.955 27.245 -16.785 ;
      RECT 27.155 -15.75 27.245 -14.742 ;
      RECT 27.105 -15.515 27.245 -15.345 ;
      RECT 27.155 -14.328 27.245 -13.32 ;
      RECT 27.105 -13.725 27.245 -13.555 ;
      RECT 27.155 -12.52 27.245 -11.512 ;
      RECT 27.105 -12.285 27.245 -12.115 ;
      RECT 27.155 -11.098 27.245 -10.09 ;
      RECT 27.105 -10.495 27.245 -10.325 ;
      RECT 27.155 -9.29 27.245 -8.282 ;
      RECT 27.105 -9.055 27.245 -8.885 ;
      RECT 27.155 -7.868 27.245 -6.86 ;
      RECT 27.105 -7.265 27.245 -7.095 ;
      RECT 27.155 -6.06 27.245 -5.052 ;
      RECT 27.105 -5.825 27.245 -5.655 ;
      RECT 27.155 -4.638 27.245 -3.63 ;
      RECT 27.105 -4.035 27.245 -3.865 ;
      RECT 27.155 -2.83 27.245 -1.822 ;
      RECT 27.105 -2.595 27.245 -2.425 ;
      RECT 27.155 -1.408 27.245 -0.4 ;
      RECT 27.105 -0.805 27.245 -0.635 ;
      RECT 27.155 0.4 27.245 1.408 ;
      RECT 27.105 0.635 27.245 0.805 ;
      RECT 26.755 -101.538 26.845 -100.531 ;
      RECT 26.755 -101.225 26.895 -101.055 ;
      RECT 26.755 -99.729 26.845 -98.722 ;
      RECT 26.755 -99.205 26.895 -99.035 ;
      RECT 26.755 -98.308 26.845 -97.301 ;
      RECT 26.755 -97.995 26.895 -97.825 ;
      RECT 26.755 -96.499 26.845 -95.492 ;
      RECT 26.755 -95.975 26.895 -95.805 ;
      RECT 26.755 -95.078 26.845 -94.071 ;
      RECT 26.755 -94.765 26.895 -94.595 ;
      RECT 26.755 -93.269 26.845 -92.262 ;
      RECT 26.755 -92.745 26.895 -92.575 ;
      RECT 26.755 -91.848 26.845 -90.841 ;
      RECT 26.755 -91.535 26.895 -91.365 ;
      RECT 26.755 -90.039 26.845 -89.032 ;
      RECT 26.755 -89.515 26.895 -89.345 ;
      RECT 26.755 -88.618 26.845 -87.611 ;
      RECT 26.755 -88.305 26.895 -88.135 ;
      RECT 26.755 -86.809 26.845 -85.802 ;
      RECT 26.755 -86.285 26.895 -86.115 ;
      RECT 26.755 -85.388 26.845 -84.381 ;
      RECT 26.755 -85.075 26.895 -84.905 ;
      RECT 26.755 -83.579 26.845 -82.572 ;
      RECT 26.755 -83.055 26.895 -82.885 ;
      RECT 26.755 -82.158 26.845 -81.151 ;
      RECT 26.755 -81.845 26.895 -81.675 ;
      RECT 26.755 -80.349 26.845 -79.342 ;
      RECT 26.755 -79.825 26.895 -79.655 ;
      RECT 26.755 -78.928 26.845 -77.921 ;
      RECT 26.755 -78.615 26.895 -78.445 ;
      RECT 26.755 -77.119 26.845 -76.112 ;
      RECT 26.755 -76.595 26.895 -76.425 ;
      RECT 26.755 -75.698 26.845 -74.691 ;
      RECT 26.755 -75.385 26.895 -75.215 ;
      RECT 26.755 -73.889 26.845 -72.882 ;
      RECT 26.755 -73.365 26.895 -73.195 ;
      RECT 26.755 -72.468 26.845 -71.461 ;
      RECT 26.755 -72.155 26.895 -71.985 ;
      RECT 26.755 -70.659 26.845 -69.652 ;
      RECT 26.755 -70.135 26.895 -69.965 ;
      RECT 26.755 -69.238 26.845 -68.231 ;
      RECT 26.755 -68.925 26.895 -68.755 ;
      RECT 26.755 -67.429 26.845 -66.422 ;
      RECT 26.755 -66.905 26.895 -66.735 ;
      RECT 26.755 -66.008 26.845 -65.001 ;
      RECT 26.755 -65.695 26.895 -65.525 ;
      RECT 26.755 -64.199 26.845 -63.192 ;
      RECT 26.755 -63.675 26.895 -63.505 ;
      RECT 26.755 -62.778 26.845 -61.771 ;
      RECT 26.755 -62.465 26.895 -62.295 ;
      RECT 26.755 -60.969 26.845 -59.962 ;
      RECT 26.755 -60.445 26.895 -60.275 ;
      RECT 26.755 -59.548 26.845 -58.541 ;
      RECT 26.755 -59.235 26.895 -59.065 ;
      RECT 26.755 -57.739 26.845 -56.732 ;
      RECT 26.755 -57.215 26.895 -57.045 ;
      RECT 26.755 -56.318 26.845 -55.311 ;
      RECT 26.755 -56.005 26.895 -55.835 ;
      RECT 26.755 -54.509 26.845 -53.502 ;
      RECT 26.755 -53.985 26.895 -53.815 ;
      RECT 26.755 -53.088 26.845 -52.081 ;
      RECT 26.755 -52.775 26.895 -52.605 ;
      RECT 26.755 -51.279 26.845 -50.272 ;
      RECT 26.755 -50.755 26.895 -50.585 ;
      RECT 26.755 -49.858 26.845 -48.851 ;
      RECT 26.755 -49.545 26.895 -49.375 ;
      RECT 26.755 -48.049 26.845 -47.042 ;
      RECT 26.755 -47.525 26.895 -47.355 ;
      RECT 26.755 -46.628 26.845 -45.621 ;
      RECT 26.755 -46.315 26.895 -46.145 ;
      RECT 26.755 -44.819 26.845 -43.812 ;
      RECT 26.755 -44.295 26.895 -44.125 ;
      RECT 26.755 -43.398 26.845 -42.391 ;
      RECT 26.755 -43.085 26.895 -42.915 ;
      RECT 26.755 -41.589 26.845 -40.582 ;
      RECT 26.755 -41.065 26.895 -40.895 ;
      RECT 26.755 -40.168 26.845 -39.161 ;
      RECT 26.755 -39.855 26.895 -39.685 ;
      RECT 26.755 -38.359 26.845 -37.352 ;
      RECT 26.755 -37.835 26.895 -37.665 ;
      RECT 26.755 -36.938 26.845 -35.931 ;
      RECT 26.755 -36.625 26.895 -36.455 ;
      RECT 26.755 -35.129 26.845 -34.122 ;
      RECT 26.755 -34.605 26.895 -34.435 ;
      RECT 26.755 -33.708 26.845 -32.701 ;
      RECT 26.755 -33.395 26.895 -33.225 ;
      RECT 26.755 -31.899 26.845 -30.892 ;
      RECT 26.755 -31.375 26.895 -31.205 ;
      RECT 26.755 -30.478 26.845 -29.471 ;
      RECT 26.755 -30.165 26.895 -29.995 ;
      RECT 26.755 -28.669 26.845 -27.662 ;
      RECT 26.755 -28.145 26.895 -27.975 ;
      RECT 26.755 -27.248 26.845 -26.241 ;
      RECT 26.755 -26.935 26.895 -26.765 ;
      RECT 26.755 -25.439 26.845 -24.432 ;
      RECT 26.755 -24.915 26.895 -24.745 ;
      RECT 26.755 -24.018 26.845 -23.011 ;
      RECT 26.755 -23.705 26.895 -23.535 ;
      RECT 26.755 -22.209 26.845 -21.202 ;
      RECT 26.755 -21.685 26.895 -21.515 ;
      RECT 26.755 -20.788 26.845 -19.781 ;
      RECT 26.755 -20.475 26.895 -20.305 ;
      RECT 26.755 -18.979 26.845 -17.972 ;
      RECT 26.755 -18.455 26.895 -18.285 ;
      RECT 26.755 -17.558 26.845 -16.551 ;
      RECT 26.755 -17.245 26.895 -17.075 ;
      RECT 26.755 -15.749 26.845 -14.742 ;
      RECT 26.755 -15.225 26.895 -15.055 ;
      RECT 26.755 -14.328 26.845 -13.321 ;
      RECT 26.755 -14.015 26.895 -13.845 ;
      RECT 26.755 -12.519 26.845 -11.512 ;
      RECT 26.755 -11.995 26.895 -11.825 ;
      RECT 26.755 -11.098 26.845 -10.091 ;
      RECT 26.755 -10.785 26.895 -10.615 ;
      RECT 26.755 -9.289 26.845 -8.282 ;
      RECT 26.755 -8.765 26.895 -8.595 ;
      RECT 26.755 -7.868 26.845 -6.861 ;
      RECT 26.755 -7.555 26.895 -7.385 ;
      RECT 26.755 -6.059 26.845 -5.052 ;
      RECT 26.755 -5.535 26.895 -5.365 ;
      RECT 26.755 -4.638 26.845 -3.631 ;
      RECT 26.755 -4.325 26.895 -4.155 ;
      RECT 26.755 -2.829 26.845 -1.822 ;
      RECT 26.755 -2.305 26.895 -2.135 ;
      RECT 26.755 -1.408 26.845 -0.401 ;
      RECT 26.755 -1.095 26.895 -0.925 ;
      RECT 26.755 0.401 26.845 1.408 ;
      RECT 26.755 0.925 26.895 1.095 ;
      RECT 24.905 -111.685 26.385 -111.585 ;
      RECT 24.905 -112.055 25.005 -111.585 ;
      RECT 24.71 -114.395 26.285 -114.275 ;
      RECT 26.185 -114.895 26.285 -114.275 ;
      RECT 25.59 -114.895 25.69 -114.275 ;
      RECT 24.71 -114.85 24.81 -114.275 ;
      RECT 25.955 -101.538 26.045 -100.53 ;
      RECT 25.905 -100.935 26.045 -100.765 ;
      RECT 25.955 -99.73 26.045 -98.722 ;
      RECT 25.905 -99.495 26.045 -99.325 ;
      RECT 25.955 -98.308 26.045 -97.3 ;
      RECT 25.905 -97.705 26.045 -97.535 ;
      RECT 25.955 -96.5 26.045 -95.492 ;
      RECT 25.905 -96.265 26.045 -96.095 ;
      RECT 25.955 -95.078 26.045 -94.07 ;
      RECT 25.905 -94.475 26.045 -94.305 ;
      RECT 25.955 -93.27 26.045 -92.262 ;
      RECT 25.905 -93.035 26.045 -92.865 ;
      RECT 25.955 -91.848 26.045 -90.84 ;
      RECT 25.905 -91.245 26.045 -91.075 ;
      RECT 25.955 -90.04 26.045 -89.032 ;
      RECT 25.905 -89.805 26.045 -89.635 ;
      RECT 25.955 -88.618 26.045 -87.61 ;
      RECT 25.905 -88.015 26.045 -87.845 ;
      RECT 25.955 -86.81 26.045 -85.802 ;
      RECT 25.905 -86.575 26.045 -86.405 ;
      RECT 25.955 -85.388 26.045 -84.38 ;
      RECT 25.905 -84.785 26.045 -84.615 ;
      RECT 25.955 -83.58 26.045 -82.572 ;
      RECT 25.905 -83.345 26.045 -83.175 ;
      RECT 25.955 -82.158 26.045 -81.15 ;
      RECT 25.905 -81.555 26.045 -81.385 ;
      RECT 25.955 -80.35 26.045 -79.342 ;
      RECT 25.905 -80.115 26.045 -79.945 ;
      RECT 25.955 -78.928 26.045 -77.92 ;
      RECT 25.905 -78.325 26.045 -78.155 ;
      RECT 25.955 -77.12 26.045 -76.112 ;
      RECT 25.905 -76.885 26.045 -76.715 ;
      RECT 25.955 -75.698 26.045 -74.69 ;
      RECT 25.905 -75.095 26.045 -74.925 ;
      RECT 25.955 -73.89 26.045 -72.882 ;
      RECT 25.905 -73.655 26.045 -73.485 ;
      RECT 25.955 -72.468 26.045 -71.46 ;
      RECT 25.905 -71.865 26.045 -71.695 ;
      RECT 25.955 -70.66 26.045 -69.652 ;
      RECT 25.905 -70.425 26.045 -70.255 ;
      RECT 25.955 -69.238 26.045 -68.23 ;
      RECT 25.905 -68.635 26.045 -68.465 ;
      RECT 25.955 -67.43 26.045 -66.422 ;
      RECT 25.905 -67.195 26.045 -67.025 ;
      RECT 25.955 -66.008 26.045 -65 ;
      RECT 25.905 -65.405 26.045 -65.235 ;
      RECT 25.955 -64.2 26.045 -63.192 ;
      RECT 25.905 -63.965 26.045 -63.795 ;
      RECT 25.955 -62.778 26.045 -61.77 ;
      RECT 25.905 -62.175 26.045 -62.005 ;
      RECT 25.955 -60.97 26.045 -59.962 ;
      RECT 25.905 -60.735 26.045 -60.565 ;
      RECT 25.955 -59.548 26.045 -58.54 ;
      RECT 25.905 -58.945 26.045 -58.775 ;
      RECT 25.955 -57.74 26.045 -56.732 ;
      RECT 25.905 -57.505 26.045 -57.335 ;
      RECT 25.955 -56.318 26.045 -55.31 ;
      RECT 25.905 -55.715 26.045 -55.545 ;
      RECT 25.955 -54.51 26.045 -53.502 ;
      RECT 25.905 -54.275 26.045 -54.105 ;
      RECT 25.955 -53.088 26.045 -52.08 ;
      RECT 25.905 -52.485 26.045 -52.315 ;
      RECT 25.955 -51.28 26.045 -50.272 ;
      RECT 25.905 -51.045 26.045 -50.875 ;
      RECT 25.955 -49.858 26.045 -48.85 ;
      RECT 25.905 -49.255 26.045 -49.085 ;
      RECT 25.955 -48.05 26.045 -47.042 ;
      RECT 25.905 -47.815 26.045 -47.645 ;
      RECT 25.955 -46.628 26.045 -45.62 ;
      RECT 25.905 -46.025 26.045 -45.855 ;
      RECT 25.955 -44.82 26.045 -43.812 ;
      RECT 25.905 -44.585 26.045 -44.415 ;
      RECT 25.955 -43.398 26.045 -42.39 ;
      RECT 25.905 -42.795 26.045 -42.625 ;
      RECT 25.955 -41.59 26.045 -40.582 ;
      RECT 25.905 -41.355 26.045 -41.185 ;
      RECT 25.955 -40.168 26.045 -39.16 ;
      RECT 25.905 -39.565 26.045 -39.395 ;
      RECT 25.955 -38.36 26.045 -37.352 ;
      RECT 25.905 -38.125 26.045 -37.955 ;
      RECT 25.955 -36.938 26.045 -35.93 ;
      RECT 25.905 -36.335 26.045 -36.165 ;
      RECT 25.955 -35.13 26.045 -34.122 ;
      RECT 25.905 -34.895 26.045 -34.725 ;
      RECT 25.955 -33.708 26.045 -32.7 ;
      RECT 25.905 -33.105 26.045 -32.935 ;
      RECT 25.955 -31.9 26.045 -30.892 ;
      RECT 25.905 -31.665 26.045 -31.495 ;
      RECT 25.955 -30.478 26.045 -29.47 ;
      RECT 25.905 -29.875 26.045 -29.705 ;
      RECT 25.955 -28.67 26.045 -27.662 ;
      RECT 25.905 -28.435 26.045 -28.265 ;
      RECT 25.955 -27.248 26.045 -26.24 ;
      RECT 25.905 -26.645 26.045 -26.475 ;
      RECT 25.955 -25.44 26.045 -24.432 ;
      RECT 25.905 -25.205 26.045 -25.035 ;
      RECT 25.955 -24.018 26.045 -23.01 ;
      RECT 25.905 -23.415 26.045 -23.245 ;
      RECT 25.955 -22.21 26.045 -21.202 ;
      RECT 25.905 -21.975 26.045 -21.805 ;
      RECT 25.955 -20.788 26.045 -19.78 ;
      RECT 25.905 -20.185 26.045 -20.015 ;
      RECT 25.955 -18.98 26.045 -17.972 ;
      RECT 25.905 -18.745 26.045 -18.575 ;
      RECT 25.955 -17.558 26.045 -16.55 ;
      RECT 25.905 -16.955 26.045 -16.785 ;
      RECT 25.955 -15.75 26.045 -14.742 ;
      RECT 25.905 -15.515 26.045 -15.345 ;
      RECT 25.955 -14.328 26.045 -13.32 ;
      RECT 25.905 -13.725 26.045 -13.555 ;
      RECT 25.955 -12.52 26.045 -11.512 ;
      RECT 25.905 -12.285 26.045 -12.115 ;
      RECT 25.955 -11.098 26.045 -10.09 ;
      RECT 25.905 -10.495 26.045 -10.325 ;
      RECT 25.955 -9.29 26.045 -8.282 ;
      RECT 25.905 -9.055 26.045 -8.885 ;
      RECT 25.955 -7.868 26.045 -6.86 ;
      RECT 25.905 -7.265 26.045 -7.095 ;
      RECT 25.955 -6.06 26.045 -5.052 ;
      RECT 25.905 -5.825 26.045 -5.655 ;
      RECT 25.955 -4.638 26.045 -3.63 ;
      RECT 25.905 -4.035 26.045 -3.865 ;
      RECT 25.955 -2.83 26.045 -1.822 ;
      RECT 25.905 -2.595 26.045 -2.425 ;
      RECT 25.955 -1.408 26.045 -0.4 ;
      RECT 25.905 -0.805 26.045 -0.635 ;
      RECT 25.955 0.4 26.045 1.408 ;
      RECT 25.905 0.635 26.045 0.805 ;
      RECT 25.83 -114.685 26.005 -114.515 ;
      RECT 25.905 -114.895 26.005 -114.515 ;
      RECT 24.945 -113.555 25.045 -113.09 ;
      RECT 25.31 -113.555 25.41 -113.1 ;
      RECT 24.945 -113.555 25.79 -113.385 ;
      RECT 25.555 -101.538 25.645 -100.531 ;
      RECT 25.555 -101.225 25.695 -101.055 ;
      RECT 25.555 -99.729 25.645 -98.722 ;
      RECT 25.555 -99.205 25.695 -99.035 ;
      RECT 25.555 -98.308 25.645 -97.301 ;
      RECT 25.555 -97.995 25.695 -97.825 ;
      RECT 25.555 -96.499 25.645 -95.492 ;
      RECT 25.555 -95.975 25.695 -95.805 ;
      RECT 25.555 -95.078 25.645 -94.071 ;
      RECT 25.555 -94.765 25.695 -94.595 ;
      RECT 25.555 -93.269 25.645 -92.262 ;
      RECT 25.555 -92.745 25.695 -92.575 ;
      RECT 25.555 -91.848 25.645 -90.841 ;
      RECT 25.555 -91.535 25.695 -91.365 ;
      RECT 25.555 -90.039 25.645 -89.032 ;
      RECT 25.555 -89.515 25.695 -89.345 ;
      RECT 25.555 -88.618 25.645 -87.611 ;
      RECT 25.555 -88.305 25.695 -88.135 ;
      RECT 25.555 -86.809 25.645 -85.802 ;
      RECT 25.555 -86.285 25.695 -86.115 ;
      RECT 25.555 -85.388 25.645 -84.381 ;
      RECT 25.555 -85.075 25.695 -84.905 ;
      RECT 25.555 -83.579 25.645 -82.572 ;
      RECT 25.555 -83.055 25.695 -82.885 ;
      RECT 25.555 -82.158 25.645 -81.151 ;
      RECT 25.555 -81.845 25.695 -81.675 ;
      RECT 25.555 -80.349 25.645 -79.342 ;
      RECT 25.555 -79.825 25.695 -79.655 ;
      RECT 25.555 -78.928 25.645 -77.921 ;
      RECT 25.555 -78.615 25.695 -78.445 ;
      RECT 25.555 -77.119 25.645 -76.112 ;
      RECT 25.555 -76.595 25.695 -76.425 ;
      RECT 25.555 -75.698 25.645 -74.691 ;
      RECT 25.555 -75.385 25.695 -75.215 ;
      RECT 25.555 -73.889 25.645 -72.882 ;
      RECT 25.555 -73.365 25.695 -73.195 ;
      RECT 25.555 -72.468 25.645 -71.461 ;
      RECT 25.555 -72.155 25.695 -71.985 ;
      RECT 25.555 -70.659 25.645 -69.652 ;
      RECT 25.555 -70.135 25.695 -69.965 ;
      RECT 25.555 -69.238 25.645 -68.231 ;
      RECT 25.555 -68.925 25.695 -68.755 ;
      RECT 25.555 -67.429 25.645 -66.422 ;
      RECT 25.555 -66.905 25.695 -66.735 ;
      RECT 25.555 -66.008 25.645 -65.001 ;
      RECT 25.555 -65.695 25.695 -65.525 ;
      RECT 25.555 -64.199 25.645 -63.192 ;
      RECT 25.555 -63.675 25.695 -63.505 ;
      RECT 25.555 -62.778 25.645 -61.771 ;
      RECT 25.555 -62.465 25.695 -62.295 ;
      RECT 25.555 -60.969 25.645 -59.962 ;
      RECT 25.555 -60.445 25.695 -60.275 ;
      RECT 25.555 -59.548 25.645 -58.541 ;
      RECT 25.555 -59.235 25.695 -59.065 ;
      RECT 25.555 -57.739 25.645 -56.732 ;
      RECT 25.555 -57.215 25.695 -57.045 ;
      RECT 25.555 -56.318 25.645 -55.311 ;
      RECT 25.555 -56.005 25.695 -55.835 ;
      RECT 25.555 -54.509 25.645 -53.502 ;
      RECT 25.555 -53.985 25.695 -53.815 ;
      RECT 25.555 -53.088 25.645 -52.081 ;
      RECT 25.555 -52.775 25.695 -52.605 ;
      RECT 25.555 -51.279 25.645 -50.272 ;
      RECT 25.555 -50.755 25.695 -50.585 ;
      RECT 25.555 -49.858 25.645 -48.851 ;
      RECT 25.555 -49.545 25.695 -49.375 ;
      RECT 25.555 -48.049 25.645 -47.042 ;
      RECT 25.555 -47.525 25.695 -47.355 ;
      RECT 25.555 -46.628 25.645 -45.621 ;
      RECT 25.555 -46.315 25.695 -46.145 ;
      RECT 25.555 -44.819 25.645 -43.812 ;
      RECT 25.555 -44.295 25.695 -44.125 ;
      RECT 25.555 -43.398 25.645 -42.391 ;
      RECT 25.555 -43.085 25.695 -42.915 ;
      RECT 25.555 -41.589 25.645 -40.582 ;
      RECT 25.555 -41.065 25.695 -40.895 ;
      RECT 25.555 -40.168 25.645 -39.161 ;
      RECT 25.555 -39.855 25.695 -39.685 ;
      RECT 25.555 -38.359 25.645 -37.352 ;
      RECT 25.555 -37.835 25.695 -37.665 ;
      RECT 25.555 -36.938 25.645 -35.931 ;
      RECT 25.555 -36.625 25.695 -36.455 ;
      RECT 25.555 -35.129 25.645 -34.122 ;
      RECT 25.555 -34.605 25.695 -34.435 ;
      RECT 25.555 -33.708 25.645 -32.701 ;
      RECT 25.555 -33.395 25.695 -33.225 ;
      RECT 25.555 -31.899 25.645 -30.892 ;
      RECT 25.555 -31.375 25.695 -31.205 ;
      RECT 25.555 -30.478 25.645 -29.471 ;
      RECT 25.555 -30.165 25.695 -29.995 ;
      RECT 25.555 -28.669 25.645 -27.662 ;
      RECT 25.555 -28.145 25.695 -27.975 ;
      RECT 25.555 -27.248 25.645 -26.241 ;
      RECT 25.555 -26.935 25.695 -26.765 ;
      RECT 25.555 -25.439 25.645 -24.432 ;
      RECT 25.555 -24.915 25.695 -24.745 ;
      RECT 25.555 -24.018 25.645 -23.011 ;
      RECT 25.555 -23.705 25.695 -23.535 ;
      RECT 25.555 -22.209 25.645 -21.202 ;
      RECT 25.555 -21.685 25.695 -21.515 ;
      RECT 25.555 -20.788 25.645 -19.781 ;
      RECT 25.555 -20.475 25.695 -20.305 ;
      RECT 25.555 -18.979 25.645 -17.972 ;
      RECT 25.555 -18.455 25.695 -18.285 ;
      RECT 25.555 -17.558 25.645 -16.551 ;
      RECT 25.555 -17.245 25.695 -17.075 ;
      RECT 25.555 -15.749 25.645 -14.742 ;
      RECT 25.555 -15.225 25.695 -15.055 ;
      RECT 25.555 -14.328 25.645 -13.321 ;
      RECT 25.555 -14.015 25.695 -13.845 ;
      RECT 25.555 -12.519 25.645 -11.512 ;
      RECT 25.555 -11.995 25.695 -11.825 ;
      RECT 25.555 -11.098 25.645 -10.091 ;
      RECT 25.555 -10.785 25.695 -10.615 ;
      RECT 25.555 -9.289 25.645 -8.282 ;
      RECT 25.555 -8.765 25.695 -8.595 ;
      RECT 25.555 -7.868 25.645 -6.861 ;
      RECT 25.555 -7.555 25.695 -7.385 ;
      RECT 25.555 -6.059 25.645 -5.052 ;
      RECT 25.555 -5.535 25.695 -5.365 ;
      RECT 25.555 -4.638 25.645 -3.631 ;
      RECT 25.555 -4.325 25.695 -4.155 ;
      RECT 25.555 -2.829 25.645 -1.822 ;
      RECT 25.555 -2.305 25.695 -2.135 ;
      RECT 25.555 -1.408 25.645 -0.401 ;
      RECT 25.555 -1.095 25.695 -0.925 ;
      RECT 25.555 0.401 25.645 1.408 ;
      RECT 25.555 0.925 25.695 1.095 ;
      RECT 25.24 -114.685 25.41 -114.515 ;
      RECT 25.31 -114.895 25.41 -114.515 ;
      RECT 24.755 -101.538 24.845 -100.53 ;
      RECT 24.705 -100.935 24.845 -100.765 ;
      RECT 24.755 -99.73 24.845 -98.722 ;
      RECT 24.705 -99.495 24.845 -99.325 ;
      RECT 24.755 -98.308 24.845 -97.3 ;
      RECT 24.705 -97.705 24.845 -97.535 ;
      RECT 24.755 -96.5 24.845 -95.492 ;
      RECT 24.705 -96.265 24.845 -96.095 ;
      RECT 24.755 -95.078 24.845 -94.07 ;
      RECT 24.705 -94.475 24.845 -94.305 ;
      RECT 24.755 -93.27 24.845 -92.262 ;
      RECT 24.705 -93.035 24.845 -92.865 ;
      RECT 24.755 -91.848 24.845 -90.84 ;
      RECT 24.705 -91.245 24.845 -91.075 ;
      RECT 24.755 -90.04 24.845 -89.032 ;
      RECT 24.705 -89.805 24.845 -89.635 ;
      RECT 24.755 -88.618 24.845 -87.61 ;
      RECT 24.705 -88.015 24.845 -87.845 ;
      RECT 24.755 -86.81 24.845 -85.802 ;
      RECT 24.705 -86.575 24.845 -86.405 ;
      RECT 24.755 -85.388 24.845 -84.38 ;
      RECT 24.705 -84.785 24.845 -84.615 ;
      RECT 24.755 -83.58 24.845 -82.572 ;
      RECT 24.705 -83.345 24.845 -83.175 ;
      RECT 24.755 -82.158 24.845 -81.15 ;
      RECT 24.705 -81.555 24.845 -81.385 ;
      RECT 24.755 -80.35 24.845 -79.342 ;
      RECT 24.705 -80.115 24.845 -79.945 ;
      RECT 24.755 -78.928 24.845 -77.92 ;
      RECT 24.705 -78.325 24.845 -78.155 ;
      RECT 24.755 -77.12 24.845 -76.112 ;
      RECT 24.705 -76.885 24.845 -76.715 ;
      RECT 24.755 -75.698 24.845 -74.69 ;
      RECT 24.705 -75.095 24.845 -74.925 ;
      RECT 24.755 -73.89 24.845 -72.882 ;
      RECT 24.705 -73.655 24.845 -73.485 ;
      RECT 24.755 -72.468 24.845 -71.46 ;
      RECT 24.705 -71.865 24.845 -71.695 ;
      RECT 24.755 -70.66 24.845 -69.652 ;
      RECT 24.705 -70.425 24.845 -70.255 ;
      RECT 24.755 -69.238 24.845 -68.23 ;
      RECT 24.705 -68.635 24.845 -68.465 ;
      RECT 24.755 -67.43 24.845 -66.422 ;
      RECT 24.705 -67.195 24.845 -67.025 ;
      RECT 24.755 -66.008 24.845 -65 ;
      RECT 24.705 -65.405 24.845 -65.235 ;
      RECT 24.755 -64.2 24.845 -63.192 ;
      RECT 24.705 -63.965 24.845 -63.795 ;
      RECT 24.755 -62.778 24.845 -61.77 ;
      RECT 24.705 -62.175 24.845 -62.005 ;
      RECT 24.755 -60.97 24.845 -59.962 ;
      RECT 24.705 -60.735 24.845 -60.565 ;
      RECT 24.755 -59.548 24.845 -58.54 ;
      RECT 24.705 -58.945 24.845 -58.775 ;
      RECT 24.755 -57.74 24.845 -56.732 ;
      RECT 24.705 -57.505 24.845 -57.335 ;
      RECT 24.755 -56.318 24.845 -55.31 ;
      RECT 24.705 -55.715 24.845 -55.545 ;
      RECT 24.755 -54.51 24.845 -53.502 ;
      RECT 24.705 -54.275 24.845 -54.105 ;
      RECT 24.755 -53.088 24.845 -52.08 ;
      RECT 24.705 -52.485 24.845 -52.315 ;
      RECT 24.755 -51.28 24.845 -50.272 ;
      RECT 24.705 -51.045 24.845 -50.875 ;
      RECT 24.755 -49.858 24.845 -48.85 ;
      RECT 24.705 -49.255 24.845 -49.085 ;
      RECT 24.755 -48.05 24.845 -47.042 ;
      RECT 24.705 -47.815 24.845 -47.645 ;
      RECT 24.755 -46.628 24.845 -45.62 ;
      RECT 24.705 -46.025 24.845 -45.855 ;
      RECT 24.755 -44.82 24.845 -43.812 ;
      RECT 24.705 -44.585 24.845 -44.415 ;
      RECT 24.755 -43.398 24.845 -42.39 ;
      RECT 24.705 -42.795 24.845 -42.625 ;
      RECT 24.755 -41.59 24.845 -40.582 ;
      RECT 24.705 -41.355 24.845 -41.185 ;
      RECT 24.755 -40.168 24.845 -39.16 ;
      RECT 24.705 -39.565 24.845 -39.395 ;
      RECT 24.755 -38.36 24.845 -37.352 ;
      RECT 24.705 -38.125 24.845 -37.955 ;
      RECT 24.755 -36.938 24.845 -35.93 ;
      RECT 24.705 -36.335 24.845 -36.165 ;
      RECT 24.755 -35.13 24.845 -34.122 ;
      RECT 24.705 -34.895 24.845 -34.725 ;
      RECT 24.755 -33.708 24.845 -32.7 ;
      RECT 24.705 -33.105 24.845 -32.935 ;
      RECT 24.755 -31.9 24.845 -30.892 ;
      RECT 24.705 -31.665 24.845 -31.495 ;
      RECT 24.755 -30.478 24.845 -29.47 ;
      RECT 24.705 -29.875 24.845 -29.705 ;
      RECT 24.755 -28.67 24.845 -27.662 ;
      RECT 24.705 -28.435 24.845 -28.265 ;
      RECT 24.755 -27.248 24.845 -26.24 ;
      RECT 24.705 -26.645 24.845 -26.475 ;
      RECT 24.755 -25.44 24.845 -24.432 ;
      RECT 24.705 -25.205 24.845 -25.035 ;
      RECT 24.755 -24.018 24.845 -23.01 ;
      RECT 24.705 -23.415 24.845 -23.245 ;
      RECT 24.755 -22.21 24.845 -21.202 ;
      RECT 24.705 -21.975 24.845 -21.805 ;
      RECT 24.755 -20.788 24.845 -19.78 ;
      RECT 24.705 -20.185 24.845 -20.015 ;
      RECT 24.755 -18.98 24.845 -17.972 ;
      RECT 24.705 -18.745 24.845 -18.575 ;
      RECT 24.755 -17.558 24.845 -16.55 ;
      RECT 24.705 -16.955 24.845 -16.785 ;
      RECT 24.755 -15.75 24.845 -14.742 ;
      RECT 24.705 -15.515 24.845 -15.345 ;
      RECT 24.755 -14.328 24.845 -13.32 ;
      RECT 24.705 -13.725 24.845 -13.555 ;
      RECT 24.755 -12.52 24.845 -11.512 ;
      RECT 24.705 -12.285 24.845 -12.115 ;
      RECT 24.755 -11.098 24.845 -10.09 ;
      RECT 24.705 -10.495 24.845 -10.325 ;
      RECT 24.755 -9.29 24.845 -8.282 ;
      RECT 24.705 -9.055 24.845 -8.885 ;
      RECT 24.755 -7.868 24.845 -6.86 ;
      RECT 24.705 -7.265 24.845 -7.095 ;
      RECT 24.755 -6.06 24.845 -5.052 ;
      RECT 24.705 -5.825 24.845 -5.655 ;
      RECT 24.755 -4.638 24.845 -3.63 ;
      RECT 24.705 -4.035 24.845 -3.865 ;
      RECT 24.755 -2.83 24.845 -1.822 ;
      RECT 24.705 -2.595 24.845 -2.425 ;
      RECT 24.755 -1.408 24.845 -0.4 ;
      RECT 24.705 -0.805 24.845 -0.635 ;
      RECT 24.755 0.4 24.845 1.408 ;
      RECT 24.705 0.635 24.845 0.805 ;
      RECT 24.355 -101.538 24.445 -100.531 ;
      RECT 24.355 -101.225 24.495 -101.055 ;
      RECT 24.355 -99.729 24.445 -98.722 ;
      RECT 24.355 -99.205 24.495 -99.035 ;
      RECT 24.355 -98.308 24.445 -97.301 ;
      RECT 24.355 -97.995 24.495 -97.825 ;
      RECT 24.355 -96.499 24.445 -95.492 ;
      RECT 24.355 -95.975 24.495 -95.805 ;
      RECT 24.355 -95.078 24.445 -94.071 ;
      RECT 24.355 -94.765 24.495 -94.595 ;
      RECT 24.355 -93.269 24.445 -92.262 ;
      RECT 24.355 -92.745 24.495 -92.575 ;
      RECT 24.355 -91.848 24.445 -90.841 ;
      RECT 24.355 -91.535 24.495 -91.365 ;
      RECT 24.355 -90.039 24.445 -89.032 ;
      RECT 24.355 -89.515 24.495 -89.345 ;
      RECT 24.355 -88.618 24.445 -87.611 ;
      RECT 24.355 -88.305 24.495 -88.135 ;
      RECT 24.355 -86.809 24.445 -85.802 ;
      RECT 24.355 -86.285 24.495 -86.115 ;
      RECT 24.355 -85.388 24.445 -84.381 ;
      RECT 24.355 -85.075 24.495 -84.905 ;
      RECT 24.355 -83.579 24.445 -82.572 ;
      RECT 24.355 -83.055 24.495 -82.885 ;
      RECT 24.355 -82.158 24.445 -81.151 ;
      RECT 24.355 -81.845 24.495 -81.675 ;
      RECT 24.355 -80.349 24.445 -79.342 ;
      RECT 24.355 -79.825 24.495 -79.655 ;
      RECT 24.355 -78.928 24.445 -77.921 ;
      RECT 24.355 -78.615 24.495 -78.445 ;
      RECT 24.355 -77.119 24.445 -76.112 ;
      RECT 24.355 -76.595 24.495 -76.425 ;
      RECT 24.355 -75.698 24.445 -74.691 ;
      RECT 24.355 -75.385 24.495 -75.215 ;
      RECT 24.355 -73.889 24.445 -72.882 ;
      RECT 24.355 -73.365 24.495 -73.195 ;
      RECT 24.355 -72.468 24.445 -71.461 ;
      RECT 24.355 -72.155 24.495 -71.985 ;
      RECT 24.355 -70.659 24.445 -69.652 ;
      RECT 24.355 -70.135 24.495 -69.965 ;
      RECT 24.355 -69.238 24.445 -68.231 ;
      RECT 24.355 -68.925 24.495 -68.755 ;
      RECT 24.355 -67.429 24.445 -66.422 ;
      RECT 24.355 -66.905 24.495 -66.735 ;
      RECT 24.355 -66.008 24.445 -65.001 ;
      RECT 24.355 -65.695 24.495 -65.525 ;
      RECT 24.355 -64.199 24.445 -63.192 ;
      RECT 24.355 -63.675 24.495 -63.505 ;
      RECT 24.355 -62.778 24.445 -61.771 ;
      RECT 24.355 -62.465 24.495 -62.295 ;
      RECT 24.355 -60.969 24.445 -59.962 ;
      RECT 24.355 -60.445 24.495 -60.275 ;
      RECT 24.355 -59.548 24.445 -58.541 ;
      RECT 24.355 -59.235 24.495 -59.065 ;
      RECT 24.355 -57.739 24.445 -56.732 ;
      RECT 24.355 -57.215 24.495 -57.045 ;
      RECT 24.355 -56.318 24.445 -55.311 ;
      RECT 24.355 -56.005 24.495 -55.835 ;
      RECT 24.355 -54.509 24.445 -53.502 ;
      RECT 24.355 -53.985 24.495 -53.815 ;
      RECT 24.355 -53.088 24.445 -52.081 ;
      RECT 24.355 -52.775 24.495 -52.605 ;
      RECT 24.355 -51.279 24.445 -50.272 ;
      RECT 24.355 -50.755 24.495 -50.585 ;
      RECT 24.355 -49.858 24.445 -48.851 ;
      RECT 24.355 -49.545 24.495 -49.375 ;
      RECT 24.355 -48.049 24.445 -47.042 ;
      RECT 24.355 -47.525 24.495 -47.355 ;
      RECT 24.355 -46.628 24.445 -45.621 ;
      RECT 24.355 -46.315 24.495 -46.145 ;
      RECT 24.355 -44.819 24.445 -43.812 ;
      RECT 24.355 -44.295 24.495 -44.125 ;
      RECT 24.355 -43.398 24.445 -42.391 ;
      RECT 24.355 -43.085 24.495 -42.915 ;
      RECT 24.355 -41.589 24.445 -40.582 ;
      RECT 24.355 -41.065 24.495 -40.895 ;
      RECT 24.355 -40.168 24.445 -39.161 ;
      RECT 24.355 -39.855 24.495 -39.685 ;
      RECT 24.355 -38.359 24.445 -37.352 ;
      RECT 24.355 -37.835 24.495 -37.665 ;
      RECT 24.355 -36.938 24.445 -35.931 ;
      RECT 24.355 -36.625 24.495 -36.455 ;
      RECT 24.355 -35.129 24.445 -34.122 ;
      RECT 24.355 -34.605 24.495 -34.435 ;
      RECT 24.355 -33.708 24.445 -32.701 ;
      RECT 24.355 -33.395 24.495 -33.225 ;
      RECT 24.355 -31.899 24.445 -30.892 ;
      RECT 24.355 -31.375 24.495 -31.205 ;
      RECT 24.355 -30.478 24.445 -29.471 ;
      RECT 24.355 -30.165 24.495 -29.995 ;
      RECT 24.355 -28.669 24.445 -27.662 ;
      RECT 24.355 -28.145 24.495 -27.975 ;
      RECT 24.355 -27.248 24.445 -26.241 ;
      RECT 24.355 -26.935 24.495 -26.765 ;
      RECT 24.355 -25.439 24.445 -24.432 ;
      RECT 24.355 -24.915 24.495 -24.745 ;
      RECT 24.355 -24.018 24.445 -23.011 ;
      RECT 24.355 -23.705 24.495 -23.535 ;
      RECT 24.355 -22.209 24.445 -21.202 ;
      RECT 24.355 -21.685 24.495 -21.515 ;
      RECT 24.355 -20.788 24.445 -19.781 ;
      RECT 24.355 -20.475 24.495 -20.305 ;
      RECT 24.355 -18.979 24.445 -17.972 ;
      RECT 24.355 -18.455 24.495 -18.285 ;
      RECT 24.355 -17.558 24.445 -16.551 ;
      RECT 24.355 -17.245 24.495 -17.075 ;
      RECT 24.355 -15.749 24.445 -14.742 ;
      RECT 24.355 -15.225 24.495 -15.055 ;
      RECT 24.355 -14.328 24.445 -13.321 ;
      RECT 24.355 -14.015 24.495 -13.845 ;
      RECT 24.355 -12.519 24.445 -11.512 ;
      RECT 24.355 -11.995 24.495 -11.825 ;
      RECT 24.355 -11.098 24.445 -10.091 ;
      RECT 24.355 -10.785 24.495 -10.615 ;
      RECT 24.355 -9.289 24.445 -8.282 ;
      RECT 24.355 -8.765 24.495 -8.595 ;
      RECT 24.355 -7.868 24.445 -6.861 ;
      RECT 24.355 -7.555 24.495 -7.385 ;
      RECT 24.355 -6.059 24.445 -5.052 ;
      RECT 24.355 -5.535 24.495 -5.365 ;
      RECT 24.355 -4.638 24.445 -3.631 ;
      RECT 24.355 -4.325 24.495 -4.155 ;
      RECT 24.355 -2.829 24.445 -1.822 ;
      RECT 24.355 -2.305 24.495 -2.135 ;
      RECT 24.355 -1.408 24.445 -0.401 ;
      RECT 24.355 -1.095 24.495 -0.925 ;
      RECT 24.355 0.401 24.445 1.408 ;
      RECT 24.355 0.925 24.495 1.095 ;
      RECT 20.185 -108.935 23.965 -108.815 ;
      RECT 21.505 -109.475 21.605 -108.815 ;
      RECT 20.945 -109.475 21.045 -108.815 ;
      RECT 20.385 -109.475 20.485 -108.815 ;
      RECT 23.555 -101.538 23.645 -100.53 ;
      RECT 23.505 -100.935 23.645 -100.765 ;
      RECT 23.555 -99.73 23.645 -98.722 ;
      RECT 23.505 -99.495 23.645 -99.325 ;
      RECT 23.555 -98.308 23.645 -97.3 ;
      RECT 23.505 -97.705 23.645 -97.535 ;
      RECT 23.555 -96.5 23.645 -95.492 ;
      RECT 23.505 -96.265 23.645 -96.095 ;
      RECT 23.555 -95.078 23.645 -94.07 ;
      RECT 23.505 -94.475 23.645 -94.305 ;
      RECT 23.555 -93.27 23.645 -92.262 ;
      RECT 23.505 -93.035 23.645 -92.865 ;
      RECT 23.555 -91.848 23.645 -90.84 ;
      RECT 23.505 -91.245 23.645 -91.075 ;
      RECT 23.555 -90.04 23.645 -89.032 ;
      RECT 23.505 -89.805 23.645 -89.635 ;
      RECT 23.555 -88.618 23.645 -87.61 ;
      RECT 23.505 -88.015 23.645 -87.845 ;
      RECT 23.555 -86.81 23.645 -85.802 ;
      RECT 23.505 -86.575 23.645 -86.405 ;
      RECT 23.555 -85.388 23.645 -84.38 ;
      RECT 23.505 -84.785 23.645 -84.615 ;
      RECT 23.555 -83.58 23.645 -82.572 ;
      RECT 23.505 -83.345 23.645 -83.175 ;
      RECT 23.555 -82.158 23.645 -81.15 ;
      RECT 23.505 -81.555 23.645 -81.385 ;
      RECT 23.555 -80.35 23.645 -79.342 ;
      RECT 23.505 -80.115 23.645 -79.945 ;
      RECT 23.555 -78.928 23.645 -77.92 ;
      RECT 23.505 -78.325 23.645 -78.155 ;
      RECT 23.555 -77.12 23.645 -76.112 ;
      RECT 23.505 -76.885 23.645 -76.715 ;
      RECT 23.555 -75.698 23.645 -74.69 ;
      RECT 23.505 -75.095 23.645 -74.925 ;
      RECT 23.555 -73.89 23.645 -72.882 ;
      RECT 23.505 -73.655 23.645 -73.485 ;
      RECT 23.555 -72.468 23.645 -71.46 ;
      RECT 23.505 -71.865 23.645 -71.695 ;
      RECT 23.555 -70.66 23.645 -69.652 ;
      RECT 23.505 -70.425 23.645 -70.255 ;
      RECT 23.555 -69.238 23.645 -68.23 ;
      RECT 23.505 -68.635 23.645 -68.465 ;
      RECT 23.555 -67.43 23.645 -66.422 ;
      RECT 23.505 -67.195 23.645 -67.025 ;
      RECT 23.555 -66.008 23.645 -65 ;
      RECT 23.505 -65.405 23.645 -65.235 ;
      RECT 23.555 -64.2 23.645 -63.192 ;
      RECT 23.505 -63.965 23.645 -63.795 ;
      RECT 23.555 -62.778 23.645 -61.77 ;
      RECT 23.505 -62.175 23.645 -62.005 ;
      RECT 23.555 -60.97 23.645 -59.962 ;
      RECT 23.505 -60.735 23.645 -60.565 ;
      RECT 23.555 -59.548 23.645 -58.54 ;
      RECT 23.505 -58.945 23.645 -58.775 ;
      RECT 23.555 -57.74 23.645 -56.732 ;
      RECT 23.505 -57.505 23.645 -57.335 ;
      RECT 23.555 -56.318 23.645 -55.31 ;
      RECT 23.505 -55.715 23.645 -55.545 ;
      RECT 23.555 -54.51 23.645 -53.502 ;
      RECT 23.505 -54.275 23.645 -54.105 ;
      RECT 23.555 -53.088 23.645 -52.08 ;
      RECT 23.505 -52.485 23.645 -52.315 ;
      RECT 23.555 -51.28 23.645 -50.272 ;
      RECT 23.505 -51.045 23.645 -50.875 ;
      RECT 23.555 -49.858 23.645 -48.85 ;
      RECT 23.505 -49.255 23.645 -49.085 ;
      RECT 23.555 -48.05 23.645 -47.042 ;
      RECT 23.505 -47.815 23.645 -47.645 ;
      RECT 23.555 -46.628 23.645 -45.62 ;
      RECT 23.505 -46.025 23.645 -45.855 ;
      RECT 23.555 -44.82 23.645 -43.812 ;
      RECT 23.505 -44.585 23.645 -44.415 ;
      RECT 23.555 -43.398 23.645 -42.39 ;
      RECT 23.505 -42.795 23.645 -42.625 ;
      RECT 23.555 -41.59 23.645 -40.582 ;
      RECT 23.505 -41.355 23.645 -41.185 ;
      RECT 23.555 -40.168 23.645 -39.16 ;
      RECT 23.505 -39.565 23.645 -39.395 ;
      RECT 23.555 -38.36 23.645 -37.352 ;
      RECT 23.505 -38.125 23.645 -37.955 ;
      RECT 23.555 -36.938 23.645 -35.93 ;
      RECT 23.505 -36.335 23.645 -36.165 ;
      RECT 23.555 -35.13 23.645 -34.122 ;
      RECT 23.505 -34.895 23.645 -34.725 ;
      RECT 23.555 -33.708 23.645 -32.7 ;
      RECT 23.505 -33.105 23.645 -32.935 ;
      RECT 23.555 -31.9 23.645 -30.892 ;
      RECT 23.505 -31.665 23.645 -31.495 ;
      RECT 23.555 -30.478 23.645 -29.47 ;
      RECT 23.505 -29.875 23.645 -29.705 ;
      RECT 23.555 -28.67 23.645 -27.662 ;
      RECT 23.505 -28.435 23.645 -28.265 ;
      RECT 23.555 -27.248 23.645 -26.24 ;
      RECT 23.505 -26.645 23.645 -26.475 ;
      RECT 23.555 -25.44 23.645 -24.432 ;
      RECT 23.505 -25.205 23.645 -25.035 ;
      RECT 23.555 -24.018 23.645 -23.01 ;
      RECT 23.505 -23.415 23.645 -23.245 ;
      RECT 23.555 -22.21 23.645 -21.202 ;
      RECT 23.505 -21.975 23.645 -21.805 ;
      RECT 23.555 -20.788 23.645 -19.78 ;
      RECT 23.505 -20.185 23.645 -20.015 ;
      RECT 23.555 -18.98 23.645 -17.972 ;
      RECT 23.505 -18.745 23.645 -18.575 ;
      RECT 23.555 -17.558 23.645 -16.55 ;
      RECT 23.505 -16.955 23.645 -16.785 ;
      RECT 23.555 -15.75 23.645 -14.742 ;
      RECT 23.505 -15.515 23.645 -15.345 ;
      RECT 23.555 -14.328 23.645 -13.32 ;
      RECT 23.505 -13.725 23.645 -13.555 ;
      RECT 23.555 -12.52 23.645 -11.512 ;
      RECT 23.505 -12.285 23.645 -12.115 ;
      RECT 23.555 -11.098 23.645 -10.09 ;
      RECT 23.505 -10.495 23.645 -10.325 ;
      RECT 23.555 -9.29 23.645 -8.282 ;
      RECT 23.505 -9.055 23.645 -8.885 ;
      RECT 23.555 -7.868 23.645 -6.86 ;
      RECT 23.505 -7.265 23.645 -7.095 ;
      RECT 23.555 -6.06 23.645 -5.052 ;
      RECT 23.505 -5.825 23.645 -5.655 ;
      RECT 23.555 -4.638 23.645 -3.63 ;
      RECT 23.505 -4.035 23.645 -3.865 ;
      RECT 23.555 -2.83 23.645 -1.822 ;
      RECT 23.505 -2.595 23.645 -2.425 ;
      RECT 23.555 -1.408 23.645 -0.4 ;
      RECT 23.505 -0.805 23.645 -0.635 ;
      RECT 23.555 0.4 23.645 1.408 ;
      RECT 23.505 0.635 23.645 0.805 ;
      RECT 22.125 -111.685 23.605 -111.585 ;
      RECT 22.125 -112.195 22.225 -111.585 ;
      RECT 22.345 -109.15 23.605 -109.05 ;
      RECT 23.505 -109.475 23.605 -109.05 ;
      RECT 22.945 -109.475 23.045 -109.05 ;
      RECT 22.385 -109.475 22.485 -109.05 ;
      RECT 23.155 -101.538 23.245 -100.531 ;
      RECT 23.155 -101.225 23.295 -101.055 ;
      RECT 23.155 -99.729 23.245 -98.722 ;
      RECT 23.155 -99.205 23.295 -99.035 ;
      RECT 23.155 -98.308 23.245 -97.301 ;
      RECT 23.155 -97.995 23.295 -97.825 ;
      RECT 23.155 -96.499 23.245 -95.492 ;
      RECT 23.155 -95.975 23.295 -95.805 ;
      RECT 23.155 -95.078 23.245 -94.071 ;
      RECT 23.155 -94.765 23.295 -94.595 ;
      RECT 23.155 -93.269 23.245 -92.262 ;
      RECT 23.155 -92.745 23.295 -92.575 ;
      RECT 23.155 -91.848 23.245 -90.841 ;
      RECT 23.155 -91.535 23.295 -91.365 ;
      RECT 23.155 -90.039 23.245 -89.032 ;
      RECT 23.155 -89.515 23.295 -89.345 ;
      RECT 23.155 -88.618 23.245 -87.611 ;
      RECT 23.155 -88.305 23.295 -88.135 ;
      RECT 23.155 -86.809 23.245 -85.802 ;
      RECT 23.155 -86.285 23.295 -86.115 ;
      RECT 23.155 -85.388 23.245 -84.381 ;
      RECT 23.155 -85.075 23.295 -84.905 ;
      RECT 23.155 -83.579 23.245 -82.572 ;
      RECT 23.155 -83.055 23.295 -82.885 ;
      RECT 23.155 -82.158 23.245 -81.151 ;
      RECT 23.155 -81.845 23.295 -81.675 ;
      RECT 23.155 -80.349 23.245 -79.342 ;
      RECT 23.155 -79.825 23.295 -79.655 ;
      RECT 23.155 -78.928 23.245 -77.921 ;
      RECT 23.155 -78.615 23.295 -78.445 ;
      RECT 23.155 -77.119 23.245 -76.112 ;
      RECT 23.155 -76.595 23.295 -76.425 ;
      RECT 23.155 -75.698 23.245 -74.691 ;
      RECT 23.155 -75.385 23.295 -75.215 ;
      RECT 23.155 -73.889 23.245 -72.882 ;
      RECT 23.155 -73.365 23.295 -73.195 ;
      RECT 23.155 -72.468 23.245 -71.461 ;
      RECT 23.155 -72.155 23.295 -71.985 ;
      RECT 23.155 -70.659 23.245 -69.652 ;
      RECT 23.155 -70.135 23.295 -69.965 ;
      RECT 23.155 -69.238 23.245 -68.231 ;
      RECT 23.155 -68.925 23.295 -68.755 ;
      RECT 23.155 -67.429 23.245 -66.422 ;
      RECT 23.155 -66.905 23.295 -66.735 ;
      RECT 23.155 -66.008 23.245 -65.001 ;
      RECT 23.155 -65.695 23.295 -65.525 ;
      RECT 23.155 -64.199 23.245 -63.192 ;
      RECT 23.155 -63.675 23.295 -63.505 ;
      RECT 23.155 -62.778 23.245 -61.771 ;
      RECT 23.155 -62.465 23.295 -62.295 ;
      RECT 23.155 -60.969 23.245 -59.962 ;
      RECT 23.155 -60.445 23.295 -60.275 ;
      RECT 23.155 -59.548 23.245 -58.541 ;
      RECT 23.155 -59.235 23.295 -59.065 ;
      RECT 23.155 -57.739 23.245 -56.732 ;
      RECT 23.155 -57.215 23.295 -57.045 ;
      RECT 23.155 -56.318 23.245 -55.311 ;
      RECT 23.155 -56.005 23.295 -55.835 ;
      RECT 23.155 -54.509 23.245 -53.502 ;
      RECT 23.155 -53.985 23.295 -53.815 ;
      RECT 23.155 -53.088 23.245 -52.081 ;
      RECT 23.155 -52.775 23.295 -52.605 ;
      RECT 23.155 -51.279 23.245 -50.272 ;
      RECT 23.155 -50.755 23.295 -50.585 ;
      RECT 23.155 -49.858 23.245 -48.851 ;
      RECT 23.155 -49.545 23.295 -49.375 ;
      RECT 23.155 -48.049 23.245 -47.042 ;
      RECT 23.155 -47.525 23.295 -47.355 ;
      RECT 23.155 -46.628 23.245 -45.621 ;
      RECT 23.155 -46.315 23.295 -46.145 ;
      RECT 23.155 -44.819 23.245 -43.812 ;
      RECT 23.155 -44.295 23.295 -44.125 ;
      RECT 23.155 -43.398 23.245 -42.391 ;
      RECT 23.155 -43.085 23.295 -42.915 ;
      RECT 23.155 -41.589 23.245 -40.582 ;
      RECT 23.155 -41.065 23.295 -40.895 ;
      RECT 23.155 -40.168 23.245 -39.161 ;
      RECT 23.155 -39.855 23.295 -39.685 ;
      RECT 23.155 -38.359 23.245 -37.352 ;
      RECT 23.155 -37.835 23.295 -37.665 ;
      RECT 23.155 -36.938 23.245 -35.931 ;
      RECT 23.155 -36.625 23.295 -36.455 ;
      RECT 23.155 -35.129 23.245 -34.122 ;
      RECT 23.155 -34.605 23.295 -34.435 ;
      RECT 23.155 -33.708 23.245 -32.701 ;
      RECT 23.155 -33.395 23.295 -33.225 ;
      RECT 23.155 -31.899 23.245 -30.892 ;
      RECT 23.155 -31.375 23.295 -31.205 ;
      RECT 23.155 -30.478 23.245 -29.471 ;
      RECT 23.155 -30.165 23.295 -29.995 ;
      RECT 23.155 -28.669 23.245 -27.662 ;
      RECT 23.155 -28.145 23.295 -27.975 ;
      RECT 23.155 -27.248 23.245 -26.241 ;
      RECT 23.155 -26.935 23.295 -26.765 ;
      RECT 23.155 -25.439 23.245 -24.432 ;
      RECT 23.155 -24.915 23.295 -24.745 ;
      RECT 23.155 -24.018 23.245 -23.011 ;
      RECT 23.155 -23.705 23.295 -23.535 ;
      RECT 23.155 -22.209 23.245 -21.202 ;
      RECT 23.155 -21.685 23.295 -21.515 ;
      RECT 23.155 -20.788 23.245 -19.781 ;
      RECT 23.155 -20.475 23.295 -20.305 ;
      RECT 23.155 -18.979 23.245 -17.972 ;
      RECT 23.155 -18.455 23.295 -18.285 ;
      RECT 23.155 -17.558 23.245 -16.551 ;
      RECT 23.155 -17.245 23.295 -17.075 ;
      RECT 23.155 -15.749 23.245 -14.742 ;
      RECT 23.155 -15.225 23.295 -15.055 ;
      RECT 23.155 -14.328 23.245 -13.321 ;
      RECT 23.155 -14.015 23.295 -13.845 ;
      RECT 23.155 -12.519 23.245 -11.512 ;
      RECT 23.155 -11.995 23.295 -11.825 ;
      RECT 23.155 -11.098 23.245 -10.091 ;
      RECT 23.155 -10.785 23.295 -10.615 ;
      RECT 23.155 -9.289 23.245 -8.282 ;
      RECT 23.155 -8.765 23.295 -8.595 ;
      RECT 23.155 -7.868 23.245 -6.861 ;
      RECT 23.155 -7.555 23.295 -7.385 ;
      RECT 23.155 -6.059 23.245 -5.052 ;
      RECT 23.155 -5.535 23.295 -5.365 ;
      RECT 23.155 -4.638 23.245 -3.631 ;
      RECT 23.155 -4.325 23.295 -4.155 ;
      RECT 23.155 -2.829 23.245 -1.822 ;
      RECT 23.155 -2.305 23.295 -2.135 ;
      RECT 23.155 -1.408 23.245 -0.401 ;
      RECT 23.155 -1.095 23.295 -0.925 ;
      RECT 23.155 0.401 23.245 1.408 ;
      RECT 23.155 0.925 23.295 1.095 ;
      RECT 22.485 -111.495 22.655 -111.385 ;
      RECT 19.335 -111.495 22.655 -111.395 ;
      RECT 22.355 -101.538 22.445 -100.53 ;
      RECT 22.305 -100.935 22.445 -100.765 ;
      RECT 22.355 -99.73 22.445 -98.722 ;
      RECT 22.305 -99.495 22.445 -99.325 ;
      RECT 22.355 -98.308 22.445 -97.3 ;
      RECT 22.305 -97.705 22.445 -97.535 ;
      RECT 22.355 -96.5 22.445 -95.492 ;
      RECT 22.305 -96.265 22.445 -96.095 ;
      RECT 22.355 -95.078 22.445 -94.07 ;
      RECT 22.305 -94.475 22.445 -94.305 ;
      RECT 22.355 -93.27 22.445 -92.262 ;
      RECT 22.305 -93.035 22.445 -92.865 ;
      RECT 22.355 -91.848 22.445 -90.84 ;
      RECT 22.305 -91.245 22.445 -91.075 ;
      RECT 22.355 -90.04 22.445 -89.032 ;
      RECT 22.305 -89.805 22.445 -89.635 ;
      RECT 22.355 -88.618 22.445 -87.61 ;
      RECT 22.305 -88.015 22.445 -87.845 ;
      RECT 22.355 -86.81 22.445 -85.802 ;
      RECT 22.305 -86.575 22.445 -86.405 ;
      RECT 22.355 -85.388 22.445 -84.38 ;
      RECT 22.305 -84.785 22.445 -84.615 ;
      RECT 22.355 -83.58 22.445 -82.572 ;
      RECT 22.305 -83.345 22.445 -83.175 ;
      RECT 22.355 -82.158 22.445 -81.15 ;
      RECT 22.305 -81.555 22.445 -81.385 ;
      RECT 22.355 -80.35 22.445 -79.342 ;
      RECT 22.305 -80.115 22.445 -79.945 ;
      RECT 22.355 -78.928 22.445 -77.92 ;
      RECT 22.305 -78.325 22.445 -78.155 ;
      RECT 22.355 -77.12 22.445 -76.112 ;
      RECT 22.305 -76.885 22.445 -76.715 ;
      RECT 22.355 -75.698 22.445 -74.69 ;
      RECT 22.305 -75.095 22.445 -74.925 ;
      RECT 22.355 -73.89 22.445 -72.882 ;
      RECT 22.305 -73.655 22.445 -73.485 ;
      RECT 22.355 -72.468 22.445 -71.46 ;
      RECT 22.305 -71.865 22.445 -71.695 ;
      RECT 22.355 -70.66 22.445 -69.652 ;
      RECT 22.305 -70.425 22.445 -70.255 ;
      RECT 22.355 -69.238 22.445 -68.23 ;
      RECT 22.305 -68.635 22.445 -68.465 ;
      RECT 22.355 -67.43 22.445 -66.422 ;
      RECT 22.305 -67.195 22.445 -67.025 ;
      RECT 22.355 -66.008 22.445 -65 ;
      RECT 22.305 -65.405 22.445 -65.235 ;
      RECT 22.355 -64.2 22.445 -63.192 ;
      RECT 22.305 -63.965 22.445 -63.795 ;
      RECT 22.355 -62.778 22.445 -61.77 ;
      RECT 22.305 -62.175 22.445 -62.005 ;
      RECT 22.355 -60.97 22.445 -59.962 ;
      RECT 22.305 -60.735 22.445 -60.565 ;
      RECT 22.355 -59.548 22.445 -58.54 ;
      RECT 22.305 -58.945 22.445 -58.775 ;
      RECT 22.355 -57.74 22.445 -56.732 ;
      RECT 22.305 -57.505 22.445 -57.335 ;
      RECT 22.355 -56.318 22.445 -55.31 ;
      RECT 22.305 -55.715 22.445 -55.545 ;
      RECT 22.355 -54.51 22.445 -53.502 ;
      RECT 22.305 -54.275 22.445 -54.105 ;
      RECT 22.355 -53.088 22.445 -52.08 ;
      RECT 22.305 -52.485 22.445 -52.315 ;
      RECT 22.355 -51.28 22.445 -50.272 ;
      RECT 22.305 -51.045 22.445 -50.875 ;
      RECT 22.355 -49.858 22.445 -48.85 ;
      RECT 22.305 -49.255 22.445 -49.085 ;
      RECT 22.355 -48.05 22.445 -47.042 ;
      RECT 22.305 -47.815 22.445 -47.645 ;
      RECT 22.355 -46.628 22.445 -45.62 ;
      RECT 22.305 -46.025 22.445 -45.855 ;
      RECT 22.355 -44.82 22.445 -43.812 ;
      RECT 22.305 -44.585 22.445 -44.415 ;
      RECT 22.355 -43.398 22.445 -42.39 ;
      RECT 22.305 -42.795 22.445 -42.625 ;
      RECT 22.355 -41.59 22.445 -40.582 ;
      RECT 22.305 -41.355 22.445 -41.185 ;
      RECT 22.355 -40.168 22.445 -39.16 ;
      RECT 22.305 -39.565 22.445 -39.395 ;
      RECT 22.355 -38.36 22.445 -37.352 ;
      RECT 22.305 -38.125 22.445 -37.955 ;
      RECT 22.355 -36.938 22.445 -35.93 ;
      RECT 22.305 -36.335 22.445 -36.165 ;
      RECT 22.355 -35.13 22.445 -34.122 ;
      RECT 22.305 -34.895 22.445 -34.725 ;
      RECT 22.355 -33.708 22.445 -32.7 ;
      RECT 22.305 -33.105 22.445 -32.935 ;
      RECT 22.355 -31.9 22.445 -30.892 ;
      RECT 22.305 -31.665 22.445 -31.495 ;
      RECT 22.355 -30.478 22.445 -29.47 ;
      RECT 22.305 -29.875 22.445 -29.705 ;
      RECT 22.355 -28.67 22.445 -27.662 ;
      RECT 22.305 -28.435 22.445 -28.265 ;
      RECT 22.355 -27.248 22.445 -26.24 ;
      RECT 22.305 -26.645 22.445 -26.475 ;
      RECT 22.355 -25.44 22.445 -24.432 ;
      RECT 22.305 -25.205 22.445 -25.035 ;
      RECT 22.355 -24.018 22.445 -23.01 ;
      RECT 22.305 -23.415 22.445 -23.245 ;
      RECT 22.355 -22.21 22.445 -21.202 ;
      RECT 22.305 -21.975 22.445 -21.805 ;
      RECT 22.355 -20.788 22.445 -19.78 ;
      RECT 22.305 -20.185 22.445 -20.015 ;
      RECT 22.355 -18.98 22.445 -17.972 ;
      RECT 22.305 -18.745 22.445 -18.575 ;
      RECT 22.355 -17.558 22.445 -16.55 ;
      RECT 22.305 -16.955 22.445 -16.785 ;
      RECT 22.355 -15.75 22.445 -14.742 ;
      RECT 22.305 -15.515 22.445 -15.345 ;
      RECT 22.355 -14.328 22.445 -13.32 ;
      RECT 22.305 -13.725 22.445 -13.555 ;
      RECT 22.355 -12.52 22.445 -11.512 ;
      RECT 22.305 -12.285 22.445 -12.115 ;
      RECT 22.355 -11.098 22.445 -10.09 ;
      RECT 22.305 -10.495 22.445 -10.325 ;
      RECT 22.355 -9.29 22.445 -8.282 ;
      RECT 22.305 -9.055 22.445 -8.885 ;
      RECT 22.355 -7.868 22.445 -6.86 ;
      RECT 22.305 -7.265 22.445 -7.095 ;
      RECT 22.355 -6.06 22.445 -5.052 ;
      RECT 22.305 -5.825 22.445 -5.655 ;
      RECT 22.355 -4.638 22.445 -3.63 ;
      RECT 22.305 -4.035 22.445 -3.865 ;
      RECT 22.355 -2.83 22.445 -1.822 ;
      RECT 22.305 -2.595 22.445 -2.425 ;
      RECT 22.355 -1.408 22.445 -0.4 ;
      RECT 22.305 -0.805 22.445 -0.635 ;
      RECT 22.355 0.4 22.445 1.408 ;
      RECT 22.305 0.635 22.445 0.805 ;
      RECT 21.955 -101.538 22.045 -100.531 ;
      RECT 21.955 -101.225 22.095 -101.055 ;
      RECT 21.955 -99.729 22.045 -98.722 ;
      RECT 21.955 -99.205 22.095 -99.035 ;
      RECT 21.955 -98.308 22.045 -97.301 ;
      RECT 21.955 -97.995 22.095 -97.825 ;
      RECT 21.955 -96.499 22.045 -95.492 ;
      RECT 21.955 -95.975 22.095 -95.805 ;
      RECT 21.955 -95.078 22.045 -94.071 ;
      RECT 21.955 -94.765 22.095 -94.595 ;
      RECT 21.955 -93.269 22.045 -92.262 ;
      RECT 21.955 -92.745 22.095 -92.575 ;
      RECT 21.955 -91.848 22.045 -90.841 ;
      RECT 21.955 -91.535 22.095 -91.365 ;
      RECT 21.955 -90.039 22.045 -89.032 ;
      RECT 21.955 -89.515 22.095 -89.345 ;
      RECT 21.955 -88.618 22.045 -87.611 ;
      RECT 21.955 -88.305 22.095 -88.135 ;
      RECT 21.955 -86.809 22.045 -85.802 ;
      RECT 21.955 -86.285 22.095 -86.115 ;
      RECT 21.955 -85.388 22.045 -84.381 ;
      RECT 21.955 -85.075 22.095 -84.905 ;
      RECT 21.955 -83.579 22.045 -82.572 ;
      RECT 21.955 -83.055 22.095 -82.885 ;
      RECT 21.955 -82.158 22.045 -81.151 ;
      RECT 21.955 -81.845 22.095 -81.675 ;
      RECT 21.955 -80.349 22.045 -79.342 ;
      RECT 21.955 -79.825 22.095 -79.655 ;
      RECT 21.955 -78.928 22.045 -77.921 ;
      RECT 21.955 -78.615 22.095 -78.445 ;
      RECT 21.955 -77.119 22.045 -76.112 ;
      RECT 21.955 -76.595 22.095 -76.425 ;
      RECT 21.955 -75.698 22.045 -74.691 ;
      RECT 21.955 -75.385 22.095 -75.215 ;
      RECT 21.955 -73.889 22.045 -72.882 ;
      RECT 21.955 -73.365 22.095 -73.195 ;
      RECT 21.955 -72.468 22.045 -71.461 ;
      RECT 21.955 -72.155 22.095 -71.985 ;
      RECT 21.955 -70.659 22.045 -69.652 ;
      RECT 21.955 -70.135 22.095 -69.965 ;
      RECT 21.955 -69.238 22.045 -68.231 ;
      RECT 21.955 -68.925 22.095 -68.755 ;
      RECT 21.955 -67.429 22.045 -66.422 ;
      RECT 21.955 -66.905 22.095 -66.735 ;
      RECT 21.955 -66.008 22.045 -65.001 ;
      RECT 21.955 -65.695 22.095 -65.525 ;
      RECT 21.955 -64.199 22.045 -63.192 ;
      RECT 21.955 -63.675 22.095 -63.505 ;
      RECT 21.955 -62.778 22.045 -61.771 ;
      RECT 21.955 -62.465 22.095 -62.295 ;
      RECT 21.955 -60.969 22.045 -59.962 ;
      RECT 21.955 -60.445 22.095 -60.275 ;
      RECT 21.955 -59.548 22.045 -58.541 ;
      RECT 21.955 -59.235 22.095 -59.065 ;
      RECT 21.955 -57.739 22.045 -56.732 ;
      RECT 21.955 -57.215 22.095 -57.045 ;
      RECT 21.955 -56.318 22.045 -55.311 ;
      RECT 21.955 -56.005 22.095 -55.835 ;
      RECT 21.955 -54.509 22.045 -53.502 ;
      RECT 21.955 -53.985 22.095 -53.815 ;
      RECT 21.955 -53.088 22.045 -52.081 ;
      RECT 21.955 -52.775 22.095 -52.605 ;
      RECT 21.955 -51.279 22.045 -50.272 ;
      RECT 21.955 -50.755 22.095 -50.585 ;
      RECT 21.955 -49.858 22.045 -48.851 ;
      RECT 21.955 -49.545 22.095 -49.375 ;
      RECT 21.955 -48.049 22.045 -47.042 ;
      RECT 21.955 -47.525 22.095 -47.355 ;
      RECT 21.955 -46.628 22.045 -45.621 ;
      RECT 21.955 -46.315 22.095 -46.145 ;
      RECT 21.955 -44.819 22.045 -43.812 ;
      RECT 21.955 -44.295 22.095 -44.125 ;
      RECT 21.955 -43.398 22.045 -42.391 ;
      RECT 21.955 -43.085 22.095 -42.915 ;
      RECT 21.955 -41.589 22.045 -40.582 ;
      RECT 21.955 -41.065 22.095 -40.895 ;
      RECT 21.955 -40.168 22.045 -39.161 ;
      RECT 21.955 -39.855 22.095 -39.685 ;
      RECT 21.955 -38.359 22.045 -37.352 ;
      RECT 21.955 -37.835 22.095 -37.665 ;
      RECT 21.955 -36.938 22.045 -35.931 ;
      RECT 21.955 -36.625 22.095 -36.455 ;
      RECT 21.955 -35.129 22.045 -34.122 ;
      RECT 21.955 -34.605 22.095 -34.435 ;
      RECT 21.955 -33.708 22.045 -32.701 ;
      RECT 21.955 -33.395 22.095 -33.225 ;
      RECT 21.955 -31.899 22.045 -30.892 ;
      RECT 21.955 -31.375 22.095 -31.205 ;
      RECT 21.955 -30.478 22.045 -29.471 ;
      RECT 21.955 -30.165 22.095 -29.995 ;
      RECT 21.955 -28.669 22.045 -27.662 ;
      RECT 21.955 -28.145 22.095 -27.975 ;
      RECT 21.955 -27.248 22.045 -26.241 ;
      RECT 21.955 -26.935 22.095 -26.765 ;
      RECT 21.955 -25.439 22.045 -24.432 ;
      RECT 21.955 -24.915 22.095 -24.745 ;
      RECT 21.955 -24.018 22.045 -23.011 ;
      RECT 21.955 -23.705 22.095 -23.535 ;
      RECT 21.955 -22.209 22.045 -21.202 ;
      RECT 21.955 -21.685 22.095 -21.515 ;
      RECT 21.955 -20.788 22.045 -19.781 ;
      RECT 21.955 -20.475 22.095 -20.305 ;
      RECT 21.955 -18.979 22.045 -17.972 ;
      RECT 21.955 -18.455 22.095 -18.285 ;
      RECT 21.955 -17.558 22.045 -16.551 ;
      RECT 21.955 -17.245 22.095 -17.075 ;
      RECT 21.955 -15.749 22.045 -14.742 ;
      RECT 21.955 -15.225 22.095 -15.055 ;
      RECT 21.955 -14.328 22.045 -13.321 ;
      RECT 21.955 -14.015 22.095 -13.845 ;
      RECT 21.955 -12.519 22.045 -11.512 ;
      RECT 21.955 -11.995 22.095 -11.825 ;
      RECT 21.955 -11.098 22.045 -10.091 ;
      RECT 21.955 -10.785 22.095 -10.615 ;
      RECT 21.955 -9.289 22.045 -8.282 ;
      RECT 21.955 -8.765 22.095 -8.595 ;
      RECT 21.955 -7.868 22.045 -6.861 ;
      RECT 21.955 -7.555 22.095 -7.385 ;
      RECT 21.955 -6.059 22.045 -5.052 ;
      RECT 21.955 -5.535 22.095 -5.365 ;
      RECT 21.955 -4.638 22.045 -3.631 ;
      RECT 21.955 -4.325 22.095 -4.155 ;
      RECT 21.955 -2.829 22.045 -1.822 ;
      RECT 21.955 -2.305 22.095 -2.135 ;
      RECT 21.955 -1.408 22.045 -0.401 ;
      RECT 21.955 -1.095 22.095 -0.925 ;
      RECT 21.955 0.401 22.045 1.408 ;
      RECT 21.955 0.925 22.095 1.095 ;
      RECT 20.105 -111.685 21.585 -111.585 ;
      RECT 20.105 -112.055 20.205 -111.585 ;
      RECT 19.91 -114.395 21.485 -114.275 ;
      RECT 21.385 -114.895 21.485 -114.275 ;
      RECT 20.79 -114.895 20.89 -114.275 ;
      RECT 19.91 -114.85 20.01 -114.275 ;
      RECT 21.155 -101.538 21.245 -100.53 ;
      RECT 21.105 -100.935 21.245 -100.765 ;
      RECT 21.155 -99.73 21.245 -98.722 ;
      RECT 21.105 -99.495 21.245 -99.325 ;
      RECT 21.155 -98.308 21.245 -97.3 ;
      RECT 21.105 -97.705 21.245 -97.535 ;
      RECT 21.155 -96.5 21.245 -95.492 ;
      RECT 21.105 -96.265 21.245 -96.095 ;
      RECT 21.155 -95.078 21.245 -94.07 ;
      RECT 21.105 -94.475 21.245 -94.305 ;
      RECT 21.155 -93.27 21.245 -92.262 ;
      RECT 21.105 -93.035 21.245 -92.865 ;
      RECT 21.155 -91.848 21.245 -90.84 ;
      RECT 21.105 -91.245 21.245 -91.075 ;
      RECT 21.155 -90.04 21.245 -89.032 ;
      RECT 21.105 -89.805 21.245 -89.635 ;
      RECT 21.155 -88.618 21.245 -87.61 ;
      RECT 21.105 -88.015 21.245 -87.845 ;
      RECT 21.155 -86.81 21.245 -85.802 ;
      RECT 21.105 -86.575 21.245 -86.405 ;
      RECT 21.155 -85.388 21.245 -84.38 ;
      RECT 21.105 -84.785 21.245 -84.615 ;
      RECT 21.155 -83.58 21.245 -82.572 ;
      RECT 21.105 -83.345 21.245 -83.175 ;
      RECT 21.155 -82.158 21.245 -81.15 ;
      RECT 21.105 -81.555 21.245 -81.385 ;
      RECT 21.155 -80.35 21.245 -79.342 ;
      RECT 21.105 -80.115 21.245 -79.945 ;
      RECT 21.155 -78.928 21.245 -77.92 ;
      RECT 21.105 -78.325 21.245 -78.155 ;
      RECT 21.155 -77.12 21.245 -76.112 ;
      RECT 21.105 -76.885 21.245 -76.715 ;
      RECT 21.155 -75.698 21.245 -74.69 ;
      RECT 21.105 -75.095 21.245 -74.925 ;
      RECT 21.155 -73.89 21.245 -72.882 ;
      RECT 21.105 -73.655 21.245 -73.485 ;
      RECT 21.155 -72.468 21.245 -71.46 ;
      RECT 21.105 -71.865 21.245 -71.695 ;
      RECT 21.155 -70.66 21.245 -69.652 ;
      RECT 21.105 -70.425 21.245 -70.255 ;
      RECT 21.155 -69.238 21.245 -68.23 ;
      RECT 21.105 -68.635 21.245 -68.465 ;
      RECT 21.155 -67.43 21.245 -66.422 ;
      RECT 21.105 -67.195 21.245 -67.025 ;
      RECT 21.155 -66.008 21.245 -65 ;
      RECT 21.105 -65.405 21.245 -65.235 ;
      RECT 21.155 -64.2 21.245 -63.192 ;
      RECT 21.105 -63.965 21.245 -63.795 ;
      RECT 21.155 -62.778 21.245 -61.77 ;
      RECT 21.105 -62.175 21.245 -62.005 ;
      RECT 21.155 -60.97 21.245 -59.962 ;
      RECT 21.105 -60.735 21.245 -60.565 ;
      RECT 21.155 -59.548 21.245 -58.54 ;
      RECT 21.105 -58.945 21.245 -58.775 ;
      RECT 21.155 -57.74 21.245 -56.732 ;
      RECT 21.105 -57.505 21.245 -57.335 ;
      RECT 21.155 -56.318 21.245 -55.31 ;
      RECT 21.105 -55.715 21.245 -55.545 ;
      RECT 21.155 -54.51 21.245 -53.502 ;
      RECT 21.105 -54.275 21.245 -54.105 ;
      RECT 21.155 -53.088 21.245 -52.08 ;
      RECT 21.105 -52.485 21.245 -52.315 ;
      RECT 21.155 -51.28 21.245 -50.272 ;
      RECT 21.105 -51.045 21.245 -50.875 ;
      RECT 21.155 -49.858 21.245 -48.85 ;
      RECT 21.105 -49.255 21.245 -49.085 ;
      RECT 21.155 -48.05 21.245 -47.042 ;
      RECT 21.105 -47.815 21.245 -47.645 ;
      RECT 21.155 -46.628 21.245 -45.62 ;
      RECT 21.105 -46.025 21.245 -45.855 ;
      RECT 21.155 -44.82 21.245 -43.812 ;
      RECT 21.105 -44.585 21.245 -44.415 ;
      RECT 21.155 -43.398 21.245 -42.39 ;
      RECT 21.105 -42.795 21.245 -42.625 ;
      RECT 21.155 -41.59 21.245 -40.582 ;
      RECT 21.105 -41.355 21.245 -41.185 ;
      RECT 21.155 -40.168 21.245 -39.16 ;
      RECT 21.105 -39.565 21.245 -39.395 ;
      RECT 21.155 -38.36 21.245 -37.352 ;
      RECT 21.105 -38.125 21.245 -37.955 ;
      RECT 21.155 -36.938 21.245 -35.93 ;
      RECT 21.105 -36.335 21.245 -36.165 ;
      RECT 21.155 -35.13 21.245 -34.122 ;
      RECT 21.105 -34.895 21.245 -34.725 ;
      RECT 21.155 -33.708 21.245 -32.7 ;
      RECT 21.105 -33.105 21.245 -32.935 ;
      RECT 21.155 -31.9 21.245 -30.892 ;
      RECT 21.105 -31.665 21.245 -31.495 ;
      RECT 21.155 -30.478 21.245 -29.47 ;
      RECT 21.105 -29.875 21.245 -29.705 ;
      RECT 21.155 -28.67 21.245 -27.662 ;
      RECT 21.105 -28.435 21.245 -28.265 ;
      RECT 21.155 -27.248 21.245 -26.24 ;
      RECT 21.105 -26.645 21.245 -26.475 ;
      RECT 21.155 -25.44 21.245 -24.432 ;
      RECT 21.105 -25.205 21.245 -25.035 ;
      RECT 21.155 -24.018 21.245 -23.01 ;
      RECT 21.105 -23.415 21.245 -23.245 ;
      RECT 21.155 -22.21 21.245 -21.202 ;
      RECT 21.105 -21.975 21.245 -21.805 ;
      RECT 21.155 -20.788 21.245 -19.78 ;
      RECT 21.105 -20.185 21.245 -20.015 ;
      RECT 21.155 -18.98 21.245 -17.972 ;
      RECT 21.105 -18.745 21.245 -18.575 ;
      RECT 21.155 -17.558 21.245 -16.55 ;
      RECT 21.105 -16.955 21.245 -16.785 ;
      RECT 21.155 -15.75 21.245 -14.742 ;
      RECT 21.105 -15.515 21.245 -15.345 ;
      RECT 21.155 -14.328 21.245 -13.32 ;
      RECT 21.105 -13.725 21.245 -13.555 ;
      RECT 21.155 -12.52 21.245 -11.512 ;
      RECT 21.105 -12.285 21.245 -12.115 ;
      RECT 21.155 -11.098 21.245 -10.09 ;
      RECT 21.105 -10.495 21.245 -10.325 ;
      RECT 21.155 -9.29 21.245 -8.282 ;
      RECT 21.105 -9.055 21.245 -8.885 ;
      RECT 21.155 -7.868 21.245 -6.86 ;
      RECT 21.105 -7.265 21.245 -7.095 ;
      RECT 21.155 -6.06 21.245 -5.052 ;
      RECT 21.105 -5.825 21.245 -5.655 ;
      RECT 21.155 -4.638 21.245 -3.63 ;
      RECT 21.105 -4.035 21.245 -3.865 ;
      RECT 21.155 -2.83 21.245 -1.822 ;
      RECT 21.105 -2.595 21.245 -2.425 ;
      RECT 21.155 -1.408 21.245 -0.4 ;
      RECT 21.105 -0.805 21.245 -0.635 ;
      RECT 21.155 0.4 21.245 1.408 ;
      RECT 21.105 0.635 21.245 0.805 ;
      RECT 21.03 -114.685 21.205 -114.515 ;
      RECT 21.105 -114.895 21.205 -114.515 ;
      RECT 20.145 -113.555 20.245 -113.09 ;
      RECT 20.51 -113.555 20.61 -113.1 ;
      RECT 20.145 -113.555 20.99 -113.385 ;
      RECT 20.755 -101.538 20.845 -100.531 ;
      RECT 20.755 -101.225 20.895 -101.055 ;
      RECT 20.755 -99.729 20.845 -98.722 ;
      RECT 20.755 -99.205 20.895 -99.035 ;
      RECT 20.755 -98.308 20.845 -97.301 ;
      RECT 20.755 -97.995 20.895 -97.825 ;
      RECT 20.755 -96.499 20.845 -95.492 ;
      RECT 20.755 -95.975 20.895 -95.805 ;
      RECT 20.755 -95.078 20.845 -94.071 ;
      RECT 20.755 -94.765 20.895 -94.595 ;
      RECT 20.755 -93.269 20.845 -92.262 ;
      RECT 20.755 -92.745 20.895 -92.575 ;
      RECT 20.755 -91.848 20.845 -90.841 ;
      RECT 20.755 -91.535 20.895 -91.365 ;
      RECT 20.755 -90.039 20.845 -89.032 ;
      RECT 20.755 -89.515 20.895 -89.345 ;
      RECT 20.755 -88.618 20.845 -87.611 ;
      RECT 20.755 -88.305 20.895 -88.135 ;
      RECT 20.755 -86.809 20.845 -85.802 ;
      RECT 20.755 -86.285 20.895 -86.115 ;
      RECT 20.755 -85.388 20.845 -84.381 ;
      RECT 20.755 -85.075 20.895 -84.905 ;
      RECT 20.755 -83.579 20.845 -82.572 ;
      RECT 20.755 -83.055 20.895 -82.885 ;
      RECT 20.755 -82.158 20.845 -81.151 ;
      RECT 20.755 -81.845 20.895 -81.675 ;
      RECT 20.755 -80.349 20.845 -79.342 ;
      RECT 20.755 -79.825 20.895 -79.655 ;
      RECT 20.755 -78.928 20.845 -77.921 ;
      RECT 20.755 -78.615 20.895 -78.445 ;
      RECT 20.755 -77.119 20.845 -76.112 ;
      RECT 20.755 -76.595 20.895 -76.425 ;
      RECT 20.755 -75.698 20.845 -74.691 ;
      RECT 20.755 -75.385 20.895 -75.215 ;
      RECT 20.755 -73.889 20.845 -72.882 ;
      RECT 20.755 -73.365 20.895 -73.195 ;
      RECT 20.755 -72.468 20.845 -71.461 ;
      RECT 20.755 -72.155 20.895 -71.985 ;
      RECT 20.755 -70.659 20.845 -69.652 ;
      RECT 20.755 -70.135 20.895 -69.965 ;
      RECT 20.755 -69.238 20.845 -68.231 ;
      RECT 20.755 -68.925 20.895 -68.755 ;
      RECT 20.755 -67.429 20.845 -66.422 ;
      RECT 20.755 -66.905 20.895 -66.735 ;
      RECT 20.755 -66.008 20.845 -65.001 ;
      RECT 20.755 -65.695 20.895 -65.525 ;
      RECT 20.755 -64.199 20.845 -63.192 ;
      RECT 20.755 -63.675 20.895 -63.505 ;
      RECT 20.755 -62.778 20.845 -61.771 ;
      RECT 20.755 -62.465 20.895 -62.295 ;
      RECT 20.755 -60.969 20.845 -59.962 ;
      RECT 20.755 -60.445 20.895 -60.275 ;
      RECT 20.755 -59.548 20.845 -58.541 ;
      RECT 20.755 -59.235 20.895 -59.065 ;
      RECT 20.755 -57.739 20.845 -56.732 ;
      RECT 20.755 -57.215 20.895 -57.045 ;
      RECT 20.755 -56.318 20.845 -55.311 ;
      RECT 20.755 -56.005 20.895 -55.835 ;
      RECT 20.755 -54.509 20.845 -53.502 ;
      RECT 20.755 -53.985 20.895 -53.815 ;
      RECT 20.755 -53.088 20.845 -52.081 ;
      RECT 20.755 -52.775 20.895 -52.605 ;
      RECT 20.755 -51.279 20.845 -50.272 ;
      RECT 20.755 -50.755 20.895 -50.585 ;
      RECT 20.755 -49.858 20.845 -48.851 ;
      RECT 20.755 -49.545 20.895 -49.375 ;
      RECT 20.755 -48.049 20.845 -47.042 ;
      RECT 20.755 -47.525 20.895 -47.355 ;
      RECT 20.755 -46.628 20.845 -45.621 ;
      RECT 20.755 -46.315 20.895 -46.145 ;
      RECT 20.755 -44.819 20.845 -43.812 ;
      RECT 20.755 -44.295 20.895 -44.125 ;
      RECT 20.755 -43.398 20.845 -42.391 ;
      RECT 20.755 -43.085 20.895 -42.915 ;
      RECT 20.755 -41.589 20.845 -40.582 ;
      RECT 20.755 -41.065 20.895 -40.895 ;
      RECT 20.755 -40.168 20.845 -39.161 ;
      RECT 20.755 -39.855 20.895 -39.685 ;
      RECT 20.755 -38.359 20.845 -37.352 ;
      RECT 20.755 -37.835 20.895 -37.665 ;
      RECT 20.755 -36.938 20.845 -35.931 ;
      RECT 20.755 -36.625 20.895 -36.455 ;
      RECT 20.755 -35.129 20.845 -34.122 ;
      RECT 20.755 -34.605 20.895 -34.435 ;
      RECT 20.755 -33.708 20.845 -32.701 ;
      RECT 20.755 -33.395 20.895 -33.225 ;
      RECT 20.755 -31.899 20.845 -30.892 ;
      RECT 20.755 -31.375 20.895 -31.205 ;
      RECT 20.755 -30.478 20.845 -29.471 ;
      RECT 20.755 -30.165 20.895 -29.995 ;
      RECT 20.755 -28.669 20.845 -27.662 ;
      RECT 20.755 -28.145 20.895 -27.975 ;
      RECT 20.755 -27.248 20.845 -26.241 ;
      RECT 20.755 -26.935 20.895 -26.765 ;
      RECT 20.755 -25.439 20.845 -24.432 ;
      RECT 20.755 -24.915 20.895 -24.745 ;
      RECT 20.755 -24.018 20.845 -23.011 ;
      RECT 20.755 -23.705 20.895 -23.535 ;
      RECT 20.755 -22.209 20.845 -21.202 ;
      RECT 20.755 -21.685 20.895 -21.515 ;
      RECT 20.755 -20.788 20.845 -19.781 ;
      RECT 20.755 -20.475 20.895 -20.305 ;
      RECT 20.755 -18.979 20.845 -17.972 ;
      RECT 20.755 -18.455 20.895 -18.285 ;
      RECT 20.755 -17.558 20.845 -16.551 ;
      RECT 20.755 -17.245 20.895 -17.075 ;
      RECT 20.755 -15.749 20.845 -14.742 ;
      RECT 20.755 -15.225 20.895 -15.055 ;
      RECT 20.755 -14.328 20.845 -13.321 ;
      RECT 20.755 -14.015 20.895 -13.845 ;
      RECT 20.755 -12.519 20.845 -11.512 ;
      RECT 20.755 -11.995 20.895 -11.825 ;
      RECT 20.755 -11.098 20.845 -10.091 ;
      RECT 20.755 -10.785 20.895 -10.615 ;
      RECT 20.755 -9.289 20.845 -8.282 ;
      RECT 20.755 -8.765 20.895 -8.595 ;
      RECT 20.755 -7.868 20.845 -6.861 ;
      RECT 20.755 -7.555 20.895 -7.385 ;
      RECT 20.755 -6.059 20.845 -5.052 ;
      RECT 20.755 -5.535 20.895 -5.365 ;
      RECT 20.755 -4.638 20.845 -3.631 ;
      RECT 20.755 -4.325 20.895 -4.155 ;
      RECT 20.755 -2.829 20.845 -1.822 ;
      RECT 20.755 -2.305 20.895 -2.135 ;
      RECT 20.755 -1.408 20.845 -0.401 ;
      RECT 20.755 -1.095 20.895 -0.925 ;
      RECT 20.755 0.401 20.845 1.408 ;
      RECT 20.755 0.925 20.895 1.095 ;
      RECT 20.44 -114.685 20.61 -114.515 ;
      RECT 20.51 -114.895 20.61 -114.515 ;
      RECT 19.955 -101.538 20.045 -100.53 ;
      RECT 19.905 -100.935 20.045 -100.765 ;
      RECT 19.955 -99.73 20.045 -98.722 ;
      RECT 19.905 -99.495 20.045 -99.325 ;
      RECT 19.955 -98.308 20.045 -97.3 ;
      RECT 19.905 -97.705 20.045 -97.535 ;
      RECT 19.955 -96.5 20.045 -95.492 ;
      RECT 19.905 -96.265 20.045 -96.095 ;
      RECT 19.955 -95.078 20.045 -94.07 ;
      RECT 19.905 -94.475 20.045 -94.305 ;
      RECT 19.955 -93.27 20.045 -92.262 ;
      RECT 19.905 -93.035 20.045 -92.865 ;
      RECT 19.955 -91.848 20.045 -90.84 ;
      RECT 19.905 -91.245 20.045 -91.075 ;
      RECT 19.955 -90.04 20.045 -89.032 ;
      RECT 19.905 -89.805 20.045 -89.635 ;
      RECT 19.955 -88.618 20.045 -87.61 ;
      RECT 19.905 -88.015 20.045 -87.845 ;
      RECT 19.955 -86.81 20.045 -85.802 ;
      RECT 19.905 -86.575 20.045 -86.405 ;
      RECT 19.955 -85.388 20.045 -84.38 ;
      RECT 19.905 -84.785 20.045 -84.615 ;
      RECT 19.955 -83.58 20.045 -82.572 ;
      RECT 19.905 -83.345 20.045 -83.175 ;
      RECT 19.955 -82.158 20.045 -81.15 ;
      RECT 19.905 -81.555 20.045 -81.385 ;
      RECT 19.955 -80.35 20.045 -79.342 ;
      RECT 19.905 -80.115 20.045 -79.945 ;
      RECT 19.955 -78.928 20.045 -77.92 ;
      RECT 19.905 -78.325 20.045 -78.155 ;
      RECT 19.955 -77.12 20.045 -76.112 ;
      RECT 19.905 -76.885 20.045 -76.715 ;
      RECT 19.955 -75.698 20.045 -74.69 ;
      RECT 19.905 -75.095 20.045 -74.925 ;
      RECT 19.955 -73.89 20.045 -72.882 ;
      RECT 19.905 -73.655 20.045 -73.485 ;
      RECT 19.955 -72.468 20.045 -71.46 ;
      RECT 19.905 -71.865 20.045 -71.695 ;
      RECT 19.955 -70.66 20.045 -69.652 ;
      RECT 19.905 -70.425 20.045 -70.255 ;
      RECT 19.955 -69.238 20.045 -68.23 ;
      RECT 19.905 -68.635 20.045 -68.465 ;
      RECT 19.955 -67.43 20.045 -66.422 ;
      RECT 19.905 -67.195 20.045 -67.025 ;
      RECT 19.955 -66.008 20.045 -65 ;
      RECT 19.905 -65.405 20.045 -65.235 ;
      RECT 19.955 -64.2 20.045 -63.192 ;
      RECT 19.905 -63.965 20.045 -63.795 ;
      RECT 19.955 -62.778 20.045 -61.77 ;
      RECT 19.905 -62.175 20.045 -62.005 ;
      RECT 19.955 -60.97 20.045 -59.962 ;
      RECT 19.905 -60.735 20.045 -60.565 ;
      RECT 19.955 -59.548 20.045 -58.54 ;
      RECT 19.905 -58.945 20.045 -58.775 ;
      RECT 19.955 -57.74 20.045 -56.732 ;
      RECT 19.905 -57.505 20.045 -57.335 ;
      RECT 19.955 -56.318 20.045 -55.31 ;
      RECT 19.905 -55.715 20.045 -55.545 ;
      RECT 19.955 -54.51 20.045 -53.502 ;
      RECT 19.905 -54.275 20.045 -54.105 ;
      RECT 19.955 -53.088 20.045 -52.08 ;
      RECT 19.905 -52.485 20.045 -52.315 ;
      RECT 19.955 -51.28 20.045 -50.272 ;
      RECT 19.905 -51.045 20.045 -50.875 ;
      RECT 19.955 -49.858 20.045 -48.85 ;
      RECT 19.905 -49.255 20.045 -49.085 ;
      RECT 19.955 -48.05 20.045 -47.042 ;
      RECT 19.905 -47.815 20.045 -47.645 ;
      RECT 19.955 -46.628 20.045 -45.62 ;
      RECT 19.905 -46.025 20.045 -45.855 ;
      RECT 19.955 -44.82 20.045 -43.812 ;
      RECT 19.905 -44.585 20.045 -44.415 ;
      RECT 19.955 -43.398 20.045 -42.39 ;
      RECT 19.905 -42.795 20.045 -42.625 ;
      RECT 19.955 -41.59 20.045 -40.582 ;
      RECT 19.905 -41.355 20.045 -41.185 ;
      RECT 19.955 -40.168 20.045 -39.16 ;
      RECT 19.905 -39.565 20.045 -39.395 ;
      RECT 19.955 -38.36 20.045 -37.352 ;
      RECT 19.905 -38.125 20.045 -37.955 ;
      RECT 19.955 -36.938 20.045 -35.93 ;
      RECT 19.905 -36.335 20.045 -36.165 ;
      RECT 19.955 -35.13 20.045 -34.122 ;
      RECT 19.905 -34.895 20.045 -34.725 ;
      RECT 19.955 -33.708 20.045 -32.7 ;
      RECT 19.905 -33.105 20.045 -32.935 ;
      RECT 19.955 -31.9 20.045 -30.892 ;
      RECT 19.905 -31.665 20.045 -31.495 ;
      RECT 19.955 -30.478 20.045 -29.47 ;
      RECT 19.905 -29.875 20.045 -29.705 ;
      RECT 19.955 -28.67 20.045 -27.662 ;
      RECT 19.905 -28.435 20.045 -28.265 ;
      RECT 19.955 -27.248 20.045 -26.24 ;
      RECT 19.905 -26.645 20.045 -26.475 ;
      RECT 19.955 -25.44 20.045 -24.432 ;
      RECT 19.905 -25.205 20.045 -25.035 ;
      RECT 19.955 -24.018 20.045 -23.01 ;
      RECT 19.905 -23.415 20.045 -23.245 ;
      RECT 19.955 -22.21 20.045 -21.202 ;
      RECT 19.905 -21.975 20.045 -21.805 ;
      RECT 19.955 -20.788 20.045 -19.78 ;
      RECT 19.905 -20.185 20.045 -20.015 ;
      RECT 19.955 -18.98 20.045 -17.972 ;
      RECT 19.905 -18.745 20.045 -18.575 ;
      RECT 19.955 -17.558 20.045 -16.55 ;
      RECT 19.905 -16.955 20.045 -16.785 ;
      RECT 19.955 -15.75 20.045 -14.742 ;
      RECT 19.905 -15.515 20.045 -15.345 ;
      RECT 19.955 -14.328 20.045 -13.32 ;
      RECT 19.905 -13.725 20.045 -13.555 ;
      RECT 19.955 -12.52 20.045 -11.512 ;
      RECT 19.905 -12.285 20.045 -12.115 ;
      RECT 19.955 -11.098 20.045 -10.09 ;
      RECT 19.905 -10.495 20.045 -10.325 ;
      RECT 19.955 -9.29 20.045 -8.282 ;
      RECT 19.905 -9.055 20.045 -8.885 ;
      RECT 19.955 -7.868 20.045 -6.86 ;
      RECT 19.905 -7.265 20.045 -7.095 ;
      RECT 19.955 -6.06 20.045 -5.052 ;
      RECT 19.905 -5.825 20.045 -5.655 ;
      RECT 19.955 -4.638 20.045 -3.63 ;
      RECT 19.905 -4.035 20.045 -3.865 ;
      RECT 19.955 -2.83 20.045 -1.822 ;
      RECT 19.905 -2.595 20.045 -2.425 ;
      RECT 19.955 -1.408 20.045 -0.4 ;
      RECT 19.905 -0.805 20.045 -0.635 ;
      RECT 19.955 0.4 20.045 1.408 ;
      RECT 19.905 0.635 20.045 0.805 ;
      RECT 19.555 -101.538 19.645 -100.531 ;
      RECT 19.555 -101.225 19.695 -101.055 ;
      RECT 19.555 -99.729 19.645 -98.722 ;
      RECT 19.555 -99.205 19.695 -99.035 ;
      RECT 19.555 -98.308 19.645 -97.301 ;
      RECT 19.555 -97.995 19.695 -97.825 ;
      RECT 19.555 -96.499 19.645 -95.492 ;
      RECT 19.555 -95.975 19.695 -95.805 ;
      RECT 19.555 -95.078 19.645 -94.071 ;
      RECT 19.555 -94.765 19.695 -94.595 ;
      RECT 19.555 -93.269 19.645 -92.262 ;
      RECT 19.555 -92.745 19.695 -92.575 ;
      RECT 19.555 -91.848 19.645 -90.841 ;
      RECT 19.555 -91.535 19.695 -91.365 ;
      RECT 19.555 -90.039 19.645 -89.032 ;
      RECT 19.555 -89.515 19.695 -89.345 ;
      RECT 19.555 -88.618 19.645 -87.611 ;
      RECT 19.555 -88.305 19.695 -88.135 ;
      RECT 19.555 -86.809 19.645 -85.802 ;
      RECT 19.555 -86.285 19.695 -86.115 ;
      RECT 19.555 -85.388 19.645 -84.381 ;
      RECT 19.555 -85.075 19.695 -84.905 ;
      RECT 19.555 -83.579 19.645 -82.572 ;
      RECT 19.555 -83.055 19.695 -82.885 ;
      RECT 19.555 -82.158 19.645 -81.151 ;
      RECT 19.555 -81.845 19.695 -81.675 ;
      RECT 19.555 -80.349 19.645 -79.342 ;
      RECT 19.555 -79.825 19.695 -79.655 ;
      RECT 19.555 -78.928 19.645 -77.921 ;
      RECT 19.555 -78.615 19.695 -78.445 ;
      RECT 19.555 -77.119 19.645 -76.112 ;
      RECT 19.555 -76.595 19.695 -76.425 ;
      RECT 19.555 -75.698 19.645 -74.691 ;
      RECT 19.555 -75.385 19.695 -75.215 ;
      RECT 19.555 -73.889 19.645 -72.882 ;
      RECT 19.555 -73.365 19.695 -73.195 ;
      RECT 19.555 -72.468 19.645 -71.461 ;
      RECT 19.555 -72.155 19.695 -71.985 ;
      RECT 19.555 -70.659 19.645 -69.652 ;
      RECT 19.555 -70.135 19.695 -69.965 ;
      RECT 19.555 -69.238 19.645 -68.231 ;
      RECT 19.555 -68.925 19.695 -68.755 ;
      RECT 19.555 -67.429 19.645 -66.422 ;
      RECT 19.555 -66.905 19.695 -66.735 ;
      RECT 19.555 -66.008 19.645 -65.001 ;
      RECT 19.555 -65.695 19.695 -65.525 ;
      RECT 19.555 -64.199 19.645 -63.192 ;
      RECT 19.555 -63.675 19.695 -63.505 ;
      RECT 19.555 -62.778 19.645 -61.771 ;
      RECT 19.555 -62.465 19.695 -62.295 ;
      RECT 19.555 -60.969 19.645 -59.962 ;
      RECT 19.555 -60.445 19.695 -60.275 ;
      RECT 19.555 -59.548 19.645 -58.541 ;
      RECT 19.555 -59.235 19.695 -59.065 ;
      RECT 19.555 -57.739 19.645 -56.732 ;
      RECT 19.555 -57.215 19.695 -57.045 ;
      RECT 19.555 -56.318 19.645 -55.311 ;
      RECT 19.555 -56.005 19.695 -55.835 ;
      RECT 19.555 -54.509 19.645 -53.502 ;
      RECT 19.555 -53.985 19.695 -53.815 ;
      RECT 19.555 -53.088 19.645 -52.081 ;
      RECT 19.555 -52.775 19.695 -52.605 ;
      RECT 19.555 -51.279 19.645 -50.272 ;
      RECT 19.555 -50.755 19.695 -50.585 ;
      RECT 19.555 -49.858 19.645 -48.851 ;
      RECT 19.555 -49.545 19.695 -49.375 ;
      RECT 19.555 -48.049 19.645 -47.042 ;
      RECT 19.555 -47.525 19.695 -47.355 ;
      RECT 19.555 -46.628 19.645 -45.621 ;
      RECT 19.555 -46.315 19.695 -46.145 ;
      RECT 19.555 -44.819 19.645 -43.812 ;
      RECT 19.555 -44.295 19.695 -44.125 ;
      RECT 19.555 -43.398 19.645 -42.391 ;
      RECT 19.555 -43.085 19.695 -42.915 ;
      RECT 19.555 -41.589 19.645 -40.582 ;
      RECT 19.555 -41.065 19.695 -40.895 ;
      RECT 19.555 -40.168 19.645 -39.161 ;
      RECT 19.555 -39.855 19.695 -39.685 ;
      RECT 19.555 -38.359 19.645 -37.352 ;
      RECT 19.555 -37.835 19.695 -37.665 ;
      RECT 19.555 -36.938 19.645 -35.931 ;
      RECT 19.555 -36.625 19.695 -36.455 ;
      RECT 19.555 -35.129 19.645 -34.122 ;
      RECT 19.555 -34.605 19.695 -34.435 ;
      RECT 19.555 -33.708 19.645 -32.701 ;
      RECT 19.555 -33.395 19.695 -33.225 ;
      RECT 19.555 -31.899 19.645 -30.892 ;
      RECT 19.555 -31.375 19.695 -31.205 ;
      RECT 19.555 -30.478 19.645 -29.471 ;
      RECT 19.555 -30.165 19.695 -29.995 ;
      RECT 19.555 -28.669 19.645 -27.662 ;
      RECT 19.555 -28.145 19.695 -27.975 ;
      RECT 19.555 -27.248 19.645 -26.241 ;
      RECT 19.555 -26.935 19.695 -26.765 ;
      RECT 19.555 -25.439 19.645 -24.432 ;
      RECT 19.555 -24.915 19.695 -24.745 ;
      RECT 19.555 -24.018 19.645 -23.011 ;
      RECT 19.555 -23.705 19.695 -23.535 ;
      RECT 19.555 -22.209 19.645 -21.202 ;
      RECT 19.555 -21.685 19.695 -21.515 ;
      RECT 19.555 -20.788 19.645 -19.781 ;
      RECT 19.555 -20.475 19.695 -20.305 ;
      RECT 19.555 -18.979 19.645 -17.972 ;
      RECT 19.555 -18.455 19.695 -18.285 ;
      RECT 19.555 -17.558 19.645 -16.551 ;
      RECT 19.555 -17.245 19.695 -17.075 ;
      RECT 19.555 -15.749 19.645 -14.742 ;
      RECT 19.555 -15.225 19.695 -15.055 ;
      RECT 19.555 -14.328 19.645 -13.321 ;
      RECT 19.555 -14.015 19.695 -13.845 ;
      RECT 19.555 -12.519 19.645 -11.512 ;
      RECT 19.555 -11.995 19.695 -11.825 ;
      RECT 19.555 -11.098 19.645 -10.091 ;
      RECT 19.555 -10.785 19.695 -10.615 ;
      RECT 19.555 -9.289 19.645 -8.282 ;
      RECT 19.555 -8.765 19.695 -8.595 ;
      RECT 19.555 -7.868 19.645 -6.861 ;
      RECT 19.555 -7.555 19.695 -7.385 ;
      RECT 19.555 -6.059 19.645 -5.052 ;
      RECT 19.555 -5.535 19.695 -5.365 ;
      RECT 19.555 -4.638 19.645 -3.631 ;
      RECT 19.555 -4.325 19.695 -4.155 ;
      RECT 19.555 -2.829 19.645 -1.822 ;
      RECT 19.555 -2.305 19.695 -2.135 ;
      RECT 19.555 -1.408 19.645 -0.401 ;
      RECT 19.555 -1.095 19.695 -0.925 ;
      RECT 19.555 0.401 19.645 1.408 ;
      RECT 19.555 0.925 19.695 1.095 ;
      RECT 15.385 -108.935 19.165 -108.815 ;
      RECT 16.705 -109.475 16.805 -108.815 ;
      RECT 16.145 -109.475 16.245 -108.815 ;
      RECT 15.585 -109.475 15.685 -108.815 ;
      RECT 18.755 -101.538 18.845 -100.53 ;
      RECT 18.705 -100.935 18.845 -100.765 ;
      RECT 18.755 -99.73 18.845 -98.722 ;
      RECT 18.705 -99.495 18.845 -99.325 ;
      RECT 18.755 -98.308 18.845 -97.3 ;
      RECT 18.705 -97.705 18.845 -97.535 ;
      RECT 18.755 -96.5 18.845 -95.492 ;
      RECT 18.705 -96.265 18.845 -96.095 ;
      RECT 18.755 -95.078 18.845 -94.07 ;
      RECT 18.705 -94.475 18.845 -94.305 ;
      RECT 18.755 -93.27 18.845 -92.262 ;
      RECT 18.705 -93.035 18.845 -92.865 ;
      RECT 18.755 -91.848 18.845 -90.84 ;
      RECT 18.705 -91.245 18.845 -91.075 ;
      RECT 18.755 -90.04 18.845 -89.032 ;
      RECT 18.705 -89.805 18.845 -89.635 ;
      RECT 18.755 -88.618 18.845 -87.61 ;
      RECT 18.705 -88.015 18.845 -87.845 ;
      RECT 18.755 -86.81 18.845 -85.802 ;
      RECT 18.705 -86.575 18.845 -86.405 ;
      RECT 18.755 -85.388 18.845 -84.38 ;
      RECT 18.705 -84.785 18.845 -84.615 ;
      RECT 18.755 -83.58 18.845 -82.572 ;
      RECT 18.705 -83.345 18.845 -83.175 ;
      RECT 18.755 -82.158 18.845 -81.15 ;
      RECT 18.705 -81.555 18.845 -81.385 ;
      RECT 18.755 -80.35 18.845 -79.342 ;
      RECT 18.705 -80.115 18.845 -79.945 ;
      RECT 18.755 -78.928 18.845 -77.92 ;
      RECT 18.705 -78.325 18.845 -78.155 ;
      RECT 18.755 -77.12 18.845 -76.112 ;
      RECT 18.705 -76.885 18.845 -76.715 ;
      RECT 18.755 -75.698 18.845 -74.69 ;
      RECT 18.705 -75.095 18.845 -74.925 ;
      RECT 18.755 -73.89 18.845 -72.882 ;
      RECT 18.705 -73.655 18.845 -73.485 ;
      RECT 18.755 -72.468 18.845 -71.46 ;
      RECT 18.705 -71.865 18.845 -71.695 ;
      RECT 18.755 -70.66 18.845 -69.652 ;
      RECT 18.705 -70.425 18.845 -70.255 ;
      RECT 18.755 -69.238 18.845 -68.23 ;
      RECT 18.705 -68.635 18.845 -68.465 ;
      RECT 18.755 -67.43 18.845 -66.422 ;
      RECT 18.705 -67.195 18.845 -67.025 ;
      RECT 18.755 -66.008 18.845 -65 ;
      RECT 18.705 -65.405 18.845 -65.235 ;
      RECT 18.755 -64.2 18.845 -63.192 ;
      RECT 18.705 -63.965 18.845 -63.795 ;
      RECT 18.755 -62.778 18.845 -61.77 ;
      RECT 18.705 -62.175 18.845 -62.005 ;
      RECT 18.755 -60.97 18.845 -59.962 ;
      RECT 18.705 -60.735 18.845 -60.565 ;
      RECT 18.755 -59.548 18.845 -58.54 ;
      RECT 18.705 -58.945 18.845 -58.775 ;
      RECT 18.755 -57.74 18.845 -56.732 ;
      RECT 18.705 -57.505 18.845 -57.335 ;
      RECT 18.755 -56.318 18.845 -55.31 ;
      RECT 18.705 -55.715 18.845 -55.545 ;
      RECT 18.755 -54.51 18.845 -53.502 ;
      RECT 18.705 -54.275 18.845 -54.105 ;
      RECT 18.755 -53.088 18.845 -52.08 ;
      RECT 18.705 -52.485 18.845 -52.315 ;
      RECT 18.755 -51.28 18.845 -50.272 ;
      RECT 18.705 -51.045 18.845 -50.875 ;
      RECT 18.755 -49.858 18.845 -48.85 ;
      RECT 18.705 -49.255 18.845 -49.085 ;
      RECT 18.755 -48.05 18.845 -47.042 ;
      RECT 18.705 -47.815 18.845 -47.645 ;
      RECT 18.755 -46.628 18.845 -45.62 ;
      RECT 18.705 -46.025 18.845 -45.855 ;
      RECT 18.755 -44.82 18.845 -43.812 ;
      RECT 18.705 -44.585 18.845 -44.415 ;
      RECT 18.755 -43.398 18.845 -42.39 ;
      RECT 18.705 -42.795 18.845 -42.625 ;
      RECT 18.755 -41.59 18.845 -40.582 ;
      RECT 18.705 -41.355 18.845 -41.185 ;
      RECT 18.755 -40.168 18.845 -39.16 ;
      RECT 18.705 -39.565 18.845 -39.395 ;
      RECT 18.755 -38.36 18.845 -37.352 ;
      RECT 18.705 -38.125 18.845 -37.955 ;
      RECT 18.755 -36.938 18.845 -35.93 ;
      RECT 18.705 -36.335 18.845 -36.165 ;
      RECT 18.755 -35.13 18.845 -34.122 ;
      RECT 18.705 -34.895 18.845 -34.725 ;
      RECT 18.755 -33.708 18.845 -32.7 ;
      RECT 18.705 -33.105 18.845 -32.935 ;
      RECT 18.755 -31.9 18.845 -30.892 ;
      RECT 18.705 -31.665 18.845 -31.495 ;
      RECT 18.755 -30.478 18.845 -29.47 ;
      RECT 18.705 -29.875 18.845 -29.705 ;
      RECT 18.755 -28.67 18.845 -27.662 ;
      RECT 18.705 -28.435 18.845 -28.265 ;
      RECT 18.755 -27.248 18.845 -26.24 ;
      RECT 18.705 -26.645 18.845 -26.475 ;
      RECT 18.755 -25.44 18.845 -24.432 ;
      RECT 18.705 -25.205 18.845 -25.035 ;
      RECT 18.755 -24.018 18.845 -23.01 ;
      RECT 18.705 -23.415 18.845 -23.245 ;
      RECT 18.755 -22.21 18.845 -21.202 ;
      RECT 18.705 -21.975 18.845 -21.805 ;
      RECT 18.755 -20.788 18.845 -19.78 ;
      RECT 18.705 -20.185 18.845 -20.015 ;
      RECT 18.755 -18.98 18.845 -17.972 ;
      RECT 18.705 -18.745 18.845 -18.575 ;
      RECT 18.755 -17.558 18.845 -16.55 ;
      RECT 18.705 -16.955 18.845 -16.785 ;
      RECT 18.755 -15.75 18.845 -14.742 ;
      RECT 18.705 -15.515 18.845 -15.345 ;
      RECT 18.755 -14.328 18.845 -13.32 ;
      RECT 18.705 -13.725 18.845 -13.555 ;
      RECT 18.755 -12.52 18.845 -11.512 ;
      RECT 18.705 -12.285 18.845 -12.115 ;
      RECT 18.755 -11.098 18.845 -10.09 ;
      RECT 18.705 -10.495 18.845 -10.325 ;
      RECT 18.755 -9.29 18.845 -8.282 ;
      RECT 18.705 -9.055 18.845 -8.885 ;
      RECT 18.755 -7.868 18.845 -6.86 ;
      RECT 18.705 -7.265 18.845 -7.095 ;
      RECT 18.755 -6.06 18.845 -5.052 ;
      RECT 18.705 -5.825 18.845 -5.655 ;
      RECT 18.755 -4.638 18.845 -3.63 ;
      RECT 18.705 -4.035 18.845 -3.865 ;
      RECT 18.755 -2.83 18.845 -1.822 ;
      RECT 18.705 -2.595 18.845 -2.425 ;
      RECT 18.755 -1.408 18.845 -0.4 ;
      RECT 18.705 -0.805 18.845 -0.635 ;
      RECT 18.755 0.4 18.845 1.408 ;
      RECT 18.705 0.635 18.845 0.805 ;
      RECT 17.325 -111.685 18.805 -111.585 ;
      RECT 17.325 -112.195 17.425 -111.585 ;
      RECT 17.545 -109.15 18.805 -109.05 ;
      RECT 18.705 -109.475 18.805 -109.05 ;
      RECT 18.145 -109.475 18.245 -109.05 ;
      RECT 17.585 -109.475 17.685 -109.05 ;
      RECT 18.355 -101.538 18.445 -100.531 ;
      RECT 18.355 -101.225 18.495 -101.055 ;
      RECT 18.355 -99.729 18.445 -98.722 ;
      RECT 18.355 -99.205 18.495 -99.035 ;
      RECT 18.355 -98.308 18.445 -97.301 ;
      RECT 18.355 -97.995 18.495 -97.825 ;
      RECT 18.355 -96.499 18.445 -95.492 ;
      RECT 18.355 -95.975 18.495 -95.805 ;
      RECT 18.355 -95.078 18.445 -94.071 ;
      RECT 18.355 -94.765 18.495 -94.595 ;
      RECT 18.355 -93.269 18.445 -92.262 ;
      RECT 18.355 -92.745 18.495 -92.575 ;
      RECT 18.355 -91.848 18.445 -90.841 ;
      RECT 18.355 -91.535 18.495 -91.365 ;
      RECT 18.355 -90.039 18.445 -89.032 ;
      RECT 18.355 -89.515 18.495 -89.345 ;
      RECT 18.355 -88.618 18.445 -87.611 ;
      RECT 18.355 -88.305 18.495 -88.135 ;
      RECT 18.355 -86.809 18.445 -85.802 ;
      RECT 18.355 -86.285 18.495 -86.115 ;
      RECT 18.355 -85.388 18.445 -84.381 ;
      RECT 18.355 -85.075 18.495 -84.905 ;
      RECT 18.355 -83.579 18.445 -82.572 ;
      RECT 18.355 -83.055 18.495 -82.885 ;
      RECT 18.355 -82.158 18.445 -81.151 ;
      RECT 18.355 -81.845 18.495 -81.675 ;
      RECT 18.355 -80.349 18.445 -79.342 ;
      RECT 18.355 -79.825 18.495 -79.655 ;
      RECT 18.355 -78.928 18.445 -77.921 ;
      RECT 18.355 -78.615 18.495 -78.445 ;
      RECT 18.355 -77.119 18.445 -76.112 ;
      RECT 18.355 -76.595 18.495 -76.425 ;
      RECT 18.355 -75.698 18.445 -74.691 ;
      RECT 18.355 -75.385 18.495 -75.215 ;
      RECT 18.355 -73.889 18.445 -72.882 ;
      RECT 18.355 -73.365 18.495 -73.195 ;
      RECT 18.355 -72.468 18.445 -71.461 ;
      RECT 18.355 -72.155 18.495 -71.985 ;
      RECT 18.355 -70.659 18.445 -69.652 ;
      RECT 18.355 -70.135 18.495 -69.965 ;
      RECT 18.355 -69.238 18.445 -68.231 ;
      RECT 18.355 -68.925 18.495 -68.755 ;
      RECT 18.355 -67.429 18.445 -66.422 ;
      RECT 18.355 -66.905 18.495 -66.735 ;
      RECT 18.355 -66.008 18.445 -65.001 ;
      RECT 18.355 -65.695 18.495 -65.525 ;
      RECT 18.355 -64.199 18.445 -63.192 ;
      RECT 18.355 -63.675 18.495 -63.505 ;
      RECT 18.355 -62.778 18.445 -61.771 ;
      RECT 18.355 -62.465 18.495 -62.295 ;
      RECT 18.355 -60.969 18.445 -59.962 ;
      RECT 18.355 -60.445 18.495 -60.275 ;
      RECT 18.355 -59.548 18.445 -58.541 ;
      RECT 18.355 -59.235 18.495 -59.065 ;
      RECT 18.355 -57.739 18.445 -56.732 ;
      RECT 18.355 -57.215 18.495 -57.045 ;
      RECT 18.355 -56.318 18.445 -55.311 ;
      RECT 18.355 -56.005 18.495 -55.835 ;
      RECT 18.355 -54.509 18.445 -53.502 ;
      RECT 18.355 -53.985 18.495 -53.815 ;
      RECT 18.355 -53.088 18.445 -52.081 ;
      RECT 18.355 -52.775 18.495 -52.605 ;
      RECT 18.355 -51.279 18.445 -50.272 ;
      RECT 18.355 -50.755 18.495 -50.585 ;
      RECT 18.355 -49.858 18.445 -48.851 ;
      RECT 18.355 -49.545 18.495 -49.375 ;
      RECT 18.355 -48.049 18.445 -47.042 ;
      RECT 18.355 -47.525 18.495 -47.355 ;
      RECT 18.355 -46.628 18.445 -45.621 ;
      RECT 18.355 -46.315 18.495 -46.145 ;
      RECT 18.355 -44.819 18.445 -43.812 ;
      RECT 18.355 -44.295 18.495 -44.125 ;
      RECT 18.355 -43.398 18.445 -42.391 ;
      RECT 18.355 -43.085 18.495 -42.915 ;
      RECT 18.355 -41.589 18.445 -40.582 ;
      RECT 18.355 -41.065 18.495 -40.895 ;
      RECT 18.355 -40.168 18.445 -39.161 ;
      RECT 18.355 -39.855 18.495 -39.685 ;
      RECT 18.355 -38.359 18.445 -37.352 ;
      RECT 18.355 -37.835 18.495 -37.665 ;
      RECT 18.355 -36.938 18.445 -35.931 ;
      RECT 18.355 -36.625 18.495 -36.455 ;
      RECT 18.355 -35.129 18.445 -34.122 ;
      RECT 18.355 -34.605 18.495 -34.435 ;
      RECT 18.355 -33.708 18.445 -32.701 ;
      RECT 18.355 -33.395 18.495 -33.225 ;
      RECT 18.355 -31.899 18.445 -30.892 ;
      RECT 18.355 -31.375 18.495 -31.205 ;
      RECT 18.355 -30.478 18.445 -29.471 ;
      RECT 18.355 -30.165 18.495 -29.995 ;
      RECT 18.355 -28.669 18.445 -27.662 ;
      RECT 18.355 -28.145 18.495 -27.975 ;
      RECT 18.355 -27.248 18.445 -26.241 ;
      RECT 18.355 -26.935 18.495 -26.765 ;
      RECT 18.355 -25.439 18.445 -24.432 ;
      RECT 18.355 -24.915 18.495 -24.745 ;
      RECT 18.355 -24.018 18.445 -23.011 ;
      RECT 18.355 -23.705 18.495 -23.535 ;
      RECT 18.355 -22.209 18.445 -21.202 ;
      RECT 18.355 -21.685 18.495 -21.515 ;
      RECT 18.355 -20.788 18.445 -19.781 ;
      RECT 18.355 -20.475 18.495 -20.305 ;
      RECT 18.355 -18.979 18.445 -17.972 ;
      RECT 18.355 -18.455 18.495 -18.285 ;
      RECT 18.355 -17.558 18.445 -16.551 ;
      RECT 18.355 -17.245 18.495 -17.075 ;
      RECT 18.355 -15.749 18.445 -14.742 ;
      RECT 18.355 -15.225 18.495 -15.055 ;
      RECT 18.355 -14.328 18.445 -13.321 ;
      RECT 18.355 -14.015 18.495 -13.845 ;
      RECT 18.355 -12.519 18.445 -11.512 ;
      RECT 18.355 -11.995 18.495 -11.825 ;
      RECT 18.355 -11.098 18.445 -10.091 ;
      RECT 18.355 -10.785 18.495 -10.615 ;
      RECT 18.355 -9.289 18.445 -8.282 ;
      RECT 18.355 -8.765 18.495 -8.595 ;
      RECT 18.355 -7.868 18.445 -6.861 ;
      RECT 18.355 -7.555 18.495 -7.385 ;
      RECT 18.355 -6.059 18.445 -5.052 ;
      RECT 18.355 -5.535 18.495 -5.365 ;
      RECT 18.355 -4.638 18.445 -3.631 ;
      RECT 18.355 -4.325 18.495 -4.155 ;
      RECT 18.355 -2.829 18.445 -1.822 ;
      RECT 18.355 -2.305 18.495 -2.135 ;
      RECT 18.355 -1.408 18.445 -0.401 ;
      RECT 18.355 -1.095 18.495 -0.925 ;
      RECT 18.355 0.401 18.445 1.408 ;
      RECT 18.355 0.925 18.495 1.095 ;
      RECT 17.685 -111.495 17.855 -111.385 ;
      RECT 14.535 -111.495 17.855 -111.395 ;
      RECT 17.555 -101.538 17.645 -100.53 ;
      RECT 17.505 -100.935 17.645 -100.765 ;
      RECT 17.555 -99.73 17.645 -98.722 ;
      RECT 17.505 -99.495 17.645 -99.325 ;
      RECT 17.555 -98.308 17.645 -97.3 ;
      RECT 17.505 -97.705 17.645 -97.535 ;
      RECT 17.555 -96.5 17.645 -95.492 ;
      RECT 17.505 -96.265 17.645 -96.095 ;
      RECT 17.555 -95.078 17.645 -94.07 ;
      RECT 17.505 -94.475 17.645 -94.305 ;
      RECT 17.555 -93.27 17.645 -92.262 ;
      RECT 17.505 -93.035 17.645 -92.865 ;
      RECT 17.555 -91.848 17.645 -90.84 ;
      RECT 17.505 -91.245 17.645 -91.075 ;
      RECT 17.555 -90.04 17.645 -89.032 ;
      RECT 17.505 -89.805 17.645 -89.635 ;
      RECT 17.555 -88.618 17.645 -87.61 ;
      RECT 17.505 -88.015 17.645 -87.845 ;
      RECT 17.555 -86.81 17.645 -85.802 ;
      RECT 17.505 -86.575 17.645 -86.405 ;
      RECT 17.555 -85.388 17.645 -84.38 ;
      RECT 17.505 -84.785 17.645 -84.615 ;
      RECT 17.555 -83.58 17.645 -82.572 ;
      RECT 17.505 -83.345 17.645 -83.175 ;
      RECT 17.555 -82.158 17.645 -81.15 ;
      RECT 17.505 -81.555 17.645 -81.385 ;
      RECT 17.555 -80.35 17.645 -79.342 ;
      RECT 17.505 -80.115 17.645 -79.945 ;
      RECT 17.555 -78.928 17.645 -77.92 ;
      RECT 17.505 -78.325 17.645 -78.155 ;
      RECT 17.555 -77.12 17.645 -76.112 ;
      RECT 17.505 -76.885 17.645 -76.715 ;
      RECT 17.555 -75.698 17.645 -74.69 ;
      RECT 17.505 -75.095 17.645 -74.925 ;
      RECT 17.555 -73.89 17.645 -72.882 ;
      RECT 17.505 -73.655 17.645 -73.485 ;
      RECT 17.555 -72.468 17.645 -71.46 ;
      RECT 17.505 -71.865 17.645 -71.695 ;
      RECT 17.555 -70.66 17.645 -69.652 ;
      RECT 17.505 -70.425 17.645 -70.255 ;
      RECT 17.555 -69.238 17.645 -68.23 ;
      RECT 17.505 -68.635 17.645 -68.465 ;
      RECT 17.555 -67.43 17.645 -66.422 ;
      RECT 17.505 -67.195 17.645 -67.025 ;
      RECT 17.555 -66.008 17.645 -65 ;
      RECT 17.505 -65.405 17.645 -65.235 ;
      RECT 17.555 -64.2 17.645 -63.192 ;
      RECT 17.505 -63.965 17.645 -63.795 ;
      RECT 17.555 -62.778 17.645 -61.77 ;
      RECT 17.505 -62.175 17.645 -62.005 ;
      RECT 17.555 -60.97 17.645 -59.962 ;
      RECT 17.505 -60.735 17.645 -60.565 ;
      RECT 17.555 -59.548 17.645 -58.54 ;
      RECT 17.505 -58.945 17.645 -58.775 ;
      RECT 17.555 -57.74 17.645 -56.732 ;
      RECT 17.505 -57.505 17.645 -57.335 ;
      RECT 17.555 -56.318 17.645 -55.31 ;
      RECT 17.505 -55.715 17.645 -55.545 ;
      RECT 17.555 -54.51 17.645 -53.502 ;
      RECT 17.505 -54.275 17.645 -54.105 ;
      RECT 17.555 -53.088 17.645 -52.08 ;
      RECT 17.505 -52.485 17.645 -52.315 ;
      RECT 17.555 -51.28 17.645 -50.272 ;
      RECT 17.505 -51.045 17.645 -50.875 ;
      RECT 17.555 -49.858 17.645 -48.85 ;
      RECT 17.505 -49.255 17.645 -49.085 ;
      RECT 17.555 -48.05 17.645 -47.042 ;
      RECT 17.505 -47.815 17.645 -47.645 ;
      RECT 17.555 -46.628 17.645 -45.62 ;
      RECT 17.505 -46.025 17.645 -45.855 ;
      RECT 17.555 -44.82 17.645 -43.812 ;
      RECT 17.505 -44.585 17.645 -44.415 ;
      RECT 17.555 -43.398 17.645 -42.39 ;
      RECT 17.505 -42.795 17.645 -42.625 ;
      RECT 17.555 -41.59 17.645 -40.582 ;
      RECT 17.505 -41.355 17.645 -41.185 ;
      RECT 17.555 -40.168 17.645 -39.16 ;
      RECT 17.505 -39.565 17.645 -39.395 ;
      RECT 17.555 -38.36 17.645 -37.352 ;
      RECT 17.505 -38.125 17.645 -37.955 ;
      RECT 17.555 -36.938 17.645 -35.93 ;
      RECT 17.505 -36.335 17.645 -36.165 ;
      RECT 17.555 -35.13 17.645 -34.122 ;
      RECT 17.505 -34.895 17.645 -34.725 ;
      RECT 17.555 -33.708 17.645 -32.7 ;
      RECT 17.505 -33.105 17.645 -32.935 ;
      RECT 17.555 -31.9 17.645 -30.892 ;
      RECT 17.505 -31.665 17.645 -31.495 ;
      RECT 17.555 -30.478 17.645 -29.47 ;
      RECT 17.505 -29.875 17.645 -29.705 ;
      RECT 17.555 -28.67 17.645 -27.662 ;
      RECT 17.505 -28.435 17.645 -28.265 ;
      RECT 17.555 -27.248 17.645 -26.24 ;
      RECT 17.505 -26.645 17.645 -26.475 ;
      RECT 17.555 -25.44 17.645 -24.432 ;
      RECT 17.505 -25.205 17.645 -25.035 ;
      RECT 17.555 -24.018 17.645 -23.01 ;
      RECT 17.505 -23.415 17.645 -23.245 ;
      RECT 17.555 -22.21 17.645 -21.202 ;
      RECT 17.505 -21.975 17.645 -21.805 ;
      RECT 17.555 -20.788 17.645 -19.78 ;
      RECT 17.505 -20.185 17.645 -20.015 ;
      RECT 17.555 -18.98 17.645 -17.972 ;
      RECT 17.505 -18.745 17.645 -18.575 ;
      RECT 17.555 -17.558 17.645 -16.55 ;
      RECT 17.505 -16.955 17.645 -16.785 ;
      RECT 17.555 -15.75 17.645 -14.742 ;
      RECT 17.505 -15.515 17.645 -15.345 ;
      RECT 17.555 -14.328 17.645 -13.32 ;
      RECT 17.505 -13.725 17.645 -13.555 ;
      RECT 17.555 -12.52 17.645 -11.512 ;
      RECT 17.505 -12.285 17.645 -12.115 ;
      RECT 17.555 -11.098 17.645 -10.09 ;
      RECT 17.505 -10.495 17.645 -10.325 ;
      RECT 17.555 -9.29 17.645 -8.282 ;
      RECT 17.505 -9.055 17.645 -8.885 ;
      RECT 17.555 -7.868 17.645 -6.86 ;
      RECT 17.505 -7.265 17.645 -7.095 ;
      RECT 17.555 -6.06 17.645 -5.052 ;
      RECT 17.505 -5.825 17.645 -5.655 ;
      RECT 17.555 -4.638 17.645 -3.63 ;
      RECT 17.505 -4.035 17.645 -3.865 ;
      RECT 17.555 -2.83 17.645 -1.822 ;
      RECT 17.505 -2.595 17.645 -2.425 ;
      RECT 17.555 -1.408 17.645 -0.4 ;
      RECT 17.505 -0.805 17.645 -0.635 ;
      RECT 17.555 0.4 17.645 1.408 ;
      RECT 17.505 0.635 17.645 0.805 ;
      RECT 17.155 -101.538 17.245 -100.531 ;
      RECT 17.155 -101.225 17.295 -101.055 ;
      RECT 17.155 -99.729 17.245 -98.722 ;
      RECT 17.155 -99.205 17.295 -99.035 ;
      RECT 17.155 -98.308 17.245 -97.301 ;
      RECT 17.155 -97.995 17.295 -97.825 ;
      RECT 17.155 -96.499 17.245 -95.492 ;
      RECT 17.155 -95.975 17.295 -95.805 ;
      RECT 17.155 -95.078 17.245 -94.071 ;
      RECT 17.155 -94.765 17.295 -94.595 ;
      RECT 17.155 -93.269 17.245 -92.262 ;
      RECT 17.155 -92.745 17.295 -92.575 ;
      RECT 17.155 -91.848 17.245 -90.841 ;
      RECT 17.155 -91.535 17.295 -91.365 ;
      RECT 17.155 -90.039 17.245 -89.032 ;
      RECT 17.155 -89.515 17.295 -89.345 ;
      RECT 17.155 -88.618 17.245 -87.611 ;
      RECT 17.155 -88.305 17.295 -88.135 ;
      RECT 17.155 -86.809 17.245 -85.802 ;
      RECT 17.155 -86.285 17.295 -86.115 ;
      RECT 17.155 -85.388 17.245 -84.381 ;
      RECT 17.155 -85.075 17.295 -84.905 ;
      RECT 17.155 -83.579 17.245 -82.572 ;
      RECT 17.155 -83.055 17.295 -82.885 ;
      RECT 17.155 -82.158 17.245 -81.151 ;
      RECT 17.155 -81.845 17.295 -81.675 ;
      RECT 17.155 -80.349 17.245 -79.342 ;
      RECT 17.155 -79.825 17.295 -79.655 ;
      RECT 17.155 -78.928 17.245 -77.921 ;
      RECT 17.155 -78.615 17.295 -78.445 ;
      RECT 17.155 -77.119 17.245 -76.112 ;
      RECT 17.155 -76.595 17.295 -76.425 ;
      RECT 17.155 -75.698 17.245 -74.691 ;
      RECT 17.155 -75.385 17.295 -75.215 ;
      RECT 17.155 -73.889 17.245 -72.882 ;
      RECT 17.155 -73.365 17.295 -73.195 ;
      RECT 17.155 -72.468 17.245 -71.461 ;
      RECT 17.155 -72.155 17.295 -71.985 ;
      RECT 17.155 -70.659 17.245 -69.652 ;
      RECT 17.155 -70.135 17.295 -69.965 ;
      RECT 17.155 -69.238 17.245 -68.231 ;
      RECT 17.155 -68.925 17.295 -68.755 ;
      RECT 17.155 -67.429 17.245 -66.422 ;
      RECT 17.155 -66.905 17.295 -66.735 ;
      RECT 17.155 -66.008 17.245 -65.001 ;
      RECT 17.155 -65.695 17.295 -65.525 ;
      RECT 17.155 -64.199 17.245 -63.192 ;
      RECT 17.155 -63.675 17.295 -63.505 ;
      RECT 17.155 -62.778 17.245 -61.771 ;
      RECT 17.155 -62.465 17.295 -62.295 ;
      RECT 17.155 -60.969 17.245 -59.962 ;
      RECT 17.155 -60.445 17.295 -60.275 ;
      RECT 17.155 -59.548 17.245 -58.541 ;
      RECT 17.155 -59.235 17.295 -59.065 ;
      RECT 17.155 -57.739 17.245 -56.732 ;
      RECT 17.155 -57.215 17.295 -57.045 ;
      RECT 17.155 -56.318 17.245 -55.311 ;
      RECT 17.155 -56.005 17.295 -55.835 ;
      RECT 17.155 -54.509 17.245 -53.502 ;
      RECT 17.155 -53.985 17.295 -53.815 ;
      RECT 17.155 -53.088 17.245 -52.081 ;
      RECT 17.155 -52.775 17.295 -52.605 ;
      RECT 17.155 -51.279 17.245 -50.272 ;
      RECT 17.155 -50.755 17.295 -50.585 ;
      RECT 17.155 -49.858 17.245 -48.851 ;
      RECT 17.155 -49.545 17.295 -49.375 ;
      RECT 17.155 -48.049 17.245 -47.042 ;
      RECT 17.155 -47.525 17.295 -47.355 ;
      RECT 17.155 -46.628 17.245 -45.621 ;
      RECT 17.155 -46.315 17.295 -46.145 ;
      RECT 17.155 -44.819 17.245 -43.812 ;
      RECT 17.155 -44.295 17.295 -44.125 ;
      RECT 17.155 -43.398 17.245 -42.391 ;
      RECT 17.155 -43.085 17.295 -42.915 ;
      RECT 17.155 -41.589 17.245 -40.582 ;
      RECT 17.155 -41.065 17.295 -40.895 ;
      RECT 17.155 -40.168 17.245 -39.161 ;
      RECT 17.155 -39.855 17.295 -39.685 ;
      RECT 17.155 -38.359 17.245 -37.352 ;
      RECT 17.155 -37.835 17.295 -37.665 ;
      RECT 17.155 -36.938 17.245 -35.931 ;
      RECT 17.155 -36.625 17.295 -36.455 ;
      RECT 17.155 -35.129 17.245 -34.122 ;
      RECT 17.155 -34.605 17.295 -34.435 ;
      RECT 17.155 -33.708 17.245 -32.701 ;
      RECT 17.155 -33.395 17.295 -33.225 ;
      RECT 17.155 -31.899 17.245 -30.892 ;
      RECT 17.155 -31.375 17.295 -31.205 ;
      RECT 17.155 -30.478 17.245 -29.471 ;
      RECT 17.155 -30.165 17.295 -29.995 ;
      RECT 17.155 -28.669 17.245 -27.662 ;
      RECT 17.155 -28.145 17.295 -27.975 ;
      RECT 17.155 -27.248 17.245 -26.241 ;
      RECT 17.155 -26.935 17.295 -26.765 ;
      RECT 17.155 -25.439 17.245 -24.432 ;
      RECT 17.155 -24.915 17.295 -24.745 ;
      RECT 17.155 -24.018 17.245 -23.011 ;
      RECT 17.155 -23.705 17.295 -23.535 ;
      RECT 17.155 -22.209 17.245 -21.202 ;
      RECT 17.155 -21.685 17.295 -21.515 ;
      RECT 17.155 -20.788 17.245 -19.781 ;
      RECT 17.155 -20.475 17.295 -20.305 ;
      RECT 17.155 -18.979 17.245 -17.972 ;
      RECT 17.155 -18.455 17.295 -18.285 ;
      RECT 17.155 -17.558 17.245 -16.551 ;
      RECT 17.155 -17.245 17.295 -17.075 ;
      RECT 17.155 -15.749 17.245 -14.742 ;
      RECT 17.155 -15.225 17.295 -15.055 ;
      RECT 17.155 -14.328 17.245 -13.321 ;
      RECT 17.155 -14.015 17.295 -13.845 ;
      RECT 17.155 -12.519 17.245 -11.512 ;
      RECT 17.155 -11.995 17.295 -11.825 ;
      RECT 17.155 -11.098 17.245 -10.091 ;
      RECT 17.155 -10.785 17.295 -10.615 ;
      RECT 17.155 -9.289 17.245 -8.282 ;
      RECT 17.155 -8.765 17.295 -8.595 ;
      RECT 17.155 -7.868 17.245 -6.861 ;
      RECT 17.155 -7.555 17.295 -7.385 ;
      RECT 17.155 -6.059 17.245 -5.052 ;
      RECT 17.155 -5.535 17.295 -5.365 ;
      RECT 17.155 -4.638 17.245 -3.631 ;
      RECT 17.155 -4.325 17.295 -4.155 ;
      RECT 17.155 -2.829 17.245 -1.822 ;
      RECT 17.155 -2.305 17.295 -2.135 ;
      RECT 17.155 -1.408 17.245 -0.401 ;
      RECT 17.155 -1.095 17.295 -0.925 ;
      RECT 17.155 0.401 17.245 1.408 ;
      RECT 17.155 0.925 17.295 1.095 ;
      RECT 15.305 -111.685 16.785 -111.585 ;
      RECT 15.305 -112.055 15.405 -111.585 ;
      RECT 15.11 -114.395 16.685 -114.275 ;
      RECT 16.585 -114.895 16.685 -114.275 ;
      RECT 15.99 -114.895 16.09 -114.275 ;
      RECT 15.11 -114.85 15.21 -114.275 ;
      RECT 16.355 -101.538 16.445 -100.53 ;
      RECT 16.305 -100.935 16.445 -100.765 ;
      RECT 16.355 -99.73 16.445 -98.722 ;
      RECT 16.305 -99.495 16.445 -99.325 ;
      RECT 16.355 -98.308 16.445 -97.3 ;
      RECT 16.305 -97.705 16.445 -97.535 ;
      RECT 16.355 -96.5 16.445 -95.492 ;
      RECT 16.305 -96.265 16.445 -96.095 ;
      RECT 16.355 -95.078 16.445 -94.07 ;
      RECT 16.305 -94.475 16.445 -94.305 ;
      RECT 16.355 -93.27 16.445 -92.262 ;
      RECT 16.305 -93.035 16.445 -92.865 ;
      RECT 16.355 -91.848 16.445 -90.84 ;
      RECT 16.305 -91.245 16.445 -91.075 ;
      RECT 16.355 -90.04 16.445 -89.032 ;
      RECT 16.305 -89.805 16.445 -89.635 ;
      RECT 16.355 -88.618 16.445 -87.61 ;
      RECT 16.305 -88.015 16.445 -87.845 ;
      RECT 16.355 -86.81 16.445 -85.802 ;
      RECT 16.305 -86.575 16.445 -86.405 ;
      RECT 16.355 -85.388 16.445 -84.38 ;
      RECT 16.305 -84.785 16.445 -84.615 ;
      RECT 16.355 -83.58 16.445 -82.572 ;
      RECT 16.305 -83.345 16.445 -83.175 ;
      RECT 16.355 -82.158 16.445 -81.15 ;
      RECT 16.305 -81.555 16.445 -81.385 ;
      RECT 16.355 -80.35 16.445 -79.342 ;
      RECT 16.305 -80.115 16.445 -79.945 ;
      RECT 16.355 -78.928 16.445 -77.92 ;
      RECT 16.305 -78.325 16.445 -78.155 ;
      RECT 16.355 -77.12 16.445 -76.112 ;
      RECT 16.305 -76.885 16.445 -76.715 ;
      RECT 16.355 -75.698 16.445 -74.69 ;
      RECT 16.305 -75.095 16.445 -74.925 ;
      RECT 16.355 -73.89 16.445 -72.882 ;
      RECT 16.305 -73.655 16.445 -73.485 ;
      RECT 16.355 -72.468 16.445 -71.46 ;
      RECT 16.305 -71.865 16.445 -71.695 ;
      RECT 16.355 -70.66 16.445 -69.652 ;
      RECT 16.305 -70.425 16.445 -70.255 ;
      RECT 16.355 -69.238 16.445 -68.23 ;
      RECT 16.305 -68.635 16.445 -68.465 ;
      RECT 16.355 -67.43 16.445 -66.422 ;
      RECT 16.305 -67.195 16.445 -67.025 ;
      RECT 16.355 -66.008 16.445 -65 ;
      RECT 16.305 -65.405 16.445 -65.235 ;
      RECT 16.355 -64.2 16.445 -63.192 ;
      RECT 16.305 -63.965 16.445 -63.795 ;
      RECT 16.355 -62.778 16.445 -61.77 ;
      RECT 16.305 -62.175 16.445 -62.005 ;
      RECT 16.355 -60.97 16.445 -59.962 ;
      RECT 16.305 -60.735 16.445 -60.565 ;
      RECT 16.355 -59.548 16.445 -58.54 ;
      RECT 16.305 -58.945 16.445 -58.775 ;
      RECT 16.355 -57.74 16.445 -56.732 ;
      RECT 16.305 -57.505 16.445 -57.335 ;
      RECT 16.355 -56.318 16.445 -55.31 ;
      RECT 16.305 -55.715 16.445 -55.545 ;
      RECT 16.355 -54.51 16.445 -53.502 ;
      RECT 16.305 -54.275 16.445 -54.105 ;
      RECT 16.355 -53.088 16.445 -52.08 ;
      RECT 16.305 -52.485 16.445 -52.315 ;
      RECT 16.355 -51.28 16.445 -50.272 ;
      RECT 16.305 -51.045 16.445 -50.875 ;
      RECT 16.355 -49.858 16.445 -48.85 ;
      RECT 16.305 -49.255 16.445 -49.085 ;
      RECT 16.355 -48.05 16.445 -47.042 ;
      RECT 16.305 -47.815 16.445 -47.645 ;
      RECT 16.355 -46.628 16.445 -45.62 ;
      RECT 16.305 -46.025 16.445 -45.855 ;
      RECT 16.355 -44.82 16.445 -43.812 ;
      RECT 16.305 -44.585 16.445 -44.415 ;
      RECT 16.355 -43.398 16.445 -42.39 ;
      RECT 16.305 -42.795 16.445 -42.625 ;
      RECT 16.355 -41.59 16.445 -40.582 ;
      RECT 16.305 -41.355 16.445 -41.185 ;
      RECT 16.355 -40.168 16.445 -39.16 ;
      RECT 16.305 -39.565 16.445 -39.395 ;
      RECT 16.355 -38.36 16.445 -37.352 ;
      RECT 16.305 -38.125 16.445 -37.955 ;
      RECT 16.355 -36.938 16.445 -35.93 ;
      RECT 16.305 -36.335 16.445 -36.165 ;
      RECT 16.355 -35.13 16.445 -34.122 ;
      RECT 16.305 -34.895 16.445 -34.725 ;
      RECT 16.355 -33.708 16.445 -32.7 ;
      RECT 16.305 -33.105 16.445 -32.935 ;
      RECT 16.355 -31.9 16.445 -30.892 ;
      RECT 16.305 -31.665 16.445 -31.495 ;
      RECT 16.355 -30.478 16.445 -29.47 ;
      RECT 16.305 -29.875 16.445 -29.705 ;
      RECT 16.355 -28.67 16.445 -27.662 ;
      RECT 16.305 -28.435 16.445 -28.265 ;
      RECT 16.355 -27.248 16.445 -26.24 ;
      RECT 16.305 -26.645 16.445 -26.475 ;
      RECT 16.355 -25.44 16.445 -24.432 ;
      RECT 16.305 -25.205 16.445 -25.035 ;
      RECT 16.355 -24.018 16.445 -23.01 ;
      RECT 16.305 -23.415 16.445 -23.245 ;
      RECT 16.355 -22.21 16.445 -21.202 ;
      RECT 16.305 -21.975 16.445 -21.805 ;
      RECT 16.355 -20.788 16.445 -19.78 ;
      RECT 16.305 -20.185 16.445 -20.015 ;
      RECT 16.355 -18.98 16.445 -17.972 ;
      RECT 16.305 -18.745 16.445 -18.575 ;
      RECT 16.355 -17.558 16.445 -16.55 ;
      RECT 16.305 -16.955 16.445 -16.785 ;
      RECT 16.355 -15.75 16.445 -14.742 ;
      RECT 16.305 -15.515 16.445 -15.345 ;
      RECT 16.355 -14.328 16.445 -13.32 ;
      RECT 16.305 -13.725 16.445 -13.555 ;
      RECT 16.355 -12.52 16.445 -11.512 ;
      RECT 16.305 -12.285 16.445 -12.115 ;
      RECT 16.355 -11.098 16.445 -10.09 ;
      RECT 16.305 -10.495 16.445 -10.325 ;
      RECT 16.355 -9.29 16.445 -8.282 ;
      RECT 16.305 -9.055 16.445 -8.885 ;
      RECT 16.355 -7.868 16.445 -6.86 ;
      RECT 16.305 -7.265 16.445 -7.095 ;
      RECT 16.355 -6.06 16.445 -5.052 ;
      RECT 16.305 -5.825 16.445 -5.655 ;
      RECT 16.355 -4.638 16.445 -3.63 ;
      RECT 16.305 -4.035 16.445 -3.865 ;
      RECT 16.355 -2.83 16.445 -1.822 ;
      RECT 16.305 -2.595 16.445 -2.425 ;
      RECT 16.355 -1.408 16.445 -0.4 ;
      RECT 16.305 -0.805 16.445 -0.635 ;
      RECT 16.355 0.4 16.445 1.408 ;
      RECT 16.305 0.635 16.445 0.805 ;
      RECT 16.23 -114.685 16.405 -114.515 ;
      RECT 16.305 -114.895 16.405 -114.515 ;
      RECT 15.345 -113.555 15.445 -113.09 ;
      RECT 15.71 -113.555 15.81 -113.1 ;
      RECT 15.345 -113.555 16.19 -113.385 ;
      RECT 15.955 -101.538 16.045 -100.531 ;
      RECT 15.955 -101.225 16.095 -101.055 ;
      RECT 15.955 -99.729 16.045 -98.722 ;
      RECT 15.955 -99.205 16.095 -99.035 ;
      RECT 15.955 -98.308 16.045 -97.301 ;
      RECT 15.955 -97.995 16.095 -97.825 ;
      RECT 15.955 -96.499 16.045 -95.492 ;
      RECT 15.955 -95.975 16.095 -95.805 ;
      RECT 15.955 -95.078 16.045 -94.071 ;
      RECT 15.955 -94.765 16.095 -94.595 ;
      RECT 15.955 -93.269 16.045 -92.262 ;
      RECT 15.955 -92.745 16.095 -92.575 ;
      RECT 15.955 -91.848 16.045 -90.841 ;
      RECT 15.955 -91.535 16.095 -91.365 ;
      RECT 15.955 -90.039 16.045 -89.032 ;
      RECT 15.955 -89.515 16.095 -89.345 ;
      RECT 15.955 -88.618 16.045 -87.611 ;
      RECT 15.955 -88.305 16.095 -88.135 ;
      RECT 15.955 -86.809 16.045 -85.802 ;
      RECT 15.955 -86.285 16.095 -86.115 ;
      RECT 15.955 -85.388 16.045 -84.381 ;
      RECT 15.955 -85.075 16.095 -84.905 ;
      RECT 15.955 -83.579 16.045 -82.572 ;
      RECT 15.955 -83.055 16.095 -82.885 ;
      RECT 15.955 -82.158 16.045 -81.151 ;
      RECT 15.955 -81.845 16.095 -81.675 ;
      RECT 15.955 -80.349 16.045 -79.342 ;
      RECT 15.955 -79.825 16.095 -79.655 ;
      RECT 15.955 -78.928 16.045 -77.921 ;
      RECT 15.955 -78.615 16.095 -78.445 ;
      RECT 15.955 -77.119 16.045 -76.112 ;
      RECT 15.955 -76.595 16.095 -76.425 ;
      RECT 15.955 -75.698 16.045 -74.691 ;
      RECT 15.955 -75.385 16.095 -75.215 ;
      RECT 15.955 -73.889 16.045 -72.882 ;
      RECT 15.955 -73.365 16.095 -73.195 ;
      RECT 15.955 -72.468 16.045 -71.461 ;
      RECT 15.955 -72.155 16.095 -71.985 ;
      RECT 15.955 -70.659 16.045 -69.652 ;
      RECT 15.955 -70.135 16.095 -69.965 ;
      RECT 15.955 -69.238 16.045 -68.231 ;
      RECT 15.955 -68.925 16.095 -68.755 ;
      RECT 15.955 -67.429 16.045 -66.422 ;
      RECT 15.955 -66.905 16.095 -66.735 ;
      RECT 15.955 -66.008 16.045 -65.001 ;
      RECT 15.955 -65.695 16.095 -65.525 ;
      RECT 15.955 -64.199 16.045 -63.192 ;
      RECT 15.955 -63.675 16.095 -63.505 ;
      RECT 15.955 -62.778 16.045 -61.771 ;
      RECT 15.955 -62.465 16.095 -62.295 ;
      RECT 15.955 -60.969 16.045 -59.962 ;
      RECT 15.955 -60.445 16.095 -60.275 ;
      RECT 15.955 -59.548 16.045 -58.541 ;
      RECT 15.955 -59.235 16.095 -59.065 ;
      RECT 15.955 -57.739 16.045 -56.732 ;
      RECT 15.955 -57.215 16.095 -57.045 ;
      RECT 15.955 -56.318 16.045 -55.311 ;
      RECT 15.955 -56.005 16.095 -55.835 ;
      RECT 15.955 -54.509 16.045 -53.502 ;
      RECT 15.955 -53.985 16.095 -53.815 ;
      RECT 15.955 -53.088 16.045 -52.081 ;
      RECT 15.955 -52.775 16.095 -52.605 ;
      RECT 15.955 -51.279 16.045 -50.272 ;
      RECT 15.955 -50.755 16.095 -50.585 ;
      RECT 15.955 -49.858 16.045 -48.851 ;
      RECT 15.955 -49.545 16.095 -49.375 ;
      RECT 15.955 -48.049 16.045 -47.042 ;
      RECT 15.955 -47.525 16.095 -47.355 ;
      RECT 15.955 -46.628 16.045 -45.621 ;
      RECT 15.955 -46.315 16.095 -46.145 ;
      RECT 15.955 -44.819 16.045 -43.812 ;
      RECT 15.955 -44.295 16.095 -44.125 ;
      RECT 15.955 -43.398 16.045 -42.391 ;
      RECT 15.955 -43.085 16.095 -42.915 ;
      RECT 15.955 -41.589 16.045 -40.582 ;
      RECT 15.955 -41.065 16.095 -40.895 ;
      RECT 15.955 -40.168 16.045 -39.161 ;
      RECT 15.955 -39.855 16.095 -39.685 ;
      RECT 15.955 -38.359 16.045 -37.352 ;
      RECT 15.955 -37.835 16.095 -37.665 ;
      RECT 15.955 -36.938 16.045 -35.931 ;
      RECT 15.955 -36.625 16.095 -36.455 ;
      RECT 15.955 -35.129 16.045 -34.122 ;
      RECT 15.955 -34.605 16.095 -34.435 ;
      RECT 15.955 -33.708 16.045 -32.701 ;
      RECT 15.955 -33.395 16.095 -33.225 ;
      RECT 15.955 -31.899 16.045 -30.892 ;
      RECT 15.955 -31.375 16.095 -31.205 ;
      RECT 15.955 -30.478 16.045 -29.471 ;
      RECT 15.955 -30.165 16.095 -29.995 ;
      RECT 15.955 -28.669 16.045 -27.662 ;
      RECT 15.955 -28.145 16.095 -27.975 ;
      RECT 15.955 -27.248 16.045 -26.241 ;
      RECT 15.955 -26.935 16.095 -26.765 ;
      RECT 15.955 -25.439 16.045 -24.432 ;
      RECT 15.955 -24.915 16.095 -24.745 ;
      RECT 15.955 -24.018 16.045 -23.011 ;
      RECT 15.955 -23.705 16.095 -23.535 ;
      RECT 15.955 -22.209 16.045 -21.202 ;
      RECT 15.955 -21.685 16.095 -21.515 ;
      RECT 15.955 -20.788 16.045 -19.781 ;
      RECT 15.955 -20.475 16.095 -20.305 ;
      RECT 15.955 -18.979 16.045 -17.972 ;
      RECT 15.955 -18.455 16.095 -18.285 ;
      RECT 15.955 -17.558 16.045 -16.551 ;
      RECT 15.955 -17.245 16.095 -17.075 ;
      RECT 15.955 -15.749 16.045 -14.742 ;
      RECT 15.955 -15.225 16.095 -15.055 ;
      RECT 15.955 -14.328 16.045 -13.321 ;
      RECT 15.955 -14.015 16.095 -13.845 ;
      RECT 15.955 -12.519 16.045 -11.512 ;
      RECT 15.955 -11.995 16.095 -11.825 ;
      RECT 15.955 -11.098 16.045 -10.091 ;
      RECT 15.955 -10.785 16.095 -10.615 ;
      RECT 15.955 -9.289 16.045 -8.282 ;
      RECT 15.955 -8.765 16.095 -8.595 ;
      RECT 15.955 -7.868 16.045 -6.861 ;
      RECT 15.955 -7.555 16.095 -7.385 ;
      RECT 15.955 -6.059 16.045 -5.052 ;
      RECT 15.955 -5.535 16.095 -5.365 ;
      RECT 15.955 -4.638 16.045 -3.631 ;
      RECT 15.955 -4.325 16.095 -4.155 ;
      RECT 15.955 -2.829 16.045 -1.822 ;
      RECT 15.955 -2.305 16.095 -2.135 ;
      RECT 15.955 -1.408 16.045 -0.401 ;
      RECT 15.955 -1.095 16.095 -0.925 ;
      RECT 15.955 0.401 16.045 1.408 ;
      RECT 15.955 0.925 16.095 1.095 ;
      RECT 15.64 -114.685 15.81 -114.515 ;
      RECT 15.71 -114.895 15.81 -114.515 ;
      RECT 15.155 -101.538 15.245 -100.53 ;
      RECT 15.105 -100.935 15.245 -100.765 ;
      RECT 15.155 -99.73 15.245 -98.722 ;
      RECT 15.105 -99.495 15.245 -99.325 ;
      RECT 15.155 -98.308 15.245 -97.3 ;
      RECT 15.105 -97.705 15.245 -97.535 ;
      RECT 15.155 -96.5 15.245 -95.492 ;
      RECT 15.105 -96.265 15.245 -96.095 ;
      RECT 15.155 -95.078 15.245 -94.07 ;
      RECT 15.105 -94.475 15.245 -94.305 ;
      RECT 15.155 -93.27 15.245 -92.262 ;
      RECT 15.105 -93.035 15.245 -92.865 ;
      RECT 15.155 -91.848 15.245 -90.84 ;
      RECT 15.105 -91.245 15.245 -91.075 ;
      RECT 15.155 -90.04 15.245 -89.032 ;
      RECT 15.105 -89.805 15.245 -89.635 ;
      RECT 15.155 -88.618 15.245 -87.61 ;
      RECT 15.105 -88.015 15.245 -87.845 ;
      RECT 15.155 -86.81 15.245 -85.802 ;
      RECT 15.105 -86.575 15.245 -86.405 ;
      RECT 15.155 -85.388 15.245 -84.38 ;
      RECT 15.105 -84.785 15.245 -84.615 ;
      RECT 15.155 -83.58 15.245 -82.572 ;
      RECT 15.105 -83.345 15.245 -83.175 ;
      RECT 15.155 -82.158 15.245 -81.15 ;
      RECT 15.105 -81.555 15.245 -81.385 ;
      RECT 15.155 -80.35 15.245 -79.342 ;
      RECT 15.105 -80.115 15.245 -79.945 ;
      RECT 15.155 -78.928 15.245 -77.92 ;
      RECT 15.105 -78.325 15.245 -78.155 ;
      RECT 15.155 -77.12 15.245 -76.112 ;
      RECT 15.105 -76.885 15.245 -76.715 ;
      RECT 15.155 -75.698 15.245 -74.69 ;
      RECT 15.105 -75.095 15.245 -74.925 ;
      RECT 15.155 -73.89 15.245 -72.882 ;
      RECT 15.105 -73.655 15.245 -73.485 ;
      RECT 15.155 -72.468 15.245 -71.46 ;
      RECT 15.105 -71.865 15.245 -71.695 ;
      RECT 15.155 -70.66 15.245 -69.652 ;
      RECT 15.105 -70.425 15.245 -70.255 ;
      RECT 15.155 -69.238 15.245 -68.23 ;
      RECT 15.105 -68.635 15.245 -68.465 ;
      RECT 15.155 -67.43 15.245 -66.422 ;
      RECT 15.105 -67.195 15.245 -67.025 ;
      RECT 15.155 -66.008 15.245 -65 ;
      RECT 15.105 -65.405 15.245 -65.235 ;
      RECT 15.155 -64.2 15.245 -63.192 ;
      RECT 15.105 -63.965 15.245 -63.795 ;
      RECT 15.155 -62.778 15.245 -61.77 ;
      RECT 15.105 -62.175 15.245 -62.005 ;
      RECT 15.155 -60.97 15.245 -59.962 ;
      RECT 15.105 -60.735 15.245 -60.565 ;
      RECT 15.155 -59.548 15.245 -58.54 ;
      RECT 15.105 -58.945 15.245 -58.775 ;
      RECT 15.155 -57.74 15.245 -56.732 ;
      RECT 15.105 -57.505 15.245 -57.335 ;
      RECT 15.155 -56.318 15.245 -55.31 ;
      RECT 15.105 -55.715 15.245 -55.545 ;
      RECT 15.155 -54.51 15.245 -53.502 ;
      RECT 15.105 -54.275 15.245 -54.105 ;
      RECT 15.155 -53.088 15.245 -52.08 ;
      RECT 15.105 -52.485 15.245 -52.315 ;
      RECT 15.155 -51.28 15.245 -50.272 ;
      RECT 15.105 -51.045 15.245 -50.875 ;
      RECT 15.155 -49.858 15.245 -48.85 ;
      RECT 15.105 -49.255 15.245 -49.085 ;
      RECT 15.155 -48.05 15.245 -47.042 ;
      RECT 15.105 -47.815 15.245 -47.645 ;
      RECT 15.155 -46.628 15.245 -45.62 ;
      RECT 15.105 -46.025 15.245 -45.855 ;
      RECT 15.155 -44.82 15.245 -43.812 ;
      RECT 15.105 -44.585 15.245 -44.415 ;
      RECT 15.155 -43.398 15.245 -42.39 ;
      RECT 15.105 -42.795 15.245 -42.625 ;
      RECT 15.155 -41.59 15.245 -40.582 ;
      RECT 15.105 -41.355 15.245 -41.185 ;
      RECT 15.155 -40.168 15.245 -39.16 ;
      RECT 15.105 -39.565 15.245 -39.395 ;
      RECT 15.155 -38.36 15.245 -37.352 ;
      RECT 15.105 -38.125 15.245 -37.955 ;
      RECT 15.155 -36.938 15.245 -35.93 ;
      RECT 15.105 -36.335 15.245 -36.165 ;
      RECT 15.155 -35.13 15.245 -34.122 ;
      RECT 15.105 -34.895 15.245 -34.725 ;
      RECT 15.155 -33.708 15.245 -32.7 ;
      RECT 15.105 -33.105 15.245 -32.935 ;
      RECT 15.155 -31.9 15.245 -30.892 ;
      RECT 15.105 -31.665 15.245 -31.495 ;
      RECT 15.155 -30.478 15.245 -29.47 ;
      RECT 15.105 -29.875 15.245 -29.705 ;
      RECT 15.155 -28.67 15.245 -27.662 ;
      RECT 15.105 -28.435 15.245 -28.265 ;
      RECT 15.155 -27.248 15.245 -26.24 ;
      RECT 15.105 -26.645 15.245 -26.475 ;
      RECT 15.155 -25.44 15.245 -24.432 ;
      RECT 15.105 -25.205 15.245 -25.035 ;
      RECT 15.155 -24.018 15.245 -23.01 ;
      RECT 15.105 -23.415 15.245 -23.245 ;
      RECT 15.155 -22.21 15.245 -21.202 ;
      RECT 15.105 -21.975 15.245 -21.805 ;
      RECT 15.155 -20.788 15.245 -19.78 ;
      RECT 15.105 -20.185 15.245 -20.015 ;
      RECT 15.155 -18.98 15.245 -17.972 ;
      RECT 15.105 -18.745 15.245 -18.575 ;
      RECT 15.155 -17.558 15.245 -16.55 ;
      RECT 15.105 -16.955 15.245 -16.785 ;
      RECT 15.155 -15.75 15.245 -14.742 ;
      RECT 15.105 -15.515 15.245 -15.345 ;
      RECT 15.155 -14.328 15.245 -13.32 ;
      RECT 15.105 -13.725 15.245 -13.555 ;
      RECT 15.155 -12.52 15.245 -11.512 ;
      RECT 15.105 -12.285 15.245 -12.115 ;
      RECT 15.155 -11.098 15.245 -10.09 ;
      RECT 15.105 -10.495 15.245 -10.325 ;
      RECT 15.155 -9.29 15.245 -8.282 ;
      RECT 15.105 -9.055 15.245 -8.885 ;
      RECT 15.155 -7.868 15.245 -6.86 ;
      RECT 15.105 -7.265 15.245 -7.095 ;
      RECT 15.155 -6.06 15.245 -5.052 ;
      RECT 15.105 -5.825 15.245 -5.655 ;
      RECT 15.155 -4.638 15.245 -3.63 ;
      RECT 15.105 -4.035 15.245 -3.865 ;
      RECT 15.155 -2.83 15.245 -1.822 ;
      RECT 15.105 -2.595 15.245 -2.425 ;
      RECT 15.155 -1.408 15.245 -0.4 ;
      RECT 15.105 -0.805 15.245 -0.635 ;
      RECT 15.155 0.4 15.245 1.408 ;
      RECT 15.105 0.635 15.245 0.805 ;
      RECT 14.755 -101.538 14.845 -100.531 ;
      RECT 14.755 -101.225 14.895 -101.055 ;
      RECT 14.755 -99.729 14.845 -98.722 ;
      RECT 14.755 -99.205 14.895 -99.035 ;
      RECT 14.755 -98.308 14.845 -97.301 ;
      RECT 14.755 -97.995 14.895 -97.825 ;
      RECT 14.755 -96.499 14.845 -95.492 ;
      RECT 14.755 -95.975 14.895 -95.805 ;
      RECT 14.755 -95.078 14.845 -94.071 ;
      RECT 14.755 -94.765 14.895 -94.595 ;
      RECT 14.755 -93.269 14.845 -92.262 ;
      RECT 14.755 -92.745 14.895 -92.575 ;
      RECT 14.755 -91.848 14.845 -90.841 ;
      RECT 14.755 -91.535 14.895 -91.365 ;
      RECT 14.755 -90.039 14.845 -89.032 ;
      RECT 14.755 -89.515 14.895 -89.345 ;
      RECT 14.755 -88.618 14.845 -87.611 ;
      RECT 14.755 -88.305 14.895 -88.135 ;
      RECT 14.755 -86.809 14.845 -85.802 ;
      RECT 14.755 -86.285 14.895 -86.115 ;
      RECT 14.755 -85.388 14.845 -84.381 ;
      RECT 14.755 -85.075 14.895 -84.905 ;
      RECT 14.755 -83.579 14.845 -82.572 ;
      RECT 14.755 -83.055 14.895 -82.885 ;
      RECT 14.755 -82.158 14.845 -81.151 ;
      RECT 14.755 -81.845 14.895 -81.675 ;
      RECT 14.755 -80.349 14.845 -79.342 ;
      RECT 14.755 -79.825 14.895 -79.655 ;
      RECT 14.755 -78.928 14.845 -77.921 ;
      RECT 14.755 -78.615 14.895 -78.445 ;
      RECT 14.755 -77.119 14.845 -76.112 ;
      RECT 14.755 -76.595 14.895 -76.425 ;
      RECT 14.755 -75.698 14.845 -74.691 ;
      RECT 14.755 -75.385 14.895 -75.215 ;
      RECT 14.755 -73.889 14.845 -72.882 ;
      RECT 14.755 -73.365 14.895 -73.195 ;
      RECT 14.755 -72.468 14.845 -71.461 ;
      RECT 14.755 -72.155 14.895 -71.985 ;
      RECT 14.755 -70.659 14.845 -69.652 ;
      RECT 14.755 -70.135 14.895 -69.965 ;
      RECT 14.755 -69.238 14.845 -68.231 ;
      RECT 14.755 -68.925 14.895 -68.755 ;
      RECT 14.755 -67.429 14.845 -66.422 ;
      RECT 14.755 -66.905 14.895 -66.735 ;
      RECT 14.755 -66.008 14.845 -65.001 ;
      RECT 14.755 -65.695 14.895 -65.525 ;
      RECT 14.755 -64.199 14.845 -63.192 ;
      RECT 14.755 -63.675 14.895 -63.505 ;
      RECT 14.755 -62.778 14.845 -61.771 ;
      RECT 14.755 -62.465 14.895 -62.295 ;
      RECT 14.755 -60.969 14.845 -59.962 ;
      RECT 14.755 -60.445 14.895 -60.275 ;
      RECT 14.755 -59.548 14.845 -58.541 ;
      RECT 14.755 -59.235 14.895 -59.065 ;
      RECT 14.755 -57.739 14.845 -56.732 ;
      RECT 14.755 -57.215 14.895 -57.045 ;
      RECT 14.755 -56.318 14.845 -55.311 ;
      RECT 14.755 -56.005 14.895 -55.835 ;
      RECT 14.755 -54.509 14.845 -53.502 ;
      RECT 14.755 -53.985 14.895 -53.815 ;
      RECT 14.755 -53.088 14.845 -52.081 ;
      RECT 14.755 -52.775 14.895 -52.605 ;
      RECT 14.755 -51.279 14.845 -50.272 ;
      RECT 14.755 -50.755 14.895 -50.585 ;
      RECT 14.755 -49.858 14.845 -48.851 ;
      RECT 14.755 -49.545 14.895 -49.375 ;
      RECT 14.755 -48.049 14.845 -47.042 ;
      RECT 14.755 -47.525 14.895 -47.355 ;
      RECT 14.755 -46.628 14.845 -45.621 ;
      RECT 14.755 -46.315 14.895 -46.145 ;
      RECT 14.755 -44.819 14.845 -43.812 ;
      RECT 14.755 -44.295 14.895 -44.125 ;
      RECT 14.755 -43.398 14.845 -42.391 ;
      RECT 14.755 -43.085 14.895 -42.915 ;
      RECT 14.755 -41.589 14.845 -40.582 ;
      RECT 14.755 -41.065 14.895 -40.895 ;
      RECT 14.755 -40.168 14.845 -39.161 ;
      RECT 14.755 -39.855 14.895 -39.685 ;
      RECT 14.755 -38.359 14.845 -37.352 ;
      RECT 14.755 -37.835 14.895 -37.665 ;
      RECT 14.755 -36.938 14.845 -35.931 ;
      RECT 14.755 -36.625 14.895 -36.455 ;
      RECT 14.755 -35.129 14.845 -34.122 ;
      RECT 14.755 -34.605 14.895 -34.435 ;
      RECT 14.755 -33.708 14.845 -32.701 ;
      RECT 14.755 -33.395 14.895 -33.225 ;
      RECT 14.755 -31.899 14.845 -30.892 ;
      RECT 14.755 -31.375 14.895 -31.205 ;
      RECT 14.755 -30.478 14.845 -29.471 ;
      RECT 14.755 -30.165 14.895 -29.995 ;
      RECT 14.755 -28.669 14.845 -27.662 ;
      RECT 14.755 -28.145 14.895 -27.975 ;
      RECT 14.755 -27.248 14.845 -26.241 ;
      RECT 14.755 -26.935 14.895 -26.765 ;
      RECT 14.755 -25.439 14.845 -24.432 ;
      RECT 14.755 -24.915 14.895 -24.745 ;
      RECT 14.755 -24.018 14.845 -23.011 ;
      RECT 14.755 -23.705 14.895 -23.535 ;
      RECT 14.755 -22.209 14.845 -21.202 ;
      RECT 14.755 -21.685 14.895 -21.515 ;
      RECT 14.755 -20.788 14.845 -19.781 ;
      RECT 14.755 -20.475 14.895 -20.305 ;
      RECT 14.755 -18.979 14.845 -17.972 ;
      RECT 14.755 -18.455 14.895 -18.285 ;
      RECT 14.755 -17.558 14.845 -16.551 ;
      RECT 14.755 -17.245 14.895 -17.075 ;
      RECT 14.755 -15.749 14.845 -14.742 ;
      RECT 14.755 -15.225 14.895 -15.055 ;
      RECT 14.755 -14.328 14.845 -13.321 ;
      RECT 14.755 -14.015 14.895 -13.845 ;
      RECT 14.755 -12.519 14.845 -11.512 ;
      RECT 14.755 -11.995 14.895 -11.825 ;
      RECT 14.755 -11.098 14.845 -10.091 ;
      RECT 14.755 -10.785 14.895 -10.615 ;
      RECT 14.755 -9.289 14.845 -8.282 ;
      RECT 14.755 -8.765 14.895 -8.595 ;
      RECT 14.755 -7.868 14.845 -6.861 ;
      RECT 14.755 -7.555 14.895 -7.385 ;
      RECT 14.755 -6.059 14.845 -5.052 ;
      RECT 14.755 -5.535 14.895 -5.365 ;
      RECT 14.755 -4.638 14.845 -3.631 ;
      RECT 14.755 -4.325 14.895 -4.155 ;
      RECT 14.755 -2.829 14.845 -1.822 ;
      RECT 14.755 -2.305 14.895 -2.135 ;
      RECT 14.755 -1.408 14.845 -0.401 ;
      RECT 14.755 -1.095 14.895 -0.925 ;
      RECT 14.755 0.401 14.845 1.408 ;
      RECT 14.755 0.925 14.895 1.095 ;
      RECT 10.585 -108.935 14.365 -108.815 ;
      RECT 11.905 -109.475 12.005 -108.815 ;
      RECT 11.345 -109.475 11.445 -108.815 ;
      RECT 10.785 -109.475 10.885 -108.815 ;
      RECT 13.955 -101.538 14.045 -100.53 ;
      RECT 13.905 -100.935 14.045 -100.765 ;
      RECT 13.955 -99.73 14.045 -98.722 ;
      RECT 13.905 -99.495 14.045 -99.325 ;
      RECT 13.955 -98.308 14.045 -97.3 ;
      RECT 13.905 -97.705 14.045 -97.535 ;
      RECT 13.955 -96.5 14.045 -95.492 ;
      RECT 13.905 -96.265 14.045 -96.095 ;
      RECT 13.955 -95.078 14.045 -94.07 ;
      RECT 13.905 -94.475 14.045 -94.305 ;
      RECT 13.955 -93.27 14.045 -92.262 ;
      RECT 13.905 -93.035 14.045 -92.865 ;
      RECT 13.955 -91.848 14.045 -90.84 ;
      RECT 13.905 -91.245 14.045 -91.075 ;
      RECT 13.955 -90.04 14.045 -89.032 ;
      RECT 13.905 -89.805 14.045 -89.635 ;
      RECT 13.955 -88.618 14.045 -87.61 ;
      RECT 13.905 -88.015 14.045 -87.845 ;
      RECT 13.955 -86.81 14.045 -85.802 ;
      RECT 13.905 -86.575 14.045 -86.405 ;
      RECT 13.955 -85.388 14.045 -84.38 ;
      RECT 13.905 -84.785 14.045 -84.615 ;
      RECT 13.955 -83.58 14.045 -82.572 ;
      RECT 13.905 -83.345 14.045 -83.175 ;
      RECT 13.955 -82.158 14.045 -81.15 ;
      RECT 13.905 -81.555 14.045 -81.385 ;
      RECT 13.955 -80.35 14.045 -79.342 ;
      RECT 13.905 -80.115 14.045 -79.945 ;
      RECT 13.955 -78.928 14.045 -77.92 ;
      RECT 13.905 -78.325 14.045 -78.155 ;
      RECT 13.955 -77.12 14.045 -76.112 ;
      RECT 13.905 -76.885 14.045 -76.715 ;
      RECT 13.955 -75.698 14.045 -74.69 ;
      RECT 13.905 -75.095 14.045 -74.925 ;
      RECT 13.955 -73.89 14.045 -72.882 ;
      RECT 13.905 -73.655 14.045 -73.485 ;
      RECT 13.955 -72.468 14.045 -71.46 ;
      RECT 13.905 -71.865 14.045 -71.695 ;
      RECT 13.955 -70.66 14.045 -69.652 ;
      RECT 13.905 -70.425 14.045 -70.255 ;
      RECT 13.955 -69.238 14.045 -68.23 ;
      RECT 13.905 -68.635 14.045 -68.465 ;
      RECT 13.955 -67.43 14.045 -66.422 ;
      RECT 13.905 -67.195 14.045 -67.025 ;
      RECT 13.955 -66.008 14.045 -65 ;
      RECT 13.905 -65.405 14.045 -65.235 ;
      RECT 13.955 -64.2 14.045 -63.192 ;
      RECT 13.905 -63.965 14.045 -63.795 ;
      RECT 13.955 -62.778 14.045 -61.77 ;
      RECT 13.905 -62.175 14.045 -62.005 ;
      RECT 13.955 -60.97 14.045 -59.962 ;
      RECT 13.905 -60.735 14.045 -60.565 ;
      RECT 13.955 -59.548 14.045 -58.54 ;
      RECT 13.905 -58.945 14.045 -58.775 ;
      RECT 13.955 -57.74 14.045 -56.732 ;
      RECT 13.905 -57.505 14.045 -57.335 ;
      RECT 13.955 -56.318 14.045 -55.31 ;
      RECT 13.905 -55.715 14.045 -55.545 ;
      RECT 13.955 -54.51 14.045 -53.502 ;
      RECT 13.905 -54.275 14.045 -54.105 ;
      RECT 13.955 -53.088 14.045 -52.08 ;
      RECT 13.905 -52.485 14.045 -52.315 ;
      RECT 13.955 -51.28 14.045 -50.272 ;
      RECT 13.905 -51.045 14.045 -50.875 ;
      RECT 13.955 -49.858 14.045 -48.85 ;
      RECT 13.905 -49.255 14.045 -49.085 ;
      RECT 13.955 -48.05 14.045 -47.042 ;
      RECT 13.905 -47.815 14.045 -47.645 ;
      RECT 13.955 -46.628 14.045 -45.62 ;
      RECT 13.905 -46.025 14.045 -45.855 ;
      RECT 13.955 -44.82 14.045 -43.812 ;
      RECT 13.905 -44.585 14.045 -44.415 ;
      RECT 13.955 -43.398 14.045 -42.39 ;
      RECT 13.905 -42.795 14.045 -42.625 ;
      RECT 13.955 -41.59 14.045 -40.582 ;
      RECT 13.905 -41.355 14.045 -41.185 ;
      RECT 13.955 -40.168 14.045 -39.16 ;
      RECT 13.905 -39.565 14.045 -39.395 ;
      RECT 13.955 -38.36 14.045 -37.352 ;
      RECT 13.905 -38.125 14.045 -37.955 ;
      RECT 13.955 -36.938 14.045 -35.93 ;
      RECT 13.905 -36.335 14.045 -36.165 ;
      RECT 13.955 -35.13 14.045 -34.122 ;
      RECT 13.905 -34.895 14.045 -34.725 ;
      RECT 13.955 -33.708 14.045 -32.7 ;
      RECT 13.905 -33.105 14.045 -32.935 ;
      RECT 13.955 -31.9 14.045 -30.892 ;
      RECT 13.905 -31.665 14.045 -31.495 ;
      RECT 13.955 -30.478 14.045 -29.47 ;
      RECT 13.905 -29.875 14.045 -29.705 ;
      RECT 13.955 -28.67 14.045 -27.662 ;
      RECT 13.905 -28.435 14.045 -28.265 ;
      RECT 13.955 -27.248 14.045 -26.24 ;
      RECT 13.905 -26.645 14.045 -26.475 ;
      RECT 13.955 -25.44 14.045 -24.432 ;
      RECT 13.905 -25.205 14.045 -25.035 ;
      RECT 13.955 -24.018 14.045 -23.01 ;
      RECT 13.905 -23.415 14.045 -23.245 ;
      RECT 13.955 -22.21 14.045 -21.202 ;
      RECT 13.905 -21.975 14.045 -21.805 ;
      RECT 13.955 -20.788 14.045 -19.78 ;
      RECT 13.905 -20.185 14.045 -20.015 ;
      RECT 13.955 -18.98 14.045 -17.972 ;
      RECT 13.905 -18.745 14.045 -18.575 ;
      RECT 13.955 -17.558 14.045 -16.55 ;
      RECT 13.905 -16.955 14.045 -16.785 ;
      RECT 13.955 -15.75 14.045 -14.742 ;
      RECT 13.905 -15.515 14.045 -15.345 ;
      RECT 13.955 -14.328 14.045 -13.32 ;
      RECT 13.905 -13.725 14.045 -13.555 ;
      RECT 13.955 -12.52 14.045 -11.512 ;
      RECT 13.905 -12.285 14.045 -12.115 ;
      RECT 13.955 -11.098 14.045 -10.09 ;
      RECT 13.905 -10.495 14.045 -10.325 ;
      RECT 13.955 -9.29 14.045 -8.282 ;
      RECT 13.905 -9.055 14.045 -8.885 ;
      RECT 13.955 -7.868 14.045 -6.86 ;
      RECT 13.905 -7.265 14.045 -7.095 ;
      RECT 13.955 -6.06 14.045 -5.052 ;
      RECT 13.905 -5.825 14.045 -5.655 ;
      RECT 13.955 -4.638 14.045 -3.63 ;
      RECT 13.905 -4.035 14.045 -3.865 ;
      RECT 13.955 -2.83 14.045 -1.822 ;
      RECT 13.905 -2.595 14.045 -2.425 ;
      RECT 13.955 -1.408 14.045 -0.4 ;
      RECT 13.905 -0.805 14.045 -0.635 ;
      RECT 13.955 0.4 14.045 1.408 ;
      RECT 13.905 0.635 14.045 0.805 ;
      RECT 12.525 -111.685 14.005 -111.585 ;
      RECT 12.525 -112.195 12.625 -111.585 ;
      RECT 12.745 -109.15 14.005 -109.05 ;
      RECT 13.905 -109.475 14.005 -109.05 ;
      RECT 13.345 -109.475 13.445 -109.05 ;
      RECT 12.785 -109.475 12.885 -109.05 ;
      RECT 13.555 -101.538 13.645 -100.531 ;
      RECT 13.555 -101.225 13.695 -101.055 ;
      RECT 13.555 -99.729 13.645 -98.722 ;
      RECT 13.555 -99.205 13.695 -99.035 ;
      RECT 13.555 -98.308 13.645 -97.301 ;
      RECT 13.555 -97.995 13.695 -97.825 ;
      RECT 13.555 -96.499 13.645 -95.492 ;
      RECT 13.555 -95.975 13.695 -95.805 ;
      RECT 13.555 -95.078 13.645 -94.071 ;
      RECT 13.555 -94.765 13.695 -94.595 ;
      RECT 13.555 -93.269 13.645 -92.262 ;
      RECT 13.555 -92.745 13.695 -92.575 ;
      RECT 13.555 -91.848 13.645 -90.841 ;
      RECT 13.555 -91.535 13.695 -91.365 ;
      RECT 13.555 -90.039 13.645 -89.032 ;
      RECT 13.555 -89.515 13.695 -89.345 ;
      RECT 13.555 -88.618 13.645 -87.611 ;
      RECT 13.555 -88.305 13.695 -88.135 ;
      RECT 13.555 -86.809 13.645 -85.802 ;
      RECT 13.555 -86.285 13.695 -86.115 ;
      RECT 13.555 -85.388 13.645 -84.381 ;
      RECT 13.555 -85.075 13.695 -84.905 ;
      RECT 13.555 -83.579 13.645 -82.572 ;
      RECT 13.555 -83.055 13.695 -82.885 ;
      RECT 13.555 -82.158 13.645 -81.151 ;
      RECT 13.555 -81.845 13.695 -81.675 ;
      RECT 13.555 -80.349 13.645 -79.342 ;
      RECT 13.555 -79.825 13.695 -79.655 ;
      RECT 13.555 -78.928 13.645 -77.921 ;
      RECT 13.555 -78.615 13.695 -78.445 ;
      RECT 13.555 -77.119 13.645 -76.112 ;
      RECT 13.555 -76.595 13.695 -76.425 ;
      RECT 13.555 -75.698 13.645 -74.691 ;
      RECT 13.555 -75.385 13.695 -75.215 ;
      RECT 13.555 -73.889 13.645 -72.882 ;
      RECT 13.555 -73.365 13.695 -73.195 ;
      RECT 13.555 -72.468 13.645 -71.461 ;
      RECT 13.555 -72.155 13.695 -71.985 ;
      RECT 13.555 -70.659 13.645 -69.652 ;
      RECT 13.555 -70.135 13.695 -69.965 ;
      RECT 13.555 -69.238 13.645 -68.231 ;
      RECT 13.555 -68.925 13.695 -68.755 ;
      RECT 13.555 -67.429 13.645 -66.422 ;
      RECT 13.555 -66.905 13.695 -66.735 ;
      RECT 13.555 -66.008 13.645 -65.001 ;
      RECT 13.555 -65.695 13.695 -65.525 ;
      RECT 13.555 -64.199 13.645 -63.192 ;
      RECT 13.555 -63.675 13.695 -63.505 ;
      RECT 13.555 -62.778 13.645 -61.771 ;
      RECT 13.555 -62.465 13.695 -62.295 ;
      RECT 13.555 -60.969 13.645 -59.962 ;
      RECT 13.555 -60.445 13.695 -60.275 ;
      RECT 13.555 -59.548 13.645 -58.541 ;
      RECT 13.555 -59.235 13.695 -59.065 ;
      RECT 13.555 -57.739 13.645 -56.732 ;
      RECT 13.555 -57.215 13.695 -57.045 ;
      RECT 13.555 -56.318 13.645 -55.311 ;
      RECT 13.555 -56.005 13.695 -55.835 ;
      RECT 13.555 -54.509 13.645 -53.502 ;
      RECT 13.555 -53.985 13.695 -53.815 ;
      RECT 13.555 -53.088 13.645 -52.081 ;
      RECT 13.555 -52.775 13.695 -52.605 ;
      RECT 13.555 -51.279 13.645 -50.272 ;
      RECT 13.555 -50.755 13.695 -50.585 ;
      RECT 13.555 -49.858 13.645 -48.851 ;
      RECT 13.555 -49.545 13.695 -49.375 ;
      RECT 13.555 -48.049 13.645 -47.042 ;
      RECT 13.555 -47.525 13.695 -47.355 ;
      RECT 13.555 -46.628 13.645 -45.621 ;
      RECT 13.555 -46.315 13.695 -46.145 ;
      RECT 13.555 -44.819 13.645 -43.812 ;
      RECT 13.555 -44.295 13.695 -44.125 ;
      RECT 13.555 -43.398 13.645 -42.391 ;
      RECT 13.555 -43.085 13.695 -42.915 ;
      RECT 13.555 -41.589 13.645 -40.582 ;
      RECT 13.555 -41.065 13.695 -40.895 ;
      RECT 13.555 -40.168 13.645 -39.161 ;
      RECT 13.555 -39.855 13.695 -39.685 ;
      RECT 13.555 -38.359 13.645 -37.352 ;
      RECT 13.555 -37.835 13.695 -37.665 ;
      RECT 13.555 -36.938 13.645 -35.931 ;
      RECT 13.555 -36.625 13.695 -36.455 ;
      RECT 13.555 -35.129 13.645 -34.122 ;
      RECT 13.555 -34.605 13.695 -34.435 ;
      RECT 13.555 -33.708 13.645 -32.701 ;
      RECT 13.555 -33.395 13.695 -33.225 ;
      RECT 13.555 -31.899 13.645 -30.892 ;
      RECT 13.555 -31.375 13.695 -31.205 ;
      RECT 13.555 -30.478 13.645 -29.471 ;
      RECT 13.555 -30.165 13.695 -29.995 ;
      RECT 13.555 -28.669 13.645 -27.662 ;
      RECT 13.555 -28.145 13.695 -27.975 ;
      RECT 13.555 -27.248 13.645 -26.241 ;
      RECT 13.555 -26.935 13.695 -26.765 ;
      RECT 13.555 -25.439 13.645 -24.432 ;
      RECT 13.555 -24.915 13.695 -24.745 ;
      RECT 13.555 -24.018 13.645 -23.011 ;
      RECT 13.555 -23.705 13.695 -23.535 ;
      RECT 13.555 -22.209 13.645 -21.202 ;
      RECT 13.555 -21.685 13.695 -21.515 ;
      RECT 13.555 -20.788 13.645 -19.781 ;
      RECT 13.555 -20.475 13.695 -20.305 ;
      RECT 13.555 -18.979 13.645 -17.972 ;
      RECT 13.555 -18.455 13.695 -18.285 ;
      RECT 13.555 -17.558 13.645 -16.551 ;
      RECT 13.555 -17.245 13.695 -17.075 ;
      RECT 13.555 -15.749 13.645 -14.742 ;
      RECT 13.555 -15.225 13.695 -15.055 ;
      RECT 13.555 -14.328 13.645 -13.321 ;
      RECT 13.555 -14.015 13.695 -13.845 ;
      RECT 13.555 -12.519 13.645 -11.512 ;
      RECT 13.555 -11.995 13.695 -11.825 ;
      RECT 13.555 -11.098 13.645 -10.091 ;
      RECT 13.555 -10.785 13.695 -10.615 ;
      RECT 13.555 -9.289 13.645 -8.282 ;
      RECT 13.555 -8.765 13.695 -8.595 ;
      RECT 13.555 -7.868 13.645 -6.861 ;
      RECT 13.555 -7.555 13.695 -7.385 ;
      RECT 13.555 -6.059 13.645 -5.052 ;
      RECT 13.555 -5.535 13.695 -5.365 ;
      RECT 13.555 -4.638 13.645 -3.631 ;
      RECT 13.555 -4.325 13.695 -4.155 ;
      RECT 13.555 -2.829 13.645 -1.822 ;
      RECT 13.555 -2.305 13.695 -2.135 ;
      RECT 13.555 -1.408 13.645 -0.401 ;
      RECT 13.555 -1.095 13.695 -0.925 ;
      RECT 13.555 0.401 13.645 1.408 ;
      RECT 13.555 0.925 13.695 1.095 ;
      RECT 12.885 -111.495 13.055 -111.385 ;
      RECT 9.735 -111.495 13.055 -111.395 ;
      RECT 12.755 -101.538 12.845 -100.53 ;
      RECT 12.705 -100.935 12.845 -100.765 ;
      RECT 12.755 -99.73 12.845 -98.722 ;
      RECT 12.705 -99.495 12.845 -99.325 ;
      RECT 12.755 -98.308 12.845 -97.3 ;
      RECT 12.705 -97.705 12.845 -97.535 ;
      RECT 12.755 -96.5 12.845 -95.492 ;
      RECT 12.705 -96.265 12.845 -96.095 ;
      RECT 12.755 -95.078 12.845 -94.07 ;
      RECT 12.705 -94.475 12.845 -94.305 ;
      RECT 12.755 -93.27 12.845 -92.262 ;
      RECT 12.705 -93.035 12.845 -92.865 ;
      RECT 12.755 -91.848 12.845 -90.84 ;
      RECT 12.705 -91.245 12.845 -91.075 ;
      RECT 12.755 -90.04 12.845 -89.032 ;
      RECT 12.705 -89.805 12.845 -89.635 ;
      RECT 12.755 -88.618 12.845 -87.61 ;
      RECT 12.705 -88.015 12.845 -87.845 ;
      RECT 12.755 -86.81 12.845 -85.802 ;
      RECT 12.705 -86.575 12.845 -86.405 ;
      RECT 12.755 -85.388 12.845 -84.38 ;
      RECT 12.705 -84.785 12.845 -84.615 ;
      RECT 12.755 -83.58 12.845 -82.572 ;
      RECT 12.705 -83.345 12.845 -83.175 ;
      RECT 12.755 -82.158 12.845 -81.15 ;
      RECT 12.705 -81.555 12.845 -81.385 ;
      RECT 12.755 -80.35 12.845 -79.342 ;
      RECT 12.705 -80.115 12.845 -79.945 ;
      RECT 12.755 -78.928 12.845 -77.92 ;
      RECT 12.705 -78.325 12.845 -78.155 ;
      RECT 12.755 -77.12 12.845 -76.112 ;
      RECT 12.705 -76.885 12.845 -76.715 ;
      RECT 12.755 -75.698 12.845 -74.69 ;
      RECT 12.705 -75.095 12.845 -74.925 ;
      RECT 12.755 -73.89 12.845 -72.882 ;
      RECT 12.705 -73.655 12.845 -73.485 ;
      RECT 12.755 -72.468 12.845 -71.46 ;
      RECT 12.705 -71.865 12.845 -71.695 ;
      RECT 12.755 -70.66 12.845 -69.652 ;
      RECT 12.705 -70.425 12.845 -70.255 ;
      RECT 12.755 -69.238 12.845 -68.23 ;
      RECT 12.705 -68.635 12.845 -68.465 ;
      RECT 12.755 -67.43 12.845 -66.422 ;
      RECT 12.705 -67.195 12.845 -67.025 ;
      RECT 12.755 -66.008 12.845 -65 ;
      RECT 12.705 -65.405 12.845 -65.235 ;
      RECT 12.755 -64.2 12.845 -63.192 ;
      RECT 12.705 -63.965 12.845 -63.795 ;
      RECT 12.755 -62.778 12.845 -61.77 ;
      RECT 12.705 -62.175 12.845 -62.005 ;
      RECT 12.755 -60.97 12.845 -59.962 ;
      RECT 12.705 -60.735 12.845 -60.565 ;
      RECT 12.755 -59.548 12.845 -58.54 ;
      RECT 12.705 -58.945 12.845 -58.775 ;
      RECT 12.755 -57.74 12.845 -56.732 ;
      RECT 12.705 -57.505 12.845 -57.335 ;
      RECT 12.755 -56.318 12.845 -55.31 ;
      RECT 12.705 -55.715 12.845 -55.545 ;
      RECT 12.755 -54.51 12.845 -53.502 ;
      RECT 12.705 -54.275 12.845 -54.105 ;
      RECT 12.755 -53.088 12.845 -52.08 ;
      RECT 12.705 -52.485 12.845 -52.315 ;
      RECT 12.755 -51.28 12.845 -50.272 ;
      RECT 12.705 -51.045 12.845 -50.875 ;
      RECT 12.755 -49.858 12.845 -48.85 ;
      RECT 12.705 -49.255 12.845 -49.085 ;
      RECT 12.755 -48.05 12.845 -47.042 ;
      RECT 12.705 -47.815 12.845 -47.645 ;
      RECT 12.755 -46.628 12.845 -45.62 ;
      RECT 12.705 -46.025 12.845 -45.855 ;
      RECT 12.755 -44.82 12.845 -43.812 ;
      RECT 12.705 -44.585 12.845 -44.415 ;
      RECT 12.755 -43.398 12.845 -42.39 ;
      RECT 12.705 -42.795 12.845 -42.625 ;
      RECT 12.755 -41.59 12.845 -40.582 ;
      RECT 12.705 -41.355 12.845 -41.185 ;
      RECT 12.755 -40.168 12.845 -39.16 ;
      RECT 12.705 -39.565 12.845 -39.395 ;
      RECT 12.755 -38.36 12.845 -37.352 ;
      RECT 12.705 -38.125 12.845 -37.955 ;
      RECT 12.755 -36.938 12.845 -35.93 ;
      RECT 12.705 -36.335 12.845 -36.165 ;
      RECT 12.755 -35.13 12.845 -34.122 ;
      RECT 12.705 -34.895 12.845 -34.725 ;
      RECT 12.755 -33.708 12.845 -32.7 ;
      RECT 12.705 -33.105 12.845 -32.935 ;
      RECT 12.755 -31.9 12.845 -30.892 ;
      RECT 12.705 -31.665 12.845 -31.495 ;
      RECT 12.755 -30.478 12.845 -29.47 ;
      RECT 12.705 -29.875 12.845 -29.705 ;
      RECT 12.755 -28.67 12.845 -27.662 ;
      RECT 12.705 -28.435 12.845 -28.265 ;
      RECT 12.755 -27.248 12.845 -26.24 ;
      RECT 12.705 -26.645 12.845 -26.475 ;
      RECT 12.755 -25.44 12.845 -24.432 ;
      RECT 12.705 -25.205 12.845 -25.035 ;
      RECT 12.755 -24.018 12.845 -23.01 ;
      RECT 12.705 -23.415 12.845 -23.245 ;
      RECT 12.755 -22.21 12.845 -21.202 ;
      RECT 12.705 -21.975 12.845 -21.805 ;
      RECT 12.755 -20.788 12.845 -19.78 ;
      RECT 12.705 -20.185 12.845 -20.015 ;
      RECT 12.755 -18.98 12.845 -17.972 ;
      RECT 12.705 -18.745 12.845 -18.575 ;
      RECT 12.755 -17.558 12.845 -16.55 ;
      RECT 12.705 -16.955 12.845 -16.785 ;
      RECT 12.755 -15.75 12.845 -14.742 ;
      RECT 12.705 -15.515 12.845 -15.345 ;
      RECT 12.755 -14.328 12.845 -13.32 ;
      RECT 12.705 -13.725 12.845 -13.555 ;
      RECT 12.755 -12.52 12.845 -11.512 ;
      RECT 12.705 -12.285 12.845 -12.115 ;
      RECT 12.755 -11.098 12.845 -10.09 ;
      RECT 12.705 -10.495 12.845 -10.325 ;
      RECT 12.755 -9.29 12.845 -8.282 ;
      RECT 12.705 -9.055 12.845 -8.885 ;
      RECT 12.755 -7.868 12.845 -6.86 ;
      RECT 12.705 -7.265 12.845 -7.095 ;
      RECT 12.755 -6.06 12.845 -5.052 ;
      RECT 12.705 -5.825 12.845 -5.655 ;
      RECT 12.755 -4.638 12.845 -3.63 ;
      RECT 12.705 -4.035 12.845 -3.865 ;
      RECT 12.755 -2.83 12.845 -1.822 ;
      RECT 12.705 -2.595 12.845 -2.425 ;
      RECT 12.755 -1.408 12.845 -0.4 ;
      RECT 12.705 -0.805 12.845 -0.635 ;
      RECT 12.755 0.4 12.845 1.408 ;
      RECT 12.705 0.635 12.845 0.805 ;
      RECT 12.355 -101.538 12.445 -100.531 ;
      RECT 12.355 -101.225 12.495 -101.055 ;
      RECT 12.355 -99.729 12.445 -98.722 ;
      RECT 12.355 -99.205 12.495 -99.035 ;
      RECT 12.355 -98.308 12.445 -97.301 ;
      RECT 12.355 -97.995 12.495 -97.825 ;
      RECT 12.355 -96.499 12.445 -95.492 ;
      RECT 12.355 -95.975 12.495 -95.805 ;
      RECT 12.355 -95.078 12.445 -94.071 ;
      RECT 12.355 -94.765 12.495 -94.595 ;
      RECT 12.355 -93.269 12.445 -92.262 ;
      RECT 12.355 -92.745 12.495 -92.575 ;
      RECT 12.355 -91.848 12.445 -90.841 ;
      RECT 12.355 -91.535 12.495 -91.365 ;
      RECT 12.355 -90.039 12.445 -89.032 ;
      RECT 12.355 -89.515 12.495 -89.345 ;
      RECT 12.355 -88.618 12.445 -87.611 ;
      RECT 12.355 -88.305 12.495 -88.135 ;
      RECT 12.355 -86.809 12.445 -85.802 ;
      RECT 12.355 -86.285 12.495 -86.115 ;
      RECT 12.355 -85.388 12.445 -84.381 ;
      RECT 12.355 -85.075 12.495 -84.905 ;
      RECT 12.355 -83.579 12.445 -82.572 ;
      RECT 12.355 -83.055 12.495 -82.885 ;
      RECT 12.355 -82.158 12.445 -81.151 ;
      RECT 12.355 -81.845 12.495 -81.675 ;
      RECT 12.355 -80.349 12.445 -79.342 ;
      RECT 12.355 -79.825 12.495 -79.655 ;
      RECT 12.355 -78.928 12.445 -77.921 ;
      RECT 12.355 -78.615 12.495 -78.445 ;
      RECT 12.355 -77.119 12.445 -76.112 ;
      RECT 12.355 -76.595 12.495 -76.425 ;
      RECT 12.355 -75.698 12.445 -74.691 ;
      RECT 12.355 -75.385 12.495 -75.215 ;
      RECT 12.355 -73.889 12.445 -72.882 ;
      RECT 12.355 -73.365 12.495 -73.195 ;
      RECT 12.355 -72.468 12.445 -71.461 ;
      RECT 12.355 -72.155 12.495 -71.985 ;
      RECT 12.355 -70.659 12.445 -69.652 ;
      RECT 12.355 -70.135 12.495 -69.965 ;
      RECT 12.355 -69.238 12.445 -68.231 ;
      RECT 12.355 -68.925 12.495 -68.755 ;
      RECT 12.355 -67.429 12.445 -66.422 ;
      RECT 12.355 -66.905 12.495 -66.735 ;
      RECT 12.355 -66.008 12.445 -65.001 ;
      RECT 12.355 -65.695 12.495 -65.525 ;
      RECT 12.355 -64.199 12.445 -63.192 ;
      RECT 12.355 -63.675 12.495 -63.505 ;
      RECT 12.355 -62.778 12.445 -61.771 ;
      RECT 12.355 -62.465 12.495 -62.295 ;
      RECT 12.355 -60.969 12.445 -59.962 ;
      RECT 12.355 -60.445 12.495 -60.275 ;
      RECT 12.355 -59.548 12.445 -58.541 ;
      RECT 12.355 -59.235 12.495 -59.065 ;
      RECT 12.355 -57.739 12.445 -56.732 ;
      RECT 12.355 -57.215 12.495 -57.045 ;
      RECT 12.355 -56.318 12.445 -55.311 ;
      RECT 12.355 -56.005 12.495 -55.835 ;
      RECT 12.355 -54.509 12.445 -53.502 ;
      RECT 12.355 -53.985 12.495 -53.815 ;
      RECT 12.355 -53.088 12.445 -52.081 ;
      RECT 12.355 -52.775 12.495 -52.605 ;
      RECT 12.355 -51.279 12.445 -50.272 ;
      RECT 12.355 -50.755 12.495 -50.585 ;
      RECT 12.355 -49.858 12.445 -48.851 ;
      RECT 12.355 -49.545 12.495 -49.375 ;
      RECT 12.355 -48.049 12.445 -47.042 ;
      RECT 12.355 -47.525 12.495 -47.355 ;
      RECT 12.355 -46.628 12.445 -45.621 ;
      RECT 12.355 -46.315 12.495 -46.145 ;
      RECT 12.355 -44.819 12.445 -43.812 ;
      RECT 12.355 -44.295 12.495 -44.125 ;
      RECT 12.355 -43.398 12.445 -42.391 ;
      RECT 12.355 -43.085 12.495 -42.915 ;
      RECT 12.355 -41.589 12.445 -40.582 ;
      RECT 12.355 -41.065 12.495 -40.895 ;
      RECT 12.355 -40.168 12.445 -39.161 ;
      RECT 12.355 -39.855 12.495 -39.685 ;
      RECT 12.355 -38.359 12.445 -37.352 ;
      RECT 12.355 -37.835 12.495 -37.665 ;
      RECT 12.355 -36.938 12.445 -35.931 ;
      RECT 12.355 -36.625 12.495 -36.455 ;
      RECT 12.355 -35.129 12.445 -34.122 ;
      RECT 12.355 -34.605 12.495 -34.435 ;
      RECT 12.355 -33.708 12.445 -32.701 ;
      RECT 12.355 -33.395 12.495 -33.225 ;
      RECT 12.355 -31.899 12.445 -30.892 ;
      RECT 12.355 -31.375 12.495 -31.205 ;
      RECT 12.355 -30.478 12.445 -29.471 ;
      RECT 12.355 -30.165 12.495 -29.995 ;
      RECT 12.355 -28.669 12.445 -27.662 ;
      RECT 12.355 -28.145 12.495 -27.975 ;
      RECT 12.355 -27.248 12.445 -26.241 ;
      RECT 12.355 -26.935 12.495 -26.765 ;
      RECT 12.355 -25.439 12.445 -24.432 ;
      RECT 12.355 -24.915 12.495 -24.745 ;
      RECT 12.355 -24.018 12.445 -23.011 ;
      RECT 12.355 -23.705 12.495 -23.535 ;
      RECT 12.355 -22.209 12.445 -21.202 ;
      RECT 12.355 -21.685 12.495 -21.515 ;
      RECT 12.355 -20.788 12.445 -19.781 ;
      RECT 12.355 -20.475 12.495 -20.305 ;
      RECT 12.355 -18.979 12.445 -17.972 ;
      RECT 12.355 -18.455 12.495 -18.285 ;
      RECT 12.355 -17.558 12.445 -16.551 ;
      RECT 12.355 -17.245 12.495 -17.075 ;
      RECT 12.355 -15.749 12.445 -14.742 ;
      RECT 12.355 -15.225 12.495 -15.055 ;
      RECT 12.355 -14.328 12.445 -13.321 ;
      RECT 12.355 -14.015 12.495 -13.845 ;
      RECT 12.355 -12.519 12.445 -11.512 ;
      RECT 12.355 -11.995 12.495 -11.825 ;
      RECT 12.355 -11.098 12.445 -10.091 ;
      RECT 12.355 -10.785 12.495 -10.615 ;
      RECT 12.355 -9.289 12.445 -8.282 ;
      RECT 12.355 -8.765 12.495 -8.595 ;
      RECT 12.355 -7.868 12.445 -6.861 ;
      RECT 12.355 -7.555 12.495 -7.385 ;
      RECT 12.355 -6.059 12.445 -5.052 ;
      RECT 12.355 -5.535 12.495 -5.365 ;
      RECT 12.355 -4.638 12.445 -3.631 ;
      RECT 12.355 -4.325 12.495 -4.155 ;
      RECT 12.355 -2.829 12.445 -1.822 ;
      RECT 12.355 -2.305 12.495 -2.135 ;
      RECT 12.355 -1.408 12.445 -0.401 ;
      RECT 12.355 -1.095 12.495 -0.925 ;
      RECT 12.355 0.401 12.445 1.408 ;
      RECT 12.355 0.925 12.495 1.095 ;
      RECT 10.505 -111.685 11.985 -111.585 ;
      RECT 10.505 -112.055 10.605 -111.585 ;
      RECT 10.31 -114.395 11.885 -114.275 ;
      RECT 11.785 -114.895 11.885 -114.275 ;
      RECT 11.19 -114.895 11.29 -114.275 ;
      RECT 10.31 -114.85 10.41 -114.275 ;
      RECT 11.555 -101.538 11.645 -100.53 ;
      RECT 11.505 -100.935 11.645 -100.765 ;
      RECT 11.555 -99.73 11.645 -98.722 ;
      RECT 11.505 -99.495 11.645 -99.325 ;
      RECT 11.555 -98.308 11.645 -97.3 ;
      RECT 11.505 -97.705 11.645 -97.535 ;
      RECT 11.555 -96.5 11.645 -95.492 ;
      RECT 11.505 -96.265 11.645 -96.095 ;
      RECT 11.555 -95.078 11.645 -94.07 ;
      RECT 11.505 -94.475 11.645 -94.305 ;
      RECT 11.555 -93.27 11.645 -92.262 ;
      RECT 11.505 -93.035 11.645 -92.865 ;
      RECT 11.555 -91.848 11.645 -90.84 ;
      RECT 11.505 -91.245 11.645 -91.075 ;
      RECT 11.555 -90.04 11.645 -89.032 ;
      RECT 11.505 -89.805 11.645 -89.635 ;
      RECT 11.555 -88.618 11.645 -87.61 ;
      RECT 11.505 -88.015 11.645 -87.845 ;
      RECT 11.555 -86.81 11.645 -85.802 ;
      RECT 11.505 -86.575 11.645 -86.405 ;
      RECT 11.555 -85.388 11.645 -84.38 ;
      RECT 11.505 -84.785 11.645 -84.615 ;
      RECT 11.555 -83.58 11.645 -82.572 ;
      RECT 11.505 -83.345 11.645 -83.175 ;
      RECT 11.555 -82.158 11.645 -81.15 ;
      RECT 11.505 -81.555 11.645 -81.385 ;
      RECT 11.555 -80.35 11.645 -79.342 ;
      RECT 11.505 -80.115 11.645 -79.945 ;
      RECT 11.555 -78.928 11.645 -77.92 ;
      RECT 11.505 -78.325 11.645 -78.155 ;
      RECT 11.555 -77.12 11.645 -76.112 ;
      RECT 11.505 -76.885 11.645 -76.715 ;
      RECT 11.555 -75.698 11.645 -74.69 ;
      RECT 11.505 -75.095 11.645 -74.925 ;
      RECT 11.555 -73.89 11.645 -72.882 ;
      RECT 11.505 -73.655 11.645 -73.485 ;
      RECT 11.555 -72.468 11.645 -71.46 ;
      RECT 11.505 -71.865 11.645 -71.695 ;
      RECT 11.555 -70.66 11.645 -69.652 ;
      RECT 11.505 -70.425 11.645 -70.255 ;
      RECT 11.555 -69.238 11.645 -68.23 ;
      RECT 11.505 -68.635 11.645 -68.465 ;
      RECT 11.555 -67.43 11.645 -66.422 ;
      RECT 11.505 -67.195 11.645 -67.025 ;
      RECT 11.555 -66.008 11.645 -65 ;
      RECT 11.505 -65.405 11.645 -65.235 ;
      RECT 11.555 -64.2 11.645 -63.192 ;
      RECT 11.505 -63.965 11.645 -63.795 ;
      RECT 11.555 -62.778 11.645 -61.77 ;
      RECT 11.505 -62.175 11.645 -62.005 ;
      RECT 11.555 -60.97 11.645 -59.962 ;
      RECT 11.505 -60.735 11.645 -60.565 ;
      RECT 11.555 -59.548 11.645 -58.54 ;
      RECT 11.505 -58.945 11.645 -58.775 ;
      RECT 11.555 -57.74 11.645 -56.732 ;
      RECT 11.505 -57.505 11.645 -57.335 ;
      RECT 11.555 -56.318 11.645 -55.31 ;
      RECT 11.505 -55.715 11.645 -55.545 ;
      RECT 11.555 -54.51 11.645 -53.502 ;
      RECT 11.505 -54.275 11.645 -54.105 ;
      RECT 11.555 -53.088 11.645 -52.08 ;
      RECT 11.505 -52.485 11.645 -52.315 ;
      RECT 11.555 -51.28 11.645 -50.272 ;
      RECT 11.505 -51.045 11.645 -50.875 ;
      RECT 11.555 -49.858 11.645 -48.85 ;
      RECT 11.505 -49.255 11.645 -49.085 ;
      RECT 11.555 -48.05 11.645 -47.042 ;
      RECT 11.505 -47.815 11.645 -47.645 ;
      RECT 11.555 -46.628 11.645 -45.62 ;
      RECT 11.505 -46.025 11.645 -45.855 ;
      RECT 11.555 -44.82 11.645 -43.812 ;
      RECT 11.505 -44.585 11.645 -44.415 ;
      RECT 11.555 -43.398 11.645 -42.39 ;
      RECT 11.505 -42.795 11.645 -42.625 ;
      RECT 11.555 -41.59 11.645 -40.582 ;
      RECT 11.505 -41.355 11.645 -41.185 ;
      RECT 11.555 -40.168 11.645 -39.16 ;
      RECT 11.505 -39.565 11.645 -39.395 ;
      RECT 11.555 -38.36 11.645 -37.352 ;
      RECT 11.505 -38.125 11.645 -37.955 ;
      RECT 11.555 -36.938 11.645 -35.93 ;
      RECT 11.505 -36.335 11.645 -36.165 ;
      RECT 11.555 -35.13 11.645 -34.122 ;
      RECT 11.505 -34.895 11.645 -34.725 ;
      RECT 11.555 -33.708 11.645 -32.7 ;
      RECT 11.505 -33.105 11.645 -32.935 ;
      RECT 11.555 -31.9 11.645 -30.892 ;
      RECT 11.505 -31.665 11.645 -31.495 ;
      RECT 11.555 -30.478 11.645 -29.47 ;
      RECT 11.505 -29.875 11.645 -29.705 ;
      RECT 11.555 -28.67 11.645 -27.662 ;
      RECT 11.505 -28.435 11.645 -28.265 ;
      RECT 11.555 -27.248 11.645 -26.24 ;
      RECT 11.505 -26.645 11.645 -26.475 ;
      RECT 11.555 -25.44 11.645 -24.432 ;
      RECT 11.505 -25.205 11.645 -25.035 ;
      RECT 11.555 -24.018 11.645 -23.01 ;
      RECT 11.505 -23.415 11.645 -23.245 ;
      RECT 11.555 -22.21 11.645 -21.202 ;
      RECT 11.505 -21.975 11.645 -21.805 ;
      RECT 11.555 -20.788 11.645 -19.78 ;
      RECT 11.505 -20.185 11.645 -20.015 ;
      RECT 11.555 -18.98 11.645 -17.972 ;
      RECT 11.505 -18.745 11.645 -18.575 ;
      RECT 11.555 -17.558 11.645 -16.55 ;
      RECT 11.505 -16.955 11.645 -16.785 ;
      RECT 11.555 -15.75 11.645 -14.742 ;
      RECT 11.505 -15.515 11.645 -15.345 ;
      RECT 11.555 -14.328 11.645 -13.32 ;
      RECT 11.505 -13.725 11.645 -13.555 ;
      RECT 11.555 -12.52 11.645 -11.512 ;
      RECT 11.505 -12.285 11.645 -12.115 ;
      RECT 11.555 -11.098 11.645 -10.09 ;
      RECT 11.505 -10.495 11.645 -10.325 ;
      RECT 11.555 -9.29 11.645 -8.282 ;
      RECT 11.505 -9.055 11.645 -8.885 ;
      RECT 11.555 -7.868 11.645 -6.86 ;
      RECT 11.505 -7.265 11.645 -7.095 ;
      RECT 11.555 -6.06 11.645 -5.052 ;
      RECT 11.505 -5.825 11.645 -5.655 ;
      RECT 11.555 -4.638 11.645 -3.63 ;
      RECT 11.505 -4.035 11.645 -3.865 ;
      RECT 11.555 -2.83 11.645 -1.822 ;
      RECT 11.505 -2.595 11.645 -2.425 ;
      RECT 11.555 -1.408 11.645 -0.4 ;
      RECT 11.505 -0.805 11.645 -0.635 ;
      RECT 11.555 0.4 11.645 1.408 ;
      RECT 11.505 0.635 11.645 0.805 ;
      RECT 11.43 -114.685 11.605 -114.515 ;
      RECT 11.505 -114.895 11.605 -114.515 ;
      RECT 10.545 -113.555 10.645 -113.09 ;
      RECT 10.91 -113.555 11.01 -113.1 ;
      RECT 10.545 -113.555 11.39 -113.385 ;
      RECT 11.155 -101.538 11.245 -100.531 ;
      RECT 11.155 -101.225 11.295 -101.055 ;
      RECT 11.155 -99.729 11.245 -98.722 ;
      RECT 11.155 -99.205 11.295 -99.035 ;
      RECT 11.155 -98.308 11.245 -97.301 ;
      RECT 11.155 -97.995 11.295 -97.825 ;
      RECT 11.155 -96.499 11.245 -95.492 ;
      RECT 11.155 -95.975 11.295 -95.805 ;
      RECT 11.155 -95.078 11.245 -94.071 ;
      RECT 11.155 -94.765 11.295 -94.595 ;
      RECT 11.155 -93.269 11.245 -92.262 ;
      RECT 11.155 -92.745 11.295 -92.575 ;
      RECT 11.155 -91.848 11.245 -90.841 ;
      RECT 11.155 -91.535 11.295 -91.365 ;
      RECT 11.155 -90.039 11.245 -89.032 ;
      RECT 11.155 -89.515 11.295 -89.345 ;
      RECT 11.155 -88.618 11.245 -87.611 ;
      RECT 11.155 -88.305 11.295 -88.135 ;
      RECT 11.155 -86.809 11.245 -85.802 ;
      RECT 11.155 -86.285 11.295 -86.115 ;
      RECT 11.155 -85.388 11.245 -84.381 ;
      RECT 11.155 -85.075 11.295 -84.905 ;
      RECT 11.155 -83.579 11.245 -82.572 ;
      RECT 11.155 -83.055 11.295 -82.885 ;
      RECT 11.155 -82.158 11.245 -81.151 ;
      RECT 11.155 -81.845 11.295 -81.675 ;
      RECT 11.155 -80.349 11.245 -79.342 ;
      RECT 11.155 -79.825 11.295 -79.655 ;
      RECT 11.155 -78.928 11.245 -77.921 ;
      RECT 11.155 -78.615 11.295 -78.445 ;
      RECT 11.155 -77.119 11.245 -76.112 ;
      RECT 11.155 -76.595 11.295 -76.425 ;
      RECT 11.155 -75.698 11.245 -74.691 ;
      RECT 11.155 -75.385 11.295 -75.215 ;
      RECT 11.155 -73.889 11.245 -72.882 ;
      RECT 11.155 -73.365 11.295 -73.195 ;
      RECT 11.155 -72.468 11.245 -71.461 ;
      RECT 11.155 -72.155 11.295 -71.985 ;
      RECT 11.155 -70.659 11.245 -69.652 ;
      RECT 11.155 -70.135 11.295 -69.965 ;
      RECT 11.155 -69.238 11.245 -68.231 ;
      RECT 11.155 -68.925 11.295 -68.755 ;
      RECT 11.155 -67.429 11.245 -66.422 ;
      RECT 11.155 -66.905 11.295 -66.735 ;
      RECT 11.155 -66.008 11.245 -65.001 ;
      RECT 11.155 -65.695 11.295 -65.525 ;
      RECT 11.155 -64.199 11.245 -63.192 ;
      RECT 11.155 -63.675 11.295 -63.505 ;
      RECT 11.155 -62.778 11.245 -61.771 ;
      RECT 11.155 -62.465 11.295 -62.295 ;
      RECT 11.155 -60.969 11.245 -59.962 ;
      RECT 11.155 -60.445 11.295 -60.275 ;
      RECT 11.155 -59.548 11.245 -58.541 ;
      RECT 11.155 -59.235 11.295 -59.065 ;
      RECT 11.155 -57.739 11.245 -56.732 ;
      RECT 11.155 -57.215 11.295 -57.045 ;
      RECT 11.155 -56.318 11.245 -55.311 ;
      RECT 11.155 -56.005 11.295 -55.835 ;
      RECT 11.155 -54.509 11.245 -53.502 ;
      RECT 11.155 -53.985 11.295 -53.815 ;
      RECT 11.155 -53.088 11.245 -52.081 ;
      RECT 11.155 -52.775 11.295 -52.605 ;
      RECT 11.155 -51.279 11.245 -50.272 ;
      RECT 11.155 -50.755 11.295 -50.585 ;
      RECT 11.155 -49.858 11.245 -48.851 ;
      RECT 11.155 -49.545 11.295 -49.375 ;
      RECT 11.155 -48.049 11.245 -47.042 ;
      RECT 11.155 -47.525 11.295 -47.355 ;
      RECT 11.155 -46.628 11.245 -45.621 ;
      RECT 11.155 -46.315 11.295 -46.145 ;
      RECT 11.155 -44.819 11.245 -43.812 ;
      RECT 11.155 -44.295 11.295 -44.125 ;
      RECT 11.155 -43.398 11.245 -42.391 ;
      RECT 11.155 -43.085 11.295 -42.915 ;
      RECT 11.155 -41.589 11.245 -40.582 ;
      RECT 11.155 -41.065 11.295 -40.895 ;
      RECT 11.155 -40.168 11.245 -39.161 ;
      RECT 11.155 -39.855 11.295 -39.685 ;
      RECT 11.155 -38.359 11.245 -37.352 ;
      RECT 11.155 -37.835 11.295 -37.665 ;
      RECT 11.155 -36.938 11.245 -35.931 ;
      RECT 11.155 -36.625 11.295 -36.455 ;
      RECT 11.155 -35.129 11.245 -34.122 ;
      RECT 11.155 -34.605 11.295 -34.435 ;
      RECT 11.155 -33.708 11.245 -32.701 ;
      RECT 11.155 -33.395 11.295 -33.225 ;
      RECT 11.155 -31.899 11.245 -30.892 ;
      RECT 11.155 -31.375 11.295 -31.205 ;
      RECT 11.155 -30.478 11.245 -29.471 ;
      RECT 11.155 -30.165 11.295 -29.995 ;
      RECT 11.155 -28.669 11.245 -27.662 ;
      RECT 11.155 -28.145 11.295 -27.975 ;
      RECT 11.155 -27.248 11.245 -26.241 ;
      RECT 11.155 -26.935 11.295 -26.765 ;
      RECT 11.155 -25.439 11.245 -24.432 ;
      RECT 11.155 -24.915 11.295 -24.745 ;
      RECT 11.155 -24.018 11.245 -23.011 ;
      RECT 11.155 -23.705 11.295 -23.535 ;
      RECT 11.155 -22.209 11.245 -21.202 ;
      RECT 11.155 -21.685 11.295 -21.515 ;
      RECT 11.155 -20.788 11.245 -19.781 ;
      RECT 11.155 -20.475 11.295 -20.305 ;
      RECT 11.155 -18.979 11.245 -17.972 ;
      RECT 11.155 -18.455 11.295 -18.285 ;
      RECT 11.155 -17.558 11.245 -16.551 ;
      RECT 11.155 -17.245 11.295 -17.075 ;
      RECT 11.155 -15.749 11.245 -14.742 ;
      RECT 11.155 -15.225 11.295 -15.055 ;
      RECT 11.155 -14.328 11.245 -13.321 ;
      RECT 11.155 -14.015 11.295 -13.845 ;
      RECT 11.155 -12.519 11.245 -11.512 ;
      RECT 11.155 -11.995 11.295 -11.825 ;
      RECT 11.155 -11.098 11.245 -10.091 ;
      RECT 11.155 -10.785 11.295 -10.615 ;
      RECT 11.155 -9.289 11.245 -8.282 ;
      RECT 11.155 -8.765 11.295 -8.595 ;
      RECT 11.155 -7.868 11.245 -6.861 ;
      RECT 11.155 -7.555 11.295 -7.385 ;
      RECT 11.155 -6.059 11.245 -5.052 ;
      RECT 11.155 -5.535 11.295 -5.365 ;
      RECT 11.155 -4.638 11.245 -3.631 ;
      RECT 11.155 -4.325 11.295 -4.155 ;
      RECT 11.155 -2.829 11.245 -1.822 ;
      RECT 11.155 -2.305 11.295 -2.135 ;
      RECT 11.155 -1.408 11.245 -0.401 ;
      RECT 11.155 -1.095 11.295 -0.925 ;
      RECT 11.155 0.401 11.245 1.408 ;
      RECT 11.155 0.925 11.295 1.095 ;
      RECT 10.84 -114.685 11.01 -114.515 ;
      RECT 10.91 -114.895 11.01 -114.515 ;
      RECT 10.355 -101.538 10.445 -100.53 ;
      RECT 10.305 -100.935 10.445 -100.765 ;
      RECT 10.355 -99.73 10.445 -98.722 ;
      RECT 10.305 -99.495 10.445 -99.325 ;
      RECT 10.355 -98.308 10.445 -97.3 ;
      RECT 10.305 -97.705 10.445 -97.535 ;
      RECT 10.355 -96.5 10.445 -95.492 ;
      RECT 10.305 -96.265 10.445 -96.095 ;
      RECT 10.355 -95.078 10.445 -94.07 ;
      RECT 10.305 -94.475 10.445 -94.305 ;
      RECT 10.355 -93.27 10.445 -92.262 ;
      RECT 10.305 -93.035 10.445 -92.865 ;
      RECT 10.355 -91.848 10.445 -90.84 ;
      RECT 10.305 -91.245 10.445 -91.075 ;
      RECT 10.355 -90.04 10.445 -89.032 ;
      RECT 10.305 -89.805 10.445 -89.635 ;
      RECT 10.355 -88.618 10.445 -87.61 ;
      RECT 10.305 -88.015 10.445 -87.845 ;
      RECT 10.355 -86.81 10.445 -85.802 ;
      RECT 10.305 -86.575 10.445 -86.405 ;
      RECT 10.355 -85.388 10.445 -84.38 ;
      RECT 10.305 -84.785 10.445 -84.615 ;
      RECT 10.355 -83.58 10.445 -82.572 ;
      RECT 10.305 -83.345 10.445 -83.175 ;
      RECT 10.355 -82.158 10.445 -81.15 ;
      RECT 10.305 -81.555 10.445 -81.385 ;
      RECT 10.355 -80.35 10.445 -79.342 ;
      RECT 10.305 -80.115 10.445 -79.945 ;
      RECT 10.355 -78.928 10.445 -77.92 ;
      RECT 10.305 -78.325 10.445 -78.155 ;
      RECT 10.355 -77.12 10.445 -76.112 ;
      RECT 10.305 -76.885 10.445 -76.715 ;
      RECT 10.355 -75.698 10.445 -74.69 ;
      RECT 10.305 -75.095 10.445 -74.925 ;
      RECT 10.355 -73.89 10.445 -72.882 ;
      RECT 10.305 -73.655 10.445 -73.485 ;
      RECT 10.355 -72.468 10.445 -71.46 ;
      RECT 10.305 -71.865 10.445 -71.695 ;
      RECT 10.355 -70.66 10.445 -69.652 ;
      RECT 10.305 -70.425 10.445 -70.255 ;
      RECT 10.355 -69.238 10.445 -68.23 ;
      RECT 10.305 -68.635 10.445 -68.465 ;
      RECT 10.355 -67.43 10.445 -66.422 ;
      RECT 10.305 -67.195 10.445 -67.025 ;
      RECT 10.355 -66.008 10.445 -65 ;
      RECT 10.305 -65.405 10.445 -65.235 ;
      RECT 10.355 -64.2 10.445 -63.192 ;
      RECT 10.305 -63.965 10.445 -63.795 ;
      RECT 10.355 -62.778 10.445 -61.77 ;
      RECT 10.305 -62.175 10.445 -62.005 ;
      RECT 10.355 -60.97 10.445 -59.962 ;
      RECT 10.305 -60.735 10.445 -60.565 ;
      RECT 10.355 -59.548 10.445 -58.54 ;
      RECT 10.305 -58.945 10.445 -58.775 ;
      RECT 10.355 -57.74 10.445 -56.732 ;
      RECT 10.305 -57.505 10.445 -57.335 ;
      RECT 10.355 -56.318 10.445 -55.31 ;
      RECT 10.305 -55.715 10.445 -55.545 ;
      RECT 10.355 -54.51 10.445 -53.502 ;
      RECT 10.305 -54.275 10.445 -54.105 ;
      RECT 10.355 -53.088 10.445 -52.08 ;
      RECT 10.305 -52.485 10.445 -52.315 ;
      RECT 10.355 -51.28 10.445 -50.272 ;
      RECT 10.305 -51.045 10.445 -50.875 ;
      RECT 10.355 -49.858 10.445 -48.85 ;
      RECT 10.305 -49.255 10.445 -49.085 ;
      RECT 10.355 -48.05 10.445 -47.042 ;
      RECT 10.305 -47.815 10.445 -47.645 ;
      RECT 10.355 -46.628 10.445 -45.62 ;
      RECT 10.305 -46.025 10.445 -45.855 ;
      RECT 10.355 -44.82 10.445 -43.812 ;
      RECT 10.305 -44.585 10.445 -44.415 ;
      RECT 10.355 -43.398 10.445 -42.39 ;
      RECT 10.305 -42.795 10.445 -42.625 ;
      RECT 10.355 -41.59 10.445 -40.582 ;
      RECT 10.305 -41.355 10.445 -41.185 ;
      RECT 10.355 -40.168 10.445 -39.16 ;
      RECT 10.305 -39.565 10.445 -39.395 ;
      RECT 10.355 -38.36 10.445 -37.352 ;
      RECT 10.305 -38.125 10.445 -37.955 ;
      RECT 10.355 -36.938 10.445 -35.93 ;
      RECT 10.305 -36.335 10.445 -36.165 ;
      RECT 10.355 -35.13 10.445 -34.122 ;
      RECT 10.305 -34.895 10.445 -34.725 ;
      RECT 10.355 -33.708 10.445 -32.7 ;
      RECT 10.305 -33.105 10.445 -32.935 ;
      RECT 10.355 -31.9 10.445 -30.892 ;
      RECT 10.305 -31.665 10.445 -31.495 ;
      RECT 10.355 -30.478 10.445 -29.47 ;
      RECT 10.305 -29.875 10.445 -29.705 ;
      RECT 10.355 -28.67 10.445 -27.662 ;
      RECT 10.305 -28.435 10.445 -28.265 ;
      RECT 10.355 -27.248 10.445 -26.24 ;
      RECT 10.305 -26.645 10.445 -26.475 ;
      RECT 10.355 -25.44 10.445 -24.432 ;
      RECT 10.305 -25.205 10.445 -25.035 ;
      RECT 10.355 -24.018 10.445 -23.01 ;
      RECT 10.305 -23.415 10.445 -23.245 ;
      RECT 10.355 -22.21 10.445 -21.202 ;
      RECT 10.305 -21.975 10.445 -21.805 ;
      RECT 10.355 -20.788 10.445 -19.78 ;
      RECT 10.305 -20.185 10.445 -20.015 ;
      RECT 10.355 -18.98 10.445 -17.972 ;
      RECT 10.305 -18.745 10.445 -18.575 ;
      RECT 10.355 -17.558 10.445 -16.55 ;
      RECT 10.305 -16.955 10.445 -16.785 ;
      RECT 10.355 -15.75 10.445 -14.742 ;
      RECT 10.305 -15.515 10.445 -15.345 ;
      RECT 10.355 -14.328 10.445 -13.32 ;
      RECT 10.305 -13.725 10.445 -13.555 ;
      RECT 10.355 -12.52 10.445 -11.512 ;
      RECT 10.305 -12.285 10.445 -12.115 ;
      RECT 10.355 -11.098 10.445 -10.09 ;
      RECT 10.305 -10.495 10.445 -10.325 ;
      RECT 10.355 -9.29 10.445 -8.282 ;
      RECT 10.305 -9.055 10.445 -8.885 ;
      RECT 10.355 -7.868 10.445 -6.86 ;
      RECT 10.305 -7.265 10.445 -7.095 ;
      RECT 10.355 -6.06 10.445 -5.052 ;
      RECT 10.305 -5.825 10.445 -5.655 ;
      RECT 10.355 -4.638 10.445 -3.63 ;
      RECT 10.305 -4.035 10.445 -3.865 ;
      RECT 10.355 -2.83 10.445 -1.822 ;
      RECT 10.305 -2.595 10.445 -2.425 ;
      RECT 10.355 -1.408 10.445 -0.4 ;
      RECT 10.305 -0.805 10.445 -0.635 ;
      RECT 10.355 0.4 10.445 1.408 ;
      RECT 10.305 0.635 10.445 0.805 ;
      RECT 9.955 -101.538 10.045 -100.531 ;
      RECT 9.955 -101.225 10.095 -101.055 ;
      RECT 9.955 -99.729 10.045 -98.722 ;
      RECT 9.955 -99.205 10.095 -99.035 ;
      RECT 9.955 -98.308 10.045 -97.301 ;
      RECT 9.955 -97.995 10.095 -97.825 ;
      RECT 9.955 -96.499 10.045 -95.492 ;
      RECT 9.955 -95.975 10.095 -95.805 ;
      RECT 9.955 -95.078 10.045 -94.071 ;
      RECT 9.955 -94.765 10.095 -94.595 ;
      RECT 9.955 -93.269 10.045 -92.262 ;
      RECT 9.955 -92.745 10.095 -92.575 ;
      RECT 9.955 -91.848 10.045 -90.841 ;
      RECT 9.955 -91.535 10.095 -91.365 ;
      RECT 9.955 -90.039 10.045 -89.032 ;
      RECT 9.955 -89.515 10.095 -89.345 ;
      RECT 9.955 -88.618 10.045 -87.611 ;
      RECT 9.955 -88.305 10.095 -88.135 ;
      RECT 9.955 -86.809 10.045 -85.802 ;
      RECT 9.955 -86.285 10.095 -86.115 ;
      RECT 9.955 -85.388 10.045 -84.381 ;
      RECT 9.955 -85.075 10.095 -84.905 ;
      RECT 9.955 -83.579 10.045 -82.572 ;
      RECT 9.955 -83.055 10.095 -82.885 ;
      RECT 9.955 -82.158 10.045 -81.151 ;
      RECT 9.955 -81.845 10.095 -81.675 ;
      RECT 9.955 -80.349 10.045 -79.342 ;
      RECT 9.955 -79.825 10.095 -79.655 ;
      RECT 9.955 -78.928 10.045 -77.921 ;
      RECT 9.955 -78.615 10.095 -78.445 ;
      RECT 9.955 -77.119 10.045 -76.112 ;
      RECT 9.955 -76.595 10.095 -76.425 ;
      RECT 9.955 -75.698 10.045 -74.691 ;
      RECT 9.955 -75.385 10.095 -75.215 ;
      RECT 9.955 -73.889 10.045 -72.882 ;
      RECT 9.955 -73.365 10.095 -73.195 ;
      RECT 9.955 -72.468 10.045 -71.461 ;
      RECT 9.955 -72.155 10.095 -71.985 ;
      RECT 9.955 -70.659 10.045 -69.652 ;
      RECT 9.955 -70.135 10.095 -69.965 ;
      RECT 9.955 -69.238 10.045 -68.231 ;
      RECT 9.955 -68.925 10.095 -68.755 ;
      RECT 9.955 -67.429 10.045 -66.422 ;
      RECT 9.955 -66.905 10.095 -66.735 ;
      RECT 9.955 -66.008 10.045 -65.001 ;
      RECT 9.955 -65.695 10.095 -65.525 ;
      RECT 9.955 -64.199 10.045 -63.192 ;
      RECT 9.955 -63.675 10.095 -63.505 ;
      RECT 9.955 -62.778 10.045 -61.771 ;
      RECT 9.955 -62.465 10.095 -62.295 ;
      RECT 9.955 -60.969 10.045 -59.962 ;
      RECT 9.955 -60.445 10.095 -60.275 ;
      RECT 9.955 -59.548 10.045 -58.541 ;
      RECT 9.955 -59.235 10.095 -59.065 ;
      RECT 9.955 -57.739 10.045 -56.732 ;
      RECT 9.955 -57.215 10.095 -57.045 ;
      RECT 9.955 -56.318 10.045 -55.311 ;
      RECT 9.955 -56.005 10.095 -55.835 ;
      RECT 9.955 -54.509 10.045 -53.502 ;
      RECT 9.955 -53.985 10.095 -53.815 ;
      RECT 9.955 -53.088 10.045 -52.081 ;
      RECT 9.955 -52.775 10.095 -52.605 ;
      RECT 9.955 -51.279 10.045 -50.272 ;
      RECT 9.955 -50.755 10.095 -50.585 ;
      RECT 9.955 -49.858 10.045 -48.851 ;
      RECT 9.955 -49.545 10.095 -49.375 ;
      RECT 9.955 -48.049 10.045 -47.042 ;
      RECT 9.955 -47.525 10.095 -47.355 ;
      RECT 9.955 -46.628 10.045 -45.621 ;
      RECT 9.955 -46.315 10.095 -46.145 ;
      RECT 9.955 -44.819 10.045 -43.812 ;
      RECT 9.955 -44.295 10.095 -44.125 ;
      RECT 9.955 -43.398 10.045 -42.391 ;
      RECT 9.955 -43.085 10.095 -42.915 ;
      RECT 9.955 -41.589 10.045 -40.582 ;
      RECT 9.955 -41.065 10.095 -40.895 ;
      RECT 9.955 -40.168 10.045 -39.161 ;
      RECT 9.955 -39.855 10.095 -39.685 ;
      RECT 9.955 -38.359 10.045 -37.352 ;
      RECT 9.955 -37.835 10.095 -37.665 ;
      RECT 9.955 -36.938 10.045 -35.931 ;
      RECT 9.955 -36.625 10.095 -36.455 ;
      RECT 9.955 -35.129 10.045 -34.122 ;
      RECT 9.955 -34.605 10.095 -34.435 ;
      RECT 9.955 -33.708 10.045 -32.701 ;
      RECT 9.955 -33.395 10.095 -33.225 ;
      RECT 9.955 -31.899 10.045 -30.892 ;
      RECT 9.955 -31.375 10.095 -31.205 ;
      RECT 9.955 -30.478 10.045 -29.471 ;
      RECT 9.955 -30.165 10.095 -29.995 ;
      RECT 9.955 -28.669 10.045 -27.662 ;
      RECT 9.955 -28.145 10.095 -27.975 ;
      RECT 9.955 -27.248 10.045 -26.241 ;
      RECT 9.955 -26.935 10.095 -26.765 ;
      RECT 9.955 -25.439 10.045 -24.432 ;
      RECT 9.955 -24.915 10.095 -24.745 ;
      RECT 9.955 -24.018 10.045 -23.011 ;
      RECT 9.955 -23.705 10.095 -23.535 ;
      RECT 9.955 -22.209 10.045 -21.202 ;
      RECT 9.955 -21.685 10.095 -21.515 ;
      RECT 9.955 -20.788 10.045 -19.781 ;
      RECT 9.955 -20.475 10.095 -20.305 ;
      RECT 9.955 -18.979 10.045 -17.972 ;
      RECT 9.955 -18.455 10.095 -18.285 ;
      RECT 9.955 -17.558 10.045 -16.551 ;
      RECT 9.955 -17.245 10.095 -17.075 ;
      RECT 9.955 -15.749 10.045 -14.742 ;
      RECT 9.955 -15.225 10.095 -15.055 ;
      RECT 9.955 -14.328 10.045 -13.321 ;
      RECT 9.955 -14.015 10.095 -13.845 ;
      RECT 9.955 -12.519 10.045 -11.512 ;
      RECT 9.955 -11.995 10.095 -11.825 ;
      RECT 9.955 -11.098 10.045 -10.091 ;
      RECT 9.955 -10.785 10.095 -10.615 ;
      RECT 9.955 -9.289 10.045 -8.282 ;
      RECT 9.955 -8.765 10.095 -8.595 ;
      RECT 9.955 -7.868 10.045 -6.861 ;
      RECT 9.955 -7.555 10.095 -7.385 ;
      RECT 9.955 -6.059 10.045 -5.052 ;
      RECT 9.955 -5.535 10.095 -5.365 ;
      RECT 9.955 -4.638 10.045 -3.631 ;
      RECT 9.955 -4.325 10.095 -4.155 ;
      RECT 9.955 -2.829 10.045 -1.822 ;
      RECT 9.955 -2.305 10.095 -2.135 ;
      RECT 9.955 -1.408 10.045 -0.401 ;
      RECT 9.955 -1.095 10.095 -0.925 ;
      RECT 9.955 0.401 10.045 1.408 ;
      RECT 9.955 0.925 10.095 1.095 ;
      RECT 5.785 -108.935 9.565 -108.815 ;
      RECT 7.105 -109.475 7.205 -108.815 ;
      RECT 6.545 -109.475 6.645 -108.815 ;
      RECT 5.985 -109.475 6.085 -108.815 ;
      RECT 9.155 -101.538 9.245 -100.53 ;
      RECT 9.105 -100.935 9.245 -100.765 ;
      RECT 9.155 -99.73 9.245 -98.722 ;
      RECT 9.105 -99.495 9.245 -99.325 ;
      RECT 9.155 -98.308 9.245 -97.3 ;
      RECT 9.105 -97.705 9.245 -97.535 ;
      RECT 9.155 -96.5 9.245 -95.492 ;
      RECT 9.105 -96.265 9.245 -96.095 ;
      RECT 9.155 -95.078 9.245 -94.07 ;
      RECT 9.105 -94.475 9.245 -94.305 ;
      RECT 9.155 -93.27 9.245 -92.262 ;
      RECT 9.105 -93.035 9.245 -92.865 ;
      RECT 9.155 -91.848 9.245 -90.84 ;
      RECT 9.105 -91.245 9.245 -91.075 ;
      RECT 9.155 -90.04 9.245 -89.032 ;
      RECT 9.105 -89.805 9.245 -89.635 ;
      RECT 9.155 -88.618 9.245 -87.61 ;
      RECT 9.105 -88.015 9.245 -87.845 ;
      RECT 9.155 -86.81 9.245 -85.802 ;
      RECT 9.105 -86.575 9.245 -86.405 ;
      RECT 9.155 -85.388 9.245 -84.38 ;
      RECT 9.105 -84.785 9.245 -84.615 ;
      RECT 9.155 -83.58 9.245 -82.572 ;
      RECT 9.105 -83.345 9.245 -83.175 ;
      RECT 9.155 -82.158 9.245 -81.15 ;
      RECT 9.105 -81.555 9.245 -81.385 ;
      RECT 9.155 -80.35 9.245 -79.342 ;
      RECT 9.105 -80.115 9.245 -79.945 ;
      RECT 9.155 -78.928 9.245 -77.92 ;
      RECT 9.105 -78.325 9.245 -78.155 ;
      RECT 9.155 -77.12 9.245 -76.112 ;
      RECT 9.105 -76.885 9.245 -76.715 ;
      RECT 9.155 -75.698 9.245 -74.69 ;
      RECT 9.105 -75.095 9.245 -74.925 ;
      RECT 9.155 -73.89 9.245 -72.882 ;
      RECT 9.105 -73.655 9.245 -73.485 ;
      RECT 9.155 -72.468 9.245 -71.46 ;
      RECT 9.105 -71.865 9.245 -71.695 ;
      RECT 9.155 -70.66 9.245 -69.652 ;
      RECT 9.105 -70.425 9.245 -70.255 ;
      RECT 9.155 -69.238 9.245 -68.23 ;
      RECT 9.105 -68.635 9.245 -68.465 ;
      RECT 9.155 -67.43 9.245 -66.422 ;
      RECT 9.105 -67.195 9.245 -67.025 ;
      RECT 9.155 -66.008 9.245 -65 ;
      RECT 9.105 -65.405 9.245 -65.235 ;
      RECT 9.155 -64.2 9.245 -63.192 ;
      RECT 9.105 -63.965 9.245 -63.795 ;
      RECT 9.155 -62.778 9.245 -61.77 ;
      RECT 9.105 -62.175 9.245 -62.005 ;
      RECT 9.155 -60.97 9.245 -59.962 ;
      RECT 9.105 -60.735 9.245 -60.565 ;
      RECT 9.155 -59.548 9.245 -58.54 ;
      RECT 9.105 -58.945 9.245 -58.775 ;
      RECT 9.155 -57.74 9.245 -56.732 ;
      RECT 9.105 -57.505 9.245 -57.335 ;
      RECT 9.155 -56.318 9.245 -55.31 ;
      RECT 9.105 -55.715 9.245 -55.545 ;
      RECT 9.155 -54.51 9.245 -53.502 ;
      RECT 9.105 -54.275 9.245 -54.105 ;
      RECT 9.155 -53.088 9.245 -52.08 ;
      RECT 9.105 -52.485 9.245 -52.315 ;
      RECT 9.155 -51.28 9.245 -50.272 ;
      RECT 9.105 -51.045 9.245 -50.875 ;
      RECT 9.155 -49.858 9.245 -48.85 ;
      RECT 9.105 -49.255 9.245 -49.085 ;
      RECT 9.155 -48.05 9.245 -47.042 ;
      RECT 9.105 -47.815 9.245 -47.645 ;
      RECT 9.155 -46.628 9.245 -45.62 ;
      RECT 9.105 -46.025 9.245 -45.855 ;
      RECT 9.155 -44.82 9.245 -43.812 ;
      RECT 9.105 -44.585 9.245 -44.415 ;
      RECT 9.155 -43.398 9.245 -42.39 ;
      RECT 9.105 -42.795 9.245 -42.625 ;
      RECT 9.155 -41.59 9.245 -40.582 ;
      RECT 9.105 -41.355 9.245 -41.185 ;
      RECT 9.155 -40.168 9.245 -39.16 ;
      RECT 9.105 -39.565 9.245 -39.395 ;
      RECT 9.155 -38.36 9.245 -37.352 ;
      RECT 9.105 -38.125 9.245 -37.955 ;
      RECT 9.155 -36.938 9.245 -35.93 ;
      RECT 9.105 -36.335 9.245 -36.165 ;
      RECT 9.155 -35.13 9.245 -34.122 ;
      RECT 9.105 -34.895 9.245 -34.725 ;
      RECT 9.155 -33.708 9.245 -32.7 ;
      RECT 9.105 -33.105 9.245 -32.935 ;
      RECT 9.155 -31.9 9.245 -30.892 ;
      RECT 9.105 -31.665 9.245 -31.495 ;
      RECT 9.155 -30.478 9.245 -29.47 ;
      RECT 9.105 -29.875 9.245 -29.705 ;
      RECT 9.155 -28.67 9.245 -27.662 ;
      RECT 9.105 -28.435 9.245 -28.265 ;
      RECT 9.155 -27.248 9.245 -26.24 ;
      RECT 9.105 -26.645 9.245 -26.475 ;
      RECT 9.155 -25.44 9.245 -24.432 ;
      RECT 9.105 -25.205 9.245 -25.035 ;
      RECT 9.155 -24.018 9.245 -23.01 ;
      RECT 9.105 -23.415 9.245 -23.245 ;
      RECT 9.155 -22.21 9.245 -21.202 ;
      RECT 9.105 -21.975 9.245 -21.805 ;
      RECT 9.155 -20.788 9.245 -19.78 ;
      RECT 9.105 -20.185 9.245 -20.015 ;
      RECT 9.155 -18.98 9.245 -17.972 ;
      RECT 9.105 -18.745 9.245 -18.575 ;
      RECT 9.155 -17.558 9.245 -16.55 ;
      RECT 9.105 -16.955 9.245 -16.785 ;
      RECT 9.155 -15.75 9.245 -14.742 ;
      RECT 9.105 -15.515 9.245 -15.345 ;
      RECT 9.155 -14.328 9.245 -13.32 ;
      RECT 9.105 -13.725 9.245 -13.555 ;
      RECT 9.155 -12.52 9.245 -11.512 ;
      RECT 9.105 -12.285 9.245 -12.115 ;
      RECT 9.155 -11.098 9.245 -10.09 ;
      RECT 9.105 -10.495 9.245 -10.325 ;
      RECT 9.155 -9.29 9.245 -8.282 ;
      RECT 9.105 -9.055 9.245 -8.885 ;
      RECT 9.155 -7.868 9.245 -6.86 ;
      RECT 9.105 -7.265 9.245 -7.095 ;
      RECT 9.155 -6.06 9.245 -5.052 ;
      RECT 9.105 -5.825 9.245 -5.655 ;
      RECT 9.155 -4.638 9.245 -3.63 ;
      RECT 9.105 -4.035 9.245 -3.865 ;
      RECT 9.155 -2.83 9.245 -1.822 ;
      RECT 9.105 -2.595 9.245 -2.425 ;
      RECT 9.155 -1.408 9.245 -0.4 ;
      RECT 9.105 -0.805 9.245 -0.635 ;
      RECT 9.155 0.4 9.245 1.408 ;
      RECT 9.105 0.635 9.245 0.805 ;
      RECT 7.725 -111.685 9.205 -111.585 ;
      RECT 7.725 -112.195 7.825 -111.585 ;
      RECT 7.945 -109.15 9.205 -109.05 ;
      RECT 9.105 -109.475 9.205 -109.05 ;
      RECT 8.545 -109.475 8.645 -109.05 ;
      RECT 7.985 -109.475 8.085 -109.05 ;
      RECT 8.755 -101.538 8.845 -100.531 ;
      RECT 8.755 -101.225 8.895 -101.055 ;
      RECT 8.755 -99.729 8.845 -98.722 ;
      RECT 8.755 -99.205 8.895 -99.035 ;
      RECT 8.755 -98.308 8.845 -97.301 ;
      RECT 8.755 -97.995 8.895 -97.825 ;
      RECT 8.755 -96.499 8.845 -95.492 ;
      RECT 8.755 -95.975 8.895 -95.805 ;
      RECT 8.755 -95.078 8.845 -94.071 ;
      RECT 8.755 -94.765 8.895 -94.595 ;
      RECT 8.755 -93.269 8.845 -92.262 ;
      RECT 8.755 -92.745 8.895 -92.575 ;
      RECT 8.755 -91.848 8.845 -90.841 ;
      RECT 8.755 -91.535 8.895 -91.365 ;
      RECT 8.755 -90.039 8.845 -89.032 ;
      RECT 8.755 -89.515 8.895 -89.345 ;
      RECT 8.755 -88.618 8.845 -87.611 ;
      RECT 8.755 -88.305 8.895 -88.135 ;
      RECT 8.755 -86.809 8.845 -85.802 ;
      RECT 8.755 -86.285 8.895 -86.115 ;
      RECT 8.755 -85.388 8.845 -84.381 ;
      RECT 8.755 -85.075 8.895 -84.905 ;
      RECT 8.755 -83.579 8.845 -82.572 ;
      RECT 8.755 -83.055 8.895 -82.885 ;
      RECT 8.755 -82.158 8.845 -81.151 ;
      RECT 8.755 -81.845 8.895 -81.675 ;
      RECT 8.755 -80.349 8.845 -79.342 ;
      RECT 8.755 -79.825 8.895 -79.655 ;
      RECT 8.755 -78.928 8.845 -77.921 ;
      RECT 8.755 -78.615 8.895 -78.445 ;
      RECT 8.755 -77.119 8.845 -76.112 ;
      RECT 8.755 -76.595 8.895 -76.425 ;
      RECT 8.755 -75.698 8.845 -74.691 ;
      RECT 8.755 -75.385 8.895 -75.215 ;
      RECT 8.755 -73.889 8.845 -72.882 ;
      RECT 8.755 -73.365 8.895 -73.195 ;
      RECT 8.755 -72.468 8.845 -71.461 ;
      RECT 8.755 -72.155 8.895 -71.985 ;
      RECT 8.755 -70.659 8.845 -69.652 ;
      RECT 8.755 -70.135 8.895 -69.965 ;
      RECT 8.755 -69.238 8.845 -68.231 ;
      RECT 8.755 -68.925 8.895 -68.755 ;
      RECT 8.755 -67.429 8.845 -66.422 ;
      RECT 8.755 -66.905 8.895 -66.735 ;
      RECT 8.755 -66.008 8.845 -65.001 ;
      RECT 8.755 -65.695 8.895 -65.525 ;
      RECT 8.755 -64.199 8.845 -63.192 ;
      RECT 8.755 -63.675 8.895 -63.505 ;
      RECT 8.755 -62.778 8.845 -61.771 ;
      RECT 8.755 -62.465 8.895 -62.295 ;
      RECT 8.755 -60.969 8.845 -59.962 ;
      RECT 8.755 -60.445 8.895 -60.275 ;
      RECT 8.755 -59.548 8.845 -58.541 ;
      RECT 8.755 -59.235 8.895 -59.065 ;
      RECT 8.755 -57.739 8.845 -56.732 ;
      RECT 8.755 -57.215 8.895 -57.045 ;
      RECT 8.755 -56.318 8.845 -55.311 ;
      RECT 8.755 -56.005 8.895 -55.835 ;
      RECT 8.755 -54.509 8.845 -53.502 ;
      RECT 8.755 -53.985 8.895 -53.815 ;
      RECT 8.755 -53.088 8.845 -52.081 ;
      RECT 8.755 -52.775 8.895 -52.605 ;
      RECT 8.755 -51.279 8.845 -50.272 ;
      RECT 8.755 -50.755 8.895 -50.585 ;
      RECT 8.755 -49.858 8.845 -48.851 ;
      RECT 8.755 -49.545 8.895 -49.375 ;
      RECT 8.755 -48.049 8.845 -47.042 ;
      RECT 8.755 -47.525 8.895 -47.355 ;
      RECT 8.755 -46.628 8.845 -45.621 ;
      RECT 8.755 -46.315 8.895 -46.145 ;
      RECT 8.755 -44.819 8.845 -43.812 ;
      RECT 8.755 -44.295 8.895 -44.125 ;
      RECT 8.755 -43.398 8.845 -42.391 ;
      RECT 8.755 -43.085 8.895 -42.915 ;
      RECT 8.755 -41.589 8.845 -40.582 ;
      RECT 8.755 -41.065 8.895 -40.895 ;
      RECT 8.755 -40.168 8.845 -39.161 ;
      RECT 8.755 -39.855 8.895 -39.685 ;
      RECT 8.755 -38.359 8.845 -37.352 ;
      RECT 8.755 -37.835 8.895 -37.665 ;
      RECT 8.755 -36.938 8.845 -35.931 ;
      RECT 8.755 -36.625 8.895 -36.455 ;
      RECT 8.755 -35.129 8.845 -34.122 ;
      RECT 8.755 -34.605 8.895 -34.435 ;
      RECT 8.755 -33.708 8.845 -32.701 ;
      RECT 8.755 -33.395 8.895 -33.225 ;
      RECT 8.755 -31.899 8.845 -30.892 ;
      RECT 8.755 -31.375 8.895 -31.205 ;
      RECT 8.755 -30.478 8.845 -29.471 ;
      RECT 8.755 -30.165 8.895 -29.995 ;
      RECT 8.755 -28.669 8.845 -27.662 ;
      RECT 8.755 -28.145 8.895 -27.975 ;
      RECT 8.755 -27.248 8.845 -26.241 ;
      RECT 8.755 -26.935 8.895 -26.765 ;
      RECT 8.755 -25.439 8.845 -24.432 ;
      RECT 8.755 -24.915 8.895 -24.745 ;
      RECT 8.755 -24.018 8.845 -23.011 ;
      RECT 8.755 -23.705 8.895 -23.535 ;
      RECT 8.755 -22.209 8.845 -21.202 ;
      RECT 8.755 -21.685 8.895 -21.515 ;
      RECT 8.755 -20.788 8.845 -19.781 ;
      RECT 8.755 -20.475 8.895 -20.305 ;
      RECT 8.755 -18.979 8.845 -17.972 ;
      RECT 8.755 -18.455 8.895 -18.285 ;
      RECT 8.755 -17.558 8.845 -16.551 ;
      RECT 8.755 -17.245 8.895 -17.075 ;
      RECT 8.755 -15.749 8.845 -14.742 ;
      RECT 8.755 -15.225 8.895 -15.055 ;
      RECT 8.755 -14.328 8.845 -13.321 ;
      RECT 8.755 -14.015 8.895 -13.845 ;
      RECT 8.755 -12.519 8.845 -11.512 ;
      RECT 8.755 -11.995 8.895 -11.825 ;
      RECT 8.755 -11.098 8.845 -10.091 ;
      RECT 8.755 -10.785 8.895 -10.615 ;
      RECT 8.755 -9.289 8.845 -8.282 ;
      RECT 8.755 -8.765 8.895 -8.595 ;
      RECT 8.755 -7.868 8.845 -6.861 ;
      RECT 8.755 -7.555 8.895 -7.385 ;
      RECT 8.755 -6.059 8.845 -5.052 ;
      RECT 8.755 -5.535 8.895 -5.365 ;
      RECT 8.755 -4.638 8.845 -3.631 ;
      RECT 8.755 -4.325 8.895 -4.155 ;
      RECT 8.755 -2.829 8.845 -1.822 ;
      RECT 8.755 -2.305 8.895 -2.135 ;
      RECT 8.755 -1.408 8.845 -0.401 ;
      RECT 8.755 -1.095 8.895 -0.925 ;
      RECT 8.755 0.401 8.845 1.408 ;
      RECT 8.755 0.925 8.895 1.095 ;
      RECT 8.085 -111.495 8.255 -111.385 ;
      RECT 4.935 -111.495 8.255 -111.395 ;
      RECT 7.955 -101.538 8.045 -100.53 ;
      RECT 7.905 -100.935 8.045 -100.765 ;
      RECT 7.955 -99.73 8.045 -98.722 ;
      RECT 7.905 -99.495 8.045 -99.325 ;
      RECT 7.955 -98.308 8.045 -97.3 ;
      RECT 7.905 -97.705 8.045 -97.535 ;
      RECT 7.955 -96.5 8.045 -95.492 ;
      RECT 7.905 -96.265 8.045 -96.095 ;
      RECT 7.955 -95.078 8.045 -94.07 ;
      RECT 7.905 -94.475 8.045 -94.305 ;
      RECT 7.955 -93.27 8.045 -92.262 ;
      RECT 7.905 -93.035 8.045 -92.865 ;
      RECT 7.955 -91.848 8.045 -90.84 ;
      RECT 7.905 -91.245 8.045 -91.075 ;
      RECT 7.955 -90.04 8.045 -89.032 ;
      RECT 7.905 -89.805 8.045 -89.635 ;
      RECT 7.955 -88.618 8.045 -87.61 ;
      RECT 7.905 -88.015 8.045 -87.845 ;
      RECT 7.955 -86.81 8.045 -85.802 ;
      RECT 7.905 -86.575 8.045 -86.405 ;
      RECT 7.955 -85.388 8.045 -84.38 ;
      RECT 7.905 -84.785 8.045 -84.615 ;
      RECT 7.955 -83.58 8.045 -82.572 ;
      RECT 7.905 -83.345 8.045 -83.175 ;
      RECT 7.955 -82.158 8.045 -81.15 ;
      RECT 7.905 -81.555 8.045 -81.385 ;
      RECT 7.955 -80.35 8.045 -79.342 ;
      RECT 7.905 -80.115 8.045 -79.945 ;
      RECT 7.955 -78.928 8.045 -77.92 ;
      RECT 7.905 -78.325 8.045 -78.155 ;
      RECT 7.955 -77.12 8.045 -76.112 ;
      RECT 7.905 -76.885 8.045 -76.715 ;
      RECT 7.955 -75.698 8.045 -74.69 ;
      RECT 7.905 -75.095 8.045 -74.925 ;
      RECT 7.955 -73.89 8.045 -72.882 ;
      RECT 7.905 -73.655 8.045 -73.485 ;
      RECT 7.955 -72.468 8.045 -71.46 ;
      RECT 7.905 -71.865 8.045 -71.695 ;
      RECT 7.955 -70.66 8.045 -69.652 ;
      RECT 7.905 -70.425 8.045 -70.255 ;
      RECT 7.955 -69.238 8.045 -68.23 ;
      RECT 7.905 -68.635 8.045 -68.465 ;
      RECT 7.955 -67.43 8.045 -66.422 ;
      RECT 7.905 -67.195 8.045 -67.025 ;
      RECT 7.955 -66.008 8.045 -65 ;
      RECT 7.905 -65.405 8.045 -65.235 ;
      RECT 7.955 -64.2 8.045 -63.192 ;
      RECT 7.905 -63.965 8.045 -63.795 ;
      RECT 7.955 -62.778 8.045 -61.77 ;
      RECT 7.905 -62.175 8.045 -62.005 ;
      RECT 7.955 -60.97 8.045 -59.962 ;
      RECT 7.905 -60.735 8.045 -60.565 ;
      RECT 7.955 -59.548 8.045 -58.54 ;
      RECT 7.905 -58.945 8.045 -58.775 ;
      RECT 7.955 -57.74 8.045 -56.732 ;
      RECT 7.905 -57.505 8.045 -57.335 ;
      RECT 7.955 -56.318 8.045 -55.31 ;
      RECT 7.905 -55.715 8.045 -55.545 ;
      RECT 7.955 -54.51 8.045 -53.502 ;
      RECT 7.905 -54.275 8.045 -54.105 ;
      RECT 7.955 -53.088 8.045 -52.08 ;
      RECT 7.905 -52.485 8.045 -52.315 ;
      RECT 7.955 -51.28 8.045 -50.272 ;
      RECT 7.905 -51.045 8.045 -50.875 ;
      RECT 7.955 -49.858 8.045 -48.85 ;
      RECT 7.905 -49.255 8.045 -49.085 ;
      RECT 7.955 -48.05 8.045 -47.042 ;
      RECT 7.905 -47.815 8.045 -47.645 ;
      RECT 7.955 -46.628 8.045 -45.62 ;
      RECT 7.905 -46.025 8.045 -45.855 ;
      RECT 7.955 -44.82 8.045 -43.812 ;
      RECT 7.905 -44.585 8.045 -44.415 ;
      RECT 7.955 -43.398 8.045 -42.39 ;
      RECT 7.905 -42.795 8.045 -42.625 ;
      RECT 7.955 -41.59 8.045 -40.582 ;
      RECT 7.905 -41.355 8.045 -41.185 ;
      RECT 7.955 -40.168 8.045 -39.16 ;
      RECT 7.905 -39.565 8.045 -39.395 ;
      RECT 7.955 -38.36 8.045 -37.352 ;
      RECT 7.905 -38.125 8.045 -37.955 ;
      RECT 7.955 -36.938 8.045 -35.93 ;
      RECT 7.905 -36.335 8.045 -36.165 ;
      RECT 7.955 -35.13 8.045 -34.122 ;
      RECT 7.905 -34.895 8.045 -34.725 ;
      RECT 7.955 -33.708 8.045 -32.7 ;
      RECT 7.905 -33.105 8.045 -32.935 ;
      RECT 7.955 -31.9 8.045 -30.892 ;
      RECT 7.905 -31.665 8.045 -31.495 ;
      RECT 7.955 -30.478 8.045 -29.47 ;
      RECT 7.905 -29.875 8.045 -29.705 ;
      RECT 7.955 -28.67 8.045 -27.662 ;
      RECT 7.905 -28.435 8.045 -28.265 ;
      RECT 7.955 -27.248 8.045 -26.24 ;
      RECT 7.905 -26.645 8.045 -26.475 ;
      RECT 7.955 -25.44 8.045 -24.432 ;
      RECT 7.905 -25.205 8.045 -25.035 ;
      RECT 7.955 -24.018 8.045 -23.01 ;
      RECT 7.905 -23.415 8.045 -23.245 ;
      RECT 7.955 -22.21 8.045 -21.202 ;
      RECT 7.905 -21.975 8.045 -21.805 ;
      RECT 7.955 -20.788 8.045 -19.78 ;
      RECT 7.905 -20.185 8.045 -20.015 ;
      RECT 7.955 -18.98 8.045 -17.972 ;
      RECT 7.905 -18.745 8.045 -18.575 ;
      RECT 7.955 -17.558 8.045 -16.55 ;
      RECT 7.905 -16.955 8.045 -16.785 ;
      RECT 7.955 -15.75 8.045 -14.742 ;
      RECT 7.905 -15.515 8.045 -15.345 ;
      RECT 7.955 -14.328 8.045 -13.32 ;
      RECT 7.905 -13.725 8.045 -13.555 ;
      RECT 7.955 -12.52 8.045 -11.512 ;
      RECT 7.905 -12.285 8.045 -12.115 ;
      RECT 7.955 -11.098 8.045 -10.09 ;
      RECT 7.905 -10.495 8.045 -10.325 ;
      RECT 7.955 -9.29 8.045 -8.282 ;
      RECT 7.905 -9.055 8.045 -8.885 ;
      RECT 7.955 -7.868 8.045 -6.86 ;
      RECT 7.905 -7.265 8.045 -7.095 ;
      RECT 7.955 -6.06 8.045 -5.052 ;
      RECT 7.905 -5.825 8.045 -5.655 ;
      RECT 7.955 -4.638 8.045 -3.63 ;
      RECT 7.905 -4.035 8.045 -3.865 ;
      RECT 7.955 -2.83 8.045 -1.822 ;
      RECT 7.905 -2.595 8.045 -2.425 ;
      RECT 7.955 -1.408 8.045 -0.4 ;
      RECT 7.905 -0.805 8.045 -0.635 ;
      RECT 7.955 0.4 8.045 1.408 ;
      RECT 7.905 0.635 8.045 0.805 ;
      RECT 7.555 -101.538 7.645 -100.531 ;
      RECT 7.555 -101.225 7.695 -101.055 ;
      RECT 7.555 -99.729 7.645 -98.722 ;
      RECT 7.555 -99.205 7.695 -99.035 ;
      RECT 7.555 -98.308 7.645 -97.301 ;
      RECT 7.555 -97.995 7.695 -97.825 ;
      RECT 7.555 -96.499 7.645 -95.492 ;
      RECT 7.555 -95.975 7.695 -95.805 ;
      RECT 7.555 -95.078 7.645 -94.071 ;
      RECT 7.555 -94.765 7.695 -94.595 ;
      RECT 7.555 -93.269 7.645 -92.262 ;
      RECT 7.555 -92.745 7.695 -92.575 ;
      RECT 7.555 -91.848 7.645 -90.841 ;
      RECT 7.555 -91.535 7.695 -91.365 ;
      RECT 7.555 -90.039 7.645 -89.032 ;
      RECT 7.555 -89.515 7.695 -89.345 ;
      RECT 7.555 -88.618 7.645 -87.611 ;
      RECT 7.555 -88.305 7.695 -88.135 ;
      RECT 7.555 -86.809 7.645 -85.802 ;
      RECT 7.555 -86.285 7.695 -86.115 ;
      RECT 7.555 -85.388 7.645 -84.381 ;
      RECT 7.555 -85.075 7.695 -84.905 ;
      RECT 7.555 -83.579 7.645 -82.572 ;
      RECT 7.555 -83.055 7.695 -82.885 ;
      RECT 7.555 -82.158 7.645 -81.151 ;
      RECT 7.555 -81.845 7.695 -81.675 ;
      RECT 7.555 -80.349 7.645 -79.342 ;
      RECT 7.555 -79.825 7.695 -79.655 ;
      RECT 7.555 -78.928 7.645 -77.921 ;
      RECT 7.555 -78.615 7.695 -78.445 ;
      RECT 7.555 -77.119 7.645 -76.112 ;
      RECT 7.555 -76.595 7.695 -76.425 ;
      RECT 7.555 -75.698 7.645 -74.691 ;
      RECT 7.555 -75.385 7.695 -75.215 ;
      RECT 7.555 -73.889 7.645 -72.882 ;
      RECT 7.555 -73.365 7.695 -73.195 ;
      RECT 7.555 -72.468 7.645 -71.461 ;
      RECT 7.555 -72.155 7.695 -71.985 ;
      RECT 7.555 -70.659 7.645 -69.652 ;
      RECT 7.555 -70.135 7.695 -69.965 ;
      RECT 7.555 -69.238 7.645 -68.231 ;
      RECT 7.555 -68.925 7.695 -68.755 ;
      RECT 7.555 -67.429 7.645 -66.422 ;
      RECT 7.555 -66.905 7.695 -66.735 ;
      RECT 7.555 -66.008 7.645 -65.001 ;
      RECT 7.555 -65.695 7.695 -65.525 ;
      RECT 7.555 -64.199 7.645 -63.192 ;
      RECT 7.555 -63.675 7.695 -63.505 ;
      RECT 7.555 -62.778 7.645 -61.771 ;
      RECT 7.555 -62.465 7.695 -62.295 ;
      RECT 7.555 -60.969 7.645 -59.962 ;
      RECT 7.555 -60.445 7.695 -60.275 ;
      RECT 7.555 -59.548 7.645 -58.541 ;
      RECT 7.555 -59.235 7.695 -59.065 ;
      RECT 7.555 -57.739 7.645 -56.732 ;
      RECT 7.555 -57.215 7.695 -57.045 ;
      RECT 7.555 -56.318 7.645 -55.311 ;
      RECT 7.555 -56.005 7.695 -55.835 ;
      RECT 7.555 -54.509 7.645 -53.502 ;
      RECT 7.555 -53.985 7.695 -53.815 ;
      RECT 7.555 -53.088 7.645 -52.081 ;
      RECT 7.555 -52.775 7.695 -52.605 ;
      RECT 7.555 -51.279 7.645 -50.272 ;
      RECT 7.555 -50.755 7.695 -50.585 ;
      RECT 7.555 -49.858 7.645 -48.851 ;
      RECT 7.555 -49.545 7.695 -49.375 ;
      RECT 7.555 -48.049 7.645 -47.042 ;
      RECT 7.555 -47.525 7.695 -47.355 ;
      RECT 7.555 -46.628 7.645 -45.621 ;
      RECT 7.555 -46.315 7.695 -46.145 ;
      RECT 7.555 -44.819 7.645 -43.812 ;
      RECT 7.555 -44.295 7.695 -44.125 ;
      RECT 7.555 -43.398 7.645 -42.391 ;
      RECT 7.555 -43.085 7.695 -42.915 ;
      RECT 7.555 -41.589 7.645 -40.582 ;
      RECT 7.555 -41.065 7.695 -40.895 ;
      RECT 7.555 -40.168 7.645 -39.161 ;
      RECT 7.555 -39.855 7.695 -39.685 ;
      RECT 7.555 -38.359 7.645 -37.352 ;
      RECT 7.555 -37.835 7.695 -37.665 ;
      RECT 7.555 -36.938 7.645 -35.931 ;
      RECT 7.555 -36.625 7.695 -36.455 ;
      RECT 7.555 -35.129 7.645 -34.122 ;
      RECT 7.555 -34.605 7.695 -34.435 ;
      RECT 7.555 -33.708 7.645 -32.701 ;
      RECT 7.555 -33.395 7.695 -33.225 ;
      RECT 7.555 -31.899 7.645 -30.892 ;
      RECT 7.555 -31.375 7.695 -31.205 ;
      RECT 7.555 -30.478 7.645 -29.471 ;
      RECT 7.555 -30.165 7.695 -29.995 ;
      RECT 7.555 -28.669 7.645 -27.662 ;
      RECT 7.555 -28.145 7.695 -27.975 ;
      RECT 7.555 -27.248 7.645 -26.241 ;
      RECT 7.555 -26.935 7.695 -26.765 ;
      RECT 7.555 -25.439 7.645 -24.432 ;
      RECT 7.555 -24.915 7.695 -24.745 ;
      RECT 7.555 -24.018 7.645 -23.011 ;
      RECT 7.555 -23.705 7.695 -23.535 ;
      RECT 7.555 -22.209 7.645 -21.202 ;
      RECT 7.555 -21.685 7.695 -21.515 ;
      RECT 7.555 -20.788 7.645 -19.781 ;
      RECT 7.555 -20.475 7.695 -20.305 ;
      RECT 7.555 -18.979 7.645 -17.972 ;
      RECT 7.555 -18.455 7.695 -18.285 ;
      RECT 7.555 -17.558 7.645 -16.551 ;
      RECT 7.555 -17.245 7.695 -17.075 ;
      RECT 7.555 -15.749 7.645 -14.742 ;
      RECT 7.555 -15.225 7.695 -15.055 ;
      RECT 7.555 -14.328 7.645 -13.321 ;
      RECT 7.555 -14.015 7.695 -13.845 ;
      RECT 7.555 -12.519 7.645 -11.512 ;
      RECT 7.555 -11.995 7.695 -11.825 ;
      RECT 7.555 -11.098 7.645 -10.091 ;
      RECT 7.555 -10.785 7.695 -10.615 ;
      RECT 7.555 -9.289 7.645 -8.282 ;
      RECT 7.555 -8.765 7.695 -8.595 ;
      RECT 7.555 -7.868 7.645 -6.861 ;
      RECT 7.555 -7.555 7.695 -7.385 ;
      RECT 7.555 -6.059 7.645 -5.052 ;
      RECT 7.555 -5.535 7.695 -5.365 ;
      RECT 7.555 -4.638 7.645 -3.631 ;
      RECT 7.555 -4.325 7.695 -4.155 ;
      RECT 7.555 -2.829 7.645 -1.822 ;
      RECT 7.555 -2.305 7.695 -2.135 ;
      RECT 7.555 -1.408 7.645 -0.401 ;
      RECT 7.555 -1.095 7.695 -0.925 ;
      RECT 7.555 0.401 7.645 1.408 ;
      RECT 7.555 0.925 7.695 1.095 ;
      RECT 5.705 -111.685 7.185 -111.585 ;
      RECT 5.705 -112.055 5.805 -111.585 ;
      RECT 5.51 -114.395 7.085 -114.275 ;
      RECT 6.985 -114.895 7.085 -114.275 ;
      RECT 6.39 -114.895 6.49 -114.275 ;
      RECT 5.51 -114.85 5.61 -114.275 ;
      RECT 6.755 -101.538 6.845 -100.53 ;
      RECT 6.705 -100.935 6.845 -100.765 ;
      RECT 6.755 -99.73 6.845 -98.722 ;
      RECT 6.705 -99.495 6.845 -99.325 ;
      RECT 6.755 -98.308 6.845 -97.3 ;
      RECT 6.705 -97.705 6.845 -97.535 ;
      RECT 6.755 -96.5 6.845 -95.492 ;
      RECT 6.705 -96.265 6.845 -96.095 ;
      RECT 6.755 -95.078 6.845 -94.07 ;
      RECT 6.705 -94.475 6.845 -94.305 ;
      RECT 6.755 -93.27 6.845 -92.262 ;
      RECT 6.705 -93.035 6.845 -92.865 ;
      RECT 6.755 -91.848 6.845 -90.84 ;
      RECT 6.705 -91.245 6.845 -91.075 ;
      RECT 6.755 -90.04 6.845 -89.032 ;
      RECT 6.705 -89.805 6.845 -89.635 ;
      RECT 6.755 -88.618 6.845 -87.61 ;
      RECT 6.705 -88.015 6.845 -87.845 ;
      RECT 6.755 -86.81 6.845 -85.802 ;
      RECT 6.705 -86.575 6.845 -86.405 ;
      RECT 6.755 -85.388 6.845 -84.38 ;
      RECT 6.705 -84.785 6.845 -84.615 ;
      RECT 6.755 -83.58 6.845 -82.572 ;
      RECT 6.705 -83.345 6.845 -83.175 ;
      RECT 6.755 -82.158 6.845 -81.15 ;
      RECT 6.705 -81.555 6.845 -81.385 ;
      RECT 6.755 -80.35 6.845 -79.342 ;
      RECT 6.705 -80.115 6.845 -79.945 ;
      RECT 6.755 -78.928 6.845 -77.92 ;
      RECT 6.705 -78.325 6.845 -78.155 ;
      RECT 6.755 -77.12 6.845 -76.112 ;
      RECT 6.705 -76.885 6.845 -76.715 ;
      RECT 6.755 -75.698 6.845 -74.69 ;
      RECT 6.705 -75.095 6.845 -74.925 ;
      RECT 6.755 -73.89 6.845 -72.882 ;
      RECT 6.705 -73.655 6.845 -73.485 ;
      RECT 6.755 -72.468 6.845 -71.46 ;
      RECT 6.705 -71.865 6.845 -71.695 ;
      RECT 6.755 -70.66 6.845 -69.652 ;
      RECT 6.705 -70.425 6.845 -70.255 ;
      RECT 6.755 -69.238 6.845 -68.23 ;
      RECT 6.705 -68.635 6.845 -68.465 ;
      RECT 6.755 -67.43 6.845 -66.422 ;
      RECT 6.705 -67.195 6.845 -67.025 ;
      RECT 6.755 -66.008 6.845 -65 ;
      RECT 6.705 -65.405 6.845 -65.235 ;
      RECT 6.755 -64.2 6.845 -63.192 ;
      RECT 6.705 -63.965 6.845 -63.795 ;
      RECT 6.755 -62.778 6.845 -61.77 ;
      RECT 6.705 -62.175 6.845 -62.005 ;
      RECT 6.755 -60.97 6.845 -59.962 ;
      RECT 6.705 -60.735 6.845 -60.565 ;
      RECT 6.755 -59.548 6.845 -58.54 ;
      RECT 6.705 -58.945 6.845 -58.775 ;
      RECT 6.755 -57.74 6.845 -56.732 ;
      RECT 6.705 -57.505 6.845 -57.335 ;
      RECT 6.755 -56.318 6.845 -55.31 ;
      RECT 6.705 -55.715 6.845 -55.545 ;
      RECT 6.755 -54.51 6.845 -53.502 ;
      RECT 6.705 -54.275 6.845 -54.105 ;
      RECT 6.755 -53.088 6.845 -52.08 ;
      RECT 6.705 -52.485 6.845 -52.315 ;
      RECT 6.755 -51.28 6.845 -50.272 ;
      RECT 6.705 -51.045 6.845 -50.875 ;
      RECT 6.755 -49.858 6.845 -48.85 ;
      RECT 6.705 -49.255 6.845 -49.085 ;
      RECT 6.755 -48.05 6.845 -47.042 ;
      RECT 6.705 -47.815 6.845 -47.645 ;
      RECT 6.755 -46.628 6.845 -45.62 ;
      RECT 6.705 -46.025 6.845 -45.855 ;
      RECT 6.755 -44.82 6.845 -43.812 ;
      RECT 6.705 -44.585 6.845 -44.415 ;
      RECT 6.755 -43.398 6.845 -42.39 ;
      RECT 6.705 -42.795 6.845 -42.625 ;
      RECT 6.755 -41.59 6.845 -40.582 ;
      RECT 6.705 -41.355 6.845 -41.185 ;
      RECT 6.755 -40.168 6.845 -39.16 ;
      RECT 6.705 -39.565 6.845 -39.395 ;
      RECT 6.755 -38.36 6.845 -37.352 ;
      RECT 6.705 -38.125 6.845 -37.955 ;
      RECT 6.755 -36.938 6.845 -35.93 ;
      RECT 6.705 -36.335 6.845 -36.165 ;
      RECT 6.755 -35.13 6.845 -34.122 ;
      RECT 6.705 -34.895 6.845 -34.725 ;
      RECT 6.755 -33.708 6.845 -32.7 ;
      RECT 6.705 -33.105 6.845 -32.935 ;
      RECT 6.755 -31.9 6.845 -30.892 ;
      RECT 6.705 -31.665 6.845 -31.495 ;
      RECT 6.755 -30.478 6.845 -29.47 ;
      RECT 6.705 -29.875 6.845 -29.705 ;
      RECT 6.755 -28.67 6.845 -27.662 ;
      RECT 6.705 -28.435 6.845 -28.265 ;
      RECT 6.755 -27.248 6.845 -26.24 ;
      RECT 6.705 -26.645 6.845 -26.475 ;
      RECT 6.755 -25.44 6.845 -24.432 ;
      RECT 6.705 -25.205 6.845 -25.035 ;
      RECT 6.755 -24.018 6.845 -23.01 ;
      RECT 6.705 -23.415 6.845 -23.245 ;
      RECT 6.755 -22.21 6.845 -21.202 ;
      RECT 6.705 -21.975 6.845 -21.805 ;
      RECT 6.755 -20.788 6.845 -19.78 ;
      RECT 6.705 -20.185 6.845 -20.015 ;
      RECT 6.755 -18.98 6.845 -17.972 ;
      RECT 6.705 -18.745 6.845 -18.575 ;
      RECT 6.755 -17.558 6.845 -16.55 ;
      RECT 6.705 -16.955 6.845 -16.785 ;
      RECT 6.755 -15.75 6.845 -14.742 ;
      RECT 6.705 -15.515 6.845 -15.345 ;
      RECT 6.755 -14.328 6.845 -13.32 ;
      RECT 6.705 -13.725 6.845 -13.555 ;
      RECT 6.755 -12.52 6.845 -11.512 ;
      RECT 6.705 -12.285 6.845 -12.115 ;
      RECT 6.755 -11.098 6.845 -10.09 ;
      RECT 6.705 -10.495 6.845 -10.325 ;
      RECT 6.755 -9.29 6.845 -8.282 ;
      RECT 6.705 -9.055 6.845 -8.885 ;
      RECT 6.755 -7.868 6.845 -6.86 ;
      RECT 6.705 -7.265 6.845 -7.095 ;
      RECT 6.755 -6.06 6.845 -5.052 ;
      RECT 6.705 -5.825 6.845 -5.655 ;
      RECT 6.755 -4.638 6.845 -3.63 ;
      RECT 6.705 -4.035 6.845 -3.865 ;
      RECT 6.755 -2.83 6.845 -1.822 ;
      RECT 6.705 -2.595 6.845 -2.425 ;
      RECT 6.755 -1.408 6.845 -0.4 ;
      RECT 6.705 -0.805 6.845 -0.635 ;
      RECT 6.755 0.4 6.845 1.408 ;
      RECT 6.705 0.635 6.845 0.805 ;
      RECT 6.63 -114.685 6.805 -114.515 ;
      RECT 6.705 -114.895 6.805 -114.515 ;
      RECT 5.745 -113.555 5.845 -113.09 ;
      RECT 6.11 -113.555 6.21 -113.1 ;
      RECT 5.745 -113.555 6.59 -113.385 ;
      RECT 6.355 -101.538 6.445 -100.531 ;
      RECT 6.355 -101.225 6.495 -101.055 ;
      RECT 6.355 -99.729 6.445 -98.722 ;
      RECT 6.355 -99.205 6.495 -99.035 ;
      RECT 6.355 -98.308 6.445 -97.301 ;
      RECT 6.355 -97.995 6.495 -97.825 ;
      RECT 6.355 -96.499 6.445 -95.492 ;
      RECT 6.355 -95.975 6.495 -95.805 ;
      RECT 6.355 -95.078 6.445 -94.071 ;
      RECT 6.355 -94.765 6.495 -94.595 ;
      RECT 6.355 -93.269 6.445 -92.262 ;
      RECT 6.355 -92.745 6.495 -92.575 ;
      RECT 6.355 -91.848 6.445 -90.841 ;
      RECT 6.355 -91.535 6.495 -91.365 ;
      RECT 6.355 -90.039 6.445 -89.032 ;
      RECT 6.355 -89.515 6.495 -89.345 ;
      RECT 6.355 -88.618 6.445 -87.611 ;
      RECT 6.355 -88.305 6.495 -88.135 ;
      RECT 6.355 -86.809 6.445 -85.802 ;
      RECT 6.355 -86.285 6.495 -86.115 ;
      RECT 6.355 -85.388 6.445 -84.381 ;
      RECT 6.355 -85.075 6.495 -84.905 ;
      RECT 6.355 -83.579 6.445 -82.572 ;
      RECT 6.355 -83.055 6.495 -82.885 ;
      RECT 6.355 -82.158 6.445 -81.151 ;
      RECT 6.355 -81.845 6.495 -81.675 ;
      RECT 6.355 -80.349 6.445 -79.342 ;
      RECT 6.355 -79.825 6.495 -79.655 ;
      RECT 6.355 -78.928 6.445 -77.921 ;
      RECT 6.355 -78.615 6.495 -78.445 ;
      RECT 6.355 -77.119 6.445 -76.112 ;
      RECT 6.355 -76.595 6.495 -76.425 ;
      RECT 6.355 -75.698 6.445 -74.691 ;
      RECT 6.355 -75.385 6.495 -75.215 ;
      RECT 6.355 -73.889 6.445 -72.882 ;
      RECT 6.355 -73.365 6.495 -73.195 ;
      RECT 6.355 -72.468 6.445 -71.461 ;
      RECT 6.355 -72.155 6.495 -71.985 ;
      RECT 6.355 -70.659 6.445 -69.652 ;
      RECT 6.355 -70.135 6.495 -69.965 ;
      RECT 6.355 -69.238 6.445 -68.231 ;
      RECT 6.355 -68.925 6.495 -68.755 ;
      RECT 6.355 -67.429 6.445 -66.422 ;
      RECT 6.355 -66.905 6.495 -66.735 ;
      RECT 6.355 -66.008 6.445 -65.001 ;
      RECT 6.355 -65.695 6.495 -65.525 ;
      RECT 6.355 -64.199 6.445 -63.192 ;
      RECT 6.355 -63.675 6.495 -63.505 ;
      RECT 6.355 -62.778 6.445 -61.771 ;
      RECT 6.355 -62.465 6.495 -62.295 ;
      RECT 6.355 -60.969 6.445 -59.962 ;
      RECT 6.355 -60.445 6.495 -60.275 ;
      RECT 6.355 -59.548 6.445 -58.541 ;
      RECT 6.355 -59.235 6.495 -59.065 ;
      RECT 6.355 -57.739 6.445 -56.732 ;
      RECT 6.355 -57.215 6.495 -57.045 ;
      RECT 6.355 -56.318 6.445 -55.311 ;
      RECT 6.355 -56.005 6.495 -55.835 ;
      RECT 6.355 -54.509 6.445 -53.502 ;
      RECT 6.355 -53.985 6.495 -53.815 ;
      RECT 6.355 -53.088 6.445 -52.081 ;
      RECT 6.355 -52.775 6.495 -52.605 ;
      RECT 6.355 -51.279 6.445 -50.272 ;
      RECT 6.355 -50.755 6.495 -50.585 ;
      RECT 6.355 -49.858 6.445 -48.851 ;
      RECT 6.355 -49.545 6.495 -49.375 ;
      RECT 6.355 -48.049 6.445 -47.042 ;
      RECT 6.355 -47.525 6.495 -47.355 ;
      RECT 6.355 -46.628 6.445 -45.621 ;
      RECT 6.355 -46.315 6.495 -46.145 ;
      RECT 6.355 -44.819 6.445 -43.812 ;
      RECT 6.355 -44.295 6.495 -44.125 ;
      RECT 6.355 -43.398 6.445 -42.391 ;
      RECT 6.355 -43.085 6.495 -42.915 ;
      RECT 6.355 -41.589 6.445 -40.582 ;
      RECT 6.355 -41.065 6.495 -40.895 ;
      RECT 6.355 -40.168 6.445 -39.161 ;
      RECT 6.355 -39.855 6.495 -39.685 ;
      RECT 6.355 -38.359 6.445 -37.352 ;
      RECT 6.355 -37.835 6.495 -37.665 ;
      RECT 6.355 -36.938 6.445 -35.931 ;
      RECT 6.355 -36.625 6.495 -36.455 ;
      RECT 6.355 -35.129 6.445 -34.122 ;
      RECT 6.355 -34.605 6.495 -34.435 ;
      RECT 6.355 -33.708 6.445 -32.701 ;
      RECT 6.355 -33.395 6.495 -33.225 ;
      RECT 6.355 -31.899 6.445 -30.892 ;
      RECT 6.355 -31.375 6.495 -31.205 ;
      RECT 6.355 -30.478 6.445 -29.471 ;
      RECT 6.355 -30.165 6.495 -29.995 ;
      RECT 6.355 -28.669 6.445 -27.662 ;
      RECT 6.355 -28.145 6.495 -27.975 ;
      RECT 6.355 -27.248 6.445 -26.241 ;
      RECT 6.355 -26.935 6.495 -26.765 ;
      RECT 6.355 -25.439 6.445 -24.432 ;
      RECT 6.355 -24.915 6.495 -24.745 ;
      RECT 6.355 -24.018 6.445 -23.011 ;
      RECT 6.355 -23.705 6.495 -23.535 ;
      RECT 6.355 -22.209 6.445 -21.202 ;
      RECT 6.355 -21.685 6.495 -21.515 ;
      RECT 6.355 -20.788 6.445 -19.781 ;
      RECT 6.355 -20.475 6.495 -20.305 ;
      RECT 6.355 -18.979 6.445 -17.972 ;
      RECT 6.355 -18.455 6.495 -18.285 ;
      RECT 6.355 -17.558 6.445 -16.551 ;
      RECT 6.355 -17.245 6.495 -17.075 ;
      RECT 6.355 -15.749 6.445 -14.742 ;
      RECT 6.355 -15.225 6.495 -15.055 ;
      RECT 6.355 -14.328 6.445 -13.321 ;
      RECT 6.355 -14.015 6.495 -13.845 ;
      RECT 6.355 -12.519 6.445 -11.512 ;
      RECT 6.355 -11.995 6.495 -11.825 ;
      RECT 6.355 -11.098 6.445 -10.091 ;
      RECT 6.355 -10.785 6.495 -10.615 ;
      RECT 6.355 -9.289 6.445 -8.282 ;
      RECT 6.355 -8.765 6.495 -8.595 ;
      RECT 6.355 -7.868 6.445 -6.861 ;
      RECT 6.355 -7.555 6.495 -7.385 ;
      RECT 6.355 -6.059 6.445 -5.052 ;
      RECT 6.355 -5.535 6.495 -5.365 ;
      RECT 6.355 -4.638 6.445 -3.631 ;
      RECT 6.355 -4.325 6.495 -4.155 ;
      RECT 6.355 -2.829 6.445 -1.822 ;
      RECT 6.355 -2.305 6.495 -2.135 ;
      RECT 6.355 -1.408 6.445 -0.401 ;
      RECT 6.355 -1.095 6.495 -0.925 ;
      RECT 6.355 0.401 6.445 1.408 ;
      RECT 6.355 0.925 6.495 1.095 ;
      RECT 6.04 -114.685 6.21 -114.515 ;
      RECT 6.11 -114.895 6.21 -114.515 ;
      RECT 5.555 -101.538 5.645 -100.53 ;
      RECT 5.505 -100.935 5.645 -100.765 ;
      RECT 5.555 -99.73 5.645 -98.722 ;
      RECT 5.505 -99.495 5.645 -99.325 ;
      RECT 5.555 -98.308 5.645 -97.3 ;
      RECT 5.505 -97.705 5.645 -97.535 ;
      RECT 5.555 -96.5 5.645 -95.492 ;
      RECT 5.505 -96.265 5.645 -96.095 ;
      RECT 5.555 -95.078 5.645 -94.07 ;
      RECT 5.505 -94.475 5.645 -94.305 ;
      RECT 5.555 -93.27 5.645 -92.262 ;
      RECT 5.505 -93.035 5.645 -92.865 ;
      RECT 5.555 -91.848 5.645 -90.84 ;
      RECT 5.505 -91.245 5.645 -91.075 ;
      RECT 5.555 -90.04 5.645 -89.032 ;
      RECT 5.505 -89.805 5.645 -89.635 ;
      RECT 5.555 -88.618 5.645 -87.61 ;
      RECT 5.505 -88.015 5.645 -87.845 ;
      RECT 5.555 -86.81 5.645 -85.802 ;
      RECT 5.505 -86.575 5.645 -86.405 ;
      RECT 5.555 -85.388 5.645 -84.38 ;
      RECT 5.505 -84.785 5.645 -84.615 ;
      RECT 5.555 -83.58 5.645 -82.572 ;
      RECT 5.505 -83.345 5.645 -83.175 ;
      RECT 5.555 -82.158 5.645 -81.15 ;
      RECT 5.505 -81.555 5.645 -81.385 ;
      RECT 5.555 -80.35 5.645 -79.342 ;
      RECT 5.505 -80.115 5.645 -79.945 ;
      RECT 5.555 -78.928 5.645 -77.92 ;
      RECT 5.505 -78.325 5.645 -78.155 ;
      RECT 5.555 -77.12 5.645 -76.112 ;
      RECT 5.505 -76.885 5.645 -76.715 ;
      RECT 5.555 -75.698 5.645 -74.69 ;
      RECT 5.505 -75.095 5.645 -74.925 ;
      RECT 5.555 -73.89 5.645 -72.882 ;
      RECT 5.505 -73.655 5.645 -73.485 ;
      RECT 5.555 -72.468 5.645 -71.46 ;
      RECT 5.505 -71.865 5.645 -71.695 ;
      RECT 5.555 -70.66 5.645 -69.652 ;
      RECT 5.505 -70.425 5.645 -70.255 ;
      RECT 5.555 -69.238 5.645 -68.23 ;
      RECT 5.505 -68.635 5.645 -68.465 ;
      RECT 5.555 -67.43 5.645 -66.422 ;
      RECT 5.505 -67.195 5.645 -67.025 ;
      RECT 5.555 -66.008 5.645 -65 ;
      RECT 5.505 -65.405 5.645 -65.235 ;
      RECT 5.555 -64.2 5.645 -63.192 ;
      RECT 5.505 -63.965 5.645 -63.795 ;
      RECT 5.555 -62.778 5.645 -61.77 ;
      RECT 5.505 -62.175 5.645 -62.005 ;
      RECT 5.555 -60.97 5.645 -59.962 ;
      RECT 5.505 -60.735 5.645 -60.565 ;
      RECT 5.555 -59.548 5.645 -58.54 ;
      RECT 5.505 -58.945 5.645 -58.775 ;
      RECT 5.555 -57.74 5.645 -56.732 ;
      RECT 5.505 -57.505 5.645 -57.335 ;
      RECT 5.555 -56.318 5.645 -55.31 ;
      RECT 5.505 -55.715 5.645 -55.545 ;
      RECT 5.555 -54.51 5.645 -53.502 ;
      RECT 5.505 -54.275 5.645 -54.105 ;
      RECT 5.555 -53.088 5.645 -52.08 ;
      RECT 5.505 -52.485 5.645 -52.315 ;
      RECT 5.555 -51.28 5.645 -50.272 ;
      RECT 5.505 -51.045 5.645 -50.875 ;
      RECT 5.555 -49.858 5.645 -48.85 ;
      RECT 5.505 -49.255 5.645 -49.085 ;
      RECT 5.555 -48.05 5.645 -47.042 ;
      RECT 5.505 -47.815 5.645 -47.645 ;
      RECT 5.555 -46.628 5.645 -45.62 ;
      RECT 5.505 -46.025 5.645 -45.855 ;
      RECT 5.555 -44.82 5.645 -43.812 ;
      RECT 5.505 -44.585 5.645 -44.415 ;
      RECT 5.555 -43.398 5.645 -42.39 ;
      RECT 5.505 -42.795 5.645 -42.625 ;
      RECT 5.555 -41.59 5.645 -40.582 ;
      RECT 5.505 -41.355 5.645 -41.185 ;
      RECT 5.555 -40.168 5.645 -39.16 ;
      RECT 5.505 -39.565 5.645 -39.395 ;
      RECT 5.555 -38.36 5.645 -37.352 ;
      RECT 5.505 -38.125 5.645 -37.955 ;
      RECT 5.555 -36.938 5.645 -35.93 ;
      RECT 5.505 -36.335 5.645 -36.165 ;
      RECT 5.555 -35.13 5.645 -34.122 ;
      RECT 5.505 -34.895 5.645 -34.725 ;
      RECT 5.555 -33.708 5.645 -32.7 ;
      RECT 5.505 -33.105 5.645 -32.935 ;
      RECT 5.555 -31.9 5.645 -30.892 ;
      RECT 5.505 -31.665 5.645 -31.495 ;
      RECT 5.555 -30.478 5.645 -29.47 ;
      RECT 5.505 -29.875 5.645 -29.705 ;
      RECT 5.555 -28.67 5.645 -27.662 ;
      RECT 5.505 -28.435 5.645 -28.265 ;
      RECT 5.555 -27.248 5.645 -26.24 ;
      RECT 5.505 -26.645 5.645 -26.475 ;
      RECT 5.555 -25.44 5.645 -24.432 ;
      RECT 5.505 -25.205 5.645 -25.035 ;
      RECT 5.555 -24.018 5.645 -23.01 ;
      RECT 5.505 -23.415 5.645 -23.245 ;
      RECT 5.555 -22.21 5.645 -21.202 ;
      RECT 5.505 -21.975 5.645 -21.805 ;
      RECT 5.555 -20.788 5.645 -19.78 ;
      RECT 5.505 -20.185 5.645 -20.015 ;
      RECT 5.555 -18.98 5.645 -17.972 ;
      RECT 5.505 -18.745 5.645 -18.575 ;
      RECT 5.555 -17.558 5.645 -16.55 ;
      RECT 5.505 -16.955 5.645 -16.785 ;
      RECT 5.555 -15.75 5.645 -14.742 ;
      RECT 5.505 -15.515 5.645 -15.345 ;
      RECT 5.555 -14.328 5.645 -13.32 ;
      RECT 5.505 -13.725 5.645 -13.555 ;
      RECT 5.555 -12.52 5.645 -11.512 ;
      RECT 5.505 -12.285 5.645 -12.115 ;
      RECT 5.555 -11.098 5.645 -10.09 ;
      RECT 5.505 -10.495 5.645 -10.325 ;
      RECT 5.555 -9.29 5.645 -8.282 ;
      RECT 5.505 -9.055 5.645 -8.885 ;
      RECT 5.555 -7.868 5.645 -6.86 ;
      RECT 5.505 -7.265 5.645 -7.095 ;
      RECT 5.555 -6.06 5.645 -5.052 ;
      RECT 5.505 -5.825 5.645 -5.655 ;
      RECT 5.555 -4.638 5.645 -3.63 ;
      RECT 5.505 -4.035 5.645 -3.865 ;
      RECT 5.555 -2.83 5.645 -1.822 ;
      RECT 5.505 -2.595 5.645 -2.425 ;
      RECT 5.555 -1.408 5.645 -0.4 ;
      RECT 5.505 -0.805 5.645 -0.635 ;
      RECT 5.555 0.4 5.645 1.408 ;
      RECT 5.505 0.635 5.645 0.805 ;
      RECT 5.155 -101.538 5.245 -100.531 ;
      RECT 5.155 -101.225 5.295 -101.055 ;
      RECT 5.155 -99.729 5.245 -98.722 ;
      RECT 5.155 -99.205 5.295 -99.035 ;
      RECT 5.155 -98.308 5.245 -97.301 ;
      RECT 5.155 -97.995 5.295 -97.825 ;
      RECT 5.155 -96.499 5.245 -95.492 ;
      RECT 5.155 -95.975 5.295 -95.805 ;
      RECT 5.155 -95.078 5.245 -94.071 ;
      RECT 5.155 -94.765 5.295 -94.595 ;
      RECT 5.155 -93.269 5.245 -92.262 ;
      RECT 5.155 -92.745 5.295 -92.575 ;
      RECT 5.155 -91.848 5.245 -90.841 ;
      RECT 5.155 -91.535 5.295 -91.365 ;
      RECT 5.155 -90.039 5.245 -89.032 ;
      RECT 5.155 -89.515 5.295 -89.345 ;
      RECT 5.155 -88.618 5.245 -87.611 ;
      RECT 5.155 -88.305 5.295 -88.135 ;
      RECT 5.155 -86.809 5.245 -85.802 ;
      RECT 5.155 -86.285 5.295 -86.115 ;
      RECT 5.155 -85.388 5.245 -84.381 ;
      RECT 5.155 -85.075 5.295 -84.905 ;
      RECT 5.155 -83.579 5.245 -82.572 ;
      RECT 5.155 -83.055 5.295 -82.885 ;
      RECT 5.155 -82.158 5.245 -81.151 ;
      RECT 5.155 -81.845 5.295 -81.675 ;
      RECT 5.155 -80.349 5.245 -79.342 ;
      RECT 5.155 -79.825 5.295 -79.655 ;
      RECT 5.155 -78.928 5.245 -77.921 ;
      RECT 5.155 -78.615 5.295 -78.445 ;
      RECT 5.155 -77.119 5.245 -76.112 ;
      RECT 5.155 -76.595 5.295 -76.425 ;
      RECT 5.155 -75.698 5.245 -74.691 ;
      RECT 5.155 -75.385 5.295 -75.215 ;
      RECT 5.155 -73.889 5.245 -72.882 ;
      RECT 5.155 -73.365 5.295 -73.195 ;
      RECT 5.155 -72.468 5.245 -71.461 ;
      RECT 5.155 -72.155 5.295 -71.985 ;
      RECT 5.155 -70.659 5.245 -69.652 ;
      RECT 5.155 -70.135 5.295 -69.965 ;
      RECT 5.155 -69.238 5.245 -68.231 ;
      RECT 5.155 -68.925 5.295 -68.755 ;
      RECT 5.155 -67.429 5.245 -66.422 ;
      RECT 5.155 -66.905 5.295 -66.735 ;
      RECT 5.155 -66.008 5.245 -65.001 ;
      RECT 5.155 -65.695 5.295 -65.525 ;
      RECT 5.155 -64.199 5.245 -63.192 ;
      RECT 5.155 -63.675 5.295 -63.505 ;
      RECT 5.155 -62.778 5.245 -61.771 ;
      RECT 5.155 -62.465 5.295 -62.295 ;
      RECT 5.155 -60.969 5.245 -59.962 ;
      RECT 5.155 -60.445 5.295 -60.275 ;
      RECT 5.155 -59.548 5.245 -58.541 ;
      RECT 5.155 -59.235 5.295 -59.065 ;
      RECT 5.155 -57.739 5.245 -56.732 ;
      RECT 5.155 -57.215 5.295 -57.045 ;
      RECT 5.155 -56.318 5.245 -55.311 ;
      RECT 5.155 -56.005 5.295 -55.835 ;
      RECT 5.155 -54.509 5.245 -53.502 ;
      RECT 5.155 -53.985 5.295 -53.815 ;
      RECT 5.155 -53.088 5.245 -52.081 ;
      RECT 5.155 -52.775 5.295 -52.605 ;
      RECT 5.155 -51.279 5.245 -50.272 ;
      RECT 5.155 -50.755 5.295 -50.585 ;
      RECT 5.155 -49.858 5.245 -48.851 ;
      RECT 5.155 -49.545 5.295 -49.375 ;
      RECT 5.155 -48.049 5.245 -47.042 ;
      RECT 5.155 -47.525 5.295 -47.355 ;
      RECT 5.155 -46.628 5.245 -45.621 ;
      RECT 5.155 -46.315 5.295 -46.145 ;
      RECT 5.155 -44.819 5.245 -43.812 ;
      RECT 5.155 -44.295 5.295 -44.125 ;
      RECT 5.155 -43.398 5.245 -42.391 ;
      RECT 5.155 -43.085 5.295 -42.915 ;
      RECT 5.155 -41.589 5.245 -40.582 ;
      RECT 5.155 -41.065 5.295 -40.895 ;
      RECT 5.155 -40.168 5.245 -39.161 ;
      RECT 5.155 -39.855 5.295 -39.685 ;
      RECT 5.155 -38.359 5.245 -37.352 ;
      RECT 5.155 -37.835 5.295 -37.665 ;
      RECT 5.155 -36.938 5.245 -35.931 ;
      RECT 5.155 -36.625 5.295 -36.455 ;
      RECT 5.155 -35.129 5.245 -34.122 ;
      RECT 5.155 -34.605 5.295 -34.435 ;
      RECT 5.155 -33.708 5.245 -32.701 ;
      RECT 5.155 -33.395 5.295 -33.225 ;
      RECT 5.155 -31.899 5.245 -30.892 ;
      RECT 5.155 -31.375 5.295 -31.205 ;
      RECT 5.155 -30.478 5.245 -29.471 ;
      RECT 5.155 -30.165 5.295 -29.995 ;
      RECT 5.155 -28.669 5.245 -27.662 ;
      RECT 5.155 -28.145 5.295 -27.975 ;
      RECT 5.155 -27.248 5.245 -26.241 ;
      RECT 5.155 -26.935 5.295 -26.765 ;
      RECT 5.155 -25.439 5.245 -24.432 ;
      RECT 5.155 -24.915 5.295 -24.745 ;
      RECT 5.155 -24.018 5.245 -23.011 ;
      RECT 5.155 -23.705 5.295 -23.535 ;
      RECT 5.155 -22.209 5.245 -21.202 ;
      RECT 5.155 -21.685 5.295 -21.515 ;
      RECT 5.155 -20.788 5.245 -19.781 ;
      RECT 5.155 -20.475 5.295 -20.305 ;
      RECT 5.155 -18.979 5.245 -17.972 ;
      RECT 5.155 -18.455 5.295 -18.285 ;
      RECT 5.155 -17.558 5.245 -16.551 ;
      RECT 5.155 -17.245 5.295 -17.075 ;
      RECT 5.155 -15.749 5.245 -14.742 ;
      RECT 5.155 -15.225 5.295 -15.055 ;
      RECT 5.155 -14.328 5.245 -13.321 ;
      RECT 5.155 -14.015 5.295 -13.845 ;
      RECT 5.155 -12.519 5.245 -11.512 ;
      RECT 5.155 -11.995 5.295 -11.825 ;
      RECT 5.155 -11.098 5.245 -10.091 ;
      RECT 5.155 -10.785 5.295 -10.615 ;
      RECT 5.155 -9.289 5.245 -8.282 ;
      RECT 5.155 -8.765 5.295 -8.595 ;
      RECT 5.155 -7.868 5.245 -6.861 ;
      RECT 5.155 -7.555 5.295 -7.385 ;
      RECT 5.155 -6.059 5.245 -5.052 ;
      RECT 5.155 -5.535 5.295 -5.365 ;
      RECT 5.155 -4.638 5.245 -3.631 ;
      RECT 5.155 -4.325 5.295 -4.155 ;
      RECT 5.155 -2.829 5.245 -1.822 ;
      RECT 5.155 -2.305 5.295 -2.135 ;
      RECT 5.155 -1.408 5.245 -0.401 ;
      RECT 5.155 -1.095 5.295 -0.925 ;
      RECT 5.155 0.401 5.245 1.408 ;
      RECT 5.155 0.925 5.295 1.095 ;
      RECT 0.985 -108.935 4.765 -108.815 ;
      RECT 2.305 -109.475 2.405 -108.815 ;
      RECT 1.745 -109.475 1.845 -108.815 ;
      RECT 1.185 -109.475 1.285 -108.815 ;
      RECT 4.355 -101.538 4.445 -100.53 ;
      RECT 4.305 -100.935 4.445 -100.765 ;
      RECT 4.355 -99.73 4.445 -98.722 ;
      RECT 4.305 -99.495 4.445 -99.325 ;
      RECT 4.355 -98.308 4.445 -97.3 ;
      RECT 4.305 -97.705 4.445 -97.535 ;
      RECT 4.355 -96.5 4.445 -95.492 ;
      RECT 4.305 -96.265 4.445 -96.095 ;
      RECT 4.355 -95.078 4.445 -94.07 ;
      RECT 4.305 -94.475 4.445 -94.305 ;
      RECT 4.355 -93.27 4.445 -92.262 ;
      RECT 4.305 -93.035 4.445 -92.865 ;
      RECT 4.355 -91.848 4.445 -90.84 ;
      RECT 4.305 -91.245 4.445 -91.075 ;
      RECT 4.355 -90.04 4.445 -89.032 ;
      RECT 4.305 -89.805 4.445 -89.635 ;
      RECT 4.355 -88.618 4.445 -87.61 ;
      RECT 4.305 -88.015 4.445 -87.845 ;
      RECT 4.355 -86.81 4.445 -85.802 ;
      RECT 4.305 -86.575 4.445 -86.405 ;
      RECT 4.355 -85.388 4.445 -84.38 ;
      RECT 4.305 -84.785 4.445 -84.615 ;
      RECT 4.355 -83.58 4.445 -82.572 ;
      RECT 4.305 -83.345 4.445 -83.175 ;
      RECT 4.355 -82.158 4.445 -81.15 ;
      RECT 4.305 -81.555 4.445 -81.385 ;
      RECT 4.355 -80.35 4.445 -79.342 ;
      RECT 4.305 -80.115 4.445 -79.945 ;
      RECT 4.355 -78.928 4.445 -77.92 ;
      RECT 4.305 -78.325 4.445 -78.155 ;
      RECT 4.355 -77.12 4.445 -76.112 ;
      RECT 4.305 -76.885 4.445 -76.715 ;
      RECT 4.355 -75.698 4.445 -74.69 ;
      RECT 4.305 -75.095 4.445 -74.925 ;
      RECT 4.355 -73.89 4.445 -72.882 ;
      RECT 4.305 -73.655 4.445 -73.485 ;
      RECT 4.355 -72.468 4.445 -71.46 ;
      RECT 4.305 -71.865 4.445 -71.695 ;
      RECT 4.355 -70.66 4.445 -69.652 ;
      RECT 4.305 -70.425 4.445 -70.255 ;
      RECT 4.355 -69.238 4.445 -68.23 ;
      RECT 4.305 -68.635 4.445 -68.465 ;
      RECT 4.355 -67.43 4.445 -66.422 ;
      RECT 4.305 -67.195 4.445 -67.025 ;
      RECT 4.355 -66.008 4.445 -65 ;
      RECT 4.305 -65.405 4.445 -65.235 ;
      RECT 4.355 -64.2 4.445 -63.192 ;
      RECT 4.305 -63.965 4.445 -63.795 ;
      RECT 4.355 -62.778 4.445 -61.77 ;
      RECT 4.305 -62.175 4.445 -62.005 ;
      RECT 4.355 -60.97 4.445 -59.962 ;
      RECT 4.305 -60.735 4.445 -60.565 ;
      RECT 4.355 -59.548 4.445 -58.54 ;
      RECT 4.305 -58.945 4.445 -58.775 ;
      RECT 4.355 -57.74 4.445 -56.732 ;
      RECT 4.305 -57.505 4.445 -57.335 ;
      RECT 4.355 -56.318 4.445 -55.31 ;
      RECT 4.305 -55.715 4.445 -55.545 ;
      RECT 4.355 -54.51 4.445 -53.502 ;
      RECT 4.305 -54.275 4.445 -54.105 ;
      RECT 4.355 -53.088 4.445 -52.08 ;
      RECT 4.305 -52.485 4.445 -52.315 ;
      RECT 4.355 -51.28 4.445 -50.272 ;
      RECT 4.305 -51.045 4.445 -50.875 ;
      RECT 4.355 -49.858 4.445 -48.85 ;
      RECT 4.305 -49.255 4.445 -49.085 ;
      RECT 4.355 -48.05 4.445 -47.042 ;
      RECT 4.305 -47.815 4.445 -47.645 ;
      RECT 4.355 -46.628 4.445 -45.62 ;
      RECT 4.305 -46.025 4.445 -45.855 ;
      RECT 4.355 -44.82 4.445 -43.812 ;
      RECT 4.305 -44.585 4.445 -44.415 ;
      RECT 4.355 -43.398 4.445 -42.39 ;
      RECT 4.305 -42.795 4.445 -42.625 ;
      RECT 4.355 -41.59 4.445 -40.582 ;
      RECT 4.305 -41.355 4.445 -41.185 ;
      RECT 4.355 -40.168 4.445 -39.16 ;
      RECT 4.305 -39.565 4.445 -39.395 ;
      RECT 4.355 -38.36 4.445 -37.352 ;
      RECT 4.305 -38.125 4.445 -37.955 ;
      RECT 4.355 -36.938 4.445 -35.93 ;
      RECT 4.305 -36.335 4.445 -36.165 ;
      RECT 4.355 -35.13 4.445 -34.122 ;
      RECT 4.305 -34.895 4.445 -34.725 ;
      RECT 4.355 -33.708 4.445 -32.7 ;
      RECT 4.305 -33.105 4.445 -32.935 ;
      RECT 4.355 -31.9 4.445 -30.892 ;
      RECT 4.305 -31.665 4.445 -31.495 ;
      RECT 4.355 -30.478 4.445 -29.47 ;
      RECT 4.305 -29.875 4.445 -29.705 ;
      RECT 4.355 -28.67 4.445 -27.662 ;
      RECT 4.305 -28.435 4.445 -28.265 ;
      RECT 4.355 -27.248 4.445 -26.24 ;
      RECT 4.305 -26.645 4.445 -26.475 ;
      RECT 4.355 -25.44 4.445 -24.432 ;
      RECT 4.305 -25.205 4.445 -25.035 ;
      RECT 4.355 -24.018 4.445 -23.01 ;
      RECT 4.305 -23.415 4.445 -23.245 ;
      RECT 4.355 -22.21 4.445 -21.202 ;
      RECT 4.305 -21.975 4.445 -21.805 ;
      RECT 4.355 -20.788 4.445 -19.78 ;
      RECT 4.305 -20.185 4.445 -20.015 ;
      RECT 4.355 -18.98 4.445 -17.972 ;
      RECT 4.305 -18.745 4.445 -18.575 ;
      RECT 4.355 -17.558 4.445 -16.55 ;
      RECT 4.305 -16.955 4.445 -16.785 ;
      RECT 4.355 -15.75 4.445 -14.742 ;
      RECT 4.305 -15.515 4.445 -15.345 ;
      RECT 4.355 -14.328 4.445 -13.32 ;
      RECT 4.305 -13.725 4.445 -13.555 ;
      RECT 4.355 -12.52 4.445 -11.512 ;
      RECT 4.305 -12.285 4.445 -12.115 ;
      RECT 4.355 -11.098 4.445 -10.09 ;
      RECT 4.305 -10.495 4.445 -10.325 ;
      RECT 4.355 -9.29 4.445 -8.282 ;
      RECT 4.305 -9.055 4.445 -8.885 ;
      RECT 4.355 -7.868 4.445 -6.86 ;
      RECT 4.305 -7.265 4.445 -7.095 ;
      RECT 4.355 -6.06 4.445 -5.052 ;
      RECT 4.305 -5.825 4.445 -5.655 ;
      RECT 4.355 -4.638 4.445 -3.63 ;
      RECT 4.305 -4.035 4.445 -3.865 ;
      RECT 4.355 -2.83 4.445 -1.822 ;
      RECT 4.305 -2.595 4.445 -2.425 ;
      RECT 4.355 -1.408 4.445 -0.4 ;
      RECT 4.305 -0.805 4.445 -0.635 ;
      RECT 4.355 0.4 4.445 1.408 ;
      RECT 4.305 0.635 4.445 0.805 ;
      RECT 2.925 -111.685 4.405 -111.585 ;
      RECT 2.925 -112.195 3.025 -111.585 ;
      RECT 3.145 -109.15 4.405 -109.05 ;
      RECT 4.305 -109.475 4.405 -109.05 ;
      RECT 3.745 -109.475 3.845 -109.05 ;
      RECT 3.185 -109.475 3.285 -109.05 ;
      RECT 3.955 -101.538 4.045 -100.531 ;
      RECT 3.955 -101.225 4.095 -101.055 ;
      RECT 3.955 -99.729 4.045 -98.722 ;
      RECT 3.955 -99.205 4.095 -99.035 ;
      RECT 3.955 -98.308 4.045 -97.301 ;
      RECT 3.955 -97.995 4.095 -97.825 ;
      RECT 3.955 -96.499 4.045 -95.492 ;
      RECT 3.955 -95.975 4.095 -95.805 ;
      RECT 3.955 -95.078 4.045 -94.071 ;
      RECT 3.955 -94.765 4.095 -94.595 ;
      RECT 3.955 -93.269 4.045 -92.262 ;
      RECT 3.955 -92.745 4.095 -92.575 ;
      RECT 3.955 -91.848 4.045 -90.841 ;
      RECT 3.955 -91.535 4.095 -91.365 ;
      RECT 3.955 -90.039 4.045 -89.032 ;
      RECT 3.955 -89.515 4.095 -89.345 ;
      RECT 3.955 -88.618 4.045 -87.611 ;
      RECT 3.955 -88.305 4.095 -88.135 ;
      RECT 3.955 -86.809 4.045 -85.802 ;
      RECT 3.955 -86.285 4.095 -86.115 ;
      RECT 3.955 -85.388 4.045 -84.381 ;
      RECT 3.955 -85.075 4.095 -84.905 ;
      RECT 3.955 -83.579 4.045 -82.572 ;
      RECT 3.955 -83.055 4.095 -82.885 ;
      RECT 3.955 -82.158 4.045 -81.151 ;
      RECT 3.955 -81.845 4.095 -81.675 ;
      RECT 3.955 -80.349 4.045 -79.342 ;
      RECT 3.955 -79.825 4.095 -79.655 ;
      RECT 3.955 -78.928 4.045 -77.921 ;
      RECT 3.955 -78.615 4.095 -78.445 ;
      RECT 3.955 -77.119 4.045 -76.112 ;
      RECT 3.955 -76.595 4.095 -76.425 ;
      RECT 3.955 -75.698 4.045 -74.691 ;
      RECT 3.955 -75.385 4.095 -75.215 ;
      RECT 3.955 -73.889 4.045 -72.882 ;
      RECT 3.955 -73.365 4.095 -73.195 ;
      RECT 3.955 -72.468 4.045 -71.461 ;
      RECT 3.955 -72.155 4.095 -71.985 ;
      RECT 3.955 -70.659 4.045 -69.652 ;
      RECT 3.955 -70.135 4.095 -69.965 ;
      RECT 3.955 -69.238 4.045 -68.231 ;
      RECT 3.955 -68.925 4.095 -68.755 ;
      RECT 3.955 -67.429 4.045 -66.422 ;
      RECT 3.955 -66.905 4.095 -66.735 ;
      RECT 3.955 -66.008 4.045 -65.001 ;
      RECT 3.955 -65.695 4.095 -65.525 ;
      RECT 3.955 -64.199 4.045 -63.192 ;
      RECT 3.955 -63.675 4.095 -63.505 ;
      RECT 3.955 -62.778 4.045 -61.771 ;
      RECT 3.955 -62.465 4.095 -62.295 ;
      RECT 3.955 -60.969 4.045 -59.962 ;
      RECT 3.955 -60.445 4.095 -60.275 ;
      RECT 3.955 -59.548 4.045 -58.541 ;
      RECT 3.955 -59.235 4.095 -59.065 ;
      RECT 3.955 -57.739 4.045 -56.732 ;
      RECT 3.955 -57.215 4.095 -57.045 ;
      RECT 3.955 -56.318 4.045 -55.311 ;
      RECT 3.955 -56.005 4.095 -55.835 ;
      RECT 3.955 -54.509 4.045 -53.502 ;
      RECT 3.955 -53.985 4.095 -53.815 ;
      RECT 3.955 -53.088 4.045 -52.081 ;
      RECT 3.955 -52.775 4.095 -52.605 ;
      RECT 3.955 -51.279 4.045 -50.272 ;
      RECT 3.955 -50.755 4.095 -50.585 ;
      RECT 3.955 -49.858 4.045 -48.851 ;
      RECT 3.955 -49.545 4.095 -49.375 ;
      RECT 3.955 -48.049 4.045 -47.042 ;
      RECT 3.955 -47.525 4.095 -47.355 ;
      RECT 3.955 -46.628 4.045 -45.621 ;
      RECT 3.955 -46.315 4.095 -46.145 ;
      RECT 3.955 -44.819 4.045 -43.812 ;
      RECT 3.955 -44.295 4.095 -44.125 ;
      RECT 3.955 -43.398 4.045 -42.391 ;
      RECT 3.955 -43.085 4.095 -42.915 ;
      RECT 3.955 -41.589 4.045 -40.582 ;
      RECT 3.955 -41.065 4.095 -40.895 ;
      RECT 3.955 -40.168 4.045 -39.161 ;
      RECT 3.955 -39.855 4.095 -39.685 ;
      RECT 3.955 -38.359 4.045 -37.352 ;
      RECT 3.955 -37.835 4.095 -37.665 ;
      RECT 3.955 -36.938 4.045 -35.931 ;
      RECT 3.955 -36.625 4.095 -36.455 ;
      RECT 3.955 -35.129 4.045 -34.122 ;
      RECT 3.955 -34.605 4.095 -34.435 ;
      RECT 3.955 -33.708 4.045 -32.701 ;
      RECT 3.955 -33.395 4.095 -33.225 ;
      RECT 3.955 -31.899 4.045 -30.892 ;
      RECT 3.955 -31.375 4.095 -31.205 ;
      RECT 3.955 -30.478 4.045 -29.471 ;
      RECT 3.955 -30.165 4.095 -29.995 ;
      RECT 3.955 -28.669 4.045 -27.662 ;
      RECT 3.955 -28.145 4.095 -27.975 ;
      RECT 3.955 -27.248 4.045 -26.241 ;
      RECT 3.955 -26.935 4.095 -26.765 ;
      RECT 3.955 -25.439 4.045 -24.432 ;
      RECT 3.955 -24.915 4.095 -24.745 ;
      RECT 3.955 -24.018 4.045 -23.011 ;
      RECT 3.955 -23.705 4.095 -23.535 ;
      RECT 3.955 -22.209 4.045 -21.202 ;
      RECT 3.955 -21.685 4.095 -21.515 ;
      RECT 3.955 -20.788 4.045 -19.781 ;
      RECT 3.955 -20.475 4.095 -20.305 ;
      RECT 3.955 -18.979 4.045 -17.972 ;
      RECT 3.955 -18.455 4.095 -18.285 ;
      RECT 3.955 -17.558 4.045 -16.551 ;
      RECT 3.955 -17.245 4.095 -17.075 ;
      RECT 3.955 -15.749 4.045 -14.742 ;
      RECT 3.955 -15.225 4.095 -15.055 ;
      RECT 3.955 -14.328 4.045 -13.321 ;
      RECT 3.955 -14.015 4.095 -13.845 ;
      RECT 3.955 -12.519 4.045 -11.512 ;
      RECT 3.955 -11.995 4.095 -11.825 ;
      RECT 3.955 -11.098 4.045 -10.091 ;
      RECT 3.955 -10.785 4.095 -10.615 ;
      RECT 3.955 -9.289 4.045 -8.282 ;
      RECT 3.955 -8.765 4.095 -8.595 ;
      RECT 3.955 -7.868 4.045 -6.861 ;
      RECT 3.955 -7.555 4.095 -7.385 ;
      RECT 3.955 -6.059 4.045 -5.052 ;
      RECT 3.955 -5.535 4.095 -5.365 ;
      RECT 3.955 -4.638 4.045 -3.631 ;
      RECT 3.955 -4.325 4.095 -4.155 ;
      RECT 3.955 -2.829 4.045 -1.822 ;
      RECT 3.955 -2.305 4.095 -2.135 ;
      RECT 3.955 -1.408 4.045 -0.401 ;
      RECT 3.955 -1.095 4.095 -0.925 ;
      RECT 3.955 0.401 4.045 1.408 ;
      RECT 3.955 0.925 4.095 1.095 ;
      RECT 3.285 -111.495 3.455 -111.385 ;
      RECT 0.135 -111.495 3.455 -111.395 ;
      RECT 3.155 -101.538 3.245 -100.53 ;
      RECT 3.105 -100.935 3.245 -100.765 ;
      RECT 3.155 -99.73 3.245 -98.722 ;
      RECT 3.105 -99.495 3.245 -99.325 ;
      RECT 3.155 -98.308 3.245 -97.3 ;
      RECT 3.105 -97.705 3.245 -97.535 ;
      RECT 3.155 -96.5 3.245 -95.492 ;
      RECT 3.105 -96.265 3.245 -96.095 ;
      RECT 3.155 -95.078 3.245 -94.07 ;
      RECT 3.105 -94.475 3.245 -94.305 ;
      RECT 3.155 -93.27 3.245 -92.262 ;
      RECT 3.105 -93.035 3.245 -92.865 ;
      RECT 3.155 -91.848 3.245 -90.84 ;
      RECT 3.105 -91.245 3.245 -91.075 ;
      RECT 3.155 -90.04 3.245 -89.032 ;
      RECT 3.105 -89.805 3.245 -89.635 ;
      RECT 3.155 -88.618 3.245 -87.61 ;
      RECT 3.105 -88.015 3.245 -87.845 ;
      RECT 3.155 -86.81 3.245 -85.802 ;
      RECT 3.105 -86.575 3.245 -86.405 ;
      RECT 3.155 -85.388 3.245 -84.38 ;
      RECT 3.105 -84.785 3.245 -84.615 ;
      RECT 3.155 -83.58 3.245 -82.572 ;
      RECT 3.105 -83.345 3.245 -83.175 ;
      RECT 3.155 -82.158 3.245 -81.15 ;
      RECT 3.105 -81.555 3.245 -81.385 ;
      RECT 3.155 -80.35 3.245 -79.342 ;
      RECT 3.105 -80.115 3.245 -79.945 ;
      RECT 3.155 -78.928 3.245 -77.92 ;
      RECT 3.105 -78.325 3.245 -78.155 ;
      RECT 3.155 -77.12 3.245 -76.112 ;
      RECT 3.105 -76.885 3.245 -76.715 ;
      RECT 3.155 -75.698 3.245 -74.69 ;
      RECT 3.105 -75.095 3.245 -74.925 ;
      RECT 3.155 -73.89 3.245 -72.882 ;
      RECT 3.105 -73.655 3.245 -73.485 ;
      RECT 3.155 -72.468 3.245 -71.46 ;
      RECT 3.105 -71.865 3.245 -71.695 ;
      RECT 3.155 -70.66 3.245 -69.652 ;
      RECT 3.105 -70.425 3.245 -70.255 ;
      RECT 3.155 -69.238 3.245 -68.23 ;
      RECT 3.105 -68.635 3.245 -68.465 ;
      RECT 3.155 -67.43 3.245 -66.422 ;
      RECT 3.105 -67.195 3.245 -67.025 ;
      RECT 3.155 -66.008 3.245 -65 ;
      RECT 3.105 -65.405 3.245 -65.235 ;
      RECT 3.155 -64.2 3.245 -63.192 ;
      RECT 3.105 -63.965 3.245 -63.795 ;
      RECT 3.155 -62.778 3.245 -61.77 ;
      RECT 3.105 -62.175 3.245 -62.005 ;
      RECT 3.155 -60.97 3.245 -59.962 ;
      RECT 3.105 -60.735 3.245 -60.565 ;
      RECT 3.155 -59.548 3.245 -58.54 ;
      RECT 3.105 -58.945 3.245 -58.775 ;
      RECT 3.155 -57.74 3.245 -56.732 ;
      RECT 3.105 -57.505 3.245 -57.335 ;
      RECT 3.155 -56.318 3.245 -55.31 ;
      RECT 3.105 -55.715 3.245 -55.545 ;
      RECT 3.155 -54.51 3.245 -53.502 ;
      RECT 3.105 -54.275 3.245 -54.105 ;
      RECT 3.155 -53.088 3.245 -52.08 ;
      RECT 3.105 -52.485 3.245 -52.315 ;
      RECT 3.155 -51.28 3.245 -50.272 ;
      RECT 3.105 -51.045 3.245 -50.875 ;
      RECT 3.155 -49.858 3.245 -48.85 ;
      RECT 3.105 -49.255 3.245 -49.085 ;
      RECT 3.155 -48.05 3.245 -47.042 ;
      RECT 3.105 -47.815 3.245 -47.645 ;
      RECT 3.155 -46.628 3.245 -45.62 ;
      RECT 3.105 -46.025 3.245 -45.855 ;
      RECT 3.155 -44.82 3.245 -43.812 ;
      RECT 3.105 -44.585 3.245 -44.415 ;
      RECT 3.155 -43.398 3.245 -42.39 ;
      RECT 3.105 -42.795 3.245 -42.625 ;
      RECT 3.155 -41.59 3.245 -40.582 ;
      RECT 3.105 -41.355 3.245 -41.185 ;
      RECT 3.155 -40.168 3.245 -39.16 ;
      RECT 3.105 -39.565 3.245 -39.395 ;
      RECT 3.155 -38.36 3.245 -37.352 ;
      RECT 3.105 -38.125 3.245 -37.955 ;
      RECT 3.155 -36.938 3.245 -35.93 ;
      RECT 3.105 -36.335 3.245 -36.165 ;
      RECT 3.155 -35.13 3.245 -34.122 ;
      RECT 3.105 -34.895 3.245 -34.725 ;
      RECT 3.155 -33.708 3.245 -32.7 ;
      RECT 3.105 -33.105 3.245 -32.935 ;
      RECT 3.155 -31.9 3.245 -30.892 ;
      RECT 3.105 -31.665 3.245 -31.495 ;
      RECT 3.155 -30.478 3.245 -29.47 ;
      RECT 3.105 -29.875 3.245 -29.705 ;
      RECT 3.155 -28.67 3.245 -27.662 ;
      RECT 3.105 -28.435 3.245 -28.265 ;
      RECT 3.155 -27.248 3.245 -26.24 ;
      RECT 3.105 -26.645 3.245 -26.475 ;
      RECT 3.155 -25.44 3.245 -24.432 ;
      RECT 3.105 -25.205 3.245 -25.035 ;
      RECT 3.155 -24.018 3.245 -23.01 ;
      RECT 3.105 -23.415 3.245 -23.245 ;
      RECT 3.155 -22.21 3.245 -21.202 ;
      RECT 3.105 -21.975 3.245 -21.805 ;
      RECT 3.155 -20.788 3.245 -19.78 ;
      RECT 3.105 -20.185 3.245 -20.015 ;
      RECT 3.155 -18.98 3.245 -17.972 ;
      RECT 3.105 -18.745 3.245 -18.575 ;
      RECT 3.155 -17.558 3.245 -16.55 ;
      RECT 3.105 -16.955 3.245 -16.785 ;
      RECT 3.155 -15.75 3.245 -14.742 ;
      RECT 3.105 -15.515 3.245 -15.345 ;
      RECT 3.155 -14.328 3.245 -13.32 ;
      RECT 3.105 -13.725 3.245 -13.555 ;
      RECT 3.155 -12.52 3.245 -11.512 ;
      RECT 3.105 -12.285 3.245 -12.115 ;
      RECT 3.155 -11.098 3.245 -10.09 ;
      RECT 3.105 -10.495 3.245 -10.325 ;
      RECT 3.155 -9.29 3.245 -8.282 ;
      RECT 3.105 -9.055 3.245 -8.885 ;
      RECT 3.155 -7.868 3.245 -6.86 ;
      RECT 3.105 -7.265 3.245 -7.095 ;
      RECT 3.155 -6.06 3.245 -5.052 ;
      RECT 3.105 -5.825 3.245 -5.655 ;
      RECT 3.155 -4.638 3.245 -3.63 ;
      RECT 3.105 -4.035 3.245 -3.865 ;
      RECT 3.155 -2.83 3.245 -1.822 ;
      RECT 3.105 -2.595 3.245 -2.425 ;
      RECT 3.155 -1.408 3.245 -0.4 ;
      RECT 3.105 -0.805 3.245 -0.635 ;
      RECT 3.155 0.4 3.245 1.408 ;
      RECT 3.105 0.635 3.245 0.805 ;
      RECT 2.755 -101.538 2.845 -100.531 ;
      RECT 2.755 -101.225 2.895 -101.055 ;
      RECT 2.755 -99.729 2.845 -98.722 ;
      RECT 2.755 -99.205 2.895 -99.035 ;
      RECT 2.755 -98.308 2.845 -97.301 ;
      RECT 2.755 -97.995 2.895 -97.825 ;
      RECT 2.755 -96.499 2.845 -95.492 ;
      RECT 2.755 -95.975 2.895 -95.805 ;
      RECT 2.755 -95.078 2.845 -94.071 ;
      RECT 2.755 -94.765 2.895 -94.595 ;
      RECT 2.755 -93.269 2.845 -92.262 ;
      RECT 2.755 -92.745 2.895 -92.575 ;
      RECT 2.755 -91.848 2.845 -90.841 ;
      RECT 2.755 -91.535 2.895 -91.365 ;
      RECT 2.755 -90.039 2.845 -89.032 ;
      RECT 2.755 -89.515 2.895 -89.345 ;
      RECT 2.755 -88.618 2.845 -87.611 ;
      RECT 2.755 -88.305 2.895 -88.135 ;
      RECT 2.755 -86.809 2.845 -85.802 ;
      RECT 2.755 -86.285 2.895 -86.115 ;
      RECT 2.755 -85.388 2.845 -84.381 ;
      RECT 2.755 -85.075 2.895 -84.905 ;
      RECT 2.755 -83.579 2.845 -82.572 ;
      RECT 2.755 -83.055 2.895 -82.885 ;
      RECT 2.755 -82.158 2.845 -81.151 ;
      RECT 2.755 -81.845 2.895 -81.675 ;
      RECT 2.755 -80.349 2.845 -79.342 ;
      RECT 2.755 -79.825 2.895 -79.655 ;
      RECT 2.755 -78.928 2.845 -77.921 ;
      RECT 2.755 -78.615 2.895 -78.445 ;
      RECT 2.755 -77.119 2.845 -76.112 ;
      RECT 2.755 -76.595 2.895 -76.425 ;
      RECT 2.755 -75.698 2.845 -74.691 ;
      RECT 2.755 -75.385 2.895 -75.215 ;
      RECT 2.755 -73.889 2.845 -72.882 ;
      RECT 2.755 -73.365 2.895 -73.195 ;
      RECT 2.755 -72.468 2.845 -71.461 ;
      RECT 2.755 -72.155 2.895 -71.985 ;
      RECT 2.755 -70.659 2.845 -69.652 ;
      RECT 2.755 -70.135 2.895 -69.965 ;
      RECT 2.755 -69.238 2.845 -68.231 ;
      RECT 2.755 -68.925 2.895 -68.755 ;
      RECT 2.755 -67.429 2.845 -66.422 ;
      RECT 2.755 -66.905 2.895 -66.735 ;
      RECT 2.755 -66.008 2.845 -65.001 ;
      RECT 2.755 -65.695 2.895 -65.525 ;
      RECT 2.755 -64.199 2.845 -63.192 ;
      RECT 2.755 -63.675 2.895 -63.505 ;
      RECT 2.755 -62.778 2.845 -61.771 ;
      RECT 2.755 -62.465 2.895 -62.295 ;
      RECT 2.755 -60.969 2.845 -59.962 ;
      RECT 2.755 -60.445 2.895 -60.275 ;
      RECT 2.755 -59.548 2.845 -58.541 ;
      RECT 2.755 -59.235 2.895 -59.065 ;
      RECT 2.755 -57.739 2.845 -56.732 ;
      RECT 2.755 -57.215 2.895 -57.045 ;
      RECT 2.755 -56.318 2.845 -55.311 ;
      RECT 2.755 -56.005 2.895 -55.835 ;
      RECT 2.755 -54.509 2.845 -53.502 ;
      RECT 2.755 -53.985 2.895 -53.815 ;
      RECT 2.755 -53.088 2.845 -52.081 ;
      RECT 2.755 -52.775 2.895 -52.605 ;
      RECT 2.755 -51.279 2.845 -50.272 ;
      RECT 2.755 -50.755 2.895 -50.585 ;
      RECT 2.755 -49.858 2.845 -48.851 ;
      RECT 2.755 -49.545 2.895 -49.375 ;
      RECT 2.755 -48.049 2.845 -47.042 ;
      RECT 2.755 -47.525 2.895 -47.355 ;
      RECT 2.755 -46.628 2.845 -45.621 ;
      RECT 2.755 -46.315 2.895 -46.145 ;
      RECT 2.755 -44.819 2.845 -43.812 ;
      RECT 2.755 -44.295 2.895 -44.125 ;
      RECT 2.755 -43.398 2.845 -42.391 ;
      RECT 2.755 -43.085 2.895 -42.915 ;
      RECT 2.755 -41.589 2.845 -40.582 ;
      RECT 2.755 -41.065 2.895 -40.895 ;
      RECT 2.755 -40.168 2.845 -39.161 ;
      RECT 2.755 -39.855 2.895 -39.685 ;
      RECT 2.755 -38.359 2.845 -37.352 ;
      RECT 2.755 -37.835 2.895 -37.665 ;
      RECT 2.755 -36.938 2.845 -35.931 ;
      RECT 2.755 -36.625 2.895 -36.455 ;
      RECT 2.755 -35.129 2.845 -34.122 ;
      RECT 2.755 -34.605 2.895 -34.435 ;
      RECT 2.755 -33.708 2.845 -32.701 ;
      RECT 2.755 -33.395 2.895 -33.225 ;
      RECT 2.755 -31.899 2.845 -30.892 ;
      RECT 2.755 -31.375 2.895 -31.205 ;
      RECT 2.755 -30.478 2.845 -29.471 ;
      RECT 2.755 -30.165 2.895 -29.995 ;
      RECT 2.755 -28.669 2.845 -27.662 ;
      RECT 2.755 -28.145 2.895 -27.975 ;
      RECT 2.755 -27.248 2.845 -26.241 ;
      RECT 2.755 -26.935 2.895 -26.765 ;
      RECT 2.755 -25.439 2.845 -24.432 ;
      RECT 2.755 -24.915 2.895 -24.745 ;
      RECT 2.755 -24.018 2.845 -23.011 ;
      RECT 2.755 -23.705 2.895 -23.535 ;
      RECT 2.755 -22.209 2.845 -21.202 ;
      RECT 2.755 -21.685 2.895 -21.515 ;
      RECT 2.755 -20.788 2.845 -19.781 ;
      RECT 2.755 -20.475 2.895 -20.305 ;
      RECT 2.755 -18.979 2.845 -17.972 ;
      RECT 2.755 -18.455 2.895 -18.285 ;
      RECT 2.755 -17.558 2.845 -16.551 ;
      RECT 2.755 -17.245 2.895 -17.075 ;
      RECT 2.755 -15.749 2.845 -14.742 ;
      RECT 2.755 -15.225 2.895 -15.055 ;
      RECT 2.755 -14.328 2.845 -13.321 ;
      RECT 2.755 -14.015 2.895 -13.845 ;
      RECT 2.755 -12.519 2.845 -11.512 ;
      RECT 2.755 -11.995 2.895 -11.825 ;
      RECT 2.755 -11.098 2.845 -10.091 ;
      RECT 2.755 -10.785 2.895 -10.615 ;
      RECT 2.755 -9.289 2.845 -8.282 ;
      RECT 2.755 -8.765 2.895 -8.595 ;
      RECT 2.755 -7.868 2.845 -6.861 ;
      RECT 2.755 -7.555 2.895 -7.385 ;
      RECT 2.755 -6.059 2.845 -5.052 ;
      RECT 2.755 -5.535 2.895 -5.365 ;
      RECT 2.755 -4.638 2.845 -3.631 ;
      RECT 2.755 -4.325 2.895 -4.155 ;
      RECT 2.755 -2.829 2.845 -1.822 ;
      RECT 2.755 -2.305 2.895 -2.135 ;
      RECT 2.755 -1.408 2.845 -0.401 ;
      RECT 2.755 -1.095 2.895 -0.925 ;
      RECT 2.755 0.401 2.845 1.408 ;
      RECT 2.755 0.925 2.895 1.095 ;
      RECT 0.905 -111.685 2.385 -111.585 ;
      RECT 0.905 -112.055 1.005 -111.585 ;
      RECT 0.71 -114.395 2.285 -114.275 ;
      RECT 2.185 -114.895 2.285 -114.275 ;
      RECT 1.59 -114.895 1.69 -114.275 ;
      RECT 0.71 -114.85 0.81 -114.275 ;
      RECT 1.955 -101.538 2.045 -100.53 ;
      RECT 1.905 -100.935 2.045 -100.765 ;
      RECT 1.955 -99.73 2.045 -98.722 ;
      RECT 1.905 -99.495 2.045 -99.325 ;
      RECT 1.955 -98.308 2.045 -97.3 ;
      RECT 1.905 -97.705 2.045 -97.535 ;
      RECT 1.955 -96.5 2.045 -95.492 ;
      RECT 1.905 -96.265 2.045 -96.095 ;
      RECT 1.955 -95.078 2.045 -94.07 ;
      RECT 1.905 -94.475 2.045 -94.305 ;
      RECT 1.955 -93.27 2.045 -92.262 ;
      RECT 1.905 -93.035 2.045 -92.865 ;
      RECT 1.955 -91.848 2.045 -90.84 ;
      RECT 1.905 -91.245 2.045 -91.075 ;
      RECT 1.955 -90.04 2.045 -89.032 ;
      RECT 1.905 -89.805 2.045 -89.635 ;
      RECT 1.955 -88.618 2.045 -87.61 ;
      RECT 1.905 -88.015 2.045 -87.845 ;
      RECT 1.955 -86.81 2.045 -85.802 ;
      RECT 1.905 -86.575 2.045 -86.405 ;
      RECT 1.955 -85.388 2.045 -84.38 ;
      RECT 1.905 -84.785 2.045 -84.615 ;
      RECT 1.955 -83.58 2.045 -82.572 ;
      RECT 1.905 -83.345 2.045 -83.175 ;
      RECT 1.955 -82.158 2.045 -81.15 ;
      RECT 1.905 -81.555 2.045 -81.385 ;
      RECT 1.955 -80.35 2.045 -79.342 ;
      RECT 1.905 -80.115 2.045 -79.945 ;
      RECT 1.955 -78.928 2.045 -77.92 ;
      RECT 1.905 -78.325 2.045 -78.155 ;
      RECT 1.955 -77.12 2.045 -76.112 ;
      RECT 1.905 -76.885 2.045 -76.715 ;
      RECT 1.955 -75.698 2.045 -74.69 ;
      RECT 1.905 -75.095 2.045 -74.925 ;
      RECT 1.955 -73.89 2.045 -72.882 ;
      RECT 1.905 -73.655 2.045 -73.485 ;
      RECT 1.955 -72.468 2.045 -71.46 ;
      RECT 1.905 -71.865 2.045 -71.695 ;
      RECT 1.955 -70.66 2.045 -69.652 ;
      RECT 1.905 -70.425 2.045 -70.255 ;
      RECT 1.955 -69.238 2.045 -68.23 ;
      RECT 1.905 -68.635 2.045 -68.465 ;
      RECT 1.955 -67.43 2.045 -66.422 ;
      RECT 1.905 -67.195 2.045 -67.025 ;
      RECT 1.955 -66.008 2.045 -65 ;
      RECT 1.905 -65.405 2.045 -65.235 ;
      RECT 1.955 -64.2 2.045 -63.192 ;
      RECT 1.905 -63.965 2.045 -63.795 ;
      RECT 1.955 -62.778 2.045 -61.77 ;
      RECT 1.905 -62.175 2.045 -62.005 ;
      RECT 1.955 -60.97 2.045 -59.962 ;
      RECT 1.905 -60.735 2.045 -60.565 ;
      RECT 1.955 -59.548 2.045 -58.54 ;
      RECT 1.905 -58.945 2.045 -58.775 ;
      RECT 1.955 -57.74 2.045 -56.732 ;
      RECT 1.905 -57.505 2.045 -57.335 ;
      RECT 1.955 -56.318 2.045 -55.31 ;
      RECT 1.905 -55.715 2.045 -55.545 ;
      RECT 1.955 -54.51 2.045 -53.502 ;
      RECT 1.905 -54.275 2.045 -54.105 ;
      RECT 1.955 -53.088 2.045 -52.08 ;
      RECT 1.905 -52.485 2.045 -52.315 ;
      RECT 1.955 -51.28 2.045 -50.272 ;
      RECT 1.905 -51.045 2.045 -50.875 ;
      RECT 1.955 -49.858 2.045 -48.85 ;
      RECT 1.905 -49.255 2.045 -49.085 ;
      RECT 1.955 -48.05 2.045 -47.042 ;
      RECT 1.905 -47.815 2.045 -47.645 ;
      RECT 1.955 -46.628 2.045 -45.62 ;
      RECT 1.905 -46.025 2.045 -45.855 ;
      RECT 1.955 -44.82 2.045 -43.812 ;
      RECT 1.905 -44.585 2.045 -44.415 ;
      RECT 1.955 -43.398 2.045 -42.39 ;
      RECT 1.905 -42.795 2.045 -42.625 ;
      RECT 1.955 -41.59 2.045 -40.582 ;
      RECT 1.905 -41.355 2.045 -41.185 ;
      RECT 1.955 -40.168 2.045 -39.16 ;
      RECT 1.905 -39.565 2.045 -39.395 ;
      RECT 1.955 -38.36 2.045 -37.352 ;
      RECT 1.905 -38.125 2.045 -37.955 ;
      RECT 1.955 -36.938 2.045 -35.93 ;
      RECT 1.905 -36.335 2.045 -36.165 ;
      RECT 1.955 -35.13 2.045 -34.122 ;
      RECT 1.905 -34.895 2.045 -34.725 ;
      RECT 1.955 -33.708 2.045 -32.7 ;
      RECT 1.905 -33.105 2.045 -32.935 ;
      RECT 1.955 -31.9 2.045 -30.892 ;
      RECT 1.905 -31.665 2.045 -31.495 ;
      RECT 1.955 -30.478 2.045 -29.47 ;
      RECT 1.905 -29.875 2.045 -29.705 ;
      RECT 1.955 -28.67 2.045 -27.662 ;
      RECT 1.905 -28.435 2.045 -28.265 ;
      RECT 1.955 -27.248 2.045 -26.24 ;
      RECT 1.905 -26.645 2.045 -26.475 ;
      RECT 1.955 -25.44 2.045 -24.432 ;
      RECT 1.905 -25.205 2.045 -25.035 ;
      RECT 1.955 -24.018 2.045 -23.01 ;
      RECT 1.905 -23.415 2.045 -23.245 ;
      RECT 1.955 -22.21 2.045 -21.202 ;
      RECT 1.905 -21.975 2.045 -21.805 ;
      RECT 1.955 -20.788 2.045 -19.78 ;
      RECT 1.905 -20.185 2.045 -20.015 ;
      RECT 1.955 -18.98 2.045 -17.972 ;
      RECT 1.905 -18.745 2.045 -18.575 ;
      RECT 1.955 -17.558 2.045 -16.55 ;
      RECT 1.905 -16.955 2.045 -16.785 ;
      RECT 1.955 -15.75 2.045 -14.742 ;
      RECT 1.905 -15.515 2.045 -15.345 ;
      RECT 1.955 -14.328 2.045 -13.32 ;
      RECT 1.905 -13.725 2.045 -13.555 ;
      RECT 1.955 -12.52 2.045 -11.512 ;
      RECT 1.905 -12.285 2.045 -12.115 ;
      RECT 1.955 -11.098 2.045 -10.09 ;
      RECT 1.905 -10.495 2.045 -10.325 ;
      RECT 1.955 -9.29 2.045 -8.282 ;
      RECT 1.905 -9.055 2.045 -8.885 ;
      RECT 1.955 -7.868 2.045 -6.86 ;
      RECT 1.905 -7.265 2.045 -7.095 ;
      RECT 1.955 -6.06 2.045 -5.052 ;
      RECT 1.905 -5.825 2.045 -5.655 ;
      RECT 1.955 -4.638 2.045 -3.63 ;
      RECT 1.905 -4.035 2.045 -3.865 ;
      RECT 1.955 -2.83 2.045 -1.822 ;
      RECT 1.905 -2.595 2.045 -2.425 ;
      RECT 1.955 -1.408 2.045 -0.4 ;
      RECT 1.905 -0.805 2.045 -0.635 ;
      RECT 1.955 0.4 2.045 1.408 ;
      RECT 1.905 0.635 2.045 0.805 ;
      RECT 1.83 -114.685 2.005 -114.515 ;
      RECT 1.905 -114.895 2.005 -114.515 ;
      RECT 0.945 -113.555 1.045 -113.09 ;
      RECT 1.31 -113.555 1.41 -113.1 ;
      RECT 0.945 -113.555 1.79 -113.385 ;
      RECT 1.555 -101.538 1.645 -100.531 ;
      RECT 1.555 -101.225 1.695 -101.055 ;
      RECT 1.555 -99.729 1.645 -98.722 ;
      RECT 1.555 -99.205 1.695 -99.035 ;
      RECT 1.555 -98.308 1.645 -97.301 ;
      RECT 1.555 -97.995 1.695 -97.825 ;
      RECT 1.555 -96.499 1.645 -95.492 ;
      RECT 1.555 -95.975 1.695 -95.805 ;
      RECT 1.555 -95.078 1.645 -94.071 ;
      RECT 1.555 -94.765 1.695 -94.595 ;
      RECT 1.555 -93.269 1.645 -92.262 ;
      RECT 1.555 -92.745 1.695 -92.575 ;
      RECT 1.555 -91.848 1.645 -90.841 ;
      RECT 1.555 -91.535 1.695 -91.365 ;
      RECT 1.555 -90.039 1.645 -89.032 ;
      RECT 1.555 -89.515 1.695 -89.345 ;
      RECT 1.555 -88.618 1.645 -87.611 ;
      RECT 1.555 -88.305 1.695 -88.135 ;
      RECT 1.555 -86.809 1.645 -85.802 ;
      RECT 1.555 -86.285 1.695 -86.115 ;
      RECT 1.555 -85.388 1.645 -84.381 ;
      RECT 1.555 -85.075 1.695 -84.905 ;
      RECT 1.555 -83.579 1.645 -82.572 ;
      RECT 1.555 -83.055 1.695 -82.885 ;
      RECT 1.555 -82.158 1.645 -81.151 ;
      RECT 1.555 -81.845 1.695 -81.675 ;
      RECT 1.555 -80.349 1.645 -79.342 ;
      RECT 1.555 -79.825 1.695 -79.655 ;
      RECT 1.555 -78.928 1.645 -77.921 ;
      RECT 1.555 -78.615 1.695 -78.445 ;
      RECT 1.555 -77.119 1.645 -76.112 ;
      RECT 1.555 -76.595 1.695 -76.425 ;
      RECT 1.555 -75.698 1.645 -74.691 ;
      RECT 1.555 -75.385 1.695 -75.215 ;
      RECT 1.555 -73.889 1.645 -72.882 ;
      RECT 1.555 -73.365 1.695 -73.195 ;
      RECT 1.555 -72.468 1.645 -71.461 ;
      RECT 1.555 -72.155 1.695 -71.985 ;
      RECT 1.555 -70.659 1.645 -69.652 ;
      RECT 1.555 -70.135 1.695 -69.965 ;
      RECT 1.555 -69.238 1.645 -68.231 ;
      RECT 1.555 -68.925 1.695 -68.755 ;
      RECT 1.555 -67.429 1.645 -66.422 ;
      RECT 1.555 -66.905 1.695 -66.735 ;
      RECT 1.555 -66.008 1.645 -65.001 ;
      RECT 1.555 -65.695 1.695 -65.525 ;
      RECT 1.555 -64.199 1.645 -63.192 ;
      RECT 1.555 -63.675 1.695 -63.505 ;
      RECT 1.555 -62.778 1.645 -61.771 ;
      RECT 1.555 -62.465 1.695 -62.295 ;
      RECT 1.555 -60.969 1.645 -59.962 ;
      RECT 1.555 -60.445 1.695 -60.275 ;
      RECT 1.555 -59.548 1.645 -58.541 ;
      RECT 1.555 -59.235 1.695 -59.065 ;
      RECT 1.555 -57.739 1.645 -56.732 ;
      RECT 1.555 -57.215 1.695 -57.045 ;
      RECT 1.555 -56.318 1.645 -55.311 ;
      RECT 1.555 -56.005 1.695 -55.835 ;
      RECT 1.555 -54.509 1.645 -53.502 ;
      RECT 1.555 -53.985 1.695 -53.815 ;
      RECT 1.555 -53.088 1.645 -52.081 ;
      RECT 1.555 -52.775 1.695 -52.605 ;
      RECT 1.555 -51.279 1.645 -50.272 ;
      RECT 1.555 -50.755 1.695 -50.585 ;
      RECT 1.555 -49.858 1.645 -48.851 ;
      RECT 1.555 -49.545 1.695 -49.375 ;
      RECT 1.555 -48.049 1.645 -47.042 ;
      RECT 1.555 -47.525 1.695 -47.355 ;
      RECT 1.555 -46.628 1.645 -45.621 ;
      RECT 1.555 -46.315 1.695 -46.145 ;
      RECT 1.555 -44.819 1.645 -43.812 ;
      RECT 1.555 -44.295 1.695 -44.125 ;
      RECT 1.555 -43.398 1.645 -42.391 ;
      RECT 1.555 -43.085 1.695 -42.915 ;
      RECT 1.555 -41.589 1.645 -40.582 ;
      RECT 1.555 -41.065 1.695 -40.895 ;
      RECT 1.555 -40.168 1.645 -39.161 ;
      RECT 1.555 -39.855 1.695 -39.685 ;
      RECT 1.555 -38.359 1.645 -37.352 ;
      RECT 1.555 -37.835 1.695 -37.665 ;
      RECT 1.555 -36.938 1.645 -35.931 ;
      RECT 1.555 -36.625 1.695 -36.455 ;
      RECT 1.555 -35.129 1.645 -34.122 ;
      RECT 1.555 -34.605 1.695 -34.435 ;
      RECT 1.555 -33.708 1.645 -32.701 ;
      RECT 1.555 -33.395 1.695 -33.225 ;
      RECT 1.555 -31.899 1.645 -30.892 ;
      RECT 1.555 -31.375 1.695 -31.205 ;
      RECT 1.555 -30.478 1.645 -29.471 ;
      RECT 1.555 -30.165 1.695 -29.995 ;
      RECT 1.555 -28.669 1.645 -27.662 ;
      RECT 1.555 -28.145 1.695 -27.975 ;
      RECT 1.555 -27.248 1.645 -26.241 ;
      RECT 1.555 -26.935 1.695 -26.765 ;
      RECT 1.555 -25.439 1.645 -24.432 ;
      RECT 1.555 -24.915 1.695 -24.745 ;
      RECT 1.555 -24.018 1.645 -23.011 ;
      RECT 1.555 -23.705 1.695 -23.535 ;
      RECT 1.555 -22.209 1.645 -21.202 ;
      RECT 1.555 -21.685 1.695 -21.515 ;
      RECT 1.555 -20.788 1.645 -19.781 ;
      RECT 1.555 -20.475 1.695 -20.305 ;
      RECT 1.555 -18.979 1.645 -17.972 ;
      RECT 1.555 -18.455 1.695 -18.285 ;
      RECT 1.555 -17.558 1.645 -16.551 ;
      RECT 1.555 -17.245 1.695 -17.075 ;
      RECT 1.555 -15.749 1.645 -14.742 ;
      RECT 1.555 -15.225 1.695 -15.055 ;
      RECT 1.555 -14.328 1.645 -13.321 ;
      RECT 1.555 -14.015 1.695 -13.845 ;
      RECT 1.555 -12.519 1.645 -11.512 ;
      RECT 1.555 -11.995 1.695 -11.825 ;
      RECT 1.555 -11.098 1.645 -10.091 ;
      RECT 1.555 -10.785 1.695 -10.615 ;
      RECT 1.555 -9.289 1.645 -8.282 ;
      RECT 1.555 -8.765 1.695 -8.595 ;
      RECT 1.555 -7.868 1.645 -6.861 ;
      RECT 1.555 -7.555 1.695 -7.385 ;
      RECT 1.555 -6.059 1.645 -5.052 ;
      RECT 1.555 -5.535 1.695 -5.365 ;
      RECT 1.555 -4.638 1.645 -3.631 ;
      RECT 1.555 -4.325 1.695 -4.155 ;
      RECT 1.555 -2.829 1.645 -1.822 ;
      RECT 1.555 -2.305 1.695 -2.135 ;
      RECT 1.555 -1.408 1.645 -0.401 ;
      RECT 1.555 -1.095 1.695 -0.925 ;
      RECT 1.555 0.401 1.645 1.408 ;
      RECT 1.555 0.925 1.695 1.095 ;
      RECT 1.24 -114.685 1.41 -114.515 ;
      RECT 1.31 -114.895 1.41 -114.515 ;
      RECT 0.755 -101.538 0.845 -100.53 ;
      RECT 0.705 -100.935 0.845 -100.765 ;
      RECT 0.755 -99.73 0.845 -98.722 ;
      RECT 0.705 -99.495 0.845 -99.325 ;
      RECT 0.755 -98.308 0.845 -97.3 ;
      RECT 0.705 -97.705 0.845 -97.535 ;
      RECT 0.755 -96.5 0.845 -95.492 ;
      RECT 0.705 -96.265 0.845 -96.095 ;
      RECT 0.755 -95.078 0.845 -94.07 ;
      RECT 0.705 -94.475 0.845 -94.305 ;
      RECT 0.755 -93.27 0.845 -92.262 ;
      RECT 0.705 -93.035 0.845 -92.865 ;
      RECT 0.755 -91.848 0.845 -90.84 ;
      RECT 0.705 -91.245 0.845 -91.075 ;
      RECT 0.755 -90.04 0.845 -89.032 ;
      RECT 0.705 -89.805 0.845 -89.635 ;
      RECT 0.755 -88.618 0.845 -87.61 ;
      RECT 0.705 -88.015 0.845 -87.845 ;
      RECT 0.755 -86.81 0.845 -85.802 ;
      RECT 0.705 -86.575 0.845 -86.405 ;
      RECT 0.755 -85.388 0.845 -84.38 ;
      RECT 0.705 -84.785 0.845 -84.615 ;
      RECT 0.755 -83.58 0.845 -82.572 ;
      RECT 0.705 -83.345 0.845 -83.175 ;
      RECT 0.755 -82.158 0.845 -81.15 ;
      RECT 0.705 -81.555 0.845 -81.385 ;
      RECT 0.755 -80.35 0.845 -79.342 ;
      RECT 0.705 -80.115 0.845 -79.945 ;
      RECT 0.755 -78.928 0.845 -77.92 ;
      RECT 0.705 -78.325 0.845 -78.155 ;
      RECT 0.755 -77.12 0.845 -76.112 ;
      RECT 0.705 -76.885 0.845 -76.715 ;
      RECT 0.755 -75.698 0.845 -74.69 ;
      RECT 0.705 -75.095 0.845 -74.925 ;
      RECT 0.755 -73.89 0.845 -72.882 ;
      RECT 0.705 -73.655 0.845 -73.485 ;
      RECT 0.755 -72.468 0.845 -71.46 ;
      RECT 0.705 -71.865 0.845 -71.695 ;
      RECT 0.755 -70.66 0.845 -69.652 ;
      RECT 0.705 -70.425 0.845 -70.255 ;
      RECT 0.755 -69.238 0.845 -68.23 ;
      RECT 0.705 -68.635 0.845 -68.465 ;
      RECT 0.755 -67.43 0.845 -66.422 ;
      RECT 0.705 -67.195 0.845 -67.025 ;
      RECT 0.755 -66.008 0.845 -65 ;
      RECT 0.705 -65.405 0.845 -65.235 ;
      RECT 0.755 -64.2 0.845 -63.192 ;
      RECT 0.705 -63.965 0.845 -63.795 ;
      RECT 0.755 -62.778 0.845 -61.77 ;
      RECT 0.705 -62.175 0.845 -62.005 ;
      RECT 0.755 -60.97 0.845 -59.962 ;
      RECT 0.705 -60.735 0.845 -60.565 ;
      RECT 0.755 -59.548 0.845 -58.54 ;
      RECT 0.705 -58.945 0.845 -58.775 ;
      RECT 0.755 -57.74 0.845 -56.732 ;
      RECT 0.705 -57.505 0.845 -57.335 ;
      RECT 0.755 -56.318 0.845 -55.31 ;
      RECT 0.705 -55.715 0.845 -55.545 ;
      RECT 0.755 -54.51 0.845 -53.502 ;
      RECT 0.705 -54.275 0.845 -54.105 ;
      RECT 0.755 -53.088 0.845 -52.08 ;
      RECT 0.705 -52.485 0.845 -52.315 ;
      RECT 0.755 -51.28 0.845 -50.272 ;
      RECT 0.705 -51.045 0.845 -50.875 ;
      RECT 0.755 -49.858 0.845 -48.85 ;
      RECT 0.705 -49.255 0.845 -49.085 ;
      RECT 0.755 -48.05 0.845 -47.042 ;
      RECT 0.705 -47.815 0.845 -47.645 ;
      RECT 0.755 -46.628 0.845 -45.62 ;
      RECT 0.705 -46.025 0.845 -45.855 ;
      RECT 0.755 -44.82 0.845 -43.812 ;
      RECT 0.705 -44.585 0.845 -44.415 ;
      RECT 0.755 -43.398 0.845 -42.39 ;
      RECT 0.705 -42.795 0.845 -42.625 ;
      RECT 0.755 -41.59 0.845 -40.582 ;
      RECT 0.705 -41.355 0.845 -41.185 ;
      RECT 0.755 -40.168 0.845 -39.16 ;
      RECT 0.705 -39.565 0.845 -39.395 ;
      RECT 0.755 -38.36 0.845 -37.352 ;
      RECT 0.705 -38.125 0.845 -37.955 ;
      RECT 0.755 -36.938 0.845 -35.93 ;
      RECT 0.705 -36.335 0.845 -36.165 ;
      RECT 0.755 -35.13 0.845 -34.122 ;
      RECT 0.705 -34.895 0.845 -34.725 ;
      RECT 0.755 -33.708 0.845 -32.7 ;
      RECT 0.705 -33.105 0.845 -32.935 ;
      RECT 0.755 -31.9 0.845 -30.892 ;
      RECT 0.705 -31.665 0.845 -31.495 ;
      RECT 0.755 -30.478 0.845 -29.47 ;
      RECT 0.705 -29.875 0.845 -29.705 ;
      RECT 0.755 -28.67 0.845 -27.662 ;
      RECT 0.705 -28.435 0.845 -28.265 ;
      RECT 0.755 -27.248 0.845 -26.24 ;
      RECT 0.705 -26.645 0.845 -26.475 ;
      RECT 0.755 -25.44 0.845 -24.432 ;
      RECT 0.705 -25.205 0.845 -25.035 ;
      RECT 0.755 -24.018 0.845 -23.01 ;
      RECT 0.705 -23.415 0.845 -23.245 ;
      RECT 0.755 -22.21 0.845 -21.202 ;
      RECT 0.705 -21.975 0.845 -21.805 ;
      RECT 0.755 -20.788 0.845 -19.78 ;
      RECT 0.705 -20.185 0.845 -20.015 ;
      RECT 0.755 -18.98 0.845 -17.972 ;
      RECT 0.705 -18.745 0.845 -18.575 ;
      RECT 0.755 -17.558 0.845 -16.55 ;
      RECT 0.705 -16.955 0.845 -16.785 ;
      RECT 0.755 -15.75 0.845 -14.742 ;
      RECT 0.705 -15.515 0.845 -15.345 ;
      RECT 0.755 -14.328 0.845 -13.32 ;
      RECT 0.705 -13.725 0.845 -13.555 ;
      RECT 0.755 -12.52 0.845 -11.512 ;
      RECT 0.705 -12.285 0.845 -12.115 ;
      RECT 0.755 -11.098 0.845 -10.09 ;
      RECT 0.705 -10.495 0.845 -10.325 ;
      RECT 0.755 -9.29 0.845 -8.282 ;
      RECT 0.705 -9.055 0.845 -8.885 ;
      RECT 0.755 -7.868 0.845 -6.86 ;
      RECT 0.705 -7.265 0.845 -7.095 ;
      RECT 0.755 -6.06 0.845 -5.052 ;
      RECT 0.705 -5.825 0.845 -5.655 ;
      RECT 0.755 -4.638 0.845 -3.63 ;
      RECT 0.705 -4.035 0.845 -3.865 ;
      RECT 0.755 -2.83 0.845 -1.822 ;
      RECT 0.705 -2.595 0.845 -2.425 ;
      RECT 0.755 -1.408 0.845 -0.4 ;
      RECT 0.705 -0.805 0.845 -0.635 ;
      RECT 0.755 0.4 0.845 1.408 ;
      RECT 0.705 0.635 0.845 0.805 ;
      RECT 0.355 -101.538 0.445 -100.531 ;
      RECT 0.355 -101.225 0.495 -101.055 ;
      RECT 0.355 -99.729 0.445 -98.722 ;
      RECT 0.355 -99.205 0.495 -99.035 ;
      RECT 0.355 -98.308 0.445 -97.301 ;
      RECT 0.355 -97.995 0.495 -97.825 ;
      RECT 0.355 -96.499 0.445 -95.492 ;
      RECT 0.355 -95.975 0.495 -95.805 ;
      RECT 0.355 -95.078 0.445 -94.071 ;
      RECT 0.355 -94.765 0.495 -94.595 ;
      RECT 0.355 -93.269 0.445 -92.262 ;
      RECT 0.355 -92.745 0.495 -92.575 ;
      RECT 0.355 -91.848 0.445 -90.841 ;
      RECT 0.355 -91.535 0.495 -91.365 ;
      RECT 0.355 -90.039 0.445 -89.032 ;
      RECT 0.355 -89.515 0.495 -89.345 ;
      RECT 0.355 -88.618 0.445 -87.611 ;
      RECT 0.355 -88.305 0.495 -88.135 ;
      RECT 0.355 -86.809 0.445 -85.802 ;
      RECT 0.355 -86.285 0.495 -86.115 ;
      RECT 0.355 -85.388 0.445 -84.381 ;
      RECT 0.355 -85.075 0.495 -84.905 ;
      RECT 0.355 -83.579 0.445 -82.572 ;
      RECT 0.355 -83.055 0.495 -82.885 ;
      RECT 0.355 -82.158 0.445 -81.151 ;
      RECT 0.355 -81.845 0.495 -81.675 ;
      RECT 0.355 -80.349 0.445 -79.342 ;
      RECT 0.355 -79.825 0.495 -79.655 ;
      RECT 0.355 -78.928 0.445 -77.921 ;
      RECT 0.355 -78.615 0.495 -78.445 ;
      RECT 0.355 -77.119 0.445 -76.112 ;
      RECT 0.355 -76.595 0.495 -76.425 ;
      RECT 0.355 -75.698 0.445 -74.691 ;
      RECT 0.355 -75.385 0.495 -75.215 ;
      RECT 0.355 -73.889 0.445 -72.882 ;
      RECT 0.355 -73.365 0.495 -73.195 ;
      RECT 0.355 -72.468 0.445 -71.461 ;
      RECT 0.355 -72.155 0.495 -71.985 ;
      RECT 0.355 -70.659 0.445 -69.652 ;
      RECT 0.355 -70.135 0.495 -69.965 ;
      RECT 0.355 -69.238 0.445 -68.231 ;
      RECT 0.355 -68.925 0.495 -68.755 ;
      RECT 0.355 -67.429 0.445 -66.422 ;
      RECT 0.355 -66.905 0.495 -66.735 ;
      RECT 0.355 -66.008 0.445 -65.001 ;
      RECT 0.355 -65.695 0.495 -65.525 ;
      RECT 0.355 -64.199 0.445 -63.192 ;
      RECT 0.355 -63.675 0.495 -63.505 ;
      RECT 0.355 -62.778 0.445 -61.771 ;
      RECT 0.355 -62.465 0.495 -62.295 ;
      RECT 0.355 -60.969 0.445 -59.962 ;
      RECT 0.355 -60.445 0.495 -60.275 ;
      RECT 0.355 -59.548 0.445 -58.541 ;
      RECT 0.355 -59.235 0.495 -59.065 ;
      RECT 0.355 -57.739 0.445 -56.732 ;
      RECT 0.355 -57.215 0.495 -57.045 ;
      RECT 0.355 -56.318 0.445 -55.311 ;
      RECT 0.355 -56.005 0.495 -55.835 ;
      RECT 0.355 -54.509 0.445 -53.502 ;
      RECT 0.355 -53.985 0.495 -53.815 ;
      RECT 0.355 -53.088 0.445 -52.081 ;
      RECT 0.355 -52.775 0.495 -52.605 ;
      RECT 0.355 -51.279 0.445 -50.272 ;
      RECT 0.355 -50.755 0.495 -50.585 ;
      RECT 0.355 -49.858 0.445 -48.851 ;
      RECT 0.355 -49.545 0.495 -49.375 ;
      RECT 0.355 -48.049 0.445 -47.042 ;
      RECT 0.355 -47.525 0.495 -47.355 ;
      RECT 0.355 -46.628 0.445 -45.621 ;
      RECT 0.355 -46.315 0.495 -46.145 ;
      RECT 0.355 -44.819 0.445 -43.812 ;
      RECT 0.355 -44.295 0.495 -44.125 ;
      RECT 0.355 -43.398 0.445 -42.391 ;
      RECT 0.355 -43.085 0.495 -42.915 ;
      RECT 0.355 -41.589 0.445 -40.582 ;
      RECT 0.355 -41.065 0.495 -40.895 ;
      RECT 0.355 -40.168 0.445 -39.161 ;
      RECT 0.355 -39.855 0.495 -39.685 ;
      RECT 0.355 -38.359 0.445 -37.352 ;
      RECT 0.355 -37.835 0.495 -37.665 ;
      RECT 0.355 -36.938 0.445 -35.931 ;
      RECT 0.355 -36.625 0.495 -36.455 ;
      RECT 0.355 -35.129 0.445 -34.122 ;
      RECT 0.355 -34.605 0.495 -34.435 ;
      RECT 0.355 -33.708 0.445 -32.701 ;
      RECT 0.355 -33.395 0.495 -33.225 ;
      RECT 0.355 -31.899 0.445 -30.892 ;
      RECT 0.355 -31.375 0.495 -31.205 ;
      RECT 0.355 -30.478 0.445 -29.471 ;
      RECT 0.355 -30.165 0.495 -29.995 ;
      RECT 0.355 -28.669 0.445 -27.662 ;
      RECT 0.355 -28.145 0.495 -27.975 ;
      RECT 0.355 -27.248 0.445 -26.241 ;
      RECT 0.355 -26.935 0.495 -26.765 ;
      RECT 0.355 -25.439 0.445 -24.432 ;
      RECT 0.355 -24.915 0.495 -24.745 ;
      RECT 0.355 -24.018 0.445 -23.011 ;
      RECT 0.355 -23.705 0.495 -23.535 ;
      RECT 0.355 -22.209 0.445 -21.202 ;
      RECT 0.355 -21.685 0.495 -21.515 ;
      RECT 0.355 -20.788 0.445 -19.781 ;
      RECT 0.355 -20.475 0.495 -20.305 ;
      RECT 0.355 -18.979 0.445 -17.972 ;
      RECT 0.355 -18.455 0.495 -18.285 ;
      RECT 0.355 -17.558 0.445 -16.551 ;
      RECT 0.355 -17.245 0.495 -17.075 ;
      RECT 0.355 -15.749 0.445 -14.742 ;
      RECT 0.355 -15.225 0.495 -15.055 ;
      RECT 0.355 -14.328 0.445 -13.321 ;
      RECT 0.355 -14.015 0.495 -13.845 ;
      RECT 0.355 -12.519 0.445 -11.512 ;
      RECT 0.355 -11.995 0.495 -11.825 ;
      RECT 0.355 -11.098 0.445 -10.091 ;
      RECT 0.355 -10.785 0.495 -10.615 ;
      RECT 0.355 -9.289 0.445 -8.282 ;
      RECT 0.355 -8.765 0.495 -8.595 ;
      RECT 0.355 -7.868 0.445 -6.861 ;
      RECT 0.355 -7.555 0.495 -7.385 ;
      RECT 0.355 -6.059 0.445 -5.052 ;
      RECT 0.355 -5.535 0.495 -5.365 ;
      RECT 0.355 -4.638 0.445 -3.631 ;
      RECT 0.355 -4.325 0.495 -4.155 ;
      RECT 0.355 -2.829 0.445 -1.822 ;
      RECT 0.355 -2.305 0.495 -2.135 ;
      RECT 0.355 -1.408 0.445 -0.401 ;
      RECT 0.355 -1.095 0.495 -0.925 ;
      RECT 0.355 0.401 0.445 1.408 ;
      RECT 0.355 0.925 0.495 1.095 ;
      RECT -5.785 4.135 -5.615 4.76 ;
      RECT -6.345 4.135 -6.245 4.76 ;
      RECT -6.345 4.135 -0.425 4.235 ;
      RECT -1.985 -108.545 -1.885 -107.055 ;
      RECT -3.285 -108.545 -3.185 -107.055 ;
      RECT -4.585 -108.545 -4.485 -107.055 ;
      RECT -5.885 -108.545 -5.785 -107.055 ;
      RECT -7.185 -108.545 -7.085 -107.055 ;
      RECT -8.485 -108.545 -8.385 -107.055 ;
      RECT -9.785 -108.545 -9.685 -107.055 ;
      RECT -11.085 -108.545 -10.985 -107.055 ;
      RECT -1.205 -108.545 -1.105 -107.235 ;
      RECT -2.505 -108.545 -2.405 -107.235 ;
      RECT -3.805 -108.545 -3.705 -107.235 ;
      RECT -5.105 -108.545 -5.005 -107.235 ;
      RECT -6.405 -108.545 -6.305 -107.235 ;
      RECT -7.705 -108.545 -7.605 -107.235 ;
      RECT -9.005 -108.545 -8.905 -107.235 ;
      RECT -10.305 -108.545 -10.205 -107.235 ;
      RECT -39.505 -108.545 -0.765 -107.865 ;
      RECT -11.705 -109.175 -11.605 -107.865 ;
      RECT -12.305 -109.175 -12.205 -107.865 ;
      RECT -1.205 -102.895 -1.105 -100.595 ;
      RECT -1.725 -102.895 -1.625 -100.595 ;
      RECT -2.505 -102.895 -2.405 -100.595 ;
      RECT -3.025 -102.895 -2.925 -100.595 ;
      RECT -3.805 -102.895 -3.705 -100.595 ;
      RECT -4.325 -102.895 -4.225 -100.595 ;
      RECT -5.105 -102.895 -5.005 -100.595 ;
      RECT -5.625 -102.895 -5.525 -100.595 ;
      RECT -6.405 -102.895 -6.305 -100.595 ;
      RECT -6.925 -102.895 -6.825 -100.595 ;
      RECT -7.705 -102.895 -7.605 -100.595 ;
      RECT -8.225 -102.895 -8.125 -100.595 ;
      RECT -9.005 -102.895 -8.905 -100.595 ;
      RECT -9.525 -102.895 -9.425 -100.595 ;
      RECT -10.305 -102.895 -10.205 -100.595 ;
      RECT -10.825 -102.895 -10.725 -100.595 ;
      RECT -11.605 -102.085 -11.505 -100.595 ;
      RECT -12.125 -102.085 -12.025 -100.595 ;
      RECT -12.905 -102.085 -12.805 -100.595 ;
      RECT -13.425 -102.085 -13.325 -100.595 ;
      RECT -14.205 -102.085 -14.105 -100.595 ;
      RECT -14.725 -102.085 -14.625 -100.595 ;
      RECT -15.505 -102.085 -15.405 -100.595 ;
      RECT -16.025 -102.085 -15.925 -100.595 ;
      RECT -16.805 -102.085 -16.705 -100.595 ;
      RECT -17.325 -102.085 -17.225 -100.595 ;
      RECT -18.105 -102.085 -18.005 -100.595 ;
      RECT -18.625 -102.085 -18.525 -100.595 ;
      RECT -19.405 -102.085 -19.305 -100.595 ;
      RECT -19.925 -102.085 -19.825 -100.595 ;
      RECT -20.705 -102.085 -20.605 -100.595 ;
      RECT -21.225 -102.085 -21.125 -100.595 ;
      RECT -22.005 -102.085 -21.905 -100.595 ;
      RECT -22.525 -102.085 -22.425 -100.595 ;
      RECT -23.305 -102.085 -23.205 -100.595 ;
      RECT -23.825 -102.085 -23.725 -100.595 ;
      RECT -24.605 -102.085 -24.505 -100.595 ;
      RECT -25.125 -102.085 -25.025 -100.595 ;
      RECT -25.905 -102.085 -25.805 -100.595 ;
      RECT -26.425 -102.085 -26.325 -100.595 ;
      RECT -27.205 -102.085 -27.105 -100.595 ;
      RECT -27.725 -102.085 -27.625 -100.595 ;
      RECT -28.505 -102.085 -28.405 -100.595 ;
      RECT -29.025 -102.085 -28.925 -100.595 ;
      RECT -29.805 -102.085 -29.705 -100.595 ;
      RECT -30.325 -102.085 -30.225 -100.595 ;
      RECT -31.105 -102.085 -31.005 -100.595 ;
      RECT -31.625 -102.085 -31.525 -100.595 ;
      RECT -37.505 -102.085 -0.765 -101.405 ;
      RECT -1.985 -96.435 -1.885 -94.135 ;
      RECT -3.285 -96.435 -3.185 -94.135 ;
      RECT -4.585 -96.435 -4.485 -94.135 ;
      RECT -5.885 -96.435 -5.785 -94.135 ;
      RECT -7.185 -96.435 -7.085 -94.135 ;
      RECT -8.485 -96.435 -8.385 -94.135 ;
      RECT -9.785 -96.435 -9.685 -94.135 ;
      RECT -11.085 -96.435 -10.985 -94.135 ;
      RECT -12.385 -96.435 -12.285 -94.135 ;
      RECT -13.685 -96.435 -13.585 -94.135 ;
      RECT -14.985 -96.435 -14.885 -94.135 ;
      RECT -16.285 -96.435 -16.185 -94.135 ;
      RECT -17.585 -96.435 -17.485 -94.135 ;
      RECT -18.885 -96.435 -18.785 -94.135 ;
      RECT -20.185 -96.435 -20.085 -94.135 ;
      RECT -21.485 -96.435 -21.385 -94.135 ;
      RECT -22.785 -96.435 -22.685 -94.135 ;
      RECT -24.085 -96.435 -23.985 -94.135 ;
      RECT -25.385 -96.435 -25.285 -94.135 ;
      RECT -26.685 -96.435 -26.585 -94.135 ;
      RECT -27.985 -96.435 -27.885 -94.135 ;
      RECT -29.285 -96.435 -29.185 -94.135 ;
      RECT -30.585 -96.435 -30.485 -94.135 ;
      RECT -31.885 -96.435 -31.785 -94.135 ;
      RECT -1.205 -96.255 -1.105 -94.315 ;
      RECT -2.505 -96.255 -2.405 -94.315 ;
      RECT -3.805 -96.255 -3.705 -94.315 ;
      RECT -5.105 -96.255 -5.005 -94.315 ;
      RECT -6.405 -96.255 -6.305 -94.315 ;
      RECT -7.705 -96.255 -7.605 -94.315 ;
      RECT -9.005 -96.255 -8.905 -94.315 ;
      RECT -10.305 -96.255 -10.205 -94.315 ;
      RECT -11.605 -96.255 -11.505 -94.315 ;
      RECT -12.905 -96.255 -12.805 -94.315 ;
      RECT -14.205 -96.255 -14.105 -94.315 ;
      RECT -15.505 -96.255 -15.405 -94.315 ;
      RECT -16.805 -96.255 -16.705 -94.315 ;
      RECT -18.105 -96.255 -18.005 -94.315 ;
      RECT -19.405 -96.255 -19.305 -94.315 ;
      RECT -20.705 -96.255 -20.605 -94.315 ;
      RECT -22.005 -96.255 -21.905 -94.315 ;
      RECT -23.305 -96.255 -23.205 -94.315 ;
      RECT -24.605 -96.255 -24.505 -94.315 ;
      RECT -25.905 -96.255 -25.805 -94.315 ;
      RECT -27.205 -96.255 -27.105 -94.315 ;
      RECT -28.505 -96.255 -28.405 -94.315 ;
      RECT -29.805 -96.255 -29.705 -94.315 ;
      RECT -31.105 -96.255 -31.005 -94.315 ;
      RECT -39.505 -95.625 -0.765 -94.945 ;
      RECT -1.205 -89.975 -1.105 -87.675 ;
      RECT -1.725 -89.975 -1.625 -87.675 ;
      RECT -2.505 -89.975 -2.405 -87.675 ;
      RECT -3.025 -89.975 -2.925 -87.675 ;
      RECT -3.805 -89.975 -3.705 -87.675 ;
      RECT -4.325 -89.975 -4.225 -87.675 ;
      RECT -5.105 -89.975 -5.005 -87.675 ;
      RECT -5.625 -89.975 -5.525 -87.675 ;
      RECT -6.405 -89.975 -6.305 -87.675 ;
      RECT -6.925 -89.975 -6.825 -87.675 ;
      RECT -7.705 -89.975 -7.605 -87.675 ;
      RECT -8.225 -89.975 -8.125 -87.675 ;
      RECT -9.005 -89.975 -8.905 -87.675 ;
      RECT -9.525 -89.975 -9.425 -87.675 ;
      RECT -10.305 -89.975 -10.205 -87.675 ;
      RECT -10.825 -89.975 -10.725 -87.675 ;
      RECT -11.605 -89.975 -11.505 -87.675 ;
      RECT -12.125 -89.975 -12.025 -87.675 ;
      RECT -12.905 -89.975 -12.805 -87.675 ;
      RECT -13.425 -89.975 -13.325 -87.675 ;
      RECT -14.205 -89.975 -14.105 -87.675 ;
      RECT -14.725 -89.975 -14.625 -87.675 ;
      RECT -15.505 -89.975 -15.405 -87.675 ;
      RECT -16.025 -89.975 -15.925 -87.675 ;
      RECT -16.805 -89.975 -16.705 -87.675 ;
      RECT -17.325 -89.975 -17.225 -87.675 ;
      RECT -18.105 -89.975 -18.005 -87.675 ;
      RECT -18.625 -89.975 -18.525 -87.675 ;
      RECT -19.405 -89.975 -19.305 -87.675 ;
      RECT -19.925 -89.975 -19.825 -87.675 ;
      RECT -20.705 -89.975 -20.605 -87.675 ;
      RECT -21.225 -89.975 -21.125 -87.675 ;
      RECT -22.005 -89.975 -21.905 -87.675 ;
      RECT -22.525 -89.975 -22.425 -87.675 ;
      RECT -23.305 -89.975 -23.205 -87.675 ;
      RECT -23.825 -89.975 -23.725 -87.675 ;
      RECT -24.605 -89.975 -24.505 -87.675 ;
      RECT -25.125 -89.975 -25.025 -87.675 ;
      RECT -25.905 -89.975 -25.805 -87.675 ;
      RECT -26.425 -89.975 -26.325 -87.675 ;
      RECT -27.205 -89.975 -27.105 -87.675 ;
      RECT -27.725 -89.975 -27.625 -87.675 ;
      RECT -28.505 -89.975 -28.405 -87.675 ;
      RECT -29.025 -89.975 -28.925 -87.675 ;
      RECT -29.805 -89.975 -29.705 -87.675 ;
      RECT -30.325 -89.975 -30.225 -87.675 ;
      RECT -31.105 -89.975 -31.005 -87.675 ;
      RECT -31.625 -89.975 -31.525 -87.675 ;
      RECT -37.505 -89.165 -0.765 -88.485 ;
      RECT -1.985 -83.515 -1.885 -81.215 ;
      RECT -3.285 -83.515 -3.185 -81.215 ;
      RECT -4.585 -83.515 -4.485 -81.215 ;
      RECT -5.885 -83.515 -5.785 -81.215 ;
      RECT -7.185 -83.515 -7.085 -81.215 ;
      RECT -8.485 -83.515 -8.385 -81.215 ;
      RECT -9.785 -83.515 -9.685 -81.215 ;
      RECT -11.085 -83.515 -10.985 -81.215 ;
      RECT -12.385 -83.515 -12.285 -81.215 ;
      RECT -13.685 -83.515 -13.585 -81.215 ;
      RECT -14.985 -83.515 -14.885 -81.215 ;
      RECT -16.285 -83.515 -16.185 -81.215 ;
      RECT -17.585 -83.515 -17.485 -81.215 ;
      RECT -18.885 -83.515 -18.785 -81.215 ;
      RECT -20.185 -83.515 -20.085 -81.215 ;
      RECT -21.485 -83.515 -21.385 -81.215 ;
      RECT -22.785 -83.515 -22.685 -81.215 ;
      RECT -24.085 -83.515 -23.985 -81.215 ;
      RECT -25.385 -83.515 -25.285 -81.215 ;
      RECT -26.685 -83.515 -26.585 -81.215 ;
      RECT -27.985 -83.515 -27.885 -81.215 ;
      RECT -29.285 -83.515 -29.185 -81.215 ;
      RECT -30.585 -83.515 -30.485 -81.215 ;
      RECT -31.885 -83.515 -31.785 -81.215 ;
      RECT -1.205 -83.335 -1.105 -81.395 ;
      RECT -2.505 -83.335 -2.405 -81.395 ;
      RECT -3.805 -83.335 -3.705 -81.395 ;
      RECT -5.105 -83.335 -5.005 -81.395 ;
      RECT -6.405 -83.335 -6.305 -81.395 ;
      RECT -7.705 -83.335 -7.605 -81.395 ;
      RECT -9.005 -83.335 -8.905 -81.395 ;
      RECT -10.305 -83.335 -10.205 -81.395 ;
      RECT -11.605 -83.335 -11.505 -81.395 ;
      RECT -12.905 -83.335 -12.805 -81.395 ;
      RECT -14.205 -83.335 -14.105 -81.395 ;
      RECT -15.505 -83.335 -15.405 -81.395 ;
      RECT -16.805 -83.335 -16.705 -81.395 ;
      RECT -18.105 -83.335 -18.005 -81.395 ;
      RECT -19.405 -83.335 -19.305 -81.395 ;
      RECT -20.705 -83.335 -20.605 -81.395 ;
      RECT -22.005 -83.335 -21.905 -81.395 ;
      RECT -23.305 -83.335 -23.205 -81.395 ;
      RECT -24.605 -83.335 -24.505 -81.395 ;
      RECT -25.905 -83.335 -25.805 -81.395 ;
      RECT -27.205 -83.335 -27.105 -81.395 ;
      RECT -28.505 -83.335 -28.405 -81.395 ;
      RECT -29.805 -83.335 -29.705 -81.395 ;
      RECT -31.105 -83.335 -31.005 -81.395 ;
      RECT -39.505 -82.705 -0.765 -82.025 ;
      RECT -1.205 -77.055 -1.105 -74.755 ;
      RECT -1.725 -77.055 -1.625 -74.755 ;
      RECT -2.505 -77.055 -2.405 -74.755 ;
      RECT -3.025 -77.055 -2.925 -74.755 ;
      RECT -3.805 -77.055 -3.705 -74.755 ;
      RECT -4.325 -77.055 -4.225 -74.755 ;
      RECT -5.105 -77.055 -5.005 -74.755 ;
      RECT -5.625 -77.055 -5.525 -74.755 ;
      RECT -6.405 -77.055 -6.305 -74.755 ;
      RECT -6.925 -77.055 -6.825 -74.755 ;
      RECT -7.705 -77.055 -7.605 -74.755 ;
      RECT -8.225 -77.055 -8.125 -74.755 ;
      RECT -9.005 -77.055 -8.905 -74.755 ;
      RECT -9.525 -77.055 -9.425 -74.755 ;
      RECT -10.305 -77.055 -10.205 -74.755 ;
      RECT -10.825 -77.055 -10.725 -74.755 ;
      RECT -11.605 -77.055 -11.505 -74.755 ;
      RECT -12.125 -77.055 -12.025 -74.755 ;
      RECT -12.905 -77.055 -12.805 -74.755 ;
      RECT -13.425 -77.055 -13.325 -74.755 ;
      RECT -14.205 -77.055 -14.105 -74.755 ;
      RECT -14.725 -77.055 -14.625 -74.755 ;
      RECT -15.505 -77.055 -15.405 -74.755 ;
      RECT -16.025 -77.055 -15.925 -74.755 ;
      RECT -16.805 -77.055 -16.705 -74.755 ;
      RECT -17.325 -77.055 -17.225 -74.755 ;
      RECT -18.105 -77.055 -18.005 -74.755 ;
      RECT -18.625 -77.055 -18.525 -74.755 ;
      RECT -19.405 -77.055 -19.305 -74.755 ;
      RECT -19.925 -77.055 -19.825 -74.755 ;
      RECT -20.705 -77.055 -20.605 -74.755 ;
      RECT -21.225 -77.055 -21.125 -74.755 ;
      RECT -22.005 -77.055 -21.905 -74.755 ;
      RECT -22.525 -77.055 -22.425 -74.755 ;
      RECT -23.305 -77.055 -23.205 -74.755 ;
      RECT -23.825 -77.055 -23.725 -74.755 ;
      RECT -24.605 -77.055 -24.505 -74.755 ;
      RECT -25.125 -77.055 -25.025 -74.755 ;
      RECT -25.905 -77.055 -25.805 -74.755 ;
      RECT -26.425 -77.055 -26.325 -74.755 ;
      RECT -27.205 -77.055 -27.105 -74.755 ;
      RECT -27.725 -77.055 -27.625 -74.755 ;
      RECT -28.505 -77.055 -28.405 -74.755 ;
      RECT -29.025 -77.055 -28.925 -74.755 ;
      RECT -29.805 -77.055 -29.705 -74.755 ;
      RECT -30.325 -77.055 -30.225 -74.755 ;
      RECT -31.105 -77.055 -31.005 -74.755 ;
      RECT -31.625 -77.055 -31.525 -74.755 ;
      RECT -37.505 -76.245 -0.765 -75.565 ;
      RECT -1.985 -70.595 -1.885 -68.295 ;
      RECT -3.285 -70.595 -3.185 -68.295 ;
      RECT -4.585 -70.595 -4.485 -68.295 ;
      RECT -5.885 -70.595 -5.785 -68.295 ;
      RECT -7.185 -70.595 -7.085 -68.295 ;
      RECT -8.485 -70.595 -8.385 -68.295 ;
      RECT -9.785 -70.595 -9.685 -68.295 ;
      RECT -11.085 -70.595 -10.985 -68.295 ;
      RECT -12.385 -70.595 -12.285 -68.295 ;
      RECT -13.685 -70.595 -13.585 -68.295 ;
      RECT -14.985 -70.595 -14.885 -68.295 ;
      RECT -16.285 -70.595 -16.185 -68.295 ;
      RECT -17.585 -70.595 -17.485 -68.295 ;
      RECT -18.885 -70.595 -18.785 -68.295 ;
      RECT -20.185 -70.595 -20.085 -68.295 ;
      RECT -21.485 -70.595 -21.385 -68.295 ;
      RECT -22.785 -70.595 -22.685 -68.295 ;
      RECT -24.085 -70.595 -23.985 -68.295 ;
      RECT -25.385 -70.595 -25.285 -68.295 ;
      RECT -26.685 -70.595 -26.585 -68.295 ;
      RECT -27.985 -70.595 -27.885 -68.295 ;
      RECT -29.285 -70.595 -29.185 -68.295 ;
      RECT -30.585 -70.595 -30.485 -68.295 ;
      RECT -31.885 -70.595 -31.785 -68.295 ;
      RECT -1.205 -70.415 -1.105 -68.475 ;
      RECT -2.505 -70.415 -2.405 -68.475 ;
      RECT -3.805 -70.415 -3.705 -68.475 ;
      RECT -5.105 -70.415 -5.005 -68.475 ;
      RECT -6.405 -70.415 -6.305 -68.475 ;
      RECT -7.705 -70.415 -7.605 -68.475 ;
      RECT -9.005 -70.415 -8.905 -68.475 ;
      RECT -10.305 -70.415 -10.205 -68.475 ;
      RECT -11.605 -70.415 -11.505 -68.475 ;
      RECT -12.905 -70.415 -12.805 -68.475 ;
      RECT -14.205 -70.415 -14.105 -68.475 ;
      RECT -15.505 -70.415 -15.405 -68.475 ;
      RECT -16.805 -70.415 -16.705 -68.475 ;
      RECT -18.105 -70.415 -18.005 -68.475 ;
      RECT -19.405 -70.415 -19.305 -68.475 ;
      RECT -20.705 -70.415 -20.605 -68.475 ;
      RECT -22.005 -70.415 -21.905 -68.475 ;
      RECT -23.305 -70.415 -23.205 -68.475 ;
      RECT -24.605 -70.415 -24.505 -68.475 ;
      RECT -25.905 -70.415 -25.805 -68.475 ;
      RECT -27.205 -70.415 -27.105 -68.475 ;
      RECT -28.505 -70.415 -28.405 -68.475 ;
      RECT -29.805 -70.415 -29.705 -68.475 ;
      RECT -31.105 -70.415 -31.005 -68.475 ;
      RECT -39.505 -69.785 -0.765 -69.105 ;
      RECT -1.205 -64.135 -1.105 -61.835 ;
      RECT -1.725 -64.135 -1.625 -61.835 ;
      RECT -2.505 -64.135 -2.405 -61.835 ;
      RECT -3.025 -64.135 -2.925 -61.835 ;
      RECT -3.805 -64.135 -3.705 -61.835 ;
      RECT -4.325 -64.135 -4.225 -61.835 ;
      RECT -5.105 -64.135 -5.005 -61.835 ;
      RECT -5.625 -64.135 -5.525 -61.835 ;
      RECT -6.405 -64.135 -6.305 -61.835 ;
      RECT -6.925 -64.135 -6.825 -61.835 ;
      RECT -7.705 -64.135 -7.605 -61.835 ;
      RECT -8.225 -64.135 -8.125 -61.835 ;
      RECT -9.005 -64.135 -8.905 -61.835 ;
      RECT -9.525 -64.135 -9.425 -61.835 ;
      RECT -10.305 -64.135 -10.205 -61.835 ;
      RECT -10.825 -64.135 -10.725 -61.835 ;
      RECT -11.605 -64.135 -11.505 -61.835 ;
      RECT -12.125 -64.135 -12.025 -61.835 ;
      RECT -12.905 -64.135 -12.805 -61.835 ;
      RECT -13.425 -64.135 -13.325 -61.835 ;
      RECT -14.205 -64.135 -14.105 -61.835 ;
      RECT -14.725 -64.135 -14.625 -61.835 ;
      RECT -15.505 -64.135 -15.405 -61.835 ;
      RECT -16.025 -64.135 -15.925 -61.835 ;
      RECT -16.805 -64.135 -16.705 -61.835 ;
      RECT -17.325 -64.135 -17.225 -61.835 ;
      RECT -18.105 -64.135 -18.005 -61.835 ;
      RECT -18.625 -64.135 -18.525 -61.835 ;
      RECT -19.405 -64.135 -19.305 -61.835 ;
      RECT -19.925 -64.135 -19.825 -61.835 ;
      RECT -20.705 -64.135 -20.605 -61.835 ;
      RECT -21.225 -64.135 -21.125 -61.835 ;
      RECT -22.005 -64.135 -21.905 -61.835 ;
      RECT -22.525 -64.135 -22.425 -61.835 ;
      RECT -23.305 -64.135 -23.205 -61.835 ;
      RECT -23.825 -64.135 -23.725 -61.835 ;
      RECT -24.605 -64.135 -24.505 -61.835 ;
      RECT -25.125 -64.135 -25.025 -61.835 ;
      RECT -25.905 -64.135 -25.805 -61.835 ;
      RECT -26.425 -64.135 -26.325 -61.835 ;
      RECT -27.205 -64.135 -27.105 -61.835 ;
      RECT -27.725 -64.135 -27.625 -61.835 ;
      RECT -28.505 -64.135 -28.405 -61.835 ;
      RECT -29.025 -64.135 -28.925 -61.835 ;
      RECT -29.805 -64.135 -29.705 -61.835 ;
      RECT -30.325 -64.135 -30.225 -61.835 ;
      RECT -31.105 -64.135 -31.005 -61.835 ;
      RECT -31.625 -64.135 -31.525 -61.835 ;
      RECT -37.505 -63.325 -0.765 -62.645 ;
      RECT -1.985 -57.675 -1.885 -55.375 ;
      RECT -3.285 -57.675 -3.185 -55.375 ;
      RECT -4.585 -57.675 -4.485 -55.375 ;
      RECT -5.885 -57.675 -5.785 -55.375 ;
      RECT -7.185 -57.675 -7.085 -55.375 ;
      RECT -8.485 -57.675 -8.385 -55.375 ;
      RECT -9.785 -57.675 -9.685 -55.375 ;
      RECT -11.085 -57.675 -10.985 -55.375 ;
      RECT -12.385 -57.675 -12.285 -55.375 ;
      RECT -13.685 -57.675 -13.585 -55.375 ;
      RECT -14.985 -57.675 -14.885 -55.375 ;
      RECT -16.285 -57.675 -16.185 -55.375 ;
      RECT -17.585 -57.675 -17.485 -55.375 ;
      RECT -18.885 -57.675 -18.785 -55.375 ;
      RECT -20.185 -57.675 -20.085 -55.375 ;
      RECT -21.485 -57.675 -21.385 -55.375 ;
      RECT -22.785 -57.675 -22.685 -55.375 ;
      RECT -24.085 -57.675 -23.985 -55.375 ;
      RECT -25.385 -57.675 -25.285 -55.375 ;
      RECT -26.685 -57.675 -26.585 -55.375 ;
      RECT -27.985 -57.675 -27.885 -55.375 ;
      RECT -29.285 -57.675 -29.185 -55.375 ;
      RECT -30.585 -57.675 -30.485 -55.375 ;
      RECT -31.885 -57.675 -31.785 -55.375 ;
      RECT -1.205 -57.495 -1.105 -55.555 ;
      RECT -2.505 -57.495 -2.405 -55.555 ;
      RECT -3.805 -57.495 -3.705 -55.555 ;
      RECT -5.105 -57.495 -5.005 -55.555 ;
      RECT -6.405 -57.495 -6.305 -55.555 ;
      RECT -7.705 -57.495 -7.605 -55.555 ;
      RECT -9.005 -57.495 -8.905 -55.555 ;
      RECT -10.305 -57.495 -10.205 -55.555 ;
      RECT -11.605 -57.495 -11.505 -55.555 ;
      RECT -12.905 -57.495 -12.805 -55.555 ;
      RECT -14.205 -57.495 -14.105 -55.555 ;
      RECT -15.505 -57.495 -15.405 -55.555 ;
      RECT -16.805 -57.495 -16.705 -55.555 ;
      RECT -18.105 -57.495 -18.005 -55.555 ;
      RECT -19.405 -57.495 -19.305 -55.555 ;
      RECT -20.705 -57.495 -20.605 -55.555 ;
      RECT -22.005 -57.495 -21.905 -55.555 ;
      RECT -23.305 -57.495 -23.205 -55.555 ;
      RECT -24.605 -57.495 -24.505 -55.555 ;
      RECT -25.905 -57.495 -25.805 -55.555 ;
      RECT -27.205 -57.495 -27.105 -55.555 ;
      RECT -28.505 -57.495 -28.405 -55.555 ;
      RECT -29.805 -57.495 -29.705 -55.555 ;
      RECT -31.105 -57.495 -31.005 -55.555 ;
      RECT -39.505 -56.865 -0.765 -56.185 ;
      RECT -1.205 -51.215 -1.105 -48.915 ;
      RECT -1.725 -51.215 -1.625 -48.915 ;
      RECT -2.505 -51.215 -2.405 -48.915 ;
      RECT -3.025 -51.215 -2.925 -48.915 ;
      RECT -3.805 -51.215 -3.705 -48.915 ;
      RECT -4.325 -51.215 -4.225 -48.915 ;
      RECT -5.105 -51.215 -5.005 -48.915 ;
      RECT -5.625 -51.215 -5.525 -48.915 ;
      RECT -6.405 -51.215 -6.305 -48.915 ;
      RECT -6.925 -51.215 -6.825 -48.915 ;
      RECT -7.705 -51.215 -7.605 -48.915 ;
      RECT -8.225 -51.215 -8.125 -48.915 ;
      RECT -9.005 -51.215 -8.905 -48.915 ;
      RECT -9.525 -51.215 -9.425 -48.915 ;
      RECT -10.305 -51.215 -10.205 -48.915 ;
      RECT -10.825 -51.215 -10.725 -48.915 ;
      RECT -11.605 -51.215 -11.505 -48.915 ;
      RECT -12.125 -51.215 -12.025 -48.915 ;
      RECT -12.905 -51.215 -12.805 -48.915 ;
      RECT -13.425 -51.215 -13.325 -48.915 ;
      RECT -14.205 -51.215 -14.105 -48.915 ;
      RECT -14.725 -51.215 -14.625 -48.915 ;
      RECT -15.505 -51.215 -15.405 -48.915 ;
      RECT -16.025 -51.215 -15.925 -48.915 ;
      RECT -16.805 -51.215 -16.705 -48.915 ;
      RECT -17.325 -51.215 -17.225 -48.915 ;
      RECT -18.105 -51.215 -18.005 -48.915 ;
      RECT -18.625 -51.215 -18.525 -48.915 ;
      RECT -19.405 -51.215 -19.305 -48.915 ;
      RECT -19.925 -51.215 -19.825 -48.915 ;
      RECT -20.705 -51.215 -20.605 -48.915 ;
      RECT -21.225 -51.215 -21.125 -48.915 ;
      RECT -22.005 -51.215 -21.905 -48.915 ;
      RECT -22.525 -51.215 -22.425 -48.915 ;
      RECT -23.305 -51.215 -23.205 -48.915 ;
      RECT -23.825 -51.215 -23.725 -48.915 ;
      RECT -24.605 -51.215 -24.505 -48.915 ;
      RECT -25.125 -51.215 -25.025 -48.915 ;
      RECT -25.905 -51.215 -25.805 -48.915 ;
      RECT -26.425 -51.215 -26.325 -48.915 ;
      RECT -27.205 -51.215 -27.105 -48.915 ;
      RECT -27.725 -51.215 -27.625 -48.915 ;
      RECT -28.505 -51.215 -28.405 -48.915 ;
      RECT -29.025 -51.215 -28.925 -48.915 ;
      RECT -29.805 -51.215 -29.705 -48.915 ;
      RECT -30.325 -51.215 -30.225 -48.915 ;
      RECT -31.105 -51.215 -31.005 -48.915 ;
      RECT -31.625 -51.215 -31.525 -48.915 ;
      RECT -37.505 -50.405 -0.765 -49.725 ;
      RECT -1.985 -44.755 -1.885 -42.455 ;
      RECT -3.285 -44.755 -3.185 -42.455 ;
      RECT -4.585 -44.755 -4.485 -42.455 ;
      RECT -5.885 -44.755 -5.785 -42.455 ;
      RECT -7.185 -44.755 -7.085 -42.455 ;
      RECT -8.485 -44.755 -8.385 -42.455 ;
      RECT -9.785 -44.755 -9.685 -42.455 ;
      RECT -11.085 -44.755 -10.985 -42.455 ;
      RECT -12.385 -44.755 -12.285 -42.455 ;
      RECT -13.685 -44.755 -13.585 -42.455 ;
      RECT -14.985 -44.755 -14.885 -42.455 ;
      RECT -16.285 -44.755 -16.185 -42.455 ;
      RECT -17.585 -44.755 -17.485 -42.455 ;
      RECT -18.885 -44.755 -18.785 -42.455 ;
      RECT -20.185 -44.755 -20.085 -42.455 ;
      RECT -21.485 -44.755 -21.385 -42.455 ;
      RECT -22.785 -44.755 -22.685 -42.455 ;
      RECT -24.085 -44.755 -23.985 -42.455 ;
      RECT -25.385 -44.755 -25.285 -42.455 ;
      RECT -26.685 -44.755 -26.585 -42.455 ;
      RECT -27.985 -44.755 -27.885 -42.455 ;
      RECT -29.285 -44.755 -29.185 -42.455 ;
      RECT -30.585 -44.755 -30.485 -42.455 ;
      RECT -31.885 -44.755 -31.785 -42.455 ;
      RECT -1.205 -44.575 -1.105 -42.635 ;
      RECT -2.505 -44.575 -2.405 -42.635 ;
      RECT -3.805 -44.575 -3.705 -42.635 ;
      RECT -5.105 -44.575 -5.005 -42.635 ;
      RECT -6.405 -44.575 -6.305 -42.635 ;
      RECT -7.705 -44.575 -7.605 -42.635 ;
      RECT -9.005 -44.575 -8.905 -42.635 ;
      RECT -10.305 -44.575 -10.205 -42.635 ;
      RECT -11.605 -44.575 -11.505 -42.635 ;
      RECT -12.905 -44.575 -12.805 -42.635 ;
      RECT -14.205 -44.575 -14.105 -42.635 ;
      RECT -15.505 -44.575 -15.405 -42.635 ;
      RECT -16.805 -44.575 -16.705 -42.635 ;
      RECT -18.105 -44.575 -18.005 -42.635 ;
      RECT -19.405 -44.575 -19.305 -42.635 ;
      RECT -20.705 -44.575 -20.605 -42.635 ;
      RECT -22.005 -44.575 -21.905 -42.635 ;
      RECT -23.305 -44.575 -23.205 -42.635 ;
      RECT -24.605 -44.575 -24.505 -42.635 ;
      RECT -25.905 -44.575 -25.805 -42.635 ;
      RECT -27.205 -44.575 -27.105 -42.635 ;
      RECT -28.505 -44.575 -28.405 -42.635 ;
      RECT -29.805 -44.575 -29.705 -42.635 ;
      RECT -31.105 -44.575 -31.005 -42.635 ;
      RECT -39.505 -43.945 -0.765 -43.265 ;
      RECT -1.205 -38.295 -1.105 -35.995 ;
      RECT -1.725 -38.295 -1.625 -35.995 ;
      RECT -2.505 -38.295 -2.405 -35.995 ;
      RECT -3.025 -38.295 -2.925 -35.995 ;
      RECT -3.805 -38.295 -3.705 -35.995 ;
      RECT -4.325 -38.295 -4.225 -35.995 ;
      RECT -5.105 -38.295 -5.005 -35.995 ;
      RECT -5.625 -38.295 -5.525 -35.995 ;
      RECT -6.405 -38.295 -6.305 -35.995 ;
      RECT -6.925 -38.295 -6.825 -35.995 ;
      RECT -7.705 -38.295 -7.605 -35.995 ;
      RECT -8.225 -38.295 -8.125 -35.995 ;
      RECT -9.005 -38.295 -8.905 -35.995 ;
      RECT -9.525 -38.295 -9.425 -35.995 ;
      RECT -10.305 -38.295 -10.205 -35.995 ;
      RECT -10.825 -38.295 -10.725 -35.995 ;
      RECT -11.605 -38.295 -11.505 -35.995 ;
      RECT -12.125 -38.295 -12.025 -35.995 ;
      RECT -12.905 -38.295 -12.805 -35.995 ;
      RECT -13.425 -38.295 -13.325 -35.995 ;
      RECT -14.205 -38.295 -14.105 -35.995 ;
      RECT -14.725 -38.295 -14.625 -35.995 ;
      RECT -15.505 -38.295 -15.405 -35.995 ;
      RECT -16.025 -38.295 -15.925 -35.995 ;
      RECT -16.805 -38.295 -16.705 -35.995 ;
      RECT -17.325 -38.295 -17.225 -35.995 ;
      RECT -18.105 -38.295 -18.005 -35.995 ;
      RECT -18.625 -38.295 -18.525 -35.995 ;
      RECT -19.405 -38.295 -19.305 -35.995 ;
      RECT -19.925 -38.295 -19.825 -35.995 ;
      RECT -20.705 -38.295 -20.605 -35.995 ;
      RECT -21.225 -38.295 -21.125 -35.995 ;
      RECT -22.005 -38.295 -21.905 -35.995 ;
      RECT -22.525 -38.295 -22.425 -35.995 ;
      RECT -23.305 -38.295 -23.205 -35.995 ;
      RECT -23.825 -38.295 -23.725 -35.995 ;
      RECT -24.605 -38.295 -24.505 -35.995 ;
      RECT -25.125 -38.295 -25.025 -35.995 ;
      RECT -25.905 -38.295 -25.805 -35.995 ;
      RECT -26.425 -38.295 -26.325 -35.995 ;
      RECT -27.205 -38.295 -27.105 -35.995 ;
      RECT -27.725 -38.295 -27.625 -35.995 ;
      RECT -28.505 -38.295 -28.405 -35.995 ;
      RECT -29.025 -38.295 -28.925 -35.995 ;
      RECT -29.805 -38.295 -29.705 -35.995 ;
      RECT -30.325 -38.295 -30.225 -35.995 ;
      RECT -31.105 -38.295 -31.005 -35.995 ;
      RECT -31.625 -38.295 -31.525 -35.995 ;
      RECT -37.505 -37.485 -0.765 -36.805 ;
      RECT -1.985 -31.835 -1.885 -29.535 ;
      RECT -3.285 -31.835 -3.185 -29.535 ;
      RECT -4.585 -31.835 -4.485 -29.535 ;
      RECT -5.885 -31.835 -5.785 -29.535 ;
      RECT -7.185 -31.835 -7.085 -29.535 ;
      RECT -8.485 -31.835 -8.385 -29.535 ;
      RECT -9.785 -31.835 -9.685 -29.535 ;
      RECT -11.085 -31.835 -10.985 -29.535 ;
      RECT -12.385 -31.835 -12.285 -29.535 ;
      RECT -13.685 -31.835 -13.585 -29.535 ;
      RECT -14.985 -31.835 -14.885 -29.535 ;
      RECT -16.285 -31.835 -16.185 -29.535 ;
      RECT -17.585 -31.835 -17.485 -29.535 ;
      RECT -18.885 -31.835 -18.785 -29.535 ;
      RECT -20.185 -31.835 -20.085 -29.535 ;
      RECT -21.485 -31.835 -21.385 -29.535 ;
      RECT -22.785 -31.835 -22.685 -29.535 ;
      RECT -24.085 -31.835 -23.985 -29.535 ;
      RECT -25.385 -31.835 -25.285 -29.535 ;
      RECT -26.685 -31.835 -26.585 -29.535 ;
      RECT -27.985 -31.835 -27.885 -29.535 ;
      RECT -29.285 -31.835 -29.185 -29.535 ;
      RECT -30.585 -31.835 -30.485 -29.535 ;
      RECT -31.885 -31.835 -31.785 -29.535 ;
      RECT -1.205 -31.655 -1.105 -29.715 ;
      RECT -2.505 -31.655 -2.405 -29.715 ;
      RECT -3.805 -31.655 -3.705 -29.715 ;
      RECT -5.105 -31.655 -5.005 -29.715 ;
      RECT -6.405 -31.655 -6.305 -29.715 ;
      RECT -7.705 -31.655 -7.605 -29.715 ;
      RECT -9.005 -31.655 -8.905 -29.715 ;
      RECT -10.305 -31.655 -10.205 -29.715 ;
      RECT -11.605 -31.655 -11.505 -29.715 ;
      RECT -12.905 -31.655 -12.805 -29.715 ;
      RECT -14.205 -31.655 -14.105 -29.715 ;
      RECT -15.505 -31.655 -15.405 -29.715 ;
      RECT -16.805 -31.655 -16.705 -29.715 ;
      RECT -18.105 -31.655 -18.005 -29.715 ;
      RECT -19.405 -31.655 -19.305 -29.715 ;
      RECT -20.705 -31.655 -20.605 -29.715 ;
      RECT -22.005 -31.655 -21.905 -29.715 ;
      RECT -23.305 -31.655 -23.205 -29.715 ;
      RECT -24.605 -31.655 -24.505 -29.715 ;
      RECT -25.905 -31.655 -25.805 -29.715 ;
      RECT -27.205 -31.655 -27.105 -29.715 ;
      RECT -28.505 -31.655 -28.405 -29.715 ;
      RECT -29.805 -31.655 -29.705 -29.715 ;
      RECT -31.105 -31.655 -31.005 -29.715 ;
      RECT -39.505 -31.025 -0.765 -30.345 ;
      RECT -1.205 -25.375 -1.105 -23.075 ;
      RECT -1.725 -25.375 -1.625 -23.075 ;
      RECT -2.505 -25.375 -2.405 -23.075 ;
      RECT -3.025 -25.375 -2.925 -23.075 ;
      RECT -3.805 -25.375 -3.705 -23.075 ;
      RECT -4.325 -25.375 -4.225 -23.075 ;
      RECT -5.105 -25.375 -5.005 -23.075 ;
      RECT -5.625 -25.375 -5.525 -23.075 ;
      RECT -6.405 -25.375 -6.305 -23.075 ;
      RECT -6.925 -25.375 -6.825 -23.075 ;
      RECT -7.705 -25.375 -7.605 -23.075 ;
      RECT -8.225 -25.375 -8.125 -23.075 ;
      RECT -9.005 -25.375 -8.905 -23.075 ;
      RECT -9.525 -25.375 -9.425 -23.075 ;
      RECT -10.305 -25.375 -10.205 -23.075 ;
      RECT -10.825 -25.375 -10.725 -23.075 ;
      RECT -11.605 -25.375 -11.505 -23.075 ;
      RECT -12.125 -25.375 -12.025 -23.075 ;
      RECT -12.905 -25.375 -12.805 -23.075 ;
      RECT -13.425 -25.375 -13.325 -23.075 ;
      RECT -14.205 -25.375 -14.105 -23.075 ;
      RECT -14.725 -25.375 -14.625 -23.075 ;
      RECT -15.505 -25.375 -15.405 -23.075 ;
      RECT -16.025 -25.375 -15.925 -23.075 ;
      RECT -16.805 -25.375 -16.705 -23.075 ;
      RECT -17.325 -25.375 -17.225 -23.075 ;
      RECT -18.105 -25.375 -18.005 -23.075 ;
      RECT -18.625 -25.375 -18.525 -23.075 ;
      RECT -19.405 -25.375 -19.305 -23.075 ;
      RECT -19.925 -25.375 -19.825 -23.075 ;
      RECT -20.705 -25.375 -20.605 -23.075 ;
      RECT -21.225 -25.375 -21.125 -23.075 ;
      RECT -22.005 -25.375 -21.905 -23.075 ;
      RECT -22.525 -25.375 -22.425 -23.075 ;
      RECT -23.305 -25.375 -23.205 -23.075 ;
      RECT -23.825 -25.375 -23.725 -23.075 ;
      RECT -24.605 -25.375 -24.505 -23.075 ;
      RECT -25.125 -25.375 -25.025 -23.075 ;
      RECT -25.905 -25.375 -25.805 -23.075 ;
      RECT -26.425 -25.375 -26.325 -23.075 ;
      RECT -27.205 -25.375 -27.105 -23.075 ;
      RECT -27.725 -25.375 -27.625 -23.075 ;
      RECT -28.505 -25.375 -28.405 -23.075 ;
      RECT -29.025 -25.375 -28.925 -23.075 ;
      RECT -29.805 -25.375 -29.705 -23.075 ;
      RECT -30.325 -25.375 -30.225 -23.075 ;
      RECT -31.105 -25.375 -31.005 -23.075 ;
      RECT -31.625 -25.375 -31.525 -23.075 ;
      RECT -37.505 -24.565 -0.765 -23.885 ;
      RECT -1.985 -18.915 -1.885 -16.615 ;
      RECT -3.285 -18.915 -3.185 -16.615 ;
      RECT -4.585 -18.915 -4.485 -16.615 ;
      RECT -5.885 -18.915 -5.785 -16.615 ;
      RECT -7.185 -18.915 -7.085 -16.615 ;
      RECT -8.485 -18.915 -8.385 -16.615 ;
      RECT -9.785 -18.915 -9.685 -16.615 ;
      RECT -11.085 -18.915 -10.985 -16.615 ;
      RECT -12.385 -18.915 -12.285 -16.615 ;
      RECT -13.685 -18.915 -13.585 -16.615 ;
      RECT -14.985 -18.915 -14.885 -16.615 ;
      RECT -16.285 -18.915 -16.185 -16.615 ;
      RECT -17.585 -18.915 -17.485 -16.615 ;
      RECT -18.885 -18.915 -18.785 -16.615 ;
      RECT -20.185 -18.915 -20.085 -16.615 ;
      RECT -21.485 -18.915 -21.385 -16.615 ;
      RECT -22.785 -18.915 -22.685 -16.615 ;
      RECT -24.085 -18.915 -23.985 -16.615 ;
      RECT -25.385 -18.915 -25.285 -16.615 ;
      RECT -26.685 -18.915 -26.585 -16.615 ;
      RECT -27.985 -18.915 -27.885 -16.615 ;
      RECT -29.285 -18.915 -29.185 -16.615 ;
      RECT -30.585 -18.915 -30.485 -16.615 ;
      RECT -31.885 -18.915 -31.785 -16.615 ;
      RECT -1.205 -18.735 -1.105 -16.795 ;
      RECT -2.505 -18.735 -2.405 -16.795 ;
      RECT -3.805 -18.735 -3.705 -16.795 ;
      RECT -5.105 -18.735 -5.005 -16.795 ;
      RECT -6.405 -18.735 -6.305 -16.795 ;
      RECT -7.705 -18.735 -7.605 -16.795 ;
      RECT -9.005 -18.735 -8.905 -16.795 ;
      RECT -10.305 -18.735 -10.205 -16.795 ;
      RECT -11.605 -18.735 -11.505 -16.795 ;
      RECT -12.905 -18.735 -12.805 -16.795 ;
      RECT -14.205 -18.735 -14.105 -16.795 ;
      RECT -15.505 -18.735 -15.405 -16.795 ;
      RECT -16.805 -18.735 -16.705 -16.795 ;
      RECT -18.105 -18.735 -18.005 -16.795 ;
      RECT -19.405 -18.735 -19.305 -16.795 ;
      RECT -20.705 -18.735 -20.605 -16.795 ;
      RECT -22.005 -18.735 -21.905 -16.795 ;
      RECT -23.305 -18.735 -23.205 -16.795 ;
      RECT -24.605 -18.735 -24.505 -16.795 ;
      RECT -25.905 -18.735 -25.805 -16.795 ;
      RECT -27.205 -18.735 -27.105 -16.795 ;
      RECT -28.505 -18.735 -28.405 -16.795 ;
      RECT -29.805 -18.735 -29.705 -16.795 ;
      RECT -31.105 -18.735 -31.005 -16.795 ;
      RECT -39.505 -18.105 -0.765 -17.425 ;
      RECT -1.205 -12.455 -1.105 -10.155 ;
      RECT -1.725 -12.455 -1.625 -10.155 ;
      RECT -2.505 -12.455 -2.405 -10.155 ;
      RECT -3.025 -12.455 -2.925 -10.155 ;
      RECT -3.805 -12.455 -3.705 -10.155 ;
      RECT -4.325 -12.455 -4.225 -10.155 ;
      RECT -5.105 -12.455 -5.005 -10.155 ;
      RECT -5.625 -12.455 -5.525 -10.155 ;
      RECT -6.405 -12.455 -6.305 -10.155 ;
      RECT -6.925 -12.455 -6.825 -10.155 ;
      RECT -7.705 -12.455 -7.605 -10.155 ;
      RECT -8.225 -12.455 -8.125 -10.155 ;
      RECT -9.005 -12.455 -8.905 -10.155 ;
      RECT -9.525 -12.455 -9.425 -10.155 ;
      RECT -10.305 -12.455 -10.205 -10.155 ;
      RECT -10.825 -12.455 -10.725 -10.155 ;
      RECT -11.605 -12.455 -11.505 -10.155 ;
      RECT -12.125 -12.455 -12.025 -10.155 ;
      RECT -12.905 -12.455 -12.805 -10.155 ;
      RECT -13.425 -12.455 -13.325 -10.155 ;
      RECT -14.205 -12.455 -14.105 -10.155 ;
      RECT -14.725 -12.455 -14.625 -10.155 ;
      RECT -15.505 -12.455 -15.405 -10.155 ;
      RECT -16.025 -12.455 -15.925 -10.155 ;
      RECT -16.805 -12.455 -16.705 -10.155 ;
      RECT -17.325 -12.455 -17.225 -10.155 ;
      RECT -18.105 -12.455 -18.005 -10.155 ;
      RECT -18.625 -12.455 -18.525 -10.155 ;
      RECT -19.405 -12.455 -19.305 -10.155 ;
      RECT -19.925 -12.455 -19.825 -10.155 ;
      RECT -20.705 -12.455 -20.605 -10.155 ;
      RECT -21.225 -12.455 -21.125 -10.155 ;
      RECT -22.005 -12.455 -21.905 -10.155 ;
      RECT -22.525 -12.455 -22.425 -10.155 ;
      RECT -23.305 -12.455 -23.205 -10.155 ;
      RECT -23.825 -12.455 -23.725 -10.155 ;
      RECT -24.605 -12.455 -24.505 -10.155 ;
      RECT -25.125 -12.455 -25.025 -10.155 ;
      RECT -25.905 -12.455 -25.805 -10.155 ;
      RECT -26.425 -12.455 -26.325 -10.155 ;
      RECT -27.205 -12.455 -27.105 -10.155 ;
      RECT -27.725 -12.455 -27.625 -10.155 ;
      RECT -28.505 -12.455 -28.405 -10.155 ;
      RECT -29.025 -12.455 -28.925 -10.155 ;
      RECT -29.805 -12.455 -29.705 -10.155 ;
      RECT -30.325 -12.455 -30.225 -10.155 ;
      RECT -31.105 -12.455 -31.005 -10.155 ;
      RECT -31.625 -12.455 -31.525 -10.155 ;
      RECT -37.505 -11.645 -0.765 -10.965 ;
      RECT -1.985 -5.995 -1.885 -3.695 ;
      RECT -3.285 -5.995 -3.185 -3.695 ;
      RECT -4.585 -5.995 -4.485 -3.695 ;
      RECT -5.885 -5.995 -5.785 -3.695 ;
      RECT -7.185 -5.995 -7.085 -3.695 ;
      RECT -8.485 -5.995 -8.385 -3.695 ;
      RECT -9.785 -5.995 -9.685 -3.695 ;
      RECT -11.085 -5.995 -10.985 -3.695 ;
      RECT -12.385 -5.995 -12.285 -3.695 ;
      RECT -13.685 -5.995 -13.585 -3.695 ;
      RECT -14.985 -5.995 -14.885 -3.695 ;
      RECT -16.285 -5.995 -16.185 -3.695 ;
      RECT -17.585 -5.995 -17.485 -3.695 ;
      RECT -18.885 -5.995 -18.785 -3.695 ;
      RECT -20.185 -5.995 -20.085 -3.695 ;
      RECT -21.485 -5.995 -21.385 -3.695 ;
      RECT -22.785 -5.995 -22.685 -3.695 ;
      RECT -24.085 -5.995 -23.985 -3.695 ;
      RECT -25.385 -5.995 -25.285 -3.695 ;
      RECT -26.685 -5.995 -26.585 -3.695 ;
      RECT -27.985 -5.995 -27.885 -3.695 ;
      RECT -29.285 -5.995 -29.185 -3.695 ;
      RECT -30.585 -5.995 -30.485 -3.695 ;
      RECT -31.885 -5.995 -31.785 -3.695 ;
      RECT -1.205 -5.815 -1.105 -3.875 ;
      RECT -2.505 -5.815 -2.405 -3.875 ;
      RECT -3.805 -5.815 -3.705 -3.875 ;
      RECT -5.105 -5.815 -5.005 -3.875 ;
      RECT -6.405 -5.815 -6.305 -3.875 ;
      RECT -7.705 -5.815 -7.605 -3.875 ;
      RECT -9.005 -5.815 -8.905 -3.875 ;
      RECT -10.305 -5.815 -10.205 -3.875 ;
      RECT -11.605 -5.815 -11.505 -3.875 ;
      RECT -12.905 -5.815 -12.805 -3.875 ;
      RECT -14.205 -5.815 -14.105 -3.875 ;
      RECT -15.505 -5.815 -15.405 -3.875 ;
      RECT -16.805 -5.815 -16.705 -3.875 ;
      RECT -18.105 -5.815 -18.005 -3.875 ;
      RECT -19.405 -5.815 -19.305 -3.875 ;
      RECT -20.705 -5.815 -20.605 -3.875 ;
      RECT -22.005 -5.815 -21.905 -3.875 ;
      RECT -23.305 -5.815 -23.205 -3.875 ;
      RECT -24.605 -5.815 -24.505 -3.875 ;
      RECT -25.905 -5.815 -25.805 -3.875 ;
      RECT -27.205 -5.815 -27.105 -3.875 ;
      RECT -28.505 -5.815 -28.405 -3.875 ;
      RECT -29.805 -5.815 -29.705 -3.875 ;
      RECT -31.105 -5.815 -31.005 -3.875 ;
      RECT -39.505 -5.185 -0.765 -4.505 ;
      RECT -32.505 1.275 -32.405 2.645 ;
      RECT -33.105 1.275 -33.005 2.645 ;
      RECT -33.705 1.275 -33.605 2.645 ;
      RECT -34.305 1.275 -34.205 2.645 ;
      RECT -34.905 1.275 -34.805 2.645 ;
      RECT -35.505 1.275 -35.405 2.645 ;
      RECT -6.065 1.275 -5.965 2.59 ;
      RECT -6.625 1.275 -6.525 2.59 ;
      RECT -37.505 1.275 -0.765 1.955 ;
      RECT -1.205 0.465 -1.105 1.955 ;
      RECT -1.725 0.465 -1.625 1.955 ;
      RECT -2.505 0.465 -2.405 1.955 ;
      RECT -3.025 0.465 -2.925 1.955 ;
      RECT -3.805 0.465 -3.705 1.955 ;
      RECT -4.325 0.465 -4.225 1.955 ;
      RECT -5.105 0.465 -5.005 1.955 ;
      RECT -5.625 0.465 -5.525 1.955 ;
      RECT -6.405 0.465 -6.305 1.955 ;
      RECT -6.925 0.465 -6.825 1.955 ;
      RECT -7.705 0.465 -7.605 1.955 ;
      RECT -8.225 0.465 -8.125 1.955 ;
      RECT -9.005 0.465 -8.905 1.955 ;
      RECT -9.525 0.465 -9.425 1.955 ;
      RECT -10.305 0.465 -10.205 1.955 ;
      RECT -10.825 0.465 -10.725 1.955 ;
      RECT -11.605 0.465 -11.505 1.955 ;
      RECT -12.125 0.465 -12.025 1.955 ;
      RECT -12.905 0.465 -12.805 1.955 ;
      RECT -13.425 0.465 -13.325 1.955 ;
      RECT -14.205 0.465 -14.105 1.955 ;
      RECT -14.725 0.465 -14.625 1.955 ;
      RECT -15.505 0.465 -15.405 1.955 ;
      RECT -16.025 0.465 -15.925 1.955 ;
      RECT -16.805 0.465 -16.705 1.955 ;
      RECT -17.325 0.465 -17.225 1.955 ;
      RECT -18.105 0.465 -18.005 1.955 ;
      RECT -18.625 0.465 -18.525 1.955 ;
      RECT -19.405 0.465 -19.305 1.955 ;
      RECT -19.925 0.465 -19.825 1.955 ;
      RECT -20.705 0.465 -20.605 1.955 ;
      RECT -21.225 0.465 -21.125 1.955 ;
      RECT -22.005 0.465 -21.905 1.955 ;
      RECT -22.525 0.465 -22.425 1.955 ;
      RECT -23.305 0.465 -23.205 1.955 ;
      RECT -23.825 0.465 -23.725 1.955 ;
      RECT -24.605 0.465 -24.505 1.955 ;
      RECT -25.125 0.465 -25.025 1.955 ;
      RECT -25.905 0.465 -25.805 1.955 ;
      RECT -26.425 0.465 -26.325 1.955 ;
      RECT -27.205 0.465 -27.105 1.955 ;
      RECT -27.725 0.465 -27.625 1.955 ;
      RECT -28.505 0.465 -28.405 1.955 ;
      RECT -29.025 0.465 -28.925 1.955 ;
      RECT -29.805 0.465 -29.705 1.955 ;
      RECT -30.325 0.465 -30.225 1.955 ;
      RECT -31.105 0.465 -31.005 1.955 ;
      RECT -31.625 0.465 -31.525 1.955 ;
      RECT -6.345 2.91 -5.615 3.03 ;
      RECT -5.785 2.22 -5.615 3.03 ;
      RECT -6.345 2.22 -6.245 3.03 ;
      RECT -6.665 -103.115 -6.565 -102.295 ;
      RECT -7.185 -103.115 -7.085 -102.295 ;
      RECT -7.185 -103.115 -6.14 -103.015 ;
      RECT -7.185 -100.475 -6.14 -100.375 ;
      RECT -6.665 -101.195 -6.565 -100.375 ;
      RECT -7.185 -101.195 -7.085 -100.375 ;
      RECT -6.665 -90.195 -6.565 -89.375 ;
      RECT -7.185 -90.195 -7.085 -89.375 ;
      RECT -7.185 -90.195 -6.14 -90.095 ;
      RECT -7.185 -87.555 -6.14 -87.455 ;
      RECT -6.665 -88.275 -6.565 -87.455 ;
      RECT -7.185 -88.275 -7.085 -87.455 ;
      RECT -6.665 -77.275 -6.565 -76.455 ;
      RECT -7.185 -77.275 -7.085 -76.455 ;
      RECT -7.185 -77.275 -6.14 -77.175 ;
      RECT -7.185 -74.635 -6.14 -74.535 ;
      RECT -6.665 -75.355 -6.565 -74.535 ;
      RECT -7.185 -75.355 -7.085 -74.535 ;
      RECT -6.665 -64.355 -6.565 -63.535 ;
      RECT -7.185 -64.355 -7.085 -63.535 ;
      RECT -7.185 -64.355 -6.14 -64.255 ;
      RECT -7.185 -61.715 -6.14 -61.615 ;
      RECT -6.665 -62.435 -6.565 -61.615 ;
      RECT -7.185 -62.435 -7.085 -61.615 ;
      RECT -6.665 -51.435 -6.565 -50.615 ;
      RECT -7.185 -51.435 -7.085 -50.615 ;
      RECT -7.185 -51.435 -6.14 -51.335 ;
      RECT -7.185 -48.795 -6.14 -48.695 ;
      RECT -6.665 -49.515 -6.565 -48.695 ;
      RECT -7.185 -49.515 -7.085 -48.695 ;
      RECT -6.665 -38.515 -6.565 -37.695 ;
      RECT -7.185 -38.515 -7.085 -37.695 ;
      RECT -7.185 -38.515 -6.14 -38.415 ;
      RECT -7.185 -35.875 -6.14 -35.775 ;
      RECT -6.665 -36.595 -6.565 -35.775 ;
      RECT -7.185 -36.595 -7.085 -35.775 ;
      RECT -6.665 -25.595 -6.565 -24.775 ;
      RECT -7.185 -25.595 -7.085 -24.775 ;
      RECT -7.185 -25.595 -6.14 -25.495 ;
      RECT -7.185 -22.955 -6.14 -22.855 ;
      RECT -6.665 -23.675 -6.565 -22.855 ;
      RECT -7.185 -23.675 -7.085 -22.855 ;
      RECT -6.665 -12.675 -6.565 -11.855 ;
      RECT -7.185 -12.675 -7.085 -11.855 ;
      RECT -7.185 -12.675 -6.14 -12.575 ;
      RECT -7.185 -10.035 -6.14 -9.935 ;
      RECT -6.665 -10.755 -6.565 -9.935 ;
      RECT -7.185 -10.755 -7.085 -9.935 ;
      RECT -6.665 0.245 -6.565 1.065 ;
      RECT -7.185 0.245 -7.085 1.065 ;
      RECT -7.185 0.245 -6.14 0.345 ;
      RECT -7.965 -103.115 -7.865 -102.295 ;
      RECT -8.485 -103.115 -8.385 -102.295 ;
      RECT -8.485 -103.115 -7.44 -103.015 ;
      RECT -8.485 -100.475 -7.44 -100.375 ;
      RECT -7.965 -101.195 -7.865 -100.375 ;
      RECT -8.485 -101.195 -8.385 -100.375 ;
      RECT -7.965 -90.195 -7.865 -89.375 ;
      RECT -8.485 -90.195 -8.385 -89.375 ;
      RECT -8.485 -90.195 -7.44 -90.095 ;
      RECT -8.485 -87.555 -7.44 -87.455 ;
      RECT -7.965 -88.275 -7.865 -87.455 ;
      RECT -8.485 -88.275 -8.385 -87.455 ;
      RECT -7.965 -77.275 -7.865 -76.455 ;
      RECT -8.485 -77.275 -8.385 -76.455 ;
      RECT -8.485 -77.275 -7.44 -77.175 ;
      RECT -8.485 -74.635 -7.44 -74.535 ;
      RECT -7.965 -75.355 -7.865 -74.535 ;
      RECT -8.485 -75.355 -8.385 -74.535 ;
      RECT -7.965 -64.355 -7.865 -63.535 ;
      RECT -8.485 -64.355 -8.385 -63.535 ;
      RECT -8.485 -64.355 -7.44 -64.255 ;
      RECT -8.485 -61.715 -7.44 -61.615 ;
      RECT -7.965 -62.435 -7.865 -61.615 ;
      RECT -8.485 -62.435 -8.385 -61.615 ;
      RECT -7.965 -51.435 -7.865 -50.615 ;
      RECT -8.485 -51.435 -8.385 -50.615 ;
      RECT -8.485 -51.435 -7.44 -51.335 ;
      RECT -8.485 -48.795 -7.44 -48.695 ;
      RECT -7.965 -49.515 -7.865 -48.695 ;
      RECT -8.485 -49.515 -8.385 -48.695 ;
      RECT -7.965 -38.515 -7.865 -37.695 ;
      RECT -8.485 -38.515 -8.385 -37.695 ;
      RECT -8.485 -38.515 -7.44 -38.415 ;
      RECT -8.485 -35.875 -7.44 -35.775 ;
      RECT -7.965 -36.595 -7.865 -35.775 ;
      RECT -8.485 -36.595 -8.385 -35.775 ;
      RECT -7.965 -25.595 -7.865 -24.775 ;
      RECT -8.485 -25.595 -8.385 -24.775 ;
      RECT -8.485 -25.595 -7.44 -25.495 ;
      RECT -8.485 -22.955 -7.44 -22.855 ;
      RECT -7.965 -23.675 -7.865 -22.855 ;
      RECT -8.485 -23.675 -8.385 -22.855 ;
      RECT -7.965 -12.675 -7.865 -11.855 ;
      RECT -8.485 -12.675 -8.385 -11.855 ;
      RECT -8.485 -12.675 -7.44 -12.575 ;
      RECT -8.485 -10.035 -7.44 -9.935 ;
      RECT -7.965 -10.755 -7.865 -9.935 ;
      RECT -8.485 -10.755 -8.385 -9.935 ;
      RECT -7.965 0.245 -7.865 1.065 ;
      RECT -8.485 0.245 -8.385 1.065 ;
      RECT -8.485 0.245 -7.44 0.345 ;
      RECT -9.265 -103.115 -9.165 -102.295 ;
      RECT -9.785 -103.115 -9.685 -102.295 ;
      RECT -9.785 -103.115 -8.74 -103.015 ;
      RECT -9.785 -100.475 -8.74 -100.375 ;
      RECT -9.265 -101.195 -9.165 -100.375 ;
      RECT -9.785 -101.195 -9.685 -100.375 ;
      RECT -9.265 -90.195 -9.165 -89.375 ;
      RECT -9.785 -90.195 -9.685 -89.375 ;
      RECT -9.785 -90.195 -8.74 -90.095 ;
      RECT -9.785 -87.555 -8.74 -87.455 ;
      RECT -9.265 -88.275 -9.165 -87.455 ;
      RECT -9.785 -88.275 -9.685 -87.455 ;
      RECT -9.265 -77.275 -9.165 -76.455 ;
      RECT -9.785 -77.275 -9.685 -76.455 ;
      RECT -9.785 -77.275 -8.74 -77.175 ;
      RECT -9.785 -74.635 -8.74 -74.535 ;
      RECT -9.265 -75.355 -9.165 -74.535 ;
      RECT -9.785 -75.355 -9.685 -74.535 ;
      RECT -9.265 -64.355 -9.165 -63.535 ;
      RECT -9.785 -64.355 -9.685 -63.535 ;
      RECT -9.785 -64.355 -8.74 -64.255 ;
      RECT -9.785 -61.715 -8.74 -61.615 ;
      RECT -9.265 -62.435 -9.165 -61.615 ;
      RECT -9.785 -62.435 -9.685 -61.615 ;
      RECT -9.265 -51.435 -9.165 -50.615 ;
      RECT -9.785 -51.435 -9.685 -50.615 ;
      RECT -9.785 -51.435 -8.74 -51.335 ;
      RECT -9.785 -48.795 -8.74 -48.695 ;
      RECT -9.265 -49.515 -9.165 -48.695 ;
      RECT -9.785 -49.515 -9.685 -48.695 ;
      RECT -9.265 -38.515 -9.165 -37.695 ;
      RECT -9.785 -38.515 -9.685 -37.695 ;
      RECT -9.785 -38.515 -8.74 -38.415 ;
      RECT -9.785 -35.875 -8.74 -35.775 ;
      RECT -9.265 -36.595 -9.165 -35.775 ;
      RECT -9.785 -36.595 -9.685 -35.775 ;
      RECT -9.265 -25.595 -9.165 -24.775 ;
      RECT -9.785 -25.595 -9.685 -24.775 ;
      RECT -9.785 -25.595 -8.74 -25.495 ;
      RECT -9.785 -22.955 -8.74 -22.855 ;
      RECT -9.265 -23.675 -9.165 -22.855 ;
      RECT -9.785 -23.675 -9.685 -22.855 ;
      RECT -9.265 -12.675 -9.165 -11.855 ;
      RECT -9.785 -12.675 -9.685 -11.855 ;
      RECT -9.785 -12.675 -8.74 -12.575 ;
      RECT -9.785 -10.035 -8.74 -9.935 ;
      RECT -9.265 -10.755 -9.165 -9.935 ;
      RECT -9.785 -10.755 -9.685 -9.935 ;
      RECT -9.265 0.245 -9.165 1.065 ;
      RECT -9.785 0.245 -9.685 1.065 ;
      RECT -9.785 0.245 -8.74 0.345 ;
      RECT -10.565 -103.115 -10.465 -102.295 ;
      RECT -11.085 -103.115 -10.985 -102.295 ;
      RECT -11.085 -103.115 -10.04 -103.015 ;
      RECT -11.085 -100.475 -10.04 -100.375 ;
      RECT -10.565 -101.195 -10.465 -100.375 ;
      RECT -11.085 -101.195 -10.985 -100.375 ;
      RECT -10.565 -90.195 -10.465 -89.375 ;
      RECT -11.085 -90.195 -10.985 -89.375 ;
      RECT -11.085 -90.195 -10.04 -90.095 ;
      RECT -11.085 -87.555 -10.04 -87.455 ;
      RECT -10.565 -88.275 -10.465 -87.455 ;
      RECT -11.085 -88.275 -10.985 -87.455 ;
      RECT -10.565 -77.275 -10.465 -76.455 ;
      RECT -11.085 -77.275 -10.985 -76.455 ;
      RECT -11.085 -77.275 -10.04 -77.175 ;
      RECT -11.085 -74.635 -10.04 -74.535 ;
      RECT -10.565 -75.355 -10.465 -74.535 ;
      RECT -11.085 -75.355 -10.985 -74.535 ;
      RECT -10.565 -64.355 -10.465 -63.535 ;
      RECT -11.085 -64.355 -10.985 -63.535 ;
      RECT -11.085 -64.355 -10.04 -64.255 ;
      RECT -11.085 -61.715 -10.04 -61.615 ;
      RECT -10.565 -62.435 -10.465 -61.615 ;
      RECT -11.085 -62.435 -10.985 -61.615 ;
      RECT -10.565 -51.435 -10.465 -50.615 ;
      RECT -11.085 -51.435 -10.985 -50.615 ;
      RECT -11.085 -51.435 -10.04 -51.335 ;
      RECT -11.085 -48.795 -10.04 -48.695 ;
      RECT -10.565 -49.515 -10.465 -48.695 ;
      RECT -11.085 -49.515 -10.985 -48.695 ;
      RECT -10.565 -38.515 -10.465 -37.695 ;
      RECT -11.085 -38.515 -10.985 -37.695 ;
      RECT -11.085 -38.515 -10.04 -38.415 ;
      RECT -11.085 -35.875 -10.04 -35.775 ;
      RECT -10.565 -36.595 -10.465 -35.775 ;
      RECT -11.085 -36.595 -10.985 -35.775 ;
      RECT -10.565 -25.595 -10.465 -24.775 ;
      RECT -11.085 -25.595 -10.985 -24.775 ;
      RECT -11.085 -25.595 -10.04 -25.495 ;
      RECT -11.085 -22.955 -10.04 -22.855 ;
      RECT -10.565 -23.675 -10.465 -22.855 ;
      RECT -11.085 -23.675 -10.985 -22.855 ;
      RECT -10.565 -12.675 -10.465 -11.855 ;
      RECT -11.085 -12.675 -10.985 -11.855 ;
      RECT -11.085 -12.675 -10.04 -12.575 ;
      RECT -11.085 -10.035 -10.04 -9.935 ;
      RECT -10.565 -10.755 -10.465 -9.935 ;
      RECT -11.085 -10.755 -10.985 -9.935 ;
      RECT -10.565 0.245 -10.465 1.065 ;
      RECT -11.085 0.245 -10.985 1.065 ;
      RECT -11.085 0.245 -10.04 0.345 ;
      RECT -11.705 -111.525 -11.605 -110.155 ;
      RECT -12.305 -111.525 -12.205 -110.155 ;
      RECT -37.505 -111.525 -11.145 -110.845 ;
      RECT -12.385 -100.475 -11.34 -100.375 ;
      RECT -11.865 -101.195 -11.765 -100.375 ;
      RECT -12.385 -101.195 -12.285 -100.375 ;
      RECT -11.865 -90.195 -11.765 -89.375 ;
      RECT -12.385 -90.195 -12.285 -89.375 ;
      RECT -12.385 -90.195 -11.34 -90.095 ;
      RECT -12.385 -87.555 -11.34 -87.455 ;
      RECT -11.865 -88.275 -11.765 -87.455 ;
      RECT -12.385 -88.275 -12.285 -87.455 ;
      RECT -11.865 -77.275 -11.765 -76.455 ;
      RECT -12.385 -77.275 -12.285 -76.455 ;
      RECT -12.385 -77.275 -11.34 -77.175 ;
      RECT -12.385 -74.635 -11.34 -74.535 ;
      RECT -11.865 -75.355 -11.765 -74.535 ;
      RECT -12.385 -75.355 -12.285 -74.535 ;
      RECT -11.865 -64.355 -11.765 -63.535 ;
      RECT -12.385 -64.355 -12.285 -63.535 ;
      RECT -12.385 -64.355 -11.34 -64.255 ;
      RECT -12.385 -61.715 -11.34 -61.615 ;
      RECT -11.865 -62.435 -11.765 -61.615 ;
      RECT -12.385 -62.435 -12.285 -61.615 ;
      RECT -11.865 -51.435 -11.765 -50.615 ;
      RECT -12.385 -51.435 -12.285 -50.615 ;
      RECT -12.385 -51.435 -11.34 -51.335 ;
      RECT -12.385 -48.795 -11.34 -48.695 ;
      RECT -11.865 -49.515 -11.765 -48.695 ;
      RECT -12.385 -49.515 -12.285 -48.695 ;
      RECT -11.865 -38.515 -11.765 -37.695 ;
      RECT -12.385 -38.515 -12.285 -37.695 ;
      RECT -12.385 -38.515 -11.34 -38.415 ;
      RECT -12.385 -35.875 -11.34 -35.775 ;
      RECT -11.865 -36.595 -11.765 -35.775 ;
      RECT -12.385 -36.595 -12.285 -35.775 ;
      RECT -11.865 -25.595 -11.765 -24.775 ;
      RECT -12.385 -25.595 -12.285 -24.775 ;
      RECT -12.385 -25.595 -11.34 -25.495 ;
      RECT -12.385 -22.955 -11.34 -22.855 ;
      RECT -11.865 -23.675 -11.765 -22.855 ;
      RECT -12.385 -23.675 -12.285 -22.855 ;
      RECT -11.865 -12.675 -11.765 -11.855 ;
      RECT -12.385 -12.675 -12.285 -11.855 ;
      RECT -12.385 -12.675 -11.34 -12.575 ;
      RECT -12.385 -10.035 -11.34 -9.935 ;
      RECT -11.865 -10.755 -11.765 -9.935 ;
      RECT -12.385 -10.755 -12.285 -9.935 ;
      RECT -11.865 0.245 -11.765 1.065 ;
      RECT -12.385 0.245 -12.285 1.065 ;
      RECT -12.385 0.245 -11.34 0.345 ;
      RECT -13.685 -100.475 -12.64 -100.375 ;
      RECT -13.165 -101.195 -13.065 -100.375 ;
      RECT -13.685 -101.195 -13.585 -100.375 ;
      RECT -13.165 -90.195 -13.065 -89.375 ;
      RECT -13.685 -90.195 -13.585 -89.375 ;
      RECT -13.685 -90.195 -12.64 -90.095 ;
      RECT -13.685 -87.555 -12.64 -87.455 ;
      RECT -13.165 -88.275 -13.065 -87.455 ;
      RECT -13.685 -88.275 -13.585 -87.455 ;
      RECT -13.165 -77.275 -13.065 -76.455 ;
      RECT -13.685 -77.275 -13.585 -76.455 ;
      RECT -13.685 -77.275 -12.64 -77.175 ;
      RECT -13.685 -74.635 -12.64 -74.535 ;
      RECT -13.165 -75.355 -13.065 -74.535 ;
      RECT -13.685 -75.355 -13.585 -74.535 ;
      RECT -13.165 -64.355 -13.065 -63.535 ;
      RECT -13.685 -64.355 -13.585 -63.535 ;
      RECT -13.685 -64.355 -12.64 -64.255 ;
      RECT -13.685 -61.715 -12.64 -61.615 ;
      RECT -13.165 -62.435 -13.065 -61.615 ;
      RECT -13.685 -62.435 -13.585 -61.615 ;
      RECT -13.165 -51.435 -13.065 -50.615 ;
      RECT -13.685 -51.435 -13.585 -50.615 ;
      RECT -13.685 -51.435 -12.64 -51.335 ;
      RECT -13.685 -48.795 -12.64 -48.695 ;
      RECT -13.165 -49.515 -13.065 -48.695 ;
      RECT -13.685 -49.515 -13.585 -48.695 ;
      RECT -13.165 -38.515 -13.065 -37.695 ;
      RECT -13.685 -38.515 -13.585 -37.695 ;
      RECT -13.685 -38.515 -12.64 -38.415 ;
      RECT -13.685 -35.875 -12.64 -35.775 ;
      RECT -13.165 -36.595 -13.065 -35.775 ;
      RECT -13.685 -36.595 -13.585 -35.775 ;
      RECT -13.165 -25.595 -13.065 -24.775 ;
      RECT -13.685 -25.595 -13.585 -24.775 ;
      RECT -13.685 -25.595 -12.64 -25.495 ;
      RECT -13.685 -22.955 -12.64 -22.855 ;
      RECT -13.165 -23.675 -13.065 -22.855 ;
      RECT -13.685 -23.675 -13.585 -22.855 ;
      RECT -13.165 -12.675 -13.065 -11.855 ;
      RECT -13.685 -12.675 -13.585 -11.855 ;
      RECT -13.685 -12.675 -12.64 -12.575 ;
      RECT -13.685 -10.035 -12.64 -9.935 ;
      RECT -13.165 -10.755 -13.065 -9.935 ;
      RECT -13.685 -10.755 -13.585 -9.935 ;
      RECT -13.165 0.245 -13.065 1.065 ;
      RECT -13.685 0.245 -13.585 1.065 ;
      RECT -13.685 0.245 -12.64 0.345 ;
      RECT -14.985 -100.475 -13.94 -100.375 ;
      RECT -14.465 -101.195 -14.365 -100.375 ;
      RECT -14.985 -101.195 -14.885 -100.375 ;
      RECT -14.465 -90.195 -14.365 -89.375 ;
      RECT -14.985 -90.195 -14.885 -89.375 ;
      RECT -14.985 -90.195 -13.94 -90.095 ;
      RECT -14.985 -87.555 -13.94 -87.455 ;
      RECT -14.465 -88.275 -14.365 -87.455 ;
      RECT -14.985 -88.275 -14.885 -87.455 ;
      RECT -14.465 -77.275 -14.365 -76.455 ;
      RECT -14.985 -77.275 -14.885 -76.455 ;
      RECT -14.985 -77.275 -13.94 -77.175 ;
      RECT -14.985 -74.635 -13.94 -74.535 ;
      RECT -14.465 -75.355 -14.365 -74.535 ;
      RECT -14.985 -75.355 -14.885 -74.535 ;
      RECT -14.465 -64.355 -14.365 -63.535 ;
      RECT -14.985 -64.355 -14.885 -63.535 ;
      RECT -14.985 -64.355 -13.94 -64.255 ;
      RECT -14.985 -61.715 -13.94 -61.615 ;
      RECT -14.465 -62.435 -14.365 -61.615 ;
      RECT -14.985 -62.435 -14.885 -61.615 ;
      RECT -14.465 -51.435 -14.365 -50.615 ;
      RECT -14.985 -51.435 -14.885 -50.615 ;
      RECT -14.985 -51.435 -13.94 -51.335 ;
      RECT -14.985 -48.795 -13.94 -48.695 ;
      RECT -14.465 -49.515 -14.365 -48.695 ;
      RECT -14.985 -49.515 -14.885 -48.695 ;
      RECT -14.465 -38.515 -14.365 -37.695 ;
      RECT -14.985 -38.515 -14.885 -37.695 ;
      RECT -14.985 -38.515 -13.94 -38.415 ;
      RECT -14.985 -35.875 -13.94 -35.775 ;
      RECT -14.465 -36.595 -14.365 -35.775 ;
      RECT -14.985 -36.595 -14.885 -35.775 ;
      RECT -14.465 -25.595 -14.365 -24.775 ;
      RECT -14.985 -25.595 -14.885 -24.775 ;
      RECT -14.985 -25.595 -13.94 -25.495 ;
      RECT -14.985 -22.955 -13.94 -22.855 ;
      RECT -14.465 -23.675 -14.365 -22.855 ;
      RECT -14.985 -23.675 -14.885 -22.855 ;
      RECT -14.465 -12.675 -14.365 -11.855 ;
      RECT -14.985 -12.675 -14.885 -11.855 ;
      RECT -14.985 -12.675 -13.94 -12.575 ;
      RECT -14.985 -10.035 -13.94 -9.935 ;
      RECT -14.465 -10.755 -14.365 -9.935 ;
      RECT -14.985 -10.755 -14.885 -9.935 ;
      RECT -14.465 0.245 -14.365 1.065 ;
      RECT -14.985 0.245 -14.885 1.065 ;
      RECT -14.985 0.245 -13.94 0.345 ;
      RECT -16.285 -100.475 -15.24 -100.375 ;
      RECT -15.765 -101.195 -15.665 -100.375 ;
      RECT -16.285 -101.195 -16.185 -100.375 ;
      RECT -15.765 -90.195 -15.665 -89.375 ;
      RECT -16.285 -90.195 -16.185 -89.375 ;
      RECT -16.285 -90.195 -15.24 -90.095 ;
      RECT -16.285 -87.555 -15.24 -87.455 ;
      RECT -15.765 -88.275 -15.665 -87.455 ;
      RECT -16.285 -88.275 -16.185 -87.455 ;
      RECT -15.765 -77.275 -15.665 -76.455 ;
      RECT -16.285 -77.275 -16.185 -76.455 ;
      RECT -16.285 -77.275 -15.24 -77.175 ;
      RECT -16.285 -74.635 -15.24 -74.535 ;
      RECT -15.765 -75.355 -15.665 -74.535 ;
      RECT -16.285 -75.355 -16.185 -74.535 ;
      RECT -15.765 -64.355 -15.665 -63.535 ;
      RECT -16.285 -64.355 -16.185 -63.535 ;
      RECT -16.285 -64.355 -15.24 -64.255 ;
      RECT -16.285 -61.715 -15.24 -61.615 ;
      RECT -15.765 -62.435 -15.665 -61.615 ;
      RECT -16.285 -62.435 -16.185 -61.615 ;
      RECT -15.765 -51.435 -15.665 -50.615 ;
      RECT -16.285 -51.435 -16.185 -50.615 ;
      RECT -16.285 -51.435 -15.24 -51.335 ;
      RECT -16.285 -48.795 -15.24 -48.695 ;
      RECT -15.765 -49.515 -15.665 -48.695 ;
      RECT -16.285 -49.515 -16.185 -48.695 ;
      RECT -15.765 -38.515 -15.665 -37.695 ;
      RECT -16.285 -38.515 -16.185 -37.695 ;
      RECT -16.285 -38.515 -15.24 -38.415 ;
      RECT -16.285 -35.875 -15.24 -35.775 ;
      RECT -15.765 -36.595 -15.665 -35.775 ;
      RECT -16.285 -36.595 -16.185 -35.775 ;
      RECT -15.765 -25.595 -15.665 -24.775 ;
      RECT -16.285 -25.595 -16.185 -24.775 ;
      RECT -16.285 -25.595 -15.24 -25.495 ;
      RECT -16.285 -22.955 -15.24 -22.855 ;
      RECT -15.765 -23.675 -15.665 -22.855 ;
      RECT -16.285 -23.675 -16.185 -22.855 ;
      RECT -15.765 -12.675 -15.665 -11.855 ;
      RECT -16.285 -12.675 -16.185 -11.855 ;
      RECT -16.285 -12.675 -15.24 -12.575 ;
      RECT -16.285 -10.035 -15.24 -9.935 ;
      RECT -15.765 -10.755 -15.665 -9.935 ;
      RECT -16.285 -10.755 -16.185 -9.935 ;
      RECT -15.765 0.245 -15.665 1.065 ;
      RECT -16.285 0.245 -16.185 1.065 ;
      RECT -16.285 0.245 -15.24 0.345 ;
      RECT -17.585 -100.475 -16.54 -100.375 ;
      RECT -17.065 -101.195 -16.965 -100.375 ;
      RECT -17.585 -101.195 -17.485 -100.375 ;
      RECT -17.065 -90.195 -16.965 -89.375 ;
      RECT -17.585 -90.195 -17.485 -89.375 ;
      RECT -17.585 -90.195 -16.54 -90.095 ;
      RECT -17.585 -87.555 -16.54 -87.455 ;
      RECT -17.065 -88.275 -16.965 -87.455 ;
      RECT -17.585 -88.275 -17.485 -87.455 ;
      RECT -17.065 -77.275 -16.965 -76.455 ;
      RECT -17.585 -77.275 -17.485 -76.455 ;
      RECT -17.585 -77.275 -16.54 -77.175 ;
      RECT -17.585 -74.635 -16.54 -74.535 ;
      RECT -17.065 -75.355 -16.965 -74.535 ;
      RECT -17.585 -75.355 -17.485 -74.535 ;
      RECT -17.065 -64.355 -16.965 -63.535 ;
      RECT -17.585 -64.355 -17.485 -63.535 ;
      RECT -17.585 -64.355 -16.54 -64.255 ;
      RECT -17.585 -61.715 -16.54 -61.615 ;
      RECT -17.065 -62.435 -16.965 -61.615 ;
      RECT -17.585 -62.435 -17.485 -61.615 ;
      RECT -17.065 -51.435 -16.965 -50.615 ;
      RECT -17.585 -51.435 -17.485 -50.615 ;
      RECT -17.585 -51.435 -16.54 -51.335 ;
      RECT -17.585 -48.795 -16.54 -48.695 ;
      RECT -17.065 -49.515 -16.965 -48.695 ;
      RECT -17.585 -49.515 -17.485 -48.695 ;
      RECT -17.065 -38.515 -16.965 -37.695 ;
      RECT -17.585 -38.515 -17.485 -37.695 ;
      RECT -17.585 -38.515 -16.54 -38.415 ;
      RECT -17.585 -35.875 -16.54 -35.775 ;
      RECT -17.065 -36.595 -16.965 -35.775 ;
      RECT -17.585 -36.595 -17.485 -35.775 ;
      RECT -17.065 -25.595 -16.965 -24.775 ;
      RECT -17.585 -25.595 -17.485 -24.775 ;
      RECT -17.585 -25.595 -16.54 -25.495 ;
      RECT -17.585 -22.955 -16.54 -22.855 ;
      RECT -17.065 -23.675 -16.965 -22.855 ;
      RECT -17.585 -23.675 -17.485 -22.855 ;
      RECT -17.065 -12.675 -16.965 -11.855 ;
      RECT -17.585 -12.675 -17.485 -11.855 ;
      RECT -17.585 -12.675 -16.54 -12.575 ;
      RECT -17.585 -10.035 -16.54 -9.935 ;
      RECT -17.065 -10.755 -16.965 -9.935 ;
      RECT -17.585 -10.755 -17.485 -9.935 ;
      RECT -17.065 0.245 -16.965 1.065 ;
      RECT -17.585 0.245 -17.485 1.065 ;
      RECT -17.585 0.245 -16.54 0.345 ;
      RECT -18.885 -100.475 -17.84 -100.375 ;
      RECT -18.365 -101.195 -18.265 -100.375 ;
      RECT -18.885 -101.195 -18.785 -100.375 ;
      RECT -18.365 -90.195 -18.265 -89.375 ;
      RECT -18.885 -90.195 -18.785 -89.375 ;
      RECT -18.885 -90.195 -17.84 -90.095 ;
      RECT -18.885 -87.555 -17.84 -87.455 ;
      RECT -18.365 -88.275 -18.265 -87.455 ;
      RECT -18.885 -88.275 -18.785 -87.455 ;
      RECT -18.365 -77.275 -18.265 -76.455 ;
      RECT -18.885 -77.275 -18.785 -76.455 ;
      RECT -18.885 -77.275 -17.84 -77.175 ;
      RECT -18.885 -74.635 -17.84 -74.535 ;
      RECT -18.365 -75.355 -18.265 -74.535 ;
      RECT -18.885 -75.355 -18.785 -74.535 ;
      RECT -18.365 -64.355 -18.265 -63.535 ;
      RECT -18.885 -64.355 -18.785 -63.535 ;
      RECT -18.885 -64.355 -17.84 -64.255 ;
      RECT -18.885 -61.715 -17.84 -61.615 ;
      RECT -18.365 -62.435 -18.265 -61.615 ;
      RECT -18.885 -62.435 -18.785 -61.615 ;
      RECT -18.365 -51.435 -18.265 -50.615 ;
      RECT -18.885 -51.435 -18.785 -50.615 ;
      RECT -18.885 -51.435 -17.84 -51.335 ;
      RECT -18.885 -48.795 -17.84 -48.695 ;
      RECT -18.365 -49.515 -18.265 -48.695 ;
      RECT -18.885 -49.515 -18.785 -48.695 ;
      RECT -18.365 -38.515 -18.265 -37.695 ;
      RECT -18.885 -38.515 -18.785 -37.695 ;
      RECT -18.885 -38.515 -17.84 -38.415 ;
      RECT -18.885 -35.875 -17.84 -35.775 ;
      RECT -18.365 -36.595 -18.265 -35.775 ;
      RECT -18.885 -36.595 -18.785 -35.775 ;
      RECT -18.365 -25.595 -18.265 -24.775 ;
      RECT -18.885 -25.595 -18.785 -24.775 ;
      RECT -18.885 -25.595 -17.84 -25.495 ;
      RECT -18.885 -22.955 -17.84 -22.855 ;
      RECT -18.365 -23.675 -18.265 -22.855 ;
      RECT -18.885 -23.675 -18.785 -22.855 ;
      RECT -18.365 -12.675 -18.265 -11.855 ;
      RECT -18.885 -12.675 -18.785 -11.855 ;
      RECT -18.885 -12.675 -17.84 -12.575 ;
      RECT -18.885 -10.035 -17.84 -9.935 ;
      RECT -18.365 -10.755 -18.265 -9.935 ;
      RECT -18.885 -10.755 -18.785 -9.935 ;
      RECT -18.365 0.245 -18.265 1.065 ;
      RECT -18.885 0.245 -18.785 1.065 ;
      RECT -18.885 0.245 -17.84 0.345 ;
      RECT -20.185 -100.475 -19.14 -100.375 ;
      RECT -19.665 -101.195 -19.565 -100.375 ;
      RECT -20.185 -101.195 -20.085 -100.375 ;
      RECT -19.665 -90.195 -19.565 -89.375 ;
      RECT -20.185 -90.195 -20.085 -89.375 ;
      RECT -20.185 -90.195 -19.14 -90.095 ;
      RECT -20.185 -87.555 -19.14 -87.455 ;
      RECT -19.665 -88.275 -19.565 -87.455 ;
      RECT -20.185 -88.275 -20.085 -87.455 ;
      RECT -19.665 -77.275 -19.565 -76.455 ;
      RECT -20.185 -77.275 -20.085 -76.455 ;
      RECT -20.185 -77.275 -19.14 -77.175 ;
      RECT -20.185 -74.635 -19.14 -74.535 ;
      RECT -19.665 -75.355 -19.565 -74.535 ;
      RECT -20.185 -75.355 -20.085 -74.535 ;
      RECT -19.665 -64.355 -19.565 -63.535 ;
      RECT -20.185 -64.355 -20.085 -63.535 ;
      RECT -20.185 -64.355 -19.14 -64.255 ;
      RECT -20.185 -61.715 -19.14 -61.615 ;
      RECT -19.665 -62.435 -19.565 -61.615 ;
      RECT -20.185 -62.435 -20.085 -61.615 ;
      RECT -19.665 -51.435 -19.565 -50.615 ;
      RECT -20.185 -51.435 -20.085 -50.615 ;
      RECT -20.185 -51.435 -19.14 -51.335 ;
      RECT -20.185 -48.795 -19.14 -48.695 ;
      RECT -19.665 -49.515 -19.565 -48.695 ;
      RECT -20.185 -49.515 -20.085 -48.695 ;
      RECT -19.665 -38.515 -19.565 -37.695 ;
      RECT -20.185 -38.515 -20.085 -37.695 ;
      RECT -20.185 -38.515 -19.14 -38.415 ;
      RECT -20.185 -35.875 -19.14 -35.775 ;
      RECT -19.665 -36.595 -19.565 -35.775 ;
      RECT -20.185 -36.595 -20.085 -35.775 ;
      RECT -19.665 -25.595 -19.565 -24.775 ;
      RECT -20.185 -25.595 -20.085 -24.775 ;
      RECT -20.185 -25.595 -19.14 -25.495 ;
      RECT -20.185 -22.955 -19.14 -22.855 ;
      RECT -19.665 -23.675 -19.565 -22.855 ;
      RECT -20.185 -23.675 -20.085 -22.855 ;
      RECT -19.665 -12.675 -19.565 -11.855 ;
      RECT -20.185 -12.675 -20.085 -11.855 ;
      RECT -20.185 -12.675 -19.14 -12.575 ;
      RECT -20.185 -10.035 -19.14 -9.935 ;
      RECT -19.665 -10.755 -19.565 -9.935 ;
      RECT -20.185 -10.755 -20.085 -9.935 ;
      RECT -19.665 0.245 -19.565 1.065 ;
      RECT -20.185 0.245 -20.085 1.065 ;
      RECT -20.185 0.245 -19.14 0.345 ;
      RECT -21.485 -100.475 -20.44 -100.375 ;
      RECT -20.965 -101.195 -20.865 -100.375 ;
      RECT -21.485 -101.195 -21.385 -100.375 ;
      RECT -20.965 -90.195 -20.865 -89.375 ;
      RECT -21.485 -90.195 -21.385 -89.375 ;
      RECT -21.485 -90.195 -20.44 -90.095 ;
      RECT -21.485 -87.555 -20.44 -87.455 ;
      RECT -20.965 -88.275 -20.865 -87.455 ;
      RECT -21.485 -88.275 -21.385 -87.455 ;
      RECT -20.965 -77.275 -20.865 -76.455 ;
      RECT -21.485 -77.275 -21.385 -76.455 ;
      RECT -21.485 -77.275 -20.44 -77.175 ;
      RECT -21.485 -74.635 -20.44 -74.535 ;
      RECT -20.965 -75.355 -20.865 -74.535 ;
      RECT -21.485 -75.355 -21.385 -74.535 ;
      RECT -20.965 -64.355 -20.865 -63.535 ;
      RECT -21.485 -64.355 -21.385 -63.535 ;
      RECT -21.485 -64.355 -20.44 -64.255 ;
      RECT -21.485 -61.715 -20.44 -61.615 ;
      RECT -20.965 -62.435 -20.865 -61.615 ;
      RECT -21.485 -62.435 -21.385 -61.615 ;
      RECT -20.965 -51.435 -20.865 -50.615 ;
      RECT -21.485 -51.435 -21.385 -50.615 ;
      RECT -21.485 -51.435 -20.44 -51.335 ;
      RECT -21.485 -48.795 -20.44 -48.695 ;
      RECT -20.965 -49.515 -20.865 -48.695 ;
      RECT -21.485 -49.515 -21.385 -48.695 ;
      RECT -20.965 -38.515 -20.865 -37.695 ;
      RECT -21.485 -38.515 -21.385 -37.695 ;
      RECT -21.485 -38.515 -20.44 -38.415 ;
      RECT -21.485 -35.875 -20.44 -35.775 ;
      RECT -20.965 -36.595 -20.865 -35.775 ;
      RECT -21.485 -36.595 -21.385 -35.775 ;
      RECT -20.965 -25.595 -20.865 -24.775 ;
      RECT -21.485 -25.595 -21.385 -24.775 ;
      RECT -21.485 -25.595 -20.44 -25.495 ;
      RECT -21.485 -22.955 -20.44 -22.855 ;
      RECT -20.965 -23.675 -20.865 -22.855 ;
      RECT -21.485 -23.675 -21.385 -22.855 ;
      RECT -20.965 -12.675 -20.865 -11.855 ;
      RECT -21.485 -12.675 -21.385 -11.855 ;
      RECT -21.485 -12.675 -20.44 -12.575 ;
      RECT -21.485 -10.035 -20.44 -9.935 ;
      RECT -20.965 -10.755 -20.865 -9.935 ;
      RECT -21.485 -10.755 -21.385 -9.935 ;
      RECT -20.965 0.245 -20.865 1.065 ;
      RECT -21.485 0.245 -21.385 1.065 ;
      RECT -21.485 0.245 -20.44 0.345 ;
      RECT -22.785 -100.475 -21.74 -100.375 ;
      RECT -22.265 -101.195 -22.165 -100.375 ;
      RECT -22.785 -101.195 -22.685 -100.375 ;
      RECT -22.265 -90.195 -22.165 -89.375 ;
      RECT -22.785 -90.195 -22.685 -89.375 ;
      RECT -22.785 -90.195 -21.74 -90.095 ;
      RECT -22.785 -87.555 -21.74 -87.455 ;
      RECT -22.265 -88.275 -22.165 -87.455 ;
      RECT -22.785 -88.275 -22.685 -87.455 ;
      RECT -22.265 -77.275 -22.165 -76.455 ;
      RECT -22.785 -77.275 -22.685 -76.455 ;
      RECT -22.785 -77.275 -21.74 -77.175 ;
      RECT -22.785 -74.635 -21.74 -74.535 ;
      RECT -22.265 -75.355 -22.165 -74.535 ;
      RECT -22.785 -75.355 -22.685 -74.535 ;
      RECT -22.265 -64.355 -22.165 -63.535 ;
      RECT -22.785 -64.355 -22.685 -63.535 ;
      RECT -22.785 -64.355 -21.74 -64.255 ;
      RECT -22.785 -61.715 -21.74 -61.615 ;
      RECT -22.265 -62.435 -22.165 -61.615 ;
      RECT -22.785 -62.435 -22.685 -61.615 ;
      RECT -22.265 -51.435 -22.165 -50.615 ;
      RECT -22.785 -51.435 -22.685 -50.615 ;
      RECT -22.785 -51.435 -21.74 -51.335 ;
      RECT -22.785 -48.795 -21.74 -48.695 ;
      RECT -22.265 -49.515 -22.165 -48.695 ;
      RECT -22.785 -49.515 -22.685 -48.695 ;
      RECT -22.265 -38.515 -22.165 -37.695 ;
      RECT -22.785 -38.515 -22.685 -37.695 ;
      RECT -22.785 -38.515 -21.74 -38.415 ;
      RECT -22.785 -35.875 -21.74 -35.775 ;
      RECT -22.265 -36.595 -22.165 -35.775 ;
      RECT -22.785 -36.595 -22.685 -35.775 ;
      RECT -22.265 -25.595 -22.165 -24.775 ;
      RECT -22.785 -25.595 -22.685 -24.775 ;
      RECT -22.785 -25.595 -21.74 -25.495 ;
      RECT -22.785 -22.955 -21.74 -22.855 ;
      RECT -22.265 -23.675 -22.165 -22.855 ;
      RECT -22.785 -23.675 -22.685 -22.855 ;
      RECT -22.265 -12.675 -22.165 -11.855 ;
      RECT -22.785 -12.675 -22.685 -11.855 ;
      RECT -22.785 -12.675 -21.74 -12.575 ;
      RECT -22.785 -10.035 -21.74 -9.935 ;
      RECT -22.265 -10.755 -22.165 -9.935 ;
      RECT -22.785 -10.755 -22.685 -9.935 ;
      RECT -22.265 0.245 -22.165 1.065 ;
      RECT -22.785 0.245 -22.685 1.065 ;
      RECT -22.785 0.245 -21.74 0.345 ;
      RECT -24.085 -100.475 -23.04 -100.375 ;
      RECT -23.565 -101.195 -23.465 -100.375 ;
      RECT -24.085 -101.195 -23.985 -100.375 ;
      RECT -23.565 -90.195 -23.465 -89.375 ;
      RECT -24.085 -90.195 -23.985 -89.375 ;
      RECT -24.085 -90.195 -23.04 -90.095 ;
      RECT -24.085 -87.555 -23.04 -87.455 ;
      RECT -23.565 -88.275 -23.465 -87.455 ;
      RECT -24.085 -88.275 -23.985 -87.455 ;
      RECT -23.565 -77.275 -23.465 -76.455 ;
      RECT -24.085 -77.275 -23.985 -76.455 ;
      RECT -24.085 -77.275 -23.04 -77.175 ;
      RECT -24.085 -74.635 -23.04 -74.535 ;
      RECT -23.565 -75.355 -23.465 -74.535 ;
      RECT -24.085 -75.355 -23.985 -74.535 ;
      RECT -23.565 -64.355 -23.465 -63.535 ;
      RECT -24.085 -64.355 -23.985 -63.535 ;
      RECT -24.085 -64.355 -23.04 -64.255 ;
      RECT -24.085 -61.715 -23.04 -61.615 ;
      RECT -23.565 -62.435 -23.465 -61.615 ;
      RECT -24.085 -62.435 -23.985 -61.615 ;
      RECT -23.565 -51.435 -23.465 -50.615 ;
      RECT -24.085 -51.435 -23.985 -50.615 ;
      RECT -24.085 -51.435 -23.04 -51.335 ;
      RECT -24.085 -48.795 -23.04 -48.695 ;
      RECT -23.565 -49.515 -23.465 -48.695 ;
      RECT -24.085 -49.515 -23.985 -48.695 ;
      RECT -23.565 -38.515 -23.465 -37.695 ;
      RECT -24.085 -38.515 -23.985 -37.695 ;
      RECT -24.085 -38.515 -23.04 -38.415 ;
      RECT -24.085 -35.875 -23.04 -35.775 ;
      RECT -23.565 -36.595 -23.465 -35.775 ;
      RECT -24.085 -36.595 -23.985 -35.775 ;
      RECT -23.565 -25.595 -23.465 -24.775 ;
      RECT -24.085 -25.595 -23.985 -24.775 ;
      RECT -24.085 -25.595 -23.04 -25.495 ;
      RECT -24.085 -22.955 -23.04 -22.855 ;
      RECT -23.565 -23.675 -23.465 -22.855 ;
      RECT -24.085 -23.675 -23.985 -22.855 ;
      RECT -23.565 -12.675 -23.465 -11.855 ;
      RECT -24.085 -12.675 -23.985 -11.855 ;
      RECT -24.085 -12.675 -23.04 -12.575 ;
      RECT -24.085 -10.035 -23.04 -9.935 ;
      RECT -23.565 -10.755 -23.465 -9.935 ;
      RECT -24.085 -10.755 -23.985 -9.935 ;
      RECT -23.565 0.245 -23.465 1.065 ;
      RECT -24.085 0.245 -23.985 1.065 ;
      RECT -24.085 0.245 -23.04 0.345 ;
      RECT -25.385 -100.475 -24.34 -100.375 ;
      RECT -24.865 -101.195 -24.765 -100.375 ;
      RECT -25.385 -101.195 -25.285 -100.375 ;
      RECT -24.865 -90.195 -24.765 -89.375 ;
      RECT -25.385 -90.195 -25.285 -89.375 ;
      RECT -25.385 -90.195 -24.34 -90.095 ;
      RECT -25.385 -87.555 -24.34 -87.455 ;
      RECT -24.865 -88.275 -24.765 -87.455 ;
      RECT -25.385 -88.275 -25.285 -87.455 ;
      RECT -24.865 -77.275 -24.765 -76.455 ;
      RECT -25.385 -77.275 -25.285 -76.455 ;
      RECT -25.385 -77.275 -24.34 -77.175 ;
      RECT -25.385 -74.635 -24.34 -74.535 ;
      RECT -24.865 -75.355 -24.765 -74.535 ;
      RECT -25.385 -75.355 -25.285 -74.535 ;
      RECT -24.865 -64.355 -24.765 -63.535 ;
      RECT -25.385 -64.355 -25.285 -63.535 ;
      RECT -25.385 -64.355 -24.34 -64.255 ;
      RECT -25.385 -61.715 -24.34 -61.615 ;
      RECT -24.865 -62.435 -24.765 -61.615 ;
      RECT -25.385 -62.435 -25.285 -61.615 ;
      RECT -24.865 -51.435 -24.765 -50.615 ;
      RECT -25.385 -51.435 -25.285 -50.615 ;
      RECT -25.385 -51.435 -24.34 -51.335 ;
      RECT -25.385 -48.795 -24.34 -48.695 ;
      RECT -24.865 -49.515 -24.765 -48.695 ;
      RECT -25.385 -49.515 -25.285 -48.695 ;
      RECT -24.865 -38.515 -24.765 -37.695 ;
      RECT -25.385 -38.515 -25.285 -37.695 ;
      RECT -25.385 -38.515 -24.34 -38.415 ;
      RECT -25.385 -35.875 -24.34 -35.775 ;
      RECT -24.865 -36.595 -24.765 -35.775 ;
      RECT -25.385 -36.595 -25.285 -35.775 ;
      RECT -24.865 -25.595 -24.765 -24.775 ;
      RECT -25.385 -25.595 -25.285 -24.775 ;
      RECT -25.385 -25.595 -24.34 -25.495 ;
      RECT -25.385 -22.955 -24.34 -22.855 ;
      RECT -24.865 -23.675 -24.765 -22.855 ;
      RECT -25.385 -23.675 -25.285 -22.855 ;
      RECT -24.865 -12.675 -24.765 -11.855 ;
      RECT -25.385 -12.675 -25.285 -11.855 ;
      RECT -25.385 -12.675 -24.34 -12.575 ;
      RECT -25.385 -10.035 -24.34 -9.935 ;
      RECT -24.865 -10.755 -24.765 -9.935 ;
      RECT -25.385 -10.755 -25.285 -9.935 ;
      RECT -24.865 0.245 -24.765 1.065 ;
      RECT -25.385 0.245 -25.285 1.065 ;
      RECT -25.385 0.245 -24.34 0.345 ;
      RECT -26.685 -100.475 -25.64 -100.375 ;
      RECT -26.165 -101.195 -26.065 -100.375 ;
      RECT -26.685 -101.195 -26.585 -100.375 ;
      RECT -26.165 -90.195 -26.065 -89.375 ;
      RECT -26.685 -90.195 -26.585 -89.375 ;
      RECT -26.685 -90.195 -25.64 -90.095 ;
      RECT -26.685 -87.555 -25.64 -87.455 ;
      RECT -26.165 -88.275 -26.065 -87.455 ;
      RECT -26.685 -88.275 -26.585 -87.455 ;
      RECT -26.165 -77.275 -26.065 -76.455 ;
      RECT -26.685 -77.275 -26.585 -76.455 ;
      RECT -26.685 -77.275 -25.64 -77.175 ;
      RECT -26.685 -74.635 -25.64 -74.535 ;
      RECT -26.165 -75.355 -26.065 -74.535 ;
      RECT -26.685 -75.355 -26.585 -74.535 ;
      RECT -26.165 -64.355 -26.065 -63.535 ;
      RECT -26.685 -64.355 -26.585 -63.535 ;
      RECT -26.685 -64.355 -25.64 -64.255 ;
      RECT -26.685 -61.715 -25.64 -61.615 ;
      RECT -26.165 -62.435 -26.065 -61.615 ;
      RECT -26.685 -62.435 -26.585 -61.615 ;
      RECT -26.165 -51.435 -26.065 -50.615 ;
      RECT -26.685 -51.435 -26.585 -50.615 ;
      RECT -26.685 -51.435 -25.64 -51.335 ;
      RECT -26.685 -48.795 -25.64 -48.695 ;
      RECT -26.165 -49.515 -26.065 -48.695 ;
      RECT -26.685 -49.515 -26.585 -48.695 ;
      RECT -26.165 -38.515 -26.065 -37.695 ;
      RECT -26.685 -38.515 -26.585 -37.695 ;
      RECT -26.685 -38.515 -25.64 -38.415 ;
      RECT -26.685 -35.875 -25.64 -35.775 ;
      RECT -26.165 -36.595 -26.065 -35.775 ;
      RECT -26.685 -36.595 -26.585 -35.775 ;
      RECT -26.165 -25.595 -26.065 -24.775 ;
      RECT -26.685 -25.595 -26.585 -24.775 ;
      RECT -26.685 -25.595 -25.64 -25.495 ;
      RECT -26.685 -22.955 -25.64 -22.855 ;
      RECT -26.165 -23.675 -26.065 -22.855 ;
      RECT -26.685 -23.675 -26.585 -22.855 ;
      RECT -26.165 -12.675 -26.065 -11.855 ;
      RECT -26.685 -12.675 -26.585 -11.855 ;
      RECT -26.685 -12.675 -25.64 -12.575 ;
      RECT -26.685 -10.035 -25.64 -9.935 ;
      RECT -26.165 -10.755 -26.065 -9.935 ;
      RECT -26.685 -10.755 -26.585 -9.935 ;
      RECT -26.165 0.245 -26.065 1.065 ;
      RECT -26.685 0.245 -26.585 1.065 ;
      RECT -26.685 0.245 -25.64 0.345 ;
      RECT -27.985 -100.475 -26.94 -100.375 ;
      RECT -27.465 -101.195 -27.365 -100.375 ;
      RECT -27.985 -101.195 -27.885 -100.375 ;
      RECT -27.465 -90.195 -27.365 -89.375 ;
      RECT -27.985 -90.195 -27.885 -89.375 ;
      RECT -27.985 -90.195 -26.94 -90.095 ;
      RECT -27.985 -87.555 -26.94 -87.455 ;
      RECT -27.465 -88.275 -27.365 -87.455 ;
      RECT -27.985 -88.275 -27.885 -87.455 ;
      RECT -27.465 -77.275 -27.365 -76.455 ;
      RECT -27.985 -77.275 -27.885 -76.455 ;
      RECT -27.985 -77.275 -26.94 -77.175 ;
      RECT -27.985 -74.635 -26.94 -74.535 ;
      RECT -27.465 -75.355 -27.365 -74.535 ;
      RECT -27.985 -75.355 -27.885 -74.535 ;
      RECT -27.465 -64.355 -27.365 -63.535 ;
      RECT -27.985 -64.355 -27.885 -63.535 ;
      RECT -27.985 -64.355 -26.94 -64.255 ;
      RECT -27.985 -61.715 -26.94 -61.615 ;
      RECT -27.465 -62.435 -27.365 -61.615 ;
      RECT -27.985 -62.435 -27.885 -61.615 ;
      RECT -27.465 -51.435 -27.365 -50.615 ;
      RECT -27.985 -51.435 -27.885 -50.615 ;
      RECT -27.985 -51.435 -26.94 -51.335 ;
      RECT -27.985 -48.795 -26.94 -48.695 ;
      RECT -27.465 -49.515 -27.365 -48.695 ;
      RECT -27.985 -49.515 -27.885 -48.695 ;
      RECT -27.465 -38.515 -27.365 -37.695 ;
      RECT -27.985 -38.515 -27.885 -37.695 ;
      RECT -27.985 -38.515 -26.94 -38.415 ;
      RECT -27.985 -35.875 -26.94 -35.775 ;
      RECT -27.465 -36.595 -27.365 -35.775 ;
      RECT -27.985 -36.595 -27.885 -35.775 ;
      RECT -27.465 -25.595 -27.365 -24.775 ;
      RECT -27.985 -25.595 -27.885 -24.775 ;
      RECT -27.985 -25.595 -26.94 -25.495 ;
      RECT -27.985 -22.955 -26.94 -22.855 ;
      RECT -27.465 -23.675 -27.365 -22.855 ;
      RECT -27.985 -23.675 -27.885 -22.855 ;
      RECT -27.465 -12.675 -27.365 -11.855 ;
      RECT -27.985 -12.675 -27.885 -11.855 ;
      RECT -27.985 -12.675 -26.94 -12.575 ;
      RECT -27.985 -10.035 -26.94 -9.935 ;
      RECT -27.465 -10.755 -27.365 -9.935 ;
      RECT -27.985 -10.755 -27.885 -9.935 ;
      RECT -27.465 0.245 -27.365 1.065 ;
      RECT -27.985 0.245 -27.885 1.065 ;
      RECT -27.985 0.245 -26.94 0.345 ;
      RECT -29.285 -100.475 -28.24 -100.375 ;
      RECT -28.765 -101.195 -28.665 -100.375 ;
      RECT -29.285 -101.195 -29.185 -100.375 ;
      RECT -28.765 -90.195 -28.665 -89.375 ;
      RECT -29.285 -90.195 -29.185 -89.375 ;
      RECT -29.285 -90.195 -28.24 -90.095 ;
      RECT -29.285 -87.555 -28.24 -87.455 ;
      RECT -28.765 -88.275 -28.665 -87.455 ;
      RECT -29.285 -88.275 -29.185 -87.455 ;
      RECT -28.765 -77.275 -28.665 -76.455 ;
      RECT -29.285 -77.275 -29.185 -76.455 ;
      RECT -29.285 -77.275 -28.24 -77.175 ;
      RECT -29.285 -74.635 -28.24 -74.535 ;
      RECT -28.765 -75.355 -28.665 -74.535 ;
      RECT -29.285 -75.355 -29.185 -74.535 ;
      RECT -28.765 -64.355 -28.665 -63.535 ;
      RECT -29.285 -64.355 -29.185 -63.535 ;
      RECT -29.285 -64.355 -28.24 -64.255 ;
      RECT -29.285 -61.715 -28.24 -61.615 ;
      RECT -28.765 -62.435 -28.665 -61.615 ;
      RECT -29.285 -62.435 -29.185 -61.615 ;
      RECT -28.765 -51.435 -28.665 -50.615 ;
      RECT -29.285 -51.435 -29.185 -50.615 ;
      RECT -29.285 -51.435 -28.24 -51.335 ;
      RECT -29.285 -48.795 -28.24 -48.695 ;
      RECT -28.765 -49.515 -28.665 -48.695 ;
      RECT -29.285 -49.515 -29.185 -48.695 ;
      RECT -28.765 -38.515 -28.665 -37.695 ;
      RECT -29.285 -38.515 -29.185 -37.695 ;
      RECT -29.285 -38.515 -28.24 -38.415 ;
      RECT -29.285 -35.875 -28.24 -35.775 ;
      RECT -28.765 -36.595 -28.665 -35.775 ;
      RECT -29.285 -36.595 -29.185 -35.775 ;
      RECT -28.765 -25.595 -28.665 -24.775 ;
      RECT -29.285 -25.595 -29.185 -24.775 ;
      RECT -29.285 -25.595 -28.24 -25.495 ;
      RECT -29.285 -22.955 -28.24 -22.855 ;
      RECT -28.765 -23.675 -28.665 -22.855 ;
      RECT -29.285 -23.675 -29.185 -22.855 ;
      RECT -28.765 -12.675 -28.665 -11.855 ;
      RECT -29.285 -12.675 -29.185 -11.855 ;
      RECT -29.285 -12.675 -28.24 -12.575 ;
      RECT -29.285 -10.035 -28.24 -9.935 ;
      RECT -28.765 -10.755 -28.665 -9.935 ;
      RECT -29.285 -10.755 -29.185 -9.935 ;
      RECT -28.765 0.245 -28.665 1.065 ;
      RECT -29.285 0.245 -29.185 1.065 ;
      RECT -29.285 0.245 -28.24 0.345 ;
      RECT -30.585 -100.475 -29.54 -100.375 ;
      RECT -30.065 -101.195 -29.965 -100.375 ;
      RECT -30.585 -101.195 -30.485 -100.375 ;
      RECT -30.065 -90.195 -29.965 -89.375 ;
      RECT -30.585 -90.195 -30.485 -89.375 ;
      RECT -30.585 -90.195 -29.54 -90.095 ;
      RECT -30.585 -87.555 -29.54 -87.455 ;
      RECT -30.065 -88.275 -29.965 -87.455 ;
      RECT -30.585 -88.275 -30.485 -87.455 ;
      RECT -30.065 -77.275 -29.965 -76.455 ;
      RECT -30.585 -77.275 -30.485 -76.455 ;
      RECT -30.585 -77.275 -29.54 -77.175 ;
      RECT -30.585 -74.635 -29.54 -74.535 ;
      RECT -30.065 -75.355 -29.965 -74.535 ;
      RECT -30.585 -75.355 -30.485 -74.535 ;
      RECT -30.065 -64.355 -29.965 -63.535 ;
      RECT -30.585 -64.355 -30.485 -63.535 ;
      RECT -30.585 -64.355 -29.54 -64.255 ;
      RECT -30.585 -61.715 -29.54 -61.615 ;
      RECT -30.065 -62.435 -29.965 -61.615 ;
      RECT -30.585 -62.435 -30.485 -61.615 ;
      RECT -30.065 -51.435 -29.965 -50.615 ;
      RECT -30.585 -51.435 -30.485 -50.615 ;
      RECT -30.585 -51.435 -29.54 -51.335 ;
      RECT -30.585 -48.795 -29.54 -48.695 ;
      RECT -30.065 -49.515 -29.965 -48.695 ;
      RECT -30.585 -49.515 -30.485 -48.695 ;
      RECT -30.065 -38.515 -29.965 -37.695 ;
      RECT -30.585 -38.515 -30.485 -37.695 ;
      RECT -30.585 -38.515 -29.54 -38.415 ;
      RECT -30.585 -35.875 -29.54 -35.775 ;
      RECT -30.065 -36.595 -29.965 -35.775 ;
      RECT -30.585 -36.595 -30.485 -35.775 ;
      RECT -30.065 -25.595 -29.965 -24.775 ;
      RECT -30.585 -25.595 -30.485 -24.775 ;
      RECT -30.585 -25.595 -29.54 -25.495 ;
      RECT -30.585 -22.955 -29.54 -22.855 ;
      RECT -30.065 -23.675 -29.965 -22.855 ;
      RECT -30.585 -23.675 -30.485 -22.855 ;
      RECT -30.065 -12.675 -29.965 -11.855 ;
      RECT -30.585 -12.675 -30.485 -11.855 ;
      RECT -30.585 -12.675 -29.54 -12.575 ;
      RECT -30.585 -10.035 -29.54 -9.935 ;
      RECT -30.065 -10.755 -29.965 -9.935 ;
      RECT -30.585 -10.755 -30.485 -9.935 ;
      RECT -30.065 0.245 -29.965 1.065 ;
      RECT -30.585 0.245 -30.485 1.065 ;
      RECT -30.585 0.245 -29.54 0.345 ;
      RECT -31.885 -100.475 -30.84 -100.375 ;
      RECT -31.365 -101.195 -31.265 -100.375 ;
      RECT -31.885 -101.195 -31.785 -100.375 ;
      RECT -31.365 -90.195 -31.265 -89.375 ;
      RECT -31.885 -90.195 -31.785 -89.375 ;
      RECT -31.885 -90.195 -30.84 -90.095 ;
      RECT -31.885 -87.555 -30.84 -87.455 ;
      RECT -31.365 -88.275 -31.265 -87.455 ;
      RECT -31.885 -88.275 -31.785 -87.455 ;
      RECT -31.365 -77.275 -31.265 -76.455 ;
      RECT -31.885 -77.275 -31.785 -76.455 ;
      RECT -31.885 -77.275 -30.84 -77.175 ;
      RECT -31.885 -74.635 -30.84 -74.535 ;
      RECT -31.365 -75.355 -31.265 -74.535 ;
      RECT -31.885 -75.355 -31.785 -74.535 ;
      RECT -31.365 -64.355 -31.265 -63.535 ;
      RECT -31.885 -64.355 -31.785 -63.535 ;
      RECT -31.885 -64.355 -30.84 -64.255 ;
      RECT -31.885 -61.715 -30.84 -61.615 ;
      RECT -31.365 -62.435 -31.265 -61.615 ;
      RECT -31.885 -62.435 -31.785 -61.615 ;
      RECT -31.365 -51.435 -31.265 -50.615 ;
      RECT -31.885 -51.435 -31.785 -50.615 ;
      RECT -31.885 -51.435 -30.84 -51.335 ;
      RECT -31.885 -48.795 -30.84 -48.695 ;
      RECT -31.365 -49.515 -31.265 -48.695 ;
      RECT -31.885 -49.515 -31.785 -48.695 ;
      RECT -31.365 -38.515 -31.265 -37.695 ;
      RECT -31.885 -38.515 -31.785 -37.695 ;
      RECT -31.885 -38.515 -30.84 -38.415 ;
      RECT -31.885 -35.875 -30.84 -35.775 ;
      RECT -31.365 -36.595 -31.265 -35.775 ;
      RECT -31.885 -36.595 -31.785 -35.775 ;
      RECT -31.365 -25.595 -31.265 -24.775 ;
      RECT -31.885 -25.595 -31.785 -24.775 ;
      RECT -31.885 -25.595 -30.84 -25.495 ;
      RECT -31.885 -22.955 -30.84 -22.855 ;
      RECT -31.365 -23.675 -31.265 -22.855 ;
      RECT -31.885 -23.675 -31.785 -22.855 ;
      RECT -31.365 -12.675 -31.265 -11.855 ;
      RECT -31.885 -12.675 -31.785 -11.855 ;
      RECT -31.885 -12.675 -30.84 -12.575 ;
      RECT -31.885 -10.035 -30.84 -9.935 ;
      RECT -31.365 -10.755 -31.265 -9.935 ;
      RECT -31.885 -10.755 -31.785 -9.935 ;
      RECT -31.365 0.245 -31.265 1.065 ;
      RECT -31.885 0.245 -31.785 1.065 ;
      RECT -31.885 0.245 -30.84 0.345 ;
      RECT -39.505 5.615 -31.945 6.295 ;
      RECT -32.505 4.985 -32.405 6.295 ;
      RECT -33.105 4.985 -33.005 6.295 ;
      RECT -33.705 4.985 -33.605 6.295 ;
      RECT -34.305 4.985 -34.205 6.295 ;
      RECT -34.905 4.985 -34.805 6.295 ;
      RECT -35.505 4.985 -35.405 6.295 ;
      RECT -36.377 -120.365 155.517 -117.645 ;
      RECT -0.605 1.935 154.095 2.035 ;
      RECT 153.55 -101.06 153.65 -100.525 ;
      RECT 153.55 -99.735 153.65 -99.2 ;
      RECT 153.55 -97.83 153.65 -97.295 ;
      RECT 153.55 -96.505 153.65 -95.97 ;
      RECT 153.55 -94.6 153.65 -94.065 ;
      RECT 153.55 -93.275 153.65 -92.74 ;
      RECT 153.55 -91.37 153.65 -90.835 ;
      RECT 153.55 -90.045 153.65 -89.51 ;
      RECT 153.55 -88.14 153.65 -87.605 ;
      RECT 153.55 -86.815 153.65 -86.28 ;
      RECT 153.55 -84.91 153.65 -84.375 ;
      RECT 153.55 -83.585 153.65 -83.05 ;
      RECT 153.55 -81.68 153.65 -81.145 ;
      RECT 153.55 -80.355 153.65 -79.82 ;
      RECT 153.55 -78.45 153.65 -77.915 ;
      RECT 153.55 -77.125 153.65 -76.59 ;
      RECT 153.55 -75.22 153.65 -74.685 ;
      RECT 153.55 -73.895 153.65 -73.36 ;
      RECT 153.55 -71.99 153.65 -71.455 ;
      RECT 153.55 -70.665 153.65 -70.13 ;
      RECT 153.55 -68.76 153.65 -68.225 ;
      RECT 153.55 -67.435 153.65 -66.9 ;
      RECT 153.55 -65.53 153.65 -64.995 ;
      RECT 153.55 -64.205 153.65 -63.67 ;
      RECT 153.55 -62.3 153.65 -61.765 ;
      RECT 153.55 -60.975 153.65 -60.44 ;
      RECT 153.55 -59.07 153.65 -58.535 ;
      RECT 153.55 -57.745 153.65 -57.21 ;
      RECT 153.55 -55.84 153.65 -55.305 ;
      RECT 153.55 -54.515 153.65 -53.98 ;
      RECT 153.55 -52.61 153.65 -52.075 ;
      RECT 153.55 -51.285 153.65 -50.75 ;
      RECT 153.55 -49.38 153.65 -48.845 ;
      RECT 153.55 -48.055 153.65 -47.52 ;
      RECT 153.55 -46.15 153.65 -45.615 ;
      RECT 153.55 -44.825 153.65 -44.29 ;
      RECT 153.55 -42.92 153.65 -42.385 ;
      RECT 153.55 -41.595 153.65 -41.06 ;
      RECT 153.55 -39.69 153.65 -39.155 ;
      RECT 153.55 -38.365 153.65 -37.83 ;
      RECT 153.55 -36.46 153.65 -35.925 ;
      RECT 153.55 -35.135 153.65 -34.6 ;
      RECT 153.55 -33.23 153.65 -32.695 ;
      RECT 153.55 -31.905 153.65 -31.37 ;
      RECT 153.55 -30 153.65 -29.465 ;
      RECT 153.55 -28.675 153.65 -28.14 ;
      RECT 153.55 -26.77 153.65 -26.235 ;
      RECT 153.55 -25.445 153.65 -24.91 ;
      RECT 153.55 -23.54 153.65 -23.005 ;
      RECT 153.55 -22.215 153.65 -21.68 ;
      RECT 153.55 -20.31 153.65 -19.775 ;
      RECT 153.55 -18.985 153.65 -18.45 ;
      RECT 153.55 -17.08 153.65 -16.545 ;
      RECT 153.55 -15.755 153.65 -15.22 ;
      RECT 153.55 -13.85 153.65 -13.315 ;
      RECT 153.55 -12.525 153.65 -11.99 ;
      RECT 153.55 -10.62 153.65 -10.085 ;
      RECT 153.55 -9.295 153.65 -8.76 ;
      RECT 153.55 -7.39 153.65 -6.855 ;
      RECT 153.55 -6.065 153.65 -5.53 ;
      RECT 153.55 -4.16 153.65 -3.625 ;
      RECT 153.55 -2.835 153.65 -2.3 ;
      RECT 153.55 -0.93 153.65 -0.395 ;
      RECT 153.55 0.395 153.65 0.93 ;
      RECT 153.425 -104.945 153.525 -103.985 ;
      RECT 153.05 -100.19 153.4 -100.07 ;
      RECT 153.05 -96.96 153.4 -96.84 ;
      RECT 153.05 -93.73 153.4 -93.61 ;
      RECT 153.05 -90.5 153.4 -90.38 ;
      RECT 153.05 -87.27 153.4 -87.15 ;
      RECT 153.05 -84.04 153.4 -83.92 ;
      RECT 153.05 -80.81 153.4 -80.69 ;
      RECT 153.05 -77.58 153.4 -77.46 ;
      RECT 153.05 -74.35 153.4 -74.23 ;
      RECT 153.05 -71.12 153.4 -71 ;
      RECT 153.05 -67.89 153.4 -67.77 ;
      RECT 153.05 -64.66 153.4 -64.54 ;
      RECT 153.05 -61.43 153.4 -61.31 ;
      RECT 153.05 -58.2 153.4 -58.08 ;
      RECT 153.05 -54.97 153.4 -54.85 ;
      RECT 153.05 -51.74 153.4 -51.62 ;
      RECT 153.05 -48.51 153.4 -48.39 ;
      RECT 153.05 -45.28 153.4 -45.16 ;
      RECT 153.05 -42.05 153.4 -41.93 ;
      RECT 153.05 -38.82 153.4 -38.7 ;
      RECT 153.05 -35.59 153.4 -35.47 ;
      RECT 153.05 -32.36 153.4 -32.24 ;
      RECT 153.05 -29.13 153.4 -29.01 ;
      RECT 153.05 -25.9 153.4 -25.78 ;
      RECT 153.05 -22.67 153.4 -22.55 ;
      RECT 153.05 -19.44 153.4 -19.32 ;
      RECT 153.05 -16.21 153.4 -16.09 ;
      RECT 153.05 -12.98 153.4 -12.86 ;
      RECT 153.05 -9.75 153.4 -9.63 ;
      RECT 153.05 -6.52 153.4 -6.4 ;
      RECT 153.05 -3.29 153.4 -3.17 ;
      RECT 153.05 -0.06 153.4 0.06 ;
      RECT 153.165 -104.945 153.265 -103.985 ;
      RECT 153.165 2.175 153.265 3.135 ;
      RECT 152.875 -112.255 152.975 -111.775 ;
      RECT 152.875 -110.765 152.975 -110.295 ;
      RECT 152.565 -100.19 152.915 -100.07 ;
      RECT 152.565 -96.96 152.915 -96.84 ;
      RECT 152.565 -93.73 152.915 -93.61 ;
      RECT 152.565 -90.5 152.915 -90.38 ;
      RECT 152.565 -87.27 152.915 -87.15 ;
      RECT 152.565 -84.04 152.915 -83.92 ;
      RECT 152.565 -80.81 152.915 -80.69 ;
      RECT 152.565 -77.58 152.915 -77.46 ;
      RECT 152.565 -74.35 152.915 -74.23 ;
      RECT 152.565 -71.12 152.915 -71 ;
      RECT 152.565 -67.89 152.915 -67.77 ;
      RECT 152.565 -64.66 152.915 -64.54 ;
      RECT 152.565 -61.43 152.915 -61.31 ;
      RECT 152.565 -58.2 152.915 -58.08 ;
      RECT 152.565 -54.97 152.915 -54.85 ;
      RECT 152.565 -51.74 152.915 -51.62 ;
      RECT 152.565 -48.51 152.915 -48.39 ;
      RECT 152.565 -45.28 152.915 -45.16 ;
      RECT 152.565 -42.05 152.915 -41.93 ;
      RECT 152.565 -38.82 152.915 -38.7 ;
      RECT 152.565 -35.59 152.915 -35.47 ;
      RECT 152.565 -32.36 152.915 -32.24 ;
      RECT 152.565 -29.13 152.915 -29.01 ;
      RECT 152.565 -25.9 152.915 -25.78 ;
      RECT 152.565 -22.67 152.915 -22.55 ;
      RECT 152.565 -19.44 152.915 -19.32 ;
      RECT 152.565 -16.21 152.915 -16.09 ;
      RECT 152.565 -12.98 152.915 -12.86 ;
      RECT 152.565 -9.75 152.915 -9.63 ;
      RECT 152.565 -6.52 152.915 -6.4 ;
      RECT 152.565 -3.29 152.915 -3.17 ;
      RECT 152.565 -0.06 152.915 0.06 ;
      RECT 152.735 -104.945 152.835 -103.985 ;
      RECT 152.735 2.175 152.835 3.135 ;
      RECT 148.835 -108.655 152.615 -108.535 ;
      RECT 152.475 -104.945 152.575 -103.985 ;
      RECT 152.35 -101.06 152.45 -100.525 ;
      RECT 152.35 -99.735 152.45 -99.2 ;
      RECT 152.35 -97.83 152.45 -97.295 ;
      RECT 152.35 -96.505 152.45 -95.97 ;
      RECT 152.35 -94.6 152.45 -94.065 ;
      RECT 152.35 -93.275 152.45 -92.74 ;
      RECT 152.35 -91.37 152.45 -90.835 ;
      RECT 152.35 -90.045 152.45 -89.51 ;
      RECT 152.35 -88.14 152.45 -87.605 ;
      RECT 152.35 -86.815 152.45 -86.28 ;
      RECT 152.35 -84.91 152.45 -84.375 ;
      RECT 152.35 -83.585 152.45 -83.05 ;
      RECT 152.35 -81.68 152.45 -81.145 ;
      RECT 152.35 -80.355 152.45 -79.82 ;
      RECT 152.35 -78.45 152.45 -77.915 ;
      RECT 152.35 -77.125 152.45 -76.59 ;
      RECT 152.35 -75.22 152.45 -74.685 ;
      RECT 152.35 -73.895 152.45 -73.36 ;
      RECT 152.35 -71.99 152.45 -71.455 ;
      RECT 152.35 -70.665 152.45 -70.13 ;
      RECT 152.35 -68.76 152.45 -68.225 ;
      RECT 152.35 -67.435 152.45 -66.9 ;
      RECT 152.35 -65.53 152.45 -64.995 ;
      RECT 152.35 -64.205 152.45 -63.67 ;
      RECT 152.35 -62.3 152.45 -61.765 ;
      RECT 152.35 -60.975 152.45 -60.44 ;
      RECT 152.35 -59.07 152.45 -58.535 ;
      RECT 152.35 -57.745 152.45 -57.21 ;
      RECT 152.35 -55.84 152.45 -55.305 ;
      RECT 152.35 -54.515 152.45 -53.98 ;
      RECT 152.35 -52.61 152.45 -52.075 ;
      RECT 152.35 -51.285 152.45 -50.75 ;
      RECT 152.35 -49.38 152.45 -48.845 ;
      RECT 152.35 -48.055 152.45 -47.52 ;
      RECT 152.35 -46.15 152.45 -45.615 ;
      RECT 152.35 -44.825 152.45 -44.29 ;
      RECT 152.35 -42.92 152.45 -42.385 ;
      RECT 152.35 -41.595 152.45 -41.06 ;
      RECT 152.35 -39.69 152.45 -39.155 ;
      RECT 152.35 -38.365 152.45 -37.83 ;
      RECT 152.35 -36.46 152.45 -35.925 ;
      RECT 152.35 -35.135 152.45 -34.6 ;
      RECT 152.35 -33.23 152.45 -32.695 ;
      RECT 152.35 -31.905 152.45 -31.37 ;
      RECT 152.35 -30 152.45 -29.465 ;
      RECT 152.35 -28.675 152.45 -28.14 ;
      RECT 152.35 -26.77 152.45 -26.235 ;
      RECT 152.35 -25.445 152.45 -24.91 ;
      RECT 152.35 -23.54 152.45 -23.005 ;
      RECT 152.35 -22.215 152.45 -21.68 ;
      RECT 152.35 -20.31 152.45 -19.775 ;
      RECT 152.35 -18.985 152.45 -18.45 ;
      RECT 152.35 -17.08 152.45 -16.545 ;
      RECT 152.35 -15.755 152.45 -15.22 ;
      RECT 152.35 -13.85 152.45 -13.315 ;
      RECT 152.35 -12.525 152.45 -11.99 ;
      RECT 152.35 -10.62 152.45 -10.085 ;
      RECT 152.35 -9.295 152.45 -8.76 ;
      RECT 152.35 -7.39 152.45 -6.855 ;
      RECT 152.35 -6.065 152.45 -5.53 ;
      RECT 152.35 -4.16 152.45 -3.625 ;
      RECT 152.35 -2.835 152.45 -2.3 ;
      RECT 152.35 -0.93 152.45 -0.395 ;
      RECT 152.35 0.395 152.45 0.93 ;
      RECT 152.285 -110.75 152.405 -110.37 ;
      RECT 152.285 -112.245 152.385 -111.775 ;
      RECT 152.225 -104.945 152.325 -103.985 ;
      RECT 151.85 -100.19 152.2 -100.07 ;
      RECT 151.85 -96.96 152.2 -96.84 ;
      RECT 151.85 -93.73 152.2 -93.61 ;
      RECT 151.85 -90.5 152.2 -90.38 ;
      RECT 151.85 -87.27 152.2 -87.15 ;
      RECT 151.85 -84.04 152.2 -83.92 ;
      RECT 151.85 -80.81 152.2 -80.69 ;
      RECT 151.85 -77.58 152.2 -77.46 ;
      RECT 151.85 -74.35 152.2 -74.23 ;
      RECT 151.85 -71.12 152.2 -71 ;
      RECT 151.85 -67.89 152.2 -67.77 ;
      RECT 151.85 -64.66 152.2 -64.54 ;
      RECT 151.85 -61.43 152.2 -61.31 ;
      RECT 151.85 -58.2 152.2 -58.08 ;
      RECT 151.85 -54.97 152.2 -54.85 ;
      RECT 151.85 -51.74 152.2 -51.62 ;
      RECT 151.85 -48.51 152.2 -48.39 ;
      RECT 151.85 -45.28 152.2 -45.16 ;
      RECT 151.85 -42.05 152.2 -41.93 ;
      RECT 151.85 -38.82 152.2 -38.7 ;
      RECT 151.85 -35.59 152.2 -35.47 ;
      RECT 151.85 -32.36 152.2 -32.24 ;
      RECT 151.85 -29.13 152.2 -29.01 ;
      RECT 151.85 -25.9 152.2 -25.78 ;
      RECT 151.85 -22.67 152.2 -22.55 ;
      RECT 151.85 -19.44 152.2 -19.32 ;
      RECT 151.85 -16.21 152.2 -16.09 ;
      RECT 151.85 -12.98 152.2 -12.86 ;
      RECT 151.85 -9.75 152.2 -9.63 ;
      RECT 151.85 -6.52 152.2 -6.4 ;
      RECT 151.85 -3.29 152.2 -3.17 ;
      RECT 151.85 -0.06 152.2 0.06 ;
      RECT 151.965 -104.945 152.065 -103.985 ;
      RECT 151.965 2.175 152.065 3.135 ;
      RECT 151.695 -109.595 151.83 -109.275 ;
      RECT 151.365 -100.19 151.715 -100.07 ;
      RECT 151.365 -96.96 151.715 -96.84 ;
      RECT 151.365 -93.73 151.715 -93.61 ;
      RECT 151.365 -90.5 151.715 -90.38 ;
      RECT 151.365 -87.27 151.715 -87.15 ;
      RECT 151.365 -84.04 151.715 -83.92 ;
      RECT 151.365 -80.81 151.715 -80.69 ;
      RECT 151.365 -77.58 151.715 -77.46 ;
      RECT 151.365 -74.35 151.715 -74.23 ;
      RECT 151.365 -71.12 151.715 -71 ;
      RECT 151.365 -67.89 151.715 -67.77 ;
      RECT 151.365 -64.66 151.715 -64.54 ;
      RECT 151.365 -61.43 151.715 -61.31 ;
      RECT 151.365 -58.2 151.715 -58.08 ;
      RECT 151.365 -54.97 151.715 -54.85 ;
      RECT 151.365 -51.74 151.715 -51.62 ;
      RECT 151.365 -48.51 151.715 -48.39 ;
      RECT 151.365 -45.28 151.715 -45.16 ;
      RECT 151.365 -42.05 151.715 -41.93 ;
      RECT 151.365 -38.82 151.715 -38.7 ;
      RECT 151.365 -35.59 151.715 -35.47 ;
      RECT 151.365 -32.36 151.715 -32.24 ;
      RECT 151.365 -29.13 151.715 -29.01 ;
      RECT 151.365 -25.9 151.715 -25.78 ;
      RECT 151.365 -22.67 151.715 -22.55 ;
      RECT 151.365 -19.44 151.715 -19.32 ;
      RECT 151.365 -16.21 151.715 -16.09 ;
      RECT 151.365 -12.98 151.715 -12.86 ;
      RECT 151.365 -9.75 151.715 -9.63 ;
      RECT 151.365 -6.52 151.715 -6.4 ;
      RECT 151.365 -3.29 151.715 -3.17 ;
      RECT 151.365 -0.06 151.715 0.06 ;
      RECT 151.535 -104.945 151.635 -103.985 ;
      RECT 151.535 2.175 151.635 3.135 ;
      RECT 151.36 -109.595 151.505 -109.275 ;
      RECT 151.275 -104.945 151.375 -103.985 ;
      RECT 151.15 -101.06 151.25 -100.525 ;
      RECT 151.15 -99.735 151.25 -99.2 ;
      RECT 151.15 -97.83 151.25 -97.295 ;
      RECT 151.15 -96.505 151.25 -95.97 ;
      RECT 151.15 -94.6 151.25 -94.065 ;
      RECT 151.15 -93.275 151.25 -92.74 ;
      RECT 151.15 -91.37 151.25 -90.835 ;
      RECT 151.15 -90.045 151.25 -89.51 ;
      RECT 151.15 -88.14 151.25 -87.605 ;
      RECT 151.15 -86.815 151.25 -86.28 ;
      RECT 151.15 -84.91 151.25 -84.375 ;
      RECT 151.15 -83.585 151.25 -83.05 ;
      RECT 151.15 -81.68 151.25 -81.145 ;
      RECT 151.15 -80.355 151.25 -79.82 ;
      RECT 151.15 -78.45 151.25 -77.915 ;
      RECT 151.15 -77.125 151.25 -76.59 ;
      RECT 151.15 -75.22 151.25 -74.685 ;
      RECT 151.15 -73.895 151.25 -73.36 ;
      RECT 151.15 -71.99 151.25 -71.455 ;
      RECT 151.15 -70.665 151.25 -70.13 ;
      RECT 151.15 -68.76 151.25 -68.225 ;
      RECT 151.15 -67.435 151.25 -66.9 ;
      RECT 151.15 -65.53 151.25 -64.995 ;
      RECT 151.15 -64.205 151.25 -63.67 ;
      RECT 151.15 -62.3 151.25 -61.765 ;
      RECT 151.15 -60.975 151.25 -60.44 ;
      RECT 151.15 -59.07 151.25 -58.535 ;
      RECT 151.15 -57.745 151.25 -57.21 ;
      RECT 151.15 -55.84 151.25 -55.305 ;
      RECT 151.15 -54.515 151.25 -53.98 ;
      RECT 151.15 -52.61 151.25 -52.075 ;
      RECT 151.15 -51.285 151.25 -50.75 ;
      RECT 151.15 -49.38 151.25 -48.845 ;
      RECT 151.15 -48.055 151.25 -47.52 ;
      RECT 151.15 -46.15 151.25 -45.615 ;
      RECT 151.15 -44.825 151.25 -44.29 ;
      RECT 151.15 -42.92 151.25 -42.385 ;
      RECT 151.15 -41.595 151.25 -41.06 ;
      RECT 151.15 -39.69 151.25 -39.155 ;
      RECT 151.15 -38.365 151.25 -37.83 ;
      RECT 151.15 -36.46 151.25 -35.925 ;
      RECT 151.15 -35.135 151.25 -34.6 ;
      RECT 151.15 -33.23 151.25 -32.695 ;
      RECT 151.15 -31.905 151.25 -31.37 ;
      RECT 151.15 -30 151.25 -29.465 ;
      RECT 151.15 -28.675 151.25 -28.14 ;
      RECT 151.15 -26.77 151.25 -26.235 ;
      RECT 151.15 -25.445 151.25 -24.91 ;
      RECT 151.15 -23.54 151.25 -23.005 ;
      RECT 151.15 -22.215 151.25 -21.68 ;
      RECT 151.15 -20.31 151.25 -19.775 ;
      RECT 151.15 -18.985 151.25 -18.45 ;
      RECT 151.15 -17.08 151.25 -16.545 ;
      RECT 151.15 -15.755 151.25 -15.22 ;
      RECT 151.15 -13.85 151.25 -13.315 ;
      RECT 151.15 -12.525 151.25 -11.99 ;
      RECT 151.15 -10.62 151.25 -10.085 ;
      RECT 151.15 -9.295 151.25 -8.76 ;
      RECT 151.15 -7.39 151.25 -6.855 ;
      RECT 151.15 -6.065 151.25 -5.53 ;
      RECT 151.15 -4.16 151.25 -3.625 ;
      RECT 151.15 -2.835 151.25 -2.3 ;
      RECT 151.15 -0.93 151.25 -0.395 ;
      RECT 151.15 0.395 151.25 0.93 ;
      RECT 151.025 -108.175 151.125 -107.215 ;
      RECT 150.65 -100.19 151 -100.07 ;
      RECT 150.65 -96.96 151 -96.84 ;
      RECT 150.65 -93.73 151 -93.61 ;
      RECT 150.65 -90.5 151 -90.38 ;
      RECT 150.65 -87.27 151 -87.15 ;
      RECT 150.65 -84.04 151 -83.92 ;
      RECT 150.65 -80.81 151 -80.69 ;
      RECT 150.65 -77.58 151 -77.46 ;
      RECT 150.65 -74.35 151 -74.23 ;
      RECT 150.65 -71.12 151 -71 ;
      RECT 150.65 -67.89 151 -67.77 ;
      RECT 150.65 -64.66 151 -64.54 ;
      RECT 150.65 -61.43 151 -61.31 ;
      RECT 150.65 -58.2 151 -58.08 ;
      RECT 150.65 -54.97 151 -54.85 ;
      RECT 150.65 -51.74 151 -51.62 ;
      RECT 150.65 -48.51 151 -48.39 ;
      RECT 150.65 -45.28 151 -45.16 ;
      RECT 150.65 -42.05 151 -41.93 ;
      RECT 150.65 -38.82 151 -38.7 ;
      RECT 150.65 -35.59 151 -35.47 ;
      RECT 150.65 -32.36 151 -32.24 ;
      RECT 150.65 -29.13 151 -29.01 ;
      RECT 150.65 -25.9 151 -25.78 ;
      RECT 150.65 -22.67 151 -22.55 ;
      RECT 150.65 -19.44 151 -19.32 ;
      RECT 150.65 -16.21 151 -16.09 ;
      RECT 150.65 -12.98 151 -12.86 ;
      RECT 150.65 -9.75 151 -9.63 ;
      RECT 150.65 -6.52 151 -6.4 ;
      RECT 150.65 -3.29 151 -3.17 ;
      RECT 150.65 -0.06 151 0.06 ;
      RECT 150.855 -112.255 150.955 -111.775 ;
      RECT 150.855 -110.765 150.955 -110.295 ;
      RECT 150.765 -108.175 150.865 -107.215 ;
      RECT 150.765 2.175 150.865 3.135 ;
      RECT 150.165 -100.19 150.515 -100.07 ;
      RECT 150.165 -96.96 150.515 -96.84 ;
      RECT 150.165 -93.73 150.515 -93.61 ;
      RECT 150.165 -90.5 150.515 -90.38 ;
      RECT 150.165 -87.27 150.515 -87.15 ;
      RECT 150.165 -84.04 150.515 -83.92 ;
      RECT 150.165 -80.81 150.515 -80.69 ;
      RECT 150.165 -77.58 150.515 -77.46 ;
      RECT 150.165 -74.35 150.515 -74.23 ;
      RECT 150.165 -71.12 150.515 -71 ;
      RECT 150.165 -67.89 150.515 -67.77 ;
      RECT 150.165 -64.66 150.515 -64.54 ;
      RECT 150.165 -61.43 150.515 -61.31 ;
      RECT 150.165 -58.2 150.515 -58.08 ;
      RECT 150.165 -54.97 150.515 -54.85 ;
      RECT 150.165 -51.74 150.515 -51.62 ;
      RECT 150.165 -48.51 150.515 -48.39 ;
      RECT 150.165 -45.28 150.515 -45.16 ;
      RECT 150.165 -42.05 150.515 -41.93 ;
      RECT 150.165 -38.82 150.515 -38.7 ;
      RECT 150.165 -35.59 150.515 -35.47 ;
      RECT 150.165 -32.36 150.515 -32.24 ;
      RECT 150.165 -29.13 150.515 -29.01 ;
      RECT 150.165 -25.9 150.515 -25.78 ;
      RECT 150.165 -22.67 150.515 -22.55 ;
      RECT 150.165 -19.44 150.515 -19.32 ;
      RECT 150.165 -16.21 150.515 -16.09 ;
      RECT 150.165 -12.98 150.515 -12.86 ;
      RECT 150.165 -9.75 150.515 -9.63 ;
      RECT 150.165 -6.52 150.515 -6.4 ;
      RECT 150.165 -3.29 150.515 -3.17 ;
      RECT 150.165 -0.06 150.515 0.06 ;
      RECT 150.335 -108.175 150.435 -107.215 ;
      RECT 150.335 2.175 150.435 3.135 ;
      RECT 150.23 -110.765 150.4 -110.385 ;
      RECT 150.265 -112.245 150.365 -111.775 ;
      RECT 150.075 -108.175 150.175 -107.215 ;
      RECT 149.95 -101.06 150.05 -100.525 ;
      RECT 149.95 -99.735 150.05 -99.2 ;
      RECT 149.95 -97.83 150.05 -97.295 ;
      RECT 149.95 -96.505 150.05 -95.97 ;
      RECT 149.95 -94.6 150.05 -94.065 ;
      RECT 149.95 -93.275 150.05 -92.74 ;
      RECT 149.95 -91.37 150.05 -90.835 ;
      RECT 149.95 -90.045 150.05 -89.51 ;
      RECT 149.95 -88.14 150.05 -87.605 ;
      RECT 149.95 -86.815 150.05 -86.28 ;
      RECT 149.95 -84.91 150.05 -84.375 ;
      RECT 149.95 -83.585 150.05 -83.05 ;
      RECT 149.95 -81.68 150.05 -81.145 ;
      RECT 149.95 -80.355 150.05 -79.82 ;
      RECT 149.95 -78.45 150.05 -77.915 ;
      RECT 149.95 -77.125 150.05 -76.59 ;
      RECT 149.95 -75.22 150.05 -74.685 ;
      RECT 149.95 -73.895 150.05 -73.36 ;
      RECT 149.95 -71.99 150.05 -71.455 ;
      RECT 149.95 -70.665 150.05 -70.13 ;
      RECT 149.95 -68.76 150.05 -68.225 ;
      RECT 149.95 -67.435 150.05 -66.9 ;
      RECT 149.95 -65.53 150.05 -64.995 ;
      RECT 149.95 -64.205 150.05 -63.67 ;
      RECT 149.95 -62.3 150.05 -61.765 ;
      RECT 149.95 -60.975 150.05 -60.44 ;
      RECT 149.95 -59.07 150.05 -58.535 ;
      RECT 149.95 -57.745 150.05 -57.21 ;
      RECT 149.95 -55.84 150.05 -55.305 ;
      RECT 149.95 -54.515 150.05 -53.98 ;
      RECT 149.95 -52.61 150.05 -52.075 ;
      RECT 149.95 -51.285 150.05 -50.75 ;
      RECT 149.95 -49.38 150.05 -48.845 ;
      RECT 149.95 -48.055 150.05 -47.52 ;
      RECT 149.95 -46.15 150.05 -45.615 ;
      RECT 149.95 -44.825 150.05 -44.29 ;
      RECT 149.95 -42.92 150.05 -42.385 ;
      RECT 149.95 -41.595 150.05 -41.06 ;
      RECT 149.95 -39.69 150.05 -39.155 ;
      RECT 149.95 -38.365 150.05 -37.83 ;
      RECT 149.95 -36.46 150.05 -35.925 ;
      RECT 149.95 -35.135 150.05 -34.6 ;
      RECT 149.95 -33.23 150.05 -32.695 ;
      RECT 149.95 -31.905 150.05 -31.37 ;
      RECT 149.95 -30 150.05 -29.465 ;
      RECT 149.95 -28.675 150.05 -28.14 ;
      RECT 149.95 -26.77 150.05 -26.235 ;
      RECT 149.95 -25.445 150.05 -24.91 ;
      RECT 149.95 -23.54 150.05 -23.005 ;
      RECT 149.95 -22.215 150.05 -21.68 ;
      RECT 149.95 -20.31 150.05 -19.775 ;
      RECT 149.95 -18.985 150.05 -18.45 ;
      RECT 149.95 -17.08 150.05 -16.545 ;
      RECT 149.95 -15.755 150.05 -15.22 ;
      RECT 149.95 -13.85 150.05 -13.315 ;
      RECT 149.95 -12.525 150.05 -11.99 ;
      RECT 149.95 -10.62 150.05 -10.085 ;
      RECT 149.95 -9.295 150.05 -8.76 ;
      RECT 149.95 -7.39 150.05 -6.855 ;
      RECT 149.95 -6.065 150.05 -5.53 ;
      RECT 149.95 -4.16 150.05 -3.625 ;
      RECT 149.95 -2.835 150.05 -2.3 ;
      RECT 149.95 -0.93 150.05 -0.395 ;
      RECT 149.95 0.395 150.05 0.93 ;
      RECT 149.825 -108.175 149.925 -107.215 ;
      RECT 149.45 -100.19 149.8 -100.07 ;
      RECT 149.45 -96.96 149.8 -96.84 ;
      RECT 149.45 -93.73 149.8 -93.61 ;
      RECT 149.45 -90.5 149.8 -90.38 ;
      RECT 149.45 -87.27 149.8 -87.15 ;
      RECT 149.45 -84.04 149.8 -83.92 ;
      RECT 149.45 -80.81 149.8 -80.69 ;
      RECT 149.45 -77.58 149.8 -77.46 ;
      RECT 149.45 -74.35 149.8 -74.23 ;
      RECT 149.45 -71.12 149.8 -71 ;
      RECT 149.45 -67.89 149.8 -67.77 ;
      RECT 149.45 -64.66 149.8 -64.54 ;
      RECT 149.45 -61.43 149.8 -61.31 ;
      RECT 149.45 -58.2 149.8 -58.08 ;
      RECT 149.45 -54.97 149.8 -54.85 ;
      RECT 149.45 -51.74 149.8 -51.62 ;
      RECT 149.45 -48.51 149.8 -48.39 ;
      RECT 149.45 -45.28 149.8 -45.16 ;
      RECT 149.45 -42.05 149.8 -41.93 ;
      RECT 149.45 -38.82 149.8 -38.7 ;
      RECT 149.45 -35.59 149.8 -35.47 ;
      RECT 149.45 -32.36 149.8 -32.24 ;
      RECT 149.45 -29.13 149.8 -29.01 ;
      RECT 149.45 -25.9 149.8 -25.78 ;
      RECT 149.45 -22.67 149.8 -22.55 ;
      RECT 149.45 -19.44 149.8 -19.32 ;
      RECT 149.45 -16.21 149.8 -16.09 ;
      RECT 149.45 -12.98 149.8 -12.86 ;
      RECT 149.45 -9.75 149.8 -9.63 ;
      RECT 149.45 -6.52 149.8 -6.4 ;
      RECT 149.45 -3.29 149.8 -3.17 ;
      RECT 149.45 -0.06 149.8 0.06 ;
      RECT 149.565 -108.175 149.665 -107.215 ;
      RECT 149.565 2.175 149.665 3.135 ;
      RECT 149.465 -113.555 149.565 -113.085 ;
      RECT 148.965 -100.19 149.315 -100.07 ;
      RECT 148.965 -96.96 149.315 -96.84 ;
      RECT 148.965 -93.73 149.315 -93.61 ;
      RECT 148.965 -90.5 149.315 -90.38 ;
      RECT 148.965 -87.27 149.315 -87.15 ;
      RECT 148.965 -84.04 149.315 -83.92 ;
      RECT 148.965 -80.81 149.315 -80.69 ;
      RECT 148.965 -77.58 149.315 -77.46 ;
      RECT 148.965 -74.35 149.315 -74.23 ;
      RECT 148.965 -71.12 149.315 -71 ;
      RECT 148.965 -67.89 149.315 -67.77 ;
      RECT 148.965 -64.66 149.315 -64.54 ;
      RECT 148.965 -61.43 149.315 -61.31 ;
      RECT 148.965 -58.2 149.315 -58.08 ;
      RECT 148.965 -54.97 149.315 -54.85 ;
      RECT 148.965 -51.74 149.315 -51.62 ;
      RECT 148.965 -48.51 149.315 -48.39 ;
      RECT 148.965 -45.28 149.315 -45.16 ;
      RECT 148.965 -42.05 149.315 -41.93 ;
      RECT 148.965 -38.82 149.315 -38.7 ;
      RECT 148.965 -35.59 149.315 -35.47 ;
      RECT 148.965 -32.36 149.315 -32.24 ;
      RECT 148.965 -29.13 149.315 -29.01 ;
      RECT 148.965 -25.9 149.315 -25.78 ;
      RECT 148.965 -22.67 149.315 -22.55 ;
      RECT 148.965 -19.44 149.315 -19.32 ;
      RECT 148.965 -16.21 149.315 -16.09 ;
      RECT 148.965 -12.98 149.315 -12.86 ;
      RECT 148.965 -9.75 149.315 -9.63 ;
      RECT 148.965 -6.52 149.315 -6.4 ;
      RECT 148.965 -3.29 149.315 -3.17 ;
      RECT 148.965 -0.06 149.315 0.06 ;
      RECT 149.1 -110.735 149.25 -110.445 ;
      RECT 149.135 -108.175 149.235 -107.215 ;
      RECT 149.135 2.175 149.235 3.135 ;
      RECT 149.115 -112.19 149.215 -111.65 ;
      RECT 148.875 -113.555 148.975 -113.085 ;
      RECT 148.875 -108.175 148.975 -107.215 ;
      RECT 148.75 -101.06 148.85 -100.525 ;
      RECT 148.75 -99.735 148.85 -99.2 ;
      RECT 148.75 -97.83 148.85 -97.295 ;
      RECT 148.75 -96.505 148.85 -95.97 ;
      RECT 148.75 -94.6 148.85 -94.065 ;
      RECT 148.75 -93.275 148.85 -92.74 ;
      RECT 148.75 -91.37 148.85 -90.835 ;
      RECT 148.75 -90.045 148.85 -89.51 ;
      RECT 148.75 -88.14 148.85 -87.605 ;
      RECT 148.75 -86.815 148.85 -86.28 ;
      RECT 148.75 -84.91 148.85 -84.375 ;
      RECT 148.75 -83.585 148.85 -83.05 ;
      RECT 148.75 -81.68 148.85 -81.145 ;
      RECT 148.75 -80.355 148.85 -79.82 ;
      RECT 148.75 -78.45 148.85 -77.915 ;
      RECT 148.75 -77.125 148.85 -76.59 ;
      RECT 148.75 -75.22 148.85 -74.685 ;
      RECT 148.75 -73.895 148.85 -73.36 ;
      RECT 148.75 -71.99 148.85 -71.455 ;
      RECT 148.75 -70.665 148.85 -70.13 ;
      RECT 148.75 -68.76 148.85 -68.225 ;
      RECT 148.75 -67.435 148.85 -66.9 ;
      RECT 148.75 -65.53 148.85 -64.995 ;
      RECT 148.75 -64.205 148.85 -63.67 ;
      RECT 148.75 -62.3 148.85 -61.765 ;
      RECT 148.75 -60.975 148.85 -60.44 ;
      RECT 148.75 -59.07 148.85 -58.535 ;
      RECT 148.75 -57.745 148.85 -57.21 ;
      RECT 148.75 -55.84 148.85 -55.305 ;
      RECT 148.75 -54.515 148.85 -53.98 ;
      RECT 148.75 -52.61 148.85 -52.075 ;
      RECT 148.75 -51.285 148.85 -50.75 ;
      RECT 148.75 -49.38 148.85 -48.845 ;
      RECT 148.75 -48.055 148.85 -47.52 ;
      RECT 148.75 -46.15 148.85 -45.615 ;
      RECT 148.75 -44.825 148.85 -44.29 ;
      RECT 148.75 -42.92 148.85 -42.385 ;
      RECT 148.75 -41.595 148.85 -41.06 ;
      RECT 148.75 -39.69 148.85 -39.155 ;
      RECT 148.75 -38.365 148.85 -37.83 ;
      RECT 148.75 -36.46 148.85 -35.925 ;
      RECT 148.75 -35.135 148.85 -34.6 ;
      RECT 148.75 -33.23 148.85 -32.695 ;
      RECT 148.75 -31.905 148.85 -31.37 ;
      RECT 148.75 -30 148.85 -29.465 ;
      RECT 148.75 -28.675 148.85 -28.14 ;
      RECT 148.75 -26.77 148.85 -26.235 ;
      RECT 148.75 -25.445 148.85 -24.91 ;
      RECT 148.75 -23.54 148.85 -23.005 ;
      RECT 148.75 -22.215 148.85 -21.68 ;
      RECT 148.75 -20.31 148.85 -19.775 ;
      RECT 148.75 -18.985 148.85 -18.45 ;
      RECT 148.75 -17.08 148.85 -16.545 ;
      RECT 148.75 -15.755 148.85 -15.22 ;
      RECT 148.75 -13.85 148.85 -13.315 ;
      RECT 148.75 -12.525 148.85 -11.99 ;
      RECT 148.75 -10.62 148.85 -10.085 ;
      RECT 148.75 -9.295 148.85 -8.76 ;
      RECT 148.75 -7.39 148.85 -6.855 ;
      RECT 148.75 -6.065 148.85 -5.53 ;
      RECT 148.75 -4.16 148.85 -3.625 ;
      RECT 148.75 -2.835 148.85 -2.3 ;
      RECT 148.75 -0.93 148.85 -0.395 ;
      RECT 148.75 0.395 148.85 0.93 ;
      RECT 148.625 -104.945 148.725 -103.985 ;
      RECT 148.25 -100.19 148.6 -100.07 ;
      RECT 148.25 -96.96 148.6 -96.84 ;
      RECT 148.25 -93.73 148.6 -93.61 ;
      RECT 148.25 -90.5 148.6 -90.38 ;
      RECT 148.25 -87.27 148.6 -87.15 ;
      RECT 148.25 -84.04 148.6 -83.92 ;
      RECT 148.25 -80.81 148.6 -80.69 ;
      RECT 148.25 -77.58 148.6 -77.46 ;
      RECT 148.25 -74.35 148.6 -74.23 ;
      RECT 148.25 -71.12 148.6 -71 ;
      RECT 148.25 -67.89 148.6 -67.77 ;
      RECT 148.25 -64.66 148.6 -64.54 ;
      RECT 148.25 -61.43 148.6 -61.31 ;
      RECT 148.25 -58.2 148.6 -58.08 ;
      RECT 148.25 -54.97 148.6 -54.85 ;
      RECT 148.25 -51.74 148.6 -51.62 ;
      RECT 148.25 -48.51 148.6 -48.39 ;
      RECT 148.25 -45.28 148.6 -45.16 ;
      RECT 148.25 -42.05 148.6 -41.93 ;
      RECT 148.25 -38.82 148.6 -38.7 ;
      RECT 148.25 -35.59 148.6 -35.47 ;
      RECT 148.25 -32.36 148.6 -32.24 ;
      RECT 148.25 -29.13 148.6 -29.01 ;
      RECT 148.25 -25.9 148.6 -25.78 ;
      RECT 148.25 -22.67 148.6 -22.55 ;
      RECT 148.25 -19.44 148.6 -19.32 ;
      RECT 148.25 -16.21 148.6 -16.09 ;
      RECT 148.25 -12.98 148.6 -12.86 ;
      RECT 148.25 -9.75 148.6 -9.63 ;
      RECT 148.25 -6.52 148.6 -6.4 ;
      RECT 148.25 -3.29 148.6 -3.17 ;
      RECT 148.25 -0.06 148.6 0.06 ;
      RECT 148.365 -104.945 148.465 -103.985 ;
      RECT 148.365 2.175 148.465 3.135 ;
      RECT 148.075 -112.255 148.175 -111.775 ;
      RECT 148.075 -110.765 148.175 -110.295 ;
      RECT 147.765 -100.19 148.115 -100.07 ;
      RECT 147.765 -96.96 148.115 -96.84 ;
      RECT 147.765 -93.73 148.115 -93.61 ;
      RECT 147.765 -90.5 148.115 -90.38 ;
      RECT 147.765 -87.27 148.115 -87.15 ;
      RECT 147.765 -84.04 148.115 -83.92 ;
      RECT 147.765 -80.81 148.115 -80.69 ;
      RECT 147.765 -77.58 148.115 -77.46 ;
      RECT 147.765 -74.35 148.115 -74.23 ;
      RECT 147.765 -71.12 148.115 -71 ;
      RECT 147.765 -67.89 148.115 -67.77 ;
      RECT 147.765 -64.66 148.115 -64.54 ;
      RECT 147.765 -61.43 148.115 -61.31 ;
      RECT 147.765 -58.2 148.115 -58.08 ;
      RECT 147.765 -54.97 148.115 -54.85 ;
      RECT 147.765 -51.74 148.115 -51.62 ;
      RECT 147.765 -48.51 148.115 -48.39 ;
      RECT 147.765 -45.28 148.115 -45.16 ;
      RECT 147.765 -42.05 148.115 -41.93 ;
      RECT 147.765 -38.82 148.115 -38.7 ;
      RECT 147.765 -35.59 148.115 -35.47 ;
      RECT 147.765 -32.36 148.115 -32.24 ;
      RECT 147.765 -29.13 148.115 -29.01 ;
      RECT 147.765 -25.9 148.115 -25.78 ;
      RECT 147.765 -22.67 148.115 -22.55 ;
      RECT 147.765 -19.44 148.115 -19.32 ;
      RECT 147.765 -16.21 148.115 -16.09 ;
      RECT 147.765 -12.98 148.115 -12.86 ;
      RECT 147.765 -9.75 148.115 -9.63 ;
      RECT 147.765 -6.52 148.115 -6.4 ;
      RECT 147.765 -3.29 148.115 -3.17 ;
      RECT 147.765 -0.06 148.115 0.06 ;
      RECT 147.935 -104.945 148.035 -103.985 ;
      RECT 147.935 2.175 148.035 3.135 ;
      RECT 144.035 -108.655 147.815 -108.535 ;
      RECT 147.675 -104.945 147.775 -103.985 ;
      RECT 147.55 -101.06 147.65 -100.525 ;
      RECT 147.55 -99.735 147.65 -99.2 ;
      RECT 147.55 -97.83 147.65 -97.295 ;
      RECT 147.55 -96.505 147.65 -95.97 ;
      RECT 147.55 -94.6 147.65 -94.065 ;
      RECT 147.55 -93.275 147.65 -92.74 ;
      RECT 147.55 -91.37 147.65 -90.835 ;
      RECT 147.55 -90.045 147.65 -89.51 ;
      RECT 147.55 -88.14 147.65 -87.605 ;
      RECT 147.55 -86.815 147.65 -86.28 ;
      RECT 147.55 -84.91 147.65 -84.375 ;
      RECT 147.55 -83.585 147.65 -83.05 ;
      RECT 147.55 -81.68 147.65 -81.145 ;
      RECT 147.55 -80.355 147.65 -79.82 ;
      RECT 147.55 -78.45 147.65 -77.915 ;
      RECT 147.55 -77.125 147.65 -76.59 ;
      RECT 147.55 -75.22 147.65 -74.685 ;
      RECT 147.55 -73.895 147.65 -73.36 ;
      RECT 147.55 -71.99 147.65 -71.455 ;
      RECT 147.55 -70.665 147.65 -70.13 ;
      RECT 147.55 -68.76 147.65 -68.225 ;
      RECT 147.55 -67.435 147.65 -66.9 ;
      RECT 147.55 -65.53 147.65 -64.995 ;
      RECT 147.55 -64.205 147.65 -63.67 ;
      RECT 147.55 -62.3 147.65 -61.765 ;
      RECT 147.55 -60.975 147.65 -60.44 ;
      RECT 147.55 -59.07 147.65 -58.535 ;
      RECT 147.55 -57.745 147.65 -57.21 ;
      RECT 147.55 -55.84 147.65 -55.305 ;
      RECT 147.55 -54.515 147.65 -53.98 ;
      RECT 147.55 -52.61 147.65 -52.075 ;
      RECT 147.55 -51.285 147.65 -50.75 ;
      RECT 147.55 -49.38 147.65 -48.845 ;
      RECT 147.55 -48.055 147.65 -47.52 ;
      RECT 147.55 -46.15 147.65 -45.615 ;
      RECT 147.55 -44.825 147.65 -44.29 ;
      RECT 147.55 -42.92 147.65 -42.385 ;
      RECT 147.55 -41.595 147.65 -41.06 ;
      RECT 147.55 -39.69 147.65 -39.155 ;
      RECT 147.55 -38.365 147.65 -37.83 ;
      RECT 147.55 -36.46 147.65 -35.925 ;
      RECT 147.55 -35.135 147.65 -34.6 ;
      RECT 147.55 -33.23 147.65 -32.695 ;
      RECT 147.55 -31.905 147.65 -31.37 ;
      RECT 147.55 -30 147.65 -29.465 ;
      RECT 147.55 -28.675 147.65 -28.14 ;
      RECT 147.55 -26.77 147.65 -26.235 ;
      RECT 147.55 -25.445 147.65 -24.91 ;
      RECT 147.55 -23.54 147.65 -23.005 ;
      RECT 147.55 -22.215 147.65 -21.68 ;
      RECT 147.55 -20.31 147.65 -19.775 ;
      RECT 147.55 -18.985 147.65 -18.45 ;
      RECT 147.55 -17.08 147.65 -16.545 ;
      RECT 147.55 -15.755 147.65 -15.22 ;
      RECT 147.55 -13.85 147.65 -13.315 ;
      RECT 147.55 -12.525 147.65 -11.99 ;
      RECT 147.55 -10.62 147.65 -10.085 ;
      RECT 147.55 -9.295 147.65 -8.76 ;
      RECT 147.55 -7.39 147.65 -6.855 ;
      RECT 147.55 -6.065 147.65 -5.53 ;
      RECT 147.55 -4.16 147.65 -3.625 ;
      RECT 147.55 -2.835 147.65 -2.3 ;
      RECT 147.55 -0.93 147.65 -0.395 ;
      RECT 147.55 0.395 147.65 0.93 ;
      RECT 147.485 -110.75 147.605 -110.37 ;
      RECT 147.485 -112.245 147.585 -111.775 ;
      RECT 147.425 -104.945 147.525 -103.985 ;
      RECT 147.05 -100.19 147.4 -100.07 ;
      RECT 147.05 -96.96 147.4 -96.84 ;
      RECT 147.05 -93.73 147.4 -93.61 ;
      RECT 147.05 -90.5 147.4 -90.38 ;
      RECT 147.05 -87.27 147.4 -87.15 ;
      RECT 147.05 -84.04 147.4 -83.92 ;
      RECT 147.05 -80.81 147.4 -80.69 ;
      RECT 147.05 -77.58 147.4 -77.46 ;
      RECT 147.05 -74.35 147.4 -74.23 ;
      RECT 147.05 -71.12 147.4 -71 ;
      RECT 147.05 -67.89 147.4 -67.77 ;
      RECT 147.05 -64.66 147.4 -64.54 ;
      RECT 147.05 -61.43 147.4 -61.31 ;
      RECT 147.05 -58.2 147.4 -58.08 ;
      RECT 147.05 -54.97 147.4 -54.85 ;
      RECT 147.05 -51.74 147.4 -51.62 ;
      RECT 147.05 -48.51 147.4 -48.39 ;
      RECT 147.05 -45.28 147.4 -45.16 ;
      RECT 147.05 -42.05 147.4 -41.93 ;
      RECT 147.05 -38.82 147.4 -38.7 ;
      RECT 147.05 -35.59 147.4 -35.47 ;
      RECT 147.05 -32.36 147.4 -32.24 ;
      RECT 147.05 -29.13 147.4 -29.01 ;
      RECT 147.05 -25.9 147.4 -25.78 ;
      RECT 147.05 -22.67 147.4 -22.55 ;
      RECT 147.05 -19.44 147.4 -19.32 ;
      RECT 147.05 -16.21 147.4 -16.09 ;
      RECT 147.05 -12.98 147.4 -12.86 ;
      RECT 147.05 -9.75 147.4 -9.63 ;
      RECT 147.05 -6.52 147.4 -6.4 ;
      RECT 147.05 -3.29 147.4 -3.17 ;
      RECT 147.05 -0.06 147.4 0.06 ;
      RECT 147.165 -104.945 147.265 -103.985 ;
      RECT 147.165 2.175 147.265 3.135 ;
      RECT 146.895 -109.595 147.03 -109.275 ;
      RECT 146.565 -100.19 146.915 -100.07 ;
      RECT 146.565 -96.96 146.915 -96.84 ;
      RECT 146.565 -93.73 146.915 -93.61 ;
      RECT 146.565 -90.5 146.915 -90.38 ;
      RECT 146.565 -87.27 146.915 -87.15 ;
      RECT 146.565 -84.04 146.915 -83.92 ;
      RECT 146.565 -80.81 146.915 -80.69 ;
      RECT 146.565 -77.58 146.915 -77.46 ;
      RECT 146.565 -74.35 146.915 -74.23 ;
      RECT 146.565 -71.12 146.915 -71 ;
      RECT 146.565 -67.89 146.915 -67.77 ;
      RECT 146.565 -64.66 146.915 -64.54 ;
      RECT 146.565 -61.43 146.915 -61.31 ;
      RECT 146.565 -58.2 146.915 -58.08 ;
      RECT 146.565 -54.97 146.915 -54.85 ;
      RECT 146.565 -51.74 146.915 -51.62 ;
      RECT 146.565 -48.51 146.915 -48.39 ;
      RECT 146.565 -45.28 146.915 -45.16 ;
      RECT 146.565 -42.05 146.915 -41.93 ;
      RECT 146.565 -38.82 146.915 -38.7 ;
      RECT 146.565 -35.59 146.915 -35.47 ;
      RECT 146.565 -32.36 146.915 -32.24 ;
      RECT 146.565 -29.13 146.915 -29.01 ;
      RECT 146.565 -25.9 146.915 -25.78 ;
      RECT 146.565 -22.67 146.915 -22.55 ;
      RECT 146.565 -19.44 146.915 -19.32 ;
      RECT 146.565 -16.21 146.915 -16.09 ;
      RECT 146.565 -12.98 146.915 -12.86 ;
      RECT 146.565 -9.75 146.915 -9.63 ;
      RECT 146.565 -6.52 146.915 -6.4 ;
      RECT 146.565 -3.29 146.915 -3.17 ;
      RECT 146.565 -0.06 146.915 0.06 ;
      RECT 146.735 -104.945 146.835 -103.985 ;
      RECT 146.735 2.175 146.835 3.135 ;
      RECT 146.56 -109.595 146.705 -109.275 ;
      RECT 146.475 -104.945 146.575 -103.985 ;
      RECT 146.35 -101.06 146.45 -100.525 ;
      RECT 146.35 -99.735 146.45 -99.2 ;
      RECT 146.35 -97.83 146.45 -97.295 ;
      RECT 146.35 -96.505 146.45 -95.97 ;
      RECT 146.35 -94.6 146.45 -94.065 ;
      RECT 146.35 -93.275 146.45 -92.74 ;
      RECT 146.35 -91.37 146.45 -90.835 ;
      RECT 146.35 -90.045 146.45 -89.51 ;
      RECT 146.35 -88.14 146.45 -87.605 ;
      RECT 146.35 -86.815 146.45 -86.28 ;
      RECT 146.35 -84.91 146.45 -84.375 ;
      RECT 146.35 -83.585 146.45 -83.05 ;
      RECT 146.35 -81.68 146.45 -81.145 ;
      RECT 146.35 -80.355 146.45 -79.82 ;
      RECT 146.35 -78.45 146.45 -77.915 ;
      RECT 146.35 -77.125 146.45 -76.59 ;
      RECT 146.35 -75.22 146.45 -74.685 ;
      RECT 146.35 -73.895 146.45 -73.36 ;
      RECT 146.35 -71.99 146.45 -71.455 ;
      RECT 146.35 -70.665 146.45 -70.13 ;
      RECT 146.35 -68.76 146.45 -68.225 ;
      RECT 146.35 -67.435 146.45 -66.9 ;
      RECT 146.35 -65.53 146.45 -64.995 ;
      RECT 146.35 -64.205 146.45 -63.67 ;
      RECT 146.35 -62.3 146.45 -61.765 ;
      RECT 146.35 -60.975 146.45 -60.44 ;
      RECT 146.35 -59.07 146.45 -58.535 ;
      RECT 146.35 -57.745 146.45 -57.21 ;
      RECT 146.35 -55.84 146.45 -55.305 ;
      RECT 146.35 -54.515 146.45 -53.98 ;
      RECT 146.35 -52.61 146.45 -52.075 ;
      RECT 146.35 -51.285 146.45 -50.75 ;
      RECT 146.35 -49.38 146.45 -48.845 ;
      RECT 146.35 -48.055 146.45 -47.52 ;
      RECT 146.35 -46.15 146.45 -45.615 ;
      RECT 146.35 -44.825 146.45 -44.29 ;
      RECT 146.35 -42.92 146.45 -42.385 ;
      RECT 146.35 -41.595 146.45 -41.06 ;
      RECT 146.35 -39.69 146.45 -39.155 ;
      RECT 146.35 -38.365 146.45 -37.83 ;
      RECT 146.35 -36.46 146.45 -35.925 ;
      RECT 146.35 -35.135 146.45 -34.6 ;
      RECT 146.35 -33.23 146.45 -32.695 ;
      RECT 146.35 -31.905 146.45 -31.37 ;
      RECT 146.35 -30 146.45 -29.465 ;
      RECT 146.35 -28.675 146.45 -28.14 ;
      RECT 146.35 -26.77 146.45 -26.235 ;
      RECT 146.35 -25.445 146.45 -24.91 ;
      RECT 146.35 -23.54 146.45 -23.005 ;
      RECT 146.35 -22.215 146.45 -21.68 ;
      RECT 146.35 -20.31 146.45 -19.775 ;
      RECT 146.35 -18.985 146.45 -18.45 ;
      RECT 146.35 -17.08 146.45 -16.545 ;
      RECT 146.35 -15.755 146.45 -15.22 ;
      RECT 146.35 -13.85 146.45 -13.315 ;
      RECT 146.35 -12.525 146.45 -11.99 ;
      RECT 146.35 -10.62 146.45 -10.085 ;
      RECT 146.35 -9.295 146.45 -8.76 ;
      RECT 146.35 -7.39 146.45 -6.855 ;
      RECT 146.35 -6.065 146.45 -5.53 ;
      RECT 146.35 -4.16 146.45 -3.625 ;
      RECT 146.35 -2.835 146.45 -2.3 ;
      RECT 146.35 -0.93 146.45 -0.395 ;
      RECT 146.35 0.395 146.45 0.93 ;
      RECT 146.225 -108.175 146.325 -107.215 ;
      RECT 145.85 -100.19 146.2 -100.07 ;
      RECT 145.85 -96.96 146.2 -96.84 ;
      RECT 145.85 -93.73 146.2 -93.61 ;
      RECT 145.85 -90.5 146.2 -90.38 ;
      RECT 145.85 -87.27 146.2 -87.15 ;
      RECT 145.85 -84.04 146.2 -83.92 ;
      RECT 145.85 -80.81 146.2 -80.69 ;
      RECT 145.85 -77.58 146.2 -77.46 ;
      RECT 145.85 -74.35 146.2 -74.23 ;
      RECT 145.85 -71.12 146.2 -71 ;
      RECT 145.85 -67.89 146.2 -67.77 ;
      RECT 145.85 -64.66 146.2 -64.54 ;
      RECT 145.85 -61.43 146.2 -61.31 ;
      RECT 145.85 -58.2 146.2 -58.08 ;
      RECT 145.85 -54.97 146.2 -54.85 ;
      RECT 145.85 -51.74 146.2 -51.62 ;
      RECT 145.85 -48.51 146.2 -48.39 ;
      RECT 145.85 -45.28 146.2 -45.16 ;
      RECT 145.85 -42.05 146.2 -41.93 ;
      RECT 145.85 -38.82 146.2 -38.7 ;
      RECT 145.85 -35.59 146.2 -35.47 ;
      RECT 145.85 -32.36 146.2 -32.24 ;
      RECT 145.85 -29.13 146.2 -29.01 ;
      RECT 145.85 -25.9 146.2 -25.78 ;
      RECT 145.85 -22.67 146.2 -22.55 ;
      RECT 145.85 -19.44 146.2 -19.32 ;
      RECT 145.85 -16.21 146.2 -16.09 ;
      RECT 145.85 -12.98 146.2 -12.86 ;
      RECT 145.85 -9.75 146.2 -9.63 ;
      RECT 145.85 -6.52 146.2 -6.4 ;
      RECT 145.85 -3.29 146.2 -3.17 ;
      RECT 145.85 -0.06 146.2 0.06 ;
      RECT 146.055 -112.255 146.155 -111.775 ;
      RECT 146.055 -110.765 146.155 -110.295 ;
      RECT 145.965 -108.175 146.065 -107.215 ;
      RECT 145.965 2.175 146.065 3.135 ;
      RECT 145.365 -100.19 145.715 -100.07 ;
      RECT 145.365 -96.96 145.715 -96.84 ;
      RECT 145.365 -93.73 145.715 -93.61 ;
      RECT 145.365 -90.5 145.715 -90.38 ;
      RECT 145.365 -87.27 145.715 -87.15 ;
      RECT 145.365 -84.04 145.715 -83.92 ;
      RECT 145.365 -80.81 145.715 -80.69 ;
      RECT 145.365 -77.58 145.715 -77.46 ;
      RECT 145.365 -74.35 145.715 -74.23 ;
      RECT 145.365 -71.12 145.715 -71 ;
      RECT 145.365 -67.89 145.715 -67.77 ;
      RECT 145.365 -64.66 145.715 -64.54 ;
      RECT 145.365 -61.43 145.715 -61.31 ;
      RECT 145.365 -58.2 145.715 -58.08 ;
      RECT 145.365 -54.97 145.715 -54.85 ;
      RECT 145.365 -51.74 145.715 -51.62 ;
      RECT 145.365 -48.51 145.715 -48.39 ;
      RECT 145.365 -45.28 145.715 -45.16 ;
      RECT 145.365 -42.05 145.715 -41.93 ;
      RECT 145.365 -38.82 145.715 -38.7 ;
      RECT 145.365 -35.59 145.715 -35.47 ;
      RECT 145.365 -32.36 145.715 -32.24 ;
      RECT 145.365 -29.13 145.715 -29.01 ;
      RECT 145.365 -25.9 145.715 -25.78 ;
      RECT 145.365 -22.67 145.715 -22.55 ;
      RECT 145.365 -19.44 145.715 -19.32 ;
      RECT 145.365 -16.21 145.715 -16.09 ;
      RECT 145.365 -12.98 145.715 -12.86 ;
      RECT 145.365 -9.75 145.715 -9.63 ;
      RECT 145.365 -6.52 145.715 -6.4 ;
      RECT 145.365 -3.29 145.715 -3.17 ;
      RECT 145.365 -0.06 145.715 0.06 ;
      RECT 145.535 -108.175 145.635 -107.215 ;
      RECT 145.535 2.175 145.635 3.135 ;
      RECT 145.43 -110.765 145.6 -110.385 ;
      RECT 145.465 -112.245 145.565 -111.775 ;
      RECT 145.275 -108.175 145.375 -107.215 ;
      RECT 145.15 -101.06 145.25 -100.525 ;
      RECT 145.15 -99.735 145.25 -99.2 ;
      RECT 145.15 -97.83 145.25 -97.295 ;
      RECT 145.15 -96.505 145.25 -95.97 ;
      RECT 145.15 -94.6 145.25 -94.065 ;
      RECT 145.15 -93.275 145.25 -92.74 ;
      RECT 145.15 -91.37 145.25 -90.835 ;
      RECT 145.15 -90.045 145.25 -89.51 ;
      RECT 145.15 -88.14 145.25 -87.605 ;
      RECT 145.15 -86.815 145.25 -86.28 ;
      RECT 145.15 -84.91 145.25 -84.375 ;
      RECT 145.15 -83.585 145.25 -83.05 ;
      RECT 145.15 -81.68 145.25 -81.145 ;
      RECT 145.15 -80.355 145.25 -79.82 ;
      RECT 145.15 -78.45 145.25 -77.915 ;
      RECT 145.15 -77.125 145.25 -76.59 ;
      RECT 145.15 -75.22 145.25 -74.685 ;
      RECT 145.15 -73.895 145.25 -73.36 ;
      RECT 145.15 -71.99 145.25 -71.455 ;
      RECT 145.15 -70.665 145.25 -70.13 ;
      RECT 145.15 -68.76 145.25 -68.225 ;
      RECT 145.15 -67.435 145.25 -66.9 ;
      RECT 145.15 -65.53 145.25 -64.995 ;
      RECT 145.15 -64.205 145.25 -63.67 ;
      RECT 145.15 -62.3 145.25 -61.765 ;
      RECT 145.15 -60.975 145.25 -60.44 ;
      RECT 145.15 -59.07 145.25 -58.535 ;
      RECT 145.15 -57.745 145.25 -57.21 ;
      RECT 145.15 -55.84 145.25 -55.305 ;
      RECT 145.15 -54.515 145.25 -53.98 ;
      RECT 145.15 -52.61 145.25 -52.075 ;
      RECT 145.15 -51.285 145.25 -50.75 ;
      RECT 145.15 -49.38 145.25 -48.845 ;
      RECT 145.15 -48.055 145.25 -47.52 ;
      RECT 145.15 -46.15 145.25 -45.615 ;
      RECT 145.15 -44.825 145.25 -44.29 ;
      RECT 145.15 -42.92 145.25 -42.385 ;
      RECT 145.15 -41.595 145.25 -41.06 ;
      RECT 145.15 -39.69 145.25 -39.155 ;
      RECT 145.15 -38.365 145.25 -37.83 ;
      RECT 145.15 -36.46 145.25 -35.925 ;
      RECT 145.15 -35.135 145.25 -34.6 ;
      RECT 145.15 -33.23 145.25 -32.695 ;
      RECT 145.15 -31.905 145.25 -31.37 ;
      RECT 145.15 -30 145.25 -29.465 ;
      RECT 145.15 -28.675 145.25 -28.14 ;
      RECT 145.15 -26.77 145.25 -26.235 ;
      RECT 145.15 -25.445 145.25 -24.91 ;
      RECT 145.15 -23.54 145.25 -23.005 ;
      RECT 145.15 -22.215 145.25 -21.68 ;
      RECT 145.15 -20.31 145.25 -19.775 ;
      RECT 145.15 -18.985 145.25 -18.45 ;
      RECT 145.15 -17.08 145.25 -16.545 ;
      RECT 145.15 -15.755 145.25 -15.22 ;
      RECT 145.15 -13.85 145.25 -13.315 ;
      RECT 145.15 -12.525 145.25 -11.99 ;
      RECT 145.15 -10.62 145.25 -10.085 ;
      RECT 145.15 -9.295 145.25 -8.76 ;
      RECT 145.15 -7.39 145.25 -6.855 ;
      RECT 145.15 -6.065 145.25 -5.53 ;
      RECT 145.15 -4.16 145.25 -3.625 ;
      RECT 145.15 -2.835 145.25 -2.3 ;
      RECT 145.15 -0.93 145.25 -0.395 ;
      RECT 145.15 0.395 145.25 0.93 ;
      RECT 145.025 -108.175 145.125 -107.215 ;
      RECT 144.65 -100.19 145 -100.07 ;
      RECT 144.65 -96.96 145 -96.84 ;
      RECT 144.65 -93.73 145 -93.61 ;
      RECT 144.65 -90.5 145 -90.38 ;
      RECT 144.65 -87.27 145 -87.15 ;
      RECT 144.65 -84.04 145 -83.92 ;
      RECT 144.65 -80.81 145 -80.69 ;
      RECT 144.65 -77.58 145 -77.46 ;
      RECT 144.65 -74.35 145 -74.23 ;
      RECT 144.65 -71.12 145 -71 ;
      RECT 144.65 -67.89 145 -67.77 ;
      RECT 144.65 -64.66 145 -64.54 ;
      RECT 144.65 -61.43 145 -61.31 ;
      RECT 144.65 -58.2 145 -58.08 ;
      RECT 144.65 -54.97 145 -54.85 ;
      RECT 144.65 -51.74 145 -51.62 ;
      RECT 144.65 -48.51 145 -48.39 ;
      RECT 144.65 -45.28 145 -45.16 ;
      RECT 144.65 -42.05 145 -41.93 ;
      RECT 144.65 -38.82 145 -38.7 ;
      RECT 144.65 -35.59 145 -35.47 ;
      RECT 144.65 -32.36 145 -32.24 ;
      RECT 144.65 -29.13 145 -29.01 ;
      RECT 144.65 -25.9 145 -25.78 ;
      RECT 144.65 -22.67 145 -22.55 ;
      RECT 144.65 -19.44 145 -19.32 ;
      RECT 144.65 -16.21 145 -16.09 ;
      RECT 144.65 -12.98 145 -12.86 ;
      RECT 144.65 -9.75 145 -9.63 ;
      RECT 144.65 -6.52 145 -6.4 ;
      RECT 144.65 -3.29 145 -3.17 ;
      RECT 144.65 -0.06 145 0.06 ;
      RECT 144.765 -108.175 144.865 -107.215 ;
      RECT 144.765 2.175 144.865 3.135 ;
      RECT 144.665 -113.555 144.765 -113.085 ;
      RECT 144.165 -100.19 144.515 -100.07 ;
      RECT 144.165 -96.96 144.515 -96.84 ;
      RECT 144.165 -93.73 144.515 -93.61 ;
      RECT 144.165 -90.5 144.515 -90.38 ;
      RECT 144.165 -87.27 144.515 -87.15 ;
      RECT 144.165 -84.04 144.515 -83.92 ;
      RECT 144.165 -80.81 144.515 -80.69 ;
      RECT 144.165 -77.58 144.515 -77.46 ;
      RECT 144.165 -74.35 144.515 -74.23 ;
      RECT 144.165 -71.12 144.515 -71 ;
      RECT 144.165 -67.89 144.515 -67.77 ;
      RECT 144.165 -64.66 144.515 -64.54 ;
      RECT 144.165 -61.43 144.515 -61.31 ;
      RECT 144.165 -58.2 144.515 -58.08 ;
      RECT 144.165 -54.97 144.515 -54.85 ;
      RECT 144.165 -51.74 144.515 -51.62 ;
      RECT 144.165 -48.51 144.515 -48.39 ;
      RECT 144.165 -45.28 144.515 -45.16 ;
      RECT 144.165 -42.05 144.515 -41.93 ;
      RECT 144.165 -38.82 144.515 -38.7 ;
      RECT 144.165 -35.59 144.515 -35.47 ;
      RECT 144.165 -32.36 144.515 -32.24 ;
      RECT 144.165 -29.13 144.515 -29.01 ;
      RECT 144.165 -25.9 144.515 -25.78 ;
      RECT 144.165 -22.67 144.515 -22.55 ;
      RECT 144.165 -19.44 144.515 -19.32 ;
      RECT 144.165 -16.21 144.515 -16.09 ;
      RECT 144.165 -12.98 144.515 -12.86 ;
      RECT 144.165 -9.75 144.515 -9.63 ;
      RECT 144.165 -6.52 144.515 -6.4 ;
      RECT 144.165 -3.29 144.515 -3.17 ;
      RECT 144.165 -0.06 144.515 0.06 ;
      RECT 144.3 -110.735 144.45 -110.445 ;
      RECT 144.335 -108.175 144.435 -107.215 ;
      RECT 144.335 2.175 144.435 3.135 ;
      RECT 144.315 -112.19 144.415 -111.65 ;
      RECT 144.075 -113.555 144.175 -113.085 ;
      RECT 144.075 -108.175 144.175 -107.215 ;
      RECT 143.95 -101.06 144.05 -100.525 ;
      RECT 143.95 -99.735 144.05 -99.2 ;
      RECT 143.95 -97.83 144.05 -97.295 ;
      RECT 143.95 -96.505 144.05 -95.97 ;
      RECT 143.95 -94.6 144.05 -94.065 ;
      RECT 143.95 -93.275 144.05 -92.74 ;
      RECT 143.95 -91.37 144.05 -90.835 ;
      RECT 143.95 -90.045 144.05 -89.51 ;
      RECT 143.95 -88.14 144.05 -87.605 ;
      RECT 143.95 -86.815 144.05 -86.28 ;
      RECT 143.95 -84.91 144.05 -84.375 ;
      RECT 143.95 -83.585 144.05 -83.05 ;
      RECT 143.95 -81.68 144.05 -81.145 ;
      RECT 143.95 -80.355 144.05 -79.82 ;
      RECT 143.95 -78.45 144.05 -77.915 ;
      RECT 143.95 -77.125 144.05 -76.59 ;
      RECT 143.95 -75.22 144.05 -74.685 ;
      RECT 143.95 -73.895 144.05 -73.36 ;
      RECT 143.95 -71.99 144.05 -71.455 ;
      RECT 143.95 -70.665 144.05 -70.13 ;
      RECT 143.95 -68.76 144.05 -68.225 ;
      RECT 143.95 -67.435 144.05 -66.9 ;
      RECT 143.95 -65.53 144.05 -64.995 ;
      RECT 143.95 -64.205 144.05 -63.67 ;
      RECT 143.95 -62.3 144.05 -61.765 ;
      RECT 143.95 -60.975 144.05 -60.44 ;
      RECT 143.95 -59.07 144.05 -58.535 ;
      RECT 143.95 -57.745 144.05 -57.21 ;
      RECT 143.95 -55.84 144.05 -55.305 ;
      RECT 143.95 -54.515 144.05 -53.98 ;
      RECT 143.95 -52.61 144.05 -52.075 ;
      RECT 143.95 -51.285 144.05 -50.75 ;
      RECT 143.95 -49.38 144.05 -48.845 ;
      RECT 143.95 -48.055 144.05 -47.52 ;
      RECT 143.95 -46.15 144.05 -45.615 ;
      RECT 143.95 -44.825 144.05 -44.29 ;
      RECT 143.95 -42.92 144.05 -42.385 ;
      RECT 143.95 -41.595 144.05 -41.06 ;
      RECT 143.95 -39.69 144.05 -39.155 ;
      RECT 143.95 -38.365 144.05 -37.83 ;
      RECT 143.95 -36.46 144.05 -35.925 ;
      RECT 143.95 -35.135 144.05 -34.6 ;
      RECT 143.95 -33.23 144.05 -32.695 ;
      RECT 143.95 -31.905 144.05 -31.37 ;
      RECT 143.95 -30 144.05 -29.465 ;
      RECT 143.95 -28.675 144.05 -28.14 ;
      RECT 143.95 -26.77 144.05 -26.235 ;
      RECT 143.95 -25.445 144.05 -24.91 ;
      RECT 143.95 -23.54 144.05 -23.005 ;
      RECT 143.95 -22.215 144.05 -21.68 ;
      RECT 143.95 -20.31 144.05 -19.775 ;
      RECT 143.95 -18.985 144.05 -18.45 ;
      RECT 143.95 -17.08 144.05 -16.545 ;
      RECT 143.95 -15.755 144.05 -15.22 ;
      RECT 143.95 -13.85 144.05 -13.315 ;
      RECT 143.95 -12.525 144.05 -11.99 ;
      RECT 143.95 -10.62 144.05 -10.085 ;
      RECT 143.95 -9.295 144.05 -8.76 ;
      RECT 143.95 -7.39 144.05 -6.855 ;
      RECT 143.95 -6.065 144.05 -5.53 ;
      RECT 143.95 -4.16 144.05 -3.625 ;
      RECT 143.95 -2.835 144.05 -2.3 ;
      RECT 143.95 -0.93 144.05 -0.395 ;
      RECT 143.95 0.395 144.05 0.93 ;
      RECT 143.825 -104.945 143.925 -103.985 ;
      RECT 143.45 -100.19 143.8 -100.07 ;
      RECT 143.45 -96.96 143.8 -96.84 ;
      RECT 143.45 -93.73 143.8 -93.61 ;
      RECT 143.45 -90.5 143.8 -90.38 ;
      RECT 143.45 -87.27 143.8 -87.15 ;
      RECT 143.45 -84.04 143.8 -83.92 ;
      RECT 143.45 -80.81 143.8 -80.69 ;
      RECT 143.45 -77.58 143.8 -77.46 ;
      RECT 143.45 -74.35 143.8 -74.23 ;
      RECT 143.45 -71.12 143.8 -71 ;
      RECT 143.45 -67.89 143.8 -67.77 ;
      RECT 143.45 -64.66 143.8 -64.54 ;
      RECT 143.45 -61.43 143.8 -61.31 ;
      RECT 143.45 -58.2 143.8 -58.08 ;
      RECT 143.45 -54.97 143.8 -54.85 ;
      RECT 143.45 -51.74 143.8 -51.62 ;
      RECT 143.45 -48.51 143.8 -48.39 ;
      RECT 143.45 -45.28 143.8 -45.16 ;
      RECT 143.45 -42.05 143.8 -41.93 ;
      RECT 143.45 -38.82 143.8 -38.7 ;
      RECT 143.45 -35.59 143.8 -35.47 ;
      RECT 143.45 -32.36 143.8 -32.24 ;
      RECT 143.45 -29.13 143.8 -29.01 ;
      RECT 143.45 -25.9 143.8 -25.78 ;
      RECT 143.45 -22.67 143.8 -22.55 ;
      RECT 143.45 -19.44 143.8 -19.32 ;
      RECT 143.45 -16.21 143.8 -16.09 ;
      RECT 143.45 -12.98 143.8 -12.86 ;
      RECT 143.45 -9.75 143.8 -9.63 ;
      RECT 143.45 -6.52 143.8 -6.4 ;
      RECT 143.45 -3.29 143.8 -3.17 ;
      RECT 143.45 -0.06 143.8 0.06 ;
      RECT 143.565 -104.945 143.665 -103.985 ;
      RECT 143.565 2.175 143.665 3.135 ;
      RECT 143.275 -112.255 143.375 -111.775 ;
      RECT 143.275 -110.765 143.375 -110.295 ;
      RECT 142.965 -100.19 143.315 -100.07 ;
      RECT 142.965 -96.96 143.315 -96.84 ;
      RECT 142.965 -93.73 143.315 -93.61 ;
      RECT 142.965 -90.5 143.315 -90.38 ;
      RECT 142.965 -87.27 143.315 -87.15 ;
      RECT 142.965 -84.04 143.315 -83.92 ;
      RECT 142.965 -80.81 143.315 -80.69 ;
      RECT 142.965 -77.58 143.315 -77.46 ;
      RECT 142.965 -74.35 143.315 -74.23 ;
      RECT 142.965 -71.12 143.315 -71 ;
      RECT 142.965 -67.89 143.315 -67.77 ;
      RECT 142.965 -64.66 143.315 -64.54 ;
      RECT 142.965 -61.43 143.315 -61.31 ;
      RECT 142.965 -58.2 143.315 -58.08 ;
      RECT 142.965 -54.97 143.315 -54.85 ;
      RECT 142.965 -51.74 143.315 -51.62 ;
      RECT 142.965 -48.51 143.315 -48.39 ;
      RECT 142.965 -45.28 143.315 -45.16 ;
      RECT 142.965 -42.05 143.315 -41.93 ;
      RECT 142.965 -38.82 143.315 -38.7 ;
      RECT 142.965 -35.59 143.315 -35.47 ;
      RECT 142.965 -32.36 143.315 -32.24 ;
      RECT 142.965 -29.13 143.315 -29.01 ;
      RECT 142.965 -25.9 143.315 -25.78 ;
      RECT 142.965 -22.67 143.315 -22.55 ;
      RECT 142.965 -19.44 143.315 -19.32 ;
      RECT 142.965 -16.21 143.315 -16.09 ;
      RECT 142.965 -12.98 143.315 -12.86 ;
      RECT 142.965 -9.75 143.315 -9.63 ;
      RECT 142.965 -6.52 143.315 -6.4 ;
      RECT 142.965 -3.29 143.315 -3.17 ;
      RECT 142.965 -0.06 143.315 0.06 ;
      RECT 143.135 -104.945 143.235 -103.985 ;
      RECT 143.135 2.175 143.235 3.135 ;
      RECT 139.235 -108.655 143.015 -108.535 ;
      RECT 142.875 -104.945 142.975 -103.985 ;
      RECT 142.75 -101.06 142.85 -100.525 ;
      RECT 142.75 -99.735 142.85 -99.2 ;
      RECT 142.75 -97.83 142.85 -97.295 ;
      RECT 142.75 -96.505 142.85 -95.97 ;
      RECT 142.75 -94.6 142.85 -94.065 ;
      RECT 142.75 -93.275 142.85 -92.74 ;
      RECT 142.75 -91.37 142.85 -90.835 ;
      RECT 142.75 -90.045 142.85 -89.51 ;
      RECT 142.75 -88.14 142.85 -87.605 ;
      RECT 142.75 -86.815 142.85 -86.28 ;
      RECT 142.75 -84.91 142.85 -84.375 ;
      RECT 142.75 -83.585 142.85 -83.05 ;
      RECT 142.75 -81.68 142.85 -81.145 ;
      RECT 142.75 -80.355 142.85 -79.82 ;
      RECT 142.75 -78.45 142.85 -77.915 ;
      RECT 142.75 -77.125 142.85 -76.59 ;
      RECT 142.75 -75.22 142.85 -74.685 ;
      RECT 142.75 -73.895 142.85 -73.36 ;
      RECT 142.75 -71.99 142.85 -71.455 ;
      RECT 142.75 -70.665 142.85 -70.13 ;
      RECT 142.75 -68.76 142.85 -68.225 ;
      RECT 142.75 -67.435 142.85 -66.9 ;
      RECT 142.75 -65.53 142.85 -64.995 ;
      RECT 142.75 -64.205 142.85 -63.67 ;
      RECT 142.75 -62.3 142.85 -61.765 ;
      RECT 142.75 -60.975 142.85 -60.44 ;
      RECT 142.75 -59.07 142.85 -58.535 ;
      RECT 142.75 -57.745 142.85 -57.21 ;
      RECT 142.75 -55.84 142.85 -55.305 ;
      RECT 142.75 -54.515 142.85 -53.98 ;
      RECT 142.75 -52.61 142.85 -52.075 ;
      RECT 142.75 -51.285 142.85 -50.75 ;
      RECT 142.75 -49.38 142.85 -48.845 ;
      RECT 142.75 -48.055 142.85 -47.52 ;
      RECT 142.75 -46.15 142.85 -45.615 ;
      RECT 142.75 -44.825 142.85 -44.29 ;
      RECT 142.75 -42.92 142.85 -42.385 ;
      RECT 142.75 -41.595 142.85 -41.06 ;
      RECT 142.75 -39.69 142.85 -39.155 ;
      RECT 142.75 -38.365 142.85 -37.83 ;
      RECT 142.75 -36.46 142.85 -35.925 ;
      RECT 142.75 -35.135 142.85 -34.6 ;
      RECT 142.75 -33.23 142.85 -32.695 ;
      RECT 142.75 -31.905 142.85 -31.37 ;
      RECT 142.75 -30 142.85 -29.465 ;
      RECT 142.75 -28.675 142.85 -28.14 ;
      RECT 142.75 -26.77 142.85 -26.235 ;
      RECT 142.75 -25.445 142.85 -24.91 ;
      RECT 142.75 -23.54 142.85 -23.005 ;
      RECT 142.75 -22.215 142.85 -21.68 ;
      RECT 142.75 -20.31 142.85 -19.775 ;
      RECT 142.75 -18.985 142.85 -18.45 ;
      RECT 142.75 -17.08 142.85 -16.545 ;
      RECT 142.75 -15.755 142.85 -15.22 ;
      RECT 142.75 -13.85 142.85 -13.315 ;
      RECT 142.75 -12.525 142.85 -11.99 ;
      RECT 142.75 -10.62 142.85 -10.085 ;
      RECT 142.75 -9.295 142.85 -8.76 ;
      RECT 142.75 -7.39 142.85 -6.855 ;
      RECT 142.75 -6.065 142.85 -5.53 ;
      RECT 142.75 -4.16 142.85 -3.625 ;
      RECT 142.75 -2.835 142.85 -2.3 ;
      RECT 142.75 -0.93 142.85 -0.395 ;
      RECT 142.75 0.395 142.85 0.93 ;
      RECT 142.685 -110.75 142.805 -110.37 ;
      RECT 142.685 -112.245 142.785 -111.775 ;
      RECT 142.625 -104.945 142.725 -103.985 ;
      RECT 142.25 -100.19 142.6 -100.07 ;
      RECT 142.25 -96.96 142.6 -96.84 ;
      RECT 142.25 -93.73 142.6 -93.61 ;
      RECT 142.25 -90.5 142.6 -90.38 ;
      RECT 142.25 -87.27 142.6 -87.15 ;
      RECT 142.25 -84.04 142.6 -83.92 ;
      RECT 142.25 -80.81 142.6 -80.69 ;
      RECT 142.25 -77.58 142.6 -77.46 ;
      RECT 142.25 -74.35 142.6 -74.23 ;
      RECT 142.25 -71.12 142.6 -71 ;
      RECT 142.25 -67.89 142.6 -67.77 ;
      RECT 142.25 -64.66 142.6 -64.54 ;
      RECT 142.25 -61.43 142.6 -61.31 ;
      RECT 142.25 -58.2 142.6 -58.08 ;
      RECT 142.25 -54.97 142.6 -54.85 ;
      RECT 142.25 -51.74 142.6 -51.62 ;
      RECT 142.25 -48.51 142.6 -48.39 ;
      RECT 142.25 -45.28 142.6 -45.16 ;
      RECT 142.25 -42.05 142.6 -41.93 ;
      RECT 142.25 -38.82 142.6 -38.7 ;
      RECT 142.25 -35.59 142.6 -35.47 ;
      RECT 142.25 -32.36 142.6 -32.24 ;
      RECT 142.25 -29.13 142.6 -29.01 ;
      RECT 142.25 -25.9 142.6 -25.78 ;
      RECT 142.25 -22.67 142.6 -22.55 ;
      RECT 142.25 -19.44 142.6 -19.32 ;
      RECT 142.25 -16.21 142.6 -16.09 ;
      RECT 142.25 -12.98 142.6 -12.86 ;
      RECT 142.25 -9.75 142.6 -9.63 ;
      RECT 142.25 -6.52 142.6 -6.4 ;
      RECT 142.25 -3.29 142.6 -3.17 ;
      RECT 142.25 -0.06 142.6 0.06 ;
      RECT 142.365 -104.945 142.465 -103.985 ;
      RECT 142.365 2.175 142.465 3.135 ;
      RECT 142.095 -109.595 142.23 -109.275 ;
      RECT 141.765 -100.19 142.115 -100.07 ;
      RECT 141.765 -96.96 142.115 -96.84 ;
      RECT 141.765 -93.73 142.115 -93.61 ;
      RECT 141.765 -90.5 142.115 -90.38 ;
      RECT 141.765 -87.27 142.115 -87.15 ;
      RECT 141.765 -84.04 142.115 -83.92 ;
      RECT 141.765 -80.81 142.115 -80.69 ;
      RECT 141.765 -77.58 142.115 -77.46 ;
      RECT 141.765 -74.35 142.115 -74.23 ;
      RECT 141.765 -71.12 142.115 -71 ;
      RECT 141.765 -67.89 142.115 -67.77 ;
      RECT 141.765 -64.66 142.115 -64.54 ;
      RECT 141.765 -61.43 142.115 -61.31 ;
      RECT 141.765 -58.2 142.115 -58.08 ;
      RECT 141.765 -54.97 142.115 -54.85 ;
      RECT 141.765 -51.74 142.115 -51.62 ;
      RECT 141.765 -48.51 142.115 -48.39 ;
      RECT 141.765 -45.28 142.115 -45.16 ;
      RECT 141.765 -42.05 142.115 -41.93 ;
      RECT 141.765 -38.82 142.115 -38.7 ;
      RECT 141.765 -35.59 142.115 -35.47 ;
      RECT 141.765 -32.36 142.115 -32.24 ;
      RECT 141.765 -29.13 142.115 -29.01 ;
      RECT 141.765 -25.9 142.115 -25.78 ;
      RECT 141.765 -22.67 142.115 -22.55 ;
      RECT 141.765 -19.44 142.115 -19.32 ;
      RECT 141.765 -16.21 142.115 -16.09 ;
      RECT 141.765 -12.98 142.115 -12.86 ;
      RECT 141.765 -9.75 142.115 -9.63 ;
      RECT 141.765 -6.52 142.115 -6.4 ;
      RECT 141.765 -3.29 142.115 -3.17 ;
      RECT 141.765 -0.06 142.115 0.06 ;
      RECT 141.935 -104.945 142.035 -103.985 ;
      RECT 141.935 2.175 142.035 3.135 ;
      RECT 141.76 -109.595 141.905 -109.275 ;
      RECT 141.675 -104.945 141.775 -103.985 ;
      RECT 141.55 -101.06 141.65 -100.525 ;
      RECT 141.55 -99.735 141.65 -99.2 ;
      RECT 141.55 -97.83 141.65 -97.295 ;
      RECT 141.55 -96.505 141.65 -95.97 ;
      RECT 141.55 -94.6 141.65 -94.065 ;
      RECT 141.55 -93.275 141.65 -92.74 ;
      RECT 141.55 -91.37 141.65 -90.835 ;
      RECT 141.55 -90.045 141.65 -89.51 ;
      RECT 141.55 -88.14 141.65 -87.605 ;
      RECT 141.55 -86.815 141.65 -86.28 ;
      RECT 141.55 -84.91 141.65 -84.375 ;
      RECT 141.55 -83.585 141.65 -83.05 ;
      RECT 141.55 -81.68 141.65 -81.145 ;
      RECT 141.55 -80.355 141.65 -79.82 ;
      RECT 141.55 -78.45 141.65 -77.915 ;
      RECT 141.55 -77.125 141.65 -76.59 ;
      RECT 141.55 -75.22 141.65 -74.685 ;
      RECT 141.55 -73.895 141.65 -73.36 ;
      RECT 141.55 -71.99 141.65 -71.455 ;
      RECT 141.55 -70.665 141.65 -70.13 ;
      RECT 141.55 -68.76 141.65 -68.225 ;
      RECT 141.55 -67.435 141.65 -66.9 ;
      RECT 141.55 -65.53 141.65 -64.995 ;
      RECT 141.55 -64.205 141.65 -63.67 ;
      RECT 141.55 -62.3 141.65 -61.765 ;
      RECT 141.55 -60.975 141.65 -60.44 ;
      RECT 141.55 -59.07 141.65 -58.535 ;
      RECT 141.55 -57.745 141.65 -57.21 ;
      RECT 141.55 -55.84 141.65 -55.305 ;
      RECT 141.55 -54.515 141.65 -53.98 ;
      RECT 141.55 -52.61 141.65 -52.075 ;
      RECT 141.55 -51.285 141.65 -50.75 ;
      RECT 141.55 -49.38 141.65 -48.845 ;
      RECT 141.55 -48.055 141.65 -47.52 ;
      RECT 141.55 -46.15 141.65 -45.615 ;
      RECT 141.55 -44.825 141.65 -44.29 ;
      RECT 141.55 -42.92 141.65 -42.385 ;
      RECT 141.55 -41.595 141.65 -41.06 ;
      RECT 141.55 -39.69 141.65 -39.155 ;
      RECT 141.55 -38.365 141.65 -37.83 ;
      RECT 141.55 -36.46 141.65 -35.925 ;
      RECT 141.55 -35.135 141.65 -34.6 ;
      RECT 141.55 -33.23 141.65 -32.695 ;
      RECT 141.55 -31.905 141.65 -31.37 ;
      RECT 141.55 -30 141.65 -29.465 ;
      RECT 141.55 -28.675 141.65 -28.14 ;
      RECT 141.55 -26.77 141.65 -26.235 ;
      RECT 141.55 -25.445 141.65 -24.91 ;
      RECT 141.55 -23.54 141.65 -23.005 ;
      RECT 141.55 -22.215 141.65 -21.68 ;
      RECT 141.55 -20.31 141.65 -19.775 ;
      RECT 141.55 -18.985 141.65 -18.45 ;
      RECT 141.55 -17.08 141.65 -16.545 ;
      RECT 141.55 -15.755 141.65 -15.22 ;
      RECT 141.55 -13.85 141.65 -13.315 ;
      RECT 141.55 -12.525 141.65 -11.99 ;
      RECT 141.55 -10.62 141.65 -10.085 ;
      RECT 141.55 -9.295 141.65 -8.76 ;
      RECT 141.55 -7.39 141.65 -6.855 ;
      RECT 141.55 -6.065 141.65 -5.53 ;
      RECT 141.55 -4.16 141.65 -3.625 ;
      RECT 141.55 -2.835 141.65 -2.3 ;
      RECT 141.55 -0.93 141.65 -0.395 ;
      RECT 141.55 0.395 141.65 0.93 ;
      RECT 141.425 -108.175 141.525 -107.215 ;
      RECT 141.05 -100.19 141.4 -100.07 ;
      RECT 141.05 -96.96 141.4 -96.84 ;
      RECT 141.05 -93.73 141.4 -93.61 ;
      RECT 141.05 -90.5 141.4 -90.38 ;
      RECT 141.05 -87.27 141.4 -87.15 ;
      RECT 141.05 -84.04 141.4 -83.92 ;
      RECT 141.05 -80.81 141.4 -80.69 ;
      RECT 141.05 -77.58 141.4 -77.46 ;
      RECT 141.05 -74.35 141.4 -74.23 ;
      RECT 141.05 -71.12 141.4 -71 ;
      RECT 141.05 -67.89 141.4 -67.77 ;
      RECT 141.05 -64.66 141.4 -64.54 ;
      RECT 141.05 -61.43 141.4 -61.31 ;
      RECT 141.05 -58.2 141.4 -58.08 ;
      RECT 141.05 -54.97 141.4 -54.85 ;
      RECT 141.05 -51.74 141.4 -51.62 ;
      RECT 141.05 -48.51 141.4 -48.39 ;
      RECT 141.05 -45.28 141.4 -45.16 ;
      RECT 141.05 -42.05 141.4 -41.93 ;
      RECT 141.05 -38.82 141.4 -38.7 ;
      RECT 141.05 -35.59 141.4 -35.47 ;
      RECT 141.05 -32.36 141.4 -32.24 ;
      RECT 141.05 -29.13 141.4 -29.01 ;
      RECT 141.05 -25.9 141.4 -25.78 ;
      RECT 141.05 -22.67 141.4 -22.55 ;
      RECT 141.05 -19.44 141.4 -19.32 ;
      RECT 141.05 -16.21 141.4 -16.09 ;
      RECT 141.05 -12.98 141.4 -12.86 ;
      RECT 141.05 -9.75 141.4 -9.63 ;
      RECT 141.05 -6.52 141.4 -6.4 ;
      RECT 141.05 -3.29 141.4 -3.17 ;
      RECT 141.05 -0.06 141.4 0.06 ;
      RECT 141.255 -112.255 141.355 -111.775 ;
      RECT 141.255 -110.765 141.355 -110.295 ;
      RECT 141.165 -108.175 141.265 -107.215 ;
      RECT 141.165 2.175 141.265 3.135 ;
      RECT 140.565 -100.19 140.915 -100.07 ;
      RECT 140.565 -96.96 140.915 -96.84 ;
      RECT 140.565 -93.73 140.915 -93.61 ;
      RECT 140.565 -90.5 140.915 -90.38 ;
      RECT 140.565 -87.27 140.915 -87.15 ;
      RECT 140.565 -84.04 140.915 -83.92 ;
      RECT 140.565 -80.81 140.915 -80.69 ;
      RECT 140.565 -77.58 140.915 -77.46 ;
      RECT 140.565 -74.35 140.915 -74.23 ;
      RECT 140.565 -71.12 140.915 -71 ;
      RECT 140.565 -67.89 140.915 -67.77 ;
      RECT 140.565 -64.66 140.915 -64.54 ;
      RECT 140.565 -61.43 140.915 -61.31 ;
      RECT 140.565 -58.2 140.915 -58.08 ;
      RECT 140.565 -54.97 140.915 -54.85 ;
      RECT 140.565 -51.74 140.915 -51.62 ;
      RECT 140.565 -48.51 140.915 -48.39 ;
      RECT 140.565 -45.28 140.915 -45.16 ;
      RECT 140.565 -42.05 140.915 -41.93 ;
      RECT 140.565 -38.82 140.915 -38.7 ;
      RECT 140.565 -35.59 140.915 -35.47 ;
      RECT 140.565 -32.36 140.915 -32.24 ;
      RECT 140.565 -29.13 140.915 -29.01 ;
      RECT 140.565 -25.9 140.915 -25.78 ;
      RECT 140.565 -22.67 140.915 -22.55 ;
      RECT 140.565 -19.44 140.915 -19.32 ;
      RECT 140.565 -16.21 140.915 -16.09 ;
      RECT 140.565 -12.98 140.915 -12.86 ;
      RECT 140.565 -9.75 140.915 -9.63 ;
      RECT 140.565 -6.52 140.915 -6.4 ;
      RECT 140.565 -3.29 140.915 -3.17 ;
      RECT 140.565 -0.06 140.915 0.06 ;
      RECT 140.735 -108.175 140.835 -107.215 ;
      RECT 140.735 2.175 140.835 3.135 ;
      RECT 140.63 -110.765 140.8 -110.385 ;
      RECT 140.665 -112.245 140.765 -111.775 ;
      RECT 140.475 -108.175 140.575 -107.215 ;
      RECT 140.35 -101.06 140.45 -100.525 ;
      RECT 140.35 -99.735 140.45 -99.2 ;
      RECT 140.35 -97.83 140.45 -97.295 ;
      RECT 140.35 -96.505 140.45 -95.97 ;
      RECT 140.35 -94.6 140.45 -94.065 ;
      RECT 140.35 -93.275 140.45 -92.74 ;
      RECT 140.35 -91.37 140.45 -90.835 ;
      RECT 140.35 -90.045 140.45 -89.51 ;
      RECT 140.35 -88.14 140.45 -87.605 ;
      RECT 140.35 -86.815 140.45 -86.28 ;
      RECT 140.35 -84.91 140.45 -84.375 ;
      RECT 140.35 -83.585 140.45 -83.05 ;
      RECT 140.35 -81.68 140.45 -81.145 ;
      RECT 140.35 -80.355 140.45 -79.82 ;
      RECT 140.35 -78.45 140.45 -77.915 ;
      RECT 140.35 -77.125 140.45 -76.59 ;
      RECT 140.35 -75.22 140.45 -74.685 ;
      RECT 140.35 -73.895 140.45 -73.36 ;
      RECT 140.35 -71.99 140.45 -71.455 ;
      RECT 140.35 -70.665 140.45 -70.13 ;
      RECT 140.35 -68.76 140.45 -68.225 ;
      RECT 140.35 -67.435 140.45 -66.9 ;
      RECT 140.35 -65.53 140.45 -64.995 ;
      RECT 140.35 -64.205 140.45 -63.67 ;
      RECT 140.35 -62.3 140.45 -61.765 ;
      RECT 140.35 -60.975 140.45 -60.44 ;
      RECT 140.35 -59.07 140.45 -58.535 ;
      RECT 140.35 -57.745 140.45 -57.21 ;
      RECT 140.35 -55.84 140.45 -55.305 ;
      RECT 140.35 -54.515 140.45 -53.98 ;
      RECT 140.35 -52.61 140.45 -52.075 ;
      RECT 140.35 -51.285 140.45 -50.75 ;
      RECT 140.35 -49.38 140.45 -48.845 ;
      RECT 140.35 -48.055 140.45 -47.52 ;
      RECT 140.35 -46.15 140.45 -45.615 ;
      RECT 140.35 -44.825 140.45 -44.29 ;
      RECT 140.35 -42.92 140.45 -42.385 ;
      RECT 140.35 -41.595 140.45 -41.06 ;
      RECT 140.35 -39.69 140.45 -39.155 ;
      RECT 140.35 -38.365 140.45 -37.83 ;
      RECT 140.35 -36.46 140.45 -35.925 ;
      RECT 140.35 -35.135 140.45 -34.6 ;
      RECT 140.35 -33.23 140.45 -32.695 ;
      RECT 140.35 -31.905 140.45 -31.37 ;
      RECT 140.35 -30 140.45 -29.465 ;
      RECT 140.35 -28.675 140.45 -28.14 ;
      RECT 140.35 -26.77 140.45 -26.235 ;
      RECT 140.35 -25.445 140.45 -24.91 ;
      RECT 140.35 -23.54 140.45 -23.005 ;
      RECT 140.35 -22.215 140.45 -21.68 ;
      RECT 140.35 -20.31 140.45 -19.775 ;
      RECT 140.35 -18.985 140.45 -18.45 ;
      RECT 140.35 -17.08 140.45 -16.545 ;
      RECT 140.35 -15.755 140.45 -15.22 ;
      RECT 140.35 -13.85 140.45 -13.315 ;
      RECT 140.35 -12.525 140.45 -11.99 ;
      RECT 140.35 -10.62 140.45 -10.085 ;
      RECT 140.35 -9.295 140.45 -8.76 ;
      RECT 140.35 -7.39 140.45 -6.855 ;
      RECT 140.35 -6.065 140.45 -5.53 ;
      RECT 140.35 -4.16 140.45 -3.625 ;
      RECT 140.35 -2.835 140.45 -2.3 ;
      RECT 140.35 -0.93 140.45 -0.395 ;
      RECT 140.35 0.395 140.45 0.93 ;
      RECT 140.225 -108.175 140.325 -107.215 ;
      RECT 139.85 -100.19 140.2 -100.07 ;
      RECT 139.85 -96.96 140.2 -96.84 ;
      RECT 139.85 -93.73 140.2 -93.61 ;
      RECT 139.85 -90.5 140.2 -90.38 ;
      RECT 139.85 -87.27 140.2 -87.15 ;
      RECT 139.85 -84.04 140.2 -83.92 ;
      RECT 139.85 -80.81 140.2 -80.69 ;
      RECT 139.85 -77.58 140.2 -77.46 ;
      RECT 139.85 -74.35 140.2 -74.23 ;
      RECT 139.85 -71.12 140.2 -71 ;
      RECT 139.85 -67.89 140.2 -67.77 ;
      RECT 139.85 -64.66 140.2 -64.54 ;
      RECT 139.85 -61.43 140.2 -61.31 ;
      RECT 139.85 -58.2 140.2 -58.08 ;
      RECT 139.85 -54.97 140.2 -54.85 ;
      RECT 139.85 -51.74 140.2 -51.62 ;
      RECT 139.85 -48.51 140.2 -48.39 ;
      RECT 139.85 -45.28 140.2 -45.16 ;
      RECT 139.85 -42.05 140.2 -41.93 ;
      RECT 139.85 -38.82 140.2 -38.7 ;
      RECT 139.85 -35.59 140.2 -35.47 ;
      RECT 139.85 -32.36 140.2 -32.24 ;
      RECT 139.85 -29.13 140.2 -29.01 ;
      RECT 139.85 -25.9 140.2 -25.78 ;
      RECT 139.85 -22.67 140.2 -22.55 ;
      RECT 139.85 -19.44 140.2 -19.32 ;
      RECT 139.85 -16.21 140.2 -16.09 ;
      RECT 139.85 -12.98 140.2 -12.86 ;
      RECT 139.85 -9.75 140.2 -9.63 ;
      RECT 139.85 -6.52 140.2 -6.4 ;
      RECT 139.85 -3.29 140.2 -3.17 ;
      RECT 139.85 -0.06 140.2 0.06 ;
      RECT 139.965 -108.175 140.065 -107.215 ;
      RECT 139.965 2.175 140.065 3.135 ;
      RECT 139.865 -113.555 139.965 -113.085 ;
      RECT 139.365 -100.19 139.715 -100.07 ;
      RECT 139.365 -96.96 139.715 -96.84 ;
      RECT 139.365 -93.73 139.715 -93.61 ;
      RECT 139.365 -90.5 139.715 -90.38 ;
      RECT 139.365 -87.27 139.715 -87.15 ;
      RECT 139.365 -84.04 139.715 -83.92 ;
      RECT 139.365 -80.81 139.715 -80.69 ;
      RECT 139.365 -77.58 139.715 -77.46 ;
      RECT 139.365 -74.35 139.715 -74.23 ;
      RECT 139.365 -71.12 139.715 -71 ;
      RECT 139.365 -67.89 139.715 -67.77 ;
      RECT 139.365 -64.66 139.715 -64.54 ;
      RECT 139.365 -61.43 139.715 -61.31 ;
      RECT 139.365 -58.2 139.715 -58.08 ;
      RECT 139.365 -54.97 139.715 -54.85 ;
      RECT 139.365 -51.74 139.715 -51.62 ;
      RECT 139.365 -48.51 139.715 -48.39 ;
      RECT 139.365 -45.28 139.715 -45.16 ;
      RECT 139.365 -42.05 139.715 -41.93 ;
      RECT 139.365 -38.82 139.715 -38.7 ;
      RECT 139.365 -35.59 139.715 -35.47 ;
      RECT 139.365 -32.36 139.715 -32.24 ;
      RECT 139.365 -29.13 139.715 -29.01 ;
      RECT 139.365 -25.9 139.715 -25.78 ;
      RECT 139.365 -22.67 139.715 -22.55 ;
      RECT 139.365 -19.44 139.715 -19.32 ;
      RECT 139.365 -16.21 139.715 -16.09 ;
      RECT 139.365 -12.98 139.715 -12.86 ;
      RECT 139.365 -9.75 139.715 -9.63 ;
      RECT 139.365 -6.52 139.715 -6.4 ;
      RECT 139.365 -3.29 139.715 -3.17 ;
      RECT 139.365 -0.06 139.715 0.06 ;
      RECT 139.5 -110.735 139.65 -110.445 ;
      RECT 139.535 -108.175 139.635 -107.215 ;
      RECT 139.535 2.175 139.635 3.135 ;
      RECT 139.515 -112.19 139.615 -111.65 ;
      RECT 139.275 -113.555 139.375 -113.085 ;
      RECT 139.275 -108.175 139.375 -107.215 ;
      RECT 139.15 -101.06 139.25 -100.525 ;
      RECT 139.15 -99.735 139.25 -99.2 ;
      RECT 139.15 -97.83 139.25 -97.295 ;
      RECT 139.15 -96.505 139.25 -95.97 ;
      RECT 139.15 -94.6 139.25 -94.065 ;
      RECT 139.15 -93.275 139.25 -92.74 ;
      RECT 139.15 -91.37 139.25 -90.835 ;
      RECT 139.15 -90.045 139.25 -89.51 ;
      RECT 139.15 -88.14 139.25 -87.605 ;
      RECT 139.15 -86.815 139.25 -86.28 ;
      RECT 139.15 -84.91 139.25 -84.375 ;
      RECT 139.15 -83.585 139.25 -83.05 ;
      RECT 139.15 -81.68 139.25 -81.145 ;
      RECT 139.15 -80.355 139.25 -79.82 ;
      RECT 139.15 -78.45 139.25 -77.915 ;
      RECT 139.15 -77.125 139.25 -76.59 ;
      RECT 139.15 -75.22 139.25 -74.685 ;
      RECT 139.15 -73.895 139.25 -73.36 ;
      RECT 139.15 -71.99 139.25 -71.455 ;
      RECT 139.15 -70.665 139.25 -70.13 ;
      RECT 139.15 -68.76 139.25 -68.225 ;
      RECT 139.15 -67.435 139.25 -66.9 ;
      RECT 139.15 -65.53 139.25 -64.995 ;
      RECT 139.15 -64.205 139.25 -63.67 ;
      RECT 139.15 -62.3 139.25 -61.765 ;
      RECT 139.15 -60.975 139.25 -60.44 ;
      RECT 139.15 -59.07 139.25 -58.535 ;
      RECT 139.15 -57.745 139.25 -57.21 ;
      RECT 139.15 -55.84 139.25 -55.305 ;
      RECT 139.15 -54.515 139.25 -53.98 ;
      RECT 139.15 -52.61 139.25 -52.075 ;
      RECT 139.15 -51.285 139.25 -50.75 ;
      RECT 139.15 -49.38 139.25 -48.845 ;
      RECT 139.15 -48.055 139.25 -47.52 ;
      RECT 139.15 -46.15 139.25 -45.615 ;
      RECT 139.15 -44.825 139.25 -44.29 ;
      RECT 139.15 -42.92 139.25 -42.385 ;
      RECT 139.15 -41.595 139.25 -41.06 ;
      RECT 139.15 -39.69 139.25 -39.155 ;
      RECT 139.15 -38.365 139.25 -37.83 ;
      RECT 139.15 -36.46 139.25 -35.925 ;
      RECT 139.15 -35.135 139.25 -34.6 ;
      RECT 139.15 -33.23 139.25 -32.695 ;
      RECT 139.15 -31.905 139.25 -31.37 ;
      RECT 139.15 -30 139.25 -29.465 ;
      RECT 139.15 -28.675 139.25 -28.14 ;
      RECT 139.15 -26.77 139.25 -26.235 ;
      RECT 139.15 -25.445 139.25 -24.91 ;
      RECT 139.15 -23.54 139.25 -23.005 ;
      RECT 139.15 -22.215 139.25 -21.68 ;
      RECT 139.15 -20.31 139.25 -19.775 ;
      RECT 139.15 -18.985 139.25 -18.45 ;
      RECT 139.15 -17.08 139.25 -16.545 ;
      RECT 139.15 -15.755 139.25 -15.22 ;
      RECT 139.15 -13.85 139.25 -13.315 ;
      RECT 139.15 -12.525 139.25 -11.99 ;
      RECT 139.15 -10.62 139.25 -10.085 ;
      RECT 139.15 -9.295 139.25 -8.76 ;
      RECT 139.15 -7.39 139.25 -6.855 ;
      RECT 139.15 -6.065 139.25 -5.53 ;
      RECT 139.15 -4.16 139.25 -3.625 ;
      RECT 139.15 -2.835 139.25 -2.3 ;
      RECT 139.15 -0.93 139.25 -0.395 ;
      RECT 139.15 0.395 139.25 0.93 ;
      RECT 139.025 -104.945 139.125 -103.985 ;
      RECT 138.65 -100.19 139 -100.07 ;
      RECT 138.65 -96.96 139 -96.84 ;
      RECT 138.65 -93.73 139 -93.61 ;
      RECT 138.65 -90.5 139 -90.38 ;
      RECT 138.65 -87.27 139 -87.15 ;
      RECT 138.65 -84.04 139 -83.92 ;
      RECT 138.65 -80.81 139 -80.69 ;
      RECT 138.65 -77.58 139 -77.46 ;
      RECT 138.65 -74.35 139 -74.23 ;
      RECT 138.65 -71.12 139 -71 ;
      RECT 138.65 -67.89 139 -67.77 ;
      RECT 138.65 -64.66 139 -64.54 ;
      RECT 138.65 -61.43 139 -61.31 ;
      RECT 138.65 -58.2 139 -58.08 ;
      RECT 138.65 -54.97 139 -54.85 ;
      RECT 138.65 -51.74 139 -51.62 ;
      RECT 138.65 -48.51 139 -48.39 ;
      RECT 138.65 -45.28 139 -45.16 ;
      RECT 138.65 -42.05 139 -41.93 ;
      RECT 138.65 -38.82 139 -38.7 ;
      RECT 138.65 -35.59 139 -35.47 ;
      RECT 138.65 -32.36 139 -32.24 ;
      RECT 138.65 -29.13 139 -29.01 ;
      RECT 138.65 -25.9 139 -25.78 ;
      RECT 138.65 -22.67 139 -22.55 ;
      RECT 138.65 -19.44 139 -19.32 ;
      RECT 138.65 -16.21 139 -16.09 ;
      RECT 138.65 -12.98 139 -12.86 ;
      RECT 138.65 -9.75 139 -9.63 ;
      RECT 138.65 -6.52 139 -6.4 ;
      RECT 138.65 -3.29 139 -3.17 ;
      RECT 138.65 -0.06 139 0.06 ;
      RECT 138.765 -104.945 138.865 -103.985 ;
      RECT 138.765 2.175 138.865 3.135 ;
      RECT 138.475 -112.255 138.575 -111.775 ;
      RECT 138.475 -110.765 138.575 -110.295 ;
      RECT 138.165 -100.19 138.515 -100.07 ;
      RECT 138.165 -96.96 138.515 -96.84 ;
      RECT 138.165 -93.73 138.515 -93.61 ;
      RECT 138.165 -90.5 138.515 -90.38 ;
      RECT 138.165 -87.27 138.515 -87.15 ;
      RECT 138.165 -84.04 138.515 -83.92 ;
      RECT 138.165 -80.81 138.515 -80.69 ;
      RECT 138.165 -77.58 138.515 -77.46 ;
      RECT 138.165 -74.35 138.515 -74.23 ;
      RECT 138.165 -71.12 138.515 -71 ;
      RECT 138.165 -67.89 138.515 -67.77 ;
      RECT 138.165 -64.66 138.515 -64.54 ;
      RECT 138.165 -61.43 138.515 -61.31 ;
      RECT 138.165 -58.2 138.515 -58.08 ;
      RECT 138.165 -54.97 138.515 -54.85 ;
      RECT 138.165 -51.74 138.515 -51.62 ;
      RECT 138.165 -48.51 138.515 -48.39 ;
      RECT 138.165 -45.28 138.515 -45.16 ;
      RECT 138.165 -42.05 138.515 -41.93 ;
      RECT 138.165 -38.82 138.515 -38.7 ;
      RECT 138.165 -35.59 138.515 -35.47 ;
      RECT 138.165 -32.36 138.515 -32.24 ;
      RECT 138.165 -29.13 138.515 -29.01 ;
      RECT 138.165 -25.9 138.515 -25.78 ;
      RECT 138.165 -22.67 138.515 -22.55 ;
      RECT 138.165 -19.44 138.515 -19.32 ;
      RECT 138.165 -16.21 138.515 -16.09 ;
      RECT 138.165 -12.98 138.515 -12.86 ;
      RECT 138.165 -9.75 138.515 -9.63 ;
      RECT 138.165 -6.52 138.515 -6.4 ;
      RECT 138.165 -3.29 138.515 -3.17 ;
      RECT 138.165 -0.06 138.515 0.06 ;
      RECT 138.335 -104.945 138.435 -103.985 ;
      RECT 138.335 2.175 138.435 3.135 ;
      RECT 134.435 -108.655 138.215 -108.535 ;
      RECT 138.075 -104.945 138.175 -103.985 ;
      RECT 137.95 -101.06 138.05 -100.525 ;
      RECT 137.95 -99.735 138.05 -99.2 ;
      RECT 137.95 -97.83 138.05 -97.295 ;
      RECT 137.95 -96.505 138.05 -95.97 ;
      RECT 137.95 -94.6 138.05 -94.065 ;
      RECT 137.95 -93.275 138.05 -92.74 ;
      RECT 137.95 -91.37 138.05 -90.835 ;
      RECT 137.95 -90.045 138.05 -89.51 ;
      RECT 137.95 -88.14 138.05 -87.605 ;
      RECT 137.95 -86.815 138.05 -86.28 ;
      RECT 137.95 -84.91 138.05 -84.375 ;
      RECT 137.95 -83.585 138.05 -83.05 ;
      RECT 137.95 -81.68 138.05 -81.145 ;
      RECT 137.95 -80.355 138.05 -79.82 ;
      RECT 137.95 -78.45 138.05 -77.915 ;
      RECT 137.95 -77.125 138.05 -76.59 ;
      RECT 137.95 -75.22 138.05 -74.685 ;
      RECT 137.95 -73.895 138.05 -73.36 ;
      RECT 137.95 -71.99 138.05 -71.455 ;
      RECT 137.95 -70.665 138.05 -70.13 ;
      RECT 137.95 -68.76 138.05 -68.225 ;
      RECT 137.95 -67.435 138.05 -66.9 ;
      RECT 137.95 -65.53 138.05 -64.995 ;
      RECT 137.95 -64.205 138.05 -63.67 ;
      RECT 137.95 -62.3 138.05 -61.765 ;
      RECT 137.95 -60.975 138.05 -60.44 ;
      RECT 137.95 -59.07 138.05 -58.535 ;
      RECT 137.95 -57.745 138.05 -57.21 ;
      RECT 137.95 -55.84 138.05 -55.305 ;
      RECT 137.95 -54.515 138.05 -53.98 ;
      RECT 137.95 -52.61 138.05 -52.075 ;
      RECT 137.95 -51.285 138.05 -50.75 ;
      RECT 137.95 -49.38 138.05 -48.845 ;
      RECT 137.95 -48.055 138.05 -47.52 ;
      RECT 137.95 -46.15 138.05 -45.615 ;
      RECT 137.95 -44.825 138.05 -44.29 ;
      RECT 137.95 -42.92 138.05 -42.385 ;
      RECT 137.95 -41.595 138.05 -41.06 ;
      RECT 137.95 -39.69 138.05 -39.155 ;
      RECT 137.95 -38.365 138.05 -37.83 ;
      RECT 137.95 -36.46 138.05 -35.925 ;
      RECT 137.95 -35.135 138.05 -34.6 ;
      RECT 137.95 -33.23 138.05 -32.695 ;
      RECT 137.95 -31.905 138.05 -31.37 ;
      RECT 137.95 -30 138.05 -29.465 ;
      RECT 137.95 -28.675 138.05 -28.14 ;
      RECT 137.95 -26.77 138.05 -26.235 ;
      RECT 137.95 -25.445 138.05 -24.91 ;
      RECT 137.95 -23.54 138.05 -23.005 ;
      RECT 137.95 -22.215 138.05 -21.68 ;
      RECT 137.95 -20.31 138.05 -19.775 ;
      RECT 137.95 -18.985 138.05 -18.45 ;
      RECT 137.95 -17.08 138.05 -16.545 ;
      RECT 137.95 -15.755 138.05 -15.22 ;
      RECT 137.95 -13.85 138.05 -13.315 ;
      RECT 137.95 -12.525 138.05 -11.99 ;
      RECT 137.95 -10.62 138.05 -10.085 ;
      RECT 137.95 -9.295 138.05 -8.76 ;
      RECT 137.95 -7.39 138.05 -6.855 ;
      RECT 137.95 -6.065 138.05 -5.53 ;
      RECT 137.95 -4.16 138.05 -3.625 ;
      RECT 137.95 -2.835 138.05 -2.3 ;
      RECT 137.95 -0.93 138.05 -0.395 ;
      RECT 137.95 0.395 138.05 0.93 ;
      RECT 137.885 -110.75 138.005 -110.37 ;
      RECT 137.885 -112.245 137.985 -111.775 ;
      RECT 137.825 -104.945 137.925 -103.985 ;
      RECT 137.45 -100.19 137.8 -100.07 ;
      RECT 137.45 -96.96 137.8 -96.84 ;
      RECT 137.45 -93.73 137.8 -93.61 ;
      RECT 137.45 -90.5 137.8 -90.38 ;
      RECT 137.45 -87.27 137.8 -87.15 ;
      RECT 137.45 -84.04 137.8 -83.92 ;
      RECT 137.45 -80.81 137.8 -80.69 ;
      RECT 137.45 -77.58 137.8 -77.46 ;
      RECT 137.45 -74.35 137.8 -74.23 ;
      RECT 137.45 -71.12 137.8 -71 ;
      RECT 137.45 -67.89 137.8 -67.77 ;
      RECT 137.45 -64.66 137.8 -64.54 ;
      RECT 137.45 -61.43 137.8 -61.31 ;
      RECT 137.45 -58.2 137.8 -58.08 ;
      RECT 137.45 -54.97 137.8 -54.85 ;
      RECT 137.45 -51.74 137.8 -51.62 ;
      RECT 137.45 -48.51 137.8 -48.39 ;
      RECT 137.45 -45.28 137.8 -45.16 ;
      RECT 137.45 -42.05 137.8 -41.93 ;
      RECT 137.45 -38.82 137.8 -38.7 ;
      RECT 137.45 -35.59 137.8 -35.47 ;
      RECT 137.45 -32.36 137.8 -32.24 ;
      RECT 137.45 -29.13 137.8 -29.01 ;
      RECT 137.45 -25.9 137.8 -25.78 ;
      RECT 137.45 -22.67 137.8 -22.55 ;
      RECT 137.45 -19.44 137.8 -19.32 ;
      RECT 137.45 -16.21 137.8 -16.09 ;
      RECT 137.45 -12.98 137.8 -12.86 ;
      RECT 137.45 -9.75 137.8 -9.63 ;
      RECT 137.45 -6.52 137.8 -6.4 ;
      RECT 137.45 -3.29 137.8 -3.17 ;
      RECT 137.45 -0.06 137.8 0.06 ;
      RECT 137.565 -104.945 137.665 -103.985 ;
      RECT 137.565 2.175 137.665 3.135 ;
      RECT 137.295 -109.595 137.43 -109.275 ;
      RECT 136.965 -100.19 137.315 -100.07 ;
      RECT 136.965 -96.96 137.315 -96.84 ;
      RECT 136.965 -93.73 137.315 -93.61 ;
      RECT 136.965 -90.5 137.315 -90.38 ;
      RECT 136.965 -87.27 137.315 -87.15 ;
      RECT 136.965 -84.04 137.315 -83.92 ;
      RECT 136.965 -80.81 137.315 -80.69 ;
      RECT 136.965 -77.58 137.315 -77.46 ;
      RECT 136.965 -74.35 137.315 -74.23 ;
      RECT 136.965 -71.12 137.315 -71 ;
      RECT 136.965 -67.89 137.315 -67.77 ;
      RECT 136.965 -64.66 137.315 -64.54 ;
      RECT 136.965 -61.43 137.315 -61.31 ;
      RECT 136.965 -58.2 137.315 -58.08 ;
      RECT 136.965 -54.97 137.315 -54.85 ;
      RECT 136.965 -51.74 137.315 -51.62 ;
      RECT 136.965 -48.51 137.315 -48.39 ;
      RECT 136.965 -45.28 137.315 -45.16 ;
      RECT 136.965 -42.05 137.315 -41.93 ;
      RECT 136.965 -38.82 137.315 -38.7 ;
      RECT 136.965 -35.59 137.315 -35.47 ;
      RECT 136.965 -32.36 137.315 -32.24 ;
      RECT 136.965 -29.13 137.315 -29.01 ;
      RECT 136.965 -25.9 137.315 -25.78 ;
      RECT 136.965 -22.67 137.315 -22.55 ;
      RECT 136.965 -19.44 137.315 -19.32 ;
      RECT 136.965 -16.21 137.315 -16.09 ;
      RECT 136.965 -12.98 137.315 -12.86 ;
      RECT 136.965 -9.75 137.315 -9.63 ;
      RECT 136.965 -6.52 137.315 -6.4 ;
      RECT 136.965 -3.29 137.315 -3.17 ;
      RECT 136.965 -0.06 137.315 0.06 ;
      RECT 137.135 -104.945 137.235 -103.985 ;
      RECT 137.135 2.175 137.235 3.135 ;
      RECT 136.96 -109.595 137.105 -109.275 ;
      RECT 136.875 -104.945 136.975 -103.985 ;
      RECT 136.75 -101.06 136.85 -100.525 ;
      RECT 136.75 -99.735 136.85 -99.2 ;
      RECT 136.75 -97.83 136.85 -97.295 ;
      RECT 136.75 -96.505 136.85 -95.97 ;
      RECT 136.75 -94.6 136.85 -94.065 ;
      RECT 136.75 -93.275 136.85 -92.74 ;
      RECT 136.75 -91.37 136.85 -90.835 ;
      RECT 136.75 -90.045 136.85 -89.51 ;
      RECT 136.75 -88.14 136.85 -87.605 ;
      RECT 136.75 -86.815 136.85 -86.28 ;
      RECT 136.75 -84.91 136.85 -84.375 ;
      RECT 136.75 -83.585 136.85 -83.05 ;
      RECT 136.75 -81.68 136.85 -81.145 ;
      RECT 136.75 -80.355 136.85 -79.82 ;
      RECT 136.75 -78.45 136.85 -77.915 ;
      RECT 136.75 -77.125 136.85 -76.59 ;
      RECT 136.75 -75.22 136.85 -74.685 ;
      RECT 136.75 -73.895 136.85 -73.36 ;
      RECT 136.75 -71.99 136.85 -71.455 ;
      RECT 136.75 -70.665 136.85 -70.13 ;
      RECT 136.75 -68.76 136.85 -68.225 ;
      RECT 136.75 -67.435 136.85 -66.9 ;
      RECT 136.75 -65.53 136.85 -64.995 ;
      RECT 136.75 -64.205 136.85 -63.67 ;
      RECT 136.75 -62.3 136.85 -61.765 ;
      RECT 136.75 -60.975 136.85 -60.44 ;
      RECT 136.75 -59.07 136.85 -58.535 ;
      RECT 136.75 -57.745 136.85 -57.21 ;
      RECT 136.75 -55.84 136.85 -55.305 ;
      RECT 136.75 -54.515 136.85 -53.98 ;
      RECT 136.75 -52.61 136.85 -52.075 ;
      RECT 136.75 -51.285 136.85 -50.75 ;
      RECT 136.75 -49.38 136.85 -48.845 ;
      RECT 136.75 -48.055 136.85 -47.52 ;
      RECT 136.75 -46.15 136.85 -45.615 ;
      RECT 136.75 -44.825 136.85 -44.29 ;
      RECT 136.75 -42.92 136.85 -42.385 ;
      RECT 136.75 -41.595 136.85 -41.06 ;
      RECT 136.75 -39.69 136.85 -39.155 ;
      RECT 136.75 -38.365 136.85 -37.83 ;
      RECT 136.75 -36.46 136.85 -35.925 ;
      RECT 136.75 -35.135 136.85 -34.6 ;
      RECT 136.75 -33.23 136.85 -32.695 ;
      RECT 136.75 -31.905 136.85 -31.37 ;
      RECT 136.75 -30 136.85 -29.465 ;
      RECT 136.75 -28.675 136.85 -28.14 ;
      RECT 136.75 -26.77 136.85 -26.235 ;
      RECT 136.75 -25.445 136.85 -24.91 ;
      RECT 136.75 -23.54 136.85 -23.005 ;
      RECT 136.75 -22.215 136.85 -21.68 ;
      RECT 136.75 -20.31 136.85 -19.775 ;
      RECT 136.75 -18.985 136.85 -18.45 ;
      RECT 136.75 -17.08 136.85 -16.545 ;
      RECT 136.75 -15.755 136.85 -15.22 ;
      RECT 136.75 -13.85 136.85 -13.315 ;
      RECT 136.75 -12.525 136.85 -11.99 ;
      RECT 136.75 -10.62 136.85 -10.085 ;
      RECT 136.75 -9.295 136.85 -8.76 ;
      RECT 136.75 -7.39 136.85 -6.855 ;
      RECT 136.75 -6.065 136.85 -5.53 ;
      RECT 136.75 -4.16 136.85 -3.625 ;
      RECT 136.75 -2.835 136.85 -2.3 ;
      RECT 136.75 -0.93 136.85 -0.395 ;
      RECT 136.75 0.395 136.85 0.93 ;
      RECT 136.625 -108.175 136.725 -107.215 ;
      RECT 136.25 -100.19 136.6 -100.07 ;
      RECT 136.25 -96.96 136.6 -96.84 ;
      RECT 136.25 -93.73 136.6 -93.61 ;
      RECT 136.25 -90.5 136.6 -90.38 ;
      RECT 136.25 -87.27 136.6 -87.15 ;
      RECT 136.25 -84.04 136.6 -83.92 ;
      RECT 136.25 -80.81 136.6 -80.69 ;
      RECT 136.25 -77.58 136.6 -77.46 ;
      RECT 136.25 -74.35 136.6 -74.23 ;
      RECT 136.25 -71.12 136.6 -71 ;
      RECT 136.25 -67.89 136.6 -67.77 ;
      RECT 136.25 -64.66 136.6 -64.54 ;
      RECT 136.25 -61.43 136.6 -61.31 ;
      RECT 136.25 -58.2 136.6 -58.08 ;
      RECT 136.25 -54.97 136.6 -54.85 ;
      RECT 136.25 -51.74 136.6 -51.62 ;
      RECT 136.25 -48.51 136.6 -48.39 ;
      RECT 136.25 -45.28 136.6 -45.16 ;
      RECT 136.25 -42.05 136.6 -41.93 ;
      RECT 136.25 -38.82 136.6 -38.7 ;
      RECT 136.25 -35.59 136.6 -35.47 ;
      RECT 136.25 -32.36 136.6 -32.24 ;
      RECT 136.25 -29.13 136.6 -29.01 ;
      RECT 136.25 -25.9 136.6 -25.78 ;
      RECT 136.25 -22.67 136.6 -22.55 ;
      RECT 136.25 -19.44 136.6 -19.32 ;
      RECT 136.25 -16.21 136.6 -16.09 ;
      RECT 136.25 -12.98 136.6 -12.86 ;
      RECT 136.25 -9.75 136.6 -9.63 ;
      RECT 136.25 -6.52 136.6 -6.4 ;
      RECT 136.25 -3.29 136.6 -3.17 ;
      RECT 136.25 -0.06 136.6 0.06 ;
      RECT 136.455 -112.255 136.555 -111.775 ;
      RECT 136.455 -110.765 136.555 -110.295 ;
      RECT 136.365 -108.175 136.465 -107.215 ;
      RECT 136.365 2.175 136.465 3.135 ;
      RECT 135.765 -100.19 136.115 -100.07 ;
      RECT 135.765 -96.96 136.115 -96.84 ;
      RECT 135.765 -93.73 136.115 -93.61 ;
      RECT 135.765 -90.5 136.115 -90.38 ;
      RECT 135.765 -87.27 136.115 -87.15 ;
      RECT 135.765 -84.04 136.115 -83.92 ;
      RECT 135.765 -80.81 136.115 -80.69 ;
      RECT 135.765 -77.58 136.115 -77.46 ;
      RECT 135.765 -74.35 136.115 -74.23 ;
      RECT 135.765 -71.12 136.115 -71 ;
      RECT 135.765 -67.89 136.115 -67.77 ;
      RECT 135.765 -64.66 136.115 -64.54 ;
      RECT 135.765 -61.43 136.115 -61.31 ;
      RECT 135.765 -58.2 136.115 -58.08 ;
      RECT 135.765 -54.97 136.115 -54.85 ;
      RECT 135.765 -51.74 136.115 -51.62 ;
      RECT 135.765 -48.51 136.115 -48.39 ;
      RECT 135.765 -45.28 136.115 -45.16 ;
      RECT 135.765 -42.05 136.115 -41.93 ;
      RECT 135.765 -38.82 136.115 -38.7 ;
      RECT 135.765 -35.59 136.115 -35.47 ;
      RECT 135.765 -32.36 136.115 -32.24 ;
      RECT 135.765 -29.13 136.115 -29.01 ;
      RECT 135.765 -25.9 136.115 -25.78 ;
      RECT 135.765 -22.67 136.115 -22.55 ;
      RECT 135.765 -19.44 136.115 -19.32 ;
      RECT 135.765 -16.21 136.115 -16.09 ;
      RECT 135.765 -12.98 136.115 -12.86 ;
      RECT 135.765 -9.75 136.115 -9.63 ;
      RECT 135.765 -6.52 136.115 -6.4 ;
      RECT 135.765 -3.29 136.115 -3.17 ;
      RECT 135.765 -0.06 136.115 0.06 ;
      RECT 135.935 -108.175 136.035 -107.215 ;
      RECT 135.935 2.175 136.035 3.135 ;
      RECT 135.83 -110.765 136 -110.385 ;
      RECT 135.865 -112.245 135.965 -111.775 ;
      RECT 135.675 -108.175 135.775 -107.215 ;
      RECT 135.55 -101.06 135.65 -100.525 ;
      RECT 135.55 -99.735 135.65 -99.2 ;
      RECT 135.55 -97.83 135.65 -97.295 ;
      RECT 135.55 -96.505 135.65 -95.97 ;
      RECT 135.55 -94.6 135.65 -94.065 ;
      RECT 135.55 -93.275 135.65 -92.74 ;
      RECT 135.55 -91.37 135.65 -90.835 ;
      RECT 135.55 -90.045 135.65 -89.51 ;
      RECT 135.55 -88.14 135.65 -87.605 ;
      RECT 135.55 -86.815 135.65 -86.28 ;
      RECT 135.55 -84.91 135.65 -84.375 ;
      RECT 135.55 -83.585 135.65 -83.05 ;
      RECT 135.55 -81.68 135.65 -81.145 ;
      RECT 135.55 -80.355 135.65 -79.82 ;
      RECT 135.55 -78.45 135.65 -77.915 ;
      RECT 135.55 -77.125 135.65 -76.59 ;
      RECT 135.55 -75.22 135.65 -74.685 ;
      RECT 135.55 -73.895 135.65 -73.36 ;
      RECT 135.55 -71.99 135.65 -71.455 ;
      RECT 135.55 -70.665 135.65 -70.13 ;
      RECT 135.55 -68.76 135.65 -68.225 ;
      RECT 135.55 -67.435 135.65 -66.9 ;
      RECT 135.55 -65.53 135.65 -64.995 ;
      RECT 135.55 -64.205 135.65 -63.67 ;
      RECT 135.55 -62.3 135.65 -61.765 ;
      RECT 135.55 -60.975 135.65 -60.44 ;
      RECT 135.55 -59.07 135.65 -58.535 ;
      RECT 135.55 -57.745 135.65 -57.21 ;
      RECT 135.55 -55.84 135.65 -55.305 ;
      RECT 135.55 -54.515 135.65 -53.98 ;
      RECT 135.55 -52.61 135.65 -52.075 ;
      RECT 135.55 -51.285 135.65 -50.75 ;
      RECT 135.55 -49.38 135.65 -48.845 ;
      RECT 135.55 -48.055 135.65 -47.52 ;
      RECT 135.55 -46.15 135.65 -45.615 ;
      RECT 135.55 -44.825 135.65 -44.29 ;
      RECT 135.55 -42.92 135.65 -42.385 ;
      RECT 135.55 -41.595 135.65 -41.06 ;
      RECT 135.55 -39.69 135.65 -39.155 ;
      RECT 135.55 -38.365 135.65 -37.83 ;
      RECT 135.55 -36.46 135.65 -35.925 ;
      RECT 135.55 -35.135 135.65 -34.6 ;
      RECT 135.55 -33.23 135.65 -32.695 ;
      RECT 135.55 -31.905 135.65 -31.37 ;
      RECT 135.55 -30 135.65 -29.465 ;
      RECT 135.55 -28.675 135.65 -28.14 ;
      RECT 135.55 -26.77 135.65 -26.235 ;
      RECT 135.55 -25.445 135.65 -24.91 ;
      RECT 135.55 -23.54 135.65 -23.005 ;
      RECT 135.55 -22.215 135.65 -21.68 ;
      RECT 135.55 -20.31 135.65 -19.775 ;
      RECT 135.55 -18.985 135.65 -18.45 ;
      RECT 135.55 -17.08 135.65 -16.545 ;
      RECT 135.55 -15.755 135.65 -15.22 ;
      RECT 135.55 -13.85 135.65 -13.315 ;
      RECT 135.55 -12.525 135.65 -11.99 ;
      RECT 135.55 -10.62 135.65 -10.085 ;
      RECT 135.55 -9.295 135.65 -8.76 ;
      RECT 135.55 -7.39 135.65 -6.855 ;
      RECT 135.55 -6.065 135.65 -5.53 ;
      RECT 135.55 -4.16 135.65 -3.625 ;
      RECT 135.55 -2.835 135.65 -2.3 ;
      RECT 135.55 -0.93 135.65 -0.395 ;
      RECT 135.55 0.395 135.65 0.93 ;
      RECT 135.425 -108.175 135.525 -107.215 ;
      RECT 135.05 -100.19 135.4 -100.07 ;
      RECT 135.05 -96.96 135.4 -96.84 ;
      RECT 135.05 -93.73 135.4 -93.61 ;
      RECT 135.05 -90.5 135.4 -90.38 ;
      RECT 135.05 -87.27 135.4 -87.15 ;
      RECT 135.05 -84.04 135.4 -83.92 ;
      RECT 135.05 -80.81 135.4 -80.69 ;
      RECT 135.05 -77.58 135.4 -77.46 ;
      RECT 135.05 -74.35 135.4 -74.23 ;
      RECT 135.05 -71.12 135.4 -71 ;
      RECT 135.05 -67.89 135.4 -67.77 ;
      RECT 135.05 -64.66 135.4 -64.54 ;
      RECT 135.05 -61.43 135.4 -61.31 ;
      RECT 135.05 -58.2 135.4 -58.08 ;
      RECT 135.05 -54.97 135.4 -54.85 ;
      RECT 135.05 -51.74 135.4 -51.62 ;
      RECT 135.05 -48.51 135.4 -48.39 ;
      RECT 135.05 -45.28 135.4 -45.16 ;
      RECT 135.05 -42.05 135.4 -41.93 ;
      RECT 135.05 -38.82 135.4 -38.7 ;
      RECT 135.05 -35.59 135.4 -35.47 ;
      RECT 135.05 -32.36 135.4 -32.24 ;
      RECT 135.05 -29.13 135.4 -29.01 ;
      RECT 135.05 -25.9 135.4 -25.78 ;
      RECT 135.05 -22.67 135.4 -22.55 ;
      RECT 135.05 -19.44 135.4 -19.32 ;
      RECT 135.05 -16.21 135.4 -16.09 ;
      RECT 135.05 -12.98 135.4 -12.86 ;
      RECT 135.05 -9.75 135.4 -9.63 ;
      RECT 135.05 -6.52 135.4 -6.4 ;
      RECT 135.05 -3.29 135.4 -3.17 ;
      RECT 135.05 -0.06 135.4 0.06 ;
      RECT 135.165 -108.175 135.265 -107.215 ;
      RECT 135.165 2.175 135.265 3.135 ;
      RECT 135.065 -113.555 135.165 -113.085 ;
      RECT 134.565 -100.19 134.915 -100.07 ;
      RECT 134.565 -96.96 134.915 -96.84 ;
      RECT 134.565 -93.73 134.915 -93.61 ;
      RECT 134.565 -90.5 134.915 -90.38 ;
      RECT 134.565 -87.27 134.915 -87.15 ;
      RECT 134.565 -84.04 134.915 -83.92 ;
      RECT 134.565 -80.81 134.915 -80.69 ;
      RECT 134.565 -77.58 134.915 -77.46 ;
      RECT 134.565 -74.35 134.915 -74.23 ;
      RECT 134.565 -71.12 134.915 -71 ;
      RECT 134.565 -67.89 134.915 -67.77 ;
      RECT 134.565 -64.66 134.915 -64.54 ;
      RECT 134.565 -61.43 134.915 -61.31 ;
      RECT 134.565 -58.2 134.915 -58.08 ;
      RECT 134.565 -54.97 134.915 -54.85 ;
      RECT 134.565 -51.74 134.915 -51.62 ;
      RECT 134.565 -48.51 134.915 -48.39 ;
      RECT 134.565 -45.28 134.915 -45.16 ;
      RECT 134.565 -42.05 134.915 -41.93 ;
      RECT 134.565 -38.82 134.915 -38.7 ;
      RECT 134.565 -35.59 134.915 -35.47 ;
      RECT 134.565 -32.36 134.915 -32.24 ;
      RECT 134.565 -29.13 134.915 -29.01 ;
      RECT 134.565 -25.9 134.915 -25.78 ;
      RECT 134.565 -22.67 134.915 -22.55 ;
      RECT 134.565 -19.44 134.915 -19.32 ;
      RECT 134.565 -16.21 134.915 -16.09 ;
      RECT 134.565 -12.98 134.915 -12.86 ;
      RECT 134.565 -9.75 134.915 -9.63 ;
      RECT 134.565 -6.52 134.915 -6.4 ;
      RECT 134.565 -3.29 134.915 -3.17 ;
      RECT 134.565 -0.06 134.915 0.06 ;
      RECT 134.7 -110.735 134.85 -110.445 ;
      RECT 134.735 -108.175 134.835 -107.215 ;
      RECT 134.735 2.175 134.835 3.135 ;
      RECT 134.715 -112.19 134.815 -111.65 ;
      RECT 134.475 -113.555 134.575 -113.085 ;
      RECT 134.475 -108.175 134.575 -107.215 ;
      RECT 134.35 -101.06 134.45 -100.525 ;
      RECT 134.35 -99.735 134.45 -99.2 ;
      RECT 134.35 -97.83 134.45 -97.295 ;
      RECT 134.35 -96.505 134.45 -95.97 ;
      RECT 134.35 -94.6 134.45 -94.065 ;
      RECT 134.35 -93.275 134.45 -92.74 ;
      RECT 134.35 -91.37 134.45 -90.835 ;
      RECT 134.35 -90.045 134.45 -89.51 ;
      RECT 134.35 -88.14 134.45 -87.605 ;
      RECT 134.35 -86.815 134.45 -86.28 ;
      RECT 134.35 -84.91 134.45 -84.375 ;
      RECT 134.35 -83.585 134.45 -83.05 ;
      RECT 134.35 -81.68 134.45 -81.145 ;
      RECT 134.35 -80.355 134.45 -79.82 ;
      RECT 134.35 -78.45 134.45 -77.915 ;
      RECT 134.35 -77.125 134.45 -76.59 ;
      RECT 134.35 -75.22 134.45 -74.685 ;
      RECT 134.35 -73.895 134.45 -73.36 ;
      RECT 134.35 -71.99 134.45 -71.455 ;
      RECT 134.35 -70.665 134.45 -70.13 ;
      RECT 134.35 -68.76 134.45 -68.225 ;
      RECT 134.35 -67.435 134.45 -66.9 ;
      RECT 134.35 -65.53 134.45 -64.995 ;
      RECT 134.35 -64.205 134.45 -63.67 ;
      RECT 134.35 -62.3 134.45 -61.765 ;
      RECT 134.35 -60.975 134.45 -60.44 ;
      RECT 134.35 -59.07 134.45 -58.535 ;
      RECT 134.35 -57.745 134.45 -57.21 ;
      RECT 134.35 -55.84 134.45 -55.305 ;
      RECT 134.35 -54.515 134.45 -53.98 ;
      RECT 134.35 -52.61 134.45 -52.075 ;
      RECT 134.35 -51.285 134.45 -50.75 ;
      RECT 134.35 -49.38 134.45 -48.845 ;
      RECT 134.35 -48.055 134.45 -47.52 ;
      RECT 134.35 -46.15 134.45 -45.615 ;
      RECT 134.35 -44.825 134.45 -44.29 ;
      RECT 134.35 -42.92 134.45 -42.385 ;
      RECT 134.35 -41.595 134.45 -41.06 ;
      RECT 134.35 -39.69 134.45 -39.155 ;
      RECT 134.35 -38.365 134.45 -37.83 ;
      RECT 134.35 -36.46 134.45 -35.925 ;
      RECT 134.35 -35.135 134.45 -34.6 ;
      RECT 134.35 -33.23 134.45 -32.695 ;
      RECT 134.35 -31.905 134.45 -31.37 ;
      RECT 134.35 -30 134.45 -29.465 ;
      RECT 134.35 -28.675 134.45 -28.14 ;
      RECT 134.35 -26.77 134.45 -26.235 ;
      RECT 134.35 -25.445 134.45 -24.91 ;
      RECT 134.35 -23.54 134.45 -23.005 ;
      RECT 134.35 -22.215 134.45 -21.68 ;
      RECT 134.35 -20.31 134.45 -19.775 ;
      RECT 134.35 -18.985 134.45 -18.45 ;
      RECT 134.35 -17.08 134.45 -16.545 ;
      RECT 134.35 -15.755 134.45 -15.22 ;
      RECT 134.35 -13.85 134.45 -13.315 ;
      RECT 134.35 -12.525 134.45 -11.99 ;
      RECT 134.35 -10.62 134.45 -10.085 ;
      RECT 134.35 -9.295 134.45 -8.76 ;
      RECT 134.35 -7.39 134.45 -6.855 ;
      RECT 134.35 -6.065 134.45 -5.53 ;
      RECT 134.35 -4.16 134.45 -3.625 ;
      RECT 134.35 -2.835 134.45 -2.3 ;
      RECT 134.35 -0.93 134.45 -0.395 ;
      RECT 134.35 0.395 134.45 0.93 ;
      RECT 134.225 -104.945 134.325 -103.985 ;
      RECT 133.85 -100.19 134.2 -100.07 ;
      RECT 133.85 -96.96 134.2 -96.84 ;
      RECT 133.85 -93.73 134.2 -93.61 ;
      RECT 133.85 -90.5 134.2 -90.38 ;
      RECT 133.85 -87.27 134.2 -87.15 ;
      RECT 133.85 -84.04 134.2 -83.92 ;
      RECT 133.85 -80.81 134.2 -80.69 ;
      RECT 133.85 -77.58 134.2 -77.46 ;
      RECT 133.85 -74.35 134.2 -74.23 ;
      RECT 133.85 -71.12 134.2 -71 ;
      RECT 133.85 -67.89 134.2 -67.77 ;
      RECT 133.85 -64.66 134.2 -64.54 ;
      RECT 133.85 -61.43 134.2 -61.31 ;
      RECT 133.85 -58.2 134.2 -58.08 ;
      RECT 133.85 -54.97 134.2 -54.85 ;
      RECT 133.85 -51.74 134.2 -51.62 ;
      RECT 133.85 -48.51 134.2 -48.39 ;
      RECT 133.85 -45.28 134.2 -45.16 ;
      RECT 133.85 -42.05 134.2 -41.93 ;
      RECT 133.85 -38.82 134.2 -38.7 ;
      RECT 133.85 -35.59 134.2 -35.47 ;
      RECT 133.85 -32.36 134.2 -32.24 ;
      RECT 133.85 -29.13 134.2 -29.01 ;
      RECT 133.85 -25.9 134.2 -25.78 ;
      RECT 133.85 -22.67 134.2 -22.55 ;
      RECT 133.85 -19.44 134.2 -19.32 ;
      RECT 133.85 -16.21 134.2 -16.09 ;
      RECT 133.85 -12.98 134.2 -12.86 ;
      RECT 133.85 -9.75 134.2 -9.63 ;
      RECT 133.85 -6.52 134.2 -6.4 ;
      RECT 133.85 -3.29 134.2 -3.17 ;
      RECT 133.85 -0.06 134.2 0.06 ;
      RECT 133.965 -104.945 134.065 -103.985 ;
      RECT 133.965 2.175 134.065 3.135 ;
      RECT 133.675 -112.255 133.775 -111.775 ;
      RECT 133.675 -110.765 133.775 -110.295 ;
      RECT 133.365 -100.19 133.715 -100.07 ;
      RECT 133.365 -96.96 133.715 -96.84 ;
      RECT 133.365 -93.73 133.715 -93.61 ;
      RECT 133.365 -90.5 133.715 -90.38 ;
      RECT 133.365 -87.27 133.715 -87.15 ;
      RECT 133.365 -84.04 133.715 -83.92 ;
      RECT 133.365 -80.81 133.715 -80.69 ;
      RECT 133.365 -77.58 133.715 -77.46 ;
      RECT 133.365 -74.35 133.715 -74.23 ;
      RECT 133.365 -71.12 133.715 -71 ;
      RECT 133.365 -67.89 133.715 -67.77 ;
      RECT 133.365 -64.66 133.715 -64.54 ;
      RECT 133.365 -61.43 133.715 -61.31 ;
      RECT 133.365 -58.2 133.715 -58.08 ;
      RECT 133.365 -54.97 133.715 -54.85 ;
      RECT 133.365 -51.74 133.715 -51.62 ;
      RECT 133.365 -48.51 133.715 -48.39 ;
      RECT 133.365 -45.28 133.715 -45.16 ;
      RECT 133.365 -42.05 133.715 -41.93 ;
      RECT 133.365 -38.82 133.715 -38.7 ;
      RECT 133.365 -35.59 133.715 -35.47 ;
      RECT 133.365 -32.36 133.715 -32.24 ;
      RECT 133.365 -29.13 133.715 -29.01 ;
      RECT 133.365 -25.9 133.715 -25.78 ;
      RECT 133.365 -22.67 133.715 -22.55 ;
      RECT 133.365 -19.44 133.715 -19.32 ;
      RECT 133.365 -16.21 133.715 -16.09 ;
      RECT 133.365 -12.98 133.715 -12.86 ;
      RECT 133.365 -9.75 133.715 -9.63 ;
      RECT 133.365 -6.52 133.715 -6.4 ;
      RECT 133.365 -3.29 133.715 -3.17 ;
      RECT 133.365 -0.06 133.715 0.06 ;
      RECT 133.535 -104.945 133.635 -103.985 ;
      RECT 133.535 2.175 133.635 3.135 ;
      RECT 129.635 -108.655 133.415 -108.535 ;
      RECT 133.275 -104.945 133.375 -103.985 ;
      RECT 133.15 -101.06 133.25 -100.525 ;
      RECT 133.15 -99.735 133.25 -99.2 ;
      RECT 133.15 -97.83 133.25 -97.295 ;
      RECT 133.15 -96.505 133.25 -95.97 ;
      RECT 133.15 -94.6 133.25 -94.065 ;
      RECT 133.15 -93.275 133.25 -92.74 ;
      RECT 133.15 -91.37 133.25 -90.835 ;
      RECT 133.15 -90.045 133.25 -89.51 ;
      RECT 133.15 -88.14 133.25 -87.605 ;
      RECT 133.15 -86.815 133.25 -86.28 ;
      RECT 133.15 -84.91 133.25 -84.375 ;
      RECT 133.15 -83.585 133.25 -83.05 ;
      RECT 133.15 -81.68 133.25 -81.145 ;
      RECT 133.15 -80.355 133.25 -79.82 ;
      RECT 133.15 -78.45 133.25 -77.915 ;
      RECT 133.15 -77.125 133.25 -76.59 ;
      RECT 133.15 -75.22 133.25 -74.685 ;
      RECT 133.15 -73.895 133.25 -73.36 ;
      RECT 133.15 -71.99 133.25 -71.455 ;
      RECT 133.15 -70.665 133.25 -70.13 ;
      RECT 133.15 -68.76 133.25 -68.225 ;
      RECT 133.15 -67.435 133.25 -66.9 ;
      RECT 133.15 -65.53 133.25 -64.995 ;
      RECT 133.15 -64.205 133.25 -63.67 ;
      RECT 133.15 -62.3 133.25 -61.765 ;
      RECT 133.15 -60.975 133.25 -60.44 ;
      RECT 133.15 -59.07 133.25 -58.535 ;
      RECT 133.15 -57.745 133.25 -57.21 ;
      RECT 133.15 -55.84 133.25 -55.305 ;
      RECT 133.15 -54.515 133.25 -53.98 ;
      RECT 133.15 -52.61 133.25 -52.075 ;
      RECT 133.15 -51.285 133.25 -50.75 ;
      RECT 133.15 -49.38 133.25 -48.845 ;
      RECT 133.15 -48.055 133.25 -47.52 ;
      RECT 133.15 -46.15 133.25 -45.615 ;
      RECT 133.15 -44.825 133.25 -44.29 ;
      RECT 133.15 -42.92 133.25 -42.385 ;
      RECT 133.15 -41.595 133.25 -41.06 ;
      RECT 133.15 -39.69 133.25 -39.155 ;
      RECT 133.15 -38.365 133.25 -37.83 ;
      RECT 133.15 -36.46 133.25 -35.925 ;
      RECT 133.15 -35.135 133.25 -34.6 ;
      RECT 133.15 -33.23 133.25 -32.695 ;
      RECT 133.15 -31.905 133.25 -31.37 ;
      RECT 133.15 -30 133.25 -29.465 ;
      RECT 133.15 -28.675 133.25 -28.14 ;
      RECT 133.15 -26.77 133.25 -26.235 ;
      RECT 133.15 -25.445 133.25 -24.91 ;
      RECT 133.15 -23.54 133.25 -23.005 ;
      RECT 133.15 -22.215 133.25 -21.68 ;
      RECT 133.15 -20.31 133.25 -19.775 ;
      RECT 133.15 -18.985 133.25 -18.45 ;
      RECT 133.15 -17.08 133.25 -16.545 ;
      RECT 133.15 -15.755 133.25 -15.22 ;
      RECT 133.15 -13.85 133.25 -13.315 ;
      RECT 133.15 -12.525 133.25 -11.99 ;
      RECT 133.15 -10.62 133.25 -10.085 ;
      RECT 133.15 -9.295 133.25 -8.76 ;
      RECT 133.15 -7.39 133.25 -6.855 ;
      RECT 133.15 -6.065 133.25 -5.53 ;
      RECT 133.15 -4.16 133.25 -3.625 ;
      RECT 133.15 -2.835 133.25 -2.3 ;
      RECT 133.15 -0.93 133.25 -0.395 ;
      RECT 133.15 0.395 133.25 0.93 ;
      RECT 133.085 -110.75 133.205 -110.37 ;
      RECT 133.085 -112.245 133.185 -111.775 ;
      RECT 133.025 -104.945 133.125 -103.985 ;
      RECT 132.65 -100.19 133 -100.07 ;
      RECT 132.65 -96.96 133 -96.84 ;
      RECT 132.65 -93.73 133 -93.61 ;
      RECT 132.65 -90.5 133 -90.38 ;
      RECT 132.65 -87.27 133 -87.15 ;
      RECT 132.65 -84.04 133 -83.92 ;
      RECT 132.65 -80.81 133 -80.69 ;
      RECT 132.65 -77.58 133 -77.46 ;
      RECT 132.65 -74.35 133 -74.23 ;
      RECT 132.65 -71.12 133 -71 ;
      RECT 132.65 -67.89 133 -67.77 ;
      RECT 132.65 -64.66 133 -64.54 ;
      RECT 132.65 -61.43 133 -61.31 ;
      RECT 132.65 -58.2 133 -58.08 ;
      RECT 132.65 -54.97 133 -54.85 ;
      RECT 132.65 -51.74 133 -51.62 ;
      RECT 132.65 -48.51 133 -48.39 ;
      RECT 132.65 -45.28 133 -45.16 ;
      RECT 132.65 -42.05 133 -41.93 ;
      RECT 132.65 -38.82 133 -38.7 ;
      RECT 132.65 -35.59 133 -35.47 ;
      RECT 132.65 -32.36 133 -32.24 ;
      RECT 132.65 -29.13 133 -29.01 ;
      RECT 132.65 -25.9 133 -25.78 ;
      RECT 132.65 -22.67 133 -22.55 ;
      RECT 132.65 -19.44 133 -19.32 ;
      RECT 132.65 -16.21 133 -16.09 ;
      RECT 132.65 -12.98 133 -12.86 ;
      RECT 132.65 -9.75 133 -9.63 ;
      RECT 132.65 -6.52 133 -6.4 ;
      RECT 132.65 -3.29 133 -3.17 ;
      RECT 132.65 -0.06 133 0.06 ;
      RECT 132.765 -104.945 132.865 -103.985 ;
      RECT 132.765 2.175 132.865 3.135 ;
      RECT 132.495 -109.595 132.63 -109.275 ;
      RECT 132.165 -100.19 132.515 -100.07 ;
      RECT 132.165 -96.96 132.515 -96.84 ;
      RECT 132.165 -93.73 132.515 -93.61 ;
      RECT 132.165 -90.5 132.515 -90.38 ;
      RECT 132.165 -87.27 132.515 -87.15 ;
      RECT 132.165 -84.04 132.515 -83.92 ;
      RECT 132.165 -80.81 132.515 -80.69 ;
      RECT 132.165 -77.58 132.515 -77.46 ;
      RECT 132.165 -74.35 132.515 -74.23 ;
      RECT 132.165 -71.12 132.515 -71 ;
      RECT 132.165 -67.89 132.515 -67.77 ;
      RECT 132.165 -64.66 132.515 -64.54 ;
      RECT 132.165 -61.43 132.515 -61.31 ;
      RECT 132.165 -58.2 132.515 -58.08 ;
      RECT 132.165 -54.97 132.515 -54.85 ;
      RECT 132.165 -51.74 132.515 -51.62 ;
      RECT 132.165 -48.51 132.515 -48.39 ;
      RECT 132.165 -45.28 132.515 -45.16 ;
      RECT 132.165 -42.05 132.515 -41.93 ;
      RECT 132.165 -38.82 132.515 -38.7 ;
      RECT 132.165 -35.59 132.515 -35.47 ;
      RECT 132.165 -32.36 132.515 -32.24 ;
      RECT 132.165 -29.13 132.515 -29.01 ;
      RECT 132.165 -25.9 132.515 -25.78 ;
      RECT 132.165 -22.67 132.515 -22.55 ;
      RECT 132.165 -19.44 132.515 -19.32 ;
      RECT 132.165 -16.21 132.515 -16.09 ;
      RECT 132.165 -12.98 132.515 -12.86 ;
      RECT 132.165 -9.75 132.515 -9.63 ;
      RECT 132.165 -6.52 132.515 -6.4 ;
      RECT 132.165 -3.29 132.515 -3.17 ;
      RECT 132.165 -0.06 132.515 0.06 ;
      RECT 132.335 -104.945 132.435 -103.985 ;
      RECT 132.335 2.175 132.435 3.135 ;
      RECT 132.16 -109.595 132.305 -109.275 ;
      RECT 132.075 -104.945 132.175 -103.985 ;
      RECT 131.95 -101.06 132.05 -100.525 ;
      RECT 131.95 -99.735 132.05 -99.2 ;
      RECT 131.95 -97.83 132.05 -97.295 ;
      RECT 131.95 -96.505 132.05 -95.97 ;
      RECT 131.95 -94.6 132.05 -94.065 ;
      RECT 131.95 -93.275 132.05 -92.74 ;
      RECT 131.95 -91.37 132.05 -90.835 ;
      RECT 131.95 -90.045 132.05 -89.51 ;
      RECT 131.95 -88.14 132.05 -87.605 ;
      RECT 131.95 -86.815 132.05 -86.28 ;
      RECT 131.95 -84.91 132.05 -84.375 ;
      RECT 131.95 -83.585 132.05 -83.05 ;
      RECT 131.95 -81.68 132.05 -81.145 ;
      RECT 131.95 -80.355 132.05 -79.82 ;
      RECT 131.95 -78.45 132.05 -77.915 ;
      RECT 131.95 -77.125 132.05 -76.59 ;
      RECT 131.95 -75.22 132.05 -74.685 ;
      RECT 131.95 -73.895 132.05 -73.36 ;
      RECT 131.95 -71.99 132.05 -71.455 ;
      RECT 131.95 -70.665 132.05 -70.13 ;
      RECT 131.95 -68.76 132.05 -68.225 ;
      RECT 131.95 -67.435 132.05 -66.9 ;
      RECT 131.95 -65.53 132.05 -64.995 ;
      RECT 131.95 -64.205 132.05 -63.67 ;
      RECT 131.95 -62.3 132.05 -61.765 ;
      RECT 131.95 -60.975 132.05 -60.44 ;
      RECT 131.95 -59.07 132.05 -58.535 ;
      RECT 131.95 -57.745 132.05 -57.21 ;
      RECT 131.95 -55.84 132.05 -55.305 ;
      RECT 131.95 -54.515 132.05 -53.98 ;
      RECT 131.95 -52.61 132.05 -52.075 ;
      RECT 131.95 -51.285 132.05 -50.75 ;
      RECT 131.95 -49.38 132.05 -48.845 ;
      RECT 131.95 -48.055 132.05 -47.52 ;
      RECT 131.95 -46.15 132.05 -45.615 ;
      RECT 131.95 -44.825 132.05 -44.29 ;
      RECT 131.95 -42.92 132.05 -42.385 ;
      RECT 131.95 -41.595 132.05 -41.06 ;
      RECT 131.95 -39.69 132.05 -39.155 ;
      RECT 131.95 -38.365 132.05 -37.83 ;
      RECT 131.95 -36.46 132.05 -35.925 ;
      RECT 131.95 -35.135 132.05 -34.6 ;
      RECT 131.95 -33.23 132.05 -32.695 ;
      RECT 131.95 -31.905 132.05 -31.37 ;
      RECT 131.95 -30 132.05 -29.465 ;
      RECT 131.95 -28.675 132.05 -28.14 ;
      RECT 131.95 -26.77 132.05 -26.235 ;
      RECT 131.95 -25.445 132.05 -24.91 ;
      RECT 131.95 -23.54 132.05 -23.005 ;
      RECT 131.95 -22.215 132.05 -21.68 ;
      RECT 131.95 -20.31 132.05 -19.775 ;
      RECT 131.95 -18.985 132.05 -18.45 ;
      RECT 131.95 -17.08 132.05 -16.545 ;
      RECT 131.95 -15.755 132.05 -15.22 ;
      RECT 131.95 -13.85 132.05 -13.315 ;
      RECT 131.95 -12.525 132.05 -11.99 ;
      RECT 131.95 -10.62 132.05 -10.085 ;
      RECT 131.95 -9.295 132.05 -8.76 ;
      RECT 131.95 -7.39 132.05 -6.855 ;
      RECT 131.95 -6.065 132.05 -5.53 ;
      RECT 131.95 -4.16 132.05 -3.625 ;
      RECT 131.95 -2.835 132.05 -2.3 ;
      RECT 131.95 -0.93 132.05 -0.395 ;
      RECT 131.95 0.395 132.05 0.93 ;
      RECT 131.825 -108.175 131.925 -107.215 ;
      RECT 131.45 -100.19 131.8 -100.07 ;
      RECT 131.45 -96.96 131.8 -96.84 ;
      RECT 131.45 -93.73 131.8 -93.61 ;
      RECT 131.45 -90.5 131.8 -90.38 ;
      RECT 131.45 -87.27 131.8 -87.15 ;
      RECT 131.45 -84.04 131.8 -83.92 ;
      RECT 131.45 -80.81 131.8 -80.69 ;
      RECT 131.45 -77.58 131.8 -77.46 ;
      RECT 131.45 -74.35 131.8 -74.23 ;
      RECT 131.45 -71.12 131.8 -71 ;
      RECT 131.45 -67.89 131.8 -67.77 ;
      RECT 131.45 -64.66 131.8 -64.54 ;
      RECT 131.45 -61.43 131.8 -61.31 ;
      RECT 131.45 -58.2 131.8 -58.08 ;
      RECT 131.45 -54.97 131.8 -54.85 ;
      RECT 131.45 -51.74 131.8 -51.62 ;
      RECT 131.45 -48.51 131.8 -48.39 ;
      RECT 131.45 -45.28 131.8 -45.16 ;
      RECT 131.45 -42.05 131.8 -41.93 ;
      RECT 131.45 -38.82 131.8 -38.7 ;
      RECT 131.45 -35.59 131.8 -35.47 ;
      RECT 131.45 -32.36 131.8 -32.24 ;
      RECT 131.45 -29.13 131.8 -29.01 ;
      RECT 131.45 -25.9 131.8 -25.78 ;
      RECT 131.45 -22.67 131.8 -22.55 ;
      RECT 131.45 -19.44 131.8 -19.32 ;
      RECT 131.45 -16.21 131.8 -16.09 ;
      RECT 131.45 -12.98 131.8 -12.86 ;
      RECT 131.45 -9.75 131.8 -9.63 ;
      RECT 131.45 -6.52 131.8 -6.4 ;
      RECT 131.45 -3.29 131.8 -3.17 ;
      RECT 131.45 -0.06 131.8 0.06 ;
      RECT 131.655 -112.255 131.755 -111.775 ;
      RECT 131.655 -110.765 131.755 -110.295 ;
      RECT 131.565 -108.175 131.665 -107.215 ;
      RECT 131.565 2.175 131.665 3.135 ;
      RECT 130.965 -100.19 131.315 -100.07 ;
      RECT 130.965 -96.96 131.315 -96.84 ;
      RECT 130.965 -93.73 131.315 -93.61 ;
      RECT 130.965 -90.5 131.315 -90.38 ;
      RECT 130.965 -87.27 131.315 -87.15 ;
      RECT 130.965 -84.04 131.315 -83.92 ;
      RECT 130.965 -80.81 131.315 -80.69 ;
      RECT 130.965 -77.58 131.315 -77.46 ;
      RECT 130.965 -74.35 131.315 -74.23 ;
      RECT 130.965 -71.12 131.315 -71 ;
      RECT 130.965 -67.89 131.315 -67.77 ;
      RECT 130.965 -64.66 131.315 -64.54 ;
      RECT 130.965 -61.43 131.315 -61.31 ;
      RECT 130.965 -58.2 131.315 -58.08 ;
      RECT 130.965 -54.97 131.315 -54.85 ;
      RECT 130.965 -51.74 131.315 -51.62 ;
      RECT 130.965 -48.51 131.315 -48.39 ;
      RECT 130.965 -45.28 131.315 -45.16 ;
      RECT 130.965 -42.05 131.315 -41.93 ;
      RECT 130.965 -38.82 131.315 -38.7 ;
      RECT 130.965 -35.59 131.315 -35.47 ;
      RECT 130.965 -32.36 131.315 -32.24 ;
      RECT 130.965 -29.13 131.315 -29.01 ;
      RECT 130.965 -25.9 131.315 -25.78 ;
      RECT 130.965 -22.67 131.315 -22.55 ;
      RECT 130.965 -19.44 131.315 -19.32 ;
      RECT 130.965 -16.21 131.315 -16.09 ;
      RECT 130.965 -12.98 131.315 -12.86 ;
      RECT 130.965 -9.75 131.315 -9.63 ;
      RECT 130.965 -6.52 131.315 -6.4 ;
      RECT 130.965 -3.29 131.315 -3.17 ;
      RECT 130.965 -0.06 131.315 0.06 ;
      RECT 131.135 -108.175 131.235 -107.215 ;
      RECT 131.135 2.175 131.235 3.135 ;
      RECT 131.03 -110.765 131.2 -110.385 ;
      RECT 131.065 -112.245 131.165 -111.775 ;
      RECT 130.875 -108.175 130.975 -107.215 ;
      RECT 130.75 -101.06 130.85 -100.525 ;
      RECT 130.75 -99.735 130.85 -99.2 ;
      RECT 130.75 -97.83 130.85 -97.295 ;
      RECT 130.75 -96.505 130.85 -95.97 ;
      RECT 130.75 -94.6 130.85 -94.065 ;
      RECT 130.75 -93.275 130.85 -92.74 ;
      RECT 130.75 -91.37 130.85 -90.835 ;
      RECT 130.75 -90.045 130.85 -89.51 ;
      RECT 130.75 -88.14 130.85 -87.605 ;
      RECT 130.75 -86.815 130.85 -86.28 ;
      RECT 130.75 -84.91 130.85 -84.375 ;
      RECT 130.75 -83.585 130.85 -83.05 ;
      RECT 130.75 -81.68 130.85 -81.145 ;
      RECT 130.75 -80.355 130.85 -79.82 ;
      RECT 130.75 -78.45 130.85 -77.915 ;
      RECT 130.75 -77.125 130.85 -76.59 ;
      RECT 130.75 -75.22 130.85 -74.685 ;
      RECT 130.75 -73.895 130.85 -73.36 ;
      RECT 130.75 -71.99 130.85 -71.455 ;
      RECT 130.75 -70.665 130.85 -70.13 ;
      RECT 130.75 -68.76 130.85 -68.225 ;
      RECT 130.75 -67.435 130.85 -66.9 ;
      RECT 130.75 -65.53 130.85 -64.995 ;
      RECT 130.75 -64.205 130.85 -63.67 ;
      RECT 130.75 -62.3 130.85 -61.765 ;
      RECT 130.75 -60.975 130.85 -60.44 ;
      RECT 130.75 -59.07 130.85 -58.535 ;
      RECT 130.75 -57.745 130.85 -57.21 ;
      RECT 130.75 -55.84 130.85 -55.305 ;
      RECT 130.75 -54.515 130.85 -53.98 ;
      RECT 130.75 -52.61 130.85 -52.075 ;
      RECT 130.75 -51.285 130.85 -50.75 ;
      RECT 130.75 -49.38 130.85 -48.845 ;
      RECT 130.75 -48.055 130.85 -47.52 ;
      RECT 130.75 -46.15 130.85 -45.615 ;
      RECT 130.75 -44.825 130.85 -44.29 ;
      RECT 130.75 -42.92 130.85 -42.385 ;
      RECT 130.75 -41.595 130.85 -41.06 ;
      RECT 130.75 -39.69 130.85 -39.155 ;
      RECT 130.75 -38.365 130.85 -37.83 ;
      RECT 130.75 -36.46 130.85 -35.925 ;
      RECT 130.75 -35.135 130.85 -34.6 ;
      RECT 130.75 -33.23 130.85 -32.695 ;
      RECT 130.75 -31.905 130.85 -31.37 ;
      RECT 130.75 -30 130.85 -29.465 ;
      RECT 130.75 -28.675 130.85 -28.14 ;
      RECT 130.75 -26.77 130.85 -26.235 ;
      RECT 130.75 -25.445 130.85 -24.91 ;
      RECT 130.75 -23.54 130.85 -23.005 ;
      RECT 130.75 -22.215 130.85 -21.68 ;
      RECT 130.75 -20.31 130.85 -19.775 ;
      RECT 130.75 -18.985 130.85 -18.45 ;
      RECT 130.75 -17.08 130.85 -16.545 ;
      RECT 130.75 -15.755 130.85 -15.22 ;
      RECT 130.75 -13.85 130.85 -13.315 ;
      RECT 130.75 -12.525 130.85 -11.99 ;
      RECT 130.75 -10.62 130.85 -10.085 ;
      RECT 130.75 -9.295 130.85 -8.76 ;
      RECT 130.75 -7.39 130.85 -6.855 ;
      RECT 130.75 -6.065 130.85 -5.53 ;
      RECT 130.75 -4.16 130.85 -3.625 ;
      RECT 130.75 -2.835 130.85 -2.3 ;
      RECT 130.75 -0.93 130.85 -0.395 ;
      RECT 130.75 0.395 130.85 0.93 ;
      RECT 130.625 -108.175 130.725 -107.215 ;
      RECT 130.25 -100.19 130.6 -100.07 ;
      RECT 130.25 -96.96 130.6 -96.84 ;
      RECT 130.25 -93.73 130.6 -93.61 ;
      RECT 130.25 -90.5 130.6 -90.38 ;
      RECT 130.25 -87.27 130.6 -87.15 ;
      RECT 130.25 -84.04 130.6 -83.92 ;
      RECT 130.25 -80.81 130.6 -80.69 ;
      RECT 130.25 -77.58 130.6 -77.46 ;
      RECT 130.25 -74.35 130.6 -74.23 ;
      RECT 130.25 -71.12 130.6 -71 ;
      RECT 130.25 -67.89 130.6 -67.77 ;
      RECT 130.25 -64.66 130.6 -64.54 ;
      RECT 130.25 -61.43 130.6 -61.31 ;
      RECT 130.25 -58.2 130.6 -58.08 ;
      RECT 130.25 -54.97 130.6 -54.85 ;
      RECT 130.25 -51.74 130.6 -51.62 ;
      RECT 130.25 -48.51 130.6 -48.39 ;
      RECT 130.25 -45.28 130.6 -45.16 ;
      RECT 130.25 -42.05 130.6 -41.93 ;
      RECT 130.25 -38.82 130.6 -38.7 ;
      RECT 130.25 -35.59 130.6 -35.47 ;
      RECT 130.25 -32.36 130.6 -32.24 ;
      RECT 130.25 -29.13 130.6 -29.01 ;
      RECT 130.25 -25.9 130.6 -25.78 ;
      RECT 130.25 -22.67 130.6 -22.55 ;
      RECT 130.25 -19.44 130.6 -19.32 ;
      RECT 130.25 -16.21 130.6 -16.09 ;
      RECT 130.25 -12.98 130.6 -12.86 ;
      RECT 130.25 -9.75 130.6 -9.63 ;
      RECT 130.25 -6.52 130.6 -6.4 ;
      RECT 130.25 -3.29 130.6 -3.17 ;
      RECT 130.25 -0.06 130.6 0.06 ;
      RECT 130.365 -108.175 130.465 -107.215 ;
      RECT 130.365 2.175 130.465 3.135 ;
      RECT 130.265 -113.555 130.365 -113.085 ;
      RECT 129.765 -100.19 130.115 -100.07 ;
      RECT 129.765 -96.96 130.115 -96.84 ;
      RECT 129.765 -93.73 130.115 -93.61 ;
      RECT 129.765 -90.5 130.115 -90.38 ;
      RECT 129.765 -87.27 130.115 -87.15 ;
      RECT 129.765 -84.04 130.115 -83.92 ;
      RECT 129.765 -80.81 130.115 -80.69 ;
      RECT 129.765 -77.58 130.115 -77.46 ;
      RECT 129.765 -74.35 130.115 -74.23 ;
      RECT 129.765 -71.12 130.115 -71 ;
      RECT 129.765 -67.89 130.115 -67.77 ;
      RECT 129.765 -64.66 130.115 -64.54 ;
      RECT 129.765 -61.43 130.115 -61.31 ;
      RECT 129.765 -58.2 130.115 -58.08 ;
      RECT 129.765 -54.97 130.115 -54.85 ;
      RECT 129.765 -51.74 130.115 -51.62 ;
      RECT 129.765 -48.51 130.115 -48.39 ;
      RECT 129.765 -45.28 130.115 -45.16 ;
      RECT 129.765 -42.05 130.115 -41.93 ;
      RECT 129.765 -38.82 130.115 -38.7 ;
      RECT 129.765 -35.59 130.115 -35.47 ;
      RECT 129.765 -32.36 130.115 -32.24 ;
      RECT 129.765 -29.13 130.115 -29.01 ;
      RECT 129.765 -25.9 130.115 -25.78 ;
      RECT 129.765 -22.67 130.115 -22.55 ;
      RECT 129.765 -19.44 130.115 -19.32 ;
      RECT 129.765 -16.21 130.115 -16.09 ;
      RECT 129.765 -12.98 130.115 -12.86 ;
      RECT 129.765 -9.75 130.115 -9.63 ;
      RECT 129.765 -6.52 130.115 -6.4 ;
      RECT 129.765 -3.29 130.115 -3.17 ;
      RECT 129.765 -0.06 130.115 0.06 ;
      RECT 129.9 -110.735 130.05 -110.445 ;
      RECT 129.935 -108.175 130.035 -107.215 ;
      RECT 129.935 2.175 130.035 3.135 ;
      RECT 129.915 -112.19 130.015 -111.65 ;
      RECT 129.675 -113.555 129.775 -113.085 ;
      RECT 129.675 -108.175 129.775 -107.215 ;
      RECT 129.55 -101.06 129.65 -100.525 ;
      RECT 129.55 -99.735 129.65 -99.2 ;
      RECT 129.55 -97.83 129.65 -97.295 ;
      RECT 129.55 -96.505 129.65 -95.97 ;
      RECT 129.55 -94.6 129.65 -94.065 ;
      RECT 129.55 -93.275 129.65 -92.74 ;
      RECT 129.55 -91.37 129.65 -90.835 ;
      RECT 129.55 -90.045 129.65 -89.51 ;
      RECT 129.55 -88.14 129.65 -87.605 ;
      RECT 129.55 -86.815 129.65 -86.28 ;
      RECT 129.55 -84.91 129.65 -84.375 ;
      RECT 129.55 -83.585 129.65 -83.05 ;
      RECT 129.55 -81.68 129.65 -81.145 ;
      RECT 129.55 -80.355 129.65 -79.82 ;
      RECT 129.55 -78.45 129.65 -77.915 ;
      RECT 129.55 -77.125 129.65 -76.59 ;
      RECT 129.55 -75.22 129.65 -74.685 ;
      RECT 129.55 -73.895 129.65 -73.36 ;
      RECT 129.55 -71.99 129.65 -71.455 ;
      RECT 129.55 -70.665 129.65 -70.13 ;
      RECT 129.55 -68.76 129.65 -68.225 ;
      RECT 129.55 -67.435 129.65 -66.9 ;
      RECT 129.55 -65.53 129.65 -64.995 ;
      RECT 129.55 -64.205 129.65 -63.67 ;
      RECT 129.55 -62.3 129.65 -61.765 ;
      RECT 129.55 -60.975 129.65 -60.44 ;
      RECT 129.55 -59.07 129.65 -58.535 ;
      RECT 129.55 -57.745 129.65 -57.21 ;
      RECT 129.55 -55.84 129.65 -55.305 ;
      RECT 129.55 -54.515 129.65 -53.98 ;
      RECT 129.55 -52.61 129.65 -52.075 ;
      RECT 129.55 -51.285 129.65 -50.75 ;
      RECT 129.55 -49.38 129.65 -48.845 ;
      RECT 129.55 -48.055 129.65 -47.52 ;
      RECT 129.55 -46.15 129.65 -45.615 ;
      RECT 129.55 -44.825 129.65 -44.29 ;
      RECT 129.55 -42.92 129.65 -42.385 ;
      RECT 129.55 -41.595 129.65 -41.06 ;
      RECT 129.55 -39.69 129.65 -39.155 ;
      RECT 129.55 -38.365 129.65 -37.83 ;
      RECT 129.55 -36.46 129.65 -35.925 ;
      RECT 129.55 -35.135 129.65 -34.6 ;
      RECT 129.55 -33.23 129.65 -32.695 ;
      RECT 129.55 -31.905 129.65 -31.37 ;
      RECT 129.55 -30 129.65 -29.465 ;
      RECT 129.55 -28.675 129.65 -28.14 ;
      RECT 129.55 -26.77 129.65 -26.235 ;
      RECT 129.55 -25.445 129.65 -24.91 ;
      RECT 129.55 -23.54 129.65 -23.005 ;
      RECT 129.55 -22.215 129.65 -21.68 ;
      RECT 129.55 -20.31 129.65 -19.775 ;
      RECT 129.55 -18.985 129.65 -18.45 ;
      RECT 129.55 -17.08 129.65 -16.545 ;
      RECT 129.55 -15.755 129.65 -15.22 ;
      RECT 129.55 -13.85 129.65 -13.315 ;
      RECT 129.55 -12.525 129.65 -11.99 ;
      RECT 129.55 -10.62 129.65 -10.085 ;
      RECT 129.55 -9.295 129.65 -8.76 ;
      RECT 129.55 -7.39 129.65 -6.855 ;
      RECT 129.55 -6.065 129.65 -5.53 ;
      RECT 129.55 -4.16 129.65 -3.625 ;
      RECT 129.55 -2.835 129.65 -2.3 ;
      RECT 129.55 -0.93 129.65 -0.395 ;
      RECT 129.55 0.395 129.65 0.93 ;
      RECT 129.425 -104.945 129.525 -103.985 ;
      RECT 129.05 -100.19 129.4 -100.07 ;
      RECT 129.05 -96.96 129.4 -96.84 ;
      RECT 129.05 -93.73 129.4 -93.61 ;
      RECT 129.05 -90.5 129.4 -90.38 ;
      RECT 129.05 -87.27 129.4 -87.15 ;
      RECT 129.05 -84.04 129.4 -83.92 ;
      RECT 129.05 -80.81 129.4 -80.69 ;
      RECT 129.05 -77.58 129.4 -77.46 ;
      RECT 129.05 -74.35 129.4 -74.23 ;
      RECT 129.05 -71.12 129.4 -71 ;
      RECT 129.05 -67.89 129.4 -67.77 ;
      RECT 129.05 -64.66 129.4 -64.54 ;
      RECT 129.05 -61.43 129.4 -61.31 ;
      RECT 129.05 -58.2 129.4 -58.08 ;
      RECT 129.05 -54.97 129.4 -54.85 ;
      RECT 129.05 -51.74 129.4 -51.62 ;
      RECT 129.05 -48.51 129.4 -48.39 ;
      RECT 129.05 -45.28 129.4 -45.16 ;
      RECT 129.05 -42.05 129.4 -41.93 ;
      RECT 129.05 -38.82 129.4 -38.7 ;
      RECT 129.05 -35.59 129.4 -35.47 ;
      RECT 129.05 -32.36 129.4 -32.24 ;
      RECT 129.05 -29.13 129.4 -29.01 ;
      RECT 129.05 -25.9 129.4 -25.78 ;
      RECT 129.05 -22.67 129.4 -22.55 ;
      RECT 129.05 -19.44 129.4 -19.32 ;
      RECT 129.05 -16.21 129.4 -16.09 ;
      RECT 129.05 -12.98 129.4 -12.86 ;
      RECT 129.05 -9.75 129.4 -9.63 ;
      RECT 129.05 -6.52 129.4 -6.4 ;
      RECT 129.05 -3.29 129.4 -3.17 ;
      RECT 129.05 -0.06 129.4 0.06 ;
      RECT 129.165 -104.945 129.265 -103.985 ;
      RECT 129.165 2.175 129.265 3.135 ;
      RECT 128.875 -112.255 128.975 -111.775 ;
      RECT 128.875 -110.765 128.975 -110.295 ;
      RECT 128.565 -100.19 128.915 -100.07 ;
      RECT 128.565 -96.96 128.915 -96.84 ;
      RECT 128.565 -93.73 128.915 -93.61 ;
      RECT 128.565 -90.5 128.915 -90.38 ;
      RECT 128.565 -87.27 128.915 -87.15 ;
      RECT 128.565 -84.04 128.915 -83.92 ;
      RECT 128.565 -80.81 128.915 -80.69 ;
      RECT 128.565 -77.58 128.915 -77.46 ;
      RECT 128.565 -74.35 128.915 -74.23 ;
      RECT 128.565 -71.12 128.915 -71 ;
      RECT 128.565 -67.89 128.915 -67.77 ;
      RECT 128.565 -64.66 128.915 -64.54 ;
      RECT 128.565 -61.43 128.915 -61.31 ;
      RECT 128.565 -58.2 128.915 -58.08 ;
      RECT 128.565 -54.97 128.915 -54.85 ;
      RECT 128.565 -51.74 128.915 -51.62 ;
      RECT 128.565 -48.51 128.915 -48.39 ;
      RECT 128.565 -45.28 128.915 -45.16 ;
      RECT 128.565 -42.05 128.915 -41.93 ;
      RECT 128.565 -38.82 128.915 -38.7 ;
      RECT 128.565 -35.59 128.915 -35.47 ;
      RECT 128.565 -32.36 128.915 -32.24 ;
      RECT 128.565 -29.13 128.915 -29.01 ;
      RECT 128.565 -25.9 128.915 -25.78 ;
      RECT 128.565 -22.67 128.915 -22.55 ;
      RECT 128.565 -19.44 128.915 -19.32 ;
      RECT 128.565 -16.21 128.915 -16.09 ;
      RECT 128.565 -12.98 128.915 -12.86 ;
      RECT 128.565 -9.75 128.915 -9.63 ;
      RECT 128.565 -6.52 128.915 -6.4 ;
      RECT 128.565 -3.29 128.915 -3.17 ;
      RECT 128.565 -0.06 128.915 0.06 ;
      RECT 128.735 -104.945 128.835 -103.985 ;
      RECT 128.735 2.175 128.835 3.135 ;
      RECT 124.835 -108.655 128.615 -108.535 ;
      RECT 128.475 -104.945 128.575 -103.985 ;
      RECT 128.35 -101.06 128.45 -100.525 ;
      RECT 128.35 -99.735 128.45 -99.2 ;
      RECT 128.35 -97.83 128.45 -97.295 ;
      RECT 128.35 -96.505 128.45 -95.97 ;
      RECT 128.35 -94.6 128.45 -94.065 ;
      RECT 128.35 -93.275 128.45 -92.74 ;
      RECT 128.35 -91.37 128.45 -90.835 ;
      RECT 128.35 -90.045 128.45 -89.51 ;
      RECT 128.35 -88.14 128.45 -87.605 ;
      RECT 128.35 -86.815 128.45 -86.28 ;
      RECT 128.35 -84.91 128.45 -84.375 ;
      RECT 128.35 -83.585 128.45 -83.05 ;
      RECT 128.35 -81.68 128.45 -81.145 ;
      RECT 128.35 -80.355 128.45 -79.82 ;
      RECT 128.35 -78.45 128.45 -77.915 ;
      RECT 128.35 -77.125 128.45 -76.59 ;
      RECT 128.35 -75.22 128.45 -74.685 ;
      RECT 128.35 -73.895 128.45 -73.36 ;
      RECT 128.35 -71.99 128.45 -71.455 ;
      RECT 128.35 -70.665 128.45 -70.13 ;
      RECT 128.35 -68.76 128.45 -68.225 ;
      RECT 128.35 -67.435 128.45 -66.9 ;
      RECT 128.35 -65.53 128.45 -64.995 ;
      RECT 128.35 -64.205 128.45 -63.67 ;
      RECT 128.35 -62.3 128.45 -61.765 ;
      RECT 128.35 -60.975 128.45 -60.44 ;
      RECT 128.35 -59.07 128.45 -58.535 ;
      RECT 128.35 -57.745 128.45 -57.21 ;
      RECT 128.35 -55.84 128.45 -55.305 ;
      RECT 128.35 -54.515 128.45 -53.98 ;
      RECT 128.35 -52.61 128.45 -52.075 ;
      RECT 128.35 -51.285 128.45 -50.75 ;
      RECT 128.35 -49.38 128.45 -48.845 ;
      RECT 128.35 -48.055 128.45 -47.52 ;
      RECT 128.35 -46.15 128.45 -45.615 ;
      RECT 128.35 -44.825 128.45 -44.29 ;
      RECT 128.35 -42.92 128.45 -42.385 ;
      RECT 128.35 -41.595 128.45 -41.06 ;
      RECT 128.35 -39.69 128.45 -39.155 ;
      RECT 128.35 -38.365 128.45 -37.83 ;
      RECT 128.35 -36.46 128.45 -35.925 ;
      RECT 128.35 -35.135 128.45 -34.6 ;
      RECT 128.35 -33.23 128.45 -32.695 ;
      RECT 128.35 -31.905 128.45 -31.37 ;
      RECT 128.35 -30 128.45 -29.465 ;
      RECT 128.35 -28.675 128.45 -28.14 ;
      RECT 128.35 -26.77 128.45 -26.235 ;
      RECT 128.35 -25.445 128.45 -24.91 ;
      RECT 128.35 -23.54 128.45 -23.005 ;
      RECT 128.35 -22.215 128.45 -21.68 ;
      RECT 128.35 -20.31 128.45 -19.775 ;
      RECT 128.35 -18.985 128.45 -18.45 ;
      RECT 128.35 -17.08 128.45 -16.545 ;
      RECT 128.35 -15.755 128.45 -15.22 ;
      RECT 128.35 -13.85 128.45 -13.315 ;
      RECT 128.35 -12.525 128.45 -11.99 ;
      RECT 128.35 -10.62 128.45 -10.085 ;
      RECT 128.35 -9.295 128.45 -8.76 ;
      RECT 128.35 -7.39 128.45 -6.855 ;
      RECT 128.35 -6.065 128.45 -5.53 ;
      RECT 128.35 -4.16 128.45 -3.625 ;
      RECT 128.35 -2.835 128.45 -2.3 ;
      RECT 128.35 -0.93 128.45 -0.395 ;
      RECT 128.35 0.395 128.45 0.93 ;
      RECT 128.285 -110.75 128.405 -110.37 ;
      RECT 128.285 -112.245 128.385 -111.775 ;
      RECT 128.225 -104.945 128.325 -103.985 ;
      RECT 127.85 -100.19 128.2 -100.07 ;
      RECT 127.85 -96.96 128.2 -96.84 ;
      RECT 127.85 -93.73 128.2 -93.61 ;
      RECT 127.85 -90.5 128.2 -90.38 ;
      RECT 127.85 -87.27 128.2 -87.15 ;
      RECT 127.85 -84.04 128.2 -83.92 ;
      RECT 127.85 -80.81 128.2 -80.69 ;
      RECT 127.85 -77.58 128.2 -77.46 ;
      RECT 127.85 -74.35 128.2 -74.23 ;
      RECT 127.85 -71.12 128.2 -71 ;
      RECT 127.85 -67.89 128.2 -67.77 ;
      RECT 127.85 -64.66 128.2 -64.54 ;
      RECT 127.85 -61.43 128.2 -61.31 ;
      RECT 127.85 -58.2 128.2 -58.08 ;
      RECT 127.85 -54.97 128.2 -54.85 ;
      RECT 127.85 -51.74 128.2 -51.62 ;
      RECT 127.85 -48.51 128.2 -48.39 ;
      RECT 127.85 -45.28 128.2 -45.16 ;
      RECT 127.85 -42.05 128.2 -41.93 ;
      RECT 127.85 -38.82 128.2 -38.7 ;
      RECT 127.85 -35.59 128.2 -35.47 ;
      RECT 127.85 -32.36 128.2 -32.24 ;
      RECT 127.85 -29.13 128.2 -29.01 ;
      RECT 127.85 -25.9 128.2 -25.78 ;
      RECT 127.85 -22.67 128.2 -22.55 ;
      RECT 127.85 -19.44 128.2 -19.32 ;
      RECT 127.85 -16.21 128.2 -16.09 ;
      RECT 127.85 -12.98 128.2 -12.86 ;
      RECT 127.85 -9.75 128.2 -9.63 ;
      RECT 127.85 -6.52 128.2 -6.4 ;
      RECT 127.85 -3.29 128.2 -3.17 ;
      RECT 127.85 -0.06 128.2 0.06 ;
      RECT 127.965 -104.945 128.065 -103.985 ;
      RECT 127.965 2.175 128.065 3.135 ;
      RECT 127.695 -109.595 127.83 -109.275 ;
      RECT 127.365 -100.19 127.715 -100.07 ;
      RECT 127.365 -96.96 127.715 -96.84 ;
      RECT 127.365 -93.73 127.715 -93.61 ;
      RECT 127.365 -90.5 127.715 -90.38 ;
      RECT 127.365 -87.27 127.715 -87.15 ;
      RECT 127.365 -84.04 127.715 -83.92 ;
      RECT 127.365 -80.81 127.715 -80.69 ;
      RECT 127.365 -77.58 127.715 -77.46 ;
      RECT 127.365 -74.35 127.715 -74.23 ;
      RECT 127.365 -71.12 127.715 -71 ;
      RECT 127.365 -67.89 127.715 -67.77 ;
      RECT 127.365 -64.66 127.715 -64.54 ;
      RECT 127.365 -61.43 127.715 -61.31 ;
      RECT 127.365 -58.2 127.715 -58.08 ;
      RECT 127.365 -54.97 127.715 -54.85 ;
      RECT 127.365 -51.74 127.715 -51.62 ;
      RECT 127.365 -48.51 127.715 -48.39 ;
      RECT 127.365 -45.28 127.715 -45.16 ;
      RECT 127.365 -42.05 127.715 -41.93 ;
      RECT 127.365 -38.82 127.715 -38.7 ;
      RECT 127.365 -35.59 127.715 -35.47 ;
      RECT 127.365 -32.36 127.715 -32.24 ;
      RECT 127.365 -29.13 127.715 -29.01 ;
      RECT 127.365 -25.9 127.715 -25.78 ;
      RECT 127.365 -22.67 127.715 -22.55 ;
      RECT 127.365 -19.44 127.715 -19.32 ;
      RECT 127.365 -16.21 127.715 -16.09 ;
      RECT 127.365 -12.98 127.715 -12.86 ;
      RECT 127.365 -9.75 127.715 -9.63 ;
      RECT 127.365 -6.52 127.715 -6.4 ;
      RECT 127.365 -3.29 127.715 -3.17 ;
      RECT 127.365 -0.06 127.715 0.06 ;
      RECT 127.535 -104.945 127.635 -103.985 ;
      RECT 127.535 2.175 127.635 3.135 ;
      RECT 127.36 -109.595 127.505 -109.275 ;
      RECT 127.275 -104.945 127.375 -103.985 ;
      RECT 127.15 -101.06 127.25 -100.525 ;
      RECT 127.15 -99.735 127.25 -99.2 ;
      RECT 127.15 -97.83 127.25 -97.295 ;
      RECT 127.15 -96.505 127.25 -95.97 ;
      RECT 127.15 -94.6 127.25 -94.065 ;
      RECT 127.15 -93.275 127.25 -92.74 ;
      RECT 127.15 -91.37 127.25 -90.835 ;
      RECT 127.15 -90.045 127.25 -89.51 ;
      RECT 127.15 -88.14 127.25 -87.605 ;
      RECT 127.15 -86.815 127.25 -86.28 ;
      RECT 127.15 -84.91 127.25 -84.375 ;
      RECT 127.15 -83.585 127.25 -83.05 ;
      RECT 127.15 -81.68 127.25 -81.145 ;
      RECT 127.15 -80.355 127.25 -79.82 ;
      RECT 127.15 -78.45 127.25 -77.915 ;
      RECT 127.15 -77.125 127.25 -76.59 ;
      RECT 127.15 -75.22 127.25 -74.685 ;
      RECT 127.15 -73.895 127.25 -73.36 ;
      RECT 127.15 -71.99 127.25 -71.455 ;
      RECT 127.15 -70.665 127.25 -70.13 ;
      RECT 127.15 -68.76 127.25 -68.225 ;
      RECT 127.15 -67.435 127.25 -66.9 ;
      RECT 127.15 -65.53 127.25 -64.995 ;
      RECT 127.15 -64.205 127.25 -63.67 ;
      RECT 127.15 -62.3 127.25 -61.765 ;
      RECT 127.15 -60.975 127.25 -60.44 ;
      RECT 127.15 -59.07 127.25 -58.535 ;
      RECT 127.15 -57.745 127.25 -57.21 ;
      RECT 127.15 -55.84 127.25 -55.305 ;
      RECT 127.15 -54.515 127.25 -53.98 ;
      RECT 127.15 -52.61 127.25 -52.075 ;
      RECT 127.15 -51.285 127.25 -50.75 ;
      RECT 127.15 -49.38 127.25 -48.845 ;
      RECT 127.15 -48.055 127.25 -47.52 ;
      RECT 127.15 -46.15 127.25 -45.615 ;
      RECT 127.15 -44.825 127.25 -44.29 ;
      RECT 127.15 -42.92 127.25 -42.385 ;
      RECT 127.15 -41.595 127.25 -41.06 ;
      RECT 127.15 -39.69 127.25 -39.155 ;
      RECT 127.15 -38.365 127.25 -37.83 ;
      RECT 127.15 -36.46 127.25 -35.925 ;
      RECT 127.15 -35.135 127.25 -34.6 ;
      RECT 127.15 -33.23 127.25 -32.695 ;
      RECT 127.15 -31.905 127.25 -31.37 ;
      RECT 127.15 -30 127.25 -29.465 ;
      RECT 127.15 -28.675 127.25 -28.14 ;
      RECT 127.15 -26.77 127.25 -26.235 ;
      RECT 127.15 -25.445 127.25 -24.91 ;
      RECT 127.15 -23.54 127.25 -23.005 ;
      RECT 127.15 -22.215 127.25 -21.68 ;
      RECT 127.15 -20.31 127.25 -19.775 ;
      RECT 127.15 -18.985 127.25 -18.45 ;
      RECT 127.15 -17.08 127.25 -16.545 ;
      RECT 127.15 -15.755 127.25 -15.22 ;
      RECT 127.15 -13.85 127.25 -13.315 ;
      RECT 127.15 -12.525 127.25 -11.99 ;
      RECT 127.15 -10.62 127.25 -10.085 ;
      RECT 127.15 -9.295 127.25 -8.76 ;
      RECT 127.15 -7.39 127.25 -6.855 ;
      RECT 127.15 -6.065 127.25 -5.53 ;
      RECT 127.15 -4.16 127.25 -3.625 ;
      RECT 127.15 -2.835 127.25 -2.3 ;
      RECT 127.15 -0.93 127.25 -0.395 ;
      RECT 127.15 0.395 127.25 0.93 ;
      RECT 127.025 -108.175 127.125 -107.215 ;
      RECT 126.65 -100.19 127 -100.07 ;
      RECT 126.65 -96.96 127 -96.84 ;
      RECT 126.65 -93.73 127 -93.61 ;
      RECT 126.65 -90.5 127 -90.38 ;
      RECT 126.65 -87.27 127 -87.15 ;
      RECT 126.65 -84.04 127 -83.92 ;
      RECT 126.65 -80.81 127 -80.69 ;
      RECT 126.65 -77.58 127 -77.46 ;
      RECT 126.65 -74.35 127 -74.23 ;
      RECT 126.65 -71.12 127 -71 ;
      RECT 126.65 -67.89 127 -67.77 ;
      RECT 126.65 -64.66 127 -64.54 ;
      RECT 126.65 -61.43 127 -61.31 ;
      RECT 126.65 -58.2 127 -58.08 ;
      RECT 126.65 -54.97 127 -54.85 ;
      RECT 126.65 -51.74 127 -51.62 ;
      RECT 126.65 -48.51 127 -48.39 ;
      RECT 126.65 -45.28 127 -45.16 ;
      RECT 126.65 -42.05 127 -41.93 ;
      RECT 126.65 -38.82 127 -38.7 ;
      RECT 126.65 -35.59 127 -35.47 ;
      RECT 126.65 -32.36 127 -32.24 ;
      RECT 126.65 -29.13 127 -29.01 ;
      RECT 126.65 -25.9 127 -25.78 ;
      RECT 126.65 -22.67 127 -22.55 ;
      RECT 126.65 -19.44 127 -19.32 ;
      RECT 126.65 -16.21 127 -16.09 ;
      RECT 126.65 -12.98 127 -12.86 ;
      RECT 126.65 -9.75 127 -9.63 ;
      RECT 126.65 -6.52 127 -6.4 ;
      RECT 126.65 -3.29 127 -3.17 ;
      RECT 126.65 -0.06 127 0.06 ;
      RECT 126.855 -112.255 126.955 -111.775 ;
      RECT 126.855 -110.765 126.955 -110.295 ;
      RECT 126.765 -108.175 126.865 -107.215 ;
      RECT 126.765 2.175 126.865 3.135 ;
      RECT 126.165 -100.19 126.515 -100.07 ;
      RECT 126.165 -96.96 126.515 -96.84 ;
      RECT 126.165 -93.73 126.515 -93.61 ;
      RECT 126.165 -90.5 126.515 -90.38 ;
      RECT 126.165 -87.27 126.515 -87.15 ;
      RECT 126.165 -84.04 126.515 -83.92 ;
      RECT 126.165 -80.81 126.515 -80.69 ;
      RECT 126.165 -77.58 126.515 -77.46 ;
      RECT 126.165 -74.35 126.515 -74.23 ;
      RECT 126.165 -71.12 126.515 -71 ;
      RECT 126.165 -67.89 126.515 -67.77 ;
      RECT 126.165 -64.66 126.515 -64.54 ;
      RECT 126.165 -61.43 126.515 -61.31 ;
      RECT 126.165 -58.2 126.515 -58.08 ;
      RECT 126.165 -54.97 126.515 -54.85 ;
      RECT 126.165 -51.74 126.515 -51.62 ;
      RECT 126.165 -48.51 126.515 -48.39 ;
      RECT 126.165 -45.28 126.515 -45.16 ;
      RECT 126.165 -42.05 126.515 -41.93 ;
      RECT 126.165 -38.82 126.515 -38.7 ;
      RECT 126.165 -35.59 126.515 -35.47 ;
      RECT 126.165 -32.36 126.515 -32.24 ;
      RECT 126.165 -29.13 126.515 -29.01 ;
      RECT 126.165 -25.9 126.515 -25.78 ;
      RECT 126.165 -22.67 126.515 -22.55 ;
      RECT 126.165 -19.44 126.515 -19.32 ;
      RECT 126.165 -16.21 126.515 -16.09 ;
      RECT 126.165 -12.98 126.515 -12.86 ;
      RECT 126.165 -9.75 126.515 -9.63 ;
      RECT 126.165 -6.52 126.515 -6.4 ;
      RECT 126.165 -3.29 126.515 -3.17 ;
      RECT 126.165 -0.06 126.515 0.06 ;
      RECT 126.335 -108.175 126.435 -107.215 ;
      RECT 126.335 2.175 126.435 3.135 ;
      RECT 126.23 -110.765 126.4 -110.385 ;
      RECT 126.265 -112.245 126.365 -111.775 ;
      RECT 126.075 -108.175 126.175 -107.215 ;
      RECT 125.95 -101.06 126.05 -100.525 ;
      RECT 125.95 -99.735 126.05 -99.2 ;
      RECT 125.95 -97.83 126.05 -97.295 ;
      RECT 125.95 -96.505 126.05 -95.97 ;
      RECT 125.95 -94.6 126.05 -94.065 ;
      RECT 125.95 -93.275 126.05 -92.74 ;
      RECT 125.95 -91.37 126.05 -90.835 ;
      RECT 125.95 -90.045 126.05 -89.51 ;
      RECT 125.95 -88.14 126.05 -87.605 ;
      RECT 125.95 -86.815 126.05 -86.28 ;
      RECT 125.95 -84.91 126.05 -84.375 ;
      RECT 125.95 -83.585 126.05 -83.05 ;
      RECT 125.95 -81.68 126.05 -81.145 ;
      RECT 125.95 -80.355 126.05 -79.82 ;
      RECT 125.95 -78.45 126.05 -77.915 ;
      RECT 125.95 -77.125 126.05 -76.59 ;
      RECT 125.95 -75.22 126.05 -74.685 ;
      RECT 125.95 -73.895 126.05 -73.36 ;
      RECT 125.95 -71.99 126.05 -71.455 ;
      RECT 125.95 -70.665 126.05 -70.13 ;
      RECT 125.95 -68.76 126.05 -68.225 ;
      RECT 125.95 -67.435 126.05 -66.9 ;
      RECT 125.95 -65.53 126.05 -64.995 ;
      RECT 125.95 -64.205 126.05 -63.67 ;
      RECT 125.95 -62.3 126.05 -61.765 ;
      RECT 125.95 -60.975 126.05 -60.44 ;
      RECT 125.95 -59.07 126.05 -58.535 ;
      RECT 125.95 -57.745 126.05 -57.21 ;
      RECT 125.95 -55.84 126.05 -55.305 ;
      RECT 125.95 -54.515 126.05 -53.98 ;
      RECT 125.95 -52.61 126.05 -52.075 ;
      RECT 125.95 -51.285 126.05 -50.75 ;
      RECT 125.95 -49.38 126.05 -48.845 ;
      RECT 125.95 -48.055 126.05 -47.52 ;
      RECT 125.95 -46.15 126.05 -45.615 ;
      RECT 125.95 -44.825 126.05 -44.29 ;
      RECT 125.95 -42.92 126.05 -42.385 ;
      RECT 125.95 -41.595 126.05 -41.06 ;
      RECT 125.95 -39.69 126.05 -39.155 ;
      RECT 125.95 -38.365 126.05 -37.83 ;
      RECT 125.95 -36.46 126.05 -35.925 ;
      RECT 125.95 -35.135 126.05 -34.6 ;
      RECT 125.95 -33.23 126.05 -32.695 ;
      RECT 125.95 -31.905 126.05 -31.37 ;
      RECT 125.95 -30 126.05 -29.465 ;
      RECT 125.95 -28.675 126.05 -28.14 ;
      RECT 125.95 -26.77 126.05 -26.235 ;
      RECT 125.95 -25.445 126.05 -24.91 ;
      RECT 125.95 -23.54 126.05 -23.005 ;
      RECT 125.95 -22.215 126.05 -21.68 ;
      RECT 125.95 -20.31 126.05 -19.775 ;
      RECT 125.95 -18.985 126.05 -18.45 ;
      RECT 125.95 -17.08 126.05 -16.545 ;
      RECT 125.95 -15.755 126.05 -15.22 ;
      RECT 125.95 -13.85 126.05 -13.315 ;
      RECT 125.95 -12.525 126.05 -11.99 ;
      RECT 125.95 -10.62 126.05 -10.085 ;
      RECT 125.95 -9.295 126.05 -8.76 ;
      RECT 125.95 -7.39 126.05 -6.855 ;
      RECT 125.95 -6.065 126.05 -5.53 ;
      RECT 125.95 -4.16 126.05 -3.625 ;
      RECT 125.95 -2.835 126.05 -2.3 ;
      RECT 125.95 -0.93 126.05 -0.395 ;
      RECT 125.95 0.395 126.05 0.93 ;
      RECT 125.825 -108.175 125.925 -107.215 ;
      RECT 125.45 -100.19 125.8 -100.07 ;
      RECT 125.45 -96.96 125.8 -96.84 ;
      RECT 125.45 -93.73 125.8 -93.61 ;
      RECT 125.45 -90.5 125.8 -90.38 ;
      RECT 125.45 -87.27 125.8 -87.15 ;
      RECT 125.45 -84.04 125.8 -83.92 ;
      RECT 125.45 -80.81 125.8 -80.69 ;
      RECT 125.45 -77.58 125.8 -77.46 ;
      RECT 125.45 -74.35 125.8 -74.23 ;
      RECT 125.45 -71.12 125.8 -71 ;
      RECT 125.45 -67.89 125.8 -67.77 ;
      RECT 125.45 -64.66 125.8 -64.54 ;
      RECT 125.45 -61.43 125.8 -61.31 ;
      RECT 125.45 -58.2 125.8 -58.08 ;
      RECT 125.45 -54.97 125.8 -54.85 ;
      RECT 125.45 -51.74 125.8 -51.62 ;
      RECT 125.45 -48.51 125.8 -48.39 ;
      RECT 125.45 -45.28 125.8 -45.16 ;
      RECT 125.45 -42.05 125.8 -41.93 ;
      RECT 125.45 -38.82 125.8 -38.7 ;
      RECT 125.45 -35.59 125.8 -35.47 ;
      RECT 125.45 -32.36 125.8 -32.24 ;
      RECT 125.45 -29.13 125.8 -29.01 ;
      RECT 125.45 -25.9 125.8 -25.78 ;
      RECT 125.45 -22.67 125.8 -22.55 ;
      RECT 125.45 -19.44 125.8 -19.32 ;
      RECT 125.45 -16.21 125.8 -16.09 ;
      RECT 125.45 -12.98 125.8 -12.86 ;
      RECT 125.45 -9.75 125.8 -9.63 ;
      RECT 125.45 -6.52 125.8 -6.4 ;
      RECT 125.45 -3.29 125.8 -3.17 ;
      RECT 125.45 -0.06 125.8 0.06 ;
      RECT 125.565 -108.175 125.665 -107.215 ;
      RECT 125.565 2.175 125.665 3.135 ;
      RECT 125.465 -113.555 125.565 -113.085 ;
      RECT 124.965 -100.19 125.315 -100.07 ;
      RECT 124.965 -96.96 125.315 -96.84 ;
      RECT 124.965 -93.73 125.315 -93.61 ;
      RECT 124.965 -90.5 125.315 -90.38 ;
      RECT 124.965 -87.27 125.315 -87.15 ;
      RECT 124.965 -84.04 125.315 -83.92 ;
      RECT 124.965 -80.81 125.315 -80.69 ;
      RECT 124.965 -77.58 125.315 -77.46 ;
      RECT 124.965 -74.35 125.315 -74.23 ;
      RECT 124.965 -71.12 125.315 -71 ;
      RECT 124.965 -67.89 125.315 -67.77 ;
      RECT 124.965 -64.66 125.315 -64.54 ;
      RECT 124.965 -61.43 125.315 -61.31 ;
      RECT 124.965 -58.2 125.315 -58.08 ;
      RECT 124.965 -54.97 125.315 -54.85 ;
      RECT 124.965 -51.74 125.315 -51.62 ;
      RECT 124.965 -48.51 125.315 -48.39 ;
      RECT 124.965 -45.28 125.315 -45.16 ;
      RECT 124.965 -42.05 125.315 -41.93 ;
      RECT 124.965 -38.82 125.315 -38.7 ;
      RECT 124.965 -35.59 125.315 -35.47 ;
      RECT 124.965 -32.36 125.315 -32.24 ;
      RECT 124.965 -29.13 125.315 -29.01 ;
      RECT 124.965 -25.9 125.315 -25.78 ;
      RECT 124.965 -22.67 125.315 -22.55 ;
      RECT 124.965 -19.44 125.315 -19.32 ;
      RECT 124.965 -16.21 125.315 -16.09 ;
      RECT 124.965 -12.98 125.315 -12.86 ;
      RECT 124.965 -9.75 125.315 -9.63 ;
      RECT 124.965 -6.52 125.315 -6.4 ;
      RECT 124.965 -3.29 125.315 -3.17 ;
      RECT 124.965 -0.06 125.315 0.06 ;
      RECT 125.1 -110.735 125.25 -110.445 ;
      RECT 125.135 -108.175 125.235 -107.215 ;
      RECT 125.135 2.175 125.235 3.135 ;
      RECT 125.115 -112.19 125.215 -111.65 ;
      RECT 124.875 -113.555 124.975 -113.085 ;
      RECT 124.875 -108.175 124.975 -107.215 ;
      RECT 124.75 -101.06 124.85 -100.525 ;
      RECT 124.75 -99.735 124.85 -99.2 ;
      RECT 124.75 -97.83 124.85 -97.295 ;
      RECT 124.75 -96.505 124.85 -95.97 ;
      RECT 124.75 -94.6 124.85 -94.065 ;
      RECT 124.75 -93.275 124.85 -92.74 ;
      RECT 124.75 -91.37 124.85 -90.835 ;
      RECT 124.75 -90.045 124.85 -89.51 ;
      RECT 124.75 -88.14 124.85 -87.605 ;
      RECT 124.75 -86.815 124.85 -86.28 ;
      RECT 124.75 -84.91 124.85 -84.375 ;
      RECT 124.75 -83.585 124.85 -83.05 ;
      RECT 124.75 -81.68 124.85 -81.145 ;
      RECT 124.75 -80.355 124.85 -79.82 ;
      RECT 124.75 -78.45 124.85 -77.915 ;
      RECT 124.75 -77.125 124.85 -76.59 ;
      RECT 124.75 -75.22 124.85 -74.685 ;
      RECT 124.75 -73.895 124.85 -73.36 ;
      RECT 124.75 -71.99 124.85 -71.455 ;
      RECT 124.75 -70.665 124.85 -70.13 ;
      RECT 124.75 -68.76 124.85 -68.225 ;
      RECT 124.75 -67.435 124.85 -66.9 ;
      RECT 124.75 -65.53 124.85 -64.995 ;
      RECT 124.75 -64.205 124.85 -63.67 ;
      RECT 124.75 -62.3 124.85 -61.765 ;
      RECT 124.75 -60.975 124.85 -60.44 ;
      RECT 124.75 -59.07 124.85 -58.535 ;
      RECT 124.75 -57.745 124.85 -57.21 ;
      RECT 124.75 -55.84 124.85 -55.305 ;
      RECT 124.75 -54.515 124.85 -53.98 ;
      RECT 124.75 -52.61 124.85 -52.075 ;
      RECT 124.75 -51.285 124.85 -50.75 ;
      RECT 124.75 -49.38 124.85 -48.845 ;
      RECT 124.75 -48.055 124.85 -47.52 ;
      RECT 124.75 -46.15 124.85 -45.615 ;
      RECT 124.75 -44.825 124.85 -44.29 ;
      RECT 124.75 -42.92 124.85 -42.385 ;
      RECT 124.75 -41.595 124.85 -41.06 ;
      RECT 124.75 -39.69 124.85 -39.155 ;
      RECT 124.75 -38.365 124.85 -37.83 ;
      RECT 124.75 -36.46 124.85 -35.925 ;
      RECT 124.75 -35.135 124.85 -34.6 ;
      RECT 124.75 -33.23 124.85 -32.695 ;
      RECT 124.75 -31.905 124.85 -31.37 ;
      RECT 124.75 -30 124.85 -29.465 ;
      RECT 124.75 -28.675 124.85 -28.14 ;
      RECT 124.75 -26.77 124.85 -26.235 ;
      RECT 124.75 -25.445 124.85 -24.91 ;
      RECT 124.75 -23.54 124.85 -23.005 ;
      RECT 124.75 -22.215 124.85 -21.68 ;
      RECT 124.75 -20.31 124.85 -19.775 ;
      RECT 124.75 -18.985 124.85 -18.45 ;
      RECT 124.75 -17.08 124.85 -16.545 ;
      RECT 124.75 -15.755 124.85 -15.22 ;
      RECT 124.75 -13.85 124.85 -13.315 ;
      RECT 124.75 -12.525 124.85 -11.99 ;
      RECT 124.75 -10.62 124.85 -10.085 ;
      RECT 124.75 -9.295 124.85 -8.76 ;
      RECT 124.75 -7.39 124.85 -6.855 ;
      RECT 124.75 -6.065 124.85 -5.53 ;
      RECT 124.75 -4.16 124.85 -3.625 ;
      RECT 124.75 -2.835 124.85 -2.3 ;
      RECT 124.75 -0.93 124.85 -0.395 ;
      RECT 124.75 0.395 124.85 0.93 ;
      RECT 124.625 -104.945 124.725 -103.985 ;
      RECT 124.25 -100.19 124.6 -100.07 ;
      RECT 124.25 -96.96 124.6 -96.84 ;
      RECT 124.25 -93.73 124.6 -93.61 ;
      RECT 124.25 -90.5 124.6 -90.38 ;
      RECT 124.25 -87.27 124.6 -87.15 ;
      RECT 124.25 -84.04 124.6 -83.92 ;
      RECT 124.25 -80.81 124.6 -80.69 ;
      RECT 124.25 -77.58 124.6 -77.46 ;
      RECT 124.25 -74.35 124.6 -74.23 ;
      RECT 124.25 -71.12 124.6 -71 ;
      RECT 124.25 -67.89 124.6 -67.77 ;
      RECT 124.25 -64.66 124.6 -64.54 ;
      RECT 124.25 -61.43 124.6 -61.31 ;
      RECT 124.25 -58.2 124.6 -58.08 ;
      RECT 124.25 -54.97 124.6 -54.85 ;
      RECT 124.25 -51.74 124.6 -51.62 ;
      RECT 124.25 -48.51 124.6 -48.39 ;
      RECT 124.25 -45.28 124.6 -45.16 ;
      RECT 124.25 -42.05 124.6 -41.93 ;
      RECT 124.25 -38.82 124.6 -38.7 ;
      RECT 124.25 -35.59 124.6 -35.47 ;
      RECT 124.25 -32.36 124.6 -32.24 ;
      RECT 124.25 -29.13 124.6 -29.01 ;
      RECT 124.25 -25.9 124.6 -25.78 ;
      RECT 124.25 -22.67 124.6 -22.55 ;
      RECT 124.25 -19.44 124.6 -19.32 ;
      RECT 124.25 -16.21 124.6 -16.09 ;
      RECT 124.25 -12.98 124.6 -12.86 ;
      RECT 124.25 -9.75 124.6 -9.63 ;
      RECT 124.25 -6.52 124.6 -6.4 ;
      RECT 124.25 -3.29 124.6 -3.17 ;
      RECT 124.25 -0.06 124.6 0.06 ;
      RECT 124.365 -104.945 124.465 -103.985 ;
      RECT 124.365 2.175 124.465 3.135 ;
      RECT 124.075 -112.255 124.175 -111.775 ;
      RECT 124.075 -110.765 124.175 -110.295 ;
      RECT 123.765 -100.19 124.115 -100.07 ;
      RECT 123.765 -96.96 124.115 -96.84 ;
      RECT 123.765 -93.73 124.115 -93.61 ;
      RECT 123.765 -90.5 124.115 -90.38 ;
      RECT 123.765 -87.27 124.115 -87.15 ;
      RECT 123.765 -84.04 124.115 -83.92 ;
      RECT 123.765 -80.81 124.115 -80.69 ;
      RECT 123.765 -77.58 124.115 -77.46 ;
      RECT 123.765 -74.35 124.115 -74.23 ;
      RECT 123.765 -71.12 124.115 -71 ;
      RECT 123.765 -67.89 124.115 -67.77 ;
      RECT 123.765 -64.66 124.115 -64.54 ;
      RECT 123.765 -61.43 124.115 -61.31 ;
      RECT 123.765 -58.2 124.115 -58.08 ;
      RECT 123.765 -54.97 124.115 -54.85 ;
      RECT 123.765 -51.74 124.115 -51.62 ;
      RECT 123.765 -48.51 124.115 -48.39 ;
      RECT 123.765 -45.28 124.115 -45.16 ;
      RECT 123.765 -42.05 124.115 -41.93 ;
      RECT 123.765 -38.82 124.115 -38.7 ;
      RECT 123.765 -35.59 124.115 -35.47 ;
      RECT 123.765 -32.36 124.115 -32.24 ;
      RECT 123.765 -29.13 124.115 -29.01 ;
      RECT 123.765 -25.9 124.115 -25.78 ;
      RECT 123.765 -22.67 124.115 -22.55 ;
      RECT 123.765 -19.44 124.115 -19.32 ;
      RECT 123.765 -16.21 124.115 -16.09 ;
      RECT 123.765 -12.98 124.115 -12.86 ;
      RECT 123.765 -9.75 124.115 -9.63 ;
      RECT 123.765 -6.52 124.115 -6.4 ;
      RECT 123.765 -3.29 124.115 -3.17 ;
      RECT 123.765 -0.06 124.115 0.06 ;
      RECT 123.935 -104.945 124.035 -103.985 ;
      RECT 123.935 2.175 124.035 3.135 ;
      RECT 120.035 -108.655 123.815 -108.535 ;
      RECT 123.675 -104.945 123.775 -103.985 ;
      RECT 123.55 -101.06 123.65 -100.525 ;
      RECT 123.55 -99.735 123.65 -99.2 ;
      RECT 123.55 -97.83 123.65 -97.295 ;
      RECT 123.55 -96.505 123.65 -95.97 ;
      RECT 123.55 -94.6 123.65 -94.065 ;
      RECT 123.55 -93.275 123.65 -92.74 ;
      RECT 123.55 -91.37 123.65 -90.835 ;
      RECT 123.55 -90.045 123.65 -89.51 ;
      RECT 123.55 -88.14 123.65 -87.605 ;
      RECT 123.55 -86.815 123.65 -86.28 ;
      RECT 123.55 -84.91 123.65 -84.375 ;
      RECT 123.55 -83.585 123.65 -83.05 ;
      RECT 123.55 -81.68 123.65 -81.145 ;
      RECT 123.55 -80.355 123.65 -79.82 ;
      RECT 123.55 -78.45 123.65 -77.915 ;
      RECT 123.55 -77.125 123.65 -76.59 ;
      RECT 123.55 -75.22 123.65 -74.685 ;
      RECT 123.55 -73.895 123.65 -73.36 ;
      RECT 123.55 -71.99 123.65 -71.455 ;
      RECT 123.55 -70.665 123.65 -70.13 ;
      RECT 123.55 -68.76 123.65 -68.225 ;
      RECT 123.55 -67.435 123.65 -66.9 ;
      RECT 123.55 -65.53 123.65 -64.995 ;
      RECT 123.55 -64.205 123.65 -63.67 ;
      RECT 123.55 -62.3 123.65 -61.765 ;
      RECT 123.55 -60.975 123.65 -60.44 ;
      RECT 123.55 -59.07 123.65 -58.535 ;
      RECT 123.55 -57.745 123.65 -57.21 ;
      RECT 123.55 -55.84 123.65 -55.305 ;
      RECT 123.55 -54.515 123.65 -53.98 ;
      RECT 123.55 -52.61 123.65 -52.075 ;
      RECT 123.55 -51.285 123.65 -50.75 ;
      RECT 123.55 -49.38 123.65 -48.845 ;
      RECT 123.55 -48.055 123.65 -47.52 ;
      RECT 123.55 -46.15 123.65 -45.615 ;
      RECT 123.55 -44.825 123.65 -44.29 ;
      RECT 123.55 -42.92 123.65 -42.385 ;
      RECT 123.55 -41.595 123.65 -41.06 ;
      RECT 123.55 -39.69 123.65 -39.155 ;
      RECT 123.55 -38.365 123.65 -37.83 ;
      RECT 123.55 -36.46 123.65 -35.925 ;
      RECT 123.55 -35.135 123.65 -34.6 ;
      RECT 123.55 -33.23 123.65 -32.695 ;
      RECT 123.55 -31.905 123.65 -31.37 ;
      RECT 123.55 -30 123.65 -29.465 ;
      RECT 123.55 -28.675 123.65 -28.14 ;
      RECT 123.55 -26.77 123.65 -26.235 ;
      RECT 123.55 -25.445 123.65 -24.91 ;
      RECT 123.55 -23.54 123.65 -23.005 ;
      RECT 123.55 -22.215 123.65 -21.68 ;
      RECT 123.55 -20.31 123.65 -19.775 ;
      RECT 123.55 -18.985 123.65 -18.45 ;
      RECT 123.55 -17.08 123.65 -16.545 ;
      RECT 123.55 -15.755 123.65 -15.22 ;
      RECT 123.55 -13.85 123.65 -13.315 ;
      RECT 123.55 -12.525 123.65 -11.99 ;
      RECT 123.55 -10.62 123.65 -10.085 ;
      RECT 123.55 -9.295 123.65 -8.76 ;
      RECT 123.55 -7.39 123.65 -6.855 ;
      RECT 123.55 -6.065 123.65 -5.53 ;
      RECT 123.55 -4.16 123.65 -3.625 ;
      RECT 123.55 -2.835 123.65 -2.3 ;
      RECT 123.55 -0.93 123.65 -0.395 ;
      RECT 123.55 0.395 123.65 0.93 ;
      RECT 123.485 -110.75 123.605 -110.37 ;
      RECT 123.485 -112.245 123.585 -111.775 ;
      RECT 123.425 -104.945 123.525 -103.985 ;
      RECT 123.05 -100.19 123.4 -100.07 ;
      RECT 123.05 -96.96 123.4 -96.84 ;
      RECT 123.05 -93.73 123.4 -93.61 ;
      RECT 123.05 -90.5 123.4 -90.38 ;
      RECT 123.05 -87.27 123.4 -87.15 ;
      RECT 123.05 -84.04 123.4 -83.92 ;
      RECT 123.05 -80.81 123.4 -80.69 ;
      RECT 123.05 -77.58 123.4 -77.46 ;
      RECT 123.05 -74.35 123.4 -74.23 ;
      RECT 123.05 -71.12 123.4 -71 ;
      RECT 123.05 -67.89 123.4 -67.77 ;
      RECT 123.05 -64.66 123.4 -64.54 ;
      RECT 123.05 -61.43 123.4 -61.31 ;
      RECT 123.05 -58.2 123.4 -58.08 ;
      RECT 123.05 -54.97 123.4 -54.85 ;
      RECT 123.05 -51.74 123.4 -51.62 ;
      RECT 123.05 -48.51 123.4 -48.39 ;
      RECT 123.05 -45.28 123.4 -45.16 ;
      RECT 123.05 -42.05 123.4 -41.93 ;
      RECT 123.05 -38.82 123.4 -38.7 ;
      RECT 123.05 -35.59 123.4 -35.47 ;
      RECT 123.05 -32.36 123.4 -32.24 ;
      RECT 123.05 -29.13 123.4 -29.01 ;
      RECT 123.05 -25.9 123.4 -25.78 ;
      RECT 123.05 -22.67 123.4 -22.55 ;
      RECT 123.05 -19.44 123.4 -19.32 ;
      RECT 123.05 -16.21 123.4 -16.09 ;
      RECT 123.05 -12.98 123.4 -12.86 ;
      RECT 123.05 -9.75 123.4 -9.63 ;
      RECT 123.05 -6.52 123.4 -6.4 ;
      RECT 123.05 -3.29 123.4 -3.17 ;
      RECT 123.05 -0.06 123.4 0.06 ;
      RECT 123.165 -104.945 123.265 -103.985 ;
      RECT 123.165 2.175 123.265 3.135 ;
      RECT 122.895 -109.595 123.03 -109.275 ;
      RECT 122.565 -100.19 122.915 -100.07 ;
      RECT 122.565 -96.96 122.915 -96.84 ;
      RECT 122.565 -93.73 122.915 -93.61 ;
      RECT 122.565 -90.5 122.915 -90.38 ;
      RECT 122.565 -87.27 122.915 -87.15 ;
      RECT 122.565 -84.04 122.915 -83.92 ;
      RECT 122.565 -80.81 122.915 -80.69 ;
      RECT 122.565 -77.58 122.915 -77.46 ;
      RECT 122.565 -74.35 122.915 -74.23 ;
      RECT 122.565 -71.12 122.915 -71 ;
      RECT 122.565 -67.89 122.915 -67.77 ;
      RECT 122.565 -64.66 122.915 -64.54 ;
      RECT 122.565 -61.43 122.915 -61.31 ;
      RECT 122.565 -58.2 122.915 -58.08 ;
      RECT 122.565 -54.97 122.915 -54.85 ;
      RECT 122.565 -51.74 122.915 -51.62 ;
      RECT 122.565 -48.51 122.915 -48.39 ;
      RECT 122.565 -45.28 122.915 -45.16 ;
      RECT 122.565 -42.05 122.915 -41.93 ;
      RECT 122.565 -38.82 122.915 -38.7 ;
      RECT 122.565 -35.59 122.915 -35.47 ;
      RECT 122.565 -32.36 122.915 -32.24 ;
      RECT 122.565 -29.13 122.915 -29.01 ;
      RECT 122.565 -25.9 122.915 -25.78 ;
      RECT 122.565 -22.67 122.915 -22.55 ;
      RECT 122.565 -19.44 122.915 -19.32 ;
      RECT 122.565 -16.21 122.915 -16.09 ;
      RECT 122.565 -12.98 122.915 -12.86 ;
      RECT 122.565 -9.75 122.915 -9.63 ;
      RECT 122.565 -6.52 122.915 -6.4 ;
      RECT 122.565 -3.29 122.915 -3.17 ;
      RECT 122.565 -0.06 122.915 0.06 ;
      RECT 122.735 -104.945 122.835 -103.985 ;
      RECT 122.735 2.175 122.835 3.135 ;
      RECT 122.56 -109.595 122.705 -109.275 ;
      RECT 122.475 -104.945 122.575 -103.985 ;
      RECT 122.35 -101.06 122.45 -100.525 ;
      RECT 122.35 -99.735 122.45 -99.2 ;
      RECT 122.35 -97.83 122.45 -97.295 ;
      RECT 122.35 -96.505 122.45 -95.97 ;
      RECT 122.35 -94.6 122.45 -94.065 ;
      RECT 122.35 -93.275 122.45 -92.74 ;
      RECT 122.35 -91.37 122.45 -90.835 ;
      RECT 122.35 -90.045 122.45 -89.51 ;
      RECT 122.35 -88.14 122.45 -87.605 ;
      RECT 122.35 -86.815 122.45 -86.28 ;
      RECT 122.35 -84.91 122.45 -84.375 ;
      RECT 122.35 -83.585 122.45 -83.05 ;
      RECT 122.35 -81.68 122.45 -81.145 ;
      RECT 122.35 -80.355 122.45 -79.82 ;
      RECT 122.35 -78.45 122.45 -77.915 ;
      RECT 122.35 -77.125 122.45 -76.59 ;
      RECT 122.35 -75.22 122.45 -74.685 ;
      RECT 122.35 -73.895 122.45 -73.36 ;
      RECT 122.35 -71.99 122.45 -71.455 ;
      RECT 122.35 -70.665 122.45 -70.13 ;
      RECT 122.35 -68.76 122.45 -68.225 ;
      RECT 122.35 -67.435 122.45 -66.9 ;
      RECT 122.35 -65.53 122.45 -64.995 ;
      RECT 122.35 -64.205 122.45 -63.67 ;
      RECT 122.35 -62.3 122.45 -61.765 ;
      RECT 122.35 -60.975 122.45 -60.44 ;
      RECT 122.35 -59.07 122.45 -58.535 ;
      RECT 122.35 -57.745 122.45 -57.21 ;
      RECT 122.35 -55.84 122.45 -55.305 ;
      RECT 122.35 -54.515 122.45 -53.98 ;
      RECT 122.35 -52.61 122.45 -52.075 ;
      RECT 122.35 -51.285 122.45 -50.75 ;
      RECT 122.35 -49.38 122.45 -48.845 ;
      RECT 122.35 -48.055 122.45 -47.52 ;
      RECT 122.35 -46.15 122.45 -45.615 ;
      RECT 122.35 -44.825 122.45 -44.29 ;
      RECT 122.35 -42.92 122.45 -42.385 ;
      RECT 122.35 -41.595 122.45 -41.06 ;
      RECT 122.35 -39.69 122.45 -39.155 ;
      RECT 122.35 -38.365 122.45 -37.83 ;
      RECT 122.35 -36.46 122.45 -35.925 ;
      RECT 122.35 -35.135 122.45 -34.6 ;
      RECT 122.35 -33.23 122.45 -32.695 ;
      RECT 122.35 -31.905 122.45 -31.37 ;
      RECT 122.35 -30 122.45 -29.465 ;
      RECT 122.35 -28.675 122.45 -28.14 ;
      RECT 122.35 -26.77 122.45 -26.235 ;
      RECT 122.35 -25.445 122.45 -24.91 ;
      RECT 122.35 -23.54 122.45 -23.005 ;
      RECT 122.35 -22.215 122.45 -21.68 ;
      RECT 122.35 -20.31 122.45 -19.775 ;
      RECT 122.35 -18.985 122.45 -18.45 ;
      RECT 122.35 -17.08 122.45 -16.545 ;
      RECT 122.35 -15.755 122.45 -15.22 ;
      RECT 122.35 -13.85 122.45 -13.315 ;
      RECT 122.35 -12.525 122.45 -11.99 ;
      RECT 122.35 -10.62 122.45 -10.085 ;
      RECT 122.35 -9.295 122.45 -8.76 ;
      RECT 122.35 -7.39 122.45 -6.855 ;
      RECT 122.35 -6.065 122.45 -5.53 ;
      RECT 122.35 -4.16 122.45 -3.625 ;
      RECT 122.35 -2.835 122.45 -2.3 ;
      RECT 122.35 -0.93 122.45 -0.395 ;
      RECT 122.35 0.395 122.45 0.93 ;
      RECT 122.225 -108.175 122.325 -107.215 ;
      RECT 121.85 -100.19 122.2 -100.07 ;
      RECT 121.85 -96.96 122.2 -96.84 ;
      RECT 121.85 -93.73 122.2 -93.61 ;
      RECT 121.85 -90.5 122.2 -90.38 ;
      RECT 121.85 -87.27 122.2 -87.15 ;
      RECT 121.85 -84.04 122.2 -83.92 ;
      RECT 121.85 -80.81 122.2 -80.69 ;
      RECT 121.85 -77.58 122.2 -77.46 ;
      RECT 121.85 -74.35 122.2 -74.23 ;
      RECT 121.85 -71.12 122.2 -71 ;
      RECT 121.85 -67.89 122.2 -67.77 ;
      RECT 121.85 -64.66 122.2 -64.54 ;
      RECT 121.85 -61.43 122.2 -61.31 ;
      RECT 121.85 -58.2 122.2 -58.08 ;
      RECT 121.85 -54.97 122.2 -54.85 ;
      RECT 121.85 -51.74 122.2 -51.62 ;
      RECT 121.85 -48.51 122.2 -48.39 ;
      RECT 121.85 -45.28 122.2 -45.16 ;
      RECT 121.85 -42.05 122.2 -41.93 ;
      RECT 121.85 -38.82 122.2 -38.7 ;
      RECT 121.85 -35.59 122.2 -35.47 ;
      RECT 121.85 -32.36 122.2 -32.24 ;
      RECT 121.85 -29.13 122.2 -29.01 ;
      RECT 121.85 -25.9 122.2 -25.78 ;
      RECT 121.85 -22.67 122.2 -22.55 ;
      RECT 121.85 -19.44 122.2 -19.32 ;
      RECT 121.85 -16.21 122.2 -16.09 ;
      RECT 121.85 -12.98 122.2 -12.86 ;
      RECT 121.85 -9.75 122.2 -9.63 ;
      RECT 121.85 -6.52 122.2 -6.4 ;
      RECT 121.85 -3.29 122.2 -3.17 ;
      RECT 121.85 -0.06 122.2 0.06 ;
      RECT 122.055 -112.255 122.155 -111.775 ;
      RECT 122.055 -110.765 122.155 -110.295 ;
      RECT 121.965 -108.175 122.065 -107.215 ;
      RECT 121.965 2.175 122.065 3.135 ;
      RECT 121.365 -100.19 121.715 -100.07 ;
      RECT 121.365 -96.96 121.715 -96.84 ;
      RECT 121.365 -93.73 121.715 -93.61 ;
      RECT 121.365 -90.5 121.715 -90.38 ;
      RECT 121.365 -87.27 121.715 -87.15 ;
      RECT 121.365 -84.04 121.715 -83.92 ;
      RECT 121.365 -80.81 121.715 -80.69 ;
      RECT 121.365 -77.58 121.715 -77.46 ;
      RECT 121.365 -74.35 121.715 -74.23 ;
      RECT 121.365 -71.12 121.715 -71 ;
      RECT 121.365 -67.89 121.715 -67.77 ;
      RECT 121.365 -64.66 121.715 -64.54 ;
      RECT 121.365 -61.43 121.715 -61.31 ;
      RECT 121.365 -58.2 121.715 -58.08 ;
      RECT 121.365 -54.97 121.715 -54.85 ;
      RECT 121.365 -51.74 121.715 -51.62 ;
      RECT 121.365 -48.51 121.715 -48.39 ;
      RECT 121.365 -45.28 121.715 -45.16 ;
      RECT 121.365 -42.05 121.715 -41.93 ;
      RECT 121.365 -38.82 121.715 -38.7 ;
      RECT 121.365 -35.59 121.715 -35.47 ;
      RECT 121.365 -32.36 121.715 -32.24 ;
      RECT 121.365 -29.13 121.715 -29.01 ;
      RECT 121.365 -25.9 121.715 -25.78 ;
      RECT 121.365 -22.67 121.715 -22.55 ;
      RECT 121.365 -19.44 121.715 -19.32 ;
      RECT 121.365 -16.21 121.715 -16.09 ;
      RECT 121.365 -12.98 121.715 -12.86 ;
      RECT 121.365 -9.75 121.715 -9.63 ;
      RECT 121.365 -6.52 121.715 -6.4 ;
      RECT 121.365 -3.29 121.715 -3.17 ;
      RECT 121.365 -0.06 121.715 0.06 ;
      RECT 121.535 -108.175 121.635 -107.215 ;
      RECT 121.535 2.175 121.635 3.135 ;
      RECT 121.43 -110.765 121.6 -110.385 ;
      RECT 121.465 -112.245 121.565 -111.775 ;
      RECT 121.275 -108.175 121.375 -107.215 ;
      RECT 121.15 -101.06 121.25 -100.525 ;
      RECT 121.15 -99.735 121.25 -99.2 ;
      RECT 121.15 -97.83 121.25 -97.295 ;
      RECT 121.15 -96.505 121.25 -95.97 ;
      RECT 121.15 -94.6 121.25 -94.065 ;
      RECT 121.15 -93.275 121.25 -92.74 ;
      RECT 121.15 -91.37 121.25 -90.835 ;
      RECT 121.15 -90.045 121.25 -89.51 ;
      RECT 121.15 -88.14 121.25 -87.605 ;
      RECT 121.15 -86.815 121.25 -86.28 ;
      RECT 121.15 -84.91 121.25 -84.375 ;
      RECT 121.15 -83.585 121.25 -83.05 ;
      RECT 121.15 -81.68 121.25 -81.145 ;
      RECT 121.15 -80.355 121.25 -79.82 ;
      RECT 121.15 -78.45 121.25 -77.915 ;
      RECT 121.15 -77.125 121.25 -76.59 ;
      RECT 121.15 -75.22 121.25 -74.685 ;
      RECT 121.15 -73.895 121.25 -73.36 ;
      RECT 121.15 -71.99 121.25 -71.455 ;
      RECT 121.15 -70.665 121.25 -70.13 ;
      RECT 121.15 -68.76 121.25 -68.225 ;
      RECT 121.15 -67.435 121.25 -66.9 ;
      RECT 121.15 -65.53 121.25 -64.995 ;
      RECT 121.15 -64.205 121.25 -63.67 ;
      RECT 121.15 -62.3 121.25 -61.765 ;
      RECT 121.15 -60.975 121.25 -60.44 ;
      RECT 121.15 -59.07 121.25 -58.535 ;
      RECT 121.15 -57.745 121.25 -57.21 ;
      RECT 121.15 -55.84 121.25 -55.305 ;
      RECT 121.15 -54.515 121.25 -53.98 ;
      RECT 121.15 -52.61 121.25 -52.075 ;
      RECT 121.15 -51.285 121.25 -50.75 ;
      RECT 121.15 -49.38 121.25 -48.845 ;
      RECT 121.15 -48.055 121.25 -47.52 ;
      RECT 121.15 -46.15 121.25 -45.615 ;
      RECT 121.15 -44.825 121.25 -44.29 ;
      RECT 121.15 -42.92 121.25 -42.385 ;
      RECT 121.15 -41.595 121.25 -41.06 ;
      RECT 121.15 -39.69 121.25 -39.155 ;
      RECT 121.15 -38.365 121.25 -37.83 ;
      RECT 121.15 -36.46 121.25 -35.925 ;
      RECT 121.15 -35.135 121.25 -34.6 ;
      RECT 121.15 -33.23 121.25 -32.695 ;
      RECT 121.15 -31.905 121.25 -31.37 ;
      RECT 121.15 -30 121.25 -29.465 ;
      RECT 121.15 -28.675 121.25 -28.14 ;
      RECT 121.15 -26.77 121.25 -26.235 ;
      RECT 121.15 -25.445 121.25 -24.91 ;
      RECT 121.15 -23.54 121.25 -23.005 ;
      RECT 121.15 -22.215 121.25 -21.68 ;
      RECT 121.15 -20.31 121.25 -19.775 ;
      RECT 121.15 -18.985 121.25 -18.45 ;
      RECT 121.15 -17.08 121.25 -16.545 ;
      RECT 121.15 -15.755 121.25 -15.22 ;
      RECT 121.15 -13.85 121.25 -13.315 ;
      RECT 121.15 -12.525 121.25 -11.99 ;
      RECT 121.15 -10.62 121.25 -10.085 ;
      RECT 121.15 -9.295 121.25 -8.76 ;
      RECT 121.15 -7.39 121.25 -6.855 ;
      RECT 121.15 -6.065 121.25 -5.53 ;
      RECT 121.15 -4.16 121.25 -3.625 ;
      RECT 121.15 -2.835 121.25 -2.3 ;
      RECT 121.15 -0.93 121.25 -0.395 ;
      RECT 121.15 0.395 121.25 0.93 ;
      RECT 121.025 -108.175 121.125 -107.215 ;
      RECT 120.65 -100.19 121 -100.07 ;
      RECT 120.65 -96.96 121 -96.84 ;
      RECT 120.65 -93.73 121 -93.61 ;
      RECT 120.65 -90.5 121 -90.38 ;
      RECT 120.65 -87.27 121 -87.15 ;
      RECT 120.65 -84.04 121 -83.92 ;
      RECT 120.65 -80.81 121 -80.69 ;
      RECT 120.65 -77.58 121 -77.46 ;
      RECT 120.65 -74.35 121 -74.23 ;
      RECT 120.65 -71.12 121 -71 ;
      RECT 120.65 -67.89 121 -67.77 ;
      RECT 120.65 -64.66 121 -64.54 ;
      RECT 120.65 -61.43 121 -61.31 ;
      RECT 120.65 -58.2 121 -58.08 ;
      RECT 120.65 -54.97 121 -54.85 ;
      RECT 120.65 -51.74 121 -51.62 ;
      RECT 120.65 -48.51 121 -48.39 ;
      RECT 120.65 -45.28 121 -45.16 ;
      RECT 120.65 -42.05 121 -41.93 ;
      RECT 120.65 -38.82 121 -38.7 ;
      RECT 120.65 -35.59 121 -35.47 ;
      RECT 120.65 -32.36 121 -32.24 ;
      RECT 120.65 -29.13 121 -29.01 ;
      RECT 120.65 -25.9 121 -25.78 ;
      RECT 120.65 -22.67 121 -22.55 ;
      RECT 120.65 -19.44 121 -19.32 ;
      RECT 120.65 -16.21 121 -16.09 ;
      RECT 120.65 -12.98 121 -12.86 ;
      RECT 120.65 -9.75 121 -9.63 ;
      RECT 120.65 -6.52 121 -6.4 ;
      RECT 120.65 -3.29 121 -3.17 ;
      RECT 120.65 -0.06 121 0.06 ;
      RECT 120.765 -108.175 120.865 -107.215 ;
      RECT 120.765 2.175 120.865 3.135 ;
      RECT 120.665 -113.555 120.765 -113.085 ;
      RECT 120.165 -100.19 120.515 -100.07 ;
      RECT 120.165 -96.96 120.515 -96.84 ;
      RECT 120.165 -93.73 120.515 -93.61 ;
      RECT 120.165 -90.5 120.515 -90.38 ;
      RECT 120.165 -87.27 120.515 -87.15 ;
      RECT 120.165 -84.04 120.515 -83.92 ;
      RECT 120.165 -80.81 120.515 -80.69 ;
      RECT 120.165 -77.58 120.515 -77.46 ;
      RECT 120.165 -74.35 120.515 -74.23 ;
      RECT 120.165 -71.12 120.515 -71 ;
      RECT 120.165 -67.89 120.515 -67.77 ;
      RECT 120.165 -64.66 120.515 -64.54 ;
      RECT 120.165 -61.43 120.515 -61.31 ;
      RECT 120.165 -58.2 120.515 -58.08 ;
      RECT 120.165 -54.97 120.515 -54.85 ;
      RECT 120.165 -51.74 120.515 -51.62 ;
      RECT 120.165 -48.51 120.515 -48.39 ;
      RECT 120.165 -45.28 120.515 -45.16 ;
      RECT 120.165 -42.05 120.515 -41.93 ;
      RECT 120.165 -38.82 120.515 -38.7 ;
      RECT 120.165 -35.59 120.515 -35.47 ;
      RECT 120.165 -32.36 120.515 -32.24 ;
      RECT 120.165 -29.13 120.515 -29.01 ;
      RECT 120.165 -25.9 120.515 -25.78 ;
      RECT 120.165 -22.67 120.515 -22.55 ;
      RECT 120.165 -19.44 120.515 -19.32 ;
      RECT 120.165 -16.21 120.515 -16.09 ;
      RECT 120.165 -12.98 120.515 -12.86 ;
      RECT 120.165 -9.75 120.515 -9.63 ;
      RECT 120.165 -6.52 120.515 -6.4 ;
      RECT 120.165 -3.29 120.515 -3.17 ;
      RECT 120.165 -0.06 120.515 0.06 ;
      RECT 120.3 -110.735 120.45 -110.445 ;
      RECT 120.335 -108.175 120.435 -107.215 ;
      RECT 120.335 2.175 120.435 3.135 ;
      RECT 120.315 -112.19 120.415 -111.65 ;
      RECT 120.075 -113.555 120.175 -113.085 ;
      RECT 120.075 -108.175 120.175 -107.215 ;
      RECT 119.95 -101.06 120.05 -100.525 ;
      RECT 119.95 -99.735 120.05 -99.2 ;
      RECT 119.95 -97.83 120.05 -97.295 ;
      RECT 119.95 -96.505 120.05 -95.97 ;
      RECT 119.95 -94.6 120.05 -94.065 ;
      RECT 119.95 -93.275 120.05 -92.74 ;
      RECT 119.95 -91.37 120.05 -90.835 ;
      RECT 119.95 -90.045 120.05 -89.51 ;
      RECT 119.95 -88.14 120.05 -87.605 ;
      RECT 119.95 -86.815 120.05 -86.28 ;
      RECT 119.95 -84.91 120.05 -84.375 ;
      RECT 119.95 -83.585 120.05 -83.05 ;
      RECT 119.95 -81.68 120.05 -81.145 ;
      RECT 119.95 -80.355 120.05 -79.82 ;
      RECT 119.95 -78.45 120.05 -77.915 ;
      RECT 119.95 -77.125 120.05 -76.59 ;
      RECT 119.95 -75.22 120.05 -74.685 ;
      RECT 119.95 -73.895 120.05 -73.36 ;
      RECT 119.95 -71.99 120.05 -71.455 ;
      RECT 119.95 -70.665 120.05 -70.13 ;
      RECT 119.95 -68.76 120.05 -68.225 ;
      RECT 119.95 -67.435 120.05 -66.9 ;
      RECT 119.95 -65.53 120.05 -64.995 ;
      RECT 119.95 -64.205 120.05 -63.67 ;
      RECT 119.95 -62.3 120.05 -61.765 ;
      RECT 119.95 -60.975 120.05 -60.44 ;
      RECT 119.95 -59.07 120.05 -58.535 ;
      RECT 119.95 -57.745 120.05 -57.21 ;
      RECT 119.95 -55.84 120.05 -55.305 ;
      RECT 119.95 -54.515 120.05 -53.98 ;
      RECT 119.95 -52.61 120.05 -52.075 ;
      RECT 119.95 -51.285 120.05 -50.75 ;
      RECT 119.95 -49.38 120.05 -48.845 ;
      RECT 119.95 -48.055 120.05 -47.52 ;
      RECT 119.95 -46.15 120.05 -45.615 ;
      RECT 119.95 -44.825 120.05 -44.29 ;
      RECT 119.95 -42.92 120.05 -42.385 ;
      RECT 119.95 -41.595 120.05 -41.06 ;
      RECT 119.95 -39.69 120.05 -39.155 ;
      RECT 119.95 -38.365 120.05 -37.83 ;
      RECT 119.95 -36.46 120.05 -35.925 ;
      RECT 119.95 -35.135 120.05 -34.6 ;
      RECT 119.95 -33.23 120.05 -32.695 ;
      RECT 119.95 -31.905 120.05 -31.37 ;
      RECT 119.95 -30 120.05 -29.465 ;
      RECT 119.95 -28.675 120.05 -28.14 ;
      RECT 119.95 -26.77 120.05 -26.235 ;
      RECT 119.95 -25.445 120.05 -24.91 ;
      RECT 119.95 -23.54 120.05 -23.005 ;
      RECT 119.95 -22.215 120.05 -21.68 ;
      RECT 119.95 -20.31 120.05 -19.775 ;
      RECT 119.95 -18.985 120.05 -18.45 ;
      RECT 119.95 -17.08 120.05 -16.545 ;
      RECT 119.95 -15.755 120.05 -15.22 ;
      RECT 119.95 -13.85 120.05 -13.315 ;
      RECT 119.95 -12.525 120.05 -11.99 ;
      RECT 119.95 -10.62 120.05 -10.085 ;
      RECT 119.95 -9.295 120.05 -8.76 ;
      RECT 119.95 -7.39 120.05 -6.855 ;
      RECT 119.95 -6.065 120.05 -5.53 ;
      RECT 119.95 -4.16 120.05 -3.625 ;
      RECT 119.95 -2.835 120.05 -2.3 ;
      RECT 119.95 -0.93 120.05 -0.395 ;
      RECT 119.95 0.395 120.05 0.93 ;
      RECT 119.825 -104.945 119.925 -103.985 ;
      RECT 119.45 -100.19 119.8 -100.07 ;
      RECT 119.45 -96.96 119.8 -96.84 ;
      RECT 119.45 -93.73 119.8 -93.61 ;
      RECT 119.45 -90.5 119.8 -90.38 ;
      RECT 119.45 -87.27 119.8 -87.15 ;
      RECT 119.45 -84.04 119.8 -83.92 ;
      RECT 119.45 -80.81 119.8 -80.69 ;
      RECT 119.45 -77.58 119.8 -77.46 ;
      RECT 119.45 -74.35 119.8 -74.23 ;
      RECT 119.45 -71.12 119.8 -71 ;
      RECT 119.45 -67.89 119.8 -67.77 ;
      RECT 119.45 -64.66 119.8 -64.54 ;
      RECT 119.45 -61.43 119.8 -61.31 ;
      RECT 119.45 -58.2 119.8 -58.08 ;
      RECT 119.45 -54.97 119.8 -54.85 ;
      RECT 119.45 -51.74 119.8 -51.62 ;
      RECT 119.45 -48.51 119.8 -48.39 ;
      RECT 119.45 -45.28 119.8 -45.16 ;
      RECT 119.45 -42.05 119.8 -41.93 ;
      RECT 119.45 -38.82 119.8 -38.7 ;
      RECT 119.45 -35.59 119.8 -35.47 ;
      RECT 119.45 -32.36 119.8 -32.24 ;
      RECT 119.45 -29.13 119.8 -29.01 ;
      RECT 119.45 -25.9 119.8 -25.78 ;
      RECT 119.45 -22.67 119.8 -22.55 ;
      RECT 119.45 -19.44 119.8 -19.32 ;
      RECT 119.45 -16.21 119.8 -16.09 ;
      RECT 119.45 -12.98 119.8 -12.86 ;
      RECT 119.45 -9.75 119.8 -9.63 ;
      RECT 119.45 -6.52 119.8 -6.4 ;
      RECT 119.45 -3.29 119.8 -3.17 ;
      RECT 119.45 -0.06 119.8 0.06 ;
      RECT 119.565 -104.945 119.665 -103.985 ;
      RECT 119.565 2.175 119.665 3.135 ;
      RECT 119.275 -112.255 119.375 -111.775 ;
      RECT 119.275 -110.765 119.375 -110.295 ;
      RECT 118.965 -100.19 119.315 -100.07 ;
      RECT 118.965 -96.96 119.315 -96.84 ;
      RECT 118.965 -93.73 119.315 -93.61 ;
      RECT 118.965 -90.5 119.315 -90.38 ;
      RECT 118.965 -87.27 119.315 -87.15 ;
      RECT 118.965 -84.04 119.315 -83.92 ;
      RECT 118.965 -80.81 119.315 -80.69 ;
      RECT 118.965 -77.58 119.315 -77.46 ;
      RECT 118.965 -74.35 119.315 -74.23 ;
      RECT 118.965 -71.12 119.315 -71 ;
      RECT 118.965 -67.89 119.315 -67.77 ;
      RECT 118.965 -64.66 119.315 -64.54 ;
      RECT 118.965 -61.43 119.315 -61.31 ;
      RECT 118.965 -58.2 119.315 -58.08 ;
      RECT 118.965 -54.97 119.315 -54.85 ;
      RECT 118.965 -51.74 119.315 -51.62 ;
      RECT 118.965 -48.51 119.315 -48.39 ;
      RECT 118.965 -45.28 119.315 -45.16 ;
      RECT 118.965 -42.05 119.315 -41.93 ;
      RECT 118.965 -38.82 119.315 -38.7 ;
      RECT 118.965 -35.59 119.315 -35.47 ;
      RECT 118.965 -32.36 119.315 -32.24 ;
      RECT 118.965 -29.13 119.315 -29.01 ;
      RECT 118.965 -25.9 119.315 -25.78 ;
      RECT 118.965 -22.67 119.315 -22.55 ;
      RECT 118.965 -19.44 119.315 -19.32 ;
      RECT 118.965 -16.21 119.315 -16.09 ;
      RECT 118.965 -12.98 119.315 -12.86 ;
      RECT 118.965 -9.75 119.315 -9.63 ;
      RECT 118.965 -6.52 119.315 -6.4 ;
      RECT 118.965 -3.29 119.315 -3.17 ;
      RECT 118.965 -0.06 119.315 0.06 ;
      RECT 119.135 -104.945 119.235 -103.985 ;
      RECT 119.135 2.175 119.235 3.135 ;
      RECT 115.235 -108.655 119.015 -108.535 ;
      RECT 118.875 -104.945 118.975 -103.985 ;
      RECT 118.75 -101.06 118.85 -100.525 ;
      RECT 118.75 -99.735 118.85 -99.2 ;
      RECT 118.75 -97.83 118.85 -97.295 ;
      RECT 118.75 -96.505 118.85 -95.97 ;
      RECT 118.75 -94.6 118.85 -94.065 ;
      RECT 118.75 -93.275 118.85 -92.74 ;
      RECT 118.75 -91.37 118.85 -90.835 ;
      RECT 118.75 -90.045 118.85 -89.51 ;
      RECT 118.75 -88.14 118.85 -87.605 ;
      RECT 118.75 -86.815 118.85 -86.28 ;
      RECT 118.75 -84.91 118.85 -84.375 ;
      RECT 118.75 -83.585 118.85 -83.05 ;
      RECT 118.75 -81.68 118.85 -81.145 ;
      RECT 118.75 -80.355 118.85 -79.82 ;
      RECT 118.75 -78.45 118.85 -77.915 ;
      RECT 118.75 -77.125 118.85 -76.59 ;
      RECT 118.75 -75.22 118.85 -74.685 ;
      RECT 118.75 -73.895 118.85 -73.36 ;
      RECT 118.75 -71.99 118.85 -71.455 ;
      RECT 118.75 -70.665 118.85 -70.13 ;
      RECT 118.75 -68.76 118.85 -68.225 ;
      RECT 118.75 -67.435 118.85 -66.9 ;
      RECT 118.75 -65.53 118.85 -64.995 ;
      RECT 118.75 -64.205 118.85 -63.67 ;
      RECT 118.75 -62.3 118.85 -61.765 ;
      RECT 118.75 -60.975 118.85 -60.44 ;
      RECT 118.75 -59.07 118.85 -58.535 ;
      RECT 118.75 -57.745 118.85 -57.21 ;
      RECT 118.75 -55.84 118.85 -55.305 ;
      RECT 118.75 -54.515 118.85 -53.98 ;
      RECT 118.75 -52.61 118.85 -52.075 ;
      RECT 118.75 -51.285 118.85 -50.75 ;
      RECT 118.75 -49.38 118.85 -48.845 ;
      RECT 118.75 -48.055 118.85 -47.52 ;
      RECT 118.75 -46.15 118.85 -45.615 ;
      RECT 118.75 -44.825 118.85 -44.29 ;
      RECT 118.75 -42.92 118.85 -42.385 ;
      RECT 118.75 -41.595 118.85 -41.06 ;
      RECT 118.75 -39.69 118.85 -39.155 ;
      RECT 118.75 -38.365 118.85 -37.83 ;
      RECT 118.75 -36.46 118.85 -35.925 ;
      RECT 118.75 -35.135 118.85 -34.6 ;
      RECT 118.75 -33.23 118.85 -32.695 ;
      RECT 118.75 -31.905 118.85 -31.37 ;
      RECT 118.75 -30 118.85 -29.465 ;
      RECT 118.75 -28.675 118.85 -28.14 ;
      RECT 118.75 -26.77 118.85 -26.235 ;
      RECT 118.75 -25.445 118.85 -24.91 ;
      RECT 118.75 -23.54 118.85 -23.005 ;
      RECT 118.75 -22.215 118.85 -21.68 ;
      RECT 118.75 -20.31 118.85 -19.775 ;
      RECT 118.75 -18.985 118.85 -18.45 ;
      RECT 118.75 -17.08 118.85 -16.545 ;
      RECT 118.75 -15.755 118.85 -15.22 ;
      RECT 118.75 -13.85 118.85 -13.315 ;
      RECT 118.75 -12.525 118.85 -11.99 ;
      RECT 118.75 -10.62 118.85 -10.085 ;
      RECT 118.75 -9.295 118.85 -8.76 ;
      RECT 118.75 -7.39 118.85 -6.855 ;
      RECT 118.75 -6.065 118.85 -5.53 ;
      RECT 118.75 -4.16 118.85 -3.625 ;
      RECT 118.75 -2.835 118.85 -2.3 ;
      RECT 118.75 -0.93 118.85 -0.395 ;
      RECT 118.75 0.395 118.85 0.93 ;
      RECT 118.685 -110.75 118.805 -110.37 ;
      RECT 118.685 -112.245 118.785 -111.775 ;
      RECT 118.625 -104.945 118.725 -103.985 ;
      RECT 118.25 -100.19 118.6 -100.07 ;
      RECT 118.25 -96.96 118.6 -96.84 ;
      RECT 118.25 -93.73 118.6 -93.61 ;
      RECT 118.25 -90.5 118.6 -90.38 ;
      RECT 118.25 -87.27 118.6 -87.15 ;
      RECT 118.25 -84.04 118.6 -83.92 ;
      RECT 118.25 -80.81 118.6 -80.69 ;
      RECT 118.25 -77.58 118.6 -77.46 ;
      RECT 118.25 -74.35 118.6 -74.23 ;
      RECT 118.25 -71.12 118.6 -71 ;
      RECT 118.25 -67.89 118.6 -67.77 ;
      RECT 118.25 -64.66 118.6 -64.54 ;
      RECT 118.25 -61.43 118.6 -61.31 ;
      RECT 118.25 -58.2 118.6 -58.08 ;
      RECT 118.25 -54.97 118.6 -54.85 ;
      RECT 118.25 -51.74 118.6 -51.62 ;
      RECT 118.25 -48.51 118.6 -48.39 ;
      RECT 118.25 -45.28 118.6 -45.16 ;
      RECT 118.25 -42.05 118.6 -41.93 ;
      RECT 118.25 -38.82 118.6 -38.7 ;
      RECT 118.25 -35.59 118.6 -35.47 ;
      RECT 118.25 -32.36 118.6 -32.24 ;
      RECT 118.25 -29.13 118.6 -29.01 ;
      RECT 118.25 -25.9 118.6 -25.78 ;
      RECT 118.25 -22.67 118.6 -22.55 ;
      RECT 118.25 -19.44 118.6 -19.32 ;
      RECT 118.25 -16.21 118.6 -16.09 ;
      RECT 118.25 -12.98 118.6 -12.86 ;
      RECT 118.25 -9.75 118.6 -9.63 ;
      RECT 118.25 -6.52 118.6 -6.4 ;
      RECT 118.25 -3.29 118.6 -3.17 ;
      RECT 118.25 -0.06 118.6 0.06 ;
      RECT 118.365 -104.945 118.465 -103.985 ;
      RECT 118.365 2.175 118.465 3.135 ;
      RECT 118.095 -109.595 118.23 -109.275 ;
      RECT 117.765 -100.19 118.115 -100.07 ;
      RECT 117.765 -96.96 118.115 -96.84 ;
      RECT 117.765 -93.73 118.115 -93.61 ;
      RECT 117.765 -90.5 118.115 -90.38 ;
      RECT 117.765 -87.27 118.115 -87.15 ;
      RECT 117.765 -84.04 118.115 -83.92 ;
      RECT 117.765 -80.81 118.115 -80.69 ;
      RECT 117.765 -77.58 118.115 -77.46 ;
      RECT 117.765 -74.35 118.115 -74.23 ;
      RECT 117.765 -71.12 118.115 -71 ;
      RECT 117.765 -67.89 118.115 -67.77 ;
      RECT 117.765 -64.66 118.115 -64.54 ;
      RECT 117.765 -61.43 118.115 -61.31 ;
      RECT 117.765 -58.2 118.115 -58.08 ;
      RECT 117.765 -54.97 118.115 -54.85 ;
      RECT 117.765 -51.74 118.115 -51.62 ;
      RECT 117.765 -48.51 118.115 -48.39 ;
      RECT 117.765 -45.28 118.115 -45.16 ;
      RECT 117.765 -42.05 118.115 -41.93 ;
      RECT 117.765 -38.82 118.115 -38.7 ;
      RECT 117.765 -35.59 118.115 -35.47 ;
      RECT 117.765 -32.36 118.115 -32.24 ;
      RECT 117.765 -29.13 118.115 -29.01 ;
      RECT 117.765 -25.9 118.115 -25.78 ;
      RECT 117.765 -22.67 118.115 -22.55 ;
      RECT 117.765 -19.44 118.115 -19.32 ;
      RECT 117.765 -16.21 118.115 -16.09 ;
      RECT 117.765 -12.98 118.115 -12.86 ;
      RECT 117.765 -9.75 118.115 -9.63 ;
      RECT 117.765 -6.52 118.115 -6.4 ;
      RECT 117.765 -3.29 118.115 -3.17 ;
      RECT 117.765 -0.06 118.115 0.06 ;
      RECT 117.935 -104.945 118.035 -103.985 ;
      RECT 117.935 2.175 118.035 3.135 ;
      RECT 117.76 -109.595 117.905 -109.275 ;
      RECT 117.675 -104.945 117.775 -103.985 ;
      RECT 117.55 -101.06 117.65 -100.525 ;
      RECT 117.55 -99.735 117.65 -99.2 ;
      RECT 117.55 -97.83 117.65 -97.295 ;
      RECT 117.55 -96.505 117.65 -95.97 ;
      RECT 117.55 -94.6 117.65 -94.065 ;
      RECT 117.55 -93.275 117.65 -92.74 ;
      RECT 117.55 -91.37 117.65 -90.835 ;
      RECT 117.55 -90.045 117.65 -89.51 ;
      RECT 117.55 -88.14 117.65 -87.605 ;
      RECT 117.55 -86.815 117.65 -86.28 ;
      RECT 117.55 -84.91 117.65 -84.375 ;
      RECT 117.55 -83.585 117.65 -83.05 ;
      RECT 117.55 -81.68 117.65 -81.145 ;
      RECT 117.55 -80.355 117.65 -79.82 ;
      RECT 117.55 -78.45 117.65 -77.915 ;
      RECT 117.55 -77.125 117.65 -76.59 ;
      RECT 117.55 -75.22 117.65 -74.685 ;
      RECT 117.55 -73.895 117.65 -73.36 ;
      RECT 117.55 -71.99 117.65 -71.455 ;
      RECT 117.55 -70.665 117.65 -70.13 ;
      RECT 117.55 -68.76 117.65 -68.225 ;
      RECT 117.55 -67.435 117.65 -66.9 ;
      RECT 117.55 -65.53 117.65 -64.995 ;
      RECT 117.55 -64.205 117.65 -63.67 ;
      RECT 117.55 -62.3 117.65 -61.765 ;
      RECT 117.55 -60.975 117.65 -60.44 ;
      RECT 117.55 -59.07 117.65 -58.535 ;
      RECT 117.55 -57.745 117.65 -57.21 ;
      RECT 117.55 -55.84 117.65 -55.305 ;
      RECT 117.55 -54.515 117.65 -53.98 ;
      RECT 117.55 -52.61 117.65 -52.075 ;
      RECT 117.55 -51.285 117.65 -50.75 ;
      RECT 117.55 -49.38 117.65 -48.845 ;
      RECT 117.55 -48.055 117.65 -47.52 ;
      RECT 117.55 -46.15 117.65 -45.615 ;
      RECT 117.55 -44.825 117.65 -44.29 ;
      RECT 117.55 -42.92 117.65 -42.385 ;
      RECT 117.55 -41.595 117.65 -41.06 ;
      RECT 117.55 -39.69 117.65 -39.155 ;
      RECT 117.55 -38.365 117.65 -37.83 ;
      RECT 117.55 -36.46 117.65 -35.925 ;
      RECT 117.55 -35.135 117.65 -34.6 ;
      RECT 117.55 -33.23 117.65 -32.695 ;
      RECT 117.55 -31.905 117.65 -31.37 ;
      RECT 117.55 -30 117.65 -29.465 ;
      RECT 117.55 -28.675 117.65 -28.14 ;
      RECT 117.55 -26.77 117.65 -26.235 ;
      RECT 117.55 -25.445 117.65 -24.91 ;
      RECT 117.55 -23.54 117.65 -23.005 ;
      RECT 117.55 -22.215 117.65 -21.68 ;
      RECT 117.55 -20.31 117.65 -19.775 ;
      RECT 117.55 -18.985 117.65 -18.45 ;
      RECT 117.55 -17.08 117.65 -16.545 ;
      RECT 117.55 -15.755 117.65 -15.22 ;
      RECT 117.55 -13.85 117.65 -13.315 ;
      RECT 117.55 -12.525 117.65 -11.99 ;
      RECT 117.55 -10.62 117.65 -10.085 ;
      RECT 117.55 -9.295 117.65 -8.76 ;
      RECT 117.55 -7.39 117.65 -6.855 ;
      RECT 117.55 -6.065 117.65 -5.53 ;
      RECT 117.55 -4.16 117.65 -3.625 ;
      RECT 117.55 -2.835 117.65 -2.3 ;
      RECT 117.55 -0.93 117.65 -0.395 ;
      RECT 117.55 0.395 117.65 0.93 ;
      RECT 117.425 -108.175 117.525 -107.215 ;
      RECT 117.05 -100.19 117.4 -100.07 ;
      RECT 117.05 -96.96 117.4 -96.84 ;
      RECT 117.05 -93.73 117.4 -93.61 ;
      RECT 117.05 -90.5 117.4 -90.38 ;
      RECT 117.05 -87.27 117.4 -87.15 ;
      RECT 117.05 -84.04 117.4 -83.92 ;
      RECT 117.05 -80.81 117.4 -80.69 ;
      RECT 117.05 -77.58 117.4 -77.46 ;
      RECT 117.05 -74.35 117.4 -74.23 ;
      RECT 117.05 -71.12 117.4 -71 ;
      RECT 117.05 -67.89 117.4 -67.77 ;
      RECT 117.05 -64.66 117.4 -64.54 ;
      RECT 117.05 -61.43 117.4 -61.31 ;
      RECT 117.05 -58.2 117.4 -58.08 ;
      RECT 117.05 -54.97 117.4 -54.85 ;
      RECT 117.05 -51.74 117.4 -51.62 ;
      RECT 117.05 -48.51 117.4 -48.39 ;
      RECT 117.05 -45.28 117.4 -45.16 ;
      RECT 117.05 -42.05 117.4 -41.93 ;
      RECT 117.05 -38.82 117.4 -38.7 ;
      RECT 117.05 -35.59 117.4 -35.47 ;
      RECT 117.05 -32.36 117.4 -32.24 ;
      RECT 117.05 -29.13 117.4 -29.01 ;
      RECT 117.05 -25.9 117.4 -25.78 ;
      RECT 117.05 -22.67 117.4 -22.55 ;
      RECT 117.05 -19.44 117.4 -19.32 ;
      RECT 117.05 -16.21 117.4 -16.09 ;
      RECT 117.05 -12.98 117.4 -12.86 ;
      RECT 117.05 -9.75 117.4 -9.63 ;
      RECT 117.05 -6.52 117.4 -6.4 ;
      RECT 117.05 -3.29 117.4 -3.17 ;
      RECT 117.05 -0.06 117.4 0.06 ;
      RECT 117.255 -112.255 117.355 -111.775 ;
      RECT 117.255 -110.765 117.355 -110.295 ;
      RECT 117.165 -108.175 117.265 -107.215 ;
      RECT 117.165 2.175 117.265 3.135 ;
      RECT 116.565 -100.19 116.915 -100.07 ;
      RECT 116.565 -96.96 116.915 -96.84 ;
      RECT 116.565 -93.73 116.915 -93.61 ;
      RECT 116.565 -90.5 116.915 -90.38 ;
      RECT 116.565 -87.27 116.915 -87.15 ;
      RECT 116.565 -84.04 116.915 -83.92 ;
      RECT 116.565 -80.81 116.915 -80.69 ;
      RECT 116.565 -77.58 116.915 -77.46 ;
      RECT 116.565 -74.35 116.915 -74.23 ;
      RECT 116.565 -71.12 116.915 -71 ;
      RECT 116.565 -67.89 116.915 -67.77 ;
      RECT 116.565 -64.66 116.915 -64.54 ;
      RECT 116.565 -61.43 116.915 -61.31 ;
      RECT 116.565 -58.2 116.915 -58.08 ;
      RECT 116.565 -54.97 116.915 -54.85 ;
      RECT 116.565 -51.74 116.915 -51.62 ;
      RECT 116.565 -48.51 116.915 -48.39 ;
      RECT 116.565 -45.28 116.915 -45.16 ;
      RECT 116.565 -42.05 116.915 -41.93 ;
      RECT 116.565 -38.82 116.915 -38.7 ;
      RECT 116.565 -35.59 116.915 -35.47 ;
      RECT 116.565 -32.36 116.915 -32.24 ;
      RECT 116.565 -29.13 116.915 -29.01 ;
      RECT 116.565 -25.9 116.915 -25.78 ;
      RECT 116.565 -22.67 116.915 -22.55 ;
      RECT 116.565 -19.44 116.915 -19.32 ;
      RECT 116.565 -16.21 116.915 -16.09 ;
      RECT 116.565 -12.98 116.915 -12.86 ;
      RECT 116.565 -9.75 116.915 -9.63 ;
      RECT 116.565 -6.52 116.915 -6.4 ;
      RECT 116.565 -3.29 116.915 -3.17 ;
      RECT 116.565 -0.06 116.915 0.06 ;
      RECT 116.735 -108.175 116.835 -107.215 ;
      RECT 116.735 2.175 116.835 3.135 ;
      RECT 116.63 -110.765 116.8 -110.385 ;
      RECT 116.665 -112.245 116.765 -111.775 ;
      RECT 116.475 -108.175 116.575 -107.215 ;
      RECT 116.35 -101.06 116.45 -100.525 ;
      RECT 116.35 -99.735 116.45 -99.2 ;
      RECT 116.35 -97.83 116.45 -97.295 ;
      RECT 116.35 -96.505 116.45 -95.97 ;
      RECT 116.35 -94.6 116.45 -94.065 ;
      RECT 116.35 -93.275 116.45 -92.74 ;
      RECT 116.35 -91.37 116.45 -90.835 ;
      RECT 116.35 -90.045 116.45 -89.51 ;
      RECT 116.35 -88.14 116.45 -87.605 ;
      RECT 116.35 -86.815 116.45 -86.28 ;
      RECT 116.35 -84.91 116.45 -84.375 ;
      RECT 116.35 -83.585 116.45 -83.05 ;
      RECT 116.35 -81.68 116.45 -81.145 ;
      RECT 116.35 -80.355 116.45 -79.82 ;
      RECT 116.35 -78.45 116.45 -77.915 ;
      RECT 116.35 -77.125 116.45 -76.59 ;
      RECT 116.35 -75.22 116.45 -74.685 ;
      RECT 116.35 -73.895 116.45 -73.36 ;
      RECT 116.35 -71.99 116.45 -71.455 ;
      RECT 116.35 -70.665 116.45 -70.13 ;
      RECT 116.35 -68.76 116.45 -68.225 ;
      RECT 116.35 -67.435 116.45 -66.9 ;
      RECT 116.35 -65.53 116.45 -64.995 ;
      RECT 116.35 -64.205 116.45 -63.67 ;
      RECT 116.35 -62.3 116.45 -61.765 ;
      RECT 116.35 -60.975 116.45 -60.44 ;
      RECT 116.35 -59.07 116.45 -58.535 ;
      RECT 116.35 -57.745 116.45 -57.21 ;
      RECT 116.35 -55.84 116.45 -55.305 ;
      RECT 116.35 -54.515 116.45 -53.98 ;
      RECT 116.35 -52.61 116.45 -52.075 ;
      RECT 116.35 -51.285 116.45 -50.75 ;
      RECT 116.35 -49.38 116.45 -48.845 ;
      RECT 116.35 -48.055 116.45 -47.52 ;
      RECT 116.35 -46.15 116.45 -45.615 ;
      RECT 116.35 -44.825 116.45 -44.29 ;
      RECT 116.35 -42.92 116.45 -42.385 ;
      RECT 116.35 -41.595 116.45 -41.06 ;
      RECT 116.35 -39.69 116.45 -39.155 ;
      RECT 116.35 -38.365 116.45 -37.83 ;
      RECT 116.35 -36.46 116.45 -35.925 ;
      RECT 116.35 -35.135 116.45 -34.6 ;
      RECT 116.35 -33.23 116.45 -32.695 ;
      RECT 116.35 -31.905 116.45 -31.37 ;
      RECT 116.35 -30 116.45 -29.465 ;
      RECT 116.35 -28.675 116.45 -28.14 ;
      RECT 116.35 -26.77 116.45 -26.235 ;
      RECT 116.35 -25.445 116.45 -24.91 ;
      RECT 116.35 -23.54 116.45 -23.005 ;
      RECT 116.35 -22.215 116.45 -21.68 ;
      RECT 116.35 -20.31 116.45 -19.775 ;
      RECT 116.35 -18.985 116.45 -18.45 ;
      RECT 116.35 -17.08 116.45 -16.545 ;
      RECT 116.35 -15.755 116.45 -15.22 ;
      RECT 116.35 -13.85 116.45 -13.315 ;
      RECT 116.35 -12.525 116.45 -11.99 ;
      RECT 116.35 -10.62 116.45 -10.085 ;
      RECT 116.35 -9.295 116.45 -8.76 ;
      RECT 116.35 -7.39 116.45 -6.855 ;
      RECT 116.35 -6.065 116.45 -5.53 ;
      RECT 116.35 -4.16 116.45 -3.625 ;
      RECT 116.35 -2.835 116.45 -2.3 ;
      RECT 116.35 -0.93 116.45 -0.395 ;
      RECT 116.35 0.395 116.45 0.93 ;
      RECT 116.225 -108.175 116.325 -107.215 ;
      RECT 115.85 -100.19 116.2 -100.07 ;
      RECT 115.85 -96.96 116.2 -96.84 ;
      RECT 115.85 -93.73 116.2 -93.61 ;
      RECT 115.85 -90.5 116.2 -90.38 ;
      RECT 115.85 -87.27 116.2 -87.15 ;
      RECT 115.85 -84.04 116.2 -83.92 ;
      RECT 115.85 -80.81 116.2 -80.69 ;
      RECT 115.85 -77.58 116.2 -77.46 ;
      RECT 115.85 -74.35 116.2 -74.23 ;
      RECT 115.85 -71.12 116.2 -71 ;
      RECT 115.85 -67.89 116.2 -67.77 ;
      RECT 115.85 -64.66 116.2 -64.54 ;
      RECT 115.85 -61.43 116.2 -61.31 ;
      RECT 115.85 -58.2 116.2 -58.08 ;
      RECT 115.85 -54.97 116.2 -54.85 ;
      RECT 115.85 -51.74 116.2 -51.62 ;
      RECT 115.85 -48.51 116.2 -48.39 ;
      RECT 115.85 -45.28 116.2 -45.16 ;
      RECT 115.85 -42.05 116.2 -41.93 ;
      RECT 115.85 -38.82 116.2 -38.7 ;
      RECT 115.85 -35.59 116.2 -35.47 ;
      RECT 115.85 -32.36 116.2 -32.24 ;
      RECT 115.85 -29.13 116.2 -29.01 ;
      RECT 115.85 -25.9 116.2 -25.78 ;
      RECT 115.85 -22.67 116.2 -22.55 ;
      RECT 115.85 -19.44 116.2 -19.32 ;
      RECT 115.85 -16.21 116.2 -16.09 ;
      RECT 115.85 -12.98 116.2 -12.86 ;
      RECT 115.85 -9.75 116.2 -9.63 ;
      RECT 115.85 -6.52 116.2 -6.4 ;
      RECT 115.85 -3.29 116.2 -3.17 ;
      RECT 115.85 -0.06 116.2 0.06 ;
      RECT 115.965 -108.175 116.065 -107.215 ;
      RECT 115.965 2.175 116.065 3.135 ;
      RECT 115.865 -113.555 115.965 -113.085 ;
      RECT 115.365 -100.19 115.715 -100.07 ;
      RECT 115.365 -96.96 115.715 -96.84 ;
      RECT 115.365 -93.73 115.715 -93.61 ;
      RECT 115.365 -90.5 115.715 -90.38 ;
      RECT 115.365 -87.27 115.715 -87.15 ;
      RECT 115.365 -84.04 115.715 -83.92 ;
      RECT 115.365 -80.81 115.715 -80.69 ;
      RECT 115.365 -77.58 115.715 -77.46 ;
      RECT 115.365 -74.35 115.715 -74.23 ;
      RECT 115.365 -71.12 115.715 -71 ;
      RECT 115.365 -67.89 115.715 -67.77 ;
      RECT 115.365 -64.66 115.715 -64.54 ;
      RECT 115.365 -61.43 115.715 -61.31 ;
      RECT 115.365 -58.2 115.715 -58.08 ;
      RECT 115.365 -54.97 115.715 -54.85 ;
      RECT 115.365 -51.74 115.715 -51.62 ;
      RECT 115.365 -48.51 115.715 -48.39 ;
      RECT 115.365 -45.28 115.715 -45.16 ;
      RECT 115.365 -42.05 115.715 -41.93 ;
      RECT 115.365 -38.82 115.715 -38.7 ;
      RECT 115.365 -35.59 115.715 -35.47 ;
      RECT 115.365 -32.36 115.715 -32.24 ;
      RECT 115.365 -29.13 115.715 -29.01 ;
      RECT 115.365 -25.9 115.715 -25.78 ;
      RECT 115.365 -22.67 115.715 -22.55 ;
      RECT 115.365 -19.44 115.715 -19.32 ;
      RECT 115.365 -16.21 115.715 -16.09 ;
      RECT 115.365 -12.98 115.715 -12.86 ;
      RECT 115.365 -9.75 115.715 -9.63 ;
      RECT 115.365 -6.52 115.715 -6.4 ;
      RECT 115.365 -3.29 115.715 -3.17 ;
      RECT 115.365 -0.06 115.715 0.06 ;
      RECT 115.5 -110.735 115.65 -110.445 ;
      RECT 115.535 -108.175 115.635 -107.215 ;
      RECT 115.535 2.175 115.635 3.135 ;
      RECT 115.515 -112.19 115.615 -111.65 ;
      RECT 115.275 -113.555 115.375 -113.085 ;
      RECT 115.275 -108.175 115.375 -107.215 ;
      RECT 115.15 -101.06 115.25 -100.525 ;
      RECT 115.15 -99.735 115.25 -99.2 ;
      RECT 115.15 -97.83 115.25 -97.295 ;
      RECT 115.15 -96.505 115.25 -95.97 ;
      RECT 115.15 -94.6 115.25 -94.065 ;
      RECT 115.15 -93.275 115.25 -92.74 ;
      RECT 115.15 -91.37 115.25 -90.835 ;
      RECT 115.15 -90.045 115.25 -89.51 ;
      RECT 115.15 -88.14 115.25 -87.605 ;
      RECT 115.15 -86.815 115.25 -86.28 ;
      RECT 115.15 -84.91 115.25 -84.375 ;
      RECT 115.15 -83.585 115.25 -83.05 ;
      RECT 115.15 -81.68 115.25 -81.145 ;
      RECT 115.15 -80.355 115.25 -79.82 ;
      RECT 115.15 -78.45 115.25 -77.915 ;
      RECT 115.15 -77.125 115.25 -76.59 ;
      RECT 115.15 -75.22 115.25 -74.685 ;
      RECT 115.15 -73.895 115.25 -73.36 ;
      RECT 115.15 -71.99 115.25 -71.455 ;
      RECT 115.15 -70.665 115.25 -70.13 ;
      RECT 115.15 -68.76 115.25 -68.225 ;
      RECT 115.15 -67.435 115.25 -66.9 ;
      RECT 115.15 -65.53 115.25 -64.995 ;
      RECT 115.15 -64.205 115.25 -63.67 ;
      RECT 115.15 -62.3 115.25 -61.765 ;
      RECT 115.15 -60.975 115.25 -60.44 ;
      RECT 115.15 -59.07 115.25 -58.535 ;
      RECT 115.15 -57.745 115.25 -57.21 ;
      RECT 115.15 -55.84 115.25 -55.305 ;
      RECT 115.15 -54.515 115.25 -53.98 ;
      RECT 115.15 -52.61 115.25 -52.075 ;
      RECT 115.15 -51.285 115.25 -50.75 ;
      RECT 115.15 -49.38 115.25 -48.845 ;
      RECT 115.15 -48.055 115.25 -47.52 ;
      RECT 115.15 -46.15 115.25 -45.615 ;
      RECT 115.15 -44.825 115.25 -44.29 ;
      RECT 115.15 -42.92 115.25 -42.385 ;
      RECT 115.15 -41.595 115.25 -41.06 ;
      RECT 115.15 -39.69 115.25 -39.155 ;
      RECT 115.15 -38.365 115.25 -37.83 ;
      RECT 115.15 -36.46 115.25 -35.925 ;
      RECT 115.15 -35.135 115.25 -34.6 ;
      RECT 115.15 -33.23 115.25 -32.695 ;
      RECT 115.15 -31.905 115.25 -31.37 ;
      RECT 115.15 -30 115.25 -29.465 ;
      RECT 115.15 -28.675 115.25 -28.14 ;
      RECT 115.15 -26.77 115.25 -26.235 ;
      RECT 115.15 -25.445 115.25 -24.91 ;
      RECT 115.15 -23.54 115.25 -23.005 ;
      RECT 115.15 -22.215 115.25 -21.68 ;
      RECT 115.15 -20.31 115.25 -19.775 ;
      RECT 115.15 -18.985 115.25 -18.45 ;
      RECT 115.15 -17.08 115.25 -16.545 ;
      RECT 115.15 -15.755 115.25 -15.22 ;
      RECT 115.15 -13.85 115.25 -13.315 ;
      RECT 115.15 -12.525 115.25 -11.99 ;
      RECT 115.15 -10.62 115.25 -10.085 ;
      RECT 115.15 -9.295 115.25 -8.76 ;
      RECT 115.15 -7.39 115.25 -6.855 ;
      RECT 115.15 -6.065 115.25 -5.53 ;
      RECT 115.15 -4.16 115.25 -3.625 ;
      RECT 115.15 -2.835 115.25 -2.3 ;
      RECT 115.15 -0.93 115.25 -0.395 ;
      RECT 115.15 0.395 115.25 0.93 ;
      RECT 115.025 -104.945 115.125 -103.985 ;
      RECT 114.65 -100.19 115 -100.07 ;
      RECT 114.65 -96.96 115 -96.84 ;
      RECT 114.65 -93.73 115 -93.61 ;
      RECT 114.65 -90.5 115 -90.38 ;
      RECT 114.65 -87.27 115 -87.15 ;
      RECT 114.65 -84.04 115 -83.92 ;
      RECT 114.65 -80.81 115 -80.69 ;
      RECT 114.65 -77.58 115 -77.46 ;
      RECT 114.65 -74.35 115 -74.23 ;
      RECT 114.65 -71.12 115 -71 ;
      RECT 114.65 -67.89 115 -67.77 ;
      RECT 114.65 -64.66 115 -64.54 ;
      RECT 114.65 -61.43 115 -61.31 ;
      RECT 114.65 -58.2 115 -58.08 ;
      RECT 114.65 -54.97 115 -54.85 ;
      RECT 114.65 -51.74 115 -51.62 ;
      RECT 114.65 -48.51 115 -48.39 ;
      RECT 114.65 -45.28 115 -45.16 ;
      RECT 114.65 -42.05 115 -41.93 ;
      RECT 114.65 -38.82 115 -38.7 ;
      RECT 114.65 -35.59 115 -35.47 ;
      RECT 114.65 -32.36 115 -32.24 ;
      RECT 114.65 -29.13 115 -29.01 ;
      RECT 114.65 -25.9 115 -25.78 ;
      RECT 114.65 -22.67 115 -22.55 ;
      RECT 114.65 -19.44 115 -19.32 ;
      RECT 114.65 -16.21 115 -16.09 ;
      RECT 114.65 -12.98 115 -12.86 ;
      RECT 114.65 -9.75 115 -9.63 ;
      RECT 114.65 -6.52 115 -6.4 ;
      RECT 114.65 -3.29 115 -3.17 ;
      RECT 114.65 -0.06 115 0.06 ;
      RECT 114.765 -104.945 114.865 -103.985 ;
      RECT 114.765 2.175 114.865 3.135 ;
      RECT 114.475 -112.255 114.575 -111.775 ;
      RECT 114.475 -110.765 114.575 -110.295 ;
      RECT 114.165 -100.19 114.515 -100.07 ;
      RECT 114.165 -96.96 114.515 -96.84 ;
      RECT 114.165 -93.73 114.515 -93.61 ;
      RECT 114.165 -90.5 114.515 -90.38 ;
      RECT 114.165 -87.27 114.515 -87.15 ;
      RECT 114.165 -84.04 114.515 -83.92 ;
      RECT 114.165 -80.81 114.515 -80.69 ;
      RECT 114.165 -77.58 114.515 -77.46 ;
      RECT 114.165 -74.35 114.515 -74.23 ;
      RECT 114.165 -71.12 114.515 -71 ;
      RECT 114.165 -67.89 114.515 -67.77 ;
      RECT 114.165 -64.66 114.515 -64.54 ;
      RECT 114.165 -61.43 114.515 -61.31 ;
      RECT 114.165 -58.2 114.515 -58.08 ;
      RECT 114.165 -54.97 114.515 -54.85 ;
      RECT 114.165 -51.74 114.515 -51.62 ;
      RECT 114.165 -48.51 114.515 -48.39 ;
      RECT 114.165 -45.28 114.515 -45.16 ;
      RECT 114.165 -42.05 114.515 -41.93 ;
      RECT 114.165 -38.82 114.515 -38.7 ;
      RECT 114.165 -35.59 114.515 -35.47 ;
      RECT 114.165 -32.36 114.515 -32.24 ;
      RECT 114.165 -29.13 114.515 -29.01 ;
      RECT 114.165 -25.9 114.515 -25.78 ;
      RECT 114.165 -22.67 114.515 -22.55 ;
      RECT 114.165 -19.44 114.515 -19.32 ;
      RECT 114.165 -16.21 114.515 -16.09 ;
      RECT 114.165 -12.98 114.515 -12.86 ;
      RECT 114.165 -9.75 114.515 -9.63 ;
      RECT 114.165 -6.52 114.515 -6.4 ;
      RECT 114.165 -3.29 114.515 -3.17 ;
      RECT 114.165 -0.06 114.515 0.06 ;
      RECT 114.335 -104.945 114.435 -103.985 ;
      RECT 114.335 2.175 114.435 3.135 ;
      RECT 110.435 -108.655 114.215 -108.535 ;
      RECT 114.075 -104.945 114.175 -103.985 ;
      RECT 113.95 -101.06 114.05 -100.525 ;
      RECT 113.95 -99.735 114.05 -99.2 ;
      RECT 113.95 -97.83 114.05 -97.295 ;
      RECT 113.95 -96.505 114.05 -95.97 ;
      RECT 113.95 -94.6 114.05 -94.065 ;
      RECT 113.95 -93.275 114.05 -92.74 ;
      RECT 113.95 -91.37 114.05 -90.835 ;
      RECT 113.95 -90.045 114.05 -89.51 ;
      RECT 113.95 -88.14 114.05 -87.605 ;
      RECT 113.95 -86.815 114.05 -86.28 ;
      RECT 113.95 -84.91 114.05 -84.375 ;
      RECT 113.95 -83.585 114.05 -83.05 ;
      RECT 113.95 -81.68 114.05 -81.145 ;
      RECT 113.95 -80.355 114.05 -79.82 ;
      RECT 113.95 -78.45 114.05 -77.915 ;
      RECT 113.95 -77.125 114.05 -76.59 ;
      RECT 113.95 -75.22 114.05 -74.685 ;
      RECT 113.95 -73.895 114.05 -73.36 ;
      RECT 113.95 -71.99 114.05 -71.455 ;
      RECT 113.95 -70.665 114.05 -70.13 ;
      RECT 113.95 -68.76 114.05 -68.225 ;
      RECT 113.95 -67.435 114.05 -66.9 ;
      RECT 113.95 -65.53 114.05 -64.995 ;
      RECT 113.95 -64.205 114.05 -63.67 ;
      RECT 113.95 -62.3 114.05 -61.765 ;
      RECT 113.95 -60.975 114.05 -60.44 ;
      RECT 113.95 -59.07 114.05 -58.535 ;
      RECT 113.95 -57.745 114.05 -57.21 ;
      RECT 113.95 -55.84 114.05 -55.305 ;
      RECT 113.95 -54.515 114.05 -53.98 ;
      RECT 113.95 -52.61 114.05 -52.075 ;
      RECT 113.95 -51.285 114.05 -50.75 ;
      RECT 113.95 -49.38 114.05 -48.845 ;
      RECT 113.95 -48.055 114.05 -47.52 ;
      RECT 113.95 -46.15 114.05 -45.615 ;
      RECT 113.95 -44.825 114.05 -44.29 ;
      RECT 113.95 -42.92 114.05 -42.385 ;
      RECT 113.95 -41.595 114.05 -41.06 ;
      RECT 113.95 -39.69 114.05 -39.155 ;
      RECT 113.95 -38.365 114.05 -37.83 ;
      RECT 113.95 -36.46 114.05 -35.925 ;
      RECT 113.95 -35.135 114.05 -34.6 ;
      RECT 113.95 -33.23 114.05 -32.695 ;
      RECT 113.95 -31.905 114.05 -31.37 ;
      RECT 113.95 -30 114.05 -29.465 ;
      RECT 113.95 -28.675 114.05 -28.14 ;
      RECT 113.95 -26.77 114.05 -26.235 ;
      RECT 113.95 -25.445 114.05 -24.91 ;
      RECT 113.95 -23.54 114.05 -23.005 ;
      RECT 113.95 -22.215 114.05 -21.68 ;
      RECT 113.95 -20.31 114.05 -19.775 ;
      RECT 113.95 -18.985 114.05 -18.45 ;
      RECT 113.95 -17.08 114.05 -16.545 ;
      RECT 113.95 -15.755 114.05 -15.22 ;
      RECT 113.95 -13.85 114.05 -13.315 ;
      RECT 113.95 -12.525 114.05 -11.99 ;
      RECT 113.95 -10.62 114.05 -10.085 ;
      RECT 113.95 -9.295 114.05 -8.76 ;
      RECT 113.95 -7.39 114.05 -6.855 ;
      RECT 113.95 -6.065 114.05 -5.53 ;
      RECT 113.95 -4.16 114.05 -3.625 ;
      RECT 113.95 -2.835 114.05 -2.3 ;
      RECT 113.95 -0.93 114.05 -0.395 ;
      RECT 113.95 0.395 114.05 0.93 ;
      RECT 113.885 -110.75 114.005 -110.37 ;
      RECT 113.885 -112.245 113.985 -111.775 ;
      RECT 113.825 -104.945 113.925 -103.985 ;
      RECT 113.45 -100.19 113.8 -100.07 ;
      RECT 113.45 -96.96 113.8 -96.84 ;
      RECT 113.45 -93.73 113.8 -93.61 ;
      RECT 113.45 -90.5 113.8 -90.38 ;
      RECT 113.45 -87.27 113.8 -87.15 ;
      RECT 113.45 -84.04 113.8 -83.92 ;
      RECT 113.45 -80.81 113.8 -80.69 ;
      RECT 113.45 -77.58 113.8 -77.46 ;
      RECT 113.45 -74.35 113.8 -74.23 ;
      RECT 113.45 -71.12 113.8 -71 ;
      RECT 113.45 -67.89 113.8 -67.77 ;
      RECT 113.45 -64.66 113.8 -64.54 ;
      RECT 113.45 -61.43 113.8 -61.31 ;
      RECT 113.45 -58.2 113.8 -58.08 ;
      RECT 113.45 -54.97 113.8 -54.85 ;
      RECT 113.45 -51.74 113.8 -51.62 ;
      RECT 113.45 -48.51 113.8 -48.39 ;
      RECT 113.45 -45.28 113.8 -45.16 ;
      RECT 113.45 -42.05 113.8 -41.93 ;
      RECT 113.45 -38.82 113.8 -38.7 ;
      RECT 113.45 -35.59 113.8 -35.47 ;
      RECT 113.45 -32.36 113.8 -32.24 ;
      RECT 113.45 -29.13 113.8 -29.01 ;
      RECT 113.45 -25.9 113.8 -25.78 ;
      RECT 113.45 -22.67 113.8 -22.55 ;
      RECT 113.45 -19.44 113.8 -19.32 ;
      RECT 113.45 -16.21 113.8 -16.09 ;
      RECT 113.45 -12.98 113.8 -12.86 ;
      RECT 113.45 -9.75 113.8 -9.63 ;
      RECT 113.45 -6.52 113.8 -6.4 ;
      RECT 113.45 -3.29 113.8 -3.17 ;
      RECT 113.45 -0.06 113.8 0.06 ;
      RECT 113.565 -104.945 113.665 -103.985 ;
      RECT 113.565 2.175 113.665 3.135 ;
      RECT 113.295 -109.595 113.43 -109.275 ;
      RECT 112.965 -100.19 113.315 -100.07 ;
      RECT 112.965 -96.96 113.315 -96.84 ;
      RECT 112.965 -93.73 113.315 -93.61 ;
      RECT 112.965 -90.5 113.315 -90.38 ;
      RECT 112.965 -87.27 113.315 -87.15 ;
      RECT 112.965 -84.04 113.315 -83.92 ;
      RECT 112.965 -80.81 113.315 -80.69 ;
      RECT 112.965 -77.58 113.315 -77.46 ;
      RECT 112.965 -74.35 113.315 -74.23 ;
      RECT 112.965 -71.12 113.315 -71 ;
      RECT 112.965 -67.89 113.315 -67.77 ;
      RECT 112.965 -64.66 113.315 -64.54 ;
      RECT 112.965 -61.43 113.315 -61.31 ;
      RECT 112.965 -58.2 113.315 -58.08 ;
      RECT 112.965 -54.97 113.315 -54.85 ;
      RECT 112.965 -51.74 113.315 -51.62 ;
      RECT 112.965 -48.51 113.315 -48.39 ;
      RECT 112.965 -45.28 113.315 -45.16 ;
      RECT 112.965 -42.05 113.315 -41.93 ;
      RECT 112.965 -38.82 113.315 -38.7 ;
      RECT 112.965 -35.59 113.315 -35.47 ;
      RECT 112.965 -32.36 113.315 -32.24 ;
      RECT 112.965 -29.13 113.315 -29.01 ;
      RECT 112.965 -25.9 113.315 -25.78 ;
      RECT 112.965 -22.67 113.315 -22.55 ;
      RECT 112.965 -19.44 113.315 -19.32 ;
      RECT 112.965 -16.21 113.315 -16.09 ;
      RECT 112.965 -12.98 113.315 -12.86 ;
      RECT 112.965 -9.75 113.315 -9.63 ;
      RECT 112.965 -6.52 113.315 -6.4 ;
      RECT 112.965 -3.29 113.315 -3.17 ;
      RECT 112.965 -0.06 113.315 0.06 ;
      RECT 113.135 -104.945 113.235 -103.985 ;
      RECT 113.135 2.175 113.235 3.135 ;
      RECT 112.96 -109.595 113.105 -109.275 ;
      RECT 112.875 -104.945 112.975 -103.985 ;
      RECT 112.75 -101.06 112.85 -100.525 ;
      RECT 112.75 -99.735 112.85 -99.2 ;
      RECT 112.75 -97.83 112.85 -97.295 ;
      RECT 112.75 -96.505 112.85 -95.97 ;
      RECT 112.75 -94.6 112.85 -94.065 ;
      RECT 112.75 -93.275 112.85 -92.74 ;
      RECT 112.75 -91.37 112.85 -90.835 ;
      RECT 112.75 -90.045 112.85 -89.51 ;
      RECT 112.75 -88.14 112.85 -87.605 ;
      RECT 112.75 -86.815 112.85 -86.28 ;
      RECT 112.75 -84.91 112.85 -84.375 ;
      RECT 112.75 -83.585 112.85 -83.05 ;
      RECT 112.75 -81.68 112.85 -81.145 ;
      RECT 112.75 -80.355 112.85 -79.82 ;
      RECT 112.75 -78.45 112.85 -77.915 ;
      RECT 112.75 -77.125 112.85 -76.59 ;
      RECT 112.75 -75.22 112.85 -74.685 ;
      RECT 112.75 -73.895 112.85 -73.36 ;
      RECT 112.75 -71.99 112.85 -71.455 ;
      RECT 112.75 -70.665 112.85 -70.13 ;
      RECT 112.75 -68.76 112.85 -68.225 ;
      RECT 112.75 -67.435 112.85 -66.9 ;
      RECT 112.75 -65.53 112.85 -64.995 ;
      RECT 112.75 -64.205 112.85 -63.67 ;
      RECT 112.75 -62.3 112.85 -61.765 ;
      RECT 112.75 -60.975 112.85 -60.44 ;
      RECT 112.75 -59.07 112.85 -58.535 ;
      RECT 112.75 -57.745 112.85 -57.21 ;
      RECT 112.75 -55.84 112.85 -55.305 ;
      RECT 112.75 -54.515 112.85 -53.98 ;
      RECT 112.75 -52.61 112.85 -52.075 ;
      RECT 112.75 -51.285 112.85 -50.75 ;
      RECT 112.75 -49.38 112.85 -48.845 ;
      RECT 112.75 -48.055 112.85 -47.52 ;
      RECT 112.75 -46.15 112.85 -45.615 ;
      RECT 112.75 -44.825 112.85 -44.29 ;
      RECT 112.75 -42.92 112.85 -42.385 ;
      RECT 112.75 -41.595 112.85 -41.06 ;
      RECT 112.75 -39.69 112.85 -39.155 ;
      RECT 112.75 -38.365 112.85 -37.83 ;
      RECT 112.75 -36.46 112.85 -35.925 ;
      RECT 112.75 -35.135 112.85 -34.6 ;
      RECT 112.75 -33.23 112.85 -32.695 ;
      RECT 112.75 -31.905 112.85 -31.37 ;
      RECT 112.75 -30 112.85 -29.465 ;
      RECT 112.75 -28.675 112.85 -28.14 ;
      RECT 112.75 -26.77 112.85 -26.235 ;
      RECT 112.75 -25.445 112.85 -24.91 ;
      RECT 112.75 -23.54 112.85 -23.005 ;
      RECT 112.75 -22.215 112.85 -21.68 ;
      RECT 112.75 -20.31 112.85 -19.775 ;
      RECT 112.75 -18.985 112.85 -18.45 ;
      RECT 112.75 -17.08 112.85 -16.545 ;
      RECT 112.75 -15.755 112.85 -15.22 ;
      RECT 112.75 -13.85 112.85 -13.315 ;
      RECT 112.75 -12.525 112.85 -11.99 ;
      RECT 112.75 -10.62 112.85 -10.085 ;
      RECT 112.75 -9.295 112.85 -8.76 ;
      RECT 112.75 -7.39 112.85 -6.855 ;
      RECT 112.75 -6.065 112.85 -5.53 ;
      RECT 112.75 -4.16 112.85 -3.625 ;
      RECT 112.75 -2.835 112.85 -2.3 ;
      RECT 112.75 -0.93 112.85 -0.395 ;
      RECT 112.75 0.395 112.85 0.93 ;
      RECT 112.625 -108.175 112.725 -107.215 ;
      RECT 112.25 -100.19 112.6 -100.07 ;
      RECT 112.25 -96.96 112.6 -96.84 ;
      RECT 112.25 -93.73 112.6 -93.61 ;
      RECT 112.25 -90.5 112.6 -90.38 ;
      RECT 112.25 -87.27 112.6 -87.15 ;
      RECT 112.25 -84.04 112.6 -83.92 ;
      RECT 112.25 -80.81 112.6 -80.69 ;
      RECT 112.25 -77.58 112.6 -77.46 ;
      RECT 112.25 -74.35 112.6 -74.23 ;
      RECT 112.25 -71.12 112.6 -71 ;
      RECT 112.25 -67.89 112.6 -67.77 ;
      RECT 112.25 -64.66 112.6 -64.54 ;
      RECT 112.25 -61.43 112.6 -61.31 ;
      RECT 112.25 -58.2 112.6 -58.08 ;
      RECT 112.25 -54.97 112.6 -54.85 ;
      RECT 112.25 -51.74 112.6 -51.62 ;
      RECT 112.25 -48.51 112.6 -48.39 ;
      RECT 112.25 -45.28 112.6 -45.16 ;
      RECT 112.25 -42.05 112.6 -41.93 ;
      RECT 112.25 -38.82 112.6 -38.7 ;
      RECT 112.25 -35.59 112.6 -35.47 ;
      RECT 112.25 -32.36 112.6 -32.24 ;
      RECT 112.25 -29.13 112.6 -29.01 ;
      RECT 112.25 -25.9 112.6 -25.78 ;
      RECT 112.25 -22.67 112.6 -22.55 ;
      RECT 112.25 -19.44 112.6 -19.32 ;
      RECT 112.25 -16.21 112.6 -16.09 ;
      RECT 112.25 -12.98 112.6 -12.86 ;
      RECT 112.25 -9.75 112.6 -9.63 ;
      RECT 112.25 -6.52 112.6 -6.4 ;
      RECT 112.25 -3.29 112.6 -3.17 ;
      RECT 112.25 -0.06 112.6 0.06 ;
      RECT 112.455 -112.255 112.555 -111.775 ;
      RECT 112.455 -110.765 112.555 -110.295 ;
      RECT 112.365 -108.175 112.465 -107.215 ;
      RECT 112.365 2.175 112.465 3.135 ;
      RECT 111.765 -100.19 112.115 -100.07 ;
      RECT 111.765 -96.96 112.115 -96.84 ;
      RECT 111.765 -93.73 112.115 -93.61 ;
      RECT 111.765 -90.5 112.115 -90.38 ;
      RECT 111.765 -87.27 112.115 -87.15 ;
      RECT 111.765 -84.04 112.115 -83.92 ;
      RECT 111.765 -80.81 112.115 -80.69 ;
      RECT 111.765 -77.58 112.115 -77.46 ;
      RECT 111.765 -74.35 112.115 -74.23 ;
      RECT 111.765 -71.12 112.115 -71 ;
      RECT 111.765 -67.89 112.115 -67.77 ;
      RECT 111.765 -64.66 112.115 -64.54 ;
      RECT 111.765 -61.43 112.115 -61.31 ;
      RECT 111.765 -58.2 112.115 -58.08 ;
      RECT 111.765 -54.97 112.115 -54.85 ;
      RECT 111.765 -51.74 112.115 -51.62 ;
      RECT 111.765 -48.51 112.115 -48.39 ;
      RECT 111.765 -45.28 112.115 -45.16 ;
      RECT 111.765 -42.05 112.115 -41.93 ;
      RECT 111.765 -38.82 112.115 -38.7 ;
      RECT 111.765 -35.59 112.115 -35.47 ;
      RECT 111.765 -32.36 112.115 -32.24 ;
      RECT 111.765 -29.13 112.115 -29.01 ;
      RECT 111.765 -25.9 112.115 -25.78 ;
      RECT 111.765 -22.67 112.115 -22.55 ;
      RECT 111.765 -19.44 112.115 -19.32 ;
      RECT 111.765 -16.21 112.115 -16.09 ;
      RECT 111.765 -12.98 112.115 -12.86 ;
      RECT 111.765 -9.75 112.115 -9.63 ;
      RECT 111.765 -6.52 112.115 -6.4 ;
      RECT 111.765 -3.29 112.115 -3.17 ;
      RECT 111.765 -0.06 112.115 0.06 ;
      RECT 111.935 -108.175 112.035 -107.215 ;
      RECT 111.935 2.175 112.035 3.135 ;
      RECT 111.83 -110.765 112 -110.385 ;
      RECT 111.865 -112.245 111.965 -111.775 ;
      RECT 111.675 -108.175 111.775 -107.215 ;
      RECT 111.55 -101.06 111.65 -100.525 ;
      RECT 111.55 -99.735 111.65 -99.2 ;
      RECT 111.55 -97.83 111.65 -97.295 ;
      RECT 111.55 -96.505 111.65 -95.97 ;
      RECT 111.55 -94.6 111.65 -94.065 ;
      RECT 111.55 -93.275 111.65 -92.74 ;
      RECT 111.55 -91.37 111.65 -90.835 ;
      RECT 111.55 -90.045 111.65 -89.51 ;
      RECT 111.55 -88.14 111.65 -87.605 ;
      RECT 111.55 -86.815 111.65 -86.28 ;
      RECT 111.55 -84.91 111.65 -84.375 ;
      RECT 111.55 -83.585 111.65 -83.05 ;
      RECT 111.55 -81.68 111.65 -81.145 ;
      RECT 111.55 -80.355 111.65 -79.82 ;
      RECT 111.55 -78.45 111.65 -77.915 ;
      RECT 111.55 -77.125 111.65 -76.59 ;
      RECT 111.55 -75.22 111.65 -74.685 ;
      RECT 111.55 -73.895 111.65 -73.36 ;
      RECT 111.55 -71.99 111.65 -71.455 ;
      RECT 111.55 -70.665 111.65 -70.13 ;
      RECT 111.55 -68.76 111.65 -68.225 ;
      RECT 111.55 -67.435 111.65 -66.9 ;
      RECT 111.55 -65.53 111.65 -64.995 ;
      RECT 111.55 -64.205 111.65 -63.67 ;
      RECT 111.55 -62.3 111.65 -61.765 ;
      RECT 111.55 -60.975 111.65 -60.44 ;
      RECT 111.55 -59.07 111.65 -58.535 ;
      RECT 111.55 -57.745 111.65 -57.21 ;
      RECT 111.55 -55.84 111.65 -55.305 ;
      RECT 111.55 -54.515 111.65 -53.98 ;
      RECT 111.55 -52.61 111.65 -52.075 ;
      RECT 111.55 -51.285 111.65 -50.75 ;
      RECT 111.55 -49.38 111.65 -48.845 ;
      RECT 111.55 -48.055 111.65 -47.52 ;
      RECT 111.55 -46.15 111.65 -45.615 ;
      RECT 111.55 -44.825 111.65 -44.29 ;
      RECT 111.55 -42.92 111.65 -42.385 ;
      RECT 111.55 -41.595 111.65 -41.06 ;
      RECT 111.55 -39.69 111.65 -39.155 ;
      RECT 111.55 -38.365 111.65 -37.83 ;
      RECT 111.55 -36.46 111.65 -35.925 ;
      RECT 111.55 -35.135 111.65 -34.6 ;
      RECT 111.55 -33.23 111.65 -32.695 ;
      RECT 111.55 -31.905 111.65 -31.37 ;
      RECT 111.55 -30 111.65 -29.465 ;
      RECT 111.55 -28.675 111.65 -28.14 ;
      RECT 111.55 -26.77 111.65 -26.235 ;
      RECT 111.55 -25.445 111.65 -24.91 ;
      RECT 111.55 -23.54 111.65 -23.005 ;
      RECT 111.55 -22.215 111.65 -21.68 ;
      RECT 111.55 -20.31 111.65 -19.775 ;
      RECT 111.55 -18.985 111.65 -18.45 ;
      RECT 111.55 -17.08 111.65 -16.545 ;
      RECT 111.55 -15.755 111.65 -15.22 ;
      RECT 111.55 -13.85 111.65 -13.315 ;
      RECT 111.55 -12.525 111.65 -11.99 ;
      RECT 111.55 -10.62 111.65 -10.085 ;
      RECT 111.55 -9.295 111.65 -8.76 ;
      RECT 111.55 -7.39 111.65 -6.855 ;
      RECT 111.55 -6.065 111.65 -5.53 ;
      RECT 111.55 -4.16 111.65 -3.625 ;
      RECT 111.55 -2.835 111.65 -2.3 ;
      RECT 111.55 -0.93 111.65 -0.395 ;
      RECT 111.55 0.395 111.65 0.93 ;
      RECT 111.425 -108.175 111.525 -107.215 ;
      RECT 111.05 -100.19 111.4 -100.07 ;
      RECT 111.05 -96.96 111.4 -96.84 ;
      RECT 111.05 -93.73 111.4 -93.61 ;
      RECT 111.05 -90.5 111.4 -90.38 ;
      RECT 111.05 -87.27 111.4 -87.15 ;
      RECT 111.05 -84.04 111.4 -83.92 ;
      RECT 111.05 -80.81 111.4 -80.69 ;
      RECT 111.05 -77.58 111.4 -77.46 ;
      RECT 111.05 -74.35 111.4 -74.23 ;
      RECT 111.05 -71.12 111.4 -71 ;
      RECT 111.05 -67.89 111.4 -67.77 ;
      RECT 111.05 -64.66 111.4 -64.54 ;
      RECT 111.05 -61.43 111.4 -61.31 ;
      RECT 111.05 -58.2 111.4 -58.08 ;
      RECT 111.05 -54.97 111.4 -54.85 ;
      RECT 111.05 -51.74 111.4 -51.62 ;
      RECT 111.05 -48.51 111.4 -48.39 ;
      RECT 111.05 -45.28 111.4 -45.16 ;
      RECT 111.05 -42.05 111.4 -41.93 ;
      RECT 111.05 -38.82 111.4 -38.7 ;
      RECT 111.05 -35.59 111.4 -35.47 ;
      RECT 111.05 -32.36 111.4 -32.24 ;
      RECT 111.05 -29.13 111.4 -29.01 ;
      RECT 111.05 -25.9 111.4 -25.78 ;
      RECT 111.05 -22.67 111.4 -22.55 ;
      RECT 111.05 -19.44 111.4 -19.32 ;
      RECT 111.05 -16.21 111.4 -16.09 ;
      RECT 111.05 -12.98 111.4 -12.86 ;
      RECT 111.05 -9.75 111.4 -9.63 ;
      RECT 111.05 -6.52 111.4 -6.4 ;
      RECT 111.05 -3.29 111.4 -3.17 ;
      RECT 111.05 -0.06 111.4 0.06 ;
      RECT 111.165 -108.175 111.265 -107.215 ;
      RECT 111.165 2.175 111.265 3.135 ;
      RECT 111.065 -113.555 111.165 -113.085 ;
      RECT 110.565 -100.19 110.915 -100.07 ;
      RECT 110.565 -96.96 110.915 -96.84 ;
      RECT 110.565 -93.73 110.915 -93.61 ;
      RECT 110.565 -90.5 110.915 -90.38 ;
      RECT 110.565 -87.27 110.915 -87.15 ;
      RECT 110.565 -84.04 110.915 -83.92 ;
      RECT 110.565 -80.81 110.915 -80.69 ;
      RECT 110.565 -77.58 110.915 -77.46 ;
      RECT 110.565 -74.35 110.915 -74.23 ;
      RECT 110.565 -71.12 110.915 -71 ;
      RECT 110.565 -67.89 110.915 -67.77 ;
      RECT 110.565 -64.66 110.915 -64.54 ;
      RECT 110.565 -61.43 110.915 -61.31 ;
      RECT 110.565 -58.2 110.915 -58.08 ;
      RECT 110.565 -54.97 110.915 -54.85 ;
      RECT 110.565 -51.74 110.915 -51.62 ;
      RECT 110.565 -48.51 110.915 -48.39 ;
      RECT 110.565 -45.28 110.915 -45.16 ;
      RECT 110.565 -42.05 110.915 -41.93 ;
      RECT 110.565 -38.82 110.915 -38.7 ;
      RECT 110.565 -35.59 110.915 -35.47 ;
      RECT 110.565 -32.36 110.915 -32.24 ;
      RECT 110.565 -29.13 110.915 -29.01 ;
      RECT 110.565 -25.9 110.915 -25.78 ;
      RECT 110.565 -22.67 110.915 -22.55 ;
      RECT 110.565 -19.44 110.915 -19.32 ;
      RECT 110.565 -16.21 110.915 -16.09 ;
      RECT 110.565 -12.98 110.915 -12.86 ;
      RECT 110.565 -9.75 110.915 -9.63 ;
      RECT 110.565 -6.52 110.915 -6.4 ;
      RECT 110.565 -3.29 110.915 -3.17 ;
      RECT 110.565 -0.06 110.915 0.06 ;
      RECT 110.7 -110.735 110.85 -110.445 ;
      RECT 110.735 -108.175 110.835 -107.215 ;
      RECT 110.735 2.175 110.835 3.135 ;
      RECT 110.715 -112.19 110.815 -111.65 ;
      RECT 110.475 -113.555 110.575 -113.085 ;
      RECT 110.475 -108.175 110.575 -107.215 ;
      RECT 110.35 -101.06 110.45 -100.525 ;
      RECT 110.35 -99.735 110.45 -99.2 ;
      RECT 110.35 -97.83 110.45 -97.295 ;
      RECT 110.35 -96.505 110.45 -95.97 ;
      RECT 110.35 -94.6 110.45 -94.065 ;
      RECT 110.35 -93.275 110.45 -92.74 ;
      RECT 110.35 -91.37 110.45 -90.835 ;
      RECT 110.35 -90.045 110.45 -89.51 ;
      RECT 110.35 -88.14 110.45 -87.605 ;
      RECT 110.35 -86.815 110.45 -86.28 ;
      RECT 110.35 -84.91 110.45 -84.375 ;
      RECT 110.35 -83.585 110.45 -83.05 ;
      RECT 110.35 -81.68 110.45 -81.145 ;
      RECT 110.35 -80.355 110.45 -79.82 ;
      RECT 110.35 -78.45 110.45 -77.915 ;
      RECT 110.35 -77.125 110.45 -76.59 ;
      RECT 110.35 -75.22 110.45 -74.685 ;
      RECT 110.35 -73.895 110.45 -73.36 ;
      RECT 110.35 -71.99 110.45 -71.455 ;
      RECT 110.35 -70.665 110.45 -70.13 ;
      RECT 110.35 -68.76 110.45 -68.225 ;
      RECT 110.35 -67.435 110.45 -66.9 ;
      RECT 110.35 -65.53 110.45 -64.995 ;
      RECT 110.35 -64.205 110.45 -63.67 ;
      RECT 110.35 -62.3 110.45 -61.765 ;
      RECT 110.35 -60.975 110.45 -60.44 ;
      RECT 110.35 -59.07 110.45 -58.535 ;
      RECT 110.35 -57.745 110.45 -57.21 ;
      RECT 110.35 -55.84 110.45 -55.305 ;
      RECT 110.35 -54.515 110.45 -53.98 ;
      RECT 110.35 -52.61 110.45 -52.075 ;
      RECT 110.35 -51.285 110.45 -50.75 ;
      RECT 110.35 -49.38 110.45 -48.845 ;
      RECT 110.35 -48.055 110.45 -47.52 ;
      RECT 110.35 -46.15 110.45 -45.615 ;
      RECT 110.35 -44.825 110.45 -44.29 ;
      RECT 110.35 -42.92 110.45 -42.385 ;
      RECT 110.35 -41.595 110.45 -41.06 ;
      RECT 110.35 -39.69 110.45 -39.155 ;
      RECT 110.35 -38.365 110.45 -37.83 ;
      RECT 110.35 -36.46 110.45 -35.925 ;
      RECT 110.35 -35.135 110.45 -34.6 ;
      RECT 110.35 -33.23 110.45 -32.695 ;
      RECT 110.35 -31.905 110.45 -31.37 ;
      RECT 110.35 -30 110.45 -29.465 ;
      RECT 110.35 -28.675 110.45 -28.14 ;
      RECT 110.35 -26.77 110.45 -26.235 ;
      RECT 110.35 -25.445 110.45 -24.91 ;
      RECT 110.35 -23.54 110.45 -23.005 ;
      RECT 110.35 -22.215 110.45 -21.68 ;
      RECT 110.35 -20.31 110.45 -19.775 ;
      RECT 110.35 -18.985 110.45 -18.45 ;
      RECT 110.35 -17.08 110.45 -16.545 ;
      RECT 110.35 -15.755 110.45 -15.22 ;
      RECT 110.35 -13.85 110.45 -13.315 ;
      RECT 110.35 -12.525 110.45 -11.99 ;
      RECT 110.35 -10.62 110.45 -10.085 ;
      RECT 110.35 -9.295 110.45 -8.76 ;
      RECT 110.35 -7.39 110.45 -6.855 ;
      RECT 110.35 -6.065 110.45 -5.53 ;
      RECT 110.35 -4.16 110.45 -3.625 ;
      RECT 110.35 -2.835 110.45 -2.3 ;
      RECT 110.35 -0.93 110.45 -0.395 ;
      RECT 110.35 0.395 110.45 0.93 ;
      RECT 110.225 -104.945 110.325 -103.985 ;
      RECT 109.85 -100.19 110.2 -100.07 ;
      RECT 109.85 -96.96 110.2 -96.84 ;
      RECT 109.85 -93.73 110.2 -93.61 ;
      RECT 109.85 -90.5 110.2 -90.38 ;
      RECT 109.85 -87.27 110.2 -87.15 ;
      RECT 109.85 -84.04 110.2 -83.92 ;
      RECT 109.85 -80.81 110.2 -80.69 ;
      RECT 109.85 -77.58 110.2 -77.46 ;
      RECT 109.85 -74.35 110.2 -74.23 ;
      RECT 109.85 -71.12 110.2 -71 ;
      RECT 109.85 -67.89 110.2 -67.77 ;
      RECT 109.85 -64.66 110.2 -64.54 ;
      RECT 109.85 -61.43 110.2 -61.31 ;
      RECT 109.85 -58.2 110.2 -58.08 ;
      RECT 109.85 -54.97 110.2 -54.85 ;
      RECT 109.85 -51.74 110.2 -51.62 ;
      RECT 109.85 -48.51 110.2 -48.39 ;
      RECT 109.85 -45.28 110.2 -45.16 ;
      RECT 109.85 -42.05 110.2 -41.93 ;
      RECT 109.85 -38.82 110.2 -38.7 ;
      RECT 109.85 -35.59 110.2 -35.47 ;
      RECT 109.85 -32.36 110.2 -32.24 ;
      RECT 109.85 -29.13 110.2 -29.01 ;
      RECT 109.85 -25.9 110.2 -25.78 ;
      RECT 109.85 -22.67 110.2 -22.55 ;
      RECT 109.85 -19.44 110.2 -19.32 ;
      RECT 109.85 -16.21 110.2 -16.09 ;
      RECT 109.85 -12.98 110.2 -12.86 ;
      RECT 109.85 -9.75 110.2 -9.63 ;
      RECT 109.85 -6.52 110.2 -6.4 ;
      RECT 109.85 -3.29 110.2 -3.17 ;
      RECT 109.85 -0.06 110.2 0.06 ;
      RECT 109.965 -104.945 110.065 -103.985 ;
      RECT 109.965 2.175 110.065 3.135 ;
      RECT 109.675 -112.255 109.775 -111.775 ;
      RECT 109.675 -110.765 109.775 -110.295 ;
      RECT 109.365 -100.19 109.715 -100.07 ;
      RECT 109.365 -96.96 109.715 -96.84 ;
      RECT 109.365 -93.73 109.715 -93.61 ;
      RECT 109.365 -90.5 109.715 -90.38 ;
      RECT 109.365 -87.27 109.715 -87.15 ;
      RECT 109.365 -84.04 109.715 -83.92 ;
      RECT 109.365 -80.81 109.715 -80.69 ;
      RECT 109.365 -77.58 109.715 -77.46 ;
      RECT 109.365 -74.35 109.715 -74.23 ;
      RECT 109.365 -71.12 109.715 -71 ;
      RECT 109.365 -67.89 109.715 -67.77 ;
      RECT 109.365 -64.66 109.715 -64.54 ;
      RECT 109.365 -61.43 109.715 -61.31 ;
      RECT 109.365 -58.2 109.715 -58.08 ;
      RECT 109.365 -54.97 109.715 -54.85 ;
      RECT 109.365 -51.74 109.715 -51.62 ;
      RECT 109.365 -48.51 109.715 -48.39 ;
      RECT 109.365 -45.28 109.715 -45.16 ;
      RECT 109.365 -42.05 109.715 -41.93 ;
      RECT 109.365 -38.82 109.715 -38.7 ;
      RECT 109.365 -35.59 109.715 -35.47 ;
      RECT 109.365 -32.36 109.715 -32.24 ;
      RECT 109.365 -29.13 109.715 -29.01 ;
      RECT 109.365 -25.9 109.715 -25.78 ;
      RECT 109.365 -22.67 109.715 -22.55 ;
      RECT 109.365 -19.44 109.715 -19.32 ;
      RECT 109.365 -16.21 109.715 -16.09 ;
      RECT 109.365 -12.98 109.715 -12.86 ;
      RECT 109.365 -9.75 109.715 -9.63 ;
      RECT 109.365 -6.52 109.715 -6.4 ;
      RECT 109.365 -3.29 109.715 -3.17 ;
      RECT 109.365 -0.06 109.715 0.06 ;
      RECT 109.535 -104.945 109.635 -103.985 ;
      RECT 109.535 2.175 109.635 3.135 ;
      RECT 105.635 -108.655 109.415 -108.535 ;
      RECT 109.275 -104.945 109.375 -103.985 ;
      RECT 109.15 -101.06 109.25 -100.525 ;
      RECT 109.15 -99.735 109.25 -99.2 ;
      RECT 109.15 -97.83 109.25 -97.295 ;
      RECT 109.15 -96.505 109.25 -95.97 ;
      RECT 109.15 -94.6 109.25 -94.065 ;
      RECT 109.15 -93.275 109.25 -92.74 ;
      RECT 109.15 -91.37 109.25 -90.835 ;
      RECT 109.15 -90.045 109.25 -89.51 ;
      RECT 109.15 -88.14 109.25 -87.605 ;
      RECT 109.15 -86.815 109.25 -86.28 ;
      RECT 109.15 -84.91 109.25 -84.375 ;
      RECT 109.15 -83.585 109.25 -83.05 ;
      RECT 109.15 -81.68 109.25 -81.145 ;
      RECT 109.15 -80.355 109.25 -79.82 ;
      RECT 109.15 -78.45 109.25 -77.915 ;
      RECT 109.15 -77.125 109.25 -76.59 ;
      RECT 109.15 -75.22 109.25 -74.685 ;
      RECT 109.15 -73.895 109.25 -73.36 ;
      RECT 109.15 -71.99 109.25 -71.455 ;
      RECT 109.15 -70.665 109.25 -70.13 ;
      RECT 109.15 -68.76 109.25 -68.225 ;
      RECT 109.15 -67.435 109.25 -66.9 ;
      RECT 109.15 -65.53 109.25 -64.995 ;
      RECT 109.15 -64.205 109.25 -63.67 ;
      RECT 109.15 -62.3 109.25 -61.765 ;
      RECT 109.15 -60.975 109.25 -60.44 ;
      RECT 109.15 -59.07 109.25 -58.535 ;
      RECT 109.15 -57.745 109.25 -57.21 ;
      RECT 109.15 -55.84 109.25 -55.305 ;
      RECT 109.15 -54.515 109.25 -53.98 ;
      RECT 109.15 -52.61 109.25 -52.075 ;
      RECT 109.15 -51.285 109.25 -50.75 ;
      RECT 109.15 -49.38 109.25 -48.845 ;
      RECT 109.15 -48.055 109.25 -47.52 ;
      RECT 109.15 -46.15 109.25 -45.615 ;
      RECT 109.15 -44.825 109.25 -44.29 ;
      RECT 109.15 -42.92 109.25 -42.385 ;
      RECT 109.15 -41.595 109.25 -41.06 ;
      RECT 109.15 -39.69 109.25 -39.155 ;
      RECT 109.15 -38.365 109.25 -37.83 ;
      RECT 109.15 -36.46 109.25 -35.925 ;
      RECT 109.15 -35.135 109.25 -34.6 ;
      RECT 109.15 -33.23 109.25 -32.695 ;
      RECT 109.15 -31.905 109.25 -31.37 ;
      RECT 109.15 -30 109.25 -29.465 ;
      RECT 109.15 -28.675 109.25 -28.14 ;
      RECT 109.15 -26.77 109.25 -26.235 ;
      RECT 109.15 -25.445 109.25 -24.91 ;
      RECT 109.15 -23.54 109.25 -23.005 ;
      RECT 109.15 -22.215 109.25 -21.68 ;
      RECT 109.15 -20.31 109.25 -19.775 ;
      RECT 109.15 -18.985 109.25 -18.45 ;
      RECT 109.15 -17.08 109.25 -16.545 ;
      RECT 109.15 -15.755 109.25 -15.22 ;
      RECT 109.15 -13.85 109.25 -13.315 ;
      RECT 109.15 -12.525 109.25 -11.99 ;
      RECT 109.15 -10.62 109.25 -10.085 ;
      RECT 109.15 -9.295 109.25 -8.76 ;
      RECT 109.15 -7.39 109.25 -6.855 ;
      RECT 109.15 -6.065 109.25 -5.53 ;
      RECT 109.15 -4.16 109.25 -3.625 ;
      RECT 109.15 -2.835 109.25 -2.3 ;
      RECT 109.15 -0.93 109.25 -0.395 ;
      RECT 109.15 0.395 109.25 0.93 ;
      RECT 109.085 -110.75 109.205 -110.37 ;
      RECT 109.085 -112.245 109.185 -111.775 ;
      RECT 109.025 -104.945 109.125 -103.985 ;
      RECT 108.65 -100.19 109 -100.07 ;
      RECT 108.65 -96.96 109 -96.84 ;
      RECT 108.65 -93.73 109 -93.61 ;
      RECT 108.65 -90.5 109 -90.38 ;
      RECT 108.65 -87.27 109 -87.15 ;
      RECT 108.65 -84.04 109 -83.92 ;
      RECT 108.65 -80.81 109 -80.69 ;
      RECT 108.65 -77.58 109 -77.46 ;
      RECT 108.65 -74.35 109 -74.23 ;
      RECT 108.65 -71.12 109 -71 ;
      RECT 108.65 -67.89 109 -67.77 ;
      RECT 108.65 -64.66 109 -64.54 ;
      RECT 108.65 -61.43 109 -61.31 ;
      RECT 108.65 -58.2 109 -58.08 ;
      RECT 108.65 -54.97 109 -54.85 ;
      RECT 108.65 -51.74 109 -51.62 ;
      RECT 108.65 -48.51 109 -48.39 ;
      RECT 108.65 -45.28 109 -45.16 ;
      RECT 108.65 -42.05 109 -41.93 ;
      RECT 108.65 -38.82 109 -38.7 ;
      RECT 108.65 -35.59 109 -35.47 ;
      RECT 108.65 -32.36 109 -32.24 ;
      RECT 108.65 -29.13 109 -29.01 ;
      RECT 108.65 -25.9 109 -25.78 ;
      RECT 108.65 -22.67 109 -22.55 ;
      RECT 108.65 -19.44 109 -19.32 ;
      RECT 108.65 -16.21 109 -16.09 ;
      RECT 108.65 -12.98 109 -12.86 ;
      RECT 108.65 -9.75 109 -9.63 ;
      RECT 108.65 -6.52 109 -6.4 ;
      RECT 108.65 -3.29 109 -3.17 ;
      RECT 108.65 -0.06 109 0.06 ;
      RECT 108.765 -104.945 108.865 -103.985 ;
      RECT 108.765 2.175 108.865 3.135 ;
      RECT 108.495 -109.595 108.63 -109.275 ;
      RECT 108.165 -100.19 108.515 -100.07 ;
      RECT 108.165 -96.96 108.515 -96.84 ;
      RECT 108.165 -93.73 108.515 -93.61 ;
      RECT 108.165 -90.5 108.515 -90.38 ;
      RECT 108.165 -87.27 108.515 -87.15 ;
      RECT 108.165 -84.04 108.515 -83.92 ;
      RECT 108.165 -80.81 108.515 -80.69 ;
      RECT 108.165 -77.58 108.515 -77.46 ;
      RECT 108.165 -74.35 108.515 -74.23 ;
      RECT 108.165 -71.12 108.515 -71 ;
      RECT 108.165 -67.89 108.515 -67.77 ;
      RECT 108.165 -64.66 108.515 -64.54 ;
      RECT 108.165 -61.43 108.515 -61.31 ;
      RECT 108.165 -58.2 108.515 -58.08 ;
      RECT 108.165 -54.97 108.515 -54.85 ;
      RECT 108.165 -51.74 108.515 -51.62 ;
      RECT 108.165 -48.51 108.515 -48.39 ;
      RECT 108.165 -45.28 108.515 -45.16 ;
      RECT 108.165 -42.05 108.515 -41.93 ;
      RECT 108.165 -38.82 108.515 -38.7 ;
      RECT 108.165 -35.59 108.515 -35.47 ;
      RECT 108.165 -32.36 108.515 -32.24 ;
      RECT 108.165 -29.13 108.515 -29.01 ;
      RECT 108.165 -25.9 108.515 -25.78 ;
      RECT 108.165 -22.67 108.515 -22.55 ;
      RECT 108.165 -19.44 108.515 -19.32 ;
      RECT 108.165 -16.21 108.515 -16.09 ;
      RECT 108.165 -12.98 108.515 -12.86 ;
      RECT 108.165 -9.75 108.515 -9.63 ;
      RECT 108.165 -6.52 108.515 -6.4 ;
      RECT 108.165 -3.29 108.515 -3.17 ;
      RECT 108.165 -0.06 108.515 0.06 ;
      RECT 108.335 -104.945 108.435 -103.985 ;
      RECT 108.335 2.175 108.435 3.135 ;
      RECT 108.16 -109.595 108.305 -109.275 ;
      RECT 108.075 -104.945 108.175 -103.985 ;
      RECT 107.95 -101.06 108.05 -100.525 ;
      RECT 107.95 -99.735 108.05 -99.2 ;
      RECT 107.95 -97.83 108.05 -97.295 ;
      RECT 107.95 -96.505 108.05 -95.97 ;
      RECT 107.95 -94.6 108.05 -94.065 ;
      RECT 107.95 -93.275 108.05 -92.74 ;
      RECT 107.95 -91.37 108.05 -90.835 ;
      RECT 107.95 -90.045 108.05 -89.51 ;
      RECT 107.95 -88.14 108.05 -87.605 ;
      RECT 107.95 -86.815 108.05 -86.28 ;
      RECT 107.95 -84.91 108.05 -84.375 ;
      RECT 107.95 -83.585 108.05 -83.05 ;
      RECT 107.95 -81.68 108.05 -81.145 ;
      RECT 107.95 -80.355 108.05 -79.82 ;
      RECT 107.95 -78.45 108.05 -77.915 ;
      RECT 107.95 -77.125 108.05 -76.59 ;
      RECT 107.95 -75.22 108.05 -74.685 ;
      RECT 107.95 -73.895 108.05 -73.36 ;
      RECT 107.95 -71.99 108.05 -71.455 ;
      RECT 107.95 -70.665 108.05 -70.13 ;
      RECT 107.95 -68.76 108.05 -68.225 ;
      RECT 107.95 -67.435 108.05 -66.9 ;
      RECT 107.95 -65.53 108.05 -64.995 ;
      RECT 107.95 -64.205 108.05 -63.67 ;
      RECT 107.95 -62.3 108.05 -61.765 ;
      RECT 107.95 -60.975 108.05 -60.44 ;
      RECT 107.95 -59.07 108.05 -58.535 ;
      RECT 107.95 -57.745 108.05 -57.21 ;
      RECT 107.95 -55.84 108.05 -55.305 ;
      RECT 107.95 -54.515 108.05 -53.98 ;
      RECT 107.95 -52.61 108.05 -52.075 ;
      RECT 107.95 -51.285 108.05 -50.75 ;
      RECT 107.95 -49.38 108.05 -48.845 ;
      RECT 107.95 -48.055 108.05 -47.52 ;
      RECT 107.95 -46.15 108.05 -45.615 ;
      RECT 107.95 -44.825 108.05 -44.29 ;
      RECT 107.95 -42.92 108.05 -42.385 ;
      RECT 107.95 -41.595 108.05 -41.06 ;
      RECT 107.95 -39.69 108.05 -39.155 ;
      RECT 107.95 -38.365 108.05 -37.83 ;
      RECT 107.95 -36.46 108.05 -35.925 ;
      RECT 107.95 -35.135 108.05 -34.6 ;
      RECT 107.95 -33.23 108.05 -32.695 ;
      RECT 107.95 -31.905 108.05 -31.37 ;
      RECT 107.95 -30 108.05 -29.465 ;
      RECT 107.95 -28.675 108.05 -28.14 ;
      RECT 107.95 -26.77 108.05 -26.235 ;
      RECT 107.95 -25.445 108.05 -24.91 ;
      RECT 107.95 -23.54 108.05 -23.005 ;
      RECT 107.95 -22.215 108.05 -21.68 ;
      RECT 107.95 -20.31 108.05 -19.775 ;
      RECT 107.95 -18.985 108.05 -18.45 ;
      RECT 107.95 -17.08 108.05 -16.545 ;
      RECT 107.95 -15.755 108.05 -15.22 ;
      RECT 107.95 -13.85 108.05 -13.315 ;
      RECT 107.95 -12.525 108.05 -11.99 ;
      RECT 107.95 -10.62 108.05 -10.085 ;
      RECT 107.95 -9.295 108.05 -8.76 ;
      RECT 107.95 -7.39 108.05 -6.855 ;
      RECT 107.95 -6.065 108.05 -5.53 ;
      RECT 107.95 -4.16 108.05 -3.625 ;
      RECT 107.95 -2.835 108.05 -2.3 ;
      RECT 107.95 -0.93 108.05 -0.395 ;
      RECT 107.95 0.395 108.05 0.93 ;
      RECT 107.825 -108.175 107.925 -107.215 ;
      RECT 107.45 -100.19 107.8 -100.07 ;
      RECT 107.45 -96.96 107.8 -96.84 ;
      RECT 107.45 -93.73 107.8 -93.61 ;
      RECT 107.45 -90.5 107.8 -90.38 ;
      RECT 107.45 -87.27 107.8 -87.15 ;
      RECT 107.45 -84.04 107.8 -83.92 ;
      RECT 107.45 -80.81 107.8 -80.69 ;
      RECT 107.45 -77.58 107.8 -77.46 ;
      RECT 107.45 -74.35 107.8 -74.23 ;
      RECT 107.45 -71.12 107.8 -71 ;
      RECT 107.45 -67.89 107.8 -67.77 ;
      RECT 107.45 -64.66 107.8 -64.54 ;
      RECT 107.45 -61.43 107.8 -61.31 ;
      RECT 107.45 -58.2 107.8 -58.08 ;
      RECT 107.45 -54.97 107.8 -54.85 ;
      RECT 107.45 -51.74 107.8 -51.62 ;
      RECT 107.45 -48.51 107.8 -48.39 ;
      RECT 107.45 -45.28 107.8 -45.16 ;
      RECT 107.45 -42.05 107.8 -41.93 ;
      RECT 107.45 -38.82 107.8 -38.7 ;
      RECT 107.45 -35.59 107.8 -35.47 ;
      RECT 107.45 -32.36 107.8 -32.24 ;
      RECT 107.45 -29.13 107.8 -29.01 ;
      RECT 107.45 -25.9 107.8 -25.78 ;
      RECT 107.45 -22.67 107.8 -22.55 ;
      RECT 107.45 -19.44 107.8 -19.32 ;
      RECT 107.45 -16.21 107.8 -16.09 ;
      RECT 107.45 -12.98 107.8 -12.86 ;
      RECT 107.45 -9.75 107.8 -9.63 ;
      RECT 107.45 -6.52 107.8 -6.4 ;
      RECT 107.45 -3.29 107.8 -3.17 ;
      RECT 107.45 -0.06 107.8 0.06 ;
      RECT 107.655 -112.255 107.755 -111.775 ;
      RECT 107.655 -110.765 107.755 -110.295 ;
      RECT 107.565 -108.175 107.665 -107.215 ;
      RECT 107.565 2.175 107.665 3.135 ;
      RECT 106.965 -100.19 107.315 -100.07 ;
      RECT 106.965 -96.96 107.315 -96.84 ;
      RECT 106.965 -93.73 107.315 -93.61 ;
      RECT 106.965 -90.5 107.315 -90.38 ;
      RECT 106.965 -87.27 107.315 -87.15 ;
      RECT 106.965 -84.04 107.315 -83.92 ;
      RECT 106.965 -80.81 107.315 -80.69 ;
      RECT 106.965 -77.58 107.315 -77.46 ;
      RECT 106.965 -74.35 107.315 -74.23 ;
      RECT 106.965 -71.12 107.315 -71 ;
      RECT 106.965 -67.89 107.315 -67.77 ;
      RECT 106.965 -64.66 107.315 -64.54 ;
      RECT 106.965 -61.43 107.315 -61.31 ;
      RECT 106.965 -58.2 107.315 -58.08 ;
      RECT 106.965 -54.97 107.315 -54.85 ;
      RECT 106.965 -51.74 107.315 -51.62 ;
      RECT 106.965 -48.51 107.315 -48.39 ;
      RECT 106.965 -45.28 107.315 -45.16 ;
      RECT 106.965 -42.05 107.315 -41.93 ;
      RECT 106.965 -38.82 107.315 -38.7 ;
      RECT 106.965 -35.59 107.315 -35.47 ;
      RECT 106.965 -32.36 107.315 -32.24 ;
      RECT 106.965 -29.13 107.315 -29.01 ;
      RECT 106.965 -25.9 107.315 -25.78 ;
      RECT 106.965 -22.67 107.315 -22.55 ;
      RECT 106.965 -19.44 107.315 -19.32 ;
      RECT 106.965 -16.21 107.315 -16.09 ;
      RECT 106.965 -12.98 107.315 -12.86 ;
      RECT 106.965 -9.75 107.315 -9.63 ;
      RECT 106.965 -6.52 107.315 -6.4 ;
      RECT 106.965 -3.29 107.315 -3.17 ;
      RECT 106.965 -0.06 107.315 0.06 ;
      RECT 107.135 -108.175 107.235 -107.215 ;
      RECT 107.135 2.175 107.235 3.135 ;
      RECT 107.03 -110.765 107.2 -110.385 ;
      RECT 107.065 -112.245 107.165 -111.775 ;
      RECT 106.875 -108.175 106.975 -107.215 ;
      RECT 106.75 -101.06 106.85 -100.525 ;
      RECT 106.75 -99.735 106.85 -99.2 ;
      RECT 106.75 -97.83 106.85 -97.295 ;
      RECT 106.75 -96.505 106.85 -95.97 ;
      RECT 106.75 -94.6 106.85 -94.065 ;
      RECT 106.75 -93.275 106.85 -92.74 ;
      RECT 106.75 -91.37 106.85 -90.835 ;
      RECT 106.75 -90.045 106.85 -89.51 ;
      RECT 106.75 -88.14 106.85 -87.605 ;
      RECT 106.75 -86.815 106.85 -86.28 ;
      RECT 106.75 -84.91 106.85 -84.375 ;
      RECT 106.75 -83.585 106.85 -83.05 ;
      RECT 106.75 -81.68 106.85 -81.145 ;
      RECT 106.75 -80.355 106.85 -79.82 ;
      RECT 106.75 -78.45 106.85 -77.915 ;
      RECT 106.75 -77.125 106.85 -76.59 ;
      RECT 106.75 -75.22 106.85 -74.685 ;
      RECT 106.75 -73.895 106.85 -73.36 ;
      RECT 106.75 -71.99 106.85 -71.455 ;
      RECT 106.75 -70.665 106.85 -70.13 ;
      RECT 106.75 -68.76 106.85 -68.225 ;
      RECT 106.75 -67.435 106.85 -66.9 ;
      RECT 106.75 -65.53 106.85 -64.995 ;
      RECT 106.75 -64.205 106.85 -63.67 ;
      RECT 106.75 -62.3 106.85 -61.765 ;
      RECT 106.75 -60.975 106.85 -60.44 ;
      RECT 106.75 -59.07 106.85 -58.535 ;
      RECT 106.75 -57.745 106.85 -57.21 ;
      RECT 106.75 -55.84 106.85 -55.305 ;
      RECT 106.75 -54.515 106.85 -53.98 ;
      RECT 106.75 -52.61 106.85 -52.075 ;
      RECT 106.75 -51.285 106.85 -50.75 ;
      RECT 106.75 -49.38 106.85 -48.845 ;
      RECT 106.75 -48.055 106.85 -47.52 ;
      RECT 106.75 -46.15 106.85 -45.615 ;
      RECT 106.75 -44.825 106.85 -44.29 ;
      RECT 106.75 -42.92 106.85 -42.385 ;
      RECT 106.75 -41.595 106.85 -41.06 ;
      RECT 106.75 -39.69 106.85 -39.155 ;
      RECT 106.75 -38.365 106.85 -37.83 ;
      RECT 106.75 -36.46 106.85 -35.925 ;
      RECT 106.75 -35.135 106.85 -34.6 ;
      RECT 106.75 -33.23 106.85 -32.695 ;
      RECT 106.75 -31.905 106.85 -31.37 ;
      RECT 106.75 -30 106.85 -29.465 ;
      RECT 106.75 -28.675 106.85 -28.14 ;
      RECT 106.75 -26.77 106.85 -26.235 ;
      RECT 106.75 -25.445 106.85 -24.91 ;
      RECT 106.75 -23.54 106.85 -23.005 ;
      RECT 106.75 -22.215 106.85 -21.68 ;
      RECT 106.75 -20.31 106.85 -19.775 ;
      RECT 106.75 -18.985 106.85 -18.45 ;
      RECT 106.75 -17.08 106.85 -16.545 ;
      RECT 106.75 -15.755 106.85 -15.22 ;
      RECT 106.75 -13.85 106.85 -13.315 ;
      RECT 106.75 -12.525 106.85 -11.99 ;
      RECT 106.75 -10.62 106.85 -10.085 ;
      RECT 106.75 -9.295 106.85 -8.76 ;
      RECT 106.75 -7.39 106.85 -6.855 ;
      RECT 106.75 -6.065 106.85 -5.53 ;
      RECT 106.75 -4.16 106.85 -3.625 ;
      RECT 106.75 -2.835 106.85 -2.3 ;
      RECT 106.75 -0.93 106.85 -0.395 ;
      RECT 106.75 0.395 106.85 0.93 ;
      RECT 106.625 -108.175 106.725 -107.215 ;
      RECT 106.25 -100.19 106.6 -100.07 ;
      RECT 106.25 -96.96 106.6 -96.84 ;
      RECT 106.25 -93.73 106.6 -93.61 ;
      RECT 106.25 -90.5 106.6 -90.38 ;
      RECT 106.25 -87.27 106.6 -87.15 ;
      RECT 106.25 -84.04 106.6 -83.92 ;
      RECT 106.25 -80.81 106.6 -80.69 ;
      RECT 106.25 -77.58 106.6 -77.46 ;
      RECT 106.25 -74.35 106.6 -74.23 ;
      RECT 106.25 -71.12 106.6 -71 ;
      RECT 106.25 -67.89 106.6 -67.77 ;
      RECT 106.25 -64.66 106.6 -64.54 ;
      RECT 106.25 -61.43 106.6 -61.31 ;
      RECT 106.25 -58.2 106.6 -58.08 ;
      RECT 106.25 -54.97 106.6 -54.85 ;
      RECT 106.25 -51.74 106.6 -51.62 ;
      RECT 106.25 -48.51 106.6 -48.39 ;
      RECT 106.25 -45.28 106.6 -45.16 ;
      RECT 106.25 -42.05 106.6 -41.93 ;
      RECT 106.25 -38.82 106.6 -38.7 ;
      RECT 106.25 -35.59 106.6 -35.47 ;
      RECT 106.25 -32.36 106.6 -32.24 ;
      RECT 106.25 -29.13 106.6 -29.01 ;
      RECT 106.25 -25.9 106.6 -25.78 ;
      RECT 106.25 -22.67 106.6 -22.55 ;
      RECT 106.25 -19.44 106.6 -19.32 ;
      RECT 106.25 -16.21 106.6 -16.09 ;
      RECT 106.25 -12.98 106.6 -12.86 ;
      RECT 106.25 -9.75 106.6 -9.63 ;
      RECT 106.25 -6.52 106.6 -6.4 ;
      RECT 106.25 -3.29 106.6 -3.17 ;
      RECT 106.25 -0.06 106.6 0.06 ;
      RECT 106.365 -108.175 106.465 -107.215 ;
      RECT 106.365 2.175 106.465 3.135 ;
      RECT 106.265 -113.555 106.365 -113.085 ;
      RECT 105.765 -100.19 106.115 -100.07 ;
      RECT 105.765 -96.96 106.115 -96.84 ;
      RECT 105.765 -93.73 106.115 -93.61 ;
      RECT 105.765 -90.5 106.115 -90.38 ;
      RECT 105.765 -87.27 106.115 -87.15 ;
      RECT 105.765 -84.04 106.115 -83.92 ;
      RECT 105.765 -80.81 106.115 -80.69 ;
      RECT 105.765 -77.58 106.115 -77.46 ;
      RECT 105.765 -74.35 106.115 -74.23 ;
      RECT 105.765 -71.12 106.115 -71 ;
      RECT 105.765 -67.89 106.115 -67.77 ;
      RECT 105.765 -64.66 106.115 -64.54 ;
      RECT 105.765 -61.43 106.115 -61.31 ;
      RECT 105.765 -58.2 106.115 -58.08 ;
      RECT 105.765 -54.97 106.115 -54.85 ;
      RECT 105.765 -51.74 106.115 -51.62 ;
      RECT 105.765 -48.51 106.115 -48.39 ;
      RECT 105.765 -45.28 106.115 -45.16 ;
      RECT 105.765 -42.05 106.115 -41.93 ;
      RECT 105.765 -38.82 106.115 -38.7 ;
      RECT 105.765 -35.59 106.115 -35.47 ;
      RECT 105.765 -32.36 106.115 -32.24 ;
      RECT 105.765 -29.13 106.115 -29.01 ;
      RECT 105.765 -25.9 106.115 -25.78 ;
      RECT 105.765 -22.67 106.115 -22.55 ;
      RECT 105.765 -19.44 106.115 -19.32 ;
      RECT 105.765 -16.21 106.115 -16.09 ;
      RECT 105.765 -12.98 106.115 -12.86 ;
      RECT 105.765 -9.75 106.115 -9.63 ;
      RECT 105.765 -6.52 106.115 -6.4 ;
      RECT 105.765 -3.29 106.115 -3.17 ;
      RECT 105.765 -0.06 106.115 0.06 ;
      RECT 105.9 -110.735 106.05 -110.445 ;
      RECT 105.935 -108.175 106.035 -107.215 ;
      RECT 105.935 2.175 106.035 3.135 ;
      RECT 105.915 -112.19 106.015 -111.65 ;
      RECT 105.675 -113.555 105.775 -113.085 ;
      RECT 105.675 -108.175 105.775 -107.215 ;
      RECT 105.55 -101.06 105.65 -100.525 ;
      RECT 105.55 -99.735 105.65 -99.2 ;
      RECT 105.55 -97.83 105.65 -97.295 ;
      RECT 105.55 -96.505 105.65 -95.97 ;
      RECT 105.55 -94.6 105.65 -94.065 ;
      RECT 105.55 -93.275 105.65 -92.74 ;
      RECT 105.55 -91.37 105.65 -90.835 ;
      RECT 105.55 -90.045 105.65 -89.51 ;
      RECT 105.55 -88.14 105.65 -87.605 ;
      RECT 105.55 -86.815 105.65 -86.28 ;
      RECT 105.55 -84.91 105.65 -84.375 ;
      RECT 105.55 -83.585 105.65 -83.05 ;
      RECT 105.55 -81.68 105.65 -81.145 ;
      RECT 105.55 -80.355 105.65 -79.82 ;
      RECT 105.55 -78.45 105.65 -77.915 ;
      RECT 105.55 -77.125 105.65 -76.59 ;
      RECT 105.55 -75.22 105.65 -74.685 ;
      RECT 105.55 -73.895 105.65 -73.36 ;
      RECT 105.55 -71.99 105.65 -71.455 ;
      RECT 105.55 -70.665 105.65 -70.13 ;
      RECT 105.55 -68.76 105.65 -68.225 ;
      RECT 105.55 -67.435 105.65 -66.9 ;
      RECT 105.55 -65.53 105.65 -64.995 ;
      RECT 105.55 -64.205 105.65 -63.67 ;
      RECT 105.55 -62.3 105.65 -61.765 ;
      RECT 105.55 -60.975 105.65 -60.44 ;
      RECT 105.55 -59.07 105.65 -58.535 ;
      RECT 105.55 -57.745 105.65 -57.21 ;
      RECT 105.55 -55.84 105.65 -55.305 ;
      RECT 105.55 -54.515 105.65 -53.98 ;
      RECT 105.55 -52.61 105.65 -52.075 ;
      RECT 105.55 -51.285 105.65 -50.75 ;
      RECT 105.55 -49.38 105.65 -48.845 ;
      RECT 105.55 -48.055 105.65 -47.52 ;
      RECT 105.55 -46.15 105.65 -45.615 ;
      RECT 105.55 -44.825 105.65 -44.29 ;
      RECT 105.55 -42.92 105.65 -42.385 ;
      RECT 105.55 -41.595 105.65 -41.06 ;
      RECT 105.55 -39.69 105.65 -39.155 ;
      RECT 105.55 -38.365 105.65 -37.83 ;
      RECT 105.55 -36.46 105.65 -35.925 ;
      RECT 105.55 -35.135 105.65 -34.6 ;
      RECT 105.55 -33.23 105.65 -32.695 ;
      RECT 105.55 -31.905 105.65 -31.37 ;
      RECT 105.55 -30 105.65 -29.465 ;
      RECT 105.55 -28.675 105.65 -28.14 ;
      RECT 105.55 -26.77 105.65 -26.235 ;
      RECT 105.55 -25.445 105.65 -24.91 ;
      RECT 105.55 -23.54 105.65 -23.005 ;
      RECT 105.55 -22.215 105.65 -21.68 ;
      RECT 105.55 -20.31 105.65 -19.775 ;
      RECT 105.55 -18.985 105.65 -18.45 ;
      RECT 105.55 -17.08 105.65 -16.545 ;
      RECT 105.55 -15.755 105.65 -15.22 ;
      RECT 105.55 -13.85 105.65 -13.315 ;
      RECT 105.55 -12.525 105.65 -11.99 ;
      RECT 105.55 -10.62 105.65 -10.085 ;
      RECT 105.55 -9.295 105.65 -8.76 ;
      RECT 105.55 -7.39 105.65 -6.855 ;
      RECT 105.55 -6.065 105.65 -5.53 ;
      RECT 105.55 -4.16 105.65 -3.625 ;
      RECT 105.55 -2.835 105.65 -2.3 ;
      RECT 105.55 -0.93 105.65 -0.395 ;
      RECT 105.55 0.395 105.65 0.93 ;
      RECT 105.425 -104.945 105.525 -103.985 ;
      RECT 105.05 -100.19 105.4 -100.07 ;
      RECT 105.05 -96.96 105.4 -96.84 ;
      RECT 105.05 -93.73 105.4 -93.61 ;
      RECT 105.05 -90.5 105.4 -90.38 ;
      RECT 105.05 -87.27 105.4 -87.15 ;
      RECT 105.05 -84.04 105.4 -83.92 ;
      RECT 105.05 -80.81 105.4 -80.69 ;
      RECT 105.05 -77.58 105.4 -77.46 ;
      RECT 105.05 -74.35 105.4 -74.23 ;
      RECT 105.05 -71.12 105.4 -71 ;
      RECT 105.05 -67.89 105.4 -67.77 ;
      RECT 105.05 -64.66 105.4 -64.54 ;
      RECT 105.05 -61.43 105.4 -61.31 ;
      RECT 105.05 -58.2 105.4 -58.08 ;
      RECT 105.05 -54.97 105.4 -54.85 ;
      RECT 105.05 -51.74 105.4 -51.62 ;
      RECT 105.05 -48.51 105.4 -48.39 ;
      RECT 105.05 -45.28 105.4 -45.16 ;
      RECT 105.05 -42.05 105.4 -41.93 ;
      RECT 105.05 -38.82 105.4 -38.7 ;
      RECT 105.05 -35.59 105.4 -35.47 ;
      RECT 105.05 -32.36 105.4 -32.24 ;
      RECT 105.05 -29.13 105.4 -29.01 ;
      RECT 105.05 -25.9 105.4 -25.78 ;
      RECT 105.05 -22.67 105.4 -22.55 ;
      RECT 105.05 -19.44 105.4 -19.32 ;
      RECT 105.05 -16.21 105.4 -16.09 ;
      RECT 105.05 -12.98 105.4 -12.86 ;
      RECT 105.05 -9.75 105.4 -9.63 ;
      RECT 105.05 -6.52 105.4 -6.4 ;
      RECT 105.05 -3.29 105.4 -3.17 ;
      RECT 105.05 -0.06 105.4 0.06 ;
      RECT 105.165 -104.945 105.265 -103.985 ;
      RECT 105.165 2.175 105.265 3.135 ;
      RECT 104.875 -112.255 104.975 -111.775 ;
      RECT 104.875 -110.765 104.975 -110.295 ;
      RECT 104.565 -100.19 104.915 -100.07 ;
      RECT 104.565 -96.96 104.915 -96.84 ;
      RECT 104.565 -93.73 104.915 -93.61 ;
      RECT 104.565 -90.5 104.915 -90.38 ;
      RECT 104.565 -87.27 104.915 -87.15 ;
      RECT 104.565 -84.04 104.915 -83.92 ;
      RECT 104.565 -80.81 104.915 -80.69 ;
      RECT 104.565 -77.58 104.915 -77.46 ;
      RECT 104.565 -74.35 104.915 -74.23 ;
      RECT 104.565 -71.12 104.915 -71 ;
      RECT 104.565 -67.89 104.915 -67.77 ;
      RECT 104.565 -64.66 104.915 -64.54 ;
      RECT 104.565 -61.43 104.915 -61.31 ;
      RECT 104.565 -58.2 104.915 -58.08 ;
      RECT 104.565 -54.97 104.915 -54.85 ;
      RECT 104.565 -51.74 104.915 -51.62 ;
      RECT 104.565 -48.51 104.915 -48.39 ;
      RECT 104.565 -45.28 104.915 -45.16 ;
      RECT 104.565 -42.05 104.915 -41.93 ;
      RECT 104.565 -38.82 104.915 -38.7 ;
      RECT 104.565 -35.59 104.915 -35.47 ;
      RECT 104.565 -32.36 104.915 -32.24 ;
      RECT 104.565 -29.13 104.915 -29.01 ;
      RECT 104.565 -25.9 104.915 -25.78 ;
      RECT 104.565 -22.67 104.915 -22.55 ;
      RECT 104.565 -19.44 104.915 -19.32 ;
      RECT 104.565 -16.21 104.915 -16.09 ;
      RECT 104.565 -12.98 104.915 -12.86 ;
      RECT 104.565 -9.75 104.915 -9.63 ;
      RECT 104.565 -6.52 104.915 -6.4 ;
      RECT 104.565 -3.29 104.915 -3.17 ;
      RECT 104.565 -0.06 104.915 0.06 ;
      RECT 104.735 -104.945 104.835 -103.985 ;
      RECT 104.735 2.175 104.835 3.135 ;
      RECT 100.835 -108.655 104.615 -108.535 ;
      RECT 104.475 -104.945 104.575 -103.985 ;
      RECT 104.35 -101.06 104.45 -100.525 ;
      RECT 104.35 -99.735 104.45 -99.2 ;
      RECT 104.35 -97.83 104.45 -97.295 ;
      RECT 104.35 -96.505 104.45 -95.97 ;
      RECT 104.35 -94.6 104.45 -94.065 ;
      RECT 104.35 -93.275 104.45 -92.74 ;
      RECT 104.35 -91.37 104.45 -90.835 ;
      RECT 104.35 -90.045 104.45 -89.51 ;
      RECT 104.35 -88.14 104.45 -87.605 ;
      RECT 104.35 -86.815 104.45 -86.28 ;
      RECT 104.35 -84.91 104.45 -84.375 ;
      RECT 104.35 -83.585 104.45 -83.05 ;
      RECT 104.35 -81.68 104.45 -81.145 ;
      RECT 104.35 -80.355 104.45 -79.82 ;
      RECT 104.35 -78.45 104.45 -77.915 ;
      RECT 104.35 -77.125 104.45 -76.59 ;
      RECT 104.35 -75.22 104.45 -74.685 ;
      RECT 104.35 -73.895 104.45 -73.36 ;
      RECT 104.35 -71.99 104.45 -71.455 ;
      RECT 104.35 -70.665 104.45 -70.13 ;
      RECT 104.35 -68.76 104.45 -68.225 ;
      RECT 104.35 -67.435 104.45 -66.9 ;
      RECT 104.35 -65.53 104.45 -64.995 ;
      RECT 104.35 -64.205 104.45 -63.67 ;
      RECT 104.35 -62.3 104.45 -61.765 ;
      RECT 104.35 -60.975 104.45 -60.44 ;
      RECT 104.35 -59.07 104.45 -58.535 ;
      RECT 104.35 -57.745 104.45 -57.21 ;
      RECT 104.35 -55.84 104.45 -55.305 ;
      RECT 104.35 -54.515 104.45 -53.98 ;
      RECT 104.35 -52.61 104.45 -52.075 ;
      RECT 104.35 -51.285 104.45 -50.75 ;
      RECT 104.35 -49.38 104.45 -48.845 ;
      RECT 104.35 -48.055 104.45 -47.52 ;
      RECT 104.35 -46.15 104.45 -45.615 ;
      RECT 104.35 -44.825 104.45 -44.29 ;
      RECT 104.35 -42.92 104.45 -42.385 ;
      RECT 104.35 -41.595 104.45 -41.06 ;
      RECT 104.35 -39.69 104.45 -39.155 ;
      RECT 104.35 -38.365 104.45 -37.83 ;
      RECT 104.35 -36.46 104.45 -35.925 ;
      RECT 104.35 -35.135 104.45 -34.6 ;
      RECT 104.35 -33.23 104.45 -32.695 ;
      RECT 104.35 -31.905 104.45 -31.37 ;
      RECT 104.35 -30 104.45 -29.465 ;
      RECT 104.35 -28.675 104.45 -28.14 ;
      RECT 104.35 -26.77 104.45 -26.235 ;
      RECT 104.35 -25.445 104.45 -24.91 ;
      RECT 104.35 -23.54 104.45 -23.005 ;
      RECT 104.35 -22.215 104.45 -21.68 ;
      RECT 104.35 -20.31 104.45 -19.775 ;
      RECT 104.35 -18.985 104.45 -18.45 ;
      RECT 104.35 -17.08 104.45 -16.545 ;
      RECT 104.35 -15.755 104.45 -15.22 ;
      RECT 104.35 -13.85 104.45 -13.315 ;
      RECT 104.35 -12.525 104.45 -11.99 ;
      RECT 104.35 -10.62 104.45 -10.085 ;
      RECT 104.35 -9.295 104.45 -8.76 ;
      RECT 104.35 -7.39 104.45 -6.855 ;
      RECT 104.35 -6.065 104.45 -5.53 ;
      RECT 104.35 -4.16 104.45 -3.625 ;
      RECT 104.35 -2.835 104.45 -2.3 ;
      RECT 104.35 -0.93 104.45 -0.395 ;
      RECT 104.35 0.395 104.45 0.93 ;
      RECT 104.285 -110.75 104.405 -110.37 ;
      RECT 104.285 -112.245 104.385 -111.775 ;
      RECT 104.225 -104.945 104.325 -103.985 ;
      RECT 103.85 -100.19 104.2 -100.07 ;
      RECT 103.85 -96.96 104.2 -96.84 ;
      RECT 103.85 -93.73 104.2 -93.61 ;
      RECT 103.85 -90.5 104.2 -90.38 ;
      RECT 103.85 -87.27 104.2 -87.15 ;
      RECT 103.85 -84.04 104.2 -83.92 ;
      RECT 103.85 -80.81 104.2 -80.69 ;
      RECT 103.85 -77.58 104.2 -77.46 ;
      RECT 103.85 -74.35 104.2 -74.23 ;
      RECT 103.85 -71.12 104.2 -71 ;
      RECT 103.85 -67.89 104.2 -67.77 ;
      RECT 103.85 -64.66 104.2 -64.54 ;
      RECT 103.85 -61.43 104.2 -61.31 ;
      RECT 103.85 -58.2 104.2 -58.08 ;
      RECT 103.85 -54.97 104.2 -54.85 ;
      RECT 103.85 -51.74 104.2 -51.62 ;
      RECT 103.85 -48.51 104.2 -48.39 ;
      RECT 103.85 -45.28 104.2 -45.16 ;
      RECT 103.85 -42.05 104.2 -41.93 ;
      RECT 103.85 -38.82 104.2 -38.7 ;
      RECT 103.85 -35.59 104.2 -35.47 ;
      RECT 103.85 -32.36 104.2 -32.24 ;
      RECT 103.85 -29.13 104.2 -29.01 ;
      RECT 103.85 -25.9 104.2 -25.78 ;
      RECT 103.85 -22.67 104.2 -22.55 ;
      RECT 103.85 -19.44 104.2 -19.32 ;
      RECT 103.85 -16.21 104.2 -16.09 ;
      RECT 103.85 -12.98 104.2 -12.86 ;
      RECT 103.85 -9.75 104.2 -9.63 ;
      RECT 103.85 -6.52 104.2 -6.4 ;
      RECT 103.85 -3.29 104.2 -3.17 ;
      RECT 103.85 -0.06 104.2 0.06 ;
      RECT 103.965 -104.945 104.065 -103.985 ;
      RECT 103.965 2.175 104.065 3.135 ;
      RECT 103.695 -109.595 103.83 -109.275 ;
      RECT 103.365 -100.19 103.715 -100.07 ;
      RECT 103.365 -96.96 103.715 -96.84 ;
      RECT 103.365 -93.73 103.715 -93.61 ;
      RECT 103.365 -90.5 103.715 -90.38 ;
      RECT 103.365 -87.27 103.715 -87.15 ;
      RECT 103.365 -84.04 103.715 -83.92 ;
      RECT 103.365 -80.81 103.715 -80.69 ;
      RECT 103.365 -77.58 103.715 -77.46 ;
      RECT 103.365 -74.35 103.715 -74.23 ;
      RECT 103.365 -71.12 103.715 -71 ;
      RECT 103.365 -67.89 103.715 -67.77 ;
      RECT 103.365 -64.66 103.715 -64.54 ;
      RECT 103.365 -61.43 103.715 -61.31 ;
      RECT 103.365 -58.2 103.715 -58.08 ;
      RECT 103.365 -54.97 103.715 -54.85 ;
      RECT 103.365 -51.74 103.715 -51.62 ;
      RECT 103.365 -48.51 103.715 -48.39 ;
      RECT 103.365 -45.28 103.715 -45.16 ;
      RECT 103.365 -42.05 103.715 -41.93 ;
      RECT 103.365 -38.82 103.715 -38.7 ;
      RECT 103.365 -35.59 103.715 -35.47 ;
      RECT 103.365 -32.36 103.715 -32.24 ;
      RECT 103.365 -29.13 103.715 -29.01 ;
      RECT 103.365 -25.9 103.715 -25.78 ;
      RECT 103.365 -22.67 103.715 -22.55 ;
      RECT 103.365 -19.44 103.715 -19.32 ;
      RECT 103.365 -16.21 103.715 -16.09 ;
      RECT 103.365 -12.98 103.715 -12.86 ;
      RECT 103.365 -9.75 103.715 -9.63 ;
      RECT 103.365 -6.52 103.715 -6.4 ;
      RECT 103.365 -3.29 103.715 -3.17 ;
      RECT 103.365 -0.06 103.715 0.06 ;
      RECT 103.535 -104.945 103.635 -103.985 ;
      RECT 103.535 2.175 103.635 3.135 ;
      RECT 103.36 -109.595 103.505 -109.275 ;
      RECT 103.275 -104.945 103.375 -103.985 ;
      RECT 103.15 -101.06 103.25 -100.525 ;
      RECT 103.15 -99.735 103.25 -99.2 ;
      RECT 103.15 -97.83 103.25 -97.295 ;
      RECT 103.15 -96.505 103.25 -95.97 ;
      RECT 103.15 -94.6 103.25 -94.065 ;
      RECT 103.15 -93.275 103.25 -92.74 ;
      RECT 103.15 -91.37 103.25 -90.835 ;
      RECT 103.15 -90.045 103.25 -89.51 ;
      RECT 103.15 -88.14 103.25 -87.605 ;
      RECT 103.15 -86.815 103.25 -86.28 ;
      RECT 103.15 -84.91 103.25 -84.375 ;
      RECT 103.15 -83.585 103.25 -83.05 ;
      RECT 103.15 -81.68 103.25 -81.145 ;
      RECT 103.15 -80.355 103.25 -79.82 ;
      RECT 103.15 -78.45 103.25 -77.915 ;
      RECT 103.15 -77.125 103.25 -76.59 ;
      RECT 103.15 -75.22 103.25 -74.685 ;
      RECT 103.15 -73.895 103.25 -73.36 ;
      RECT 103.15 -71.99 103.25 -71.455 ;
      RECT 103.15 -70.665 103.25 -70.13 ;
      RECT 103.15 -68.76 103.25 -68.225 ;
      RECT 103.15 -67.435 103.25 -66.9 ;
      RECT 103.15 -65.53 103.25 -64.995 ;
      RECT 103.15 -64.205 103.25 -63.67 ;
      RECT 103.15 -62.3 103.25 -61.765 ;
      RECT 103.15 -60.975 103.25 -60.44 ;
      RECT 103.15 -59.07 103.25 -58.535 ;
      RECT 103.15 -57.745 103.25 -57.21 ;
      RECT 103.15 -55.84 103.25 -55.305 ;
      RECT 103.15 -54.515 103.25 -53.98 ;
      RECT 103.15 -52.61 103.25 -52.075 ;
      RECT 103.15 -51.285 103.25 -50.75 ;
      RECT 103.15 -49.38 103.25 -48.845 ;
      RECT 103.15 -48.055 103.25 -47.52 ;
      RECT 103.15 -46.15 103.25 -45.615 ;
      RECT 103.15 -44.825 103.25 -44.29 ;
      RECT 103.15 -42.92 103.25 -42.385 ;
      RECT 103.15 -41.595 103.25 -41.06 ;
      RECT 103.15 -39.69 103.25 -39.155 ;
      RECT 103.15 -38.365 103.25 -37.83 ;
      RECT 103.15 -36.46 103.25 -35.925 ;
      RECT 103.15 -35.135 103.25 -34.6 ;
      RECT 103.15 -33.23 103.25 -32.695 ;
      RECT 103.15 -31.905 103.25 -31.37 ;
      RECT 103.15 -30 103.25 -29.465 ;
      RECT 103.15 -28.675 103.25 -28.14 ;
      RECT 103.15 -26.77 103.25 -26.235 ;
      RECT 103.15 -25.445 103.25 -24.91 ;
      RECT 103.15 -23.54 103.25 -23.005 ;
      RECT 103.15 -22.215 103.25 -21.68 ;
      RECT 103.15 -20.31 103.25 -19.775 ;
      RECT 103.15 -18.985 103.25 -18.45 ;
      RECT 103.15 -17.08 103.25 -16.545 ;
      RECT 103.15 -15.755 103.25 -15.22 ;
      RECT 103.15 -13.85 103.25 -13.315 ;
      RECT 103.15 -12.525 103.25 -11.99 ;
      RECT 103.15 -10.62 103.25 -10.085 ;
      RECT 103.15 -9.295 103.25 -8.76 ;
      RECT 103.15 -7.39 103.25 -6.855 ;
      RECT 103.15 -6.065 103.25 -5.53 ;
      RECT 103.15 -4.16 103.25 -3.625 ;
      RECT 103.15 -2.835 103.25 -2.3 ;
      RECT 103.15 -0.93 103.25 -0.395 ;
      RECT 103.15 0.395 103.25 0.93 ;
      RECT 103.025 -108.175 103.125 -107.215 ;
      RECT 102.65 -100.19 103 -100.07 ;
      RECT 102.65 -96.96 103 -96.84 ;
      RECT 102.65 -93.73 103 -93.61 ;
      RECT 102.65 -90.5 103 -90.38 ;
      RECT 102.65 -87.27 103 -87.15 ;
      RECT 102.65 -84.04 103 -83.92 ;
      RECT 102.65 -80.81 103 -80.69 ;
      RECT 102.65 -77.58 103 -77.46 ;
      RECT 102.65 -74.35 103 -74.23 ;
      RECT 102.65 -71.12 103 -71 ;
      RECT 102.65 -67.89 103 -67.77 ;
      RECT 102.65 -64.66 103 -64.54 ;
      RECT 102.65 -61.43 103 -61.31 ;
      RECT 102.65 -58.2 103 -58.08 ;
      RECT 102.65 -54.97 103 -54.85 ;
      RECT 102.65 -51.74 103 -51.62 ;
      RECT 102.65 -48.51 103 -48.39 ;
      RECT 102.65 -45.28 103 -45.16 ;
      RECT 102.65 -42.05 103 -41.93 ;
      RECT 102.65 -38.82 103 -38.7 ;
      RECT 102.65 -35.59 103 -35.47 ;
      RECT 102.65 -32.36 103 -32.24 ;
      RECT 102.65 -29.13 103 -29.01 ;
      RECT 102.65 -25.9 103 -25.78 ;
      RECT 102.65 -22.67 103 -22.55 ;
      RECT 102.65 -19.44 103 -19.32 ;
      RECT 102.65 -16.21 103 -16.09 ;
      RECT 102.65 -12.98 103 -12.86 ;
      RECT 102.65 -9.75 103 -9.63 ;
      RECT 102.65 -6.52 103 -6.4 ;
      RECT 102.65 -3.29 103 -3.17 ;
      RECT 102.65 -0.06 103 0.06 ;
      RECT 102.855 -112.255 102.955 -111.775 ;
      RECT 102.855 -110.765 102.955 -110.295 ;
      RECT 102.765 -108.175 102.865 -107.215 ;
      RECT 102.765 2.175 102.865 3.135 ;
      RECT 102.165 -100.19 102.515 -100.07 ;
      RECT 102.165 -96.96 102.515 -96.84 ;
      RECT 102.165 -93.73 102.515 -93.61 ;
      RECT 102.165 -90.5 102.515 -90.38 ;
      RECT 102.165 -87.27 102.515 -87.15 ;
      RECT 102.165 -84.04 102.515 -83.92 ;
      RECT 102.165 -80.81 102.515 -80.69 ;
      RECT 102.165 -77.58 102.515 -77.46 ;
      RECT 102.165 -74.35 102.515 -74.23 ;
      RECT 102.165 -71.12 102.515 -71 ;
      RECT 102.165 -67.89 102.515 -67.77 ;
      RECT 102.165 -64.66 102.515 -64.54 ;
      RECT 102.165 -61.43 102.515 -61.31 ;
      RECT 102.165 -58.2 102.515 -58.08 ;
      RECT 102.165 -54.97 102.515 -54.85 ;
      RECT 102.165 -51.74 102.515 -51.62 ;
      RECT 102.165 -48.51 102.515 -48.39 ;
      RECT 102.165 -45.28 102.515 -45.16 ;
      RECT 102.165 -42.05 102.515 -41.93 ;
      RECT 102.165 -38.82 102.515 -38.7 ;
      RECT 102.165 -35.59 102.515 -35.47 ;
      RECT 102.165 -32.36 102.515 -32.24 ;
      RECT 102.165 -29.13 102.515 -29.01 ;
      RECT 102.165 -25.9 102.515 -25.78 ;
      RECT 102.165 -22.67 102.515 -22.55 ;
      RECT 102.165 -19.44 102.515 -19.32 ;
      RECT 102.165 -16.21 102.515 -16.09 ;
      RECT 102.165 -12.98 102.515 -12.86 ;
      RECT 102.165 -9.75 102.515 -9.63 ;
      RECT 102.165 -6.52 102.515 -6.4 ;
      RECT 102.165 -3.29 102.515 -3.17 ;
      RECT 102.165 -0.06 102.515 0.06 ;
      RECT 102.335 -108.175 102.435 -107.215 ;
      RECT 102.335 2.175 102.435 3.135 ;
      RECT 102.23 -110.765 102.4 -110.385 ;
      RECT 102.265 -112.245 102.365 -111.775 ;
      RECT 102.075 -108.175 102.175 -107.215 ;
      RECT 101.95 -101.06 102.05 -100.525 ;
      RECT 101.95 -99.735 102.05 -99.2 ;
      RECT 101.95 -97.83 102.05 -97.295 ;
      RECT 101.95 -96.505 102.05 -95.97 ;
      RECT 101.95 -94.6 102.05 -94.065 ;
      RECT 101.95 -93.275 102.05 -92.74 ;
      RECT 101.95 -91.37 102.05 -90.835 ;
      RECT 101.95 -90.045 102.05 -89.51 ;
      RECT 101.95 -88.14 102.05 -87.605 ;
      RECT 101.95 -86.815 102.05 -86.28 ;
      RECT 101.95 -84.91 102.05 -84.375 ;
      RECT 101.95 -83.585 102.05 -83.05 ;
      RECT 101.95 -81.68 102.05 -81.145 ;
      RECT 101.95 -80.355 102.05 -79.82 ;
      RECT 101.95 -78.45 102.05 -77.915 ;
      RECT 101.95 -77.125 102.05 -76.59 ;
      RECT 101.95 -75.22 102.05 -74.685 ;
      RECT 101.95 -73.895 102.05 -73.36 ;
      RECT 101.95 -71.99 102.05 -71.455 ;
      RECT 101.95 -70.665 102.05 -70.13 ;
      RECT 101.95 -68.76 102.05 -68.225 ;
      RECT 101.95 -67.435 102.05 -66.9 ;
      RECT 101.95 -65.53 102.05 -64.995 ;
      RECT 101.95 -64.205 102.05 -63.67 ;
      RECT 101.95 -62.3 102.05 -61.765 ;
      RECT 101.95 -60.975 102.05 -60.44 ;
      RECT 101.95 -59.07 102.05 -58.535 ;
      RECT 101.95 -57.745 102.05 -57.21 ;
      RECT 101.95 -55.84 102.05 -55.305 ;
      RECT 101.95 -54.515 102.05 -53.98 ;
      RECT 101.95 -52.61 102.05 -52.075 ;
      RECT 101.95 -51.285 102.05 -50.75 ;
      RECT 101.95 -49.38 102.05 -48.845 ;
      RECT 101.95 -48.055 102.05 -47.52 ;
      RECT 101.95 -46.15 102.05 -45.615 ;
      RECT 101.95 -44.825 102.05 -44.29 ;
      RECT 101.95 -42.92 102.05 -42.385 ;
      RECT 101.95 -41.595 102.05 -41.06 ;
      RECT 101.95 -39.69 102.05 -39.155 ;
      RECT 101.95 -38.365 102.05 -37.83 ;
      RECT 101.95 -36.46 102.05 -35.925 ;
      RECT 101.95 -35.135 102.05 -34.6 ;
      RECT 101.95 -33.23 102.05 -32.695 ;
      RECT 101.95 -31.905 102.05 -31.37 ;
      RECT 101.95 -30 102.05 -29.465 ;
      RECT 101.95 -28.675 102.05 -28.14 ;
      RECT 101.95 -26.77 102.05 -26.235 ;
      RECT 101.95 -25.445 102.05 -24.91 ;
      RECT 101.95 -23.54 102.05 -23.005 ;
      RECT 101.95 -22.215 102.05 -21.68 ;
      RECT 101.95 -20.31 102.05 -19.775 ;
      RECT 101.95 -18.985 102.05 -18.45 ;
      RECT 101.95 -17.08 102.05 -16.545 ;
      RECT 101.95 -15.755 102.05 -15.22 ;
      RECT 101.95 -13.85 102.05 -13.315 ;
      RECT 101.95 -12.525 102.05 -11.99 ;
      RECT 101.95 -10.62 102.05 -10.085 ;
      RECT 101.95 -9.295 102.05 -8.76 ;
      RECT 101.95 -7.39 102.05 -6.855 ;
      RECT 101.95 -6.065 102.05 -5.53 ;
      RECT 101.95 -4.16 102.05 -3.625 ;
      RECT 101.95 -2.835 102.05 -2.3 ;
      RECT 101.95 -0.93 102.05 -0.395 ;
      RECT 101.95 0.395 102.05 0.93 ;
      RECT 101.825 -108.175 101.925 -107.215 ;
      RECT 101.45 -100.19 101.8 -100.07 ;
      RECT 101.45 -96.96 101.8 -96.84 ;
      RECT 101.45 -93.73 101.8 -93.61 ;
      RECT 101.45 -90.5 101.8 -90.38 ;
      RECT 101.45 -87.27 101.8 -87.15 ;
      RECT 101.45 -84.04 101.8 -83.92 ;
      RECT 101.45 -80.81 101.8 -80.69 ;
      RECT 101.45 -77.58 101.8 -77.46 ;
      RECT 101.45 -74.35 101.8 -74.23 ;
      RECT 101.45 -71.12 101.8 -71 ;
      RECT 101.45 -67.89 101.8 -67.77 ;
      RECT 101.45 -64.66 101.8 -64.54 ;
      RECT 101.45 -61.43 101.8 -61.31 ;
      RECT 101.45 -58.2 101.8 -58.08 ;
      RECT 101.45 -54.97 101.8 -54.85 ;
      RECT 101.45 -51.74 101.8 -51.62 ;
      RECT 101.45 -48.51 101.8 -48.39 ;
      RECT 101.45 -45.28 101.8 -45.16 ;
      RECT 101.45 -42.05 101.8 -41.93 ;
      RECT 101.45 -38.82 101.8 -38.7 ;
      RECT 101.45 -35.59 101.8 -35.47 ;
      RECT 101.45 -32.36 101.8 -32.24 ;
      RECT 101.45 -29.13 101.8 -29.01 ;
      RECT 101.45 -25.9 101.8 -25.78 ;
      RECT 101.45 -22.67 101.8 -22.55 ;
      RECT 101.45 -19.44 101.8 -19.32 ;
      RECT 101.45 -16.21 101.8 -16.09 ;
      RECT 101.45 -12.98 101.8 -12.86 ;
      RECT 101.45 -9.75 101.8 -9.63 ;
      RECT 101.45 -6.52 101.8 -6.4 ;
      RECT 101.45 -3.29 101.8 -3.17 ;
      RECT 101.45 -0.06 101.8 0.06 ;
      RECT 101.565 -108.175 101.665 -107.215 ;
      RECT 101.565 2.175 101.665 3.135 ;
      RECT 101.465 -113.555 101.565 -113.085 ;
      RECT 100.965 -100.19 101.315 -100.07 ;
      RECT 100.965 -96.96 101.315 -96.84 ;
      RECT 100.965 -93.73 101.315 -93.61 ;
      RECT 100.965 -90.5 101.315 -90.38 ;
      RECT 100.965 -87.27 101.315 -87.15 ;
      RECT 100.965 -84.04 101.315 -83.92 ;
      RECT 100.965 -80.81 101.315 -80.69 ;
      RECT 100.965 -77.58 101.315 -77.46 ;
      RECT 100.965 -74.35 101.315 -74.23 ;
      RECT 100.965 -71.12 101.315 -71 ;
      RECT 100.965 -67.89 101.315 -67.77 ;
      RECT 100.965 -64.66 101.315 -64.54 ;
      RECT 100.965 -61.43 101.315 -61.31 ;
      RECT 100.965 -58.2 101.315 -58.08 ;
      RECT 100.965 -54.97 101.315 -54.85 ;
      RECT 100.965 -51.74 101.315 -51.62 ;
      RECT 100.965 -48.51 101.315 -48.39 ;
      RECT 100.965 -45.28 101.315 -45.16 ;
      RECT 100.965 -42.05 101.315 -41.93 ;
      RECT 100.965 -38.82 101.315 -38.7 ;
      RECT 100.965 -35.59 101.315 -35.47 ;
      RECT 100.965 -32.36 101.315 -32.24 ;
      RECT 100.965 -29.13 101.315 -29.01 ;
      RECT 100.965 -25.9 101.315 -25.78 ;
      RECT 100.965 -22.67 101.315 -22.55 ;
      RECT 100.965 -19.44 101.315 -19.32 ;
      RECT 100.965 -16.21 101.315 -16.09 ;
      RECT 100.965 -12.98 101.315 -12.86 ;
      RECT 100.965 -9.75 101.315 -9.63 ;
      RECT 100.965 -6.52 101.315 -6.4 ;
      RECT 100.965 -3.29 101.315 -3.17 ;
      RECT 100.965 -0.06 101.315 0.06 ;
      RECT 101.1 -110.735 101.25 -110.445 ;
      RECT 101.135 -108.175 101.235 -107.215 ;
      RECT 101.135 2.175 101.235 3.135 ;
      RECT 101.115 -112.19 101.215 -111.65 ;
      RECT 100.875 -113.555 100.975 -113.085 ;
      RECT 100.875 -108.175 100.975 -107.215 ;
      RECT 100.75 -101.06 100.85 -100.525 ;
      RECT 100.75 -99.735 100.85 -99.2 ;
      RECT 100.75 -97.83 100.85 -97.295 ;
      RECT 100.75 -96.505 100.85 -95.97 ;
      RECT 100.75 -94.6 100.85 -94.065 ;
      RECT 100.75 -93.275 100.85 -92.74 ;
      RECT 100.75 -91.37 100.85 -90.835 ;
      RECT 100.75 -90.045 100.85 -89.51 ;
      RECT 100.75 -88.14 100.85 -87.605 ;
      RECT 100.75 -86.815 100.85 -86.28 ;
      RECT 100.75 -84.91 100.85 -84.375 ;
      RECT 100.75 -83.585 100.85 -83.05 ;
      RECT 100.75 -81.68 100.85 -81.145 ;
      RECT 100.75 -80.355 100.85 -79.82 ;
      RECT 100.75 -78.45 100.85 -77.915 ;
      RECT 100.75 -77.125 100.85 -76.59 ;
      RECT 100.75 -75.22 100.85 -74.685 ;
      RECT 100.75 -73.895 100.85 -73.36 ;
      RECT 100.75 -71.99 100.85 -71.455 ;
      RECT 100.75 -70.665 100.85 -70.13 ;
      RECT 100.75 -68.76 100.85 -68.225 ;
      RECT 100.75 -67.435 100.85 -66.9 ;
      RECT 100.75 -65.53 100.85 -64.995 ;
      RECT 100.75 -64.205 100.85 -63.67 ;
      RECT 100.75 -62.3 100.85 -61.765 ;
      RECT 100.75 -60.975 100.85 -60.44 ;
      RECT 100.75 -59.07 100.85 -58.535 ;
      RECT 100.75 -57.745 100.85 -57.21 ;
      RECT 100.75 -55.84 100.85 -55.305 ;
      RECT 100.75 -54.515 100.85 -53.98 ;
      RECT 100.75 -52.61 100.85 -52.075 ;
      RECT 100.75 -51.285 100.85 -50.75 ;
      RECT 100.75 -49.38 100.85 -48.845 ;
      RECT 100.75 -48.055 100.85 -47.52 ;
      RECT 100.75 -46.15 100.85 -45.615 ;
      RECT 100.75 -44.825 100.85 -44.29 ;
      RECT 100.75 -42.92 100.85 -42.385 ;
      RECT 100.75 -41.595 100.85 -41.06 ;
      RECT 100.75 -39.69 100.85 -39.155 ;
      RECT 100.75 -38.365 100.85 -37.83 ;
      RECT 100.75 -36.46 100.85 -35.925 ;
      RECT 100.75 -35.135 100.85 -34.6 ;
      RECT 100.75 -33.23 100.85 -32.695 ;
      RECT 100.75 -31.905 100.85 -31.37 ;
      RECT 100.75 -30 100.85 -29.465 ;
      RECT 100.75 -28.675 100.85 -28.14 ;
      RECT 100.75 -26.77 100.85 -26.235 ;
      RECT 100.75 -25.445 100.85 -24.91 ;
      RECT 100.75 -23.54 100.85 -23.005 ;
      RECT 100.75 -22.215 100.85 -21.68 ;
      RECT 100.75 -20.31 100.85 -19.775 ;
      RECT 100.75 -18.985 100.85 -18.45 ;
      RECT 100.75 -17.08 100.85 -16.545 ;
      RECT 100.75 -15.755 100.85 -15.22 ;
      RECT 100.75 -13.85 100.85 -13.315 ;
      RECT 100.75 -12.525 100.85 -11.99 ;
      RECT 100.75 -10.62 100.85 -10.085 ;
      RECT 100.75 -9.295 100.85 -8.76 ;
      RECT 100.75 -7.39 100.85 -6.855 ;
      RECT 100.75 -6.065 100.85 -5.53 ;
      RECT 100.75 -4.16 100.85 -3.625 ;
      RECT 100.75 -2.835 100.85 -2.3 ;
      RECT 100.75 -0.93 100.85 -0.395 ;
      RECT 100.75 0.395 100.85 0.93 ;
      RECT 100.625 -104.945 100.725 -103.985 ;
      RECT 100.25 -100.19 100.6 -100.07 ;
      RECT 100.25 -96.96 100.6 -96.84 ;
      RECT 100.25 -93.73 100.6 -93.61 ;
      RECT 100.25 -90.5 100.6 -90.38 ;
      RECT 100.25 -87.27 100.6 -87.15 ;
      RECT 100.25 -84.04 100.6 -83.92 ;
      RECT 100.25 -80.81 100.6 -80.69 ;
      RECT 100.25 -77.58 100.6 -77.46 ;
      RECT 100.25 -74.35 100.6 -74.23 ;
      RECT 100.25 -71.12 100.6 -71 ;
      RECT 100.25 -67.89 100.6 -67.77 ;
      RECT 100.25 -64.66 100.6 -64.54 ;
      RECT 100.25 -61.43 100.6 -61.31 ;
      RECT 100.25 -58.2 100.6 -58.08 ;
      RECT 100.25 -54.97 100.6 -54.85 ;
      RECT 100.25 -51.74 100.6 -51.62 ;
      RECT 100.25 -48.51 100.6 -48.39 ;
      RECT 100.25 -45.28 100.6 -45.16 ;
      RECT 100.25 -42.05 100.6 -41.93 ;
      RECT 100.25 -38.82 100.6 -38.7 ;
      RECT 100.25 -35.59 100.6 -35.47 ;
      RECT 100.25 -32.36 100.6 -32.24 ;
      RECT 100.25 -29.13 100.6 -29.01 ;
      RECT 100.25 -25.9 100.6 -25.78 ;
      RECT 100.25 -22.67 100.6 -22.55 ;
      RECT 100.25 -19.44 100.6 -19.32 ;
      RECT 100.25 -16.21 100.6 -16.09 ;
      RECT 100.25 -12.98 100.6 -12.86 ;
      RECT 100.25 -9.75 100.6 -9.63 ;
      RECT 100.25 -6.52 100.6 -6.4 ;
      RECT 100.25 -3.29 100.6 -3.17 ;
      RECT 100.25 -0.06 100.6 0.06 ;
      RECT 100.365 -104.945 100.465 -103.985 ;
      RECT 100.365 2.175 100.465 3.135 ;
      RECT 100.075 -112.255 100.175 -111.775 ;
      RECT 100.075 -110.765 100.175 -110.295 ;
      RECT 99.765 -100.19 100.115 -100.07 ;
      RECT 99.765 -96.96 100.115 -96.84 ;
      RECT 99.765 -93.73 100.115 -93.61 ;
      RECT 99.765 -90.5 100.115 -90.38 ;
      RECT 99.765 -87.27 100.115 -87.15 ;
      RECT 99.765 -84.04 100.115 -83.92 ;
      RECT 99.765 -80.81 100.115 -80.69 ;
      RECT 99.765 -77.58 100.115 -77.46 ;
      RECT 99.765 -74.35 100.115 -74.23 ;
      RECT 99.765 -71.12 100.115 -71 ;
      RECT 99.765 -67.89 100.115 -67.77 ;
      RECT 99.765 -64.66 100.115 -64.54 ;
      RECT 99.765 -61.43 100.115 -61.31 ;
      RECT 99.765 -58.2 100.115 -58.08 ;
      RECT 99.765 -54.97 100.115 -54.85 ;
      RECT 99.765 -51.74 100.115 -51.62 ;
      RECT 99.765 -48.51 100.115 -48.39 ;
      RECT 99.765 -45.28 100.115 -45.16 ;
      RECT 99.765 -42.05 100.115 -41.93 ;
      RECT 99.765 -38.82 100.115 -38.7 ;
      RECT 99.765 -35.59 100.115 -35.47 ;
      RECT 99.765 -32.36 100.115 -32.24 ;
      RECT 99.765 -29.13 100.115 -29.01 ;
      RECT 99.765 -25.9 100.115 -25.78 ;
      RECT 99.765 -22.67 100.115 -22.55 ;
      RECT 99.765 -19.44 100.115 -19.32 ;
      RECT 99.765 -16.21 100.115 -16.09 ;
      RECT 99.765 -12.98 100.115 -12.86 ;
      RECT 99.765 -9.75 100.115 -9.63 ;
      RECT 99.765 -6.52 100.115 -6.4 ;
      RECT 99.765 -3.29 100.115 -3.17 ;
      RECT 99.765 -0.06 100.115 0.06 ;
      RECT 99.935 -104.945 100.035 -103.985 ;
      RECT 99.935 2.175 100.035 3.135 ;
      RECT 96.035 -108.655 99.815 -108.535 ;
      RECT 99.675 -104.945 99.775 -103.985 ;
      RECT 99.55 -101.06 99.65 -100.525 ;
      RECT 99.55 -99.735 99.65 -99.2 ;
      RECT 99.55 -97.83 99.65 -97.295 ;
      RECT 99.55 -96.505 99.65 -95.97 ;
      RECT 99.55 -94.6 99.65 -94.065 ;
      RECT 99.55 -93.275 99.65 -92.74 ;
      RECT 99.55 -91.37 99.65 -90.835 ;
      RECT 99.55 -90.045 99.65 -89.51 ;
      RECT 99.55 -88.14 99.65 -87.605 ;
      RECT 99.55 -86.815 99.65 -86.28 ;
      RECT 99.55 -84.91 99.65 -84.375 ;
      RECT 99.55 -83.585 99.65 -83.05 ;
      RECT 99.55 -81.68 99.65 -81.145 ;
      RECT 99.55 -80.355 99.65 -79.82 ;
      RECT 99.55 -78.45 99.65 -77.915 ;
      RECT 99.55 -77.125 99.65 -76.59 ;
      RECT 99.55 -75.22 99.65 -74.685 ;
      RECT 99.55 -73.895 99.65 -73.36 ;
      RECT 99.55 -71.99 99.65 -71.455 ;
      RECT 99.55 -70.665 99.65 -70.13 ;
      RECT 99.55 -68.76 99.65 -68.225 ;
      RECT 99.55 -67.435 99.65 -66.9 ;
      RECT 99.55 -65.53 99.65 -64.995 ;
      RECT 99.55 -64.205 99.65 -63.67 ;
      RECT 99.55 -62.3 99.65 -61.765 ;
      RECT 99.55 -60.975 99.65 -60.44 ;
      RECT 99.55 -59.07 99.65 -58.535 ;
      RECT 99.55 -57.745 99.65 -57.21 ;
      RECT 99.55 -55.84 99.65 -55.305 ;
      RECT 99.55 -54.515 99.65 -53.98 ;
      RECT 99.55 -52.61 99.65 -52.075 ;
      RECT 99.55 -51.285 99.65 -50.75 ;
      RECT 99.55 -49.38 99.65 -48.845 ;
      RECT 99.55 -48.055 99.65 -47.52 ;
      RECT 99.55 -46.15 99.65 -45.615 ;
      RECT 99.55 -44.825 99.65 -44.29 ;
      RECT 99.55 -42.92 99.65 -42.385 ;
      RECT 99.55 -41.595 99.65 -41.06 ;
      RECT 99.55 -39.69 99.65 -39.155 ;
      RECT 99.55 -38.365 99.65 -37.83 ;
      RECT 99.55 -36.46 99.65 -35.925 ;
      RECT 99.55 -35.135 99.65 -34.6 ;
      RECT 99.55 -33.23 99.65 -32.695 ;
      RECT 99.55 -31.905 99.65 -31.37 ;
      RECT 99.55 -30 99.65 -29.465 ;
      RECT 99.55 -28.675 99.65 -28.14 ;
      RECT 99.55 -26.77 99.65 -26.235 ;
      RECT 99.55 -25.445 99.65 -24.91 ;
      RECT 99.55 -23.54 99.65 -23.005 ;
      RECT 99.55 -22.215 99.65 -21.68 ;
      RECT 99.55 -20.31 99.65 -19.775 ;
      RECT 99.55 -18.985 99.65 -18.45 ;
      RECT 99.55 -17.08 99.65 -16.545 ;
      RECT 99.55 -15.755 99.65 -15.22 ;
      RECT 99.55 -13.85 99.65 -13.315 ;
      RECT 99.55 -12.525 99.65 -11.99 ;
      RECT 99.55 -10.62 99.65 -10.085 ;
      RECT 99.55 -9.295 99.65 -8.76 ;
      RECT 99.55 -7.39 99.65 -6.855 ;
      RECT 99.55 -6.065 99.65 -5.53 ;
      RECT 99.55 -4.16 99.65 -3.625 ;
      RECT 99.55 -2.835 99.65 -2.3 ;
      RECT 99.55 -0.93 99.65 -0.395 ;
      RECT 99.55 0.395 99.65 0.93 ;
      RECT 99.485 -110.75 99.605 -110.37 ;
      RECT 99.485 -112.245 99.585 -111.775 ;
      RECT 99.425 -104.945 99.525 -103.985 ;
      RECT 99.05 -100.19 99.4 -100.07 ;
      RECT 99.05 -96.96 99.4 -96.84 ;
      RECT 99.05 -93.73 99.4 -93.61 ;
      RECT 99.05 -90.5 99.4 -90.38 ;
      RECT 99.05 -87.27 99.4 -87.15 ;
      RECT 99.05 -84.04 99.4 -83.92 ;
      RECT 99.05 -80.81 99.4 -80.69 ;
      RECT 99.05 -77.58 99.4 -77.46 ;
      RECT 99.05 -74.35 99.4 -74.23 ;
      RECT 99.05 -71.12 99.4 -71 ;
      RECT 99.05 -67.89 99.4 -67.77 ;
      RECT 99.05 -64.66 99.4 -64.54 ;
      RECT 99.05 -61.43 99.4 -61.31 ;
      RECT 99.05 -58.2 99.4 -58.08 ;
      RECT 99.05 -54.97 99.4 -54.85 ;
      RECT 99.05 -51.74 99.4 -51.62 ;
      RECT 99.05 -48.51 99.4 -48.39 ;
      RECT 99.05 -45.28 99.4 -45.16 ;
      RECT 99.05 -42.05 99.4 -41.93 ;
      RECT 99.05 -38.82 99.4 -38.7 ;
      RECT 99.05 -35.59 99.4 -35.47 ;
      RECT 99.05 -32.36 99.4 -32.24 ;
      RECT 99.05 -29.13 99.4 -29.01 ;
      RECT 99.05 -25.9 99.4 -25.78 ;
      RECT 99.05 -22.67 99.4 -22.55 ;
      RECT 99.05 -19.44 99.4 -19.32 ;
      RECT 99.05 -16.21 99.4 -16.09 ;
      RECT 99.05 -12.98 99.4 -12.86 ;
      RECT 99.05 -9.75 99.4 -9.63 ;
      RECT 99.05 -6.52 99.4 -6.4 ;
      RECT 99.05 -3.29 99.4 -3.17 ;
      RECT 99.05 -0.06 99.4 0.06 ;
      RECT 99.165 -104.945 99.265 -103.985 ;
      RECT 99.165 2.175 99.265 3.135 ;
      RECT 98.895 -109.595 99.03 -109.275 ;
      RECT 98.565 -100.19 98.915 -100.07 ;
      RECT 98.565 -96.96 98.915 -96.84 ;
      RECT 98.565 -93.73 98.915 -93.61 ;
      RECT 98.565 -90.5 98.915 -90.38 ;
      RECT 98.565 -87.27 98.915 -87.15 ;
      RECT 98.565 -84.04 98.915 -83.92 ;
      RECT 98.565 -80.81 98.915 -80.69 ;
      RECT 98.565 -77.58 98.915 -77.46 ;
      RECT 98.565 -74.35 98.915 -74.23 ;
      RECT 98.565 -71.12 98.915 -71 ;
      RECT 98.565 -67.89 98.915 -67.77 ;
      RECT 98.565 -64.66 98.915 -64.54 ;
      RECT 98.565 -61.43 98.915 -61.31 ;
      RECT 98.565 -58.2 98.915 -58.08 ;
      RECT 98.565 -54.97 98.915 -54.85 ;
      RECT 98.565 -51.74 98.915 -51.62 ;
      RECT 98.565 -48.51 98.915 -48.39 ;
      RECT 98.565 -45.28 98.915 -45.16 ;
      RECT 98.565 -42.05 98.915 -41.93 ;
      RECT 98.565 -38.82 98.915 -38.7 ;
      RECT 98.565 -35.59 98.915 -35.47 ;
      RECT 98.565 -32.36 98.915 -32.24 ;
      RECT 98.565 -29.13 98.915 -29.01 ;
      RECT 98.565 -25.9 98.915 -25.78 ;
      RECT 98.565 -22.67 98.915 -22.55 ;
      RECT 98.565 -19.44 98.915 -19.32 ;
      RECT 98.565 -16.21 98.915 -16.09 ;
      RECT 98.565 -12.98 98.915 -12.86 ;
      RECT 98.565 -9.75 98.915 -9.63 ;
      RECT 98.565 -6.52 98.915 -6.4 ;
      RECT 98.565 -3.29 98.915 -3.17 ;
      RECT 98.565 -0.06 98.915 0.06 ;
      RECT 98.735 -104.945 98.835 -103.985 ;
      RECT 98.735 2.175 98.835 3.135 ;
      RECT 98.56 -109.595 98.705 -109.275 ;
      RECT 98.475 -104.945 98.575 -103.985 ;
      RECT 98.35 -101.06 98.45 -100.525 ;
      RECT 98.35 -99.735 98.45 -99.2 ;
      RECT 98.35 -97.83 98.45 -97.295 ;
      RECT 98.35 -96.505 98.45 -95.97 ;
      RECT 98.35 -94.6 98.45 -94.065 ;
      RECT 98.35 -93.275 98.45 -92.74 ;
      RECT 98.35 -91.37 98.45 -90.835 ;
      RECT 98.35 -90.045 98.45 -89.51 ;
      RECT 98.35 -88.14 98.45 -87.605 ;
      RECT 98.35 -86.815 98.45 -86.28 ;
      RECT 98.35 -84.91 98.45 -84.375 ;
      RECT 98.35 -83.585 98.45 -83.05 ;
      RECT 98.35 -81.68 98.45 -81.145 ;
      RECT 98.35 -80.355 98.45 -79.82 ;
      RECT 98.35 -78.45 98.45 -77.915 ;
      RECT 98.35 -77.125 98.45 -76.59 ;
      RECT 98.35 -75.22 98.45 -74.685 ;
      RECT 98.35 -73.895 98.45 -73.36 ;
      RECT 98.35 -71.99 98.45 -71.455 ;
      RECT 98.35 -70.665 98.45 -70.13 ;
      RECT 98.35 -68.76 98.45 -68.225 ;
      RECT 98.35 -67.435 98.45 -66.9 ;
      RECT 98.35 -65.53 98.45 -64.995 ;
      RECT 98.35 -64.205 98.45 -63.67 ;
      RECT 98.35 -62.3 98.45 -61.765 ;
      RECT 98.35 -60.975 98.45 -60.44 ;
      RECT 98.35 -59.07 98.45 -58.535 ;
      RECT 98.35 -57.745 98.45 -57.21 ;
      RECT 98.35 -55.84 98.45 -55.305 ;
      RECT 98.35 -54.515 98.45 -53.98 ;
      RECT 98.35 -52.61 98.45 -52.075 ;
      RECT 98.35 -51.285 98.45 -50.75 ;
      RECT 98.35 -49.38 98.45 -48.845 ;
      RECT 98.35 -48.055 98.45 -47.52 ;
      RECT 98.35 -46.15 98.45 -45.615 ;
      RECT 98.35 -44.825 98.45 -44.29 ;
      RECT 98.35 -42.92 98.45 -42.385 ;
      RECT 98.35 -41.595 98.45 -41.06 ;
      RECT 98.35 -39.69 98.45 -39.155 ;
      RECT 98.35 -38.365 98.45 -37.83 ;
      RECT 98.35 -36.46 98.45 -35.925 ;
      RECT 98.35 -35.135 98.45 -34.6 ;
      RECT 98.35 -33.23 98.45 -32.695 ;
      RECT 98.35 -31.905 98.45 -31.37 ;
      RECT 98.35 -30 98.45 -29.465 ;
      RECT 98.35 -28.675 98.45 -28.14 ;
      RECT 98.35 -26.77 98.45 -26.235 ;
      RECT 98.35 -25.445 98.45 -24.91 ;
      RECT 98.35 -23.54 98.45 -23.005 ;
      RECT 98.35 -22.215 98.45 -21.68 ;
      RECT 98.35 -20.31 98.45 -19.775 ;
      RECT 98.35 -18.985 98.45 -18.45 ;
      RECT 98.35 -17.08 98.45 -16.545 ;
      RECT 98.35 -15.755 98.45 -15.22 ;
      RECT 98.35 -13.85 98.45 -13.315 ;
      RECT 98.35 -12.525 98.45 -11.99 ;
      RECT 98.35 -10.62 98.45 -10.085 ;
      RECT 98.35 -9.295 98.45 -8.76 ;
      RECT 98.35 -7.39 98.45 -6.855 ;
      RECT 98.35 -6.065 98.45 -5.53 ;
      RECT 98.35 -4.16 98.45 -3.625 ;
      RECT 98.35 -2.835 98.45 -2.3 ;
      RECT 98.35 -0.93 98.45 -0.395 ;
      RECT 98.35 0.395 98.45 0.93 ;
      RECT 98.225 -108.175 98.325 -107.215 ;
      RECT 97.85 -100.19 98.2 -100.07 ;
      RECT 97.85 -96.96 98.2 -96.84 ;
      RECT 97.85 -93.73 98.2 -93.61 ;
      RECT 97.85 -90.5 98.2 -90.38 ;
      RECT 97.85 -87.27 98.2 -87.15 ;
      RECT 97.85 -84.04 98.2 -83.92 ;
      RECT 97.85 -80.81 98.2 -80.69 ;
      RECT 97.85 -77.58 98.2 -77.46 ;
      RECT 97.85 -74.35 98.2 -74.23 ;
      RECT 97.85 -71.12 98.2 -71 ;
      RECT 97.85 -67.89 98.2 -67.77 ;
      RECT 97.85 -64.66 98.2 -64.54 ;
      RECT 97.85 -61.43 98.2 -61.31 ;
      RECT 97.85 -58.2 98.2 -58.08 ;
      RECT 97.85 -54.97 98.2 -54.85 ;
      RECT 97.85 -51.74 98.2 -51.62 ;
      RECT 97.85 -48.51 98.2 -48.39 ;
      RECT 97.85 -45.28 98.2 -45.16 ;
      RECT 97.85 -42.05 98.2 -41.93 ;
      RECT 97.85 -38.82 98.2 -38.7 ;
      RECT 97.85 -35.59 98.2 -35.47 ;
      RECT 97.85 -32.36 98.2 -32.24 ;
      RECT 97.85 -29.13 98.2 -29.01 ;
      RECT 97.85 -25.9 98.2 -25.78 ;
      RECT 97.85 -22.67 98.2 -22.55 ;
      RECT 97.85 -19.44 98.2 -19.32 ;
      RECT 97.85 -16.21 98.2 -16.09 ;
      RECT 97.85 -12.98 98.2 -12.86 ;
      RECT 97.85 -9.75 98.2 -9.63 ;
      RECT 97.85 -6.52 98.2 -6.4 ;
      RECT 97.85 -3.29 98.2 -3.17 ;
      RECT 97.85 -0.06 98.2 0.06 ;
      RECT 98.055 -112.255 98.155 -111.775 ;
      RECT 98.055 -110.765 98.155 -110.295 ;
      RECT 97.965 -108.175 98.065 -107.215 ;
      RECT 97.965 2.175 98.065 3.135 ;
      RECT 97.365 -100.19 97.715 -100.07 ;
      RECT 97.365 -96.96 97.715 -96.84 ;
      RECT 97.365 -93.73 97.715 -93.61 ;
      RECT 97.365 -90.5 97.715 -90.38 ;
      RECT 97.365 -87.27 97.715 -87.15 ;
      RECT 97.365 -84.04 97.715 -83.92 ;
      RECT 97.365 -80.81 97.715 -80.69 ;
      RECT 97.365 -77.58 97.715 -77.46 ;
      RECT 97.365 -74.35 97.715 -74.23 ;
      RECT 97.365 -71.12 97.715 -71 ;
      RECT 97.365 -67.89 97.715 -67.77 ;
      RECT 97.365 -64.66 97.715 -64.54 ;
      RECT 97.365 -61.43 97.715 -61.31 ;
      RECT 97.365 -58.2 97.715 -58.08 ;
      RECT 97.365 -54.97 97.715 -54.85 ;
      RECT 97.365 -51.74 97.715 -51.62 ;
      RECT 97.365 -48.51 97.715 -48.39 ;
      RECT 97.365 -45.28 97.715 -45.16 ;
      RECT 97.365 -42.05 97.715 -41.93 ;
      RECT 97.365 -38.82 97.715 -38.7 ;
      RECT 97.365 -35.59 97.715 -35.47 ;
      RECT 97.365 -32.36 97.715 -32.24 ;
      RECT 97.365 -29.13 97.715 -29.01 ;
      RECT 97.365 -25.9 97.715 -25.78 ;
      RECT 97.365 -22.67 97.715 -22.55 ;
      RECT 97.365 -19.44 97.715 -19.32 ;
      RECT 97.365 -16.21 97.715 -16.09 ;
      RECT 97.365 -12.98 97.715 -12.86 ;
      RECT 97.365 -9.75 97.715 -9.63 ;
      RECT 97.365 -6.52 97.715 -6.4 ;
      RECT 97.365 -3.29 97.715 -3.17 ;
      RECT 97.365 -0.06 97.715 0.06 ;
      RECT 97.535 -108.175 97.635 -107.215 ;
      RECT 97.535 2.175 97.635 3.135 ;
      RECT 97.43 -110.765 97.6 -110.385 ;
      RECT 97.465 -112.245 97.565 -111.775 ;
      RECT 97.275 -108.175 97.375 -107.215 ;
      RECT 97.15 -101.06 97.25 -100.525 ;
      RECT 97.15 -99.735 97.25 -99.2 ;
      RECT 97.15 -97.83 97.25 -97.295 ;
      RECT 97.15 -96.505 97.25 -95.97 ;
      RECT 97.15 -94.6 97.25 -94.065 ;
      RECT 97.15 -93.275 97.25 -92.74 ;
      RECT 97.15 -91.37 97.25 -90.835 ;
      RECT 97.15 -90.045 97.25 -89.51 ;
      RECT 97.15 -88.14 97.25 -87.605 ;
      RECT 97.15 -86.815 97.25 -86.28 ;
      RECT 97.15 -84.91 97.25 -84.375 ;
      RECT 97.15 -83.585 97.25 -83.05 ;
      RECT 97.15 -81.68 97.25 -81.145 ;
      RECT 97.15 -80.355 97.25 -79.82 ;
      RECT 97.15 -78.45 97.25 -77.915 ;
      RECT 97.15 -77.125 97.25 -76.59 ;
      RECT 97.15 -75.22 97.25 -74.685 ;
      RECT 97.15 -73.895 97.25 -73.36 ;
      RECT 97.15 -71.99 97.25 -71.455 ;
      RECT 97.15 -70.665 97.25 -70.13 ;
      RECT 97.15 -68.76 97.25 -68.225 ;
      RECT 97.15 -67.435 97.25 -66.9 ;
      RECT 97.15 -65.53 97.25 -64.995 ;
      RECT 97.15 -64.205 97.25 -63.67 ;
      RECT 97.15 -62.3 97.25 -61.765 ;
      RECT 97.15 -60.975 97.25 -60.44 ;
      RECT 97.15 -59.07 97.25 -58.535 ;
      RECT 97.15 -57.745 97.25 -57.21 ;
      RECT 97.15 -55.84 97.25 -55.305 ;
      RECT 97.15 -54.515 97.25 -53.98 ;
      RECT 97.15 -52.61 97.25 -52.075 ;
      RECT 97.15 -51.285 97.25 -50.75 ;
      RECT 97.15 -49.38 97.25 -48.845 ;
      RECT 97.15 -48.055 97.25 -47.52 ;
      RECT 97.15 -46.15 97.25 -45.615 ;
      RECT 97.15 -44.825 97.25 -44.29 ;
      RECT 97.15 -42.92 97.25 -42.385 ;
      RECT 97.15 -41.595 97.25 -41.06 ;
      RECT 97.15 -39.69 97.25 -39.155 ;
      RECT 97.15 -38.365 97.25 -37.83 ;
      RECT 97.15 -36.46 97.25 -35.925 ;
      RECT 97.15 -35.135 97.25 -34.6 ;
      RECT 97.15 -33.23 97.25 -32.695 ;
      RECT 97.15 -31.905 97.25 -31.37 ;
      RECT 97.15 -30 97.25 -29.465 ;
      RECT 97.15 -28.675 97.25 -28.14 ;
      RECT 97.15 -26.77 97.25 -26.235 ;
      RECT 97.15 -25.445 97.25 -24.91 ;
      RECT 97.15 -23.54 97.25 -23.005 ;
      RECT 97.15 -22.215 97.25 -21.68 ;
      RECT 97.15 -20.31 97.25 -19.775 ;
      RECT 97.15 -18.985 97.25 -18.45 ;
      RECT 97.15 -17.08 97.25 -16.545 ;
      RECT 97.15 -15.755 97.25 -15.22 ;
      RECT 97.15 -13.85 97.25 -13.315 ;
      RECT 97.15 -12.525 97.25 -11.99 ;
      RECT 97.15 -10.62 97.25 -10.085 ;
      RECT 97.15 -9.295 97.25 -8.76 ;
      RECT 97.15 -7.39 97.25 -6.855 ;
      RECT 97.15 -6.065 97.25 -5.53 ;
      RECT 97.15 -4.16 97.25 -3.625 ;
      RECT 97.15 -2.835 97.25 -2.3 ;
      RECT 97.15 -0.93 97.25 -0.395 ;
      RECT 97.15 0.395 97.25 0.93 ;
      RECT 97.025 -108.175 97.125 -107.215 ;
      RECT 96.65 -100.19 97 -100.07 ;
      RECT 96.65 -96.96 97 -96.84 ;
      RECT 96.65 -93.73 97 -93.61 ;
      RECT 96.65 -90.5 97 -90.38 ;
      RECT 96.65 -87.27 97 -87.15 ;
      RECT 96.65 -84.04 97 -83.92 ;
      RECT 96.65 -80.81 97 -80.69 ;
      RECT 96.65 -77.58 97 -77.46 ;
      RECT 96.65 -74.35 97 -74.23 ;
      RECT 96.65 -71.12 97 -71 ;
      RECT 96.65 -67.89 97 -67.77 ;
      RECT 96.65 -64.66 97 -64.54 ;
      RECT 96.65 -61.43 97 -61.31 ;
      RECT 96.65 -58.2 97 -58.08 ;
      RECT 96.65 -54.97 97 -54.85 ;
      RECT 96.65 -51.74 97 -51.62 ;
      RECT 96.65 -48.51 97 -48.39 ;
      RECT 96.65 -45.28 97 -45.16 ;
      RECT 96.65 -42.05 97 -41.93 ;
      RECT 96.65 -38.82 97 -38.7 ;
      RECT 96.65 -35.59 97 -35.47 ;
      RECT 96.65 -32.36 97 -32.24 ;
      RECT 96.65 -29.13 97 -29.01 ;
      RECT 96.65 -25.9 97 -25.78 ;
      RECT 96.65 -22.67 97 -22.55 ;
      RECT 96.65 -19.44 97 -19.32 ;
      RECT 96.65 -16.21 97 -16.09 ;
      RECT 96.65 -12.98 97 -12.86 ;
      RECT 96.65 -9.75 97 -9.63 ;
      RECT 96.65 -6.52 97 -6.4 ;
      RECT 96.65 -3.29 97 -3.17 ;
      RECT 96.65 -0.06 97 0.06 ;
      RECT 96.765 -108.175 96.865 -107.215 ;
      RECT 96.765 2.175 96.865 3.135 ;
      RECT 96.665 -113.555 96.765 -113.085 ;
      RECT 96.165 -100.19 96.515 -100.07 ;
      RECT 96.165 -96.96 96.515 -96.84 ;
      RECT 96.165 -93.73 96.515 -93.61 ;
      RECT 96.165 -90.5 96.515 -90.38 ;
      RECT 96.165 -87.27 96.515 -87.15 ;
      RECT 96.165 -84.04 96.515 -83.92 ;
      RECT 96.165 -80.81 96.515 -80.69 ;
      RECT 96.165 -77.58 96.515 -77.46 ;
      RECT 96.165 -74.35 96.515 -74.23 ;
      RECT 96.165 -71.12 96.515 -71 ;
      RECT 96.165 -67.89 96.515 -67.77 ;
      RECT 96.165 -64.66 96.515 -64.54 ;
      RECT 96.165 -61.43 96.515 -61.31 ;
      RECT 96.165 -58.2 96.515 -58.08 ;
      RECT 96.165 -54.97 96.515 -54.85 ;
      RECT 96.165 -51.74 96.515 -51.62 ;
      RECT 96.165 -48.51 96.515 -48.39 ;
      RECT 96.165 -45.28 96.515 -45.16 ;
      RECT 96.165 -42.05 96.515 -41.93 ;
      RECT 96.165 -38.82 96.515 -38.7 ;
      RECT 96.165 -35.59 96.515 -35.47 ;
      RECT 96.165 -32.36 96.515 -32.24 ;
      RECT 96.165 -29.13 96.515 -29.01 ;
      RECT 96.165 -25.9 96.515 -25.78 ;
      RECT 96.165 -22.67 96.515 -22.55 ;
      RECT 96.165 -19.44 96.515 -19.32 ;
      RECT 96.165 -16.21 96.515 -16.09 ;
      RECT 96.165 -12.98 96.515 -12.86 ;
      RECT 96.165 -9.75 96.515 -9.63 ;
      RECT 96.165 -6.52 96.515 -6.4 ;
      RECT 96.165 -3.29 96.515 -3.17 ;
      RECT 96.165 -0.06 96.515 0.06 ;
      RECT 96.3 -110.735 96.45 -110.445 ;
      RECT 96.335 -108.175 96.435 -107.215 ;
      RECT 96.335 2.175 96.435 3.135 ;
      RECT 96.315 -112.19 96.415 -111.65 ;
      RECT 96.075 -113.555 96.175 -113.085 ;
      RECT 96.075 -108.175 96.175 -107.215 ;
      RECT 95.95 -101.06 96.05 -100.525 ;
      RECT 95.95 -99.735 96.05 -99.2 ;
      RECT 95.95 -97.83 96.05 -97.295 ;
      RECT 95.95 -96.505 96.05 -95.97 ;
      RECT 95.95 -94.6 96.05 -94.065 ;
      RECT 95.95 -93.275 96.05 -92.74 ;
      RECT 95.95 -91.37 96.05 -90.835 ;
      RECT 95.95 -90.045 96.05 -89.51 ;
      RECT 95.95 -88.14 96.05 -87.605 ;
      RECT 95.95 -86.815 96.05 -86.28 ;
      RECT 95.95 -84.91 96.05 -84.375 ;
      RECT 95.95 -83.585 96.05 -83.05 ;
      RECT 95.95 -81.68 96.05 -81.145 ;
      RECT 95.95 -80.355 96.05 -79.82 ;
      RECT 95.95 -78.45 96.05 -77.915 ;
      RECT 95.95 -77.125 96.05 -76.59 ;
      RECT 95.95 -75.22 96.05 -74.685 ;
      RECT 95.95 -73.895 96.05 -73.36 ;
      RECT 95.95 -71.99 96.05 -71.455 ;
      RECT 95.95 -70.665 96.05 -70.13 ;
      RECT 95.95 -68.76 96.05 -68.225 ;
      RECT 95.95 -67.435 96.05 -66.9 ;
      RECT 95.95 -65.53 96.05 -64.995 ;
      RECT 95.95 -64.205 96.05 -63.67 ;
      RECT 95.95 -62.3 96.05 -61.765 ;
      RECT 95.95 -60.975 96.05 -60.44 ;
      RECT 95.95 -59.07 96.05 -58.535 ;
      RECT 95.95 -57.745 96.05 -57.21 ;
      RECT 95.95 -55.84 96.05 -55.305 ;
      RECT 95.95 -54.515 96.05 -53.98 ;
      RECT 95.95 -52.61 96.05 -52.075 ;
      RECT 95.95 -51.285 96.05 -50.75 ;
      RECT 95.95 -49.38 96.05 -48.845 ;
      RECT 95.95 -48.055 96.05 -47.52 ;
      RECT 95.95 -46.15 96.05 -45.615 ;
      RECT 95.95 -44.825 96.05 -44.29 ;
      RECT 95.95 -42.92 96.05 -42.385 ;
      RECT 95.95 -41.595 96.05 -41.06 ;
      RECT 95.95 -39.69 96.05 -39.155 ;
      RECT 95.95 -38.365 96.05 -37.83 ;
      RECT 95.95 -36.46 96.05 -35.925 ;
      RECT 95.95 -35.135 96.05 -34.6 ;
      RECT 95.95 -33.23 96.05 -32.695 ;
      RECT 95.95 -31.905 96.05 -31.37 ;
      RECT 95.95 -30 96.05 -29.465 ;
      RECT 95.95 -28.675 96.05 -28.14 ;
      RECT 95.95 -26.77 96.05 -26.235 ;
      RECT 95.95 -25.445 96.05 -24.91 ;
      RECT 95.95 -23.54 96.05 -23.005 ;
      RECT 95.95 -22.215 96.05 -21.68 ;
      RECT 95.95 -20.31 96.05 -19.775 ;
      RECT 95.95 -18.985 96.05 -18.45 ;
      RECT 95.95 -17.08 96.05 -16.545 ;
      RECT 95.95 -15.755 96.05 -15.22 ;
      RECT 95.95 -13.85 96.05 -13.315 ;
      RECT 95.95 -12.525 96.05 -11.99 ;
      RECT 95.95 -10.62 96.05 -10.085 ;
      RECT 95.95 -9.295 96.05 -8.76 ;
      RECT 95.95 -7.39 96.05 -6.855 ;
      RECT 95.95 -6.065 96.05 -5.53 ;
      RECT 95.95 -4.16 96.05 -3.625 ;
      RECT 95.95 -2.835 96.05 -2.3 ;
      RECT 95.95 -0.93 96.05 -0.395 ;
      RECT 95.95 0.395 96.05 0.93 ;
      RECT 95.825 -104.945 95.925 -103.985 ;
      RECT 95.45 -100.19 95.8 -100.07 ;
      RECT 95.45 -96.96 95.8 -96.84 ;
      RECT 95.45 -93.73 95.8 -93.61 ;
      RECT 95.45 -90.5 95.8 -90.38 ;
      RECT 95.45 -87.27 95.8 -87.15 ;
      RECT 95.45 -84.04 95.8 -83.92 ;
      RECT 95.45 -80.81 95.8 -80.69 ;
      RECT 95.45 -77.58 95.8 -77.46 ;
      RECT 95.45 -74.35 95.8 -74.23 ;
      RECT 95.45 -71.12 95.8 -71 ;
      RECT 95.45 -67.89 95.8 -67.77 ;
      RECT 95.45 -64.66 95.8 -64.54 ;
      RECT 95.45 -61.43 95.8 -61.31 ;
      RECT 95.45 -58.2 95.8 -58.08 ;
      RECT 95.45 -54.97 95.8 -54.85 ;
      RECT 95.45 -51.74 95.8 -51.62 ;
      RECT 95.45 -48.51 95.8 -48.39 ;
      RECT 95.45 -45.28 95.8 -45.16 ;
      RECT 95.45 -42.05 95.8 -41.93 ;
      RECT 95.45 -38.82 95.8 -38.7 ;
      RECT 95.45 -35.59 95.8 -35.47 ;
      RECT 95.45 -32.36 95.8 -32.24 ;
      RECT 95.45 -29.13 95.8 -29.01 ;
      RECT 95.45 -25.9 95.8 -25.78 ;
      RECT 95.45 -22.67 95.8 -22.55 ;
      RECT 95.45 -19.44 95.8 -19.32 ;
      RECT 95.45 -16.21 95.8 -16.09 ;
      RECT 95.45 -12.98 95.8 -12.86 ;
      RECT 95.45 -9.75 95.8 -9.63 ;
      RECT 95.45 -6.52 95.8 -6.4 ;
      RECT 95.45 -3.29 95.8 -3.17 ;
      RECT 95.45 -0.06 95.8 0.06 ;
      RECT 95.565 -104.945 95.665 -103.985 ;
      RECT 95.565 2.175 95.665 3.135 ;
      RECT 95.275 -112.255 95.375 -111.775 ;
      RECT 95.275 -110.765 95.375 -110.295 ;
      RECT 94.965 -100.19 95.315 -100.07 ;
      RECT 94.965 -96.96 95.315 -96.84 ;
      RECT 94.965 -93.73 95.315 -93.61 ;
      RECT 94.965 -90.5 95.315 -90.38 ;
      RECT 94.965 -87.27 95.315 -87.15 ;
      RECT 94.965 -84.04 95.315 -83.92 ;
      RECT 94.965 -80.81 95.315 -80.69 ;
      RECT 94.965 -77.58 95.315 -77.46 ;
      RECT 94.965 -74.35 95.315 -74.23 ;
      RECT 94.965 -71.12 95.315 -71 ;
      RECT 94.965 -67.89 95.315 -67.77 ;
      RECT 94.965 -64.66 95.315 -64.54 ;
      RECT 94.965 -61.43 95.315 -61.31 ;
      RECT 94.965 -58.2 95.315 -58.08 ;
      RECT 94.965 -54.97 95.315 -54.85 ;
      RECT 94.965 -51.74 95.315 -51.62 ;
      RECT 94.965 -48.51 95.315 -48.39 ;
      RECT 94.965 -45.28 95.315 -45.16 ;
      RECT 94.965 -42.05 95.315 -41.93 ;
      RECT 94.965 -38.82 95.315 -38.7 ;
      RECT 94.965 -35.59 95.315 -35.47 ;
      RECT 94.965 -32.36 95.315 -32.24 ;
      RECT 94.965 -29.13 95.315 -29.01 ;
      RECT 94.965 -25.9 95.315 -25.78 ;
      RECT 94.965 -22.67 95.315 -22.55 ;
      RECT 94.965 -19.44 95.315 -19.32 ;
      RECT 94.965 -16.21 95.315 -16.09 ;
      RECT 94.965 -12.98 95.315 -12.86 ;
      RECT 94.965 -9.75 95.315 -9.63 ;
      RECT 94.965 -6.52 95.315 -6.4 ;
      RECT 94.965 -3.29 95.315 -3.17 ;
      RECT 94.965 -0.06 95.315 0.06 ;
      RECT 95.135 -104.945 95.235 -103.985 ;
      RECT 95.135 2.175 95.235 3.135 ;
      RECT 91.235 -108.655 95.015 -108.535 ;
      RECT 94.875 -104.945 94.975 -103.985 ;
      RECT 94.75 -101.06 94.85 -100.525 ;
      RECT 94.75 -99.735 94.85 -99.2 ;
      RECT 94.75 -97.83 94.85 -97.295 ;
      RECT 94.75 -96.505 94.85 -95.97 ;
      RECT 94.75 -94.6 94.85 -94.065 ;
      RECT 94.75 -93.275 94.85 -92.74 ;
      RECT 94.75 -91.37 94.85 -90.835 ;
      RECT 94.75 -90.045 94.85 -89.51 ;
      RECT 94.75 -88.14 94.85 -87.605 ;
      RECT 94.75 -86.815 94.85 -86.28 ;
      RECT 94.75 -84.91 94.85 -84.375 ;
      RECT 94.75 -83.585 94.85 -83.05 ;
      RECT 94.75 -81.68 94.85 -81.145 ;
      RECT 94.75 -80.355 94.85 -79.82 ;
      RECT 94.75 -78.45 94.85 -77.915 ;
      RECT 94.75 -77.125 94.85 -76.59 ;
      RECT 94.75 -75.22 94.85 -74.685 ;
      RECT 94.75 -73.895 94.85 -73.36 ;
      RECT 94.75 -71.99 94.85 -71.455 ;
      RECT 94.75 -70.665 94.85 -70.13 ;
      RECT 94.75 -68.76 94.85 -68.225 ;
      RECT 94.75 -67.435 94.85 -66.9 ;
      RECT 94.75 -65.53 94.85 -64.995 ;
      RECT 94.75 -64.205 94.85 -63.67 ;
      RECT 94.75 -62.3 94.85 -61.765 ;
      RECT 94.75 -60.975 94.85 -60.44 ;
      RECT 94.75 -59.07 94.85 -58.535 ;
      RECT 94.75 -57.745 94.85 -57.21 ;
      RECT 94.75 -55.84 94.85 -55.305 ;
      RECT 94.75 -54.515 94.85 -53.98 ;
      RECT 94.75 -52.61 94.85 -52.075 ;
      RECT 94.75 -51.285 94.85 -50.75 ;
      RECT 94.75 -49.38 94.85 -48.845 ;
      RECT 94.75 -48.055 94.85 -47.52 ;
      RECT 94.75 -46.15 94.85 -45.615 ;
      RECT 94.75 -44.825 94.85 -44.29 ;
      RECT 94.75 -42.92 94.85 -42.385 ;
      RECT 94.75 -41.595 94.85 -41.06 ;
      RECT 94.75 -39.69 94.85 -39.155 ;
      RECT 94.75 -38.365 94.85 -37.83 ;
      RECT 94.75 -36.46 94.85 -35.925 ;
      RECT 94.75 -35.135 94.85 -34.6 ;
      RECT 94.75 -33.23 94.85 -32.695 ;
      RECT 94.75 -31.905 94.85 -31.37 ;
      RECT 94.75 -30 94.85 -29.465 ;
      RECT 94.75 -28.675 94.85 -28.14 ;
      RECT 94.75 -26.77 94.85 -26.235 ;
      RECT 94.75 -25.445 94.85 -24.91 ;
      RECT 94.75 -23.54 94.85 -23.005 ;
      RECT 94.75 -22.215 94.85 -21.68 ;
      RECT 94.75 -20.31 94.85 -19.775 ;
      RECT 94.75 -18.985 94.85 -18.45 ;
      RECT 94.75 -17.08 94.85 -16.545 ;
      RECT 94.75 -15.755 94.85 -15.22 ;
      RECT 94.75 -13.85 94.85 -13.315 ;
      RECT 94.75 -12.525 94.85 -11.99 ;
      RECT 94.75 -10.62 94.85 -10.085 ;
      RECT 94.75 -9.295 94.85 -8.76 ;
      RECT 94.75 -7.39 94.85 -6.855 ;
      RECT 94.75 -6.065 94.85 -5.53 ;
      RECT 94.75 -4.16 94.85 -3.625 ;
      RECT 94.75 -2.835 94.85 -2.3 ;
      RECT 94.75 -0.93 94.85 -0.395 ;
      RECT 94.75 0.395 94.85 0.93 ;
      RECT 94.685 -110.75 94.805 -110.37 ;
      RECT 94.685 -112.245 94.785 -111.775 ;
      RECT 94.625 -104.945 94.725 -103.985 ;
      RECT 94.25 -100.19 94.6 -100.07 ;
      RECT 94.25 -96.96 94.6 -96.84 ;
      RECT 94.25 -93.73 94.6 -93.61 ;
      RECT 94.25 -90.5 94.6 -90.38 ;
      RECT 94.25 -87.27 94.6 -87.15 ;
      RECT 94.25 -84.04 94.6 -83.92 ;
      RECT 94.25 -80.81 94.6 -80.69 ;
      RECT 94.25 -77.58 94.6 -77.46 ;
      RECT 94.25 -74.35 94.6 -74.23 ;
      RECT 94.25 -71.12 94.6 -71 ;
      RECT 94.25 -67.89 94.6 -67.77 ;
      RECT 94.25 -64.66 94.6 -64.54 ;
      RECT 94.25 -61.43 94.6 -61.31 ;
      RECT 94.25 -58.2 94.6 -58.08 ;
      RECT 94.25 -54.97 94.6 -54.85 ;
      RECT 94.25 -51.74 94.6 -51.62 ;
      RECT 94.25 -48.51 94.6 -48.39 ;
      RECT 94.25 -45.28 94.6 -45.16 ;
      RECT 94.25 -42.05 94.6 -41.93 ;
      RECT 94.25 -38.82 94.6 -38.7 ;
      RECT 94.25 -35.59 94.6 -35.47 ;
      RECT 94.25 -32.36 94.6 -32.24 ;
      RECT 94.25 -29.13 94.6 -29.01 ;
      RECT 94.25 -25.9 94.6 -25.78 ;
      RECT 94.25 -22.67 94.6 -22.55 ;
      RECT 94.25 -19.44 94.6 -19.32 ;
      RECT 94.25 -16.21 94.6 -16.09 ;
      RECT 94.25 -12.98 94.6 -12.86 ;
      RECT 94.25 -9.75 94.6 -9.63 ;
      RECT 94.25 -6.52 94.6 -6.4 ;
      RECT 94.25 -3.29 94.6 -3.17 ;
      RECT 94.25 -0.06 94.6 0.06 ;
      RECT 94.365 -104.945 94.465 -103.985 ;
      RECT 94.365 2.175 94.465 3.135 ;
      RECT 94.095 -109.595 94.23 -109.275 ;
      RECT 93.765 -100.19 94.115 -100.07 ;
      RECT 93.765 -96.96 94.115 -96.84 ;
      RECT 93.765 -93.73 94.115 -93.61 ;
      RECT 93.765 -90.5 94.115 -90.38 ;
      RECT 93.765 -87.27 94.115 -87.15 ;
      RECT 93.765 -84.04 94.115 -83.92 ;
      RECT 93.765 -80.81 94.115 -80.69 ;
      RECT 93.765 -77.58 94.115 -77.46 ;
      RECT 93.765 -74.35 94.115 -74.23 ;
      RECT 93.765 -71.12 94.115 -71 ;
      RECT 93.765 -67.89 94.115 -67.77 ;
      RECT 93.765 -64.66 94.115 -64.54 ;
      RECT 93.765 -61.43 94.115 -61.31 ;
      RECT 93.765 -58.2 94.115 -58.08 ;
      RECT 93.765 -54.97 94.115 -54.85 ;
      RECT 93.765 -51.74 94.115 -51.62 ;
      RECT 93.765 -48.51 94.115 -48.39 ;
      RECT 93.765 -45.28 94.115 -45.16 ;
      RECT 93.765 -42.05 94.115 -41.93 ;
      RECT 93.765 -38.82 94.115 -38.7 ;
      RECT 93.765 -35.59 94.115 -35.47 ;
      RECT 93.765 -32.36 94.115 -32.24 ;
      RECT 93.765 -29.13 94.115 -29.01 ;
      RECT 93.765 -25.9 94.115 -25.78 ;
      RECT 93.765 -22.67 94.115 -22.55 ;
      RECT 93.765 -19.44 94.115 -19.32 ;
      RECT 93.765 -16.21 94.115 -16.09 ;
      RECT 93.765 -12.98 94.115 -12.86 ;
      RECT 93.765 -9.75 94.115 -9.63 ;
      RECT 93.765 -6.52 94.115 -6.4 ;
      RECT 93.765 -3.29 94.115 -3.17 ;
      RECT 93.765 -0.06 94.115 0.06 ;
      RECT 93.935 -104.945 94.035 -103.985 ;
      RECT 93.935 2.175 94.035 3.135 ;
      RECT 93.76 -109.595 93.905 -109.275 ;
      RECT 93.675 -104.945 93.775 -103.985 ;
      RECT 93.55 -101.06 93.65 -100.525 ;
      RECT 93.55 -99.735 93.65 -99.2 ;
      RECT 93.55 -97.83 93.65 -97.295 ;
      RECT 93.55 -96.505 93.65 -95.97 ;
      RECT 93.55 -94.6 93.65 -94.065 ;
      RECT 93.55 -93.275 93.65 -92.74 ;
      RECT 93.55 -91.37 93.65 -90.835 ;
      RECT 93.55 -90.045 93.65 -89.51 ;
      RECT 93.55 -88.14 93.65 -87.605 ;
      RECT 93.55 -86.815 93.65 -86.28 ;
      RECT 93.55 -84.91 93.65 -84.375 ;
      RECT 93.55 -83.585 93.65 -83.05 ;
      RECT 93.55 -81.68 93.65 -81.145 ;
      RECT 93.55 -80.355 93.65 -79.82 ;
      RECT 93.55 -78.45 93.65 -77.915 ;
      RECT 93.55 -77.125 93.65 -76.59 ;
      RECT 93.55 -75.22 93.65 -74.685 ;
      RECT 93.55 -73.895 93.65 -73.36 ;
      RECT 93.55 -71.99 93.65 -71.455 ;
      RECT 93.55 -70.665 93.65 -70.13 ;
      RECT 93.55 -68.76 93.65 -68.225 ;
      RECT 93.55 -67.435 93.65 -66.9 ;
      RECT 93.55 -65.53 93.65 -64.995 ;
      RECT 93.55 -64.205 93.65 -63.67 ;
      RECT 93.55 -62.3 93.65 -61.765 ;
      RECT 93.55 -60.975 93.65 -60.44 ;
      RECT 93.55 -59.07 93.65 -58.535 ;
      RECT 93.55 -57.745 93.65 -57.21 ;
      RECT 93.55 -55.84 93.65 -55.305 ;
      RECT 93.55 -54.515 93.65 -53.98 ;
      RECT 93.55 -52.61 93.65 -52.075 ;
      RECT 93.55 -51.285 93.65 -50.75 ;
      RECT 93.55 -49.38 93.65 -48.845 ;
      RECT 93.55 -48.055 93.65 -47.52 ;
      RECT 93.55 -46.15 93.65 -45.615 ;
      RECT 93.55 -44.825 93.65 -44.29 ;
      RECT 93.55 -42.92 93.65 -42.385 ;
      RECT 93.55 -41.595 93.65 -41.06 ;
      RECT 93.55 -39.69 93.65 -39.155 ;
      RECT 93.55 -38.365 93.65 -37.83 ;
      RECT 93.55 -36.46 93.65 -35.925 ;
      RECT 93.55 -35.135 93.65 -34.6 ;
      RECT 93.55 -33.23 93.65 -32.695 ;
      RECT 93.55 -31.905 93.65 -31.37 ;
      RECT 93.55 -30 93.65 -29.465 ;
      RECT 93.55 -28.675 93.65 -28.14 ;
      RECT 93.55 -26.77 93.65 -26.235 ;
      RECT 93.55 -25.445 93.65 -24.91 ;
      RECT 93.55 -23.54 93.65 -23.005 ;
      RECT 93.55 -22.215 93.65 -21.68 ;
      RECT 93.55 -20.31 93.65 -19.775 ;
      RECT 93.55 -18.985 93.65 -18.45 ;
      RECT 93.55 -17.08 93.65 -16.545 ;
      RECT 93.55 -15.755 93.65 -15.22 ;
      RECT 93.55 -13.85 93.65 -13.315 ;
      RECT 93.55 -12.525 93.65 -11.99 ;
      RECT 93.55 -10.62 93.65 -10.085 ;
      RECT 93.55 -9.295 93.65 -8.76 ;
      RECT 93.55 -7.39 93.65 -6.855 ;
      RECT 93.55 -6.065 93.65 -5.53 ;
      RECT 93.55 -4.16 93.65 -3.625 ;
      RECT 93.55 -2.835 93.65 -2.3 ;
      RECT 93.55 -0.93 93.65 -0.395 ;
      RECT 93.55 0.395 93.65 0.93 ;
      RECT 93.425 -108.175 93.525 -107.215 ;
      RECT 93.05 -100.19 93.4 -100.07 ;
      RECT 93.05 -96.96 93.4 -96.84 ;
      RECT 93.05 -93.73 93.4 -93.61 ;
      RECT 93.05 -90.5 93.4 -90.38 ;
      RECT 93.05 -87.27 93.4 -87.15 ;
      RECT 93.05 -84.04 93.4 -83.92 ;
      RECT 93.05 -80.81 93.4 -80.69 ;
      RECT 93.05 -77.58 93.4 -77.46 ;
      RECT 93.05 -74.35 93.4 -74.23 ;
      RECT 93.05 -71.12 93.4 -71 ;
      RECT 93.05 -67.89 93.4 -67.77 ;
      RECT 93.05 -64.66 93.4 -64.54 ;
      RECT 93.05 -61.43 93.4 -61.31 ;
      RECT 93.05 -58.2 93.4 -58.08 ;
      RECT 93.05 -54.97 93.4 -54.85 ;
      RECT 93.05 -51.74 93.4 -51.62 ;
      RECT 93.05 -48.51 93.4 -48.39 ;
      RECT 93.05 -45.28 93.4 -45.16 ;
      RECT 93.05 -42.05 93.4 -41.93 ;
      RECT 93.05 -38.82 93.4 -38.7 ;
      RECT 93.05 -35.59 93.4 -35.47 ;
      RECT 93.05 -32.36 93.4 -32.24 ;
      RECT 93.05 -29.13 93.4 -29.01 ;
      RECT 93.05 -25.9 93.4 -25.78 ;
      RECT 93.05 -22.67 93.4 -22.55 ;
      RECT 93.05 -19.44 93.4 -19.32 ;
      RECT 93.05 -16.21 93.4 -16.09 ;
      RECT 93.05 -12.98 93.4 -12.86 ;
      RECT 93.05 -9.75 93.4 -9.63 ;
      RECT 93.05 -6.52 93.4 -6.4 ;
      RECT 93.05 -3.29 93.4 -3.17 ;
      RECT 93.05 -0.06 93.4 0.06 ;
      RECT 93.255 -112.255 93.355 -111.775 ;
      RECT 93.255 -110.765 93.355 -110.295 ;
      RECT 93.165 -108.175 93.265 -107.215 ;
      RECT 93.165 2.175 93.265 3.135 ;
      RECT 92.565 -100.19 92.915 -100.07 ;
      RECT 92.565 -96.96 92.915 -96.84 ;
      RECT 92.565 -93.73 92.915 -93.61 ;
      RECT 92.565 -90.5 92.915 -90.38 ;
      RECT 92.565 -87.27 92.915 -87.15 ;
      RECT 92.565 -84.04 92.915 -83.92 ;
      RECT 92.565 -80.81 92.915 -80.69 ;
      RECT 92.565 -77.58 92.915 -77.46 ;
      RECT 92.565 -74.35 92.915 -74.23 ;
      RECT 92.565 -71.12 92.915 -71 ;
      RECT 92.565 -67.89 92.915 -67.77 ;
      RECT 92.565 -64.66 92.915 -64.54 ;
      RECT 92.565 -61.43 92.915 -61.31 ;
      RECT 92.565 -58.2 92.915 -58.08 ;
      RECT 92.565 -54.97 92.915 -54.85 ;
      RECT 92.565 -51.74 92.915 -51.62 ;
      RECT 92.565 -48.51 92.915 -48.39 ;
      RECT 92.565 -45.28 92.915 -45.16 ;
      RECT 92.565 -42.05 92.915 -41.93 ;
      RECT 92.565 -38.82 92.915 -38.7 ;
      RECT 92.565 -35.59 92.915 -35.47 ;
      RECT 92.565 -32.36 92.915 -32.24 ;
      RECT 92.565 -29.13 92.915 -29.01 ;
      RECT 92.565 -25.9 92.915 -25.78 ;
      RECT 92.565 -22.67 92.915 -22.55 ;
      RECT 92.565 -19.44 92.915 -19.32 ;
      RECT 92.565 -16.21 92.915 -16.09 ;
      RECT 92.565 -12.98 92.915 -12.86 ;
      RECT 92.565 -9.75 92.915 -9.63 ;
      RECT 92.565 -6.52 92.915 -6.4 ;
      RECT 92.565 -3.29 92.915 -3.17 ;
      RECT 92.565 -0.06 92.915 0.06 ;
      RECT 92.735 -108.175 92.835 -107.215 ;
      RECT 92.735 2.175 92.835 3.135 ;
      RECT 92.63 -110.765 92.8 -110.385 ;
      RECT 92.665 -112.245 92.765 -111.775 ;
      RECT 92.475 -108.175 92.575 -107.215 ;
      RECT 92.35 -101.06 92.45 -100.525 ;
      RECT 92.35 -99.735 92.45 -99.2 ;
      RECT 92.35 -97.83 92.45 -97.295 ;
      RECT 92.35 -96.505 92.45 -95.97 ;
      RECT 92.35 -94.6 92.45 -94.065 ;
      RECT 92.35 -93.275 92.45 -92.74 ;
      RECT 92.35 -91.37 92.45 -90.835 ;
      RECT 92.35 -90.045 92.45 -89.51 ;
      RECT 92.35 -88.14 92.45 -87.605 ;
      RECT 92.35 -86.815 92.45 -86.28 ;
      RECT 92.35 -84.91 92.45 -84.375 ;
      RECT 92.35 -83.585 92.45 -83.05 ;
      RECT 92.35 -81.68 92.45 -81.145 ;
      RECT 92.35 -80.355 92.45 -79.82 ;
      RECT 92.35 -78.45 92.45 -77.915 ;
      RECT 92.35 -77.125 92.45 -76.59 ;
      RECT 92.35 -75.22 92.45 -74.685 ;
      RECT 92.35 -73.895 92.45 -73.36 ;
      RECT 92.35 -71.99 92.45 -71.455 ;
      RECT 92.35 -70.665 92.45 -70.13 ;
      RECT 92.35 -68.76 92.45 -68.225 ;
      RECT 92.35 -67.435 92.45 -66.9 ;
      RECT 92.35 -65.53 92.45 -64.995 ;
      RECT 92.35 -64.205 92.45 -63.67 ;
      RECT 92.35 -62.3 92.45 -61.765 ;
      RECT 92.35 -60.975 92.45 -60.44 ;
      RECT 92.35 -59.07 92.45 -58.535 ;
      RECT 92.35 -57.745 92.45 -57.21 ;
      RECT 92.35 -55.84 92.45 -55.305 ;
      RECT 92.35 -54.515 92.45 -53.98 ;
      RECT 92.35 -52.61 92.45 -52.075 ;
      RECT 92.35 -51.285 92.45 -50.75 ;
      RECT 92.35 -49.38 92.45 -48.845 ;
      RECT 92.35 -48.055 92.45 -47.52 ;
      RECT 92.35 -46.15 92.45 -45.615 ;
      RECT 92.35 -44.825 92.45 -44.29 ;
      RECT 92.35 -42.92 92.45 -42.385 ;
      RECT 92.35 -41.595 92.45 -41.06 ;
      RECT 92.35 -39.69 92.45 -39.155 ;
      RECT 92.35 -38.365 92.45 -37.83 ;
      RECT 92.35 -36.46 92.45 -35.925 ;
      RECT 92.35 -35.135 92.45 -34.6 ;
      RECT 92.35 -33.23 92.45 -32.695 ;
      RECT 92.35 -31.905 92.45 -31.37 ;
      RECT 92.35 -30 92.45 -29.465 ;
      RECT 92.35 -28.675 92.45 -28.14 ;
      RECT 92.35 -26.77 92.45 -26.235 ;
      RECT 92.35 -25.445 92.45 -24.91 ;
      RECT 92.35 -23.54 92.45 -23.005 ;
      RECT 92.35 -22.215 92.45 -21.68 ;
      RECT 92.35 -20.31 92.45 -19.775 ;
      RECT 92.35 -18.985 92.45 -18.45 ;
      RECT 92.35 -17.08 92.45 -16.545 ;
      RECT 92.35 -15.755 92.45 -15.22 ;
      RECT 92.35 -13.85 92.45 -13.315 ;
      RECT 92.35 -12.525 92.45 -11.99 ;
      RECT 92.35 -10.62 92.45 -10.085 ;
      RECT 92.35 -9.295 92.45 -8.76 ;
      RECT 92.35 -7.39 92.45 -6.855 ;
      RECT 92.35 -6.065 92.45 -5.53 ;
      RECT 92.35 -4.16 92.45 -3.625 ;
      RECT 92.35 -2.835 92.45 -2.3 ;
      RECT 92.35 -0.93 92.45 -0.395 ;
      RECT 92.35 0.395 92.45 0.93 ;
      RECT 92.225 -108.175 92.325 -107.215 ;
      RECT 91.85 -100.19 92.2 -100.07 ;
      RECT 91.85 -96.96 92.2 -96.84 ;
      RECT 91.85 -93.73 92.2 -93.61 ;
      RECT 91.85 -90.5 92.2 -90.38 ;
      RECT 91.85 -87.27 92.2 -87.15 ;
      RECT 91.85 -84.04 92.2 -83.92 ;
      RECT 91.85 -80.81 92.2 -80.69 ;
      RECT 91.85 -77.58 92.2 -77.46 ;
      RECT 91.85 -74.35 92.2 -74.23 ;
      RECT 91.85 -71.12 92.2 -71 ;
      RECT 91.85 -67.89 92.2 -67.77 ;
      RECT 91.85 -64.66 92.2 -64.54 ;
      RECT 91.85 -61.43 92.2 -61.31 ;
      RECT 91.85 -58.2 92.2 -58.08 ;
      RECT 91.85 -54.97 92.2 -54.85 ;
      RECT 91.85 -51.74 92.2 -51.62 ;
      RECT 91.85 -48.51 92.2 -48.39 ;
      RECT 91.85 -45.28 92.2 -45.16 ;
      RECT 91.85 -42.05 92.2 -41.93 ;
      RECT 91.85 -38.82 92.2 -38.7 ;
      RECT 91.85 -35.59 92.2 -35.47 ;
      RECT 91.85 -32.36 92.2 -32.24 ;
      RECT 91.85 -29.13 92.2 -29.01 ;
      RECT 91.85 -25.9 92.2 -25.78 ;
      RECT 91.85 -22.67 92.2 -22.55 ;
      RECT 91.85 -19.44 92.2 -19.32 ;
      RECT 91.85 -16.21 92.2 -16.09 ;
      RECT 91.85 -12.98 92.2 -12.86 ;
      RECT 91.85 -9.75 92.2 -9.63 ;
      RECT 91.85 -6.52 92.2 -6.4 ;
      RECT 91.85 -3.29 92.2 -3.17 ;
      RECT 91.85 -0.06 92.2 0.06 ;
      RECT 91.965 -108.175 92.065 -107.215 ;
      RECT 91.965 2.175 92.065 3.135 ;
      RECT 91.865 -113.555 91.965 -113.085 ;
      RECT 91.365 -100.19 91.715 -100.07 ;
      RECT 91.365 -96.96 91.715 -96.84 ;
      RECT 91.365 -93.73 91.715 -93.61 ;
      RECT 91.365 -90.5 91.715 -90.38 ;
      RECT 91.365 -87.27 91.715 -87.15 ;
      RECT 91.365 -84.04 91.715 -83.92 ;
      RECT 91.365 -80.81 91.715 -80.69 ;
      RECT 91.365 -77.58 91.715 -77.46 ;
      RECT 91.365 -74.35 91.715 -74.23 ;
      RECT 91.365 -71.12 91.715 -71 ;
      RECT 91.365 -67.89 91.715 -67.77 ;
      RECT 91.365 -64.66 91.715 -64.54 ;
      RECT 91.365 -61.43 91.715 -61.31 ;
      RECT 91.365 -58.2 91.715 -58.08 ;
      RECT 91.365 -54.97 91.715 -54.85 ;
      RECT 91.365 -51.74 91.715 -51.62 ;
      RECT 91.365 -48.51 91.715 -48.39 ;
      RECT 91.365 -45.28 91.715 -45.16 ;
      RECT 91.365 -42.05 91.715 -41.93 ;
      RECT 91.365 -38.82 91.715 -38.7 ;
      RECT 91.365 -35.59 91.715 -35.47 ;
      RECT 91.365 -32.36 91.715 -32.24 ;
      RECT 91.365 -29.13 91.715 -29.01 ;
      RECT 91.365 -25.9 91.715 -25.78 ;
      RECT 91.365 -22.67 91.715 -22.55 ;
      RECT 91.365 -19.44 91.715 -19.32 ;
      RECT 91.365 -16.21 91.715 -16.09 ;
      RECT 91.365 -12.98 91.715 -12.86 ;
      RECT 91.365 -9.75 91.715 -9.63 ;
      RECT 91.365 -6.52 91.715 -6.4 ;
      RECT 91.365 -3.29 91.715 -3.17 ;
      RECT 91.365 -0.06 91.715 0.06 ;
      RECT 91.5 -110.735 91.65 -110.445 ;
      RECT 91.535 -108.175 91.635 -107.215 ;
      RECT 91.535 2.175 91.635 3.135 ;
      RECT 91.515 -112.19 91.615 -111.65 ;
      RECT 91.275 -113.555 91.375 -113.085 ;
      RECT 91.275 -108.175 91.375 -107.215 ;
      RECT 91.15 -101.06 91.25 -100.525 ;
      RECT 91.15 -99.735 91.25 -99.2 ;
      RECT 91.15 -97.83 91.25 -97.295 ;
      RECT 91.15 -96.505 91.25 -95.97 ;
      RECT 91.15 -94.6 91.25 -94.065 ;
      RECT 91.15 -93.275 91.25 -92.74 ;
      RECT 91.15 -91.37 91.25 -90.835 ;
      RECT 91.15 -90.045 91.25 -89.51 ;
      RECT 91.15 -88.14 91.25 -87.605 ;
      RECT 91.15 -86.815 91.25 -86.28 ;
      RECT 91.15 -84.91 91.25 -84.375 ;
      RECT 91.15 -83.585 91.25 -83.05 ;
      RECT 91.15 -81.68 91.25 -81.145 ;
      RECT 91.15 -80.355 91.25 -79.82 ;
      RECT 91.15 -78.45 91.25 -77.915 ;
      RECT 91.15 -77.125 91.25 -76.59 ;
      RECT 91.15 -75.22 91.25 -74.685 ;
      RECT 91.15 -73.895 91.25 -73.36 ;
      RECT 91.15 -71.99 91.25 -71.455 ;
      RECT 91.15 -70.665 91.25 -70.13 ;
      RECT 91.15 -68.76 91.25 -68.225 ;
      RECT 91.15 -67.435 91.25 -66.9 ;
      RECT 91.15 -65.53 91.25 -64.995 ;
      RECT 91.15 -64.205 91.25 -63.67 ;
      RECT 91.15 -62.3 91.25 -61.765 ;
      RECT 91.15 -60.975 91.25 -60.44 ;
      RECT 91.15 -59.07 91.25 -58.535 ;
      RECT 91.15 -57.745 91.25 -57.21 ;
      RECT 91.15 -55.84 91.25 -55.305 ;
      RECT 91.15 -54.515 91.25 -53.98 ;
      RECT 91.15 -52.61 91.25 -52.075 ;
      RECT 91.15 -51.285 91.25 -50.75 ;
      RECT 91.15 -49.38 91.25 -48.845 ;
      RECT 91.15 -48.055 91.25 -47.52 ;
      RECT 91.15 -46.15 91.25 -45.615 ;
      RECT 91.15 -44.825 91.25 -44.29 ;
      RECT 91.15 -42.92 91.25 -42.385 ;
      RECT 91.15 -41.595 91.25 -41.06 ;
      RECT 91.15 -39.69 91.25 -39.155 ;
      RECT 91.15 -38.365 91.25 -37.83 ;
      RECT 91.15 -36.46 91.25 -35.925 ;
      RECT 91.15 -35.135 91.25 -34.6 ;
      RECT 91.15 -33.23 91.25 -32.695 ;
      RECT 91.15 -31.905 91.25 -31.37 ;
      RECT 91.15 -30 91.25 -29.465 ;
      RECT 91.15 -28.675 91.25 -28.14 ;
      RECT 91.15 -26.77 91.25 -26.235 ;
      RECT 91.15 -25.445 91.25 -24.91 ;
      RECT 91.15 -23.54 91.25 -23.005 ;
      RECT 91.15 -22.215 91.25 -21.68 ;
      RECT 91.15 -20.31 91.25 -19.775 ;
      RECT 91.15 -18.985 91.25 -18.45 ;
      RECT 91.15 -17.08 91.25 -16.545 ;
      RECT 91.15 -15.755 91.25 -15.22 ;
      RECT 91.15 -13.85 91.25 -13.315 ;
      RECT 91.15 -12.525 91.25 -11.99 ;
      RECT 91.15 -10.62 91.25 -10.085 ;
      RECT 91.15 -9.295 91.25 -8.76 ;
      RECT 91.15 -7.39 91.25 -6.855 ;
      RECT 91.15 -6.065 91.25 -5.53 ;
      RECT 91.15 -4.16 91.25 -3.625 ;
      RECT 91.15 -2.835 91.25 -2.3 ;
      RECT 91.15 -0.93 91.25 -0.395 ;
      RECT 91.15 0.395 91.25 0.93 ;
      RECT 91.025 -104.945 91.125 -103.985 ;
      RECT 90.65 -100.19 91 -100.07 ;
      RECT 90.65 -96.96 91 -96.84 ;
      RECT 90.65 -93.73 91 -93.61 ;
      RECT 90.65 -90.5 91 -90.38 ;
      RECT 90.65 -87.27 91 -87.15 ;
      RECT 90.65 -84.04 91 -83.92 ;
      RECT 90.65 -80.81 91 -80.69 ;
      RECT 90.65 -77.58 91 -77.46 ;
      RECT 90.65 -74.35 91 -74.23 ;
      RECT 90.65 -71.12 91 -71 ;
      RECT 90.65 -67.89 91 -67.77 ;
      RECT 90.65 -64.66 91 -64.54 ;
      RECT 90.65 -61.43 91 -61.31 ;
      RECT 90.65 -58.2 91 -58.08 ;
      RECT 90.65 -54.97 91 -54.85 ;
      RECT 90.65 -51.74 91 -51.62 ;
      RECT 90.65 -48.51 91 -48.39 ;
      RECT 90.65 -45.28 91 -45.16 ;
      RECT 90.65 -42.05 91 -41.93 ;
      RECT 90.65 -38.82 91 -38.7 ;
      RECT 90.65 -35.59 91 -35.47 ;
      RECT 90.65 -32.36 91 -32.24 ;
      RECT 90.65 -29.13 91 -29.01 ;
      RECT 90.65 -25.9 91 -25.78 ;
      RECT 90.65 -22.67 91 -22.55 ;
      RECT 90.65 -19.44 91 -19.32 ;
      RECT 90.65 -16.21 91 -16.09 ;
      RECT 90.65 -12.98 91 -12.86 ;
      RECT 90.65 -9.75 91 -9.63 ;
      RECT 90.65 -6.52 91 -6.4 ;
      RECT 90.65 -3.29 91 -3.17 ;
      RECT 90.65 -0.06 91 0.06 ;
      RECT 90.765 -104.945 90.865 -103.985 ;
      RECT 90.765 2.175 90.865 3.135 ;
      RECT 90.475 -112.255 90.575 -111.775 ;
      RECT 90.475 -110.765 90.575 -110.295 ;
      RECT 90.165 -100.19 90.515 -100.07 ;
      RECT 90.165 -96.96 90.515 -96.84 ;
      RECT 90.165 -93.73 90.515 -93.61 ;
      RECT 90.165 -90.5 90.515 -90.38 ;
      RECT 90.165 -87.27 90.515 -87.15 ;
      RECT 90.165 -84.04 90.515 -83.92 ;
      RECT 90.165 -80.81 90.515 -80.69 ;
      RECT 90.165 -77.58 90.515 -77.46 ;
      RECT 90.165 -74.35 90.515 -74.23 ;
      RECT 90.165 -71.12 90.515 -71 ;
      RECT 90.165 -67.89 90.515 -67.77 ;
      RECT 90.165 -64.66 90.515 -64.54 ;
      RECT 90.165 -61.43 90.515 -61.31 ;
      RECT 90.165 -58.2 90.515 -58.08 ;
      RECT 90.165 -54.97 90.515 -54.85 ;
      RECT 90.165 -51.74 90.515 -51.62 ;
      RECT 90.165 -48.51 90.515 -48.39 ;
      RECT 90.165 -45.28 90.515 -45.16 ;
      RECT 90.165 -42.05 90.515 -41.93 ;
      RECT 90.165 -38.82 90.515 -38.7 ;
      RECT 90.165 -35.59 90.515 -35.47 ;
      RECT 90.165 -32.36 90.515 -32.24 ;
      RECT 90.165 -29.13 90.515 -29.01 ;
      RECT 90.165 -25.9 90.515 -25.78 ;
      RECT 90.165 -22.67 90.515 -22.55 ;
      RECT 90.165 -19.44 90.515 -19.32 ;
      RECT 90.165 -16.21 90.515 -16.09 ;
      RECT 90.165 -12.98 90.515 -12.86 ;
      RECT 90.165 -9.75 90.515 -9.63 ;
      RECT 90.165 -6.52 90.515 -6.4 ;
      RECT 90.165 -3.29 90.515 -3.17 ;
      RECT 90.165 -0.06 90.515 0.06 ;
      RECT 90.335 -104.945 90.435 -103.985 ;
      RECT 90.335 2.175 90.435 3.135 ;
      RECT 86.435 -108.655 90.215 -108.535 ;
      RECT 90.075 -104.945 90.175 -103.985 ;
      RECT 89.95 -101.06 90.05 -100.525 ;
      RECT 89.95 -99.735 90.05 -99.2 ;
      RECT 89.95 -97.83 90.05 -97.295 ;
      RECT 89.95 -96.505 90.05 -95.97 ;
      RECT 89.95 -94.6 90.05 -94.065 ;
      RECT 89.95 -93.275 90.05 -92.74 ;
      RECT 89.95 -91.37 90.05 -90.835 ;
      RECT 89.95 -90.045 90.05 -89.51 ;
      RECT 89.95 -88.14 90.05 -87.605 ;
      RECT 89.95 -86.815 90.05 -86.28 ;
      RECT 89.95 -84.91 90.05 -84.375 ;
      RECT 89.95 -83.585 90.05 -83.05 ;
      RECT 89.95 -81.68 90.05 -81.145 ;
      RECT 89.95 -80.355 90.05 -79.82 ;
      RECT 89.95 -78.45 90.05 -77.915 ;
      RECT 89.95 -77.125 90.05 -76.59 ;
      RECT 89.95 -75.22 90.05 -74.685 ;
      RECT 89.95 -73.895 90.05 -73.36 ;
      RECT 89.95 -71.99 90.05 -71.455 ;
      RECT 89.95 -70.665 90.05 -70.13 ;
      RECT 89.95 -68.76 90.05 -68.225 ;
      RECT 89.95 -67.435 90.05 -66.9 ;
      RECT 89.95 -65.53 90.05 -64.995 ;
      RECT 89.95 -64.205 90.05 -63.67 ;
      RECT 89.95 -62.3 90.05 -61.765 ;
      RECT 89.95 -60.975 90.05 -60.44 ;
      RECT 89.95 -59.07 90.05 -58.535 ;
      RECT 89.95 -57.745 90.05 -57.21 ;
      RECT 89.95 -55.84 90.05 -55.305 ;
      RECT 89.95 -54.515 90.05 -53.98 ;
      RECT 89.95 -52.61 90.05 -52.075 ;
      RECT 89.95 -51.285 90.05 -50.75 ;
      RECT 89.95 -49.38 90.05 -48.845 ;
      RECT 89.95 -48.055 90.05 -47.52 ;
      RECT 89.95 -46.15 90.05 -45.615 ;
      RECT 89.95 -44.825 90.05 -44.29 ;
      RECT 89.95 -42.92 90.05 -42.385 ;
      RECT 89.95 -41.595 90.05 -41.06 ;
      RECT 89.95 -39.69 90.05 -39.155 ;
      RECT 89.95 -38.365 90.05 -37.83 ;
      RECT 89.95 -36.46 90.05 -35.925 ;
      RECT 89.95 -35.135 90.05 -34.6 ;
      RECT 89.95 -33.23 90.05 -32.695 ;
      RECT 89.95 -31.905 90.05 -31.37 ;
      RECT 89.95 -30 90.05 -29.465 ;
      RECT 89.95 -28.675 90.05 -28.14 ;
      RECT 89.95 -26.77 90.05 -26.235 ;
      RECT 89.95 -25.445 90.05 -24.91 ;
      RECT 89.95 -23.54 90.05 -23.005 ;
      RECT 89.95 -22.215 90.05 -21.68 ;
      RECT 89.95 -20.31 90.05 -19.775 ;
      RECT 89.95 -18.985 90.05 -18.45 ;
      RECT 89.95 -17.08 90.05 -16.545 ;
      RECT 89.95 -15.755 90.05 -15.22 ;
      RECT 89.95 -13.85 90.05 -13.315 ;
      RECT 89.95 -12.525 90.05 -11.99 ;
      RECT 89.95 -10.62 90.05 -10.085 ;
      RECT 89.95 -9.295 90.05 -8.76 ;
      RECT 89.95 -7.39 90.05 -6.855 ;
      RECT 89.95 -6.065 90.05 -5.53 ;
      RECT 89.95 -4.16 90.05 -3.625 ;
      RECT 89.95 -2.835 90.05 -2.3 ;
      RECT 89.95 -0.93 90.05 -0.395 ;
      RECT 89.95 0.395 90.05 0.93 ;
      RECT 89.885 -110.75 90.005 -110.37 ;
      RECT 89.885 -112.245 89.985 -111.775 ;
      RECT 89.825 -104.945 89.925 -103.985 ;
      RECT 89.45 -100.19 89.8 -100.07 ;
      RECT 89.45 -96.96 89.8 -96.84 ;
      RECT 89.45 -93.73 89.8 -93.61 ;
      RECT 89.45 -90.5 89.8 -90.38 ;
      RECT 89.45 -87.27 89.8 -87.15 ;
      RECT 89.45 -84.04 89.8 -83.92 ;
      RECT 89.45 -80.81 89.8 -80.69 ;
      RECT 89.45 -77.58 89.8 -77.46 ;
      RECT 89.45 -74.35 89.8 -74.23 ;
      RECT 89.45 -71.12 89.8 -71 ;
      RECT 89.45 -67.89 89.8 -67.77 ;
      RECT 89.45 -64.66 89.8 -64.54 ;
      RECT 89.45 -61.43 89.8 -61.31 ;
      RECT 89.45 -58.2 89.8 -58.08 ;
      RECT 89.45 -54.97 89.8 -54.85 ;
      RECT 89.45 -51.74 89.8 -51.62 ;
      RECT 89.45 -48.51 89.8 -48.39 ;
      RECT 89.45 -45.28 89.8 -45.16 ;
      RECT 89.45 -42.05 89.8 -41.93 ;
      RECT 89.45 -38.82 89.8 -38.7 ;
      RECT 89.45 -35.59 89.8 -35.47 ;
      RECT 89.45 -32.36 89.8 -32.24 ;
      RECT 89.45 -29.13 89.8 -29.01 ;
      RECT 89.45 -25.9 89.8 -25.78 ;
      RECT 89.45 -22.67 89.8 -22.55 ;
      RECT 89.45 -19.44 89.8 -19.32 ;
      RECT 89.45 -16.21 89.8 -16.09 ;
      RECT 89.45 -12.98 89.8 -12.86 ;
      RECT 89.45 -9.75 89.8 -9.63 ;
      RECT 89.45 -6.52 89.8 -6.4 ;
      RECT 89.45 -3.29 89.8 -3.17 ;
      RECT 89.45 -0.06 89.8 0.06 ;
      RECT 89.565 -104.945 89.665 -103.985 ;
      RECT 89.565 2.175 89.665 3.135 ;
      RECT 89.295 -109.595 89.43 -109.275 ;
      RECT 88.965 -100.19 89.315 -100.07 ;
      RECT 88.965 -96.96 89.315 -96.84 ;
      RECT 88.965 -93.73 89.315 -93.61 ;
      RECT 88.965 -90.5 89.315 -90.38 ;
      RECT 88.965 -87.27 89.315 -87.15 ;
      RECT 88.965 -84.04 89.315 -83.92 ;
      RECT 88.965 -80.81 89.315 -80.69 ;
      RECT 88.965 -77.58 89.315 -77.46 ;
      RECT 88.965 -74.35 89.315 -74.23 ;
      RECT 88.965 -71.12 89.315 -71 ;
      RECT 88.965 -67.89 89.315 -67.77 ;
      RECT 88.965 -64.66 89.315 -64.54 ;
      RECT 88.965 -61.43 89.315 -61.31 ;
      RECT 88.965 -58.2 89.315 -58.08 ;
      RECT 88.965 -54.97 89.315 -54.85 ;
      RECT 88.965 -51.74 89.315 -51.62 ;
      RECT 88.965 -48.51 89.315 -48.39 ;
      RECT 88.965 -45.28 89.315 -45.16 ;
      RECT 88.965 -42.05 89.315 -41.93 ;
      RECT 88.965 -38.82 89.315 -38.7 ;
      RECT 88.965 -35.59 89.315 -35.47 ;
      RECT 88.965 -32.36 89.315 -32.24 ;
      RECT 88.965 -29.13 89.315 -29.01 ;
      RECT 88.965 -25.9 89.315 -25.78 ;
      RECT 88.965 -22.67 89.315 -22.55 ;
      RECT 88.965 -19.44 89.315 -19.32 ;
      RECT 88.965 -16.21 89.315 -16.09 ;
      RECT 88.965 -12.98 89.315 -12.86 ;
      RECT 88.965 -9.75 89.315 -9.63 ;
      RECT 88.965 -6.52 89.315 -6.4 ;
      RECT 88.965 -3.29 89.315 -3.17 ;
      RECT 88.965 -0.06 89.315 0.06 ;
      RECT 89.135 -104.945 89.235 -103.985 ;
      RECT 89.135 2.175 89.235 3.135 ;
      RECT 88.96 -109.595 89.105 -109.275 ;
      RECT 88.875 -104.945 88.975 -103.985 ;
      RECT 88.75 -101.06 88.85 -100.525 ;
      RECT 88.75 -99.735 88.85 -99.2 ;
      RECT 88.75 -97.83 88.85 -97.295 ;
      RECT 88.75 -96.505 88.85 -95.97 ;
      RECT 88.75 -94.6 88.85 -94.065 ;
      RECT 88.75 -93.275 88.85 -92.74 ;
      RECT 88.75 -91.37 88.85 -90.835 ;
      RECT 88.75 -90.045 88.85 -89.51 ;
      RECT 88.75 -88.14 88.85 -87.605 ;
      RECT 88.75 -86.815 88.85 -86.28 ;
      RECT 88.75 -84.91 88.85 -84.375 ;
      RECT 88.75 -83.585 88.85 -83.05 ;
      RECT 88.75 -81.68 88.85 -81.145 ;
      RECT 88.75 -80.355 88.85 -79.82 ;
      RECT 88.75 -78.45 88.85 -77.915 ;
      RECT 88.75 -77.125 88.85 -76.59 ;
      RECT 88.75 -75.22 88.85 -74.685 ;
      RECT 88.75 -73.895 88.85 -73.36 ;
      RECT 88.75 -71.99 88.85 -71.455 ;
      RECT 88.75 -70.665 88.85 -70.13 ;
      RECT 88.75 -68.76 88.85 -68.225 ;
      RECT 88.75 -67.435 88.85 -66.9 ;
      RECT 88.75 -65.53 88.85 -64.995 ;
      RECT 88.75 -64.205 88.85 -63.67 ;
      RECT 88.75 -62.3 88.85 -61.765 ;
      RECT 88.75 -60.975 88.85 -60.44 ;
      RECT 88.75 -59.07 88.85 -58.535 ;
      RECT 88.75 -57.745 88.85 -57.21 ;
      RECT 88.75 -55.84 88.85 -55.305 ;
      RECT 88.75 -54.515 88.85 -53.98 ;
      RECT 88.75 -52.61 88.85 -52.075 ;
      RECT 88.75 -51.285 88.85 -50.75 ;
      RECT 88.75 -49.38 88.85 -48.845 ;
      RECT 88.75 -48.055 88.85 -47.52 ;
      RECT 88.75 -46.15 88.85 -45.615 ;
      RECT 88.75 -44.825 88.85 -44.29 ;
      RECT 88.75 -42.92 88.85 -42.385 ;
      RECT 88.75 -41.595 88.85 -41.06 ;
      RECT 88.75 -39.69 88.85 -39.155 ;
      RECT 88.75 -38.365 88.85 -37.83 ;
      RECT 88.75 -36.46 88.85 -35.925 ;
      RECT 88.75 -35.135 88.85 -34.6 ;
      RECT 88.75 -33.23 88.85 -32.695 ;
      RECT 88.75 -31.905 88.85 -31.37 ;
      RECT 88.75 -30 88.85 -29.465 ;
      RECT 88.75 -28.675 88.85 -28.14 ;
      RECT 88.75 -26.77 88.85 -26.235 ;
      RECT 88.75 -25.445 88.85 -24.91 ;
      RECT 88.75 -23.54 88.85 -23.005 ;
      RECT 88.75 -22.215 88.85 -21.68 ;
      RECT 88.75 -20.31 88.85 -19.775 ;
      RECT 88.75 -18.985 88.85 -18.45 ;
      RECT 88.75 -17.08 88.85 -16.545 ;
      RECT 88.75 -15.755 88.85 -15.22 ;
      RECT 88.75 -13.85 88.85 -13.315 ;
      RECT 88.75 -12.525 88.85 -11.99 ;
      RECT 88.75 -10.62 88.85 -10.085 ;
      RECT 88.75 -9.295 88.85 -8.76 ;
      RECT 88.75 -7.39 88.85 -6.855 ;
      RECT 88.75 -6.065 88.85 -5.53 ;
      RECT 88.75 -4.16 88.85 -3.625 ;
      RECT 88.75 -2.835 88.85 -2.3 ;
      RECT 88.75 -0.93 88.85 -0.395 ;
      RECT 88.75 0.395 88.85 0.93 ;
      RECT 88.625 -108.175 88.725 -107.215 ;
      RECT 88.25 -100.19 88.6 -100.07 ;
      RECT 88.25 -96.96 88.6 -96.84 ;
      RECT 88.25 -93.73 88.6 -93.61 ;
      RECT 88.25 -90.5 88.6 -90.38 ;
      RECT 88.25 -87.27 88.6 -87.15 ;
      RECT 88.25 -84.04 88.6 -83.92 ;
      RECT 88.25 -80.81 88.6 -80.69 ;
      RECT 88.25 -77.58 88.6 -77.46 ;
      RECT 88.25 -74.35 88.6 -74.23 ;
      RECT 88.25 -71.12 88.6 -71 ;
      RECT 88.25 -67.89 88.6 -67.77 ;
      RECT 88.25 -64.66 88.6 -64.54 ;
      RECT 88.25 -61.43 88.6 -61.31 ;
      RECT 88.25 -58.2 88.6 -58.08 ;
      RECT 88.25 -54.97 88.6 -54.85 ;
      RECT 88.25 -51.74 88.6 -51.62 ;
      RECT 88.25 -48.51 88.6 -48.39 ;
      RECT 88.25 -45.28 88.6 -45.16 ;
      RECT 88.25 -42.05 88.6 -41.93 ;
      RECT 88.25 -38.82 88.6 -38.7 ;
      RECT 88.25 -35.59 88.6 -35.47 ;
      RECT 88.25 -32.36 88.6 -32.24 ;
      RECT 88.25 -29.13 88.6 -29.01 ;
      RECT 88.25 -25.9 88.6 -25.78 ;
      RECT 88.25 -22.67 88.6 -22.55 ;
      RECT 88.25 -19.44 88.6 -19.32 ;
      RECT 88.25 -16.21 88.6 -16.09 ;
      RECT 88.25 -12.98 88.6 -12.86 ;
      RECT 88.25 -9.75 88.6 -9.63 ;
      RECT 88.25 -6.52 88.6 -6.4 ;
      RECT 88.25 -3.29 88.6 -3.17 ;
      RECT 88.25 -0.06 88.6 0.06 ;
      RECT 88.455 -112.255 88.555 -111.775 ;
      RECT 88.455 -110.765 88.555 -110.295 ;
      RECT 88.365 -108.175 88.465 -107.215 ;
      RECT 88.365 2.175 88.465 3.135 ;
      RECT 87.765 -100.19 88.115 -100.07 ;
      RECT 87.765 -96.96 88.115 -96.84 ;
      RECT 87.765 -93.73 88.115 -93.61 ;
      RECT 87.765 -90.5 88.115 -90.38 ;
      RECT 87.765 -87.27 88.115 -87.15 ;
      RECT 87.765 -84.04 88.115 -83.92 ;
      RECT 87.765 -80.81 88.115 -80.69 ;
      RECT 87.765 -77.58 88.115 -77.46 ;
      RECT 87.765 -74.35 88.115 -74.23 ;
      RECT 87.765 -71.12 88.115 -71 ;
      RECT 87.765 -67.89 88.115 -67.77 ;
      RECT 87.765 -64.66 88.115 -64.54 ;
      RECT 87.765 -61.43 88.115 -61.31 ;
      RECT 87.765 -58.2 88.115 -58.08 ;
      RECT 87.765 -54.97 88.115 -54.85 ;
      RECT 87.765 -51.74 88.115 -51.62 ;
      RECT 87.765 -48.51 88.115 -48.39 ;
      RECT 87.765 -45.28 88.115 -45.16 ;
      RECT 87.765 -42.05 88.115 -41.93 ;
      RECT 87.765 -38.82 88.115 -38.7 ;
      RECT 87.765 -35.59 88.115 -35.47 ;
      RECT 87.765 -32.36 88.115 -32.24 ;
      RECT 87.765 -29.13 88.115 -29.01 ;
      RECT 87.765 -25.9 88.115 -25.78 ;
      RECT 87.765 -22.67 88.115 -22.55 ;
      RECT 87.765 -19.44 88.115 -19.32 ;
      RECT 87.765 -16.21 88.115 -16.09 ;
      RECT 87.765 -12.98 88.115 -12.86 ;
      RECT 87.765 -9.75 88.115 -9.63 ;
      RECT 87.765 -6.52 88.115 -6.4 ;
      RECT 87.765 -3.29 88.115 -3.17 ;
      RECT 87.765 -0.06 88.115 0.06 ;
      RECT 87.935 -108.175 88.035 -107.215 ;
      RECT 87.935 2.175 88.035 3.135 ;
      RECT 87.83 -110.765 88 -110.385 ;
      RECT 87.865 -112.245 87.965 -111.775 ;
      RECT 87.675 -108.175 87.775 -107.215 ;
      RECT 87.55 -101.06 87.65 -100.525 ;
      RECT 87.55 -99.735 87.65 -99.2 ;
      RECT 87.55 -97.83 87.65 -97.295 ;
      RECT 87.55 -96.505 87.65 -95.97 ;
      RECT 87.55 -94.6 87.65 -94.065 ;
      RECT 87.55 -93.275 87.65 -92.74 ;
      RECT 87.55 -91.37 87.65 -90.835 ;
      RECT 87.55 -90.045 87.65 -89.51 ;
      RECT 87.55 -88.14 87.65 -87.605 ;
      RECT 87.55 -86.815 87.65 -86.28 ;
      RECT 87.55 -84.91 87.65 -84.375 ;
      RECT 87.55 -83.585 87.65 -83.05 ;
      RECT 87.55 -81.68 87.65 -81.145 ;
      RECT 87.55 -80.355 87.65 -79.82 ;
      RECT 87.55 -78.45 87.65 -77.915 ;
      RECT 87.55 -77.125 87.65 -76.59 ;
      RECT 87.55 -75.22 87.65 -74.685 ;
      RECT 87.55 -73.895 87.65 -73.36 ;
      RECT 87.55 -71.99 87.65 -71.455 ;
      RECT 87.55 -70.665 87.65 -70.13 ;
      RECT 87.55 -68.76 87.65 -68.225 ;
      RECT 87.55 -67.435 87.65 -66.9 ;
      RECT 87.55 -65.53 87.65 -64.995 ;
      RECT 87.55 -64.205 87.65 -63.67 ;
      RECT 87.55 -62.3 87.65 -61.765 ;
      RECT 87.55 -60.975 87.65 -60.44 ;
      RECT 87.55 -59.07 87.65 -58.535 ;
      RECT 87.55 -57.745 87.65 -57.21 ;
      RECT 87.55 -55.84 87.65 -55.305 ;
      RECT 87.55 -54.515 87.65 -53.98 ;
      RECT 87.55 -52.61 87.65 -52.075 ;
      RECT 87.55 -51.285 87.65 -50.75 ;
      RECT 87.55 -49.38 87.65 -48.845 ;
      RECT 87.55 -48.055 87.65 -47.52 ;
      RECT 87.55 -46.15 87.65 -45.615 ;
      RECT 87.55 -44.825 87.65 -44.29 ;
      RECT 87.55 -42.92 87.65 -42.385 ;
      RECT 87.55 -41.595 87.65 -41.06 ;
      RECT 87.55 -39.69 87.65 -39.155 ;
      RECT 87.55 -38.365 87.65 -37.83 ;
      RECT 87.55 -36.46 87.65 -35.925 ;
      RECT 87.55 -35.135 87.65 -34.6 ;
      RECT 87.55 -33.23 87.65 -32.695 ;
      RECT 87.55 -31.905 87.65 -31.37 ;
      RECT 87.55 -30 87.65 -29.465 ;
      RECT 87.55 -28.675 87.65 -28.14 ;
      RECT 87.55 -26.77 87.65 -26.235 ;
      RECT 87.55 -25.445 87.65 -24.91 ;
      RECT 87.55 -23.54 87.65 -23.005 ;
      RECT 87.55 -22.215 87.65 -21.68 ;
      RECT 87.55 -20.31 87.65 -19.775 ;
      RECT 87.55 -18.985 87.65 -18.45 ;
      RECT 87.55 -17.08 87.65 -16.545 ;
      RECT 87.55 -15.755 87.65 -15.22 ;
      RECT 87.55 -13.85 87.65 -13.315 ;
      RECT 87.55 -12.525 87.65 -11.99 ;
      RECT 87.55 -10.62 87.65 -10.085 ;
      RECT 87.55 -9.295 87.65 -8.76 ;
      RECT 87.55 -7.39 87.65 -6.855 ;
      RECT 87.55 -6.065 87.65 -5.53 ;
      RECT 87.55 -4.16 87.65 -3.625 ;
      RECT 87.55 -2.835 87.65 -2.3 ;
      RECT 87.55 -0.93 87.65 -0.395 ;
      RECT 87.55 0.395 87.65 0.93 ;
      RECT 87.425 -108.175 87.525 -107.215 ;
      RECT 87.05 -100.19 87.4 -100.07 ;
      RECT 87.05 -96.96 87.4 -96.84 ;
      RECT 87.05 -93.73 87.4 -93.61 ;
      RECT 87.05 -90.5 87.4 -90.38 ;
      RECT 87.05 -87.27 87.4 -87.15 ;
      RECT 87.05 -84.04 87.4 -83.92 ;
      RECT 87.05 -80.81 87.4 -80.69 ;
      RECT 87.05 -77.58 87.4 -77.46 ;
      RECT 87.05 -74.35 87.4 -74.23 ;
      RECT 87.05 -71.12 87.4 -71 ;
      RECT 87.05 -67.89 87.4 -67.77 ;
      RECT 87.05 -64.66 87.4 -64.54 ;
      RECT 87.05 -61.43 87.4 -61.31 ;
      RECT 87.05 -58.2 87.4 -58.08 ;
      RECT 87.05 -54.97 87.4 -54.85 ;
      RECT 87.05 -51.74 87.4 -51.62 ;
      RECT 87.05 -48.51 87.4 -48.39 ;
      RECT 87.05 -45.28 87.4 -45.16 ;
      RECT 87.05 -42.05 87.4 -41.93 ;
      RECT 87.05 -38.82 87.4 -38.7 ;
      RECT 87.05 -35.59 87.4 -35.47 ;
      RECT 87.05 -32.36 87.4 -32.24 ;
      RECT 87.05 -29.13 87.4 -29.01 ;
      RECT 87.05 -25.9 87.4 -25.78 ;
      RECT 87.05 -22.67 87.4 -22.55 ;
      RECT 87.05 -19.44 87.4 -19.32 ;
      RECT 87.05 -16.21 87.4 -16.09 ;
      RECT 87.05 -12.98 87.4 -12.86 ;
      RECT 87.05 -9.75 87.4 -9.63 ;
      RECT 87.05 -6.52 87.4 -6.4 ;
      RECT 87.05 -3.29 87.4 -3.17 ;
      RECT 87.05 -0.06 87.4 0.06 ;
      RECT 87.165 -108.175 87.265 -107.215 ;
      RECT 87.165 2.175 87.265 3.135 ;
      RECT 87.065 -113.555 87.165 -113.085 ;
      RECT 86.565 -100.19 86.915 -100.07 ;
      RECT 86.565 -96.96 86.915 -96.84 ;
      RECT 86.565 -93.73 86.915 -93.61 ;
      RECT 86.565 -90.5 86.915 -90.38 ;
      RECT 86.565 -87.27 86.915 -87.15 ;
      RECT 86.565 -84.04 86.915 -83.92 ;
      RECT 86.565 -80.81 86.915 -80.69 ;
      RECT 86.565 -77.58 86.915 -77.46 ;
      RECT 86.565 -74.35 86.915 -74.23 ;
      RECT 86.565 -71.12 86.915 -71 ;
      RECT 86.565 -67.89 86.915 -67.77 ;
      RECT 86.565 -64.66 86.915 -64.54 ;
      RECT 86.565 -61.43 86.915 -61.31 ;
      RECT 86.565 -58.2 86.915 -58.08 ;
      RECT 86.565 -54.97 86.915 -54.85 ;
      RECT 86.565 -51.74 86.915 -51.62 ;
      RECT 86.565 -48.51 86.915 -48.39 ;
      RECT 86.565 -45.28 86.915 -45.16 ;
      RECT 86.565 -42.05 86.915 -41.93 ;
      RECT 86.565 -38.82 86.915 -38.7 ;
      RECT 86.565 -35.59 86.915 -35.47 ;
      RECT 86.565 -32.36 86.915 -32.24 ;
      RECT 86.565 -29.13 86.915 -29.01 ;
      RECT 86.565 -25.9 86.915 -25.78 ;
      RECT 86.565 -22.67 86.915 -22.55 ;
      RECT 86.565 -19.44 86.915 -19.32 ;
      RECT 86.565 -16.21 86.915 -16.09 ;
      RECT 86.565 -12.98 86.915 -12.86 ;
      RECT 86.565 -9.75 86.915 -9.63 ;
      RECT 86.565 -6.52 86.915 -6.4 ;
      RECT 86.565 -3.29 86.915 -3.17 ;
      RECT 86.565 -0.06 86.915 0.06 ;
      RECT 86.7 -110.735 86.85 -110.445 ;
      RECT 86.735 -108.175 86.835 -107.215 ;
      RECT 86.735 2.175 86.835 3.135 ;
      RECT 86.715 -112.19 86.815 -111.65 ;
      RECT 86.475 -113.555 86.575 -113.085 ;
      RECT 86.475 -108.175 86.575 -107.215 ;
      RECT 86.35 -101.06 86.45 -100.525 ;
      RECT 86.35 -99.735 86.45 -99.2 ;
      RECT 86.35 -97.83 86.45 -97.295 ;
      RECT 86.35 -96.505 86.45 -95.97 ;
      RECT 86.35 -94.6 86.45 -94.065 ;
      RECT 86.35 -93.275 86.45 -92.74 ;
      RECT 86.35 -91.37 86.45 -90.835 ;
      RECT 86.35 -90.045 86.45 -89.51 ;
      RECT 86.35 -88.14 86.45 -87.605 ;
      RECT 86.35 -86.815 86.45 -86.28 ;
      RECT 86.35 -84.91 86.45 -84.375 ;
      RECT 86.35 -83.585 86.45 -83.05 ;
      RECT 86.35 -81.68 86.45 -81.145 ;
      RECT 86.35 -80.355 86.45 -79.82 ;
      RECT 86.35 -78.45 86.45 -77.915 ;
      RECT 86.35 -77.125 86.45 -76.59 ;
      RECT 86.35 -75.22 86.45 -74.685 ;
      RECT 86.35 -73.895 86.45 -73.36 ;
      RECT 86.35 -71.99 86.45 -71.455 ;
      RECT 86.35 -70.665 86.45 -70.13 ;
      RECT 86.35 -68.76 86.45 -68.225 ;
      RECT 86.35 -67.435 86.45 -66.9 ;
      RECT 86.35 -65.53 86.45 -64.995 ;
      RECT 86.35 -64.205 86.45 -63.67 ;
      RECT 86.35 -62.3 86.45 -61.765 ;
      RECT 86.35 -60.975 86.45 -60.44 ;
      RECT 86.35 -59.07 86.45 -58.535 ;
      RECT 86.35 -57.745 86.45 -57.21 ;
      RECT 86.35 -55.84 86.45 -55.305 ;
      RECT 86.35 -54.515 86.45 -53.98 ;
      RECT 86.35 -52.61 86.45 -52.075 ;
      RECT 86.35 -51.285 86.45 -50.75 ;
      RECT 86.35 -49.38 86.45 -48.845 ;
      RECT 86.35 -48.055 86.45 -47.52 ;
      RECT 86.35 -46.15 86.45 -45.615 ;
      RECT 86.35 -44.825 86.45 -44.29 ;
      RECT 86.35 -42.92 86.45 -42.385 ;
      RECT 86.35 -41.595 86.45 -41.06 ;
      RECT 86.35 -39.69 86.45 -39.155 ;
      RECT 86.35 -38.365 86.45 -37.83 ;
      RECT 86.35 -36.46 86.45 -35.925 ;
      RECT 86.35 -35.135 86.45 -34.6 ;
      RECT 86.35 -33.23 86.45 -32.695 ;
      RECT 86.35 -31.905 86.45 -31.37 ;
      RECT 86.35 -30 86.45 -29.465 ;
      RECT 86.35 -28.675 86.45 -28.14 ;
      RECT 86.35 -26.77 86.45 -26.235 ;
      RECT 86.35 -25.445 86.45 -24.91 ;
      RECT 86.35 -23.54 86.45 -23.005 ;
      RECT 86.35 -22.215 86.45 -21.68 ;
      RECT 86.35 -20.31 86.45 -19.775 ;
      RECT 86.35 -18.985 86.45 -18.45 ;
      RECT 86.35 -17.08 86.45 -16.545 ;
      RECT 86.35 -15.755 86.45 -15.22 ;
      RECT 86.35 -13.85 86.45 -13.315 ;
      RECT 86.35 -12.525 86.45 -11.99 ;
      RECT 86.35 -10.62 86.45 -10.085 ;
      RECT 86.35 -9.295 86.45 -8.76 ;
      RECT 86.35 -7.39 86.45 -6.855 ;
      RECT 86.35 -6.065 86.45 -5.53 ;
      RECT 86.35 -4.16 86.45 -3.625 ;
      RECT 86.35 -2.835 86.45 -2.3 ;
      RECT 86.35 -0.93 86.45 -0.395 ;
      RECT 86.35 0.395 86.45 0.93 ;
      RECT 86.225 -104.945 86.325 -103.985 ;
      RECT 85.85 -100.19 86.2 -100.07 ;
      RECT 85.85 -96.96 86.2 -96.84 ;
      RECT 85.85 -93.73 86.2 -93.61 ;
      RECT 85.85 -90.5 86.2 -90.38 ;
      RECT 85.85 -87.27 86.2 -87.15 ;
      RECT 85.85 -84.04 86.2 -83.92 ;
      RECT 85.85 -80.81 86.2 -80.69 ;
      RECT 85.85 -77.58 86.2 -77.46 ;
      RECT 85.85 -74.35 86.2 -74.23 ;
      RECT 85.85 -71.12 86.2 -71 ;
      RECT 85.85 -67.89 86.2 -67.77 ;
      RECT 85.85 -64.66 86.2 -64.54 ;
      RECT 85.85 -61.43 86.2 -61.31 ;
      RECT 85.85 -58.2 86.2 -58.08 ;
      RECT 85.85 -54.97 86.2 -54.85 ;
      RECT 85.85 -51.74 86.2 -51.62 ;
      RECT 85.85 -48.51 86.2 -48.39 ;
      RECT 85.85 -45.28 86.2 -45.16 ;
      RECT 85.85 -42.05 86.2 -41.93 ;
      RECT 85.85 -38.82 86.2 -38.7 ;
      RECT 85.85 -35.59 86.2 -35.47 ;
      RECT 85.85 -32.36 86.2 -32.24 ;
      RECT 85.85 -29.13 86.2 -29.01 ;
      RECT 85.85 -25.9 86.2 -25.78 ;
      RECT 85.85 -22.67 86.2 -22.55 ;
      RECT 85.85 -19.44 86.2 -19.32 ;
      RECT 85.85 -16.21 86.2 -16.09 ;
      RECT 85.85 -12.98 86.2 -12.86 ;
      RECT 85.85 -9.75 86.2 -9.63 ;
      RECT 85.85 -6.52 86.2 -6.4 ;
      RECT 85.85 -3.29 86.2 -3.17 ;
      RECT 85.85 -0.06 86.2 0.06 ;
      RECT 85.965 -104.945 86.065 -103.985 ;
      RECT 85.965 2.175 86.065 3.135 ;
      RECT 85.675 -112.255 85.775 -111.775 ;
      RECT 85.675 -110.765 85.775 -110.295 ;
      RECT 85.365 -100.19 85.715 -100.07 ;
      RECT 85.365 -96.96 85.715 -96.84 ;
      RECT 85.365 -93.73 85.715 -93.61 ;
      RECT 85.365 -90.5 85.715 -90.38 ;
      RECT 85.365 -87.27 85.715 -87.15 ;
      RECT 85.365 -84.04 85.715 -83.92 ;
      RECT 85.365 -80.81 85.715 -80.69 ;
      RECT 85.365 -77.58 85.715 -77.46 ;
      RECT 85.365 -74.35 85.715 -74.23 ;
      RECT 85.365 -71.12 85.715 -71 ;
      RECT 85.365 -67.89 85.715 -67.77 ;
      RECT 85.365 -64.66 85.715 -64.54 ;
      RECT 85.365 -61.43 85.715 -61.31 ;
      RECT 85.365 -58.2 85.715 -58.08 ;
      RECT 85.365 -54.97 85.715 -54.85 ;
      RECT 85.365 -51.74 85.715 -51.62 ;
      RECT 85.365 -48.51 85.715 -48.39 ;
      RECT 85.365 -45.28 85.715 -45.16 ;
      RECT 85.365 -42.05 85.715 -41.93 ;
      RECT 85.365 -38.82 85.715 -38.7 ;
      RECT 85.365 -35.59 85.715 -35.47 ;
      RECT 85.365 -32.36 85.715 -32.24 ;
      RECT 85.365 -29.13 85.715 -29.01 ;
      RECT 85.365 -25.9 85.715 -25.78 ;
      RECT 85.365 -22.67 85.715 -22.55 ;
      RECT 85.365 -19.44 85.715 -19.32 ;
      RECT 85.365 -16.21 85.715 -16.09 ;
      RECT 85.365 -12.98 85.715 -12.86 ;
      RECT 85.365 -9.75 85.715 -9.63 ;
      RECT 85.365 -6.52 85.715 -6.4 ;
      RECT 85.365 -3.29 85.715 -3.17 ;
      RECT 85.365 -0.06 85.715 0.06 ;
      RECT 85.535 -104.945 85.635 -103.985 ;
      RECT 85.535 2.175 85.635 3.135 ;
      RECT 81.635 -108.655 85.415 -108.535 ;
      RECT 85.275 -104.945 85.375 -103.985 ;
      RECT 85.15 -101.06 85.25 -100.525 ;
      RECT 85.15 -99.735 85.25 -99.2 ;
      RECT 85.15 -97.83 85.25 -97.295 ;
      RECT 85.15 -96.505 85.25 -95.97 ;
      RECT 85.15 -94.6 85.25 -94.065 ;
      RECT 85.15 -93.275 85.25 -92.74 ;
      RECT 85.15 -91.37 85.25 -90.835 ;
      RECT 85.15 -90.045 85.25 -89.51 ;
      RECT 85.15 -88.14 85.25 -87.605 ;
      RECT 85.15 -86.815 85.25 -86.28 ;
      RECT 85.15 -84.91 85.25 -84.375 ;
      RECT 85.15 -83.585 85.25 -83.05 ;
      RECT 85.15 -81.68 85.25 -81.145 ;
      RECT 85.15 -80.355 85.25 -79.82 ;
      RECT 85.15 -78.45 85.25 -77.915 ;
      RECT 85.15 -77.125 85.25 -76.59 ;
      RECT 85.15 -75.22 85.25 -74.685 ;
      RECT 85.15 -73.895 85.25 -73.36 ;
      RECT 85.15 -71.99 85.25 -71.455 ;
      RECT 85.15 -70.665 85.25 -70.13 ;
      RECT 85.15 -68.76 85.25 -68.225 ;
      RECT 85.15 -67.435 85.25 -66.9 ;
      RECT 85.15 -65.53 85.25 -64.995 ;
      RECT 85.15 -64.205 85.25 -63.67 ;
      RECT 85.15 -62.3 85.25 -61.765 ;
      RECT 85.15 -60.975 85.25 -60.44 ;
      RECT 85.15 -59.07 85.25 -58.535 ;
      RECT 85.15 -57.745 85.25 -57.21 ;
      RECT 85.15 -55.84 85.25 -55.305 ;
      RECT 85.15 -54.515 85.25 -53.98 ;
      RECT 85.15 -52.61 85.25 -52.075 ;
      RECT 85.15 -51.285 85.25 -50.75 ;
      RECT 85.15 -49.38 85.25 -48.845 ;
      RECT 85.15 -48.055 85.25 -47.52 ;
      RECT 85.15 -46.15 85.25 -45.615 ;
      RECT 85.15 -44.825 85.25 -44.29 ;
      RECT 85.15 -42.92 85.25 -42.385 ;
      RECT 85.15 -41.595 85.25 -41.06 ;
      RECT 85.15 -39.69 85.25 -39.155 ;
      RECT 85.15 -38.365 85.25 -37.83 ;
      RECT 85.15 -36.46 85.25 -35.925 ;
      RECT 85.15 -35.135 85.25 -34.6 ;
      RECT 85.15 -33.23 85.25 -32.695 ;
      RECT 85.15 -31.905 85.25 -31.37 ;
      RECT 85.15 -30 85.25 -29.465 ;
      RECT 85.15 -28.675 85.25 -28.14 ;
      RECT 85.15 -26.77 85.25 -26.235 ;
      RECT 85.15 -25.445 85.25 -24.91 ;
      RECT 85.15 -23.54 85.25 -23.005 ;
      RECT 85.15 -22.215 85.25 -21.68 ;
      RECT 85.15 -20.31 85.25 -19.775 ;
      RECT 85.15 -18.985 85.25 -18.45 ;
      RECT 85.15 -17.08 85.25 -16.545 ;
      RECT 85.15 -15.755 85.25 -15.22 ;
      RECT 85.15 -13.85 85.25 -13.315 ;
      RECT 85.15 -12.525 85.25 -11.99 ;
      RECT 85.15 -10.62 85.25 -10.085 ;
      RECT 85.15 -9.295 85.25 -8.76 ;
      RECT 85.15 -7.39 85.25 -6.855 ;
      RECT 85.15 -6.065 85.25 -5.53 ;
      RECT 85.15 -4.16 85.25 -3.625 ;
      RECT 85.15 -2.835 85.25 -2.3 ;
      RECT 85.15 -0.93 85.25 -0.395 ;
      RECT 85.15 0.395 85.25 0.93 ;
      RECT 85.085 -110.75 85.205 -110.37 ;
      RECT 85.085 -112.245 85.185 -111.775 ;
      RECT 85.025 -104.945 85.125 -103.985 ;
      RECT 84.65 -100.19 85 -100.07 ;
      RECT 84.65 -96.96 85 -96.84 ;
      RECT 84.65 -93.73 85 -93.61 ;
      RECT 84.65 -90.5 85 -90.38 ;
      RECT 84.65 -87.27 85 -87.15 ;
      RECT 84.65 -84.04 85 -83.92 ;
      RECT 84.65 -80.81 85 -80.69 ;
      RECT 84.65 -77.58 85 -77.46 ;
      RECT 84.65 -74.35 85 -74.23 ;
      RECT 84.65 -71.12 85 -71 ;
      RECT 84.65 -67.89 85 -67.77 ;
      RECT 84.65 -64.66 85 -64.54 ;
      RECT 84.65 -61.43 85 -61.31 ;
      RECT 84.65 -58.2 85 -58.08 ;
      RECT 84.65 -54.97 85 -54.85 ;
      RECT 84.65 -51.74 85 -51.62 ;
      RECT 84.65 -48.51 85 -48.39 ;
      RECT 84.65 -45.28 85 -45.16 ;
      RECT 84.65 -42.05 85 -41.93 ;
      RECT 84.65 -38.82 85 -38.7 ;
      RECT 84.65 -35.59 85 -35.47 ;
      RECT 84.65 -32.36 85 -32.24 ;
      RECT 84.65 -29.13 85 -29.01 ;
      RECT 84.65 -25.9 85 -25.78 ;
      RECT 84.65 -22.67 85 -22.55 ;
      RECT 84.65 -19.44 85 -19.32 ;
      RECT 84.65 -16.21 85 -16.09 ;
      RECT 84.65 -12.98 85 -12.86 ;
      RECT 84.65 -9.75 85 -9.63 ;
      RECT 84.65 -6.52 85 -6.4 ;
      RECT 84.65 -3.29 85 -3.17 ;
      RECT 84.65 -0.06 85 0.06 ;
      RECT 84.765 -104.945 84.865 -103.985 ;
      RECT 84.765 2.175 84.865 3.135 ;
      RECT 84.495 -109.595 84.63 -109.275 ;
      RECT 84.165 -100.19 84.515 -100.07 ;
      RECT 84.165 -96.96 84.515 -96.84 ;
      RECT 84.165 -93.73 84.515 -93.61 ;
      RECT 84.165 -90.5 84.515 -90.38 ;
      RECT 84.165 -87.27 84.515 -87.15 ;
      RECT 84.165 -84.04 84.515 -83.92 ;
      RECT 84.165 -80.81 84.515 -80.69 ;
      RECT 84.165 -77.58 84.515 -77.46 ;
      RECT 84.165 -74.35 84.515 -74.23 ;
      RECT 84.165 -71.12 84.515 -71 ;
      RECT 84.165 -67.89 84.515 -67.77 ;
      RECT 84.165 -64.66 84.515 -64.54 ;
      RECT 84.165 -61.43 84.515 -61.31 ;
      RECT 84.165 -58.2 84.515 -58.08 ;
      RECT 84.165 -54.97 84.515 -54.85 ;
      RECT 84.165 -51.74 84.515 -51.62 ;
      RECT 84.165 -48.51 84.515 -48.39 ;
      RECT 84.165 -45.28 84.515 -45.16 ;
      RECT 84.165 -42.05 84.515 -41.93 ;
      RECT 84.165 -38.82 84.515 -38.7 ;
      RECT 84.165 -35.59 84.515 -35.47 ;
      RECT 84.165 -32.36 84.515 -32.24 ;
      RECT 84.165 -29.13 84.515 -29.01 ;
      RECT 84.165 -25.9 84.515 -25.78 ;
      RECT 84.165 -22.67 84.515 -22.55 ;
      RECT 84.165 -19.44 84.515 -19.32 ;
      RECT 84.165 -16.21 84.515 -16.09 ;
      RECT 84.165 -12.98 84.515 -12.86 ;
      RECT 84.165 -9.75 84.515 -9.63 ;
      RECT 84.165 -6.52 84.515 -6.4 ;
      RECT 84.165 -3.29 84.515 -3.17 ;
      RECT 84.165 -0.06 84.515 0.06 ;
      RECT 84.335 -104.945 84.435 -103.985 ;
      RECT 84.335 2.175 84.435 3.135 ;
      RECT 84.16 -109.595 84.305 -109.275 ;
      RECT 84.075 -104.945 84.175 -103.985 ;
      RECT 83.95 -101.06 84.05 -100.525 ;
      RECT 83.95 -99.735 84.05 -99.2 ;
      RECT 83.95 -97.83 84.05 -97.295 ;
      RECT 83.95 -96.505 84.05 -95.97 ;
      RECT 83.95 -94.6 84.05 -94.065 ;
      RECT 83.95 -93.275 84.05 -92.74 ;
      RECT 83.95 -91.37 84.05 -90.835 ;
      RECT 83.95 -90.045 84.05 -89.51 ;
      RECT 83.95 -88.14 84.05 -87.605 ;
      RECT 83.95 -86.815 84.05 -86.28 ;
      RECT 83.95 -84.91 84.05 -84.375 ;
      RECT 83.95 -83.585 84.05 -83.05 ;
      RECT 83.95 -81.68 84.05 -81.145 ;
      RECT 83.95 -80.355 84.05 -79.82 ;
      RECT 83.95 -78.45 84.05 -77.915 ;
      RECT 83.95 -77.125 84.05 -76.59 ;
      RECT 83.95 -75.22 84.05 -74.685 ;
      RECT 83.95 -73.895 84.05 -73.36 ;
      RECT 83.95 -71.99 84.05 -71.455 ;
      RECT 83.95 -70.665 84.05 -70.13 ;
      RECT 83.95 -68.76 84.05 -68.225 ;
      RECT 83.95 -67.435 84.05 -66.9 ;
      RECT 83.95 -65.53 84.05 -64.995 ;
      RECT 83.95 -64.205 84.05 -63.67 ;
      RECT 83.95 -62.3 84.05 -61.765 ;
      RECT 83.95 -60.975 84.05 -60.44 ;
      RECT 83.95 -59.07 84.05 -58.535 ;
      RECT 83.95 -57.745 84.05 -57.21 ;
      RECT 83.95 -55.84 84.05 -55.305 ;
      RECT 83.95 -54.515 84.05 -53.98 ;
      RECT 83.95 -52.61 84.05 -52.075 ;
      RECT 83.95 -51.285 84.05 -50.75 ;
      RECT 83.95 -49.38 84.05 -48.845 ;
      RECT 83.95 -48.055 84.05 -47.52 ;
      RECT 83.95 -46.15 84.05 -45.615 ;
      RECT 83.95 -44.825 84.05 -44.29 ;
      RECT 83.95 -42.92 84.05 -42.385 ;
      RECT 83.95 -41.595 84.05 -41.06 ;
      RECT 83.95 -39.69 84.05 -39.155 ;
      RECT 83.95 -38.365 84.05 -37.83 ;
      RECT 83.95 -36.46 84.05 -35.925 ;
      RECT 83.95 -35.135 84.05 -34.6 ;
      RECT 83.95 -33.23 84.05 -32.695 ;
      RECT 83.95 -31.905 84.05 -31.37 ;
      RECT 83.95 -30 84.05 -29.465 ;
      RECT 83.95 -28.675 84.05 -28.14 ;
      RECT 83.95 -26.77 84.05 -26.235 ;
      RECT 83.95 -25.445 84.05 -24.91 ;
      RECT 83.95 -23.54 84.05 -23.005 ;
      RECT 83.95 -22.215 84.05 -21.68 ;
      RECT 83.95 -20.31 84.05 -19.775 ;
      RECT 83.95 -18.985 84.05 -18.45 ;
      RECT 83.95 -17.08 84.05 -16.545 ;
      RECT 83.95 -15.755 84.05 -15.22 ;
      RECT 83.95 -13.85 84.05 -13.315 ;
      RECT 83.95 -12.525 84.05 -11.99 ;
      RECT 83.95 -10.62 84.05 -10.085 ;
      RECT 83.95 -9.295 84.05 -8.76 ;
      RECT 83.95 -7.39 84.05 -6.855 ;
      RECT 83.95 -6.065 84.05 -5.53 ;
      RECT 83.95 -4.16 84.05 -3.625 ;
      RECT 83.95 -2.835 84.05 -2.3 ;
      RECT 83.95 -0.93 84.05 -0.395 ;
      RECT 83.95 0.395 84.05 0.93 ;
      RECT 83.825 -108.175 83.925 -107.215 ;
      RECT 83.45 -100.19 83.8 -100.07 ;
      RECT 83.45 -96.96 83.8 -96.84 ;
      RECT 83.45 -93.73 83.8 -93.61 ;
      RECT 83.45 -90.5 83.8 -90.38 ;
      RECT 83.45 -87.27 83.8 -87.15 ;
      RECT 83.45 -84.04 83.8 -83.92 ;
      RECT 83.45 -80.81 83.8 -80.69 ;
      RECT 83.45 -77.58 83.8 -77.46 ;
      RECT 83.45 -74.35 83.8 -74.23 ;
      RECT 83.45 -71.12 83.8 -71 ;
      RECT 83.45 -67.89 83.8 -67.77 ;
      RECT 83.45 -64.66 83.8 -64.54 ;
      RECT 83.45 -61.43 83.8 -61.31 ;
      RECT 83.45 -58.2 83.8 -58.08 ;
      RECT 83.45 -54.97 83.8 -54.85 ;
      RECT 83.45 -51.74 83.8 -51.62 ;
      RECT 83.45 -48.51 83.8 -48.39 ;
      RECT 83.45 -45.28 83.8 -45.16 ;
      RECT 83.45 -42.05 83.8 -41.93 ;
      RECT 83.45 -38.82 83.8 -38.7 ;
      RECT 83.45 -35.59 83.8 -35.47 ;
      RECT 83.45 -32.36 83.8 -32.24 ;
      RECT 83.45 -29.13 83.8 -29.01 ;
      RECT 83.45 -25.9 83.8 -25.78 ;
      RECT 83.45 -22.67 83.8 -22.55 ;
      RECT 83.45 -19.44 83.8 -19.32 ;
      RECT 83.45 -16.21 83.8 -16.09 ;
      RECT 83.45 -12.98 83.8 -12.86 ;
      RECT 83.45 -9.75 83.8 -9.63 ;
      RECT 83.45 -6.52 83.8 -6.4 ;
      RECT 83.45 -3.29 83.8 -3.17 ;
      RECT 83.45 -0.06 83.8 0.06 ;
      RECT 83.655 -112.255 83.755 -111.775 ;
      RECT 83.655 -110.765 83.755 -110.295 ;
      RECT 83.565 -108.175 83.665 -107.215 ;
      RECT 83.565 2.175 83.665 3.135 ;
      RECT 82.965 -100.19 83.315 -100.07 ;
      RECT 82.965 -96.96 83.315 -96.84 ;
      RECT 82.965 -93.73 83.315 -93.61 ;
      RECT 82.965 -90.5 83.315 -90.38 ;
      RECT 82.965 -87.27 83.315 -87.15 ;
      RECT 82.965 -84.04 83.315 -83.92 ;
      RECT 82.965 -80.81 83.315 -80.69 ;
      RECT 82.965 -77.58 83.315 -77.46 ;
      RECT 82.965 -74.35 83.315 -74.23 ;
      RECT 82.965 -71.12 83.315 -71 ;
      RECT 82.965 -67.89 83.315 -67.77 ;
      RECT 82.965 -64.66 83.315 -64.54 ;
      RECT 82.965 -61.43 83.315 -61.31 ;
      RECT 82.965 -58.2 83.315 -58.08 ;
      RECT 82.965 -54.97 83.315 -54.85 ;
      RECT 82.965 -51.74 83.315 -51.62 ;
      RECT 82.965 -48.51 83.315 -48.39 ;
      RECT 82.965 -45.28 83.315 -45.16 ;
      RECT 82.965 -42.05 83.315 -41.93 ;
      RECT 82.965 -38.82 83.315 -38.7 ;
      RECT 82.965 -35.59 83.315 -35.47 ;
      RECT 82.965 -32.36 83.315 -32.24 ;
      RECT 82.965 -29.13 83.315 -29.01 ;
      RECT 82.965 -25.9 83.315 -25.78 ;
      RECT 82.965 -22.67 83.315 -22.55 ;
      RECT 82.965 -19.44 83.315 -19.32 ;
      RECT 82.965 -16.21 83.315 -16.09 ;
      RECT 82.965 -12.98 83.315 -12.86 ;
      RECT 82.965 -9.75 83.315 -9.63 ;
      RECT 82.965 -6.52 83.315 -6.4 ;
      RECT 82.965 -3.29 83.315 -3.17 ;
      RECT 82.965 -0.06 83.315 0.06 ;
      RECT 83.135 -108.175 83.235 -107.215 ;
      RECT 83.135 2.175 83.235 3.135 ;
      RECT 83.03 -110.765 83.2 -110.385 ;
      RECT 83.065 -112.245 83.165 -111.775 ;
      RECT 82.875 -108.175 82.975 -107.215 ;
      RECT 82.75 -101.06 82.85 -100.525 ;
      RECT 82.75 -99.735 82.85 -99.2 ;
      RECT 82.75 -97.83 82.85 -97.295 ;
      RECT 82.75 -96.505 82.85 -95.97 ;
      RECT 82.75 -94.6 82.85 -94.065 ;
      RECT 82.75 -93.275 82.85 -92.74 ;
      RECT 82.75 -91.37 82.85 -90.835 ;
      RECT 82.75 -90.045 82.85 -89.51 ;
      RECT 82.75 -88.14 82.85 -87.605 ;
      RECT 82.75 -86.815 82.85 -86.28 ;
      RECT 82.75 -84.91 82.85 -84.375 ;
      RECT 82.75 -83.585 82.85 -83.05 ;
      RECT 82.75 -81.68 82.85 -81.145 ;
      RECT 82.75 -80.355 82.85 -79.82 ;
      RECT 82.75 -78.45 82.85 -77.915 ;
      RECT 82.75 -77.125 82.85 -76.59 ;
      RECT 82.75 -75.22 82.85 -74.685 ;
      RECT 82.75 -73.895 82.85 -73.36 ;
      RECT 82.75 -71.99 82.85 -71.455 ;
      RECT 82.75 -70.665 82.85 -70.13 ;
      RECT 82.75 -68.76 82.85 -68.225 ;
      RECT 82.75 -67.435 82.85 -66.9 ;
      RECT 82.75 -65.53 82.85 -64.995 ;
      RECT 82.75 -64.205 82.85 -63.67 ;
      RECT 82.75 -62.3 82.85 -61.765 ;
      RECT 82.75 -60.975 82.85 -60.44 ;
      RECT 82.75 -59.07 82.85 -58.535 ;
      RECT 82.75 -57.745 82.85 -57.21 ;
      RECT 82.75 -55.84 82.85 -55.305 ;
      RECT 82.75 -54.515 82.85 -53.98 ;
      RECT 82.75 -52.61 82.85 -52.075 ;
      RECT 82.75 -51.285 82.85 -50.75 ;
      RECT 82.75 -49.38 82.85 -48.845 ;
      RECT 82.75 -48.055 82.85 -47.52 ;
      RECT 82.75 -46.15 82.85 -45.615 ;
      RECT 82.75 -44.825 82.85 -44.29 ;
      RECT 82.75 -42.92 82.85 -42.385 ;
      RECT 82.75 -41.595 82.85 -41.06 ;
      RECT 82.75 -39.69 82.85 -39.155 ;
      RECT 82.75 -38.365 82.85 -37.83 ;
      RECT 82.75 -36.46 82.85 -35.925 ;
      RECT 82.75 -35.135 82.85 -34.6 ;
      RECT 82.75 -33.23 82.85 -32.695 ;
      RECT 82.75 -31.905 82.85 -31.37 ;
      RECT 82.75 -30 82.85 -29.465 ;
      RECT 82.75 -28.675 82.85 -28.14 ;
      RECT 82.75 -26.77 82.85 -26.235 ;
      RECT 82.75 -25.445 82.85 -24.91 ;
      RECT 82.75 -23.54 82.85 -23.005 ;
      RECT 82.75 -22.215 82.85 -21.68 ;
      RECT 82.75 -20.31 82.85 -19.775 ;
      RECT 82.75 -18.985 82.85 -18.45 ;
      RECT 82.75 -17.08 82.85 -16.545 ;
      RECT 82.75 -15.755 82.85 -15.22 ;
      RECT 82.75 -13.85 82.85 -13.315 ;
      RECT 82.75 -12.525 82.85 -11.99 ;
      RECT 82.75 -10.62 82.85 -10.085 ;
      RECT 82.75 -9.295 82.85 -8.76 ;
      RECT 82.75 -7.39 82.85 -6.855 ;
      RECT 82.75 -6.065 82.85 -5.53 ;
      RECT 82.75 -4.16 82.85 -3.625 ;
      RECT 82.75 -2.835 82.85 -2.3 ;
      RECT 82.75 -0.93 82.85 -0.395 ;
      RECT 82.75 0.395 82.85 0.93 ;
      RECT 82.625 -108.175 82.725 -107.215 ;
      RECT 82.25 -100.19 82.6 -100.07 ;
      RECT 82.25 -96.96 82.6 -96.84 ;
      RECT 82.25 -93.73 82.6 -93.61 ;
      RECT 82.25 -90.5 82.6 -90.38 ;
      RECT 82.25 -87.27 82.6 -87.15 ;
      RECT 82.25 -84.04 82.6 -83.92 ;
      RECT 82.25 -80.81 82.6 -80.69 ;
      RECT 82.25 -77.58 82.6 -77.46 ;
      RECT 82.25 -74.35 82.6 -74.23 ;
      RECT 82.25 -71.12 82.6 -71 ;
      RECT 82.25 -67.89 82.6 -67.77 ;
      RECT 82.25 -64.66 82.6 -64.54 ;
      RECT 82.25 -61.43 82.6 -61.31 ;
      RECT 82.25 -58.2 82.6 -58.08 ;
      RECT 82.25 -54.97 82.6 -54.85 ;
      RECT 82.25 -51.74 82.6 -51.62 ;
      RECT 82.25 -48.51 82.6 -48.39 ;
      RECT 82.25 -45.28 82.6 -45.16 ;
      RECT 82.25 -42.05 82.6 -41.93 ;
      RECT 82.25 -38.82 82.6 -38.7 ;
      RECT 82.25 -35.59 82.6 -35.47 ;
      RECT 82.25 -32.36 82.6 -32.24 ;
      RECT 82.25 -29.13 82.6 -29.01 ;
      RECT 82.25 -25.9 82.6 -25.78 ;
      RECT 82.25 -22.67 82.6 -22.55 ;
      RECT 82.25 -19.44 82.6 -19.32 ;
      RECT 82.25 -16.21 82.6 -16.09 ;
      RECT 82.25 -12.98 82.6 -12.86 ;
      RECT 82.25 -9.75 82.6 -9.63 ;
      RECT 82.25 -6.52 82.6 -6.4 ;
      RECT 82.25 -3.29 82.6 -3.17 ;
      RECT 82.25 -0.06 82.6 0.06 ;
      RECT 82.365 -108.175 82.465 -107.215 ;
      RECT 82.365 2.175 82.465 3.135 ;
      RECT 82.265 -113.555 82.365 -113.085 ;
      RECT 81.765 -100.19 82.115 -100.07 ;
      RECT 81.765 -96.96 82.115 -96.84 ;
      RECT 81.765 -93.73 82.115 -93.61 ;
      RECT 81.765 -90.5 82.115 -90.38 ;
      RECT 81.765 -87.27 82.115 -87.15 ;
      RECT 81.765 -84.04 82.115 -83.92 ;
      RECT 81.765 -80.81 82.115 -80.69 ;
      RECT 81.765 -77.58 82.115 -77.46 ;
      RECT 81.765 -74.35 82.115 -74.23 ;
      RECT 81.765 -71.12 82.115 -71 ;
      RECT 81.765 -67.89 82.115 -67.77 ;
      RECT 81.765 -64.66 82.115 -64.54 ;
      RECT 81.765 -61.43 82.115 -61.31 ;
      RECT 81.765 -58.2 82.115 -58.08 ;
      RECT 81.765 -54.97 82.115 -54.85 ;
      RECT 81.765 -51.74 82.115 -51.62 ;
      RECT 81.765 -48.51 82.115 -48.39 ;
      RECT 81.765 -45.28 82.115 -45.16 ;
      RECT 81.765 -42.05 82.115 -41.93 ;
      RECT 81.765 -38.82 82.115 -38.7 ;
      RECT 81.765 -35.59 82.115 -35.47 ;
      RECT 81.765 -32.36 82.115 -32.24 ;
      RECT 81.765 -29.13 82.115 -29.01 ;
      RECT 81.765 -25.9 82.115 -25.78 ;
      RECT 81.765 -22.67 82.115 -22.55 ;
      RECT 81.765 -19.44 82.115 -19.32 ;
      RECT 81.765 -16.21 82.115 -16.09 ;
      RECT 81.765 -12.98 82.115 -12.86 ;
      RECT 81.765 -9.75 82.115 -9.63 ;
      RECT 81.765 -6.52 82.115 -6.4 ;
      RECT 81.765 -3.29 82.115 -3.17 ;
      RECT 81.765 -0.06 82.115 0.06 ;
      RECT 81.9 -110.735 82.05 -110.445 ;
      RECT 81.935 -108.175 82.035 -107.215 ;
      RECT 81.935 2.175 82.035 3.135 ;
      RECT 81.915 -112.19 82.015 -111.65 ;
      RECT 81.675 -113.555 81.775 -113.085 ;
      RECT 81.675 -108.175 81.775 -107.215 ;
      RECT 81.55 -101.06 81.65 -100.525 ;
      RECT 81.55 -99.735 81.65 -99.2 ;
      RECT 81.55 -97.83 81.65 -97.295 ;
      RECT 81.55 -96.505 81.65 -95.97 ;
      RECT 81.55 -94.6 81.65 -94.065 ;
      RECT 81.55 -93.275 81.65 -92.74 ;
      RECT 81.55 -91.37 81.65 -90.835 ;
      RECT 81.55 -90.045 81.65 -89.51 ;
      RECT 81.55 -88.14 81.65 -87.605 ;
      RECT 81.55 -86.815 81.65 -86.28 ;
      RECT 81.55 -84.91 81.65 -84.375 ;
      RECT 81.55 -83.585 81.65 -83.05 ;
      RECT 81.55 -81.68 81.65 -81.145 ;
      RECT 81.55 -80.355 81.65 -79.82 ;
      RECT 81.55 -78.45 81.65 -77.915 ;
      RECT 81.55 -77.125 81.65 -76.59 ;
      RECT 81.55 -75.22 81.65 -74.685 ;
      RECT 81.55 -73.895 81.65 -73.36 ;
      RECT 81.55 -71.99 81.65 -71.455 ;
      RECT 81.55 -70.665 81.65 -70.13 ;
      RECT 81.55 -68.76 81.65 -68.225 ;
      RECT 81.55 -67.435 81.65 -66.9 ;
      RECT 81.55 -65.53 81.65 -64.995 ;
      RECT 81.55 -64.205 81.65 -63.67 ;
      RECT 81.55 -62.3 81.65 -61.765 ;
      RECT 81.55 -60.975 81.65 -60.44 ;
      RECT 81.55 -59.07 81.65 -58.535 ;
      RECT 81.55 -57.745 81.65 -57.21 ;
      RECT 81.55 -55.84 81.65 -55.305 ;
      RECT 81.55 -54.515 81.65 -53.98 ;
      RECT 81.55 -52.61 81.65 -52.075 ;
      RECT 81.55 -51.285 81.65 -50.75 ;
      RECT 81.55 -49.38 81.65 -48.845 ;
      RECT 81.55 -48.055 81.65 -47.52 ;
      RECT 81.55 -46.15 81.65 -45.615 ;
      RECT 81.55 -44.825 81.65 -44.29 ;
      RECT 81.55 -42.92 81.65 -42.385 ;
      RECT 81.55 -41.595 81.65 -41.06 ;
      RECT 81.55 -39.69 81.65 -39.155 ;
      RECT 81.55 -38.365 81.65 -37.83 ;
      RECT 81.55 -36.46 81.65 -35.925 ;
      RECT 81.55 -35.135 81.65 -34.6 ;
      RECT 81.55 -33.23 81.65 -32.695 ;
      RECT 81.55 -31.905 81.65 -31.37 ;
      RECT 81.55 -30 81.65 -29.465 ;
      RECT 81.55 -28.675 81.65 -28.14 ;
      RECT 81.55 -26.77 81.65 -26.235 ;
      RECT 81.55 -25.445 81.65 -24.91 ;
      RECT 81.55 -23.54 81.65 -23.005 ;
      RECT 81.55 -22.215 81.65 -21.68 ;
      RECT 81.55 -20.31 81.65 -19.775 ;
      RECT 81.55 -18.985 81.65 -18.45 ;
      RECT 81.55 -17.08 81.65 -16.545 ;
      RECT 81.55 -15.755 81.65 -15.22 ;
      RECT 81.55 -13.85 81.65 -13.315 ;
      RECT 81.55 -12.525 81.65 -11.99 ;
      RECT 81.55 -10.62 81.65 -10.085 ;
      RECT 81.55 -9.295 81.65 -8.76 ;
      RECT 81.55 -7.39 81.65 -6.855 ;
      RECT 81.55 -6.065 81.65 -5.53 ;
      RECT 81.55 -4.16 81.65 -3.625 ;
      RECT 81.55 -2.835 81.65 -2.3 ;
      RECT 81.55 -0.93 81.65 -0.395 ;
      RECT 81.55 0.395 81.65 0.93 ;
      RECT 81.425 -104.945 81.525 -103.985 ;
      RECT 81.05 -100.19 81.4 -100.07 ;
      RECT 81.05 -96.96 81.4 -96.84 ;
      RECT 81.05 -93.73 81.4 -93.61 ;
      RECT 81.05 -90.5 81.4 -90.38 ;
      RECT 81.05 -87.27 81.4 -87.15 ;
      RECT 81.05 -84.04 81.4 -83.92 ;
      RECT 81.05 -80.81 81.4 -80.69 ;
      RECT 81.05 -77.58 81.4 -77.46 ;
      RECT 81.05 -74.35 81.4 -74.23 ;
      RECT 81.05 -71.12 81.4 -71 ;
      RECT 81.05 -67.89 81.4 -67.77 ;
      RECT 81.05 -64.66 81.4 -64.54 ;
      RECT 81.05 -61.43 81.4 -61.31 ;
      RECT 81.05 -58.2 81.4 -58.08 ;
      RECT 81.05 -54.97 81.4 -54.85 ;
      RECT 81.05 -51.74 81.4 -51.62 ;
      RECT 81.05 -48.51 81.4 -48.39 ;
      RECT 81.05 -45.28 81.4 -45.16 ;
      RECT 81.05 -42.05 81.4 -41.93 ;
      RECT 81.05 -38.82 81.4 -38.7 ;
      RECT 81.05 -35.59 81.4 -35.47 ;
      RECT 81.05 -32.36 81.4 -32.24 ;
      RECT 81.05 -29.13 81.4 -29.01 ;
      RECT 81.05 -25.9 81.4 -25.78 ;
      RECT 81.05 -22.67 81.4 -22.55 ;
      RECT 81.05 -19.44 81.4 -19.32 ;
      RECT 81.05 -16.21 81.4 -16.09 ;
      RECT 81.05 -12.98 81.4 -12.86 ;
      RECT 81.05 -9.75 81.4 -9.63 ;
      RECT 81.05 -6.52 81.4 -6.4 ;
      RECT 81.05 -3.29 81.4 -3.17 ;
      RECT 81.05 -0.06 81.4 0.06 ;
      RECT 81.165 -104.945 81.265 -103.985 ;
      RECT 81.165 2.175 81.265 3.135 ;
      RECT 80.875 -112.255 80.975 -111.775 ;
      RECT 80.875 -110.765 80.975 -110.295 ;
      RECT 80.565 -100.19 80.915 -100.07 ;
      RECT 80.565 -96.96 80.915 -96.84 ;
      RECT 80.565 -93.73 80.915 -93.61 ;
      RECT 80.565 -90.5 80.915 -90.38 ;
      RECT 80.565 -87.27 80.915 -87.15 ;
      RECT 80.565 -84.04 80.915 -83.92 ;
      RECT 80.565 -80.81 80.915 -80.69 ;
      RECT 80.565 -77.58 80.915 -77.46 ;
      RECT 80.565 -74.35 80.915 -74.23 ;
      RECT 80.565 -71.12 80.915 -71 ;
      RECT 80.565 -67.89 80.915 -67.77 ;
      RECT 80.565 -64.66 80.915 -64.54 ;
      RECT 80.565 -61.43 80.915 -61.31 ;
      RECT 80.565 -58.2 80.915 -58.08 ;
      RECT 80.565 -54.97 80.915 -54.85 ;
      RECT 80.565 -51.74 80.915 -51.62 ;
      RECT 80.565 -48.51 80.915 -48.39 ;
      RECT 80.565 -45.28 80.915 -45.16 ;
      RECT 80.565 -42.05 80.915 -41.93 ;
      RECT 80.565 -38.82 80.915 -38.7 ;
      RECT 80.565 -35.59 80.915 -35.47 ;
      RECT 80.565 -32.36 80.915 -32.24 ;
      RECT 80.565 -29.13 80.915 -29.01 ;
      RECT 80.565 -25.9 80.915 -25.78 ;
      RECT 80.565 -22.67 80.915 -22.55 ;
      RECT 80.565 -19.44 80.915 -19.32 ;
      RECT 80.565 -16.21 80.915 -16.09 ;
      RECT 80.565 -12.98 80.915 -12.86 ;
      RECT 80.565 -9.75 80.915 -9.63 ;
      RECT 80.565 -6.52 80.915 -6.4 ;
      RECT 80.565 -3.29 80.915 -3.17 ;
      RECT 80.565 -0.06 80.915 0.06 ;
      RECT 80.735 -104.945 80.835 -103.985 ;
      RECT 80.735 2.175 80.835 3.135 ;
      RECT 76.835 -108.655 80.615 -108.535 ;
      RECT 80.475 -104.945 80.575 -103.985 ;
      RECT 80.35 -101.06 80.45 -100.525 ;
      RECT 80.35 -99.735 80.45 -99.2 ;
      RECT 80.35 -97.83 80.45 -97.295 ;
      RECT 80.35 -96.505 80.45 -95.97 ;
      RECT 80.35 -94.6 80.45 -94.065 ;
      RECT 80.35 -93.275 80.45 -92.74 ;
      RECT 80.35 -91.37 80.45 -90.835 ;
      RECT 80.35 -90.045 80.45 -89.51 ;
      RECT 80.35 -88.14 80.45 -87.605 ;
      RECT 80.35 -86.815 80.45 -86.28 ;
      RECT 80.35 -84.91 80.45 -84.375 ;
      RECT 80.35 -83.585 80.45 -83.05 ;
      RECT 80.35 -81.68 80.45 -81.145 ;
      RECT 80.35 -80.355 80.45 -79.82 ;
      RECT 80.35 -78.45 80.45 -77.915 ;
      RECT 80.35 -77.125 80.45 -76.59 ;
      RECT 80.35 -75.22 80.45 -74.685 ;
      RECT 80.35 -73.895 80.45 -73.36 ;
      RECT 80.35 -71.99 80.45 -71.455 ;
      RECT 80.35 -70.665 80.45 -70.13 ;
      RECT 80.35 -68.76 80.45 -68.225 ;
      RECT 80.35 -67.435 80.45 -66.9 ;
      RECT 80.35 -65.53 80.45 -64.995 ;
      RECT 80.35 -64.205 80.45 -63.67 ;
      RECT 80.35 -62.3 80.45 -61.765 ;
      RECT 80.35 -60.975 80.45 -60.44 ;
      RECT 80.35 -59.07 80.45 -58.535 ;
      RECT 80.35 -57.745 80.45 -57.21 ;
      RECT 80.35 -55.84 80.45 -55.305 ;
      RECT 80.35 -54.515 80.45 -53.98 ;
      RECT 80.35 -52.61 80.45 -52.075 ;
      RECT 80.35 -51.285 80.45 -50.75 ;
      RECT 80.35 -49.38 80.45 -48.845 ;
      RECT 80.35 -48.055 80.45 -47.52 ;
      RECT 80.35 -46.15 80.45 -45.615 ;
      RECT 80.35 -44.825 80.45 -44.29 ;
      RECT 80.35 -42.92 80.45 -42.385 ;
      RECT 80.35 -41.595 80.45 -41.06 ;
      RECT 80.35 -39.69 80.45 -39.155 ;
      RECT 80.35 -38.365 80.45 -37.83 ;
      RECT 80.35 -36.46 80.45 -35.925 ;
      RECT 80.35 -35.135 80.45 -34.6 ;
      RECT 80.35 -33.23 80.45 -32.695 ;
      RECT 80.35 -31.905 80.45 -31.37 ;
      RECT 80.35 -30 80.45 -29.465 ;
      RECT 80.35 -28.675 80.45 -28.14 ;
      RECT 80.35 -26.77 80.45 -26.235 ;
      RECT 80.35 -25.445 80.45 -24.91 ;
      RECT 80.35 -23.54 80.45 -23.005 ;
      RECT 80.35 -22.215 80.45 -21.68 ;
      RECT 80.35 -20.31 80.45 -19.775 ;
      RECT 80.35 -18.985 80.45 -18.45 ;
      RECT 80.35 -17.08 80.45 -16.545 ;
      RECT 80.35 -15.755 80.45 -15.22 ;
      RECT 80.35 -13.85 80.45 -13.315 ;
      RECT 80.35 -12.525 80.45 -11.99 ;
      RECT 80.35 -10.62 80.45 -10.085 ;
      RECT 80.35 -9.295 80.45 -8.76 ;
      RECT 80.35 -7.39 80.45 -6.855 ;
      RECT 80.35 -6.065 80.45 -5.53 ;
      RECT 80.35 -4.16 80.45 -3.625 ;
      RECT 80.35 -2.835 80.45 -2.3 ;
      RECT 80.35 -0.93 80.45 -0.395 ;
      RECT 80.35 0.395 80.45 0.93 ;
      RECT 80.285 -110.75 80.405 -110.37 ;
      RECT 80.285 -112.245 80.385 -111.775 ;
      RECT 80.225 -104.945 80.325 -103.985 ;
      RECT 79.85 -100.19 80.2 -100.07 ;
      RECT 79.85 -96.96 80.2 -96.84 ;
      RECT 79.85 -93.73 80.2 -93.61 ;
      RECT 79.85 -90.5 80.2 -90.38 ;
      RECT 79.85 -87.27 80.2 -87.15 ;
      RECT 79.85 -84.04 80.2 -83.92 ;
      RECT 79.85 -80.81 80.2 -80.69 ;
      RECT 79.85 -77.58 80.2 -77.46 ;
      RECT 79.85 -74.35 80.2 -74.23 ;
      RECT 79.85 -71.12 80.2 -71 ;
      RECT 79.85 -67.89 80.2 -67.77 ;
      RECT 79.85 -64.66 80.2 -64.54 ;
      RECT 79.85 -61.43 80.2 -61.31 ;
      RECT 79.85 -58.2 80.2 -58.08 ;
      RECT 79.85 -54.97 80.2 -54.85 ;
      RECT 79.85 -51.74 80.2 -51.62 ;
      RECT 79.85 -48.51 80.2 -48.39 ;
      RECT 79.85 -45.28 80.2 -45.16 ;
      RECT 79.85 -42.05 80.2 -41.93 ;
      RECT 79.85 -38.82 80.2 -38.7 ;
      RECT 79.85 -35.59 80.2 -35.47 ;
      RECT 79.85 -32.36 80.2 -32.24 ;
      RECT 79.85 -29.13 80.2 -29.01 ;
      RECT 79.85 -25.9 80.2 -25.78 ;
      RECT 79.85 -22.67 80.2 -22.55 ;
      RECT 79.85 -19.44 80.2 -19.32 ;
      RECT 79.85 -16.21 80.2 -16.09 ;
      RECT 79.85 -12.98 80.2 -12.86 ;
      RECT 79.85 -9.75 80.2 -9.63 ;
      RECT 79.85 -6.52 80.2 -6.4 ;
      RECT 79.85 -3.29 80.2 -3.17 ;
      RECT 79.85 -0.06 80.2 0.06 ;
      RECT 79.965 -104.945 80.065 -103.985 ;
      RECT 79.965 2.175 80.065 3.135 ;
      RECT 79.695 -109.595 79.83 -109.275 ;
      RECT 79.365 -100.19 79.715 -100.07 ;
      RECT 79.365 -96.96 79.715 -96.84 ;
      RECT 79.365 -93.73 79.715 -93.61 ;
      RECT 79.365 -90.5 79.715 -90.38 ;
      RECT 79.365 -87.27 79.715 -87.15 ;
      RECT 79.365 -84.04 79.715 -83.92 ;
      RECT 79.365 -80.81 79.715 -80.69 ;
      RECT 79.365 -77.58 79.715 -77.46 ;
      RECT 79.365 -74.35 79.715 -74.23 ;
      RECT 79.365 -71.12 79.715 -71 ;
      RECT 79.365 -67.89 79.715 -67.77 ;
      RECT 79.365 -64.66 79.715 -64.54 ;
      RECT 79.365 -61.43 79.715 -61.31 ;
      RECT 79.365 -58.2 79.715 -58.08 ;
      RECT 79.365 -54.97 79.715 -54.85 ;
      RECT 79.365 -51.74 79.715 -51.62 ;
      RECT 79.365 -48.51 79.715 -48.39 ;
      RECT 79.365 -45.28 79.715 -45.16 ;
      RECT 79.365 -42.05 79.715 -41.93 ;
      RECT 79.365 -38.82 79.715 -38.7 ;
      RECT 79.365 -35.59 79.715 -35.47 ;
      RECT 79.365 -32.36 79.715 -32.24 ;
      RECT 79.365 -29.13 79.715 -29.01 ;
      RECT 79.365 -25.9 79.715 -25.78 ;
      RECT 79.365 -22.67 79.715 -22.55 ;
      RECT 79.365 -19.44 79.715 -19.32 ;
      RECT 79.365 -16.21 79.715 -16.09 ;
      RECT 79.365 -12.98 79.715 -12.86 ;
      RECT 79.365 -9.75 79.715 -9.63 ;
      RECT 79.365 -6.52 79.715 -6.4 ;
      RECT 79.365 -3.29 79.715 -3.17 ;
      RECT 79.365 -0.06 79.715 0.06 ;
      RECT 79.535 -104.945 79.635 -103.985 ;
      RECT 79.535 2.175 79.635 3.135 ;
      RECT 79.36 -109.595 79.505 -109.275 ;
      RECT 79.275 -104.945 79.375 -103.985 ;
      RECT 79.15 -101.06 79.25 -100.525 ;
      RECT 79.15 -99.735 79.25 -99.2 ;
      RECT 79.15 -97.83 79.25 -97.295 ;
      RECT 79.15 -96.505 79.25 -95.97 ;
      RECT 79.15 -94.6 79.25 -94.065 ;
      RECT 79.15 -93.275 79.25 -92.74 ;
      RECT 79.15 -91.37 79.25 -90.835 ;
      RECT 79.15 -90.045 79.25 -89.51 ;
      RECT 79.15 -88.14 79.25 -87.605 ;
      RECT 79.15 -86.815 79.25 -86.28 ;
      RECT 79.15 -84.91 79.25 -84.375 ;
      RECT 79.15 -83.585 79.25 -83.05 ;
      RECT 79.15 -81.68 79.25 -81.145 ;
      RECT 79.15 -80.355 79.25 -79.82 ;
      RECT 79.15 -78.45 79.25 -77.915 ;
      RECT 79.15 -77.125 79.25 -76.59 ;
      RECT 79.15 -75.22 79.25 -74.685 ;
      RECT 79.15 -73.895 79.25 -73.36 ;
      RECT 79.15 -71.99 79.25 -71.455 ;
      RECT 79.15 -70.665 79.25 -70.13 ;
      RECT 79.15 -68.76 79.25 -68.225 ;
      RECT 79.15 -67.435 79.25 -66.9 ;
      RECT 79.15 -65.53 79.25 -64.995 ;
      RECT 79.15 -64.205 79.25 -63.67 ;
      RECT 79.15 -62.3 79.25 -61.765 ;
      RECT 79.15 -60.975 79.25 -60.44 ;
      RECT 79.15 -59.07 79.25 -58.535 ;
      RECT 79.15 -57.745 79.25 -57.21 ;
      RECT 79.15 -55.84 79.25 -55.305 ;
      RECT 79.15 -54.515 79.25 -53.98 ;
      RECT 79.15 -52.61 79.25 -52.075 ;
      RECT 79.15 -51.285 79.25 -50.75 ;
      RECT 79.15 -49.38 79.25 -48.845 ;
      RECT 79.15 -48.055 79.25 -47.52 ;
      RECT 79.15 -46.15 79.25 -45.615 ;
      RECT 79.15 -44.825 79.25 -44.29 ;
      RECT 79.15 -42.92 79.25 -42.385 ;
      RECT 79.15 -41.595 79.25 -41.06 ;
      RECT 79.15 -39.69 79.25 -39.155 ;
      RECT 79.15 -38.365 79.25 -37.83 ;
      RECT 79.15 -36.46 79.25 -35.925 ;
      RECT 79.15 -35.135 79.25 -34.6 ;
      RECT 79.15 -33.23 79.25 -32.695 ;
      RECT 79.15 -31.905 79.25 -31.37 ;
      RECT 79.15 -30 79.25 -29.465 ;
      RECT 79.15 -28.675 79.25 -28.14 ;
      RECT 79.15 -26.77 79.25 -26.235 ;
      RECT 79.15 -25.445 79.25 -24.91 ;
      RECT 79.15 -23.54 79.25 -23.005 ;
      RECT 79.15 -22.215 79.25 -21.68 ;
      RECT 79.15 -20.31 79.25 -19.775 ;
      RECT 79.15 -18.985 79.25 -18.45 ;
      RECT 79.15 -17.08 79.25 -16.545 ;
      RECT 79.15 -15.755 79.25 -15.22 ;
      RECT 79.15 -13.85 79.25 -13.315 ;
      RECT 79.15 -12.525 79.25 -11.99 ;
      RECT 79.15 -10.62 79.25 -10.085 ;
      RECT 79.15 -9.295 79.25 -8.76 ;
      RECT 79.15 -7.39 79.25 -6.855 ;
      RECT 79.15 -6.065 79.25 -5.53 ;
      RECT 79.15 -4.16 79.25 -3.625 ;
      RECT 79.15 -2.835 79.25 -2.3 ;
      RECT 79.15 -0.93 79.25 -0.395 ;
      RECT 79.15 0.395 79.25 0.93 ;
      RECT 79.025 -108.175 79.125 -107.215 ;
      RECT 78.65 -100.19 79 -100.07 ;
      RECT 78.65 -96.96 79 -96.84 ;
      RECT 78.65 -93.73 79 -93.61 ;
      RECT 78.65 -90.5 79 -90.38 ;
      RECT 78.65 -87.27 79 -87.15 ;
      RECT 78.65 -84.04 79 -83.92 ;
      RECT 78.65 -80.81 79 -80.69 ;
      RECT 78.65 -77.58 79 -77.46 ;
      RECT 78.65 -74.35 79 -74.23 ;
      RECT 78.65 -71.12 79 -71 ;
      RECT 78.65 -67.89 79 -67.77 ;
      RECT 78.65 -64.66 79 -64.54 ;
      RECT 78.65 -61.43 79 -61.31 ;
      RECT 78.65 -58.2 79 -58.08 ;
      RECT 78.65 -54.97 79 -54.85 ;
      RECT 78.65 -51.74 79 -51.62 ;
      RECT 78.65 -48.51 79 -48.39 ;
      RECT 78.65 -45.28 79 -45.16 ;
      RECT 78.65 -42.05 79 -41.93 ;
      RECT 78.65 -38.82 79 -38.7 ;
      RECT 78.65 -35.59 79 -35.47 ;
      RECT 78.65 -32.36 79 -32.24 ;
      RECT 78.65 -29.13 79 -29.01 ;
      RECT 78.65 -25.9 79 -25.78 ;
      RECT 78.65 -22.67 79 -22.55 ;
      RECT 78.65 -19.44 79 -19.32 ;
      RECT 78.65 -16.21 79 -16.09 ;
      RECT 78.65 -12.98 79 -12.86 ;
      RECT 78.65 -9.75 79 -9.63 ;
      RECT 78.65 -6.52 79 -6.4 ;
      RECT 78.65 -3.29 79 -3.17 ;
      RECT 78.65 -0.06 79 0.06 ;
      RECT 78.855 -112.255 78.955 -111.775 ;
      RECT 78.855 -110.765 78.955 -110.295 ;
      RECT 78.765 -108.175 78.865 -107.215 ;
      RECT 78.765 2.175 78.865 3.135 ;
      RECT 78.165 -100.19 78.515 -100.07 ;
      RECT 78.165 -96.96 78.515 -96.84 ;
      RECT 78.165 -93.73 78.515 -93.61 ;
      RECT 78.165 -90.5 78.515 -90.38 ;
      RECT 78.165 -87.27 78.515 -87.15 ;
      RECT 78.165 -84.04 78.515 -83.92 ;
      RECT 78.165 -80.81 78.515 -80.69 ;
      RECT 78.165 -77.58 78.515 -77.46 ;
      RECT 78.165 -74.35 78.515 -74.23 ;
      RECT 78.165 -71.12 78.515 -71 ;
      RECT 78.165 -67.89 78.515 -67.77 ;
      RECT 78.165 -64.66 78.515 -64.54 ;
      RECT 78.165 -61.43 78.515 -61.31 ;
      RECT 78.165 -58.2 78.515 -58.08 ;
      RECT 78.165 -54.97 78.515 -54.85 ;
      RECT 78.165 -51.74 78.515 -51.62 ;
      RECT 78.165 -48.51 78.515 -48.39 ;
      RECT 78.165 -45.28 78.515 -45.16 ;
      RECT 78.165 -42.05 78.515 -41.93 ;
      RECT 78.165 -38.82 78.515 -38.7 ;
      RECT 78.165 -35.59 78.515 -35.47 ;
      RECT 78.165 -32.36 78.515 -32.24 ;
      RECT 78.165 -29.13 78.515 -29.01 ;
      RECT 78.165 -25.9 78.515 -25.78 ;
      RECT 78.165 -22.67 78.515 -22.55 ;
      RECT 78.165 -19.44 78.515 -19.32 ;
      RECT 78.165 -16.21 78.515 -16.09 ;
      RECT 78.165 -12.98 78.515 -12.86 ;
      RECT 78.165 -9.75 78.515 -9.63 ;
      RECT 78.165 -6.52 78.515 -6.4 ;
      RECT 78.165 -3.29 78.515 -3.17 ;
      RECT 78.165 -0.06 78.515 0.06 ;
      RECT 78.335 -108.175 78.435 -107.215 ;
      RECT 78.335 2.175 78.435 3.135 ;
      RECT 78.23 -110.765 78.4 -110.385 ;
      RECT 78.265 -112.245 78.365 -111.775 ;
      RECT 78.075 -108.175 78.175 -107.215 ;
      RECT 77.95 -101.06 78.05 -100.525 ;
      RECT 77.95 -99.735 78.05 -99.2 ;
      RECT 77.95 -97.83 78.05 -97.295 ;
      RECT 77.95 -96.505 78.05 -95.97 ;
      RECT 77.95 -94.6 78.05 -94.065 ;
      RECT 77.95 -93.275 78.05 -92.74 ;
      RECT 77.95 -91.37 78.05 -90.835 ;
      RECT 77.95 -90.045 78.05 -89.51 ;
      RECT 77.95 -88.14 78.05 -87.605 ;
      RECT 77.95 -86.815 78.05 -86.28 ;
      RECT 77.95 -84.91 78.05 -84.375 ;
      RECT 77.95 -83.585 78.05 -83.05 ;
      RECT 77.95 -81.68 78.05 -81.145 ;
      RECT 77.95 -80.355 78.05 -79.82 ;
      RECT 77.95 -78.45 78.05 -77.915 ;
      RECT 77.95 -77.125 78.05 -76.59 ;
      RECT 77.95 -75.22 78.05 -74.685 ;
      RECT 77.95 -73.895 78.05 -73.36 ;
      RECT 77.95 -71.99 78.05 -71.455 ;
      RECT 77.95 -70.665 78.05 -70.13 ;
      RECT 77.95 -68.76 78.05 -68.225 ;
      RECT 77.95 -67.435 78.05 -66.9 ;
      RECT 77.95 -65.53 78.05 -64.995 ;
      RECT 77.95 -64.205 78.05 -63.67 ;
      RECT 77.95 -62.3 78.05 -61.765 ;
      RECT 77.95 -60.975 78.05 -60.44 ;
      RECT 77.95 -59.07 78.05 -58.535 ;
      RECT 77.95 -57.745 78.05 -57.21 ;
      RECT 77.95 -55.84 78.05 -55.305 ;
      RECT 77.95 -54.515 78.05 -53.98 ;
      RECT 77.95 -52.61 78.05 -52.075 ;
      RECT 77.95 -51.285 78.05 -50.75 ;
      RECT 77.95 -49.38 78.05 -48.845 ;
      RECT 77.95 -48.055 78.05 -47.52 ;
      RECT 77.95 -46.15 78.05 -45.615 ;
      RECT 77.95 -44.825 78.05 -44.29 ;
      RECT 77.95 -42.92 78.05 -42.385 ;
      RECT 77.95 -41.595 78.05 -41.06 ;
      RECT 77.95 -39.69 78.05 -39.155 ;
      RECT 77.95 -38.365 78.05 -37.83 ;
      RECT 77.95 -36.46 78.05 -35.925 ;
      RECT 77.95 -35.135 78.05 -34.6 ;
      RECT 77.95 -33.23 78.05 -32.695 ;
      RECT 77.95 -31.905 78.05 -31.37 ;
      RECT 77.95 -30 78.05 -29.465 ;
      RECT 77.95 -28.675 78.05 -28.14 ;
      RECT 77.95 -26.77 78.05 -26.235 ;
      RECT 77.95 -25.445 78.05 -24.91 ;
      RECT 77.95 -23.54 78.05 -23.005 ;
      RECT 77.95 -22.215 78.05 -21.68 ;
      RECT 77.95 -20.31 78.05 -19.775 ;
      RECT 77.95 -18.985 78.05 -18.45 ;
      RECT 77.95 -17.08 78.05 -16.545 ;
      RECT 77.95 -15.755 78.05 -15.22 ;
      RECT 77.95 -13.85 78.05 -13.315 ;
      RECT 77.95 -12.525 78.05 -11.99 ;
      RECT 77.95 -10.62 78.05 -10.085 ;
      RECT 77.95 -9.295 78.05 -8.76 ;
      RECT 77.95 -7.39 78.05 -6.855 ;
      RECT 77.95 -6.065 78.05 -5.53 ;
      RECT 77.95 -4.16 78.05 -3.625 ;
      RECT 77.95 -2.835 78.05 -2.3 ;
      RECT 77.95 -0.93 78.05 -0.395 ;
      RECT 77.95 0.395 78.05 0.93 ;
      RECT 77.825 -108.175 77.925 -107.215 ;
      RECT 77.45 -100.19 77.8 -100.07 ;
      RECT 77.45 -96.96 77.8 -96.84 ;
      RECT 77.45 -93.73 77.8 -93.61 ;
      RECT 77.45 -90.5 77.8 -90.38 ;
      RECT 77.45 -87.27 77.8 -87.15 ;
      RECT 77.45 -84.04 77.8 -83.92 ;
      RECT 77.45 -80.81 77.8 -80.69 ;
      RECT 77.45 -77.58 77.8 -77.46 ;
      RECT 77.45 -74.35 77.8 -74.23 ;
      RECT 77.45 -71.12 77.8 -71 ;
      RECT 77.45 -67.89 77.8 -67.77 ;
      RECT 77.45 -64.66 77.8 -64.54 ;
      RECT 77.45 -61.43 77.8 -61.31 ;
      RECT 77.45 -58.2 77.8 -58.08 ;
      RECT 77.45 -54.97 77.8 -54.85 ;
      RECT 77.45 -51.74 77.8 -51.62 ;
      RECT 77.45 -48.51 77.8 -48.39 ;
      RECT 77.45 -45.28 77.8 -45.16 ;
      RECT 77.45 -42.05 77.8 -41.93 ;
      RECT 77.45 -38.82 77.8 -38.7 ;
      RECT 77.45 -35.59 77.8 -35.47 ;
      RECT 77.45 -32.36 77.8 -32.24 ;
      RECT 77.45 -29.13 77.8 -29.01 ;
      RECT 77.45 -25.9 77.8 -25.78 ;
      RECT 77.45 -22.67 77.8 -22.55 ;
      RECT 77.45 -19.44 77.8 -19.32 ;
      RECT 77.45 -16.21 77.8 -16.09 ;
      RECT 77.45 -12.98 77.8 -12.86 ;
      RECT 77.45 -9.75 77.8 -9.63 ;
      RECT 77.45 -6.52 77.8 -6.4 ;
      RECT 77.45 -3.29 77.8 -3.17 ;
      RECT 77.45 -0.06 77.8 0.06 ;
      RECT 77.565 -108.175 77.665 -107.215 ;
      RECT 77.565 2.175 77.665 3.135 ;
      RECT 77.465 -113.555 77.565 -113.085 ;
      RECT 76.965 -100.19 77.315 -100.07 ;
      RECT 76.965 -96.96 77.315 -96.84 ;
      RECT 76.965 -93.73 77.315 -93.61 ;
      RECT 76.965 -90.5 77.315 -90.38 ;
      RECT 76.965 -87.27 77.315 -87.15 ;
      RECT 76.965 -84.04 77.315 -83.92 ;
      RECT 76.965 -80.81 77.315 -80.69 ;
      RECT 76.965 -77.58 77.315 -77.46 ;
      RECT 76.965 -74.35 77.315 -74.23 ;
      RECT 76.965 -71.12 77.315 -71 ;
      RECT 76.965 -67.89 77.315 -67.77 ;
      RECT 76.965 -64.66 77.315 -64.54 ;
      RECT 76.965 -61.43 77.315 -61.31 ;
      RECT 76.965 -58.2 77.315 -58.08 ;
      RECT 76.965 -54.97 77.315 -54.85 ;
      RECT 76.965 -51.74 77.315 -51.62 ;
      RECT 76.965 -48.51 77.315 -48.39 ;
      RECT 76.965 -45.28 77.315 -45.16 ;
      RECT 76.965 -42.05 77.315 -41.93 ;
      RECT 76.965 -38.82 77.315 -38.7 ;
      RECT 76.965 -35.59 77.315 -35.47 ;
      RECT 76.965 -32.36 77.315 -32.24 ;
      RECT 76.965 -29.13 77.315 -29.01 ;
      RECT 76.965 -25.9 77.315 -25.78 ;
      RECT 76.965 -22.67 77.315 -22.55 ;
      RECT 76.965 -19.44 77.315 -19.32 ;
      RECT 76.965 -16.21 77.315 -16.09 ;
      RECT 76.965 -12.98 77.315 -12.86 ;
      RECT 76.965 -9.75 77.315 -9.63 ;
      RECT 76.965 -6.52 77.315 -6.4 ;
      RECT 76.965 -3.29 77.315 -3.17 ;
      RECT 76.965 -0.06 77.315 0.06 ;
      RECT 77.1 -110.735 77.25 -110.445 ;
      RECT 77.135 -108.175 77.235 -107.215 ;
      RECT 77.135 2.175 77.235 3.135 ;
      RECT 77.115 -112.19 77.215 -111.65 ;
      RECT 76.875 -113.555 76.975 -113.085 ;
      RECT 76.875 -108.175 76.975 -107.215 ;
      RECT 76.75 -101.06 76.85 -100.525 ;
      RECT 76.75 -99.735 76.85 -99.2 ;
      RECT 76.75 -97.83 76.85 -97.295 ;
      RECT 76.75 -96.505 76.85 -95.97 ;
      RECT 76.75 -94.6 76.85 -94.065 ;
      RECT 76.75 -93.275 76.85 -92.74 ;
      RECT 76.75 -91.37 76.85 -90.835 ;
      RECT 76.75 -90.045 76.85 -89.51 ;
      RECT 76.75 -88.14 76.85 -87.605 ;
      RECT 76.75 -86.815 76.85 -86.28 ;
      RECT 76.75 -84.91 76.85 -84.375 ;
      RECT 76.75 -83.585 76.85 -83.05 ;
      RECT 76.75 -81.68 76.85 -81.145 ;
      RECT 76.75 -80.355 76.85 -79.82 ;
      RECT 76.75 -78.45 76.85 -77.915 ;
      RECT 76.75 -77.125 76.85 -76.59 ;
      RECT 76.75 -75.22 76.85 -74.685 ;
      RECT 76.75 -73.895 76.85 -73.36 ;
      RECT 76.75 -71.99 76.85 -71.455 ;
      RECT 76.75 -70.665 76.85 -70.13 ;
      RECT 76.75 -68.76 76.85 -68.225 ;
      RECT 76.75 -67.435 76.85 -66.9 ;
      RECT 76.75 -65.53 76.85 -64.995 ;
      RECT 76.75 -64.205 76.85 -63.67 ;
      RECT 76.75 -62.3 76.85 -61.765 ;
      RECT 76.75 -60.975 76.85 -60.44 ;
      RECT 76.75 -59.07 76.85 -58.535 ;
      RECT 76.75 -57.745 76.85 -57.21 ;
      RECT 76.75 -55.84 76.85 -55.305 ;
      RECT 76.75 -54.515 76.85 -53.98 ;
      RECT 76.75 -52.61 76.85 -52.075 ;
      RECT 76.75 -51.285 76.85 -50.75 ;
      RECT 76.75 -49.38 76.85 -48.845 ;
      RECT 76.75 -48.055 76.85 -47.52 ;
      RECT 76.75 -46.15 76.85 -45.615 ;
      RECT 76.75 -44.825 76.85 -44.29 ;
      RECT 76.75 -42.92 76.85 -42.385 ;
      RECT 76.75 -41.595 76.85 -41.06 ;
      RECT 76.75 -39.69 76.85 -39.155 ;
      RECT 76.75 -38.365 76.85 -37.83 ;
      RECT 76.75 -36.46 76.85 -35.925 ;
      RECT 76.75 -35.135 76.85 -34.6 ;
      RECT 76.75 -33.23 76.85 -32.695 ;
      RECT 76.75 -31.905 76.85 -31.37 ;
      RECT 76.75 -30 76.85 -29.465 ;
      RECT 76.75 -28.675 76.85 -28.14 ;
      RECT 76.75 -26.77 76.85 -26.235 ;
      RECT 76.75 -25.445 76.85 -24.91 ;
      RECT 76.75 -23.54 76.85 -23.005 ;
      RECT 76.75 -22.215 76.85 -21.68 ;
      RECT 76.75 -20.31 76.85 -19.775 ;
      RECT 76.75 -18.985 76.85 -18.45 ;
      RECT 76.75 -17.08 76.85 -16.545 ;
      RECT 76.75 -15.755 76.85 -15.22 ;
      RECT 76.75 -13.85 76.85 -13.315 ;
      RECT 76.75 -12.525 76.85 -11.99 ;
      RECT 76.75 -10.62 76.85 -10.085 ;
      RECT 76.75 -9.295 76.85 -8.76 ;
      RECT 76.75 -7.39 76.85 -6.855 ;
      RECT 76.75 -6.065 76.85 -5.53 ;
      RECT 76.75 -4.16 76.85 -3.625 ;
      RECT 76.75 -2.835 76.85 -2.3 ;
      RECT 76.75 -0.93 76.85 -0.395 ;
      RECT 76.75 0.395 76.85 0.93 ;
      RECT 76.625 -104.945 76.725 -103.985 ;
      RECT 76.25 -100.19 76.6 -100.07 ;
      RECT 76.25 -96.96 76.6 -96.84 ;
      RECT 76.25 -93.73 76.6 -93.61 ;
      RECT 76.25 -90.5 76.6 -90.38 ;
      RECT 76.25 -87.27 76.6 -87.15 ;
      RECT 76.25 -84.04 76.6 -83.92 ;
      RECT 76.25 -80.81 76.6 -80.69 ;
      RECT 76.25 -77.58 76.6 -77.46 ;
      RECT 76.25 -74.35 76.6 -74.23 ;
      RECT 76.25 -71.12 76.6 -71 ;
      RECT 76.25 -67.89 76.6 -67.77 ;
      RECT 76.25 -64.66 76.6 -64.54 ;
      RECT 76.25 -61.43 76.6 -61.31 ;
      RECT 76.25 -58.2 76.6 -58.08 ;
      RECT 76.25 -54.97 76.6 -54.85 ;
      RECT 76.25 -51.74 76.6 -51.62 ;
      RECT 76.25 -48.51 76.6 -48.39 ;
      RECT 76.25 -45.28 76.6 -45.16 ;
      RECT 76.25 -42.05 76.6 -41.93 ;
      RECT 76.25 -38.82 76.6 -38.7 ;
      RECT 76.25 -35.59 76.6 -35.47 ;
      RECT 76.25 -32.36 76.6 -32.24 ;
      RECT 76.25 -29.13 76.6 -29.01 ;
      RECT 76.25 -25.9 76.6 -25.78 ;
      RECT 76.25 -22.67 76.6 -22.55 ;
      RECT 76.25 -19.44 76.6 -19.32 ;
      RECT 76.25 -16.21 76.6 -16.09 ;
      RECT 76.25 -12.98 76.6 -12.86 ;
      RECT 76.25 -9.75 76.6 -9.63 ;
      RECT 76.25 -6.52 76.6 -6.4 ;
      RECT 76.25 -3.29 76.6 -3.17 ;
      RECT 76.25 -0.06 76.6 0.06 ;
      RECT 76.365 -104.945 76.465 -103.985 ;
      RECT 76.365 2.175 76.465 3.135 ;
      RECT 76.075 -112.255 76.175 -111.775 ;
      RECT 76.075 -110.765 76.175 -110.295 ;
      RECT 75.765 -100.19 76.115 -100.07 ;
      RECT 75.765 -96.96 76.115 -96.84 ;
      RECT 75.765 -93.73 76.115 -93.61 ;
      RECT 75.765 -90.5 76.115 -90.38 ;
      RECT 75.765 -87.27 76.115 -87.15 ;
      RECT 75.765 -84.04 76.115 -83.92 ;
      RECT 75.765 -80.81 76.115 -80.69 ;
      RECT 75.765 -77.58 76.115 -77.46 ;
      RECT 75.765 -74.35 76.115 -74.23 ;
      RECT 75.765 -71.12 76.115 -71 ;
      RECT 75.765 -67.89 76.115 -67.77 ;
      RECT 75.765 -64.66 76.115 -64.54 ;
      RECT 75.765 -61.43 76.115 -61.31 ;
      RECT 75.765 -58.2 76.115 -58.08 ;
      RECT 75.765 -54.97 76.115 -54.85 ;
      RECT 75.765 -51.74 76.115 -51.62 ;
      RECT 75.765 -48.51 76.115 -48.39 ;
      RECT 75.765 -45.28 76.115 -45.16 ;
      RECT 75.765 -42.05 76.115 -41.93 ;
      RECT 75.765 -38.82 76.115 -38.7 ;
      RECT 75.765 -35.59 76.115 -35.47 ;
      RECT 75.765 -32.36 76.115 -32.24 ;
      RECT 75.765 -29.13 76.115 -29.01 ;
      RECT 75.765 -25.9 76.115 -25.78 ;
      RECT 75.765 -22.67 76.115 -22.55 ;
      RECT 75.765 -19.44 76.115 -19.32 ;
      RECT 75.765 -16.21 76.115 -16.09 ;
      RECT 75.765 -12.98 76.115 -12.86 ;
      RECT 75.765 -9.75 76.115 -9.63 ;
      RECT 75.765 -6.52 76.115 -6.4 ;
      RECT 75.765 -3.29 76.115 -3.17 ;
      RECT 75.765 -0.06 76.115 0.06 ;
      RECT 75.935 -104.945 76.035 -103.985 ;
      RECT 75.935 2.175 76.035 3.135 ;
      RECT 72.035 -108.655 75.815 -108.535 ;
      RECT 75.675 -104.945 75.775 -103.985 ;
      RECT 75.55 -101.06 75.65 -100.525 ;
      RECT 75.55 -99.735 75.65 -99.2 ;
      RECT 75.55 -97.83 75.65 -97.295 ;
      RECT 75.55 -96.505 75.65 -95.97 ;
      RECT 75.55 -94.6 75.65 -94.065 ;
      RECT 75.55 -93.275 75.65 -92.74 ;
      RECT 75.55 -91.37 75.65 -90.835 ;
      RECT 75.55 -90.045 75.65 -89.51 ;
      RECT 75.55 -88.14 75.65 -87.605 ;
      RECT 75.55 -86.815 75.65 -86.28 ;
      RECT 75.55 -84.91 75.65 -84.375 ;
      RECT 75.55 -83.585 75.65 -83.05 ;
      RECT 75.55 -81.68 75.65 -81.145 ;
      RECT 75.55 -80.355 75.65 -79.82 ;
      RECT 75.55 -78.45 75.65 -77.915 ;
      RECT 75.55 -77.125 75.65 -76.59 ;
      RECT 75.55 -75.22 75.65 -74.685 ;
      RECT 75.55 -73.895 75.65 -73.36 ;
      RECT 75.55 -71.99 75.65 -71.455 ;
      RECT 75.55 -70.665 75.65 -70.13 ;
      RECT 75.55 -68.76 75.65 -68.225 ;
      RECT 75.55 -67.435 75.65 -66.9 ;
      RECT 75.55 -65.53 75.65 -64.995 ;
      RECT 75.55 -64.205 75.65 -63.67 ;
      RECT 75.55 -62.3 75.65 -61.765 ;
      RECT 75.55 -60.975 75.65 -60.44 ;
      RECT 75.55 -59.07 75.65 -58.535 ;
      RECT 75.55 -57.745 75.65 -57.21 ;
      RECT 75.55 -55.84 75.65 -55.305 ;
      RECT 75.55 -54.515 75.65 -53.98 ;
      RECT 75.55 -52.61 75.65 -52.075 ;
      RECT 75.55 -51.285 75.65 -50.75 ;
      RECT 75.55 -49.38 75.65 -48.845 ;
      RECT 75.55 -48.055 75.65 -47.52 ;
      RECT 75.55 -46.15 75.65 -45.615 ;
      RECT 75.55 -44.825 75.65 -44.29 ;
      RECT 75.55 -42.92 75.65 -42.385 ;
      RECT 75.55 -41.595 75.65 -41.06 ;
      RECT 75.55 -39.69 75.65 -39.155 ;
      RECT 75.55 -38.365 75.65 -37.83 ;
      RECT 75.55 -36.46 75.65 -35.925 ;
      RECT 75.55 -35.135 75.65 -34.6 ;
      RECT 75.55 -33.23 75.65 -32.695 ;
      RECT 75.55 -31.905 75.65 -31.37 ;
      RECT 75.55 -30 75.65 -29.465 ;
      RECT 75.55 -28.675 75.65 -28.14 ;
      RECT 75.55 -26.77 75.65 -26.235 ;
      RECT 75.55 -25.445 75.65 -24.91 ;
      RECT 75.55 -23.54 75.65 -23.005 ;
      RECT 75.55 -22.215 75.65 -21.68 ;
      RECT 75.55 -20.31 75.65 -19.775 ;
      RECT 75.55 -18.985 75.65 -18.45 ;
      RECT 75.55 -17.08 75.65 -16.545 ;
      RECT 75.55 -15.755 75.65 -15.22 ;
      RECT 75.55 -13.85 75.65 -13.315 ;
      RECT 75.55 -12.525 75.65 -11.99 ;
      RECT 75.55 -10.62 75.65 -10.085 ;
      RECT 75.55 -9.295 75.65 -8.76 ;
      RECT 75.55 -7.39 75.65 -6.855 ;
      RECT 75.55 -6.065 75.65 -5.53 ;
      RECT 75.55 -4.16 75.65 -3.625 ;
      RECT 75.55 -2.835 75.65 -2.3 ;
      RECT 75.55 -0.93 75.65 -0.395 ;
      RECT 75.55 0.395 75.65 0.93 ;
      RECT 75.485 -110.75 75.605 -110.37 ;
      RECT 75.485 -112.245 75.585 -111.775 ;
      RECT 75.425 -104.945 75.525 -103.985 ;
      RECT 75.05 -100.19 75.4 -100.07 ;
      RECT 75.05 -96.96 75.4 -96.84 ;
      RECT 75.05 -93.73 75.4 -93.61 ;
      RECT 75.05 -90.5 75.4 -90.38 ;
      RECT 75.05 -87.27 75.4 -87.15 ;
      RECT 75.05 -84.04 75.4 -83.92 ;
      RECT 75.05 -80.81 75.4 -80.69 ;
      RECT 75.05 -77.58 75.4 -77.46 ;
      RECT 75.05 -74.35 75.4 -74.23 ;
      RECT 75.05 -71.12 75.4 -71 ;
      RECT 75.05 -67.89 75.4 -67.77 ;
      RECT 75.05 -64.66 75.4 -64.54 ;
      RECT 75.05 -61.43 75.4 -61.31 ;
      RECT 75.05 -58.2 75.4 -58.08 ;
      RECT 75.05 -54.97 75.4 -54.85 ;
      RECT 75.05 -51.74 75.4 -51.62 ;
      RECT 75.05 -48.51 75.4 -48.39 ;
      RECT 75.05 -45.28 75.4 -45.16 ;
      RECT 75.05 -42.05 75.4 -41.93 ;
      RECT 75.05 -38.82 75.4 -38.7 ;
      RECT 75.05 -35.59 75.4 -35.47 ;
      RECT 75.05 -32.36 75.4 -32.24 ;
      RECT 75.05 -29.13 75.4 -29.01 ;
      RECT 75.05 -25.9 75.4 -25.78 ;
      RECT 75.05 -22.67 75.4 -22.55 ;
      RECT 75.05 -19.44 75.4 -19.32 ;
      RECT 75.05 -16.21 75.4 -16.09 ;
      RECT 75.05 -12.98 75.4 -12.86 ;
      RECT 75.05 -9.75 75.4 -9.63 ;
      RECT 75.05 -6.52 75.4 -6.4 ;
      RECT 75.05 -3.29 75.4 -3.17 ;
      RECT 75.05 -0.06 75.4 0.06 ;
      RECT 75.165 -104.945 75.265 -103.985 ;
      RECT 75.165 2.175 75.265 3.135 ;
      RECT 74.895 -109.595 75.03 -109.275 ;
      RECT 74.565 -100.19 74.915 -100.07 ;
      RECT 74.565 -96.96 74.915 -96.84 ;
      RECT 74.565 -93.73 74.915 -93.61 ;
      RECT 74.565 -90.5 74.915 -90.38 ;
      RECT 74.565 -87.27 74.915 -87.15 ;
      RECT 74.565 -84.04 74.915 -83.92 ;
      RECT 74.565 -80.81 74.915 -80.69 ;
      RECT 74.565 -77.58 74.915 -77.46 ;
      RECT 74.565 -74.35 74.915 -74.23 ;
      RECT 74.565 -71.12 74.915 -71 ;
      RECT 74.565 -67.89 74.915 -67.77 ;
      RECT 74.565 -64.66 74.915 -64.54 ;
      RECT 74.565 -61.43 74.915 -61.31 ;
      RECT 74.565 -58.2 74.915 -58.08 ;
      RECT 74.565 -54.97 74.915 -54.85 ;
      RECT 74.565 -51.74 74.915 -51.62 ;
      RECT 74.565 -48.51 74.915 -48.39 ;
      RECT 74.565 -45.28 74.915 -45.16 ;
      RECT 74.565 -42.05 74.915 -41.93 ;
      RECT 74.565 -38.82 74.915 -38.7 ;
      RECT 74.565 -35.59 74.915 -35.47 ;
      RECT 74.565 -32.36 74.915 -32.24 ;
      RECT 74.565 -29.13 74.915 -29.01 ;
      RECT 74.565 -25.9 74.915 -25.78 ;
      RECT 74.565 -22.67 74.915 -22.55 ;
      RECT 74.565 -19.44 74.915 -19.32 ;
      RECT 74.565 -16.21 74.915 -16.09 ;
      RECT 74.565 -12.98 74.915 -12.86 ;
      RECT 74.565 -9.75 74.915 -9.63 ;
      RECT 74.565 -6.52 74.915 -6.4 ;
      RECT 74.565 -3.29 74.915 -3.17 ;
      RECT 74.565 -0.06 74.915 0.06 ;
      RECT 74.735 -104.945 74.835 -103.985 ;
      RECT 74.735 2.175 74.835 3.135 ;
      RECT 74.56 -109.595 74.705 -109.275 ;
      RECT 74.475 -104.945 74.575 -103.985 ;
      RECT 74.35 -101.06 74.45 -100.525 ;
      RECT 74.35 -99.735 74.45 -99.2 ;
      RECT 74.35 -97.83 74.45 -97.295 ;
      RECT 74.35 -96.505 74.45 -95.97 ;
      RECT 74.35 -94.6 74.45 -94.065 ;
      RECT 74.35 -93.275 74.45 -92.74 ;
      RECT 74.35 -91.37 74.45 -90.835 ;
      RECT 74.35 -90.045 74.45 -89.51 ;
      RECT 74.35 -88.14 74.45 -87.605 ;
      RECT 74.35 -86.815 74.45 -86.28 ;
      RECT 74.35 -84.91 74.45 -84.375 ;
      RECT 74.35 -83.585 74.45 -83.05 ;
      RECT 74.35 -81.68 74.45 -81.145 ;
      RECT 74.35 -80.355 74.45 -79.82 ;
      RECT 74.35 -78.45 74.45 -77.915 ;
      RECT 74.35 -77.125 74.45 -76.59 ;
      RECT 74.35 -75.22 74.45 -74.685 ;
      RECT 74.35 -73.895 74.45 -73.36 ;
      RECT 74.35 -71.99 74.45 -71.455 ;
      RECT 74.35 -70.665 74.45 -70.13 ;
      RECT 74.35 -68.76 74.45 -68.225 ;
      RECT 74.35 -67.435 74.45 -66.9 ;
      RECT 74.35 -65.53 74.45 -64.995 ;
      RECT 74.35 -64.205 74.45 -63.67 ;
      RECT 74.35 -62.3 74.45 -61.765 ;
      RECT 74.35 -60.975 74.45 -60.44 ;
      RECT 74.35 -59.07 74.45 -58.535 ;
      RECT 74.35 -57.745 74.45 -57.21 ;
      RECT 74.35 -55.84 74.45 -55.305 ;
      RECT 74.35 -54.515 74.45 -53.98 ;
      RECT 74.35 -52.61 74.45 -52.075 ;
      RECT 74.35 -51.285 74.45 -50.75 ;
      RECT 74.35 -49.38 74.45 -48.845 ;
      RECT 74.35 -48.055 74.45 -47.52 ;
      RECT 74.35 -46.15 74.45 -45.615 ;
      RECT 74.35 -44.825 74.45 -44.29 ;
      RECT 74.35 -42.92 74.45 -42.385 ;
      RECT 74.35 -41.595 74.45 -41.06 ;
      RECT 74.35 -39.69 74.45 -39.155 ;
      RECT 74.35 -38.365 74.45 -37.83 ;
      RECT 74.35 -36.46 74.45 -35.925 ;
      RECT 74.35 -35.135 74.45 -34.6 ;
      RECT 74.35 -33.23 74.45 -32.695 ;
      RECT 74.35 -31.905 74.45 -31.37 ;
      RECT 74.35 -30 74.45 -29.465 ;
      RECT 74.35 -28.675 74.45 -28.14 ;
      RECT 74.35 -26.77 74.45 -26.235 ;
      RECT 74.35 -25.445 74.45 -24.91 ;
      RECT 74.35 -23.54 74.45 -23.005 ;
      RECT 74.35 -22.215 74.45 -21.68 ;
      RECT 74.35 -20.31 74.45 -19.775 ;
      RECT 74.35 -18.985 74.45 -18.45 ;
      RECT 74.35 -17.08 74.45 -16.545 ;
      RECT 74.35 -15.755 74.45 -15.22 ;
      RECT 74.35 -13.85 74.45 -13.315 ;
      RECT 74.35 -12.525 74.45 -11.99 ;
      RECT 74.35 -10.62 74.45 -10.085 ;
      RECT 74.35 -9.295 74.45 -8.76 ;
      RECT 74.35 -7.39 74.45 -6.855 ;
      RECT 74.35 -6.065 74.45 -5.53 ;
      RECT 74.35 -4.16 74.45 -3.625 ;
      RECT 74.35 -2.835 74.45 -2.3 ;
      RECT 74.35 -0.93 74.45 -0.395 ;
      RECT 74.35 0.395 74.45 0.93 ;
      RECT 74.225 -108.175 74.325 -107.215 ;
      RECT 73.85 -100.19 74.2 -100.07 ;
      RECT 73.85 -96.96 74.2 -96.84 ;
      RECT 73.85 -93.73 74.2 -93.61 ;
      RECT 73.85 -90.5 74.2 -90.38 ;
      RECT 73.85 -87.27 74.2 -87.15 ;
      RECT 73.85 -84.04 74.2 -83.92 ;
      RECT 73.85 -80.81 74.2 -80.69 ;
      RECT 73.85 -77.58 74.2 -77.46 ;
      RECT 73.85 -74.35 74.2 -74.23 ;
      RECT 73.85 -71.12 74.2 -71 ;
      RECT 73.85 -67.89 74.2 -67.77 ;
      RECT 73.85 -64.66 74.2 -64.54 ;
      RECT 73.85 -61.43 74.2 -61.31 ;
      RECT 73.85 -58.2 74.2 -58.08 ;
      RECT 73.85 -54.97 74.2 -54.85 ;
      RECT 73.85 -51.74 74.2 -51.62 ;
      RECT 73.85 -48.51 74.2 -48.39 ;
      RECT 73.85 -45.28 74.2 -45.16 ;
      RECT 73.85 -42.05 74.2 -41.93 ;
      RECT 73.85 -38.82 74.2 -38.7 ;
      RECT 73.85 -35.59 74.2 -35.47 ;
      RECT 73.85 -32.36 74.2 -32.24 ;
      RECT 73.85 -29.13 74.2 -29.01 ;
      RECT 73.85 -25.9 74.2 -25.78 ;
      RECT 73.85 -22.67 74.2 -22.55 ;
      RECT 73.85 -19.44 74.2 -19.32 ;
      RECT 73.85 -16.21 74.2 -16.09 ;
      RECT 73.85 -12.98 74.2 -12.86 ;
      RECT 73.85 -9.75 74.2 -9.63 ;
      RECT 73.85 -6.52 74.2 -6.4 ;
      RECT 73.85 -3.29 74.2 -3.17 ;
      RECT 73.85 -0.06 74.2 0.06 ;
      RECT 74.055 -112.255 74.155 -111.775 ;
      RECT 74.055 -110.765 74.155 -110.295 ;
      RECT 73.965 -108.175 74.065 -107.215 ;
      RECT 73.965 2.175 74.065 3.135 ;
      RECT 73.365 -100.19 73.715 -100.07 ;
      RECT 73.365 -96.96 73.715 -96.84 ;
      RECT 73.365 -93.73 73.715 -93.61 ;
      RECT 73.365 -90.5 73.715 -90.38 ;
      RECT 73.365 -87.27 73.715 -87.15 ;
      RECT 73.365 -84.04 73.715 -83.92 ;
      RECT 73.365 -80.81 73.715 -80.69 ;
      RECT 73.365 -77.58 73.715 -77.46 ;
      RECT 73.365 -74.35 73.715 -74.23 ;
      RECT 73.365 -71.12 73.715 -71 ;
      RECT 73.365 -67.89 73.715 -67.77 ;
      RECT 73.365 -64.66 73.715 -64.54 ;
      RECT 73.365 -61.43 73.715 -61.31 ;
      RECT 73.365 -58.2 73.715 -58.08 ;
      RECT 73.365 -54.97 73.715 -54.85 ;
      RECT 73.365 -51.74 73.715 -51.62 ;
      RECT 73.365 -48.51 73.715 -48.39 ;
      RECT 73.365 -45.28 73.715 -45.16 ;
      RECT 73.365 -42.05 73.715 -41.93 ;
      RECT 73.365 -38.82 73.715 -38.7 ;
      RECT 73.365 -35.59 73.715 -35.47 ;
      RECT 73.365 -32.36 73.715 -32.24 ;
      RECT 73.365 -29.13 73.715 -29.01 ;
      RECT 73.365 -25.9 73.715 -25.78 ;
      RECT 73.365 -22.67 73.715 -22.55 ;
      RECT 73.365 -19.44 73.715 -19.32 ;
      RECT 73.365 -16.21 73.715 -16.09 ;
      RECT 73.365 -12.98 73.715 -12.86 ;
      RECT 73.365 -9.75 73.715 -9.63 ;
      RECT 73.365 -6.52 73.715 -6.4 ;
      RECT 73.365 -3.29 73.715 -3.17 ;
      RECT 73.365 -0.06 73.715 0.06 ;
      RECT 73.535 -108.175 73.635 -107.215 ;
      RECT 73.535 2.175 73.635 3.135 ;
      RECT 73.43 -110.765 73.6 -110.385 ;
      RECT 73.465 -112.245 73.565 -111.775 ;
      RECT 73.275 -108.175 73.375 -107.215 ;
      RECT 73.15 -101.06 73.25 -100.525 ;
      RECT 73.15 -99.735 73.25 -99.2 ;
      RECT 73.15 -97.83 73.25 -97.295 ;
      RECT 73.15 -96.505 73.25 -95.97 ;
      RECT 73.15 -94.6 73.25 -94.065 ;
      RECT 73.15 -93.275 73.25 -92.74 ;
      RECT 73.15 -91.37 73.25 -90.835 ;
      RECT 73.15 -90.045 73.25 -89.51 ;
      RECT 73.15 -88.14 73.25 -87.605 ;
      RECT 73.15 -86.815 73.25 -86.28 ;
      RECT 73.15 -84.91 73.25 -84.375 ;
      RECT 73.15 -83.585 73.25 -83.05 ;
      RECT 73.15 -81.68 73.25 -81.145 ;
      RECT 73.15 -80.355 73.25 -79.82 ;
      RECT 73.15 -78.45 73.25 -77.915 ;
      RECT 73.15 -77.125 73.25 -76.59 ;
      RECT 73.15 -75.22 73.25 -74.685 ;
      RECT 73.15 -73.895 73.25 -73.36 ;
      RECT 73.15 -71.99 73.25 -71.455 ;
      RECT 73.15 -70.665 73.25 -70.13 ;
      RECT 73.15 -68.76 73.25 -68.225 ;
      RECT 73.15 -67.435 73.25 -66.9 ;
      RECT 73.15 -65.53 73.25 -64.995 ;
      RECT 73.15 -64.205 73.25 -63.67 ;
      RECT 73.15 -62.3 73.25 -61.765 ;
      RECT 73.15 -60.975 73.25 -60.44 ;
      RECT 73.15 -59.07 73.25 -58.535 ;
      RECT 73.15 -57.745 73.25 -57.21 ;
      RECT 73.15 -55.84 73.25 -55.305 ;
      RECT 73.15 -54.515 73.25 -53.98 ;
      RECT 73.15 -52.61 73.25 -52.075 ;
      RECT 73.15 -51.285 73.25 -50.75 ;
      RECT 73.15 -49.38 73.25 -48.845 ;
      RECT 73.15 -48.055 73.25 -47.52 ;
      RECT 73.15 -46.15 73.25 -45.615 ;
      RECT 73.15 -44.825 73.25 -44.29 ;
      RECT 73.15 -42.92 73.25 -42.385 ;
      RECT 73.15 -41.595 73.25 -41.06 ;
      RECT 73.15 -39.69 73.25 -39.155 ;
      RECT 73.15 -38.365 73.25 -37.83 ;
      RECT 73.15 -36.46 73.25 -35.925 ;
      RECT 73.15 -35.135 73.25 -34.6 ;
      RECT 73.15 -33.23 73.25 -32.695 ;
      RECT 73.15 -31.905 73.25 -31.37 ;
      RECT 73.15 -30 73.25 -29.465 ;
      RECT 73.15 -28.675 73.25 -28.14 ;
      RECT 73.15 -26.77 73.25 -26.235 ;
      RECT 73.15 -25.445 73.25 -24.91 ;
      RECT 73.15 -23.54 73.25 -23.005 ;
      RECT 73.15 -22.215 73.25 -21.68 ;
      RECT 73.15 -20.31 73.25 -19.775 ;
      RECT 73.15 -18.985 73.25 -18.45 ;
      RECT 73.15 -17.08 73.25 -16.545 ;
      RECT 73.15 -15.755 73.25 -15.22 ;
      RECT 73.15 -13.85 73.25 -13.315 ;
      RECT 73.15 -12.525 73.25 -11.99 ;
      RECT 73.15 -10.62 73.25 -10.085 ;
      RECT 73.15 -9.295 73.25 -8.76 ;
      RECT 73.15 -7.39 73.25 -6.855 ;
      RECT 73.15 -6.065 73.25 -5.53 ;
      RECT 73.15 -4.16 73.25 -3.625 ;
      RECT 73.15 -2.835 73.25 -2.3 ;
      RECT 73.15 -0.93 73.25 -0.395 ;
      RECT 73.15 0.395 73.25 0.93 ;
      RECT 73.025 -108.175 73.125 -107.215 ;
      RECT 72.65 -100.19 73 -100.07 ;
      RECT 72.65 -96.96 73 -96.84 ;
      RECT 72.65 -93.73 73 -93.61 ;
      RECT 72.65 -90.5 73 -90.38 ;
      RECT 72.65 -87.27 73 -87.15 ;
      RECT 72.65 -84.04 73 -83.92 ;
      RECT 72.65 -80.81 73 -80.69 ;
      RECT 72.65 -77.58 73 -77.46 ;
      RECT 72.65 -74.35 73 -74.23 ;
      RECT 72.65 -71.12 73 -71 ;
      RECT 72.65 -67.89 73 -67.77 ;
      RECT 72.65 -64.66 73 -64.54 ;
      RECT 72.65 -61.43 73 -61.31 ;
      RECT 72.65 -58.2 73 -58.08 ;
      RECT 72.65 -54.97 73 -54.85 ;
      RECT 72.65 -51.74 73 -51.62 ;
      RECT 72.65 -48.51 73 -48.39 ;
      RECT 72.65 -45.28 73 -45.16 ;
      RECT 72.65 -42.05 73 -41.93 ;
      RECT 72.65 -38.82 73 -38.7 ;
      RECT 72.65 -35.59 73 -35.47 ;
      RECT 72.65 -32.36 73 -32.24 ;
      RECT 72.65 -29.13 73 -29.01 ;
      RECT 72.65 -25.9 73 -25.78 ;
      RECT 72.65 -22.67 73 -22.55 ;
      RECT 72.65 -19.44 73 -19.32 ;
      RECT 72.65 -16.21 73 -16.09 ;
      RECT 72.65 -12.98 73 -12.86 ;
      RECT 72.65 -9.75 73 -9.63 ;
      RECT 72.65 -6.52 73 -6.4 ;
      RECT 72.65 -3.29 73 -3.17 ;
      RECT 72.65 -0.06 73 0.06 ;
      RECT 72.765 -108.175 72.865 -107.215 ;
      RECT 72.765 2.175 72.865 3.135 ;
      RECT 72.665 -113.555 72.765 -113.085 ;
      RECT 72.165 -100.19 72.515 -100.07 ;
      RECT 72.165 -96.96 72.515 -96.84 ;
      RECT 72.165 -93.73 72.515 -93.61 ;
      RECT 72.165 -90.5 72.515 -90.38 ;
      RECT 72.165 -87.27 72.515 -87.15 ;
      RECT 72.165 -84.04 72.515 -83.92 ;
      RECT 72.165 -80.81 72.515 -80.69 ;
      RECT 72.165 -77.58 72.515 -77.46 ;
      RECT 72.165 -74.35 72.515 -74.23 ;
      RECT 72.165 -71.12 72.515 -71 ;
      RECT 72.165 -67.89 72.515 -67.77 ;
      RECT 72.165 -64.66 72.515 -64.54 ;
      RECT 72.165 -61.43 72.515 -61.31 ;
      RECT 72.165 -58.2 72.515 -58.08 ;
      RECT 72.165 -54.97 72.515 -54.85 ;
      RECT 72.165 -51.74 72.515 -51.62 ;
      RECT 72.165 -48.51 72.515 -48.39 ;
      RECT 72.165 -45.28 72.515 -45.16 ;
      RECT 72.165 -42.05 72.515 -41.93 ;
      RECT 72.165 -38.82 72.515 -38.7 ;
      RECT 72.165 -35.59 72.515 -35.47 ;
      RECT 72.165 -32.36 72.515 -32.24 ;
      RECT 72.165 -29.13 72.515 -29.01 ;
      RECT 72.165 -25.9 72.515 -25.78 ;
      RECT 72.165 -22.67 72.515 -22.55 ;
      RECT 72.165 -19.44 72.515 -19.32 ;
      RECT 72.165 -16.21 72.515 -16.09 ;
      RECT 72.165 -12.98 72.515 -12.86 ;
      RECT 72.165 -9.75 72.515 -9.63 ;
      RECT 72.165 -6.52 72.515 -6.4 ;
      RECT 72.165 -3.29 72.515 -3.17 ;
      RECT 72.165 -0.06 72.515 0.06 ;
      RECT 72.3 -110.735 72.45 -110.445 ;
      RECT 72.335 -108.175 72.435 -107.215 ;
      RECT 72.335 2.175 72.435 3.135 ;
      RECT 72.315 -112.19 72.415 -111.65 ;
      RECT 72.075 -113.555 72.175 -113.085 ;
      RECT 72.075 -108.175 72.175 -107.215 ;
      RECT 71.95 -101.06 72.05 -100.525 ;
      RECT 71.95 -99.735 72.05 -99.2 ;
      RECT 71.95 -97.83 72.05 -97.295 ;
      RECT 71.95 -96.505 72.05 -95.97 ;
      RECT 71.95 -94.6 72.05 -94.065 ;
      RECT 71.95 -93.275 72.05 -92.74 ;
      RECT 71.95 -91.37 72.05 -90.835 ;
      RECT 71.95 -90.045 72.05 -89.51 ;
      RECT 71.95 -88.14 72.05 -87.605 ;
      RECT 71.95 -86.815 72.05 -86.28 ;
      RECT 71.95 -84.91 72.05 -84.375 ;
      RECT 71.95 -83.585 72.05 -83.05 ;
      RECT 71.95 -81.68 72.05 -81.145 ;
      RECT 71.95 -80.355 72.05 -79.82 ;
      RECT 71.95 -78.45 72.05 -77.915 ;
      RECT 71.95 -77.125 72.05 -76.59 ;
      RECT 71.95 -75.22 72.05 -74.685 ;
      RECT 71.95 -73.895 72.05 -73.36 ;
      RECT 71.95 -71.99 72.05 -71.455 ;
      RECT 71.95 -70.665 72.05 -70.13 ;
      RECT 71.95 -68.76 72.05 -68.225 ;
      RECT 71.95 -67.435 72.05 -66.9 ;
      RECT 71.95 -65.53 72.05 -64.995 ;
      RECT 71.95 -64.205 72.05 -63.67 ;
      RECT 71.95 -62.3 72.05 -61.765 ;
      RECT 71.95 -60.975 72.05 -60.44 ;
      RECT 71.95 -59.07 72.05 -58.535 ;
      RECT 71.95 -57.745 72.05 -57.21 ;
      RECT 71.95 -55.84 72.05 -55.305 ;
      RECT 71.95 -54.515 72.05 -53.98 ;
      RECT 71.95 -52.61 72.05 -52.075 ;
      RECT 71.95 -51.285 72.05 -50.75 ;
      RECT 71.95 -49.38 72.05 -48.845 ;
      RECT 71.95 -48.055 72.05 -47.52 ;
      RECT 71.95 -46.15 72.05 -45.615 ;
      RECT 71.95 -44.825 72.05 -44.29 ;
      RECT 71.95 -42.92 72.05 -42.385 ;
      RECT 71.95 -41.595 72.05 -41.06 ;
      RECT 71.95 -39.69 72.05 -39.155 ;
      RECT 71.95 -38.365 72.05 -37.83 ;
      RECT 71.95 -36.46 72.05 -35.925 ;
      RECT 71.95 -35.135 72.05 -34.6 ;
      RECT 71.95 -33.23 72.05 -32.695 ;
      RECT 71.95 -31.905 72.05 -31.37 ;
      RECT 71.95 -30 72.05 -29.465 ;
      RECT 71.95 -28.675 72.05 -28.14 ;
      RECT 71.95 -26.77 72.05 -26.235 ;
      RECT 71.95 -25.445 72.05 -24.91 ;
      RECT 71.95 -23.54 72.05 -23.005 ;
      RECT 71.95 -22.215 72.05 -21.68 ;
      RECT 71.95 -20.31 72.05 -19.775 ;
      RECT 71.95 -18.985 72.05 -18.45 ;
      RECT 71.95 -17.08 72.05 -16.545 ;
      RECT 71.95 -15.755 72.05 -15.22 ;
      RECT 71.95 -13.85 72.05 -13.315 ;
      RECT 71.95 -12.525 72.05 -11.99 ;
      RECT 71.95 -10.62 72.05 -10.085 ;
      RECT 71.95 -9.295 72.05 -8.76 ;
      RECT 71.95 -7.39 72.05 -6.855 ;
      RECT 71.95 -6.065 72.05 -5.53 ;
      RECT 71.95 -4.16 72.05 -3.625 ;
      RECT 71.95 -2.835 72.05 -2.3 ;
      RECT 71.95 -0.93 72.05 -0.395 ;
      RECT 71.95 0.395 72.05 0.93 ;
      RECT 71.825 -104.945 71.925 -103.985 ;
      RECT 71.45 -100.19 71.8 -100.07 ;
      RECT 71.45 -96.96 71.8 -96.84 ;
      RECT 71.45 -93.73 71.8 -93.61 ;
      RECT 71.45 -90.5 71.8 -90.38 ;
      RECT 71.45 -87.27 71.8 -87.15 ;
      RECT 71.45 -84.04 71.8 -83.92 ;
      RECT 71.45 -80.81 71.8 -80.69 ;
      RECT 71.45 -77.58 71.8 -77.46 ;
      RECT 71.45 -74.35 71.8 -74.23 ;
      RECT 71.45 -71.12 71.8 -71 ;
      RECT 71.45 -67.89 71.8 -67.77 ;
      RECT 71.45 -64.66 71.8 -64.54 ;
      RECT 71.45 -61.43 71.8 -61.31 ;
      RECT 71.45 -58.2 71.8 -58.08 ;
      RECT 71.45 -54.97 71.8 -54.85 ;
      RECT 71.45 -51.74 71.8 -51.62 ;
      RECT 71.45 -48.51 71.8 -48.39 ;
      RECT 71.45 -45.28 71.8 -45.16 ;
      RECT 71.45 -42.05 71.8 -41.93 ;
      RECT 71.45 -38.82 71.8 -38.7 ;
      RECT 71.45 -35.59 71.8 -35.47 ;
      RECT 71.45 -32.36 71.8 -32.24 ;
      RECT 71.45 -29.13 71.8 -29.01 ;
      RECT 71.45 -25.9 71.8 -25.78 ;
      RECT 71.45 -22.67 71.8 -22.55 ;
      RECT 71.45 -19.44 71.8 -19.32 ;
      RECT 71.45 -16.21 71.8 -16.09 ;
      RECT 71.45 -12.98 71.8 -12.86 ;
      RECT 71.45 -9.75 71.8 -9.63 ;
      RECT 71.45 -6.52 71.8 -6.4 ;
      RECT 71.45 -3.29 71.8 -3.17 ;
      RECT 71.45 -0.06 71.8 0.06 ;
      RECT 71.565 -104.945 71.665 -103.985 ;
      RECT 71.565 2.175 71.665 3.135 ;
      RECT 71.275 -112.255 71.375 -111.775 ;
      RECT 71.275 -110.765 71.375 -110.295 ;
      RECT 70.965 -100.19 71.315 -100.07 ;
      RECT 70.965 -96.96 71.315 -96.84 ;
      RECT 70.965 -93.73 71.315 -93.61 ;
      RECT 70.965 -90.5 71.315 -90.38 ;
      RECT 70.965 -87.27 71.315 -87.15 ;
      RECT 70.965 -84.04 71.315 -83.92 ;
      RECT 70.965 -80.81 71.315 -80.69 ;
      RECT 70.965 -77.58 71.315 -77.46 ;
      RECT 70.965 -74.35 71.315 -74.23 ;
      RECT 70.965 -71.12 71.315 -71 ;
      RECT 70.965 -67.89 71.315 -67.77 ;
      RECT 70.965 -64.66 71.315 -64.54 ;
      RECT 70.965 -61.43 71.315 -61.31 ;
      RECT 70.965 -58.2 71.315 -58.08 ;
      RECT 70.965 -54.97 71.315 -54.85 ;
      RECT 70.965 -51.74 71.315 -51.62 ;
      RECT 70.965 -48.51 71.315 -48.39 ;
      RECT 70.965 -45.28 71.315 -45.16 ;
      RECT 70.965 -42.05 71.315 -41.93 ;
      RECT 70.965 -38.82 71.315 -38.7 ;
      RECT 70.965 -35.59 71.315 -35.47 ;
      RECT 70.965 -32.36 71.315 -32.24 ;
      RECT 70.965 -29.13 71.315 -29.01 ;
      RECT 70.965 -25.9 71.315 -25.78 ;
      RECT 70.965 -22.67 71.315 -22.55 ;
      RECT 70.965 -19.44 71.315 -19.32 ;
      RECT 70.965 -16.21 71.315 -16.09 ;
      RECT 70.965 -12.98 71.315 -12.86 ;
      RECT 70.965 -9.75 71.315 -9.63 ;
      RECT 70.965 -6.52 71.315 -6.4 ;
      RECT 70.965 -3.29 71.315 -3.17 ;
      RECT 70.965 -0.06 71.315 0.06 ;
      RECT 71.135 -104.945 71.235 -103.985 ;
      RECT 71.135 2.175 71.235 3.135 ;
      RECT 67.235 -108.655 71.015 -108.535 ;
      RECT 70.875 -104.945 70.975 -103.985 ;
      RECT 70.75 -101.06 70.85 -100.525 ;
      RECT 70.75 -99.735 70.85 -99.2 ;
      RECT 70.75 -97.83 70.85 -97.295 ;
      RECT 70.75 -96.505 70.85 -95.97 ;
      RECT 70.75 -94.6 70.85 -94.065 ;
      RECT 70.75 -93.275 70.85 -92.74 ;
      RECT 70.75 -91.37 70.85 -90.835 ;
      RECT 70.75 -90.045 70.85 -89.51 ;
      RECT 70.75 -88.14 70.85 -87.605 ;
      RECT 70.75 -86.815 70.85 -86.28 ;
      RECT 70.75 -84.91 70.85 -84.375 ;
      RECT 70.75 -83.585 70.85 -83.05 ;
      RECT 70.75 -81.68 70.85 -81.145 ;
      RECT 70.75 -80.355 70.85 -79.82 ;
      RECT 70.75 -78.45 70.85 -77.915 ;
      RECT 70.75 -77.125 70.85 -76.59 ;
      RECT 70.75 -75.22 70.85 -74.685 ;
      RECT 70.75 -73.895 70.85 -73.36 ;
      RECT 70.75 -71.99 70.85 -71.455 ;
      RECT 70.75 -70.665 70.85 -70.13 ;
      RECT 70.75 -68.76 70.85 -68.225 ;
      RECT 70.75 -67.435 70.85 -66.9 ;
      RECT 70.75 -65.53 70.85 -64.995 ;
      RECT 70.75 -64.205 70.85 -63.67 ;
      RECT 70.75 -62.3 70.85 -61.765 ;
      RECT 70.75 -60.975 70.85 -60.44 ;
      RECT 70.75 -59.07 70.85 -58.535 ;
      RECT 70.75 -57.745 70.85 -57.21 ;
      RECT 70.75 -55.84 70.85 -55.305 ;
      RECT 70.75 -54.515 70.85 -53.98 ;
      RECT 70.75 -52.61 70.85 -52.075 ;
      RECT 70.75 -51.285 70.85 -50.75 ;
      RECT 70.75 -49.38 70.85 -48.845 ;
      RECT 70.75 -48.055 70.85 -47.52 ;
      RECT 70.75 -46.15 70.85 -45.615 ;
      RECT 70.75 -44.825 70.85 -44.29 ;
      RECT 70.75 -42.92 70.85 -42.385 ;
      RECT 70.75 -41.595 70.85 -41.06 ;
      RECT 70.75 -39.69 70.85 -39.155 ;
      RECT 70.75 -38.365 70.85 -37.83 ;
      RECT 70.75 -36.46 70.85 -35.925 ;
      RECT 70.75 -35.135 70.85 -34.6 ;
      RECT 70.75 -33.23 70.85 -32.695 ;
      RECT 70.75 -31.905 70.85 -31.37 ;
      RECT 70.75 -30 70.85 -29.465 ;
      RECT 70.75 -28.675 70.85 -28.14 ;
      RECT 70.75 -26.77 70.85 -26.235 ;
      RECT 70.75 -25.445 70.85 -24.91 ;
      RECT 70.75 -23.54 70.85 -23.005 ;
      RECT 70.75 -22.215 70.85 -21.68 ;
      RECT 70.75 -20.31 70.85 -19.775 ;
      RECT 70.75 -18.985 70.85 -18.45 ;
      RECT 70.75 -17.08 70.85 -16.545 ;
      RECT 70.75 -15.755 70.85 -15.22 ;
      RECT 70.75 -13.85 70.85 -13.315 ;
      RECT 70.75 -12.525 70.85 -11.99 ;
      RECT 70.75 -10.62 70.85 -10.085 ;
      RECT 70.75 -9.295 70.85 -8.76 ;
      RECT 70.75 -7.39 70.85 -6.855 ;
      RECT 70.75 -6.065 70.85 -5.53 ;
      RECT 70.75 -4.16 70.85 -3.625 ;
      RECT 70.75 -2.835 70.85 -2.3 ;
      RECT 70.75 -0.93 70.85 -0.395 ;
      RECT 70.75 0.395 70.85 0.93 ;
      RECT 70.685 -110.75 70.805 -110.37 ;
      RECT 70.685 -112.245 70.785 -111.775 ;
      RECT 70.625 -104.945 70.725 -103.985 ;
      RECT 70.25 -100.19 70.6 -100.07 ;
      RECT 70.25 -96.96 70.6 -96.84 ;
      RECT 70.25 -93.73 70.6 -93.61 ;
      RECT 70.25 -90.5 70.6 -90.38 ;
      RECT 70.25 -87.27 70.6 -87.15 ;
      RECT 70.25 -84.04 70.6 -83.92 ;
      RECT 70.25 -80.81 70.6 -80.69 ;
      RECT 70.25 -77.58 70.6 -77.46 ;
      RECT 70.25 -74.35 70.6 -74.23 ;
      RECT 70.25 -71.12 70.6 -71 ;
      RECT 70.25 -67.89 70.6 -67.77 ;
      RECT 70.25 -64.66 70.6 -64.54 ;
      RECT 70.25 -61.43 70.6 -61.31 ;
      RECT 70.25 -58.2 70.6 -58.08 ;
      RECT 70.25 -54.97 70.6 -54.85 ;
      RECT 70.25 -51.74 70.6 -51.62 ;
      RECT 70.25 -48.51 70.6 -48.39 ;
      RECT 70.25 -45.28 70.6 -45.16 ;
      RECT 70.25 -42.05 70.6 -41.93 ;
      RECT 70.25 -38.82 70.6 -38.7 ;
      RECT 70.25 -35.59 70.6 -35.47 ;
      RECT 70.25 -32.36 70.6 -32.24 ;
      RECT 70.25 -29.13 70.6 -29.01 ;
      RECT 70.25 -25.9 70.6 -25.78 ;
      RECT 70.25 -22.67 70.6 -22.55 ;
      RECT 70.25 -19.44 70.6 -19.32 ;
      RECT 70.25 -16.21 70.6 -16.09 ;
      RECT 70.25 -12.98 70.6 -12.86 ;
      RECT 70.25 -9.75 70.6 -9.63 ;
      RECT 70.25 -6.52 70.6 -6.4 ;
      RECT 70.25 -3.29 70.6 -3.17 ;
      RECT 70.25 -0.06 70.6 0.06 ;
      RECT 70.365 -104.945 70.465 -103.985 ;
      RECT 70.365 2.175 70.465 3.135 ;
      RECT 70.095 -109.595 70.23 -109.275 ;
      RECT 69.765 -100.19 70.115 -100.07 ;
      RECT 69.765 -96.96 70.115 -96.84 ;
      RECT 69.765 -93.73 70.115 -93.61 ;
      RECT 69.765 -90.5 70.115 -90.38 ;
      RECT 69.765 -87.27 70.115 -87.15 ;
      RECT 69.765 -84.04 70.115 -83.92 ;
      RECT 69.765 -80.81 70.115 -80.69 ;
      RECT 69.765 -77.58 70.115 -77.46 ;
      RECT 69.765 -74.35 70.115 -74.23 ;
      RECT 69.765 -71.12 70.115 -71 ;
      RECT 69.765 -67.89 70.115 -67.77 ;
      RECT 69.765 -64.66 70.115 -64.54 ;
      RECT 69.765 -61.43 70.115 -61.31 ;
      RECT 69.765 -58.2 70.115 -58.08 ;
      RECT 69.765 -54.97 70.115 -54.85 ;
      RECT 69.765 -51.74 70.115 -51.62 ;
      RECT 69.765 -48.51 70.115 -48.39 ;
      RECT 69.765 -45.28 70.115 -45.16 ;
      RECT 69.765 -42.05 70.115 -41.93 ;
      RECT 69.765 -38.82 70.115 -38.7 ;
      RECT 69.765 -35.59 70.115 -35.47 ;
      RECT 69.765 -32.36 70.115 -32.24 ;
      RECT 69.765 -29.13 70.115 -29.01 ;
      RECT 69.765 -25.9 70.115 -25.78 ;
      RECT 69.765 -22.67 70.115 -22.55 ;
      RECT 69.765 -19.44 70.115 -19.32 ;
      RECT 69.765 -16.21 70.115 -16.09 ;
      RECT 69.765 -12.98 70.115 -12.86 ;
      RECT 69.765 -9.75 70.115 -9.63 ;
      RECT 69.765 -6.52 70.115 -6.4 ;
      RECT 69.765 -3.29 70.115 -3.17 ;
      RECT 69.765 -0.06 70.115 0.06 ;
      RECT 69.935 -104.945 70.035 -103.985 ;
      RECT 69.935 2.175 70.035 3.135 ;
      RECT 69.76 -109.595 69.905 -109.275 ;
      RECT 69.675 -104.945 69.775 -103.985 ;
      RECT 69.55 -101.06 69.65 -100.525 ;
      RECT 69.55 -99.735 69.65 -99.2 ;
      RECT 69.55 -97.83 69.65 -97.295 ;
      RECT 69.55 -96.505 69.65 -95.97 ;
      RECT 69.55 -94.6 69.65 -94.065 ;
      RECT 69.55 -93.275 69.65 -92.74 ;
      RECT 69.55 -91.37 69.65 -90.835 ;
      RECT 69.55 -90.045 69.65 -89.51 ;
      RECT 69.55 -88.14 69.65 -87.605 ;
      RECT 69.55 -86.815 69.65 -86.28 ;
      RECT 69.55 -84.91 69.65 -84.375 ;
      RECT 69.55 -83.585 69.65 -83.05 ;
      RECT 69.55 -81.68 69.65 -81.145 ;
      RECT 69.55 -80.355 69.65 -79.82 ;
      RECT 69.55 -78.45 69.65 -77.915 ;
      RECT 69.55 -77.125 69.65 -76.59 ;
      RECT 69.55 -75.22 69.65 -74.685 ;
      RECT 69.55 -73.895 69.65 -73.36 ;
      RECT 69.55 -71.99 69.65 -71.455 ;
      RECT 69.55 -70.665 69.65 -70.13 ;
      RECT 69.55 -68.76 69.65 -68.225 ;
      RECT 69.55 -67.435 69.65 -66.9 ;
      RECT 69.55 -65.53 69.65 -64.995 ;
      RECT 69.55 -64.205 69.65 -63.67 ;
      RECT 69.55 -62.3 69.65 -61.765 ;
      RECT 69.55 -60.975 69.65 -60.44 ;
      RECT 69.55 -59.07 69.65 -58.535 ;
      RECT 69.55 -57.745 69.65 -57.21 ;
      RECT 69.55 -55.84 69.65 -55.305 ;
      RECT 69.55 -54.515 69.65 -53.98 ;
      RECT 69.55 -52.61 69.65 -52.075 ;
      RECT 69.55 -51.285 69.65 -50.75 ;
      RECT 69.55 -49.38 69.65 -48.845 ;
      RECT 69.55 -48.055 69.65 -47.52 ;
      RECT 69.55 -46.15 69.65 -45.615 ;
      RECT 69.55 -44.825 69.65 -44.29 ;
      RECT 69.55 -42.92 69.65 -42.385 ;
      RECT 69.55 -41.595 69.65 -41.06 ;
      RECT 69.55 -39.69 69.65 -39.155 ;
      RECT 69.55 -38.365 69.65 -37.83 ;
      RECT 69.55 -36.46 69.65 -35.925 ;
      RECT 69.55 -35.135 69.65 -34.6 ;
      RECT 69.55 -33.23 69.65 -32.695 ;
      RECT 69.55 -31.905 69.65 -31.37 ;
      RECT 69.55 -30 69.65 -29.465 ;
      RECT 69.55 -28.675 69.65 -28.14 ;
      RECT 69.55 -26.77 69.65 -26.235 ;
      RECT 69.55 -25.445 69.65 -24.91 ;
      RECT 69.55 -23.54 69.65 -23.005 ;
      RECT 69.55 -22.215 69.65 -21.68 ;
      RECT 69.55 -20.31 69.65 -19.775 ;
      RECT 69.55 -18.985 69.65 -18.45 ;
      RECT 69.55 -17.08 69.65 -16.545 ;
      RECT 69.55 -15.755 69.65 -15.22 ;
      RECT 69.55 -13.85 69.65 -13.315 ;
      RECT 69.55 -12.525 69.65 -11.99 ;
      RECT 69.55 -10.62 69.65 -10.085 ;
      RECT 69.55 -9.295 69.65 -8.76 ;
      RECT 69.55 -7.39 69.65 -6.855 ;
      RECT 69.55 -6.065 69.65 -5.53 ;
      RECT 69.55 -4.16 69.65 -3.625 ;
      RECT 69.55 -2.835 69.65 -2.3 ;
      RECT 69.55 -0.93 69.65 -0.395 ;
      RECT 69.55 0.395 69.65 0.93 ;
      RECT 69.425 -108.175 69.525 -107.215 ;
      RECT 69.05 -100.19 69.4 -100.07 ;
      RECT 69.05 -96.96 69.4 -96.84 ;
      RECT 69.05 -93.73 69.4 -93.61 ;
      RECT 69.05 -90.5 69.4 -90.38 ;
      RECT 69.05 -87.27 69.4 -87.15 ;
      RECT 69.05 -84.04 69.4 -83.92 ;
      RECT 69.05 -80.81 69.4 -80.69 ;
      RECT 69.05 -77.58 69.4 -77.46 ;
      RECT 69.05 -74.35 69.4 -74.23 ;
      RECT 69.05 -71.12 69.4 -71 ;
      RECT 69.05 -67.89 69.4 -67.77 ;
      RECT 69.05 -64.66 69.4 -64.54 ;
      RECT 69.05 -61.43 69.4 -61.31 ;
      RECT 69.05 -58.2 69.4 -58.08 ;
      RECT 69.05 -54.97 69.4 -54.85 ;
      RECT 69.05 -51.74 69.4 -51.62 ;
      RECT 69.05 -48.51 69.4 -48.39 ;
      RECT 69.05 -45.28 69.4 -45.16 ;
      RECT 69.05 -42.05 69.4 -41.93 ;
      RECT 69.05 -38.82 69.4 -38.7 ;
      RECT 69.05 -35.59 69.4 -35.47 ;
      RECT 69.05 -32.36 69.4 -32.24 ;
      RECT 69.05 -29.13 69.4 -29.01 ;
      RECT 69.05 -25.9 69.4 -25.78 ;
      RECT 69.05 -22.67 69.4 -22.55 ;
      RECT 69.05 -19.44 69.4 -19.32 ;
      RECT 69.05 -16.21 69.4 -16.09 ;
      RECT 69.05 -12.98 69.4 -12.86 ;
      RECT 69.05 -9.75 69.4 -9.63 ;
      RECT 69.05 -6.52 69.4 -6.4 ;
      RECT 69.05 -3.29 69.4 -3.17 ;
      RECT 69.05 -0.06 69.4 0.06 ;
      RECT 69.255 -112.255 69.355 -111.775 ;
      RECT 69.255 -110.765 69.355 -110.295 ;
      RECT 69.165 -108.175 69.265 -107.215 ;
      RECT 69.165 2.175 69.265 3.135 ;
      RECT 68.565 -100.19 68.915 -100.07 ;
      RECT 68.565 -96.96 68.915 -96.84 ;
      RECT 68.565 -93.73 68.915 -93.61 ;
      RECT 68.565 -90.5 68.915 -90.38 ;
      RECT 68.565 -87.27 68.915 -87.15 ;
      RECT 68.565 -84.04 68.915 -83.92 ;
      RECT 68.565 -80.81 68.915 -80.69 ;
      RECT 68.565 -77.58 68.915 -77.46 ;
      RECT 68.565 -74.35 68.915 -74.23 ;
      RECT 68.565 -71.12 68.915 -71 ;
      RECT 68.565 -67.89 68.915 -67.77 ;
      RECT 68.565 -64.66 68.915 -64.54 ;
      RECT 68.565 -61.43 68.915 -61.31 ;
      RECT 68.565 -58.2 68.915 -58.08 ;
      RECT 68.565 -54.97 68.915 -54.85 ;
      RECT 68.565 -51.74 68.915 -51.62 ;
      RECT 68.565 -48.51 68.915 -48.39 ;
      RECT 68.565 -45.28 68.915 -45.16 ;
      RECT 68.565 -42.05 68.915 -41.93 ;
      RECT 68.565 -38.82 68.915 -38.7 ;
      RECT 68.565 -35.59 68.915 -35.47 ;
      RECT 68.565 -32.36 68.915 -32.24 ;
      RECT 68.565 -29.13 68.915 -29.01 ;
      RECT 68.565 -25.9 68.915 -25.78 ;
      RECT 68.565 -22.67 68.915 -22.55 ;
      RECT 68.565 -19.44 68.915 -19.32 ;
      RECT 68.565 -16.21 68.915 -16.09 ;
      RECT 68.565 -12.98 68.915 -12.86 ;
      RECT 68.565 -9.75 68.915 -9.63 ;
      RECT 68.565 -6.52 68.915 -6.4 ;
      RECT 68.565 -3.29 68.915 -3.17 ;
      RECT 68.565 -0.06 68.915 0.06 ;
      RECT 68.735 -108.175 68.835 -107.215 ;
      RECT 68.735 2.175 68.835 3.135 ;
      RECT 68.63 -110.765 68.8 -110.385 ;
      RECT 68.665 -112.245 68.765 -111.775 ;
      RECT 68.475 -108.175 68.575 -107.215 ;
      RECT 68.35 -101.06 68.45 -100.525 ;
      RECT 68.35 -99.735 68.45 -99.2 ;
      RECT 68.35 -97.83 68.45 -97.295 ;
      RECT 68.35 -96.505 68.45 -95.97 ;
      RECT 68.35 -94.6 68.45 -94.065 ;
      RECT 68.35 -93.275 68.45 -92.74 ;
      RECT 68.35 -91.37 68.45 -90.835 ;
      RECT 68.35 -90.045 68.45 -89.51 ;
      RECT 68.35 -88.14 68.45 -87.605 ;
      RECT 68.35 -86.815 68.45 -86.28 ;
      RECT 68.35 -84.91 68.45 -84.375 ;
      RECT 68.35 -83.585 68.45 -83.05 ;
      RECT 68.35 -81.68 68.45 -81.145 ;
      RECT 68.35 -80.355 68.45 -79.82 ;
      RECT 68.35 -78.45 68.45 -77.915 ;
      RECT 68.35 -77.125 68.45 -76.59 ;
      RECT 68.35 -75.22 68.45 -74.685 ;
      RECT 68.35 -73.895 68.45 -73.36 ;
      RECT 68.35 -71.99 68.45 -71.455 ;
      RECT 68.35 -70.665 68.45 -70.13 ;
      RECT 68.35 -68.76 68.45 -68.225 ;
      RECT 68.35 -67.435 68.45 -66.9 ;
      RECT 68.35 -65.53 68.45 -64.995 ;
      RECT 68.35 -64.205 68.45 -63.67 ;
      RECT 68.35 -62.3 68.45 -61.765 ;
      RECT 68.35 -60.975 68.45 -60.44 ;
      RECT 68.35 -59.07 68.45 -58.535 ;
      RECT 68.35 -57.745 68.45 -57.21 ;
      RECT 68.35 -55.84 68.45 -55.305 ;
      RECT 68.35 -54.515 68.45 -53.98 ;
      RECT 68.35 -52.61 68.45 -52.075 ;
      RECT 68.35 -51.285 68.45 -50.75 ;
      RECT 68.35 -49.38 68.45 -48.845 ;
      RECT 68.35 -48.055 68.45 -47.52 ;
      RECT 68.35 -46.15 68.45 -45.615 ;
      RECT 68.35 -44.825 68.45 -44.29 ;
      RECT 68.35 -42.92 68.45 -42.385 ;
      RECT 68.35 -41.595 68.45 -41.06 ;
      RECT 68.35 -39.69 68.45 -39.155 ;
      RECT 68.35 -38.365 68.45 -37.83 ;
      RECT 68.35 -36.46 68.45 -35.925 ;
      RECT 68.35 -35.135 68.45 -34.6 ;
      RECT 68.35 -33.23 68.45 -32.695 ;
      RECT 68.35 -31.905 68.45 -31.37 ;
      RECT 68.35 -30 68.45 -29.465 ;
      RECT 68.35 -28.675 68.45 -28.14 ;
      RECT 68.35 -26.77 68.45 -26.235 ;
      RECT 68.35 -25.445 68.45 -24.91 ;
      RECT 68.35 -23.54 68.45 -23.005 ;
      RECT 68.35 -22.215 68.45 -21.68 ;
      RECT 68.35 -20.31 68.45 -19.775 ;
      RECT 68.35 -18.985 68.45 -18.45 ;
      RECT 68.35 -17.08 68.45 -16.545 ;
      RECT 68.35 -15.755 68.45 -15.22 ;
      RECT 68.35 -13.85 68.45 -13.315 ;
      RECT 68.35 -12.525 68.45 -11.99 ;
      RECT 68.35 -10.62 68.45 -10.085 ;
      RECT 68.35 -9.295 68.45 -8.76 ;
      RECT 68.35 -7.39 68.45 -6.855 ;
      RECT 68.35 -6.065 68.45 -5.53 ;
      RECT 68.35 -4.16 68.45 -3.625 ;
      RECT 68.35 -2.835 68.45 -2.3 ;
      RECT 68.35 -0.93 68.45 -0.395 ;
      RECT 68.35 0.395 68.45 0.93 ;
      RECT 68.225 -108.175 68.325 -107.215 ;
      RECT 67.85 -100.19 68.2 -100.07 ;
      RECT 67.85 -96.96 68.2 -96.84 ;
      RECT 67.85 -93.73 68.2 -93.61 ;
      RECT 67.85 -90.5 68.2 -90.38 ;
      RECT 67.85 -87.27 68.2 -87.15 ;
      RECT 67.85 -84.04 68.2 -83.92 ;
      RECT 67.85 -80.81 68.2 -80.69 ;
      RECT 67.85 -77.58 68.2 -77.46 ;
      RECT 67.85 -74.35 68.2 -74.23 ;
      RECT 67.85 -71.12 68.2 -71 ;
      RECT 67.85 -67.89 68.2 -67.77 ;
      RECT 67.85 -64.66 68.2 -64.54 ;
      RECT 67.85 -61.43 68.2 -61.31 ;
      RECT 67.85 -58.2 68.2 -58.08 ;
      RECT 67.85 -54.97 68.2 -54.85 ;
      RECT 67.85 -51.74 68.2 -51.62 ;
      RECT 67.85 -48.51 68.2 -48.39 ;
      RECT 67.85 -45.28 68.2 -45.16 ;
      RECT 67.85 -42.05 68.2 -41.93 ;
      RECT 67.85 -38.82 68.2 -38.7 ;
      RECT 67.85 -35.59 68.2 -35.47 ;
      RECT 67.85 -32.36 68.2 -32.24 ;
      RECT 67.85 -29.13 68.2 -29.01 ;
      RECT 67.85 -25.9 68.2 -25.78 ;
      RECT 67.85 -22.67 68.2 -22.55 ;
      RECT 67.85 -19.44 68.2 -19.32 ;
      RECT 67.85 -16.21 68.2 -16.09 ;
      RECT 67.85 -12.98 68.2 -12.86 ;
      RECT 67.85 -9.75 68.2 -9.63 ;
      RECT 67.85 -6.52 68.2 -6.4 ;
      RECT 67.85 -3.29 68.2 -3.17 ;
      RECT 67.85 -0.06 68.2 0.06 ;
      RECT 67.965 -108.175 68.065 -107.215 ;
      RECT 67.965 2.175 68.065 3.135 ;
      RECT 67.865 -113.555 67.965 -113.085 ;
      RECT 67.365 -100.19 67.715 -100.07 ;
      RECT 67.365 -96.96 67.715 -96.84 ;
      RECT 67.365 -93.73 67.715 -93.61 ;
      RECT 67.365 -90.5 67.715 -90.38 ;
      RECT 67.365 -87.27 67.715 -87.15 ;
      RECT 67.365 -84.04 67.715 -83.92 ;
      RECT 67.365 -80.81 67.715 -80.69 ;
      RECT 67.365 -77.58 67.715 -77.46 ;
      RECT 67.365 -74.35 67.715 -74.23 ;
      RECT 67.365 -71.12 67.715 -71 ;
      RECT 67.365 -67.89 67.715 -67.77 ;
      RECT 67.365 -64.66 67.715 -64.54 ;
      RECT 67.365 -61.43 67.715 -61.31 ;
      RECT 67.365 -58.2 67.715 -58.08 ;
      RECT 67.365 -54.97 67.715 -54.85 ;
      RECT 67.365 -51.74 67.715 -51.62 ;
      RECT 67.365 -48.51 67.715 -48.39 ;
      RECT 67.365 -45.28 67.715 -45.16 ;
      RECT 67.365 -42.05 67.715 -41.93 ;
      RECT 67.365 -38.82 67.715 -38.7 ;
      RECT 67.365 -35.59 67.715 -35.47 ;
      RECT 67.365 -32.36 67.715 -32.24 ;
      RECT 67.365 -29.13 67.715 -29.01 ;
      RECT 67.365 -25.9 67.715 -25.78 ;
      RECT 67.365 -22.67 67.715 -22.55 ;
      RECT 67.365 -19.44 67.715 -19.32 ;
      RECT 67.365 -16.21 67.715 -16.09 ;
      RECT 67.365 -12.98 67.715 -12.86 ;
      RECT 67.365 -9.75 67.715 -9.63 ;
      RECT 67.365 -6.52 67.715 -6.4 ;
      RECT 67.365 -3.29 67.715 -3.17 ;
      RECT 67.365 -0.06 67.715 0.06 ;
      RECT 67.5 -110.735 67.65 -110.445 ;
      RECT 67.535 -108.175 67.635 -107.215 ;
      RECT 67.535 2.175 67.635 3.135 ;
      RECT 67.515 -112.19 67.615 -111.65 ;
      RECT 67.275 -113.555 67.375 -113.085 ;
      RECT 67.275 -108.175 67.375 -107.215 ;
      RECT 67.15 -101.06 67.25 -100.525 ;
      RECT 67.15 -99.735 67.25 -99.2 ;
      RECT 67.15 -97.83 67.25 -97.295 ;
      RECT 67.15 -96.505 67.25 -95.97 ;
      RECT 67.15 -94.6 67.25 -94.065 ;
      RECT 67.15 -93.275 67.25 -92.74 ;
      RECT 67.15 -91.37 67.25 -90.835 ;
      RECT 67.15 -90.045 67.25 -89.51 ;
      RECT 67.15 -88.14 67.25 -87.605 ;
      RECT 67.15 -86.815 67.25 -86.28 ;
      RECT 67.15 -84.91 67.25 -84.375 ;
      RECT 67.15 -83.585 67.25 -83.05 ;
      RECT 67.15 -81.68 67.25 -81.145 ;
      RECT 67.15 -80.355 67.25 -79.82 ;
      RECT 67.15 -78.45 67.25 -77.915 ;
      RECT 67.15 -77.125 67.25 -76.59 ;
      RECT 67.15 -75.22 67.25 -74.685 ;
      RECT 67.15 -73.895 67.25 -73.36 ;
      RECT 67.15 -71.99 67.25 -71.455 ;
      RECT 67.15 -70.665 67.25 -70.13 ;
      RECT 67.15 -68.76 67.25 -68.225 ;
      RECT 67.15 -67.435 67.25 -66.9 ;
      RECT 67.15 -65.53 67.25 -64.995 ;
      RECT 67.15 -64.205 67.25 -63.67 ;
      RECT 67.15 -62.3 67.25 -61.765 ;
      RECT 67.15 -60.975 67.25 -60.44 ;
      RECT 67.15 -59.07 67.25 -58.535 ;
      RECT 67.15 -57.745 67.25 -57.21 ;
      RECT 67.15 -55.84 67.25 -55.305 ;
      RECT 67.15 -54.515 67.25 -53.98 ;
      RECT 67.15 -52.61 67.25 -52.075 ;
      RECT 67.15 -51.285 67.25 -50.75 ;
      RECT 67.15 -49.38 67.25 -48.845 ;
      RECT 67.15 -48.055 67.25 -47.52 ;
      RECT 67.15 -46.15 67.25 -45.615 ;
      RECT 67.15 -44.825 67.25 -44.29 ;
      RECT 67.15 -42.92 67.25 -42.385 ;
      RECT 67.15 -41.595 67.25 -41.06 ;
      RECT 67.15 -39.69 67.25 -39.155 ;
      RECT 67.15 -38.365 67.25 -37.83 ;
      RECT 67.15 -36.46 67.25 -35.925 ;
      RECT 67.15 -35.135 67.25 -34.6 ;
      RECT 67.15 -33.23 67.25 -32.695 ;
      RECT 67.15 -31.905 67.25 -31.37 ;
      RECT 67.15 -30 67.25 -29.465 ;
      RECT 67.15 -28.675 67.25 -28.14 ;
      RECT 67.15 -26.77 67.25 -26.235 ;
      RECT 67.15 -25.445 67.25 -24.91 ;
      RECT 67.15 -23.54 67.25 -23.005 ;
      RECT 67.15 -22.215 67.25 -21.68 ;
      RECT 67.15 -20.31 67.25 -19.775 ;
      RECT 67.15 -18.985 67.25 -18.45 ;
      RECT 67.15 -17.08 67.25 -16.545 ;
      RECT 67.15 -15.755 67.25 -15.22 ;
      RECT 67.15 -13.85 67.25 -13.315 ;
      RECT 67.15 -12.525 67.25 -11.99 ;
      RECT 67.15 -10.62 67.25 -10.085 ;
      RECT 67.15 -9.295 67.25 -8.76 ;
      RECT 67.15 -7.39 67.25 -6.855 ;
      RECT 67.15 -6.065 67.25 -5.53 ;
      RECT 67.15 -4.16 67.25 -3.625 ;
      RECT 67.15 -2.835 67.25 -2.3 ;
      RECT 67.15 -0.93 67.25 -0.395 ;
      RECT 67.15 0.395 67.25 0.93 ;
      RECT 67.025 -104.945 67.125 -103.985 ;
      RECT 66.65 -100.19 67 -100.07 ;
      RECT 66.65 -96.96 67 -96.84 ;
      RECT 66.65 -93.73 67 -93.61 ;
      RECT 66.65 -90.5 67 -90.38 ;
      RECT 66.65 -87.27 67 -87.15 ;
      RECT 66.65 -84.04 67 -83.92 ;
      RECT 66.65 -80.81 67 -80.69 ;
      RECT 66.65 -77.58 67 -77.46 ;
      RECT 66.65 -74.35 67 -74.23 ;
      RECT 66.65 -71.12 67 -71 ;
      RECT 66.65 -67.89 67 -67.77 ;
      RECT 66.65 -64.66 67 -64.54 ;
      RECT 66.65 -61.43 67 -61.31 ;
      RECT 66.65 -58.2 67 -58.08 ;
      RECT 66.65 -54.97 67 -54.85 ;
      RECT 66.65 -51.74 67 -51.62 ;
      RECT 66.65 -48.51 67 -48.39 ;
      RECT 66.65 -45.28 67 -45.16 ;
      RECT 66.65 -42.05 67 -41.93 ;
      RECT 66.65 -38.82 67 -38.7 ;
      RECT 66.65 -35.59 67 -35.47 ;
      RECT 66.65 -32.36 67 -32.24 ;
      RECT 66.65 -29.13 67 -29.01 ;
      RECT 66.65 -25.9 67 -25.78 ;
      RECT 66.65 -22.67 67 -22.55 ;
      RECT 66.65 -19.44 67 -19.32 ;
      RECT 66.65 -16.21 67 -16.09 ;
      RECT 66.65 -12.98 67 -12.86 ;
      RECT 66.65 -9.75 67 -9.63 ;
      RECT 66.65 -6.52 67 -6.4 ;
      RECT 66.65 -3.29 67 -3.17 ;
      RECT 66.65 -0.06 67 0.06 ;
      RECT 66.765 -104.945 66.865 -103.985 ;
      RECT 66.765 2.175 66.865 3.135 ;
      RECT 66.475 -112.255 66.575 -111.775 ;
      RECT 66.475 -110.765 66.575 -110.295 ;
      RECT 66.165 -100.19 66.515 -100.07 ;
      RECT 66.165 -96.96 66.515 -96.84 ;
      RECT 66.165 -93.73 66.515 -93.61 ;
      RECT 66.165 -90.5 66.515 -90.38 ;
      RECT 66.165 -87.27 66.515 -87.15 ;
      RECT 66.165 -84.04 66.515 -83.92 ;
      RECT 66.165 -80.81 66.515 -80.69 ;
      RECT 66.165 -77.58 66.515 -77.46 ;
      RECT 66.165 -74.35 66.515 -74.23 ;
      RECT 66.165 -71.12 66.515 -71 ;
      RECT 66.165 -67.89 66.515 -67.77 ;
      RECT 66.165 -64.66 66.515 -64.54 ;
      RECT 66.165 -61.43 66.515 -61.31 ;
      RECT 66.165 -58.2 66.515 -58.08 ;
      RECT 66.165 -54.97 66.515 -54.85 ;
      RECT 66.165 -51.74 66.515 -51.62 ;
      RECT 66.165 -48.51 66.515 -48.39 ;
      RECT 66.165 -45.28 66.515 -45.16 ;
      RECT 66.165 -42.05 66.515 -41.93 ;
      RECT 66.165 -38.82 66.515 -38.7 ;
      RECT 66.165 -35.59 66.515 -35.47 ;
      RECT 66.165 -32.36 66.515 -32.24 ;
      RECT 66.165 -29.13 66.515 -29.01 ;
      RECT 66.165 -25.9 66.515 -25.78 ;
      RECT 66.165 -22.67 66.515 -22.55 ;
      RECT 66.165 -19.44 66.515 -19.32 ;
      RECT 66.165 -16.21 66.515 -16.09 ;
      RECT 66.165 -12.98 66.515 -12.86 ;
      RECT 66.165 -9.75 66.515 -9.63 ;
      RECT 66.165 -6.52 66.515 -6.4 ;
      RECT 66.165 -3.29 66.515 -3.17 ;
      RECT 66.165 -0.06 66.515 0.06 ;
      RECT 66.335 -104.945 66.435 -103.985 ;
      RECT 66.335 2.175 66.435 3.135 ;
      RECT 62.435 -108.655 66.215 -108.535 ;
      RECT 66.075 -104.945 66.175 -103.985 ;
      RECT 65.95 -101.06 66.05 -100.525 ;
      RECT 65.95 -99.735 66.05 -99.2 ;
      RECT 65.95 -97.83 66.05 -97.295 ;
      RECT 65.95 -96.505 66.05 -95.97 ;
      RECT 65.95 -94.6 66.05 -94.065 ;
      RECT 65.95 -93.275 66.05 -92.74 ;
      RECT 65.95 -91.37 66.05 -90.835 ;
      RECT 65.95 -90.045 66.05 -89.51 ;
      RECT 65.95 -88.14 66.05 -87.605 ;
      RECT 65.95 -86.815 66.05 -86.28 ;
      RECT 65.95 -84.91 66.05 -84.375 ;
      RECT 65.95 -83.585 66.05 -83.05 ;
      RECT 65.95 -81.68 66.05 -81.145 ;
      RECT 65.95 -80.355 66.05 -79.82 ;
      RECT 65.95 -78.45 66.05 -77.915 ;
      RECT 65.95 -77.125 66.05 -76.59 ;
      RECT 65.95 -75.22 66.05 -74.685 ;
      RECT 65.95 -73.895 66.05 -73.36 ;
      RECT 65.95 -71.99 66.05 -71.455 ;
      RECT 65.95 -70.665 66.05 -70.13 ;
      RECT 65.95 -68.76 66.05 -68.225 ;
      RECT 65.95 -67.435 66.05 -66.9 ;
      RECT 65.95 -65.53 66.05 -64.995 ;
      RECT 65.95 -64.205 66.05 -63.67 ;
      RECT 65.95 -62.3 66.05 -61.765 ;
      RECT 65.95 -60.975 66.05 -60.44 ;
      RECT 65.95 -59.07 66.05 -58.535 ;
      RECT 65.95 -57.745 66.05 -57.21 ;
      RECT 65.95 -55.84 66.05 -55.305 ;
      RECT 65.95 -54.515 66.05 -53.98 ;
      RECT 65.95 -52.61 66.05 -52.075 ;
      RECT 65.95 -51.285 66.05 -50.75 ;
      RECT 65.95 -49.38 66.05 -48.845 ;
      RECT 65.95 -48.055 66.05 -47.52 ;
      RECT 65.95 -46.15 66.05 -45.615 ;
      RECT 65.95 -44.825 66.05 -44.29 ;
      RECT 65.95 -42.92 66.05 -42.385 ;
      RECT 65.95 -41.595 66.05 -41.06 ;
      RECT 65.95 -39.69 66.05 -39.155 ;
      RECT 65.95 -38.365 66.05 -37.83 ;
      RECT 65.95 -36.46 66.05 -35.925 ;
      RECT 65.95 -35.135 66.05 -34.6 ;
      RECT 65.95 -33.23 66.05 -32.695 ;
      RECT 65.95 -31.905 66.05 -31.37 ;
      RECT 65.95 -30 66.05 -29.465 ;
      RECT 65.95 -28.675 66.05 -28.14 ;
      RECT 65.95 -26.77 66.05 -26.235 ;
      RECT 65.95 -25.445 66.05 -24.91 ;
      RECT 65.95 -23.54 66.05 -23.005 ;
      RECT 65.95 -22.215 66.05 -21.68 ;
      RECT 65.95 -20.31 66.05 -19.775 ;
      RECT 65.95 -18.985 66.05 -18.45 ;
      RECT 65.95 -17.08 66.05 -16.545 ;
      RECT 65.95 -15.755 66.05 -15.22 ;
      RECT 65.95 -13.85 66.05 -13.315 ;
      RECT 65.95 -12.525 66.05 -11.99 ;
      RECT 65.95 -10.62 66.05 -10.085 ;
      RECT 65.95 -9.295 66.05 -8.76 ;
      RECT 65.95 -7.39 66.05 -6.855 ;
      RECT 65.95 -6.065 66.05 -5.53 ;
      RECT 65.95 -4.16 66.05 -3.625 ;
      RECT 65.95 -2.835 66.05 -2.3 ;
      RECT 65.95 -0.93 66.05 -0.395 ;
      RECT 65.95 0.395 66.05 0.93 ;
      RECT 65.885 -110.75 66.005 -110.37 ;
      RECT 65.885 -112.245 65.985 -111.775 ;
      RECT 65.825 -104.945 65.925 -103.985 ;
      RECT 65.45 -100.19 65.8 -100.07 ;
      RECT 65.45 -96.96 65.8 -96.84 ;
      RECT 65.45 -93.73 65.8 -93.61 ;
      RECT 65.45 -90.5 65.8 -90.38 ;
      RECT 65.45 -87.27 65.8 -87.15 ;
      RECT 65.45 -84.04 65.8 -83.92 ;
      RECT 65.45 -80.81 65.8 -80.69 ;
      RECT 65.45 -77.58 65.8 -77.46 ;
      RECT 65.45 -74.35 65.8 -74.23 ;
      RECT 65.45 -71.12 65.8 -71 ;
      RECT 65.45 -67.89 65.8 -67.77 ;
      RECT 65.45 -64.66 65.8 -64.54 ;
      RECT 65.45 -61.43 65.8 -61.31 ;
      RECT 65.45 -58.2 65.8 -58.08 ;
      RECT 65.45 -54.97 65.8 -54.85 ;
      RECT 65.45 -51.74 65.8 -51.62 ;
      RECT 65.45 -48.51 65.8 -48.39 ;
      RECT 65.45 -45.28 65.8 -45.16 ;
      RECT 65.45 -42.05 65.8 -41.93 ;
      RECT 65.45 -38.82 65.8 -38.7 ;
      RECT 65.45 -35.59 65.8 -35.47 ;
      RECT 65.45 -32.36 65.8 -32.24 ;
      RECT 65.45 -29.13 65.8 -29.01 ;
      RECT 65.45 -25.9 65.8 -25.78 ;
      RECT 65.45 -22.67 65.8 -22.55 ;
      RECT 65.45 -19.44 65.8 -19.32 ;
      RECT 65.45 -16.21 65.8 -16.09 ;
      RECT 65.45 -12.98 65.8 -12.86 ;
      RECT 65.45 -9.75 65.8 -9.63 ;
      RECT 65.45 -6.52 65.8 -6.4 ;
      RECT 65.45 -3.29 65.8 -3.17 ;
      RECT 65.45 -0.06 65.8 0.06 ;
      RECT 65.565 -104.945 65.665 -103.985 ;
      RECT 65.565 2.175 65.665 3.135 ;
      RECT 65.295 -109.595 65.43 -109.275 ;
      RECT 64.965 -100.19 65.315 -100.07 ;
      RECT 64.965 -96.96 65.315 -96.84 ;
      RECT 64.965 -93.73 65.315 -93.61 ;
      RECT 64.965 -90.5 65.315 -90.38 ;
      RECT 64.965 -87.27 65.315 -87.15 ;
      RECT 64.965 -84.04 65.315 -83.92 ;
      RECT 64.965 -80.81 65.315 -80.69 ;
      RECT 64.965 -77.58 65.315 -77.46 ;
      RECT 64.965 -74.35 65.315 -74.23 ;
      RECT 64.965 -71.12 65.315 -71 ;
      RECT 64.965 -67.89 65.315 -67.77 ;
      RECT 64.965 -64.66 65.315 -64.54 ;
      RECT 64.965 -61.43 65.315 -61.31 ;
      RECT 64.965 -58.2 65.315 -58.08 ;
      RECT 64.965 -54.97 65.315 -54.85 ;
      RECT 64.965 -51.74 65.315 -51.62 ;
      RECT 64.965 -48.51 65.315 -48.39 ;
      RECT 64.965 -45.28 65.315 -45.16 ;
      RECT 64.965 -42.05 65.315 -41.93 ;
      RECT 64.965 -38.82 65.315 -38.7 ;
      RECT 64.965 -35.59 65.315 -35.47 ;
      RECT 64.965 -32.36 65.315 -32.24 ;
      RECT 64.965 -29.13 65.315 -29.01 ;
      RECT 64.965 -25.9 65.315 -25.78 ;
      RECT 64.965 -22.67 65.315 -22.55 ;
      RECT 64.965 -19.44 65.315 -19.32 ;
      RECT 64.965 -16.21 65.315 -16.09 ;
      RECT 64.965 -12.98 65.315 -12.86 ;
      RECT 64.965 -9.75 65.315 -9.63 ;
      RECT 64.965 -6.52 65.315 -6.4 ;
      RECT 64.965 -3.29 65.315 -3.17 ;
      RECT 64.965 -0.06 65.315 0.06 ;
      RECT 65.135 -104.945 65.235 -103.985 ;
      RECT 65.135 2.175 65.235 3.135 ;
      RECT 64.96 -109.595 65.105 -109.275 ;
      RECT 64.875 -104.945 64.975 -103.985 ;
      RECT 64.75 -101.06 64.85 -100.525 ;
      RECT 64.75 -99.735 64.85 -99.2 ;
      RECT 64.75 -97.83 64.85 -97.295 ;
      RECT 64.75 -96.505 64.85 -95.97 ;
      RECT 64.75 -94.6 64.85 -94.065 ;
      RECT 64.75 -93.275 64.85 -92.74 ;
      RECT 64.75 -91.37 64.85 -90.835 ;
      RECT 64.75 -90.045 64.85 -89.51 ;
      RECT 64.75 -88.14 64.85 -87.605 ;
      RECT 64.75 -86.815 64.85 -86.28 ;
      RECT 64.75 -84.91 64.85 -84.375 ;
      RECT 64.75 -83.585 64.85 -83.05 ;
      RECT 64.75 -81.68 64.85 -81.145 ;
      RECT 64.75 -80.355 64.85 -79.82 ;
      RECT 64.75 -78.45 64.85 -77.915 ;
      RECT 64.75 -77.125 64.85 -76.59 ;
      RECT 64.75 -75.22 64.85 -74.685 ;
      RECT 64.75 -73.895 64.85 -73.36 ;
      RECT 64.75 -71.99 64.85 -71.455 ;
      RECT 64.75 -70.665 64.85 -70.13 ;
      RECT 64.75 -68.76 64.85 -68.225 ;
      RECT 64.75 -67.435 64.85 -66.9 ;
      RECT 64.75 -65.53 64.85 -64.995 ;
      RECT 64.75 -64.205 64.85 -63.67 ;
      RECT 64.75 -62.3 64.85 -61.765 ;
      RECT 64.75 -60.975 64.85 -60.44 ;
      RECT 64.75 -59.07 64.85 -58.535 ;
      RECT 64.75 -57.745 64.85 -57.21 ;
      RECT 64.75 -55.84 64.85 -55.305 ;
      RECT 64.75 -54.515 64.85 -53.98 ;
      RECT 64.75 -52.61 64.85 -52.075 ;
      RECT 64.75 -51.285 64.85 -50.75 ;
      RECT 64.75 -49.38 64.85 -48.845 ;
      RECT 64.75 -48.055 64.85 -47.52 ;
      RECT 64.75 -46.15 64.85 -45.615 ;
      RECT 64.75 -44.825 64.85 -44.29 ;
      RECT 64.75 -42.92 64.85 -42.385 ;
      RECT 64.75 -41.595 64.85 -41.06 ;
      RECT 64.75 -39.69 64.85 -39.155 ;
      RECT 64.75 -38.365 64.85 -37.83 ;
      RECT 64.75 -36.46 64.85 -35.925 ;
      RECT 64.75 -35.135 64.85 -34.6 ;
      RECT 64.75 -33.23 64.85 -32.695 ;
      RECT 64.75 -31.905 64.85 -31.37 ;
      RECT 64.75 -30 64.85 -29.465 ;
      RECT 64.75 -28.675 64.85 -28.14 ;
      RECT 64.75 -26.77 64.85 -26.235 ;
      RECT 64.75 -25.445 64.85 -24.91 ;
      RECT 64.75 -23.54 64.85 -23.005 ;
      RECT 64.75 -22.215 64.85 -21.68 ;
      RECT 64.75 -20.31 64.85 -19.775 ;
      RECT 64.75 -18.985 64.85 -18.45 ;
      RECT 64.75 -17.08 64.85 -16.545 ;
      RECT 64.75 -15.755 64.85 -15.22 ;
      RECT 64.75 -13.85 64.85 -13.315 ;
      RECT 64.75 -12.525 64.85 -11.99 ;
      RECT 64.75 -10.62 64.85 -10.085 ;
      RECT 64.75 -9.295 64.85 -8.76 ;
      RECT 64.75 -7.39 64.85 -6.855 ;
      RECT 64.75 -6.065 64.85 -5.53 ;
      RECT 64.75 -4.16 64.85 -3.625 ;
      RECT 64.75 -2.835 64.85 -2.3 ;
      RECT 64.75 -0.93 64.85 -0.395 ;
      RECT 64.75 0.395 64.85 0.93 ;
      RECT 64.625 -108.175 64.725 -107.215 ;
      RECT 64.25 -100.19 64.6 -100.07 ;
      RECT 64.25 -96.96 64.6 -96.84 ;
      RECT 64.25 -93.73 64.6 -93.61 ;
      RECT 64.25 -90.5 64.6 -90.38 ;
      RECT 64.25 -87.27 64.6 -87.15 ;
      RECT 64.25 -84.04 64.6 -83.92 ;
      RECT 64.25 -80.81 64.6 -80.69 ;
      RECT 64.25 -77.58 64.6 -77.46 ;
      RECT 64.25 -74.35 64.6 -74.23 ;
      RECT 64.25 -71.12 64.6 -71 ;
      RECT 64.25 -67.89 64.6 -67.77 ;
      RECT 64.25 -64.66 64.6 -64.54 ;
      RECT 64.25 -61.43 64.6 -61.31 ;
      RECT 64.25 -58.2 64.6 -58.08 ;
      RECT 64.25 -54.97 64.6 -54.85 ;
      RECT 64.25 -51.74 64.6 -51.62 ;
      RECT 64.25 -48.51 64.6 -48.39 ;
      RECT 64.25 -45.28 64.6 -45.16 ;
      RECT 64.25 -42.05 64.6 -41.93 ;
      RECT 64.25 -38.82 64.6 -38.7 ;
      RECT 64.25 -35.59 64.6 -35.47 ;
      RECT 64.25 -32.36 64.6 -32.24 ;
      RECT 64.25 -29.13 64.6 -29.01 ;
      RECT 64.25 -25.9 64.6 -25.78 ;
      RECT 64.25 -22.67 64.6 -22.55 ;
      RECT 64.25 -19.44 64.6 -19.32 ;
      RECT 64.25 -16.21 64.6 -16.09 ;
      RECT 64.25 -12.98 64.6 -12.86 ;
      RECT 64.25 -9.75 64.6 -9.63 ;
      RECT 64.25 -6.52 64.6 -6.4 ;
      RECT 64.25 -3.29 64.6 -3.17 ;
      RECT 64.25 -0.06 64.6 0.06 ;
      RECT 64.455 -112.255 64.555 -111.775 ;
      RECT 64.455 -110.765 64.555 -110.295 ;
      RECT 64.365 -108.175 64.465 -107.215 ;
      RECT 64.365 2.175 64.465 3.135 ;
      RECT 63.765 -100.19 64.115 -100.07 ;
      RECT 63.765 -96.96 64.115 -96.84 ;
      RECT 63.765 -93.73 64.115 -93.61 ;
      RECT 63.765 -90.5 64.115 -90.38 ;
      RECT 63.765 -87.27 64.115 -87.15 ;
      RECT 63.765 -84.04 64.115 -83.92 ;
      RECT 63.765 -80.81 64.115 -80.69 ;
      RECT 63.765 -77.58 64.115 -77.46 ;
      RECT 63.765 -74.35 64.115 -74.23 ;
      RECT 63.765 -71.12 64.115 -71 ;
      RECT 63.765 -67.89 64.115 -67.77 ;
      RECT 63.765 -64.66 64.115 -64.54 ;
      RECT 63.765 -61.43 64.115 -61.31 ;
      RECT 63.765 -58.2 64.115 -58.08 ;
      RECT 63.765 -54.97 64.115 -54.85 ;
      RECT 63.765 -51.74 64.115 -51.62 ;
      RECT 63.765 -48.51 64.115 -48.39 ;
      RECT 63.765 -45.28 64.115 -45.16 ;
      RECT 63.765 -42.05 64.115 -41.93 ;
      RECT 63.765 -38.82 64.115 -38.7 ;
      RECT 63.765 -35.59 64.115 -35.47 ;
      RECT 63.765 -32.36 64.115 -32.24 ;
      RECT 63.765 -29.13 64.115 -29.01 ;
      RECT 63.765 -25.9 64.115 -25.78 ;
      RECT 63.765 -22.67 64.115 -22.55 ;
      RECT 63.765 -19.44 64.115 -19.32 ;
      RECT 63.765 -16.21 64.115 -16.09 ;
      RECT 63.765 -12.98 64.115 -12.86 ;
      RECT 63.765 -9.75 64.115 -9.63 ;
      RECT 63.765 -6.52 64.115 -6.4 ;
      RECT 63.765 -3.29 64.115 -3.17 ;
      RECT 63.765 -0.06 64.115 0.06 ;
      RECT 63.935 -108.175 64.035 -107.215 ;
      RECT 63.935 2.175 64.035 3.135 ;
      RECT 63.83 -110.765 64 -110.385 ;
      RECT 63.865 -112.245 63.965 -111.775 ;
      RECT 63.675 -108.175 63.775 -107.215 ;
      RECT 63.55 -101.06 63.65 -100.525 ;
      RECT 63.55 -99.735 63.65 -99.2 ;
      RECT 63.55 -97.83 63.65 -97.295 ;
      RECT 63.55 -96.505 63.65 -95.97 ;
      RECT 63.55 -94.6 63.65 -94.065 ;
      RECT 63.55 -93.275 63.65 -92.74 ;
      RECT 63.55 -91.37 63.65 -90.835 ;
      RECT 63.55 -90.045 63.65 -89.51 ;
      RECT 63.55 -88.14 63.65 -87.605 ;
      RECT 63.55 -86.815 63.65 -86.28 ;
      RECT 63.55 -84.91 63.65 -84.375 ;
      RECT 63.55 -83.585 63.65 -83.05 ;
      RECT 63.55 -81.68 63.65 -81.145 ;
      RECT 63.55 -80.355 63.65 -79.82 ;
      RECT 63.55 -78.45 63.65 -77.915 ;
      RECT 63.55 -77.125 63.65 -76.59 ;
      RECT 63.55 -75.22 63.65 -74.685 ;
      RECT 63.55 -73.895 63.65 -73.36 ;
      RECT 63.55 -71.99 63.65 -71.455 ;
      RECT 63.55 -70.665 63.65 -70.13 ;
      RECT 63.55 -68.76 63.65 -68.225 ;
      RECT 63.55 -67.435 63.65 -66.9 ;
      RECT 63.55 -65.53 63.65 -64.995 ;
      RECT 63.55 -64.205 63.65 -63.67 ;
      RECT 63.55 -62.3 63.65 -61.765 ;
      RECT 63.55 -60.975 63.65 -60.44 ;
      RECT 63.55 -59.07 63.65 -58.535 ;
      RECT 63.55 -57.745 63.65 -57.21 ;
      RECT 63.55 -55.84 63.65 -55.305 ;
      RECT 63.55 -54.515 63.65 -53.98 ;
      RECT 63.55 -52.61 63.65 -52.075 ;
      RECT 63.55 -51.285 63.65 -50.75 ;
      RECT 63.55 -49.38 63.65 -48.845 ;
      RECT 63.55 -48.055 63.65 -47.52 ;
      RECT 63.55 -46.15 63.65 -45.615 ;
      RECT 63.55 -44.825 63.65 -44.29 ;
      RECT 63.55 -42.92 63.65 -42.385 ;
      RECT 63.55 -41.595 63.65 -41.06 ;
      RECT 63.55 -39.69 63.65 -39.155 ;
      RECT 63.55 -38.365 63.65 -37.83 ;
      RECT 63.55 -36.46 63.65 -35.925 ;
      RECT 63.55 -35.135 63.65 -34.6 ;
      RECT 63.55 -33.23 63.65 -32.695 ;
      RECT 63.55 -31.905 63.65 -31.37 ;
      RECT 63.55 -30 63.65 -29.465 ;
      RECT 63.55 -28.675 63.65 -28.14 ;
      RECT 63.55 -26.77 63.65 -26.235 ;
      RECT 63.55 -25.445 63.65 -24.91 ;
      RECT 63.55 -23.54 63.65 -23.005 ;
      RECT 63.55 -22.215 63.65 -21.68 ;
      RECT 63.55 -20.31 63.65 -19.775 ;
      RECT 63.55 -18.985 63.65 -18.45 ;
      RECT 63.55 -17.08 63.65 -16.545 ;
      RECT 63.55 -15.755 63.65 -15.22 ;
      RECT 63.55 -13.85 63.65 -13.315 ;
      RECT 63.55 -12.525 63.65 -11.99 ;
      RECT 63.55 -10.62 63.65 -10.085 ;
      RECT 63.55 -9.295 63.65 -8.76 ;
      RECT 63.55 -7.39 63.65 -6.855 ;
      RECT 63.55 -6.065 63.65 -5.53 ;
      RECT 63.55 -4.16 63.65 -3.625 ;
      RECT 63.55 -2.835 63.65 -2.3 ;
      RECT 63.55 -0.93 63.65 -0.395 ;
      RECT 63.55 0.395 63.65 0.93 ;
      RECT 63.425 -108.175 63.525 -107.215 ;
      RECT 63.05 -100.19 63.4 -100.07 ;
      RECT 63.05 -96.96 63.4 -96.84 ;
      RECT 63.05 -93.73 63.4 -93.61 ;
      RECT 63.05 -90.5 63.4 -90.38 ;
      RECT 63.05 -87.27 63.4 -87.15 ;
      RECT 63.05 -84.04 63.4 -83.92 ;
      RECT 63.05 -80.81 63.4 -80.69 ;
      RECT 63.05 -77.58 63.4 -77.46 ;
      RECT 63.05 -74.35 63.4 -74.23 ;
      RECT 63.05 -71.12 63.4 -71 ;
      RECT 63.05 -67.89 63.4 -67.77 ;
      RECT 63.05 -64.66 63.4 -64.54 ;
      RECT 63.05 -61.43 63.4 -61.31 ;
      RECT 63.05 -58.2 63.4 -58.08 ;
      RECT 63.05 -54.97 63.4 -54.85 ;
      RECT 63.05 -51.74 63.4 -51.62 ;
      RECT 63.05 -48.51 63.4 -48.39 ;
      RECT 63.05 -45.28 63.4 -45.16 ;
      RECT 63.05 -42.05 63.4 -41.93 ;
      RECT 63.05 -38.82 63.4 -38.7 ;
      RECT 63.05 -35.59 63.4 -35.47 ;
      RECT 63.05 -32.36 63.4 -32.24 ;
      RECT 63.05 -29.13 63.4 -29.01 ;
      RECT 63.05 -25.9 63.4 -25.78 ;
      RECT 63.05 -22.67 63.4 -22.55 ;
      RECT 63.05 -19.44 63.4 -19.32 ;
      RECT 63.05 -16.21 63.4 -16.09 ;
      RECT 63.05 -12.98 63.4 -12.86 ;
      RECT 63.05 -9.75 63.4 -9.63 ;
      RECT 63.05 -6.52 63.4 -6.4 ;
      RECT 63.05 -3.29 63.4 -3.17 ;
      RECT 63.05 -0.06 63.4 0.06 ;
      RECT 63.165 -108.175 63.265 -107.215 ;
      RECT 63.165 2.175 63.265 3.135 ;
      RECT 63.065 -113.555 63.165 -113.085 ;
      RECT 62.565 -100.19 62.915 -100.07 ;
      RECT 62.565 -96.96 62.915 -96.84 ;
      RECT 62.565 -93.73 62.915 -93.61 ;
      RECT 62.565 -90.5 62.915 -90.38 ;
      RECT 62.565 -87.27 62.915 -87.15 ;
      RECT 62.565 -84.04 62.915 -83.92 ;
      RECT 62.565 -80.81 62.915 -80.69 ;
      RECT 62.565 -77.58 62.915 -77.46 ;
      RECT 62.565 -74.35 62.915 -74.23 ;
      RECT 62.565 -71.12 62.915 -71 ;
      RECT 62.565 -67.89 62.915 -67.77 ;
      RECT 62.565 -64.66 62.915 -64.54 ;
      RECT 62.565 -61.43 62.915 -61.31 ;
      RECT 62.565 -58.2 62.915 -58.08 ;
      RECT 62.565 -54.97 62.915 -54.85 ;
      RECT 62.565 -51.74 62.915 -51.62 ;
      RECT 62.565 -48.51 62.915 -48.39 ;
      RECT 62.565 -45.28 62.915 -45.16 ;
      RECT 62.565 -42.05 62.915 -41.93 ;
      RECT 62.565 -38.82 62.915 -38.7 ;
      RECT 62.565 -35.59 62.915 -35.47 ;
      RECT 62.565 -32.36 62.915 -32.24 ;
      RECT 62.565 -29.13 62.915 -29.01 ;
      RECT 62.565 -25.9 62.915 -25.78 ;
      RECT 62.565 -22.67 62.915 -22.55 ;
      RECT 62.565 -19.44 62.915 -19.32 ;
      RECT 62.565 -16.21 62.915 -16.09 ;
      RECT 62.565 -12.98 62.915 -12.86 ;
      RECT 62.565 -9.75 62.915 -9.63 ;
      RECT 62.565 -6.52 62.915 -6.4 ;
      RECT 62.565 -3.29 62.915 -3.17 ;
      RECT 62.565 -0.06 62.915 0.06 ;
      RECT 62.7 -110.735 62.85 -110.445 ;
      RECT 62.735 -108.175 62.835 -107.215 ;
      RECT 62.735 2.175 62.835 3.135 ;
      RECT 62.715 -112.19 62.815 -111.65 ;
      RECT 62.475 -113.555 62.575 -113.085 ;
      RECT 62.475 -108.175 62.575 -107.215 ;
      RECT 62.35 -101.06 62.45 -100.525 ;
      RECT 62.35 -99.735 62.45 -99.2 ;
      RECT 62.35 -97.83 62.45 -97.295 ;
      RECT 62.35 -96.505 62.45 -95.97 ;
      RECT 62.35 -94.6 62.45 -94.065 ;
      RECT 62.35 -93.275 62.45 -92.74 ;
      RECT 62.35 -91.37 62.45 -90.835 ;
      RECT 62.35 -90.045 62.45 -89.51 ;
      RECT 62.35 -88.14 62.45 -87.605 ;
      RECT 62.35 -86.815 62.45 -86.28 ;
      RECT 62.35 -84.91 62.45 -84.375 ;
      RECT 62.35 -83.585 62.45 -83.05 ;
      RECT 62.35 -81.68 62.45 -81.145 ;
      RECT 62.35 -80.355 62.45 -79.82 ;
      RECT 62.35 -78.45 62.45 -77.915 ;
      RECT 62.35 -77.125 62.45 -76.59 ;
      RECT 62.35 -75.22 62.45 -74.685 ;
      RECT 62.35 -73.895 62.45 -73.36 ;
      RECT 62.35 -71.99 62.45 -71.455 ;
      RECT 62.35 -70.665 62.45 -70.13 ;
      RECT 62.35 -68.76 62.45 -68.225 ;
      RECT 62.35 -67.435 62.45 -66.9 ;
      RECT 62.35 -65.53 62.45 -64.995 ;
      RECT 62.35 -64.205 62.45 -63.67 ;
      RECT 62.35 -62.3 62.45 -61.765 ;
      RECT 62.35 -60.975 62.45 -60.44 ;
      RECT 62.35 -59.07 62.45 -58.535 ;
      RECT 62.35 -57.745 62.45 -57.21 ;
      RECT 62.35 -55.84 62.45 -55.305 ;
      RECT 62.35 -54.515 62.45 -53.98 ;
      RECT 62.35 -52.61 62.45 -52.075 ;
      RECT 62.35 -51.285 62.45 -50.75 ;
      RECT 62.35 -49.38 62.45 -48.845 ;
      RECT 62.35 -48.055 62.45 -47.52 ;
      RECT 62.35 -46.15 62.45 -45.615 ;
      RECT 62.35 -44.825 62.45 -44.29 ;
      RECT 62.35 -42.92 62.45 -42.385 ;
      RECT 62.35 -41.595 62.45 -41.06 ;
      RECT 62.35 -39.69 62.45 -39.155 ;
      RECT 62.35 -38.365 62.45 -37.83 ;
      RECT 62.35 -36.46 62.45 -35.925 ;
      RECT 62.35 -35.135 62.45 -34.6 ;
      RECT 62.35 -33.23 62.45 -32.695 ;
      RECT 62.35 -31.905 62.45 -31.37 ;
      RECT 62.35 -30 62.45 -29.465 ;
      RECT 62.35 -28.675 62.45 -28.14 ;
      RECT 62.35 -26.77 62.45 -26.235 ;
      RECT 62.35 -25.445 62.45 -24.91 ;
      RECT 62.35 -23.54 62.45 -23.005 ;
      RECT 62.35 -22.215 62.45 -21.68 ;
      RECT 62.35 -20.31 62.45 -19.775 ;
      RECT 62.35 -18.985 62.45 -18.45 ;
      RECT 62.35 -17.08 62.45 -16.545 ;
      RECT 62.35 -15.755 62.45 -15.22 ;
      RECT 62.35 -13.85 62.45 -13.315 ;
      RECT 62.35 -12.525 62.45 -11.99 ;
      RECT 62.35 -10.62 62.45 -10.085 ;
      RECT 62.35 -9.295 62.45 -8.76 ;
      RECT 62.35 -7.39 62.45 -6.855 ;
      RECT 62.35 -6.065 62.45 -5.53 ;
      RECT 62.35 -4.16 62.45 -3.625 ;
      RECT 62.35 -2.835 62.45 -2.3 ;
      RECT 62.35 -0.93 62.45 -0.395 ;
      RECT 62.35 0.395 62.45 0.93 ;
      RECT 62.225 -104.945 62.325 -103.985 ;
      RECT 61.85 -100.19 62.2 -100.07 ;
      RECT 61.85 -96.96 62.2 -96.84 ;
      RECT 61.85 -93.73 62.2 -93.61 ;
      RECT 61.85 -90.5 62.2 -90.38 ;
      RECT 61.85 -87.27 62.2 -87.15 ;
      RECT 61.85 -84.04 62.2 -83.92 ;
      RECT 61.85 -80.81 62.2 -80.69 ;
      RECT 61.85 -77.58 62.2 -77.46 ;
      RECT 61.85 -74.35 62.2 -74.23 ;
      RECT 61.85 -71.12 62.2 -71 ;
      RECT 61.85 -67.89 62.2 -67.77 ;
      RECT 61.85 -64.66 62.2 -64.54 ;
      RECT 61.85 -61.43 62.2 -61.31 ;
      RECT 61.85 -58.2 62.2 -58.08 ;
      RECT 61.85 -54.97 62.2 -54.85 ;
      RECT 61.85 -51.74 62.2 -51.62 ;
      RECT 61.85 -48.51 62.2 -48.39 ;
      RECT 61.85 -45.28 62.2 -45.16 ;
      RECT 61.85 -42.05 62.2 -41.93 ;
      RECT 61.85 -38.82 62.2 -38.7 ;
      RECT 61.85 -35.59 62.2 -35.47 ;
      RECT 61.85 -32.36 62.2 -32.24 ;
      RECT 61.85 -29.13 62.2 -29.01 ;
      RECT 61.85 -25.9 62.2 -25.78 ;
      RECT 61.85 -22.67 62.2 -22.55 ;
      RECT 61.85 -19.44 62.2 -19.32 ;
      RECT 61.85 -16.21 62.2 -16.09 ;
      RECT 61.85 -12.98 62.2 -12.86 ;
      RECT 61.85 -9.75 62.2 -9.63 ;
      RECT 61.85 -6.52 62.2 -6.4 ;
      RECT 61.85 -3.29 62.2 -3.17 ;
      RECT 61.85 -0.06 62.2 0.06 ;
      RECT 61.965 -104.945 62.065 -103.985 ;
      RECT 61.965 2.175 62.065 3.135 ;
      RECT 61.675 -112.255 61.775 -111.775 ;
      RECT 61.675 -110.765 61.775 -110.295 ;
      RECT 61.365 -100.19 61.715 -100.07 ;
      RECT 61.365 -96.96 61.715 -96.84 ;
      RECT 61.365 -93.73 61.715 -93.61 ;
      RECT 61.365 -90.5 61.715 -90.38 ;
      RECT 61.365 -87.27 61.715 -87.15 ;
      RECT 61.365 -84.04 61.715 -83.92 ;
      RECT 61.365 -80.81 61.715 -80.69 ;
      RECT 61.365 -77.58 61.715 -77.46 ;
      RECT 61.365 -74.35 61.715 -74.23 ;
      RECT 61.365 -71.12 61.715 -71 ;
      RECT 61.365 -67.89 61.715 -67.77 ;
      RECT 61.365 -64.66 61.715 -64.54 ;
      RECT 61.365 -61.43 61.715 -61.31 ;
      RECT 61.365 -58.2 61.715 -58.08 ;
      RECT 61.365 -54.97 61.715 -54.85 ;
      RECT 61.365 -51.74 61.715 -51.62 ;
      RECT 61.365 -48.51 61.715 -48.39 ;
      RECT 61.365 -45.28 61.715 -45.16 ;
      RECT 61.365 -42.05 61.715 -41.93 ;
      RECT 61.365 -38.82 61.715 -38.7 ;
      RECT 61.365 -35.59 61.715 -35.47 ;
      RECT 61.365 -32.36 61.715 -32.24 ;
      RECT 61.365 -29.13 61.715 -29.01 ;
      RECT 61.365 -25.9 61.715 -25.78 ;
      RECT 61.365 -22.67 61.715 -22.55 ;
      RECT 61.365 -19.44 61.715 -19.32 ;
      RECT 61.365 -16.21 61.715 -16.09 ;
      RECT 61.365 -12.98 61.715 -12.86 ;
      RECT 61.365 -9.75 61.715 -9.63 ;
      RECT 61.365 -6.52 61.715 -6.4 ;
      RECT 61.365 -3.29 61.715 -3.17 ;
      RECT 61.365 -0.06 61.715 0.06 ;
      RECT 61.535 -104.945 61.635 -103.985 ;
      RECT 61.535 2.175 61.635 3.135 ;
      RECT 57.635 -108.655 61.415 -108.535 ;
      RECT 61.275 -104.945 61.375 -103.985 ;
      RECT 61.15 -101.06 61.25 -100.525 ;
      RECT 61.15 -99.735 61.25 -99.2 ;
      RECT 61.15 -97.83 61.25 -97.295 ;
      RECT 61.15 -96.505 61.25 -95.97 ;
      RECT 61.15 -94.6 61.25 -94.065 ;
      RECT 61.15 -93.275 61.25 -92.74 ;
      RECT 61.15 -91.37 61.25 -90.835 ;
      RECT 61.15 -90.045 61.25 -89.51 ;
      RECT 61.15 -88.14 61.25 -87.605 ;
      RECT 61.15 -86.815 61.25 -86.28 ;
      RECT 61.15 -84.91 61.25 -84.375 ;
      RECT 61.15 -83.585 61.25 -83.05 ;
      RECT 61.15 -81.68 61.25 -81.145 ;
      RECT 61.15 -80.355 61.25 -79.82 ;
      RECT 61.15 -78.45 61.25 -77.915 ;
      RECT 61.15 -77.125 61.25 -76.59 ;
      RECT 61.15 -75.22 61.25 -74.685 ;
      RECT 61.15 -73.895 61.25 -73.36 ;
      RECT 61.15 -71.99 61.25 -71.455 ;
      RECT 61.15 -70.665 61.25 -70.13 ;
      RECT 61.15 -68.76 61.25 -68.225 ;
      RECT 61.15 -67.435 61.25 -66.9 ;
      RECT 61.15 -65.53 61.25 -64.995 ;
      RECT 61.15 -64.205 61.25 -63.67 ;
      RECT 61.15 -62.3 61.25 -61.765 ;
      RECT 61.15 -60.975 61.25 -60.44 ;
      RECT 61.15 -59.07 61.25 -58.535 ;
      RECT 61.15 -57.745 61.25 -57.21 ;
      RECT 61.15 -55.84 61.25 -55.305 ;
      RECT 61.15 -54.515 61.25 -53.98 ;
      RECT 61.15 -52.61 61.25 -52.075 ;
      RECT 61.15 -51.285 61.25 -50.75 ;
      RECT 61.15 -49.38 61.25 -48.845 ;
      RECT 61.15 -48.055 61.25 -47.52 ;
      RECT 61.15 -46.15 61.25 -45.615 ;
      RECT 61.15 -44.825 61.25 -44.29 ;
      RECT 61.15 -42.92 61.25 -42.385 ;
      RECT 61.15 -41.595 61.25 -41.06 ;
      RECT 61.15 -39.69 61.25 -39.155 ;
      RECT 61.15 -38.365 61.25 -37.83 ;
      RECT 61.15 -36.46 61.25 -35.925 ;
      RECT 61.15 -35.135 61.25 -34.6 ;
      RECT 61.15 -33.23 61.25 -32.695 ;
      RECT 61.15 -31.905 61.25 -31.37 ;
      RECT 61.15 -30 61.25 -29.465 ;
      RECT 61.15 -28.675 61.25 -28.14 ;
      RECT 61.15 -26.77 61.25 -26.235 ;
      RECT 61.15 -25.445 61.25 -24.91 ;
      RECT 61.15 -23.54 61.25 -23.005 ;
      RECT 61.15 -22.215 61.25 -21.68 ;
      RECT 61.15 -20.31 61.25 -19.775 ;
      RECT 61.15 -18.985 61.25 -18.45 ;
      RECT 61.15 -17.08 61.25 -16.545 ;
      RECT 61.15 -15.755 61.25 -15.22 ;
      RECT 61.15 -13.85 61.25 -13.315 ;
      RECT 61.15 -12.525 61.25 -11.99 ;
      RECT 61.15 -10.62 61.25 -10.085 ;
      RECT 61.15 -9.295 61.25 -8.76 ;
      RECT 61.15 -7.39 61.25 -6.855 ;
      RECT 61.15 -6.065 61.25 -5.53 ;
      RECT 61.15 -4.16 61.25 -3.625 ;
      RECT 61.15 -2.835 61.25 -2.3 ;
      RECT 61.15 -0.93 61.25 -0.395 ;
      RECT 61.15 0.395 61.25 0.93 ;
      RECT 61.085 -110.75 61.205 -110.37 ;
      RECT 61.085 -112.245 61.185 -111.775 ;
      RECT 61.025 -104.945 61.125 -103.985 ;
      RECT 60.65 -100.19 61 -100.07 ;
      RECT 60.65 -96.96 61 -96.84 ;
      RECT 60.65 -93.73 61 -93.61 ;
      RECT 60.65 -90.5 61 -90.38 ;
      RECT 60.65 -87.27 61 -87.15 ;
      RECT 60.65 -84.04 61 -83.92 ;
      RECT 60.65 -80.81 61 -80.69 ;
      RECT 60.65 -77.58 61 -77.46 ;
      RECT 60.65 -74.35 61 -74.23 ;
      RECT 60.65 -71.12 61 -71 ;
      RECT 60.65 -67.89 61 -67.77 ;
      RECT 60.65 -64.66 61 -64.54 ;
      RECT 60.65 -61.43 61 -61.31 ;
      RECT 60.65 -58.2 61 -58.08 ;
      RECT 60.65 -54.97 61 -54.85 ;
      RECT 60.65 -51.74 61 -51.62 ;
      RECT 60.65 -48.51 61 -48.39 ;
      RECT 60.65 -45.28 61 -45.16 ;
      RECT 60.65 -42.05 61 -41.93 ;
      RECT 60.65 -38.82 61 -38.7 ;
      RECT 60.65 -35.59 61 -35.47 ;
      RECT 60.65 -32.36 61 -32.24 ;
      RECT 60.65 -29.13 61 -29.01 ;
      RECT 60.65 -25.9 61 -25.78 ;
      RECT 60.65 -22.67 61 -22.55 ;
      RECT 60.65 -19.44 61 -19.32 ;
      RECT 60.65 -16.21 61 -16.09 ;
      RECT 60.65 -12.98 61 -12.86 ;
      RECT 60.65 -9.75 61 -9.63 ;
      RECT 60.65 -6.52 61 -6.4 ;
      RECT 60.65 -3.29 61 -3.17 ;
      RECT 60.65 -0.06 61 0.06 ;
      RECT 60.765 -104.945 60.865 -103.985 ;
      RECT 60.765 2.175 60.865 3.135 ;
      RECT 60.495 -109.595 60.63 -109.275 ;
      RECT 60.165 -100.19 60.515 -100.07 ;
      RECT 60.165 -96.96 60.515 -96.84 ;
      RECT 60.165 -93.73 60.515 -93.61 ;
      RECT 60.165 -90.5 60.515 -90.38 ;
      RECT 60.165 -87.27 60.515 -87.15 ;
      RECT 60.165 -84.04 60.515 -83.92 ;
      RECT 60.165 -80.81 60.515 -80.69 ;
      RECT 60.165 -77.58 60.515 -77.46 ;
      RECT 60.165 -74.35 60.515 -74.23 ;
      RECT 60.165 -71.12 60.515 -71 ;
      RECT 60.165 -67.89 60.515 -67.77 ;
      RECT 60.165 -64.66 60.515 -64.54 ;
      RECT 60.165 -61.43 60.515 -61.31 ;
      RECT 60.165 -58.2 60.515 -58.08 ;
      RECT 60.165 -54.97 60.515 -54.85 ;
      RECT 60.165 -51.74 60.515 -51.62 ;
      RECT 60.165 -48.51 60.515 -48.39 ;
      RECT 60.165 -45.28 60.515 -45.16 ;
      RECT 60.165 -42.05 60.515 -41.93 ;
      RECT 60.165 -38.82 60.515 -38.7 ;
      RECT 60.165 -35.59 60.515 -35.47 ;
      RECT 60.165 -32.36 60.515 -32.24 ;
      RECT 60.165 -29.13 60.515 -29.01 ;
      RECT 60.165 -25.9 60.515 -25.78 ;
      RECT 60.165 -22.67 60.515 -22.55 ;
      RECT 60.165 -19.44 60.515 -19.32 ;
      RECT 60.165 -16.21 60.515 -16.09 ;
      RECT 60.165 -12.98 60.515 -12.86 ;
      RECT 60.165 -9.75 60.515 -9.63 ;
      RECT 60.165 -6.52 60.515 -6.4 ;
      RECT 60.165 -3.29 60.515 -3.17 ;
      RECT 60.165 -0.06 60.515 0.06 ;
      RECT 60.335 -104.945 60.435 -103.985 ;
      RECT 60.335 2.175 60.435 3.135 ;
      RECT 60.16 -109.595 60.305 -109.275 ;
      RECT 60.075 -104.945 60.175 -103.985 ;
      RECT 59.95 -101.06 60.05 -100.525 ;
      RECT 59.95 -99.735 60.05 -99.2 ;
      RECT 59.95 -97.83 60.05 -97.295 ;
      RECT 59.95 -96.505 60.05 -95.97 ;
      RECT 59.95 -94.6 60.05 -94.065 ;
      RECT 59.95 -93.275 60.05 -92.74 ;
      RECT 59.95 -91.37 60.05 -90.835 ;
      RECT 59.95 -90.045 60.05 -89.51 ;
      RECT 59.95 -88.14 60.05 -87.605 ;
      RECT 59.95 -86.815 60.05 -86.28 ;
      RECT 59.95 -84.91 60.05 -84.375 ;
      RECT 59.95 -83.585 60.05 -83.05 ;
      RECT 59.95 -81.68 60.05 -81.145 ;
      RECT 59.95 -80.355 60.05 -79.82 ;
      RECT 59.95 -78.45 60.05 -77.915 ;
      RECT 59.95 -77.125 60.05 -76.59 ;
      RECT 59.95 -75.22 60.05 -74.685 ;
      RECT 59.95 -73.895 60.05 -73.36 ;
      RECT 59.95 -71.99 60.05 -71.455 ;
      RECT 59.95 -70.665 60.05 -70.13 ;
      RECT 59.95 -68.76 60.05 -68.225 ;
      RECT 59.95 -67.435 60.05 -66.9 ;
      RECT 59.95 -65.53 60.05 -64.995 ;
      RECT 59.95 -64.205 60.05 -63.67 ;
      RECT 59.95 -62.3 60.05 -61.765 ;
      RECT 59.95 -60.975 60.05 -60.44 ;
      RECT 59.95 -59.07 60.05 -58.535 ;
      RECT 59.95 -57.745 60.05 -57.21 ;
      RECT 59.95 -55.84 60.05 -55.305 ;
      RECT 59.95 -54.515 60.05 -53.98 ;
      RECT 59.95 -52.61 60.05 -52.075 ;
      RECT 59.95 -51.285 60.05 -50.75 ;
      RECT 59.95 -49.38 60.05 -48.845 ;
      RECT 59.95 -48.055 60.05 -47.52 ;
      RECT 59.95 -46.15 60.05 -45.615 ;
      RECT 59.95 -44.825 60.05 -44.29 ;
      RECT 59.95 -42.92 60.05 -42.385 ;
      RECT 59.95 -41.595 60.05 -41.06 ;
      RECT 59.95 -39.69 60.05 -39.155 ;
      RECT 59.95 -38.365 60.05 -37.83 ;
      RECT 59.95 -36.46 60.05 -35.925 ;
      RECT 59.95 -35.135 60.05 -34.6 ;
      RECT 59.95 -33.23 60.05 -32.695 ;
      RECT 59.95 -31.905 60.05 -31.37 ;
      RECT 59.95 -30 60.05 -29.465 ;
      RECT 59.95 -28.675 60.05 -28.14 ;
      RECT 59.95 -26.77 60.05 -26.235 ;
      RECT 59.95 -25.445 60.05 -24.91 ;
      RECT 59.95 -23.54 60.05 -23.005 ;
      RECT 59.95 -22.215 60.05 -21.68 ;
      RECT 59.95 -20.31 60.05 -19.775 ;
      RECT 59.95 -18.985 60.05 -18.45 ;
      RECT 59.95 -17.08 60.05 -16.545 ;
      RECT 59.95 -15.755 60.05 -15.22 ;
      RECT 59.95 -13.85 60.05 -13.315 ;
      RECT 59.95 -12.525 60.05 -11.99 ;
      RECT 59.95 -10.62 60.05 -10.085 ;
      RECT 59.95 -9.295 60.05 -8.76 ;
      RECT 59.95 -7.39 60.05 -6.855 ;
      RECT 59.95 -6.065 60.05 -5.53 ;
      RECT 59.95 -4.16 60.05 -3.625 ;
      RECT 59.95 -2.835 60.05 -2.3 ;
      RECT 59.95 -0.93 60.05 -0.395 ;
      RECT 59.95 0.395 60.05 0.93 ;
      RECT 59.825 -108.175 59.925 -107.215 ;
      RECT 59.45 -100.19 59.8 -100.07 ;
      RECT 59.45 -96.96 59.8 -96.84 ;
      RECT 59.45 -93.73 59.8 -93.61 ;
      RECT 59.45 -90.5 59.8 -90.38 ;
      RECT 59.45 -87.27 59.8 -87.15 ;
      RECT 59.45 -84.04 59.8 -83.92 ;
      RECT 59.45 -80.81 59.8 -80.69 ;
      RECT 59.45 -77.58 59.8 -77.46 ;
      RECT 59.45 -74.35 59.8 -74.23 ;
      RECT 59.45 -71.12 59.8 -71 ;
      RECT 59.45 -67.89 59.8 -67.77 ;
      RECT 59.45 -64.66 59.8 -64.54 ;
      RECT 59.45 -61.43 59.8 -61.31 ;
      RECT 59.45 -58.2 59.8 -58.08 ;
      RECT 59.45 -54.97 59.8 -54.85 ;
      RECT 59.45 -51.74 59.8 -51.62 ;
      RECT 59.45 -48.51 59.8 -48.39 ;
      RECT 59.45 -45.28 59.8 -45.16 ;
      RECT 59.45 -42.05 59.8 -41.93 ;
      RECT 59.45 -38.82 59.8 -38.7 ;
      RECT 59.45 -35.59 59.8 -35.47 ;
      RECT 59.45 -32.36 59.8 -32.24 ;
      RECT 59.45 -29.13 59.8 -29.01 ;
      RECT 59.45 -25.9 59.8 -25.78 ;
      RECT 59.45 -22.67 59.8 -22.55 ;
      RECT 59.45 -19.44 59.8 -19.32 ;
      RECT 59.45 -16.21 59.8 -16.09 ;
      RECT 59.45 -12.98 59.8 -12.86 ;
      RECT 59.45 -9.75 59.8 -9.63 ;
      RECT 59.45 -6.52 59.8 -6.4 ;
      RECT 59.45 -3.29 59.8 -3.17 ;
      RECT 59.45 -0.06 59.8 0.06 ;
      RECT 59.655 -112.255 59.755 -111.775 ;
      RECT 59.655 -110.765 59.755 -110.295 ;
      RECT 59.565 -108.175 59.665 -107.215 ;
      RECT 59.565 2.175 59.665 3.135 ;
      RECT 58.965 -100.19 59.315 -100.07 ;
      RECT 58.965 -96.96 59.315 -96.84 ;
      RECT 58.965 -93.73 59.315 -93.61 ;
      RECT 58.965 -90.5 59.315 -90.38 ;
      RECT 58.965 -87.27 59.315 -87.15 ;
      RECT 58.965 -84.04 59.315 -83.92 ;
      RECT 58.965 -80.81 59.315 -80.69 ;
      RECT 58.965 -77.58 59.315 -77.46 ;
      RECT 58.965 -74.35 59.315 -74.23 ;
      RECT 58.965 -71.12 59.315 -71 ;
      RECT 58.965 -67.89 59.315 -67.77 ;
      RECT 58.965 -64.66 59.315 -64.54 ;
      RECT 58.965 -61.43 59.315 -61.31 ;
      RECT 58.965 -58.2 59.315 -58.08 ;
      RECT 58.965 -54.97 59.315 -54.85 ;
      RECT 58.965 -51.74 59.315 -51.62 ;
      RECT 58.965 -48.51 59.315 -48.39 ;
      RECT 58.965 -45.28 59.315 -45.16 ;
      RECT 58.965 -42.05 59.315 -41.93 ;
      RECT 58.965 -38.82 59.315 -38.7 ;
      RECT 58.965 -35.59 59.315 -35.47 ;
      RECT 58.965 -32.36 59.315 -32.24 ;
      RECT 58.965 -29.13 59.315 -29.01 ;
      RECT 58.965 -25.9 59.315 -25.78 ;
      RECT 58.965 -22.67 59.315 -22.55 ;
      RECT 58.965 -19.44 59.315 -19.32 ;
      RECT 58.965 -16.21 59.315 -16.09 ;
      RECT 58.965 -12.98 59.315 -12.86 ;
      RECT 58.965 -9.75 59.315 -9.63 ;
      RECT 58.965 -6.52 59.315 -6.4 ;
      RECT 58.965 -3.29 59.315 -3.17 ;
      RECT 58.965 -0.06 59.315 0.06 ;
      RECT 59.135 -108.175 59.235 -107.215 ;
      RECT 59.135 2.175 59.235 3.135 ;
      RECT 59.03 -110.765 59.2 -110.385 ;
      RECT 59.065 -112.245 59.165 -111.775 ;
      RECT 58.875 -108.175 58.975 -107.215 ;
      RECT 58.75 -101.06 58.85 -100.525 ;
      RECT 58.75 -99.735 58.85 -99.2 ;
      RECT 58.75 -97.83 58.85 -97.295 ;
      RECT 58.75 -96.505 58.85 -95.97 ;
      RECT 58.75 -94.6 58.85 -94.065 ;
      RECT 58.75 -93.275 58.85 -92.74 ;
      RECT 58.75 -91.37 58.85 -90.835 ;
      RECT 58.75 -90.045 58.85 -89.51 ;
      RECT 58.75 -88.14 58.85 -87.605 ;
      RECT 58.75 -86.815 58.85 -86.28 ;
      RECT 58.75 -84.91 58.85 -84.375 ;
      RECT 58.75 -83.585 58.85 -83.05 ;
      RECT 58.75 -81.68 58.85 -81.145 ;
      RECT 58.75 -80.355 58.85 -79.82 ;
      RECT 58.75 -78.45 58.85 -77.915 ;
      RECT 58.75 -77.125 58.85 -76.59 ;
      RECT 58.75 -75.22 58.85 -74.685 ;
      RECT 58.75 -73.895 58.85 -73.36 ;
      RECT 58.75 -71.99 58.85 -71.455 ;
      RECT 58.75 -70.665 58.85 -70.13 ;
      RECT 58.75 -68.76 58.85 -68.225 ;
      RECT 58.75 -67.435 58.85 -66.9 ;
      RECT 58.75 -65.53 58.85 -64.995 ;
      RECT 58.75 -64.205 58.85 -63.67 ;
      RECT 58.75 -62.3 58.85 -61.765 ;
      RECT 58.75 -60.975 58.85 -60.44 ;
      RECT 58.75 -59.07 58.85 -58.535 ;
      RECT 58.75 -57.745 58.85 -57.21 ;
      RECT 58.75 -55.84 58.85 -55.305 ;
      RECT 58.75 -54.515 58.85 -53.98 ;
      RECT 58.75 -52.61 58.85 -52.075 ;
      RECT 58.75 -51.285 58.85 -50.75 ;
      RECT 58.75 -49.38 58.85 -48.845 ;
      RECT 58.75 -48.055 58.85 -47.52 ;
      RECT 58.75 -46.15 58.85 -45.615 ;
      RECT 58.75 -44.825 58.85 -44.29 ;
      RECT 58.75 -42.92 58.85 -42.385 ;
      RECT 58.75 -41.595 58.85 -41.06 ;
      RECT 58.75 -39.69 58.85 -39.155 ;
      RECT 58.75 -38.365 58.85 -37.83 ;
      RECT 58.75 -36.46 58.85 -35.925 ;
      RECT 58.75 -35.135 58.85 -34.6 ;
      RECT 58.75 -33.23 58.85 -32.695 ;
      RECT 58.75 -31.905 58.85 -31.37 ;
      RECT 58.75 -30 58.85 -29.465 ;
      RECT 58.75 -28.675 58.85 -28.14 ;
      RECT 58.75 -26.77 58.85 -26.235 ;
      RECT 58.75 -25.445 58.85 -24.91 ;
      RECT 58.75 -23.54 58.85 -23.005 ;
      RECT 58.75 -22.215 58.85 -21.68 ;
      RECT 58.75 -20.31 58.85 -19.775 ;
      RECT 58.75 -18.985 58.85 -18.45 ;
      RECT 58.75 -17.08 58.85 -16.545 ;
      RECT 58.75 -15.755 58.85 -15.22 ;
      RECT 58.75 -13.85 58.85 -13.315 ;
      RECT 58.75 -12.525 58.85 -11.99 ;
      RECT 58.75 -10.62 58.85 -10.085 ;
      RECT 58.75 -9.295 58.85 -8.76 ;
      RECT 58.75 -7.39 58.85 -6.855 ;
      RECT 58.75 -6.065 58.85 -5.53 ;
      RECT 58.75 -4.16 58.85 -3.625 ;
      RECT 58.75 -2.835 58.85 -2.3 ;
      RECT 58.75 -0.93 58.85 -0.395 ;
      RECT 58.75 0.395 58.85 0.93 ;
      RECT 58.625 -108.175 58.725 -107.215 ;
      RECT 58.25 -100.19 58.6 -100.07 ;
      RECT 58.25 -96.96 58.6 -96.84 ;
      RECT 58.25 -93.73 58.6 -93.61 ;
      RECT 58.25 -90.5 58.6 -90.38 ;
      RECT 58.25 -87.27 58.6 -87.15 ;
      RECT 58.25 -84.04 58.6 -83.92 ;
      RECT 58.25 -80.81 58.6 -80.69 ;
      RECT 58.25 -77.58 58.6 -77.46 ;
      RECT 58.25 -74.35 58.6 -74.23 ;
      RECT 58.25 -71.12 58.6 -71 ;
      RECT 58.25 -67.89 58.6 -67.77 ;
      RECT 58.25 -64.66 58.6 -64.54 ;
      RECT 58.25 -61.43 58.6 -61.31 ;
      RECT 58.25 -58.2 58.6 -58.08 ;
      RECT 58.25 -54.97 58.6 -54.85 ;
      RECT 58.25 -51.74 58.6 -51.62 ;
      RECT 58.25 -48.51 58.6 -48.39 ;
      RECT 58.25 -45.28 58.6 -45.16 ;
      RECT 58.25 -42.05 58.6 -41.93 ;
      RECT 58.25 -38.82 58.6 -38.7 ;
      RECT 58.25 -35.59 58.6 -35.47 ;
      RECT 58.25 -32.36 58.6 -32.24 ;
      RECT 58.25 -29.13 58.6 -29.01 ;
      RECT 58.25 -25.9 58.6 -25.78 ;
      RECT 58.25 -22.67 58.6 -22.55 ;
      RECT 58.25 -19.44 58.6 -19.32 ;
      RECT 58.25 -16.21 58.6 -16.09 ;
      RECT 58.25 -12.98 58.6 -12.86 ;
      RECT 58.25 -9.75 58.6 -9.63 ;
      RECT 58.25 -6.52 58.6 -6.4 ;
      RECT 58.25 -3.29 58.6 -3.17 ;
      RECT 58.25 -0.06 58.6 0.06 ;
      RECT 58.365 -108.175 58.465 -107.215 ;
      RECT 58.365 2.175 58.465 3.135 ;
      RECT 58.265 -113.555 58.365 -113.085 ;
      RECT 57.765 -100.19 58.115 -100.07 ;
      RECT 57.765 -96.96 58.115 -96.84 ;
      RECT 57.765 -93.73 58.115 -93.61 ;
      RECT 57.765 -90.5 58.115 -90.38 ;
      RECT 57.765 -87.27 58.115 -87.15 ;
      RECT 57.765 -84.04 58.115 -83.92 ;
      RECT 57.765 -80.81 58.115 -80.69 ;
      RECT 57.765 -77.58 58.115 -77.46 ;
      RECT 57.765 -74.35 58.115 -74.23 ;
      RECT 57.765 -71.12 58.115 -71 ;
      RECT 57.765 -67.89 58.115 -67.77 ;
      RECT 57.765 -64.66 58.115 -64.54 ;
      RECT 57.765 -61.43 58.115 -61.31 ;
      RECT 57.765 -58.2 58.115 -58.08 ;
      RECT 57.765 -54.97 58.115 -54.85 ;
      RECT 57.765 -51.74 58.115 -51.62 ;
      RECT 57.765 -48.51 58.115 -48.39 ;
      RECT 57.765 -45.28 58.115 -45.16 ;
      RECT 57.765 -42.05 58.115 -41.93 ;
      RECT 57.765 -38.82 58.115 -38.7 ;
      RECT 57.765 -35.59 58.115 -35.47 ;
      RECT 57.765 -32.36 58.115 -32.24 ;
      RECT 57.765 -29.13 58.115 -29.01 ;
      RECT 57.765 -25.9 58.115 -25.78 ;
      RECT 57.765 -22.67 58.115 -22.55 ;
      RECT 57.765 -19.44 58.115 -19.32 ;
      RECT 57.765 -16.21 58.115 -16.09 ;
      RECT 57.765 -12.98 58.115 -12.86 ;
      RECT 57.765 -9.75 58.115 -9.63 ;
      RECT 57.765 -6.52 58.115 -6.4 ;
      RECT 57.765 -3.29 58.115 -3.17 ;
      RECT 57.765 -0.06 58.115 0.06 ;
      RECT 57.9 -110.735 58.05 -110.445 ;
      RECT 57.935 -108.175 58.035 -107.215 ;
      RECT 57.935 2.175 58.035 3.135 ;
      RECT 57.915 -112.19 58.015 -111.65 ;
      RECT 57.675 -113.555 57.775 -113.085 ;
      RECT 57.675 -108.175 57.775 -107.215 ;
      RECT 57.55 -101.06 57.65 -100.525 ;
      RECT 57.55 -99.735 57.65 -99.2 ;
      RECT 57.55 -97.83 57.65 -97.295 ;
      RECT 57.55 -96.505 57.65 -95.97 ;
      RECT 57.55 -94.6 57.65 -94.065 ;
      RECT 57.55 -93.275 57.65 -92.74 ;
      RECT 57.55 -91.37 57.65 -90.835 ;
      RECT 57.55 -90.045 57.65 -89.51 ;
      RECT 57.55 -88.14 57.65 -87.605 ;
      RECT 57.55 -86.815 57.65 -86.28 ;
      RECT 57.55 -84.91 57.65 -84.375 ;
      RECT 57.55 -83.585 57.65 -83.05 ;
      RECT 57.55 -81.68 57.65 -81.145 ;
      RECT 57.55 -80.355 57.65 -79.82 ;
      RECT 57.55 -78.45 57.65 -77.915 ;
      RECT 57.55 -77.125 57.65 -76.59 ;
      RECT 57.55 -75.22 57.65 -74.685 ;
      RECT 57.55 -73.895 57.65 -73.36 ;
      RECT 57.55 -71.99 57.65 -71.455 ;
      RECT 57.55 -70.665 57.65 -70.13 ;
      RECT 57.55 -68.76 57.65 -68.225 ;
      RECT 57.55 -67.435 57.65 -66.9 ;
      RECT 57.55 -65.53 57.65 -64.995 ;
      RECT 57.55 -64.205 57.65 -63.67 ;
      RECT 57.55 -62.3 57.65 -61.765 ;
      RECT 57.55 -60.975 57.65 -60.44 ;
      RECT 57.55 -59.07 57.65 -58.535 ;
      RECT 57.55 -57.745 57.65 -57.21 ;
      RECT 57.55 -55.84 57.65 -55.305 ;
      RECT 57.55 -54.515 57.65 -53.98 ;
      RECT 57.55 -52.61 57.65 -52.075 ;
      RECT 57.55 -51.285 57.65 -50.75 ;
      RECT 57.55 -49.38 57.65 -48.845 ;
      RECT 57.55 -48.055 57.65 -47.52 ;
      RECT 57.55 -46.15 57.65 -45.615 ;
      RECT 57.55 -44.825 57.65 -44.29 ;
      RECT 57.55 -42.92 57.65 -42.385 ;
      RECT 57.55 -41.595 57.65 -41.06 ;
      RECT 57.55 -39.69 57.65 -39.155 ;
      RECT 57.55 -38.365 57.65 -37.83 ;
      RECT 57.55 -36.46 57.65 -35.925 ;
      RECT 57.55 -35.135 57.65 -34.6 ;
      RECT 57.55 -33.23 57.65 -32.695 ;
      RECT 57.55 -31.905 57.65 -31.37 ;
      RECT 57.55 -30 57.65 -29.465 ;
      RECT 57.55 -28.675 57.65 -28.14 ;
      RECT 57.55 -26.77 57.65 -26.235 ;
      RECT 57.55 -25.445 57.65 -24.91 ;
      RECT 57.55 -23.54 57.65 -23.005 ;
      RECT 57.55 -22.215 57.65 -21.68 ;
      RECT 57.55 -20.31 57.65 -19.775 ;
      RECT 57.55 -18.985 57.65 -18.45 ;
      RECT 57.55 -17.08 57.65 -16.545 ;
      RECT 57.55 -15.755 57.65 -15.22 ;
      RECT 57.55 -13.85 57.65 -13.315 ;
      RECT 57.55 -12.525 57.65 -11.99 ;
      RECT 57.55 -10.62 57.65 -10.085 ;
      RECT 57.55 -9.295 57.65 -8.76 ;
      RECT 57.55 -7.39 57.65 -6.855 ;
      RECT 57.55 -6.065 57.65 -5.53 ;
      RECT 57.55 -4.16 57.65 -3.625 ;
      RECT 57.55 -2.835 57.65 -2.3 ;
      RECT 57.55 -0.93 57.65 -0.395 ;
      RECT 57.55 0.395 57.65 0.93 ;
      RECT 57.425 -104.945 57.525 -103.985 ;
      RECT 57.05 -100.19 57.4 -100.07 ;
      RECT 57.05 -96.96 57.4 -96.84 ;
      RECT 57.05 -93.73 57.4 -93.61 ;
      RECT 57.05 -90.5 57.4 -90.38 ;
      RECT 57.05 -87.27 57.4 -87.15 ;
      RECT 57.05 -84.04 57.4 -83.92 ;
      RECT 57.05 -80.81 57.4 -80.69 ;
      RECT 57.05 -77.58 57.4 -77.46 ;
      RECT 57.05 -74.35 57.4 -74.23 ;
      RECT 57.05 -71.12 57.4 -71 ;
      RECT 57.05 -67.89 57.4 -67.77 ;
      RECT 57.05 -64.66 57.4 -64.54 ;
      RECT 57.05 -61.43 57.4 -61.31 ;
      RECT 57.05 -58.2 57.4 -58.08 ;
      RECT 57.05 -54.97 57.4 -54.85 ;
      RECT 57.05 -51.74 57.4 -51.62 ;
      RECT 57.05 -48.51 57.4 -48.39 ;
      RECT 57.05 -45.28 57.4 -45.16 ;
      RECT 57.05 -42.05 57.4 -41.93 ;
      RECT 57.05 -38.82 57.4 -38.7 ;
      RECT 57.05 -35.59 57.4 -35.47 ;
      RECT 57.05 -32.36 57.4 -32.24 ;
      RECT 57.05 -29.13 57.4 -29.01 ;
      RECT 57.05 -25.9 57.4 -25.78 ;
      RECT 57.05 -22.67 57.4 -22.55 ;
      RECT 57.05 -19.44 57.4 -19.32 ;
      RECT 57.05 -16.21 57.4 -16.09 ;
      RECT 57.05 -12.98 57.4 -12.86 ;
      RECT 57.05 -9.75 57.4 -9.63 ;
      RECT 57.05 -6.52 57.4 -6.4 ;
      RECT 57.05 -3.29 57.4 -3.17 ;
      RECT 57.05 -0.06 57.4 0.06 ;
      RECT 57.165 -104.945 57.265 -103.985 ;
      RECT 57.165 2.175 57.265 3.135 ;
      RECT 56.875 -112.255 56.975 -111.775 ;
      RECT 56.875 -110.765 56.975 -110.295 ;
      RECT 56.565 -100.19 56.915 -100.07 ;
      RECT 56.565 -96.96 56.915 -96.84 ;
      RECT 56.565 -93.73 56.915 -93.61 ;
      RECT 56.565 -90.5 56.915 -90.38 ;
      RECT 56.565 -87.27 56.915 -87.15 ;
      RECT 56.565 -84.04 56.915 -83.92 ;
      RECT 56.565 -80.81 56.915 -80.69 ;
      RECT 56.565 -77.58 56.915 -77.46 ;
      RECT 56.565 -74.35 56.915 -74.23 ;
      RECT 56.565 -71.12 56.915 -71 ;
      RECT 56.565 -67.89 56.915 -67.77 ;
      RECT 56.565 -64.66 56.915 -64.54 ;
      RECT 56.565 -61.43 56.915 -61.31 ;
      RECT 56.565 -58.2 56.915 -58.08 ;
      RECT 56.565 -54.97 56.915 -54.85 ;
      RECT 56.565 -51.74 56.915 -51.62 ;
      RECT 56.565 -48.51 56.915 -48.39 ;
      RECT 56.565 -45.28 56.915 -45.16 ;
      RECT 56.565 -42.05 56.915 -41.93 ;
      RECT 56.565 -38.82 56.915 -38.7 ;
      RECT 56.565 -35.59 56.915 -35.47 ;
      RECT 56.565 -32.36 56.915 -32.24 ;
      RECT 56.565 -29.13 56.915 -29.01 ;
      RECT 56.565 -25.9 56.915 -25.78 ;
      RECT 56.565 -22.67 56.915 -22.55 ;
      RECT 56.565 -19.44 56.915 -19.32 ;
      RECT 56.565 -16.21 56.915 -16.09 ;
      RECT 56.565 -12.98 56.915 -12.86 ;
      RECT 56.565 -9.75 56.915 -9.63 ;
      RECT 56.565 -6.52 56.915 -6.4 ;
      RECT 56.565 -3.29 56.915 -3.17 ;
      RECT 56.565 -0.06 56.915 0.06 ;
      RECT 56.735 -104.945 56.835 -103.985 ;
      RECT 56.735 2.175 56.835 3.135 ;
      RECT 52.835 -108.655 56.615 -108.535 ;
      RECT 56.475 -104.945 56.575 -103.985 ;
      RECT 56.35 -101.06 56.45 -100.525 ;
      RECT 56.35 -99.735 56.45 -99.2 ;
      RECT 56.35 -97.83 56.45 -97.295 ;
      RECT 56.35 -96.505 56.45 -95.97 ;
      RECT 56.35 -94.6 56.45 -94.065 ;
      RECT 56.35 -93.275 56.45 -92.74 ;
      RECT 56.35 -91.37 56.45 -90.835 ;
      RECT 56.35 -90.045 56.45 -89.51 ;
      RECT 56.35 -88.14 56.45 -87.605 ;
      RECT 56.35 -86.815 56.45 -86.28 ;
      RECT 56.35 -84.91 56.45 -84.375 ;
      RECT 56.35 -83.585 56.45 -83.05 ;
      RECT 56.35 -81.68 56.45 -81.145 ;
      RECT 56.35 -80.355 56.45 -79.82 ;
      RECT 56.35 -78.45 56.45 -77.915 ;
      RECT 56.35 -77.125 56.45 -76.59 ;
      RECT 56.35 -75.22 56.45 -74.685 ;
      RECT 56.35 -73.895 56.45 -73.36 ;
      RECT 56.35 -71.99 56.45 -71.455 ;
      RECT 56.35 -70.665 56.45 -70.13 ;
      RECT 56.35 -68.76 56.45 -68.225 ;
      RECT 56.35 -67.435 56.45 -66.9 ;
      RECT 56.35 -65.53 56.45 -64.995 ;
      RECT 56.35 -64.205 56.45 -63.67 ;
      RECT 56.35 -62.3 56.45 -61.765 ;
      RECT 56.35 -60.975 56.45 -60.44 ;
      RECT 56.35 -59.07 56.45 -58.535 ;
      RECT 56.35 -57.745 56.45 -57.21 ;
      RECT 56.35 -55.84 56.45 -55.305 ;
      RECT 56.35 -54.515 56.45 -53.98 ;
      RECT 56.35 -52.61 56.45 -52.075 ;
      RECT 56.35 -51.285 56.45 -50.75 ;
      RECT 56.35 -49.38 56.45 -48.845 ;
      RECT 56.35 -48.055 56.45 -47.52 ;
      RECT 56.35 -46.15 56.45 -45.615 ;
      RECT 56.35 -44.825 56.45 -44.29 ;
      RECT 56.35 -42.92 56.45 -42.385 ;
      RECT 56.35 -41.595 56.45 -41.06 ;
      RECT 56.35 -39.69 56.45 -39.155 ;
      RECT 56.35 -38.365 56.45 -37.83 ;
      RECT 56.35 -36.46 56.45 -35.925 ;
      RECT 56.35 -35.135 56.45 -34.6 ;
      RECT 56.35 -33.23 56.45 -32.695 ;
      RECT 56.35 -31.905 56.45 -31.37 ;
      RECT 56.35 -30 56.45 -29.465 ;
      RECT 56.35 -28.675 56.45 -28.14 ;
      RECT 56.35 -26.77 56.45 -26.235 ;
      RECT 56.35 -25.445 56.45 -24.91 ;
      RECT 56.35 -23.54 56.45 -23.005 ;
      RECT 56.35 -22.215 56.45 -21.68 ;
      RECT 56.35 -20.31 56.45 -19.775 ;
      RECT 56.35 -18.985 56.45 -18.45 ;
      RECT 56.35 -17.08 56.45 -16.545 ;
      RECT 56.35 -15.755 56.45 -15.22 ;
      RECT 56.35 -13.85 56.45 -13.315 ;
      RECT 56.35 -12.525 56.45 -11.99 ;
      RECT 56.35 -10.62 56.45 -10.085 ;
      RECT 56.35 -9.295 56.45 -8.76 ;
      RECT 56.35 -7.39 56.45 -6.855 ;
      RECT 56.35 -6.065 56.45 -5.53 ;
      RECT 56.35 -4.16 56.45 -3.625 ;
      RECT 56.35 -2.835 56.45 -2.3 ;
      RECT 56.35 -0.93 56.45 -0.395 ;
      RECT 56.35 0.395 56.45 0.93 ;
      RECT 56.285 -110.75 56.405 -110.37 ;
      RECT 56.285 -112.245 56.385 -111.775 ;
      RECT 56.225 -104.945 56.325 -103.985 ;
      RECT 55.85 -100.19 56.2 -100.07 ;
      RECT 55.85 -96.96 56.2 -96.84 ;
      RECT 55.85 -93.73 56.2 -93.61 ;
      RECT 55.85 -90.5 56.2 -90.38 ;
      RECT 55.85 -87.27 56.2 -87.15 ;
      RECT 55.85 -84.04 56.2 -83.92 ;
      RECT 55.85 -80.81 56.2 -80.69 ;
      RECT 55.85 -77.58 56.2 -77.46 ;
      RECT 55.85 -74.35 56.2 -74.23 ;
      RECT 55.85 -71.12 56.2 -71 ;
      RECT 55.85 -67.89 56.2 -67.77 ;
      RECT 55.85 -64.66 56.2 -64.54 ;
      RECT 55.85 -61.43 56.2 -61.31 ;
      RECT 55.85 -58.2 56.2 -58.08 ;
      RECT 55.85 -54.97 56.2 -54.85 ;
      RECT 55.85 -51.74 56.2 -51.62 ;
      RECT 55.85 -48.51 56.2 -48.39 ;
      RECT 55.85 -45.28 56.2 -45.16 ;
      RECT 55.85 -42.05 56.2 -41.93 ;
      RECT 55.85 -38.82 56.2 -38.7 ;
      RECT 55.85 -35.59 56.2 -35.47 ;
      RECT 55.85 -32.36 56.2 -32.24 ;
      RECT 55.85 -29.13 56.2 -29.01 ;
      RECT 55.85 -25.9 56.2 -25.78 ;
      RECT 55.85 -22.67 56.2 -22.55 ;
      RECT 55.85 -19.44 56.2 -19.32 ;
      RECT 55.85 -16.21 56.2 -16.09 ;
      RECT 55.85 -12.98 56.2 -12.86 ;
      RECT 55.85 -9.75 56.2 -9.63 ;
      RECT 55.85 -6.52 56.2 -6.4 ;
      RECT 55.85 -3.29 56.2 -3.17 ;
      RECT 55.85 -0.06 56.2 0.06 ;
      RECT 55.965 -104.945 56.065 -103.985 ;
      RECT 55.965 2.175 56.065 3.135 ;
      RECT 55.695 -109.595 55.83 -109.275 ;
      RECT 55.365 -100.19 55.715 -100.07 ;
      RECT 55.365 -96.96 55.715 -96.84 ;
      RECT 55.365 -93.73 55.715 -93.61 ;
      RECT 55.365 -90.5 55.715 -90.38 ;
      RECT 55.365 -87.27 55.715 -87.15 ;
      RECT 55.365 -84.04 55.715 -83.92 ;
      RECT 55.365 -80.81 55.715 -80.69 ;
      RECT 55.365 -77.58 55.715 -77.46 ;
      RECT 55.365 -74.35 55.715 -74.23 ;
      RECT 55.365 -71.12 55.715 -71 ;
      RECT 55.365 -67.89 55.715 -67.77 ;
      RECT 55.365 -64.66 55.715 -64.54 ;
      RECT 55.365 -61.43 55.715 -61.31 ;
      RECT 55.365 -58.2 55.715 -58.08 ;
      RECT 55.365 -54.97 55.715 -54.85 ;
      RECT 55.365 -51.74 55.715 -51.62 ;
      RECT 55.365 -48.51 55.715 -48.39 ;
      RECT 55.365 -45.28 55.715 -45.16 ;
      RECT 55.365 -42.05 55.715 -41.93 ;
      RECT 55.365 -38.82 55.715 -38.7 ;
      RECT 55.365 -35.59 55.715 -35.47 ;
      RECT 55.365 -32.36 55.715 -32.24 ;
      RECT 55.365 -29.13 55.715 -29.01 ;
      RECT 55.365 -25.9 55.715 -25.78 ;
      RECT 55.365 -22.67 55.715 -22.55 ;
      RECT 55.365 -19.44 55.715 -19.32 ;
      RECT 55.365 -16.21 55.715 -16.09 ;
      RECT 55.365 -12.98 55.715 -12.86 ;
      RECT 55.365 -9.75 55.715 -9.63 ;
      RECT 55.365 -6.52 55.715 -6.4 ;
      RECT 55.365 -3.29 55.715 -3.17 ;
      RECT 55.365 -0.06 55.715 0.06 ;
      RECT 55.535 -104.945 55.635 -103.985 ;
      RECT 55.535 2.175 55.635 3.135 ;
      RECT 55.36 -109.595 55.505 -109.275 ;
      RECT 55.275 -104.945 55.375 -103.985 ;
      RECT 55.15 -101.06 55.25 -100.525 ;
      RECT 55.15 -99.735 55.25 -99.2 ;
      RECT 55.15 -97.83 55.25 -97.295 ;
      RECT 55.15 -96.505 55.25 -95.97 ;
      RECT 55.15 -94.6 55.25 -94.065 ;
      RECT 55.15 -93.275 55.25 -92.74 ;
      RECT 55.15 -91.37 55.25 -90.835 ;
      RECT 55.15 -90.045 55.25 -89.51 ;
      RECT 55.15 -88.14 55.25 -87.605 ;
      RECT 55.15 -86.815 55.25 -86.28 ;
      RECT 55.15 -84.91 55.25 -84.375 ;
      RECT 55.15 -83.585 55.25 -83.05 ;
      RECT 55.15 -81.68 55.25 -81.145 ;
      RECT 55.15 -80.355 55.25 -79.82 ;
      RECT 55.15 -78.45 55.25 -77.915 ;
      RECT 55.15 -77.125 55.25 -76.59 ;
      RECT 55.15 -75.22 55.25 -74.685 ;
      RECT 55.15 -73.895 55.25 -73.36 ;
      RECT 55.15 -71.99 55.25 -71.455 ;
      RECT 55.15 -70.665 55.25 -70.13 ;
      RECT 55.15 -68.76 55.25 -68.225 ;
      RECT 55.15 -67.435 55.25 -66.9 ;
      RECT 55.15 -65.53 55.25 -64.995 ;
      RECT 55.15 -64.205 55.25 -63.67 ;
      RECT 55.15 -62.3 55.25 -61.765 ;
      RECT 55.15 -60.975 55.25 -60.44 ;
      RECT 55.15 -59.07 55.25 -58.535 ;
      RECT 55.15 -57.745 55.25 -57.21 ;
      RECT 55.15 -55.84 55.25 -55.305 ;
      RECT 55.15 -54.515 55.25 -53.98 ;
      RECT 55.15 -52.61 55.25 -52.075 ;
      RECT 55.15 -51.285 55.25 -50.75 ;
      RECT 55.15 -49.38 55.25 -48.845 ;
      RECT 55.15 -48.055 55.25 -47.52 ;
      RECT 55.15 -46.15 55.25 -45.615 ;
      RECT 55.15 -44.825 55.25 -44.29 ;
      RECT 55.15 -42.92 55.25 -42.385 ;
      RECT 55.15 -41.595 55.25 -41.06 ;
      RECT 55.15 -39.69 55.25 -39.155 ;
      RECT 55.15 -38.365 55.25 -37.83 ;
      RECT 55.15 -36.46 55.25 -35.925 ;
      RECT 55.15 -35.135 55.25 -34.6 ;
      RECT 55.15 -33.23 55.25 -32.695 ;
      RECT 55.15 -31.905 55.25 -31.37 ;
      RECT 55.15 -30 55.25 -29.465 ;
      RECT 55.15 -28.675 55.25 -28.14 ;
      RECT 55.15 -26.77 55.25 -26.235 ;
      RECT 55.15 -25.445 55.25 -24.91 ;
      RECT 55.15 -23.54 55.25 -23.005 ;
      RECT 55.15 -22.215 55.25 -21.68 ;
      RECT 55.15 -20.31 55.25 -19.775 ;
      RECT 55.15 -18.985 55.25 -18.45 ;
      RECT 55.15 -17.08 55.25 -16.545 ;
      RECT 55.15 -15.755 55.25 -15.22 ;
      RECT 55.15 -13.85 55.25 -13.315 ;
      RECT 55.15 -12.525 55.25 -11.99 ;
      RECT 55.15 -10.62 55.25 -10.085 ;
      RECT 55.15 -9.295 55.25 -8.76 ;
      RECT 55.15 -7.39 55.25 -6.855 ;
      RECT 55.15 -6.065 55.25 -5.53 ;
      RECT 55.15 -4.16 55.25 -3.625 ;
      RECT 55.15 -2.835 55.25 -2.3 ;
      RECT 55.15 -0.93 55.25 -0.395 ;
      RECT 55.15 0.395 55.25 0.93 ;
      RECT 55.025 -108.175 55.125 -107.215 ;
      RECT 54.65 -100.19 55 -100.07 ;
      RECT 54.65 -96.96 55 -96.84 ;
      RECT 54.65 -93.73 55 -93.61 ;
      RECT 54.65 -90.5 55 -90.38 ;
      RECT 54.65 -87.27 55 -87.15 ;
      RECT 54.65 -84.04 55 -83.92 ;
      RECT 54.65 -80.81 55 -80.69 ;
      RECT 54.65 -77.58 55 -77.46 ;
      RECT 54.65 -74.35 55 -74.23 ;
      RECT 54.65 -71.12 55 -71 ;
      RECT 54.65 -67.89 55 -67.77 ;
      RECT 54.65 -64.66 55 -64.54 ;
      RECT 54.65 -61.43 55 -61.31 ;
      RECT 54.65 -58.2 55 -58.08 ;
      RECT 54.65 -54.97 55 -54.85 ;
      RECT 54.65 -51.74 55 -51.62 ;
      RECT 54.65 -48.51 55 -48.39 ;
      RECT 54.65 -45.28 55 -45.16 ;
      RECT 54.65 -42.05 55 -41.93 ;
      RECT 54.65 -38.82 55 -38.7 ;
      RECT 54.65 -35.59 55 -35.47 ;
      RECT 54.65 -32.36 55 -32.24 ;
      RECT 54.65 -29.13 55 -29.01 ;
      RECT 54.65 -25.9 55 -25.78 ;
      RECT 54.65 -22.67 55 -22.55 ;
      RECT 54.65 -19.44 55 -19.32 ;
      RECT 54.65 -16.21 55 -16.09 ;
      RECT 54.65 -12.98 55 -12.86 ;
      RECT 54.65 -9.75 55 -9.63 ;
      RECT 54.65 -6.52 55 -6.4 ;
      RECT 54.65 -3.29 55 -3.17 ;
      RECT 54.65 -0.06 55 0.06 ;
      RECT 54.855 -112.255 54.955 -111.775 ;
      RECT 54.855 -110.765 54.955 -110.295 ;
      RECT 54.765 -108.175 54.865 -107.215 ;
      RECT 54.765 2.175 54.865 3.135 ;
      RECT 54.165 -100.19 54.515 -100.07 ;
      RECT 54.165 -96.96 54.515 -96.84 ;
      RECT 54.165 -93.73 54.515 -93.61 ;
      RECT 54.165 -90.5 54.515 -90.38 ;
      RECT 54.165 -87.27 54.515 -87.15 ;
      RECT 54.165 -84.04 54.515 -83.92 ;
      RECT 54.165 -80.81 54.515 -80.69 ;
      RECT 54.165 -77.58 54.515 -77.46 ;
      RECT 54.165 -74.35 54.515 -74.23 ;
      RECT 54.165 -71.12 54.515 -71 ;
      RECT 54.165 -67.89 54.515 -67.77 ;
      RECT 54.165 -64.66 54.515 -64.54 ;
      RECT 54.165 -61.43 54.515 -61.31 ;
      RECT 54.165 -58.2 54.515 -58.08 ;
      RECT 54.165 -54.97 54.515 -54.85 ;
      RECT 54.165 -51.74 54.515 -51.62 ;
      RECT 54.165 -48.51 54.515 -48.39 ;
      RECT 54.165 -45.28 54.515 -45.16 ;
      RECT 54.165 -42.05 54.515 -41.93 ;
      RECT 54.165 -38.82 54.515 -38.7 ;
      RECT 54.165 -35.59 54.515 -35.47 ;
      RECT 54.165 -32.36 54.515 -32.24 ;
      RECT 54.165 -29.13 54.515 -29.01 ;
      RECT 54.165 -25.9 54.515 -25.78 ;
      RECT 54.165 -22.67 54.515 -22.55 ;
      RECT 54.165 -19.44 54.515 -19.32 ;
      RECT 54.165 -16.21 54.515 -16.09 ;
      RECT 54.165 -12.98 54.515 -12.86 ;
      RECT 54.165 -9.75 54.515 -9.63 ;
      RECT 54.165 -6.52 54.515 -6.4 ;
      RECT 54.165 -3.29 54.515 -3.17 ;
      RECT 54.165 -0.06 54.515 0.06 ;
      RECT 54.335 -108.175 54.435 -107.215 ;
      RECT 54.335 2.175 54.435 3.135 ;
      RECT 54.23 -110.765 54.4 -110.385 ;
      RECT 54.265 -112.245 54.365 -111.775 ;
      RECT 54.075 -108.175 54.175 -107.215 ;
      RECT 53.95 -101.06 54.05 -100.525 ;
      RECT 53.95 -99.735 54.05 -99.2 ;
      RECT 53.95 -97.83 54.05 -97.295 ;
      RECT 53.95 -96.505 54.05 -95.97 ;
      RECT 53.95 -94.6 54.05 -94.065 ;
      RECT 53.95 -93.275 54.05 -92.74 ;
      RECT 53.95 -91.37 54.05 -90.835 ;
      RECT 53.95 -90.045 54.05 -89.51 ;
      RECT 53.95 -88.14 54.05 -87.605 ;
      RECT 53.95 -86.815 54.05 -86.28 ;
      RECT 53.95 -84.91 54.05 -84.375 ;
      RECT 53.95 -83.585 54.05 -83.05 ;
      RECT 53.95 -81.68 54.05 -81.145 ;
      RECT 53.95 -80.355 54.05 -79.82 ;
      RECT 53.95 -78.45 54.05 -77.915 ;
      RECT 53.95 -77.125 54.05 -76.59 ;
      RECT 53.95 -75.22 54.05 -74.685 ;
      RECT 53.95 -73.895 54.05 -73.36 ;
      RECT 53.95 -71.99 54.05 -71.455 ;
      RECT 53.95 -70.665 54.05 -70.13 ;
      RECT 53.95 -68.76 54.05 -68.225 ;
      RECT 53.95 -67.435 54.05 -66.9 ;
      RECT 53.95 -65.53 54.05 -64.995 ;
      RECT 53.95 -64.205 54.05 -63.67 ;
      RECT 53.95 -62.3 54.05 -61.765 ;
      RECT 53.95 -60.975 54.05 -60.44 ;
      RECT 53.95 -59.07 54.05 -58.535 ;
      RECT 53.95 -57.745 54.05 -57.21 ;
      RECT 53.95 -55.84 54.05 -55.305 ;
      RECT 53.95 -54.515 54.05 -53.98 ;
      RECT 53.95 -52.61 54.05 -52.075 ;
      RECT 53.95 -51.285 54.05 -50.75 ;
      RECT 53.95 -49.38 54.05 -48.845 ;
      RECT 53.95 -48.055 54.05 -47.52 ;
      RECT 53.95 -46.15 54.05 -45.615 ;
      RECT 53.95 -44.825 54.05 -44.29 ;
      RECT 53.95 -42.92 54.05 -42.385 ;
      RECT 53.95 -41.595 54.05 -41.06 ;
      RECT 53.95 -39.69 54.05 -39.155 ;
      RECT 53.95 -38.365 54.05 -37.83 ;
      RECT 53.95 -36.46 54.05 -35.925 ;
      RECT 53.95 -35.135 54.05 -34.6 ;
      RECT 53.95 -33.23 54.05 -32.695 ;
      RECT 53.95 -31.905 54.05 -31.37 ;
      RECT 53.95 -30 54.05 -29.465 ;
      RECT 53.95 -28.675 54.05 -28.14 ;
      RECT 53.95 -26.77 54.05 -26.235 ;
      RECT 53.95 -25.445 54.05 -24.91 ;
      RECT 53.95 -23.54 54.05 -23.005 ;
      RECT 53.95 -22.215 54.05 -21.68 ;
      RECT 53.95 -20.31 54.05 -19.775 ;
      RECT 53.95 -18.985 54.05 -18.45 ;
      RECT 53.95 -17.08 54.05 -16.545 ;
      RECT 53.95 -15.755 54.05 -15.22 ;
      RECT 53.95 -13.85 54.05 -13.315 ;
      RECT 53.95 -12.525 54.05 -11.99 ;
      RECT 53.95 -10.62 54.05 -10.085 ;
      RECT 53.95 -9.295 54.05 -8.76 ;
      RECT 53.95 -7.39 54.05 -6.855 ;
      RECT 53.95 -6.065 54.05 -5.53 ;
      RECT 53.95 -4.16 54.05 -3.625 ;
      RECT 53.95 -2.835 54.05 -2.3 ;
      RECT 53.95 -0.93 54.05 -0.395 ;
      RECT 53.95 0.395 54.05 0.93 ;
      RECT 53.825 -108.175 53.925 -107.215 ;
      RECT 53.45 -100.19 53.8 -100.07 ;
      RECT 53.45 -96.96 53.8 -96.84 ;
      RECT 53.45 -93.73 53.8 -93.61 ;
      RECT 53.45 -90.5 53.8 -90.38 ;
      RECT 53.45 -87.27 53.8 -87.15 ;
      RECT 53.45 -84.04 53.8 -83.92 ;
      RECT 53.45 -80.81 53.8 -80.69 ;
      RECT 53.45 -77.58 53.8 -77.46 ;
      RECT 53.45 -74.35 53.8 -74.23 ;
      RECT 53.45 -71.12 53.8 -71 ;
      RECT 53.45 -67.89 53.8 -67.77 ;
      RECT 53.45 -64.66 53.8 -64.54 ;
      RECT 53.45 -61.43 53.8 -61.31 ;
      RECT 53.45 -58.2 53.8 -58.08 ;
      RECT 53.45 -54.97 53.8 -54.85 ;
      RECT 53.45 -51.74 53.8 -51.62 ;
      RECT 53.45 -48.51 53.8 -48.39 ;
      RECT 53.45 -45.28 53.8 -45.16 ;
      RECT 53.45 -42.05 53.8 -41.93 ;
      RECT 53.45 -38.82 53.8 -38.7 ;
      RECT 53.45 -35.59 53.8 -35.47 ;
      RECT 53.45 -32.36 53.8 -32.24 ;
      RECT 53.45 -29.13 53.8 -29.01 ;
      RECT 53.45 -25.9 53.8 -25.78 ;
      RECT 53.45 -22.67 53.8 -22.55 ;
      RECT 53.45 -19.44 53.8 -19.32 ;
      RECT 53.45 -16.21 53.8 -16.09 ;
      RECT 53.45 -12.98 53.8 -12.86 ;
      RECT 53.45 -9.75 53.8 -9.63 ;
      RECT 53.45 -6.52 53.8 -6.4 ;
      RECT 53.45 -3.29 53.8 -3.17 ;
      RECT 53.45 -0.06 53.8 0.06 ;
      RECT 53.565 -108.175 53.665 -107.215 ;
      RECT 53.565 2.175 53.665 3.135 ;
      RECT 53.465 -113.555 53.565 -113.085 ;
      RECT 52.965 -100.19 53.315 -100.07 ;
      RECT 52.965 -96.96 53.315 -96.84 ;
      RECT 52.965 -93.73 53.315 -93.61 ;
      RECT 52.965 -90.5 53.315 -90.38 ;
      RECT 52.965 -87.27 53.315 -87.15 ;
      RECT 52.965 -84.04 53.315 -83.92 ;
      RECT 52.965 -80.81 53.315 -80.69 ;
      RECT 52.965 -77.58 53.315 -77.46 ;
      RECT 52.965 -74.35 53.315 -74.23 ;
      RECT 52.965 -71.12 53.315 -71 ;
      RECT 52.965 -67.89 53.315 -67.77 ;
      RECT 52.965 -64.66 53.315 -64.54 ;
      RECT 52.965 -61.43 53.315 -61.31 ;
      RECT 52.965 -58.2 53.315 -58.08 ;
      RECT 52.965 -54.97 53.315 -54.85 ;
      RECT 52.965 -51.74 53.315 -51.62 ;
      RECT 52.965 -48.51 53.315 -48.39 ;
      RECT 52.965 -45.28 53.315 -45.16 ;
      RECT 52.965 -42.05 53.315 -41.93 ;
      RECT 52.965 -38.82 53.315 -38.7 ;
      RECT 52.965 -35.59 53.315 -35.47 ;
      RECT 52.965 -32.36 53.315 -32.24 ;
      RECT 52.965 -29.13 53.315 -29.01 ;
      RECT 52.965 -25.9 53.315 -25.78 ;
      RECT 52.965 -22.67 53.315 -22.55 ;
      RECT 52.965 -19.44 53.315 -19.32 ;
      RECT 52.965 -16.21 53.315 -16.09 ;
      RECT 52.965 -12.98 53.315 -12.86 ;
      RECT 52.965 -9.75 53.315 -9.63 ;
      RECT 52.965 -6.52 53.315 -6.4 ;
      RECT 52.965 -3.29 53.315 -3.17 ;
      RECT 52.965 -0.06 53.315 0.06 ;
      RECT 53.1 -110.735 53.25 -110.445 ;
      RECT 53.135 -108.175 53.235 -107.215 ;
      RECT 53.135 2.175 53.235 3.135 ;
      RECT 53.115 -112.19 53.215 -111.65 ;
      RECT 52.875 -113.555 52.975 -113.085 ;
      RECT 52.875 -108.175 52.975 -107.215 ;
      RECT 52.75 -101.06 52.85 -100.525 ;
      RECT 52.75 -99.735 52.85 -99.2 ;
      RECT 52.75 -97.83 52.85 -97.295 ;
      RECT 52.75 -96.505 52.85 -95.97 ;
      RECT 52.75 -94.6 52.85 -94.065 ;
      RECT 52.75 -93.275 52.85 -92.74 ;
      RECT 52.75 -91.37 52.85 -90.835 ;
      RECT 52.75 -90.045 52.85 -89.51 ;
      RECT 52.75 -88.14 52.85 -87.605 ;
      RECT 52.75 -86.815 52.85 -86.28 ;
      RECT 52.75 -84.91 52.85 -84.375 ;
      RECT 52.75 -83.585 52.85 -83.05 ;
      RECT 52.75 -81.68 52.85 -81.145 ;
      RECT 52.75 -80.355 52.85 -79.82 ;
      RECT 52.75 -78.45 52.85 -77.915 ;
      RECT 52.75 -77.125 52.85 -76.59 ;
      RECT 52.75 -75.22 52.85 -74.685 ;
      RECT 52.75 -73.895 52.85 -73.36 ;
      RECT 52.75 -71.99 52.85 -71.455 ;
      RECT 52.75 -70.665 52.85 -70.13 ;
      RECT 52.75 -68.76 52.85 -68.225 ;
      RECT 52.75 -67.435 52.85 -66.9 ;
      RECT 52.75 -65.53 52.85 -64.995 ;
      RECT 52.75 -64.205 52.85 -63.67 ;
      RECT 52.75 -62.3 52.85 -61.765 ;
      RECT 52.75 -60.975 52.85 -60.44 ;
      RECT 52.75 -59.07 52.85 -58.535 ;
      RECT 52.75 -57.745 52.85 -57.21 ;
      RECT 52.75 -55.84 52.85 -55.305 ;
      RECT 52.75 -54.515 52.85 -53.98 ;
      RECT 52.75 -52.61 52.85 -52.075 ;
      RECT 52.75 -51.285 52.85 -50.75 ;
      RECT 52.75 -49.38 52.85 -48.845 ;
      RECT 52.75 -48.055 52.85 -47.52 ;
      RECT 52.75 -46.15 52.85 -45.615 ;
      RECT 52.75 -44.825 52.85 -44.29 ;
      RECT 52.75 -42.92 52.85 -42.385 ;
      RECT 52.75 -41.595 52.85 -41.06 ;
      RECT 52.75 -39.69 52.85 -39.155 ;
      RECT 52.75 -38.365 52.85 -37.83 ;
      RECT 52.75 -36.46 52.85 -35.925 ;
      RECT 52.75 -35.135 52.85 -34.6 ;
      RECT 52.75 -33.23 52.85 -32.695 ;
      RECT 52.75 -31.905 52.85 -31.37 ;
      RECT 52.75 -30 52.85 -29.465 ;
      RECT 52.75 -28.675 52.85 -28.14 ;
      RECT 52.75 -26.77 52.85 -26.235 ;
      RECT 52.75 -25.445 52.85 -24.91 ;
      RECT 52.75 -23.54 52.85 -23.005 ;
      RECT 52.75 -22.215 52.85 -21.68 ;
      RECT 52.75 -20.31 52.85 -19.775 ;
      RECT 52.75 -18.985 52.85 -18.45 ;
      RECT 52.75 -17.08 52.85 -16.545 ;
      RECT 52.75 -15.755 52.85 -15.22 ;
      RECT 52.75 -13.85 52.85 -13.315 ;
      RECT 52.75 -12.525 52.85 -11.99 ;
      RECT 52.75 -10.62 52.85 -10.085 ;
      RECT 52.75 -9.295 52.85 -8.76 ;
      RECT 52.75 -7.39 52.85 -6.855 ;
      RECT 52.75 -6.065 52.85 -5.53 ;
      RECT 52.75 -4.16 52.85 -3.625 ;
      RECT 52.75 -2.835 52.85 -2.3 ;
      RECT 52.75 -0.93 52.85 -0.395 ;
      RECT 52.75 0.395 52.85 0.93 ;
      RECT 52.625 -104.945 52.725 -103.985 ;
      RECT 52.25 -100.19 52.6 -100.07 ;
      RECT 52.25 -96.96 52.6 -96.84 ;
      RECT 52.25 -93.73 52.6 -93.61 ;
      RECT 52.25 -90.5 52.6 -90.38 ;
      RECT 52.25 -87.27 52.6 -87.15 ;
      RECT 52.25 -84.04 52.6 -83.92 ;
      RECT 52.25 -80.81 52.6 -80.69 ;
      RECT 52.25 -77.58 52.6 -77.46 ;
      RECT 52.25 -74.35 52.6 -74.23 ;
      RECT 52.25 -71.12 52.6 -71 ;
      RECT 52.25 -67.89 52.6 -67.77 ;
      RECT 52.25 -64.66 52.6 -64.54 ;
      RECT 52.25 -61.43 52.6 -61.31 ;
      RECT 52.25 -58.2 52.6 -58.08 ;
      RECT 52.25 -54.97 52.6 -54.85 ;
      RECT 52.25 -51.74 52.6 -51.62 ;
      RECT 52.25 -48.51 52.6 -48.39 ;
      RECT 52.25 -45.28 52.6 -45.16 ;
      RECT 52.25 -42.05 52.6 -41.93 ;
      RECT 52.25 -38.82 52.6 -38.7 ;
      RECT 52.25 -35.59 52.6 -35.47 ;
      RECT 52.25 -32.36 52.6 -32.24 ;
      RECT 52.25 -29.13 52.6 -29.01 ;
      RECT 52.25 -25.9 52.6 -25.78 ;
      RECT 52.25 -22.67 52.6 -22.55 ;
      RECT 52.25 -19.44 52.6 -19.32 ;
      RECT 52.25 -16.21 52.6 -16.09 ;
      RECT 52.25 -12.98 52.6 -12.86 ;
      RECT 52.25 -9.75 52.6 -9.63 ;
      RECT 52.25 -6.52 52.6 -6.4 ;
      RECT 52.25 -3.29 52.6 -3.17 ;
      RECT 52.25 -0.06 52.6 0.06 ;
      RECT 52.365 -104.945 52.465 -103.985 ;
      RECT 52.365 2.175 52.465 3.135 ;
      RECT 52.075 -112.255 52.175 -111.775 ;
      RECT 52.075 -110.765 52.175 -110.295 ;
      RECT 51.765 -100.19 52.115 -100.07 ;
      RECT 51.765 -96.96 52.115 -96.84 ;
      RECT 51.765 -93.73 52.115 -93.61 ;
      RECT 51.765 -90.5 52.115 -90.38 ;
      RECT 51.765 -87.27 52.115 -87.15 ;
      RECT 51.765 -84.04 52.115 -83.92 ;
      RECT 51.765 -80.81 52.115 -80.69 ;
      RECT 51.765 -77.58 52.115 -77.46 ;
      RECT 51.765 -74.35 52.115 -74.23 ;
      RECT 51.765 -71.12 52.115 -71 ;
      RECT 51.765 -67.89 52.115 -67.77 ;
      RECT 51.765 -64.66 52.115 -64.54 ;
      RECT 51.765 -61.43 52.115 -61.31 ;
      RECT 51.765 -58.2 52.115 -58.08 ;
      RECT 51.765 -54.97 52.115 -54.85 ;
      RECT 51.765 -51.74 52.115 -51.62 ;
      RECT 51.765 -48.51 52.115 -48.39 ;
      RECT 51.765 -45.28 52.115 -45.16 ;
      RECT 51.765 -42.05 52.115 -41.93 ;
      RECT 51.765 -38.82 52.115 -38.7 ;
      RECT 51.765 -35.59 52.115 -35.47 ;
      RECT 51.765 -32.36 52.115 -32.24 ;
      RECT 51.765 -29.13 52.115 -29.01 ;
      RECT 51.765 -25.9 52.115 -25.78 ;
      RECT 51.765 -22.67 52.115 -22.55 ;
      RECT 51.765 -19.44 52.115 -19.32 ;
      RECT 51.765 -16.21 52.115 -16.09 ;
      RECT 51.765 -12.98 52.115 -12.86 ;
      RECT 51.765 -9.75 52.115 -9.63 ;
      RECT 51.765 -6.52 52.115 -6.4 ;
      RECT 51.765 -3.29 52.115 -3.17 ;
      RECT 51.765 -0.06 52.115 0.06 ;
      RECT 51.935 -104.945 52.035 -103.985 ;
      RECT 51.935 2.175 52.035 3.135 ;
      RECT 48.035 -108.655 51.815 -108.535 ;
      RECT 51.675 -104.945 51.775 -103.985 ;
      RECT 51.55 -101.06 51.65 -100.525 ;
      RECT 51.55 -99.735 51.65 -99.2 ;
      RECT 51.55 -97.83 51.65 -97.295 ;
      RECT 51.55 -96.505 51.65 -95.97 ;
      RECT 51.55 -94.6 51.65 -94.065 ;
      RECT 51.55 -93.275 51.65 -92.74 ;
      RECT 51.55 -91.37 51.65 -90.835 ;
      RECT 51.55 -90.045 51.65 -89.51 ;
      RECT 51.55 -88.14 51.65 -87.605 ;
      RECT 51.55 -86.815 51.65 -86.28 ;
      RECT 51.55 -84.91 51.65 -84.375 ;
      RECT 51.55 -83.585 51.65 -83.05 ;
      RECT 51.55 -81.68 51.65 -81.145 ;
      RECT 51.55 -80.355 51.65 -79.82 ;
      RECT 51.55 -78.45 51.65 -77.915 ;
      RECT 51.55 -77.125 51.65 -76.59 ;
      RECT 51.55 -75.22 51.65 -74.685 ;
      RECT 51.55 -73.895 51.65 -73.36 ;
      RECT 51.55 -71.99 51.65 -71.455 ;
      RECT 51.55 -70.665 51.65 -70.13 ;
      RECT 51.55 -68.76 51.65 -68.225 ;
      RECT 51.55 -67.435 51.65 -66.9 ;
      RECT 51.55 -65.53 51.65 -64.995 ;
      RECT 51.55 -64.205 51.65 -63.67 ;
      RECT 51.55 -62.3 51.65 -61.765 ;
      RECT 51.55 -60.975 51.65 -60.44 ;
      RECT 51.55 -59.07 51.65 -58.535 ;
      RECT 51.55 -57.745 51.65 -57.21 ;
      RECT 51.55 -55.84 51.65 -55.305 ;
      RECT 51.55 -54.515 51.65 -53.98 ;
      RECT 51.55 -52.61 51.65 -52.075 ;
      RECT 51.55 -51.285 51.65 -50.75 ;
      RECT 51.55 -49.38 51.65 -48.845 ;
      RECT 51.55 -48.055 51.65 -47.52 ;
      RECT 51.55 -46.15 51.65 -45.615 ;
      RECT 51.55 -44.825 51.65 -44.29 ;
      RECT 51.55 -42.92 51.65 -42.385 ;
      RECT 51.55 -41.595 51.65 -41.06 ;
      RECT 51.55 -39.69 51.65 -39.155 ;
      RECT 51.55 -38.365 51.65 -37.83 ;
      RECT 51.55 -36.46 51.65 -35.925 ;
      RECT 51.55 -35.135 51.65 -34.6 ;
      RECT 51.55 -33.23 51.65 -32.695 ;
      RECT 51.55 -31.905 51.65 -31.37 ;
      RECT 51.55 -30 51.65 -29.465 ;
      RECT 51.55 -28.675 51.65 -28.14 ;
      RECT 51.55 -26.77 51.65 -26.235 ;
      RECT 51.55 -25.445 51.65 -24.91 ;
      RECT 51.55 -23.54 51.65 -23.005 ;
      RECT 51.55 -22.215 51.65 -21.68 ;
      RECT 51.55 -20.31 51.65 -19.775 ;
      RECT 51.55 -18.985 51.65 -18.45 ;
      RECT 51.55 -17.08 51.65 -16.545 ;
      RECT 51.55 -15.755 51.65 -15.22 ;
      RECT 51.55 -13.85 51.65 -13.315 ;
      RECT 51.55 -12.525 51.65 -11.99 ;
      RECT 51.55 -10.62 51.65 -10.085 ;
      RECT 51.55 -9.295 51.65 -8.76 ;
      RECT 51.55 -7.39 51.65 -6.855 ;
      RECT 51.55 -6.065 51.65 -5.53 ;
      RECT 51.55 -4.16 51.65 -3.625 ;
      RECT 51.55 -2.835 51.65 -2.3 ;
      RECT 51.55 -0.93 51.65 -0.395 ;
      RECT 51.55 0.395 51.65 0.93 ;
      RECT 51.485 -110.75 51.605 -110.37 ;
      RECT 51.485 -112.245 51.585 -111.775 ;
      RECT 51.425 -104.945 51.525 -103.985 ;
      RECT 51.05 -100.19 51.4 -100.07 ;
      RECT 51.05 -96.96 51.4 -96.84 ;
      RECT 51.05 -93.73 51.4 -93.61 ;
      RECT 51.05 -90.5 51.4 -90.38 ;
      RECT 51.05 -87.27 51.4 -87.15 ;
      RECT 51.05 -84.04 51.4 -83.92 ;
      RECT 51.05 -80.81 51.4 -80.69 ;
      RECT 51.05 -77.58 51.4 -77.46 ;
      RECT 51.05 -74.35 51.4 -74.23 ;
      RECT 51.05 -71.12 51.4 -71 ;
      RECT 51.05 -67.89 51.4 -67.77 ;
      RECT 51.05 -64.66 51.4 -64.54 ;
      RECT 51.05 -61.43 51.4 -61.31 ;
      RECT 51.05 -58.2 51.4 -58.08 ;
      RECT 51.05 -54.97 51.4 -54.85 ;
      RECT 51.05 -51.74 51.4 -51.62 ;
      RECT 51.05 -48.51 51.4 -48.39 ;
      RECT 51.05 -45.28 51.4 -45.16 ;
      RECT 51.05 -42.05 51.4 -41.93 ;
      RECT 51.05 -38.82 51.4 -38.7 ;
      RECT 51.05 -35.59 51.4 -35.47 ;
      RECT 51.05 -32.36 51.4 -32.24 ;
      RECT 51.05 -29.13 51.4 -29.01 ;
      RECT 51.05 -25.9 51.4 -25.78 ;
      RECT 51.05 -22.67 51.4 -22.55 ;
      RECT 51.05 -19.44 51.4 -19.32 ;
      RECT 51.05 -16.21 51.4 -16.09 ;
      RECT 51.05 -12.98 51.4 -12.86 ;
      RECT 51.05 -9.75 51.4 -9.63 ;
      RECT 51.05 -6.52 51.4 -6.4 ;
      RECT 51.05 -3.29 51.4 -3.17 ;
      RECT 51.05 -0.06 51.4 0.06 ;
      RECT 51.165 -104.945 51.265 -103.985 ;
      RECT 51.165 2.175 51.265 3.135 ;
      RECT 50.895 -109.595 51.03 -109.275 ;
      RECT 50.565 -100.19 50.915 -100.07 ;
      RECT 50.565 -96.96 50.915 -96.84 ;
      RECT 50.565 -93.73 50.915 -93.61 ;
      RECT 50.565 -90.5 50.915 -90.38 ;
      RECT 50.565 -87.27 50.915 -87.15 ;
      RECT 50.565 -84.04 50.915 -83.92 ;
      RECT 50.565 -80.81 50.915 -80.69 ;
      RECT 50.565 -77.58 50.915 -77.46 ;
      RECT 50.565 -74.35 50.915 -74.23 ;
      RECT 50.565 -71.12 50.915 -71 ;
      RECT 50.565 -67.89 50.915 -67.77 ;
      RECT 50.565 -64.66 50.915 -64.54 ;
      RECT 50.565 -61.43 50.915 -61.31 ;
      RECT 50.565 -58.2 50.915 -58.08 ;
      RECT 50.565 -54.97 50.915 -54.85 ;
      RECT 50.565 -51.74 50.915 -51.62 ;
      RECT 50.565 -48.51 50.915 -48.39 ;
      RECT 50.565 -45.28 50.915 -45.16 ;
      RECT 50.565 -42.05 50.915 -41.93 ;
      RECT 50.565 -38.82 50.915 -38.7 ;
      RECT 50.565 -35.59 50.915 -35.47 ;
      RECT 50.565 -32.36 50.915 -32.24 ;
      RECT 50.565 -29.13 50.915 -29.01 ;
      RECT 50.565 -25.9 50.915 -25.78 ;
      RECT 50.565 -22.67 50.915 -22.55 ;
      RECT 50.565 -19.44 50.915 -19.32 ;
      RECT 50.565 -16.21 50.915 -16.09 ;
      RECT 50.565 -12.98 50.915 -12.86 ;
      RECT 50.565 -9.75 50.915 -9.63 ;
      RECT 50.565 -6.52 50.915 -6.4 ;
      RECT 50.565 -3.29 50.915 -3.17 ;
      RECT 50.565 -0.06 50.915 0.06 ;
      RECT 50.735 -104.945 50.835 -103.985 ;
      RECT 50.735 2.175 50.835 3.135 ;
      RECT 50.56 -109.595 50.705 -109.275 ;
      RECT 50.475 -104.945 50.575 -103.985 ;
      RECT 50.35 -101.06 50.45 -100.525 ;
      RECT 50.35 -99.735 50.45 -99.2 ;
      RECT 50.35 -97.83 50.45 -97.295 ;
      RECT 50.35 -96.505 50.45 -95.97 ;
      RECT 50.35 -94.6 50.45 -94.065 ;
      RECT 50.35 -93.275 50.45 -92.74 ;
      RECT 50.35 -91.37 50.45 -90.835 ;
      RECT 50.35 -90.045 50.45 -89.51 ;
      RECT 50.35 -88.14 50.45 -87.605 ;
      RECT 50.35 -86.815 50.45 -86.28 ;
      RECT 50.35 -84.91 50.45 -84.375 ;
      RECT 50.35 -83.585 50.45 -83.05 ;
      RECT 50.35 -81.68 50.45 -81.145 ;
      RECT 50.35 -80.355 50.45 -79.82 ;
      RECT 50.35 -78.45 50.45 -77.915 ;
      RECT 50.35 -77.125 50.45 -76.59 ;
      RECT 50.35 -75.22 50.45 -74.685 ;
      RECT 50.35 -73.895 50.45 -73.36 ;
      RECT 50.35 -71.99 50.45 -71.455 ;
      RECT 50.35 -70.665 50.45 -70.13 ;
      RECT 50.35 -68.76 50.45 -68.225 ;
      RECT 50.35 -67.435 50.45 -66.9 ;
      RECT 50.35 -65.53 50.45 -64.995 ;
      RECT 50.35 -64.205 50.45 -63.67 ;
      RECT 50.35 -62.3 50.45 -61.765 ;
      RECT 50.35 -60.975 50.45 -60.44 ;
      RECT 50.35 -59.07 50.45 -58.535 ;
      RECT 50.35 -57.745 50.45 -57.21 ;
      RECT 50.35 -55.84 50.45 -55.305 ;
      RECT 50.35 -54.515 50.45 -53.98 ;
      RECT 50.35 -52.61 50.45 -52.075 ;
      RECT 50.35 -51.285 50.45 -50.75 ;
      RECT 50.35 -49.38 50.45 -48.845 ;
      RECT 50.35 -48.055 50.45 -47.52 ;
      RECT 50.35 -46.15 50.45 -45.615 ;
      RECT 50.35 -44.825 50.45 -44.29 ;
      RECT 50.35 -42.92 50.45 -42.385 ;
      RECT 50.35 -41.595 50.45 -41.06 ;
      RECT 50.35 -39.69 50.45 -39.155 ;
      RECT 50.35 -38.365 50.45 -37.83 ;
      RECT 50.35 -36.46 50.45 -35.925 ;
      RECT 50.35 -35.135 50.45 -34.6 ;
      RECT 50.35 -33.23 50.45 -32.695 ;
      RECT 50.35 -31.905 50.45 -31.37 ;
      RECT 50.35 -30 50.45 -29.465 ;
      RECT 50.35 -28.675 50.45 -28.14 ;
      RECT 50.35 -26.77 50.45 -26.235 ;
      RECT 50.35 -25.445 50.45 -24.91 ;
      RECT 50.35 -23.54 50.45 -23.005 ;
      RECT 50.35 -22.215 50.45 -21.68 ;
      RECT 50.35 -20.31 50.45 -19.775 ;
      RECT 50.35 -18.985 50.45 -18.45 ;
      RECT 50.35 -17.08 50.45 -16.545 ;
      RECT 50.35 -15.755 50.45 -15.22 ;
      RECT 50.35 -13.85 50.45 -13.315 ;
      RECT 50.35 -12.525 50.45 -11.99 ;
      RECT 50.35 -10.62 50.45 -10.085 ;
      RECT 50.35 -9.295 50.45 -8.76 ;
      RECT 50.35 -7.39 50.45 -6.855 ;
      RECT 50.35 -6.065 50.45 -5.53 ;
      RECT 50.35 -4.16 50.45 -3.625 ;
      RECT 50.35 -2.835 50.45 -2.3 ;
      RECT 50.35 -0.93 50.45 -0.395 ;
      RECT 50.35 0.395 50.45 0.93 ;
      RECT 50.225 -108.175 50.325 -107.215 ;
      RECT 49.85 -100.19 50.2 -100.07 ;
      RECT 49.85 -96.96 50.2 -96.84 ;
      RECT 49.85 -93.73 50.2 -93.61 ;
      RECT 49.85 -90.5 50.2 -90.38 ;
      RECT 49.85 -87.27 50.2 -87.15 ;
      RECT 49.85 -84.04 50.2 -83.92 ;
      RECT 49.85 -80.81 50.2 -80.69 ;
      RECT 49.85 -77.58 50.2 -77.46 ;
      RECT 49.85 -74.35 50.2 -74.23 ;
      RECT 49.85 -71.12 50.2 -71 ;
      RECT 49.85 -67.89 50.2 -67.77 ;
      RECT 49.85 -64.66 50.2 -64.54 ;
      RECT 49.85 -61.43 50.2 -61.31 ;
      RECT 49.85 -58.2 50.2 -58.08 ;
      RECT 49.85 -54.97 50.2 -54.85 ;
      RECT 49.85 -51.74 50.2 -51.62 ;
      RECT 49.85 -48.51 50.2 -48.39 ;
      RECT 49.85 -45.28 50.2 -45.16 ;
      RECT 49.85 -42.05 50.2 -41.93 ;
      RECT 49.85 -38.82 50.2 -38.7 ;
      RECT 49.85 -35.59 50.2 -35.47 ;
      RECT 49.85 -32.36 50.2 -32.24 ;
      RECT 49.85 -29.13 50.2 -29.01 ;
      RECT 49.85 -25.9 50.2 -25.78 ;
      RECT 49.85 -22.67 50.2 -22.55 ;
      RECT 49.85 -19.44 50.2 -19.32 ;
      RECT 49.85 -16.21 50.2 -16.09 ;
      RECT 49.85 -12.98 50.2 -12.86 ;
      RECT 49.85 -9.75 50.2 -9.63 ;
      RECT 49.85 -6.52 50.2 -6.4 ;
      RECT 49.85 -3.29 50.2 -3.17 ;
      RECT 49.85 -0.06 50.2 0.06 ;
      RECT 50.055 -112.255 50.155 -111.775 ;
      RECT 50.055 -110.765 50.155 -110.295 ;
      RECT 49.965 -108.175 50.065 -107.215 ;
      RECT 49.965 2.175 50.065 3.135 ;
      RECT 49.365 -100.19 49.715 -100.07 ;
      RECT 49.365 -96.96 49.715 -96.84 ;
      RECT 49.365 -93.73 49.715 -93.61 ;
      RECT 49.365 -90.5 49.715 -90.38 ;
      RECT 49.365 -87.27 49.715 -87.15 ;
      RECT 49.365 -84.04 49.715 -83.92 ;
      RECT 49.365 -80.81 49.715 -80.69 ;
      RECT 49.365 -77.58 49.715 -77.46 ;
      RECT 49.365 -74.35 49.715 -74.23 ;
      RECT 49.365 -71.12 49.715 -71 ;
      RECT 49.365 -67.89 49.715 -67.77 ;
      RECT 49.365 -64.66 49.715 -64.54 ;
      RECT 49.365 -61.43 49.715 -61.31 ;
      RECT 49.365 -58.2 49.715 -58.08 ;
      RECT 49.365 -54.97 49.715 -54.85 ;
      RECT 49.365 -51.74 49.715 -51.62 ;
      RECT 49.365 -48.51 49.715 -48.39 ;
      RECT 49.365 -45.28 49.715 -45.16 ;
      RECT 49.365 -42.05 49.715 -41.93 ;
      RECT 49.365 -38.82 49.715 -38.7 ;
      RECT 49.365 -35.59 49.715 -35.47 ;
      RECT 49.365 -32.36 49.715 -32.24 ;
      RECT 49.365 -29.13 49.715 -29.01 ;
      RECT 49.365 -25.9 49.715 -25.78 ;
      RECT 49.365 -22.67 49.715 -22.55 ;
      RECT 49.365 -19.44 49.715 -19.32 ;
      RECT 49.365 -16.21 49.715 -16.09 ;
      RECT 49.365 -12.98 49.715 -12.86 ;
      RECT 49.365 -9.75 49.715 -9.63 ;
      RECT 49.365 -6.52 49.715 -6.4 ;
      RECT 49.365 -3.29 49.715 -3.17 ;
      RECT 49.365 -0.06 49.715 0.06 ;
      RECT 49.535 -108.175 49.635 -107.215 ;
      RECT 49.535 2.175 49.635 3.135 ;
      RECT 49.43 -110.765 49.6 -110.385 ;
      RECT 49.465 -112.245 49.565 -111.775 ;
      RECT 49.275 -108.175 49.375 -107.215 ;
      RECT 49.15 -101.06 49.25 -100.525 ;
      RECT 49.15 -99.735 49.25 -99.2 ;
      RECT 49.15 -97.83 49.25 -97.295 ;
      RECT 49.15 -96.505 49.25 -95.97 ;
      RECT 49.15 -94.6 49.25 -94.065 ;
      RECT 49.15 -93.275 49.25 -92.74 ;
      RECT 49.15 -91.37 49.25 -90.835 ;
      RECT 49.15 -90.045 49.25 -89.51 ;
      RECT 49.15 -88.14 49.25 -87.605 ;
      RECT 49.15 -86.815 49.25 -86.28 ;
      RECT 49.15 -84.91 49.25 -84.375 ;
      RECT 49.15 -83.585 49.25 -83.05 ;
      RECT 49.15 -81.68 49.25 -81.145 ;
      RECT 49.15 -80.355 49.25 -79.82 ;
      RECT 49.15 -78.45 49.25 -77.915 ;
      RECT 49.15 -77.125 49.25 -76.59 ;
      RECT 49.15 -75.22 49.25 -74.685 ;
      RECT 49.15 -73.895 49.25 -73.36 ;
      RECT 49.15 -71.99 49.25 -71.455 ;
      RECT 49.15 -70.665 49.25 -70.13 ;
      RECT 49.15 -68.76 49.25 -68.225 ;
      RECT 49.15 -67.435 49.25 -66.9 ;
      RECT 49.15 -65.53 49.25 -64.995 ;
      RECT 49.15 -64.205 49.25 -63.67 ;
      RECT 49.15 -62.3 49.25 -61.765 ;
      RECT 49.15 -60.975 49.25 -60.44 ;
      RECT 49.15 -59.07 49.25 -58.535 ;
      RECT 49.15 -57.745 49.25 -57.21 ;
      RECT 49.15 -55.84 49.25 -55.305 ;
      RECT 49.15 -54.515 49.25 -53.98 ;
      RECT 49.15 -52.61 49.25 -52.075 ;
      RECT 49.15 -51.285 49.25 -50.75 ;
      RECT 49.15 -49.38 49.25 -48.845 ;
      RECT 49.15 -48.055 49.25 -47.52 ;
      RECT 49.15 -46.15 49.25 -45.615 ;
      RECT 49.15 -44.825 49.25 -44.29 ;
      RECT 49.15 -42.92 49.25 -42.385 ;
      RECT 49.15 -41.595 49.25 -41.06 ;
      RECT 49.15 -39.69 49.25 -39.155 ;
      RECT 49.15 -38.365 49.25 -37.83 ;
      RECT 49.15 -36.46 49.25 -35.925 ;
      RECT 49.15 -35.135 49.25 -34.6 ;
      RECT 49.15 -33.23 49.25 -32.695 ;
      RECT 49.15 -31.905 49.25 -31.37 ;
      RECT 49.15 -30 49.25 -29.465 ;
      RECT 49.15 -28.675 49.25 -28.14 ;
      RECT 49.15 -26.77 49.25 -26.235 ;
      RECT 49.15 -25.445 49.25 -24.91 ;
      RECT 49.15 -23.54 49.25 -23.005 ;
      RECT 49.15 -22.215 49.25 -21.68 ;
      RECT 49.15 -20.31 49.25 -19.775 ;
      RECT 49.15 -18.985 49.25 -18.45 ;
      RECT 49.15 -17.08 49.25 -16.545 ;
      RECT 49.15 -15.755 49.25 -15.22 ;
      RECT 49.15 -13.85 49.25 -13.315 ;
      RECT 49.15 -12.525 49.25 -11.99 ;
      RECT 49.15 -10.62 49.25 -10.085 ;
      RECT 49.15 -9.295 49.25 -8.76 ;
      RECT 49.15 -7.39 49.25 -6.855 ;
      RECT 49.15 -6.065 49.25 -5.53 ;
      RECT 49.15 -4.16 49.25 -3.625 ;
      RECT 49.15 -2.835 49.25 -2.3 ;
      RECT 49.15 -0.93 49.25 -0.395 ;
      RECT 49.15 0.395 49.25 0.93 ;
      RECT 49.025 -108.175 49.125 -107.215 ;
      RECT 48.65 -100.19 49 -100.07 ;
      RECT 48.65 -96.96 49 -96.84 ;
      RECT 48.65 -93.73 49 -93.61 ;
      RECT 48.65 -90.5 49 -90.38 ;
      RECT 48.65 -87.27 49 -87.15 ;
      RECT 48.65 -84.04 49 -83.92 ;
      RECT 48.65 -80.81 49 -80.69 ;
      RECT 48.65 -77.58 49 -77.46 ;
      RECT 48.65 -74.35 49 -74.23 ;
      RECT 48.65 -71.12 49 -71 ;
      RECT 48.65 -67.89 49 -67.77 ;
      RECT 48.65 -64.66 49 -64.54 ;
      RECT 48.65 -61.43 49 -61.31 ;
      RECT 48.65 -58.2 49 -58.08 ;
      RECT 48.65 -54.97 49 -54.85 ;
      RECT 48.65 -51.74 49 -51.62 ;
      RECT 48.65 -48.51 49 -48.39 ;
      RECT 48.65 -45.28 49 -45.16 ;
      RECT 48.65 -42.05 49 -41.93 ;
      RECT 48.65 -38.82 49 -38.7 ;
      RECT 48.65 -35.59 49 -35.47 ;
      RECT 48.65 -32.36 49 -32.24 ;
      RECT 48.65 -29.13 49 -29.01 ;
      RECT 48.65 -25.9 49 -25.78 ;
      RECT 48.65 -22.67 49 -22.55 ;
      RECT 48.65 -19.44 49 -19.32 ;
      RECT 48.65 -16.21 49 -16.09 ;
      RECT 48.65 -12.98 49 -12.86 ;
      RECT 48.65 -9.75 49 -9.63 ;
      RECT 48.65 -6.52 49 -6.4 ;
      RECT 48.65 -3.29 49 -3.17 ;
      RECT 48.65 -0.06 49 0.06 ;
      RECT 48.765 -108.175 48.865 -107.215 ;
      RECT 48.765 2.175 48.865 3.135 ;
      RECT 48.665 -113.555 48.765 -113.085 ;
      RECT 48.165 -100.19 48.515 -100.07 ;
      RECT 48.165 -96.96 48.515 -96.84 ;
      RECT 48.165 -93.73 48.515 -93.61 ;
      RECT 48.165 -90.5 48.515 -90.38 ;
      RECT 48.165 -87.27 48.515 -87.15 ;
      RECT 48.165 -84.04 48.515 -83.92 ;
      RECT 48.165 -80.81 48.515 -80.69 ;
      RECT 48.165 -77.58 48.515 -77.46 ;
      RECT 48.165 -74.35 48.515 -74.23 ;
      RECT 48.165 -71.12 48.515 -71 ;
      RECT 48.165 -67.89 48.515 -67.77 ;
      RECT 48.165 -64.66 48.515 -64.54 ;
      RECT 48.165 -61.43 48.515 -61.31 ;
      RECT 48.165 -58.2 48.515 -58.08 ;
      RECT 48.165 -54.97 48.515 -54.85 ;
      RECT 48.165 -51.74 48.515 -51.62 ;
      RECT 48.165 -48.51 48.515 -48.39 ;
      RECT 48.165 -45.28 48.515 -45.16 ;
      RECT 48.165 -42.05 48.515 -41.93 ;
      RECT 48.165 -38.82 48.515 -38.7 ;
      RECT 48.165 -35.59 48.515 -35.47 ;
      RECT 48.165 -32.36 48.515 -32.24 ;
      RECT 48.165 -29.13 48.515 -29.01 ;
      RECT 48.165 -25.9 48.515 -25.78 ;
      RECT 48.165 -22.67 48.515 -22.55 ;
      RECT 48.165 -19.44 48.515 -19.32 ;
      RECT 48.165 -16.21 48.515 -16.09 ;
      RECT 48.165 -12.98 48.515 -12.86 ;
      RECT 48.165 -9.75 48.515 -9.63 ;
      RECT 48.165 -6.52 48.515 -6.4 ;
      RECT 48.165 -3.29 48.515 -3.17 ;
      RECT 48.165 -0.06 48.515 0.06 ;
      RECT 48.3 -110.735 48.45 -110.445 ;
      RECT 48.335 -108.175 48.435 -107.215 ;
      RECT 48.335 2.175 48.435 3.135 ;
      RECT 48.315 -112.19 48.415 -111.65 ;
      RECT 48.075 -113.555 48.175 -113.085 ;
      RECT 48.075 -108.175 48.175 -107.215 ;
      RECT 47.95 -101.06 48.05 -100.525 ;
      RECT 47.95 -99.735 48.05 -99.2 ;
      RECT 47.95 -97.83 48.05 -97.295 ;
      RECT 47.95 -96.505 48.05 -95.97 ;
      RECT 47.95 -94.6 48.05 -94.065 ;
      RECT 47.95 -93.275 48.05 -92.74 ;
      RECT 47.95 -91.37 48.05 -90.835 ;
      RECT 47.95 -90.045 48.05 -89.51 ;
      RECT 47.95 -88.14 48.05 -87.605 ;
      RECT 47.95 -86.815 48.05 -86.28 ;
      RECT 47.95 -84.91 48.05 -84.375 ;
      RECT 47.95 -83.585 48.05 -83.05 ;
      RECT 47.95 -81.68 48.05 -81.145 ;
      RECT 47.95 -80.355 48.05 -79.82 ;
      RECT 47.95 -78.45 48.05 -77.915 ;
      RECT 47.95 -77.125 48.05 -76.59 ;
      RECT 47.95 -75.22 48.05 -74.685 ;
      RECT 47.95 -73.895 48.05 -73.36 ;
      RECT 47.95 -71.99 48.05 -71.455 ;
      RECT 47.95 -70.665 48.05 -70.13 ;
      RECT 47.95 -68.76 48.05 -68.225 ;
      RECT 47.95 -67.435 48.05 -66.9 ;
      RECT 47.95 -65.53 48.05 -64.995 ;
      RECT 47.95 -64.205 48.05 -63.67 ;
      RECT 47.95 -62.3 48.05 -61.765 ;
      RECT 47.95 -60.975 48.05 -60.44 ;
      RECT 47.95 -59.07 48.05 -58.535 ;
      RECT 47.95 -57.745 48.05 -57.21 ;
      RECT 47.95 -55.84 48.05 -55.305 ;
      RECT 47.95 -54.515 48.05 -53.98 ;
      RECT 47.95 -52.61 48.05 -52.075 ;
      RECT 47.95 -51.285 48.05 -50.75 ;
      RECT 47.95 -49.38 48.05 -48.845 ;
      RECT 47.95 -48.055 48.05 -47.52 ;
      RECT 47.95 -46.15 48.05 -45.615 ;
      RECT 47.95 -44.825 48.05 -44.29 ;
      RECT 47.95 -42.92 48.05 -42.385 ;
      RECT 47.95 -41.595 48.05 -41.06 ;
      RECT 47.95 -39.69 48.05 -39.155 ;
      RECT 47.95 -38.365 48.05 -37.83 ;
      RECT 47.95 -36.46 48.05 -35.925 ;
      RECT 47.95 -35.135 48.05 -34.6 ;
      RECT 47.95 -33.23 48.05 -32.695 ;
      RECT 47.95 -31.905 48.05 -31.37 ;
      RECT 47.95 -30 48.05 -29.465 ;
      RECT 47.95 -28.675 48.05 -28.14 ;
      RECT 47.95 -26.77 48.05 -26.235 ;
      RECT 47.95 -25.445 48.05 -24.91 ;
      RECT 47.95 -23.54 48.05 -23.005 ;
      RECT 47.95 -22.215 48.05 -21.68 ;
      RECT 47.95 -20.31 48.05 -19.775 ;
      RECT 47.95 -18.985 48.05 -18.45 ;
      RECT 47.95 -17.08 48.05 -16.545 ;
      RECT 47.95 -15.755 48.05 -15.22 ;
      RECT 47.95 -13.85 48.05 -13.315 ;
      RECT 47.95 -12.525 48.05 -11.99 ;
      RECT 47.95 -10.62 48.05 -10.085 ;
      RECT 47.95 -9.295 48.05 -8.76 ;
      RECT 47.95 -7.39 48.05 -6.855 ;
      RECT 47.95 -6.065 48.05 -5.53 ;
      RECT 47.95 -4.16 48.05 -3.625 ;
      RECT 47.95 -2.835 48.05 -2.3 ;
      RECT 47.95 -0.93 48.05 -0.395 ;
      RECT 47.95 0.395 48.05 0.93 ;
      RECT 47.825 -104.945 47.925 -103.985 ;
      RECT 47.45 -100.19 47.8 -100.07 ;
      RECT 47.45 -96.96 47.8 -96.84 ;
      RECT 47.45 -93.73 47.8 -93.61 ;
      RECT 47.45 -90.5 47.8 -90.38 ;
      RECT 47.45 -87.27 47.8 -87.15 ;
      RECT 47.45 -84.04 47.8 -83.92 ;
      RECT 47.45 -80.81 47.8 -80.69 ;
      RECT 47.45 -77.58 47.8 -77.46 ;
      RECT 47.45 -74.35 47.8 -74.23 ;
      RECT 47.45 -71.12 47.8 -71 ;
      RECT 47.45 -67.89 47.8 -67.77 ;
      RECT 47.45 -64.66 47.8 -64.54 ;
      RECT 47.45 -61.43 47.8 -61.31 ;
      RECT 47.45 -58.2 47.8 -58.08 ;
      RECT 47.45 -54.97 47.8 -54.85 ;
      RECT 47.45 -51.74 47.8 -51.62 ;
      RECT 47.45 -48.51 47.8 -48.39 ;
      RECT 47.45 -45.28 47.8 -45.16 ;
      RECT 47.45 -42.05 47.8 -41.93 ;
      RECT 47.45 -38.82 47.8 -38.7 ;
      RECT 47.45 -35.59 47.8 -35.47 ;
      RECT 47.45 -32.36 47.8 -32.24 ;
      RECT 47.45 -29.13 47.8 -29.01 ;
      RECT 47.45 -25.9 47.8 -25.78 ;
      RECT 47.45 -22.67 47.8 -22.55 ;
      RECT 47.45 -19.44 47.8 -19.32 ;
      RECT 47.45 -16.21 47.8 -16.09 ;
      RECT 47.45 -12.98 47.8 -12.86 ;
      RECT 47.45 -9.75 47.8 -9.63 ;
      RECT 47.45 -6.52 47.8 -6.4 ;
      RECT 47.45 -3.29 47.8 -3.17 ;
      RECT 47.45 -0.06 47.8 0.06 ;
      RECT 47.565 -104.945 47.665 -103.985 ;
      RECT 47.565 2.175 47.665 3.135 ;
      RECT 47.275 -112.255 47.375 -111.775 ;
      RECT 47.275 -110.765 47.375 -110.295 ;
      RECT 46.965 -100.19 47.315 -100.07 ;
      RECT 46.965 -96.96 47.315 -96.84 ;
      RECT 46.965 -93.73 47.315 -93.61 ;
      RECT 46.965 -90.5 47.315 -90.38 ;
      RECT 46.965 -87.27 47.315 -87.15 ;
      RECT 46.965 -84.04 47.315 -83.92 ;
      RECT 46.965 -80.81 47.315 -80.69 ;
      RECT 46.965 -77.58 47.315 -77.46 ;
      RECT 46.965 -74.35 47.315 -74.23 ;
      RECT 46.965 -71.12 47.315 -71 ;
      RECT 46.965 -67.89 47.315 -67.77 ;
      RECT 46.965 -64.66 47.315 -64.54 ;
      RECT 46.965 -61.43 47.315 -61.31 ;
      RECT 46.965 -58.2 47.315 -58.08 ;
      RECT 46.965 -54.97 47.315 -54.85 ;
      RECT 46.965 -51.74 47.315 -51.62 ;
      RECT 46.965 -48.51 47.315 -48.39 ;
      RECT 46.965 -45.28 47.315 -45.16 ;
      RECT 46.965 -42.05 47.315 -41.93 ;
      RECT 46.965 -38.82 47.315 -38.7 ;
      RECT 46.965 -35.59 47.315 -35.47 ;
      RECT 46.965 -32.36 47.315 -32.24 ;
      RECT 46.965 -29.13 47.315 -29.01 ;
      RECT 46.965 -25.9 47.315 -25.78 ;
      RECT 46.965 -22.67 47.315 -22.55 ;
      RECT 46.965 -19.44 47.315 -19.32 ;
      RECT 46.965 -16.21 47.315 -16.09 ;
      RECT 46.965 -12.98 47.315 -12.86 ;
      RECT 46.965 -9.75 47.315 -9.63 ;
      RECT 46.965 -6.52 47.315 -6.4 ;
      RECT 46.965 -3.29 47.315 -3.17 ;
      RECT 46.965 -0.06 47.315 0.06 ;
      RECT 47.135 -104.945 47.235 -103.985 ;
      RECT 47.135 2.175 47.235 3.135 ;
      RECT 43.235 -108.655 47.015 -108.535 ;
      RECT 46.875 -104.945 46.975 -103.985 ;
      RECT 46.75 -101.06 46.85 -100.525 ;
      RECT 46.75 -99.735 46.85 -99.2 ;
      RECT 46.75 -97.83 46.85 -97.295 ;
      RECT 46.75 -96.505 46.85 -95.97 ;
      RECT 46.75 -94.6 46.85 -94.065 ;
      RECT 46.75 -93.275 46.85 -92.74 ;
      RECT 46.75 -91.37 46.85 -90.835 ;
      RECT 46.75 -90.045 46.85 -89.51 ;
      RECT 46.75 -88.14 46.85 -87.605 ;
      RECT 46.75 -86.815 46.85 -86.28 ;
      RECT 46.75 -84.91 46.85 -84.375 ;
      RECT 46.75 -83.585 46.85 -83.05 ;
      RECT 46.75 -81.68 46.85 -81.145 ;
      RECT 46.75 -80.355 46.85 -79.82 ;
      RECT 46.75 -78.45 46.85 -77.915 ;
      RECT 46.75 -77.125 46.85 -76.59 ;
      RECT 46.75 -75.22 46.85 -74.685 ;
      RECT 46.75 -73.895 46.85 -73.36 ;
      RECT 46.75 -71.99 46.85 -71.455 ;
      RECT 46.75 -70.665 46.85 -70.13 ;
      RECT 46.75 -68.76 46.85 -68.225 ;
      RECT 46.75 -67.435 46.85 -66.9 ;
      RECT 46.75 -65.53 46.85 -64.995 ;
      RECT 46.75 -64.205 46.85 -63.67 ;
      RECT 46.75 -62.3 46.85 -61.765 ;
      RECT 46.75 -60.975 46.85 -60.44 ;
      RECT 46.75 -59.07 46.85 -58.535 ;
      RECT 46.75 -57.745 46.85 -57.21 ;
      RECT 46.75 -55.84 46.85 -55.305 ;
      RECT 46.75 -54.515 46.85 -53.98 ;
      RECT 46.75 -52.61 46.85 -52.075 ;
      RECT 46.75 -51.285 46.85 -50.75 ;
      RECT 46.75 -49.38 46.85 -48.845 ;
      RECT 46.75 -48.055 46.85 -47.52 ;
      RECT 46.75 -46.15 46.85 -45.615 ;
      RECT 46.75 -44.825 46.85 -44.29 ;
      RECT 46.75 -42.92 46.85 -42.385 ;
      RECT 46.75 -41.595 46.85 -41.06 ;
      RECT 46.75 -39.69 46.85 -39.155 ;
      RECT 46.75 -38.365 46.85 -37.83 ;
      RECT 46.75 -36.46 46.85 -35.925 ;
      RECT 46.75 -35.135 46.85 -34.6 ;
      RECT 46.75 -33.23 46.85 -32.695 ;
      RECT 46.75 -31.905 46.85 -31.37 ;
      RECT 46.75 -30 46.85 -29.465 ;
      RECT 46.75 -28.675 46.85 -28.14 ;
      RECT 46.75 -26.77 46.85 -26.235 ;
      RECT 46.75 -25.445 46.85 -24.91 ;
      RECT 46.75 -23.54 46.85 -23.005 ;
      RECT 46.75 -22.215 46.85 -21.68 ;
      RECT 46.75 -20.31 46.85 -19.775 ;
      RECT 46.75 -18.985 46.85 -18.45 ;
      RECT 46.75 -17.08 46.85 -16.545 ;
      RECT 46.75 -15.755 46.85 -15.22 ;
      RECT 46.75 -13.85 46.85 -13.315 ;
      RECT 46.75 -12.525 46.85 -11.99 ;
      RECT 46.75 -10.62 46.85 -10.085 ;
      RECT 46.75 -9.295 46.85 -8.76 ;
      RECT 46.75 -7.39 46.85 -6.855 ;
      RECT 46.75 -6.065 46.85 -5.53 ;
      RECT 46.75 -4.16 46.85 -3.625 ;
      RECT 46.75 -2.835 46.85 -2.3 ;
      RECT 46.75 -0.93 46.85 -0.395 ;
      RECT 46.75 0.395 46.85 0.93 ;
      RECT 46.685 -110.75 46.805 -110.37 ;
      RECT 46.685 -112.245 46.785 -111.775 ;
      RECT 46.625 -104.945 46.725 -103.985 ;
      RECT 46.25 -100.19 46.6 -100.07 ;
      RECT 46.25 -96.96 46.6 -96.84 ;
      RECT 46.25 -93.73 46.6 -93.61 ;
      RECT 46.25 -90.5 46.6 -90.38 ;
      RECT 46.25 -87.27 46.6 -87.15 ;
      RECT 46.25 -84.04 46.6 -83.92 ;
      RECT 46.25 -80.81 46.6 -80.69 ;
      RECT 46.25 -77.58 46.6 -77.46 ;
      RECT 46.25 -74.35 46.6 -74.23 ;
      RECT 46.25 -71.12 46.6 -71 ;
      RECT 46.25 -67.89 46.6 -67.77 ;
      RECT 46.25 -64.66 46.6 -64.54 ;
      RECT 46.25 -61.43 46.6 -61.31 ;
      RECT 46.25 -58.2 46.6 -58.08 ;
      RECT 46.25 -54.97 46.6 -54.85 ;
      RECT 46.25 -51.74 46.6 -51.62 ;
      RECT 46.25 -48.51 46.6 -48.39 ;
      RECT 46.25 -45.28 46.6 -45.16 ;
      RECT 46.25 -42.05 46.6 -41.93 ;
      RECT 46.25 -38.82 46.6 -38.7 ;
      RECT 46.25 -35.59 46.6 -35.47 ;
      RECT 46.25 -32.36 46.6 -32.24 ;
      RECT 46.25 -29.13 46.6 -29.01 ;
      RECT 46.25 -25.9 46.6 -25.78 ;
      RECT 46.25 -22.67 46.6 -22.55 ;
      RECT 46.25 -19.44 46.6 -19.32 ;
      RECT 46.25 -16.21 46.6 -16.09 ;
      RECT 46.25 -12.98 46.6 -12.86 ;
      RECT 46.25 -9.75 46.6 -9.63 ;
      RECT 46.25 -6.52 46.6 -6.4 ;
      RECT 46.25 -3.29 46.6 -3.17 ;
      RECT 46.25 -0.06 46.6 0.06 ;
      RECT 46.365 -104.945 46.465 -103.985 ;
      RECT 46.365 2.175 46.465 3.135 ;
      RECT 46.095 -109.595 46.23 -109.275 ;
      RECT 45.765 -100.19 46.115 -100.07 ;
      RECT 45.765 -96.96 46.115 -96.84 ;
      RECT 45.765 -93.73 46.115 -93.61 ;
      RECT 45.765 -90.5 46.115 -90.38 ;
      RECT 45.765 -87.27 46.115 -87.15 ;
      RECT 45.765 -84.04 46.115 -83.92 ;
      RECT 45.765 -80.81 46.115 -80.69 ;
      RECT 45.765 -77.58 46.115 -77.46 ;
      RECT 45.765 -74.35 46.115 -74.23 ;
      RECT 45.765 -71.12 46.115 -71 ;
      RECT 45.765 -67.89 46.115 -67.77 ;
      RECT 45.765 -64.66 46.115 -64.54 ;
      RECT 45.765 -61.43 46.115 -61.31 ;
      RECT 45.765 -58.2 46.115 -58.08 ;
      RECT 45.765 -54.97 46.115 -54.85 ;
      RECT 45.765 -51.74 46.115 -51.62 ;
      RECT 45.765 -48.51 46.115 -48.39 ;
      RECT 45.765 -45.28 46.115 -45.16 ;
      RECT 45.765 -42.05 46.115 -41.93 ;
      RECT 45.765 -38.82 46.115 -38.7 ;
      RECT 45.765 -35.59 46.115 -35.47 ;
      RECT 45.765 -32.36 46.115 -32.24 ;
      RECT 45.765 -29.13 46.115 -29.01 ;
      RECT 45.765 -25.9 46.115 -25.78 ;
      RECT 45.765 -22.67 46.115 -22.55 ;
      RECT 45.765 -19.44 46.115 -19.32 ;
      RECT 45.765 -16.21 46.115 -16.09 ;
      RECT 45.765 -12.98 46.115 -12.86 ;
      RECT 45.765 -9.75 46.115 -9.63 ;
      RECT 45.765 -6.52 46.115 -6.4 ;
      RECT 45.765 -3.29 46.115 -3.17 ;
      RECT 45.765 -0.06 46.115 0.06 ;
      RECT 45.935 -104.945 46.035 -103.985 ;
      RECT 45.935 2.175 46.035 3.135 ;
      RECT 45.76 -109.595 45.905 -109.275 ;
      RECT 45.675 -104.945 45.775 -103.985 ;
      RECT 45.55 -101.06 45.65 -100.525 ;
      RECT 45.55 -99.735 45.65 -99.2 ;
      RECT 45.55 -97.83 45.65 -97.295 ;
      RECT 45.55 -96.505 45.65 -95.97 ;
      RECT 45.55 -94.6 45.65 -94.065 ;
      RECT 45.55 -93.275 45.65 -92.74 ;
      RECT 45.55 -91.37 45.65 -90.835 ;
      RECT 45.55 -90.045 45.65 -89.51 ;
      RECT 45.55 -88.14 45.65 -87.605 ;
      RECT 45.55 -86.815 45.65 -86.28 ;
      RECT 45.55 -84.91 45.65 -84.375 ;
      RECT 45.55 -83.585 45.65 -83.05 ;
      RECT 45.55 -81.68 45.65 -81.145 ;
      RECT 45.55 -80.355 45.65 -79.82 ;
      RECT 45.55 -78.45 45.65 -77.915 ;
      RECT 45.55 -77.125 45.65 -76.59 ;
      RECT 45.55 -75.22 45.65 -74.685 ;
      RECT 45.55 -73.895 45.65 -73.36 ;
      RECT 45.55 -71.99 45.65 -71.455 ;
      RECT 45.55 -70.665 45.65 -70.13 ;
      RECT 45.55 -68.76 45.65 -68.225 ;
      RECT 45.55 -67.435 45.65 -66.9 ;
      RECT 45.55 -65.53 45.65 -64.995 ;
      RECT 45.55 -64.205 45.65 -63.67 ;
      RECT 45.55 -62.3 45.65 -61.765 ;
      RECT 45.55 -60.975 45.65 -60.44 ;
      RECT 45.55 -59.07 45.65 -58.535 ;
      RECT 45.55 -57.745 45.65 -57.21 ;
      RECT 45.55 -55.84 45.65 -55.305 ;
      RECT 45.55 -54.515 45.65 -53.98 ;
      RECT 45.55 -52.61 45.65 -52.075 ;
      RECT 45.55 -51.285 45.65 -50.75 ;
      RECT 45.55 -49.38 45.65 -48.845 ;
      RECT 45.55 -48.055 45.65 -47.52 ;
      RECT 45.55 -46.15 45.65 -45.615 ;
      RECT 45.55 -44.825 45.65 -44.29 ;
      RECT 45.55 -42.92 45.65 -42.385 ;
      RECT 45.55 -41.595 45.65 -41.06 ;
      RECT 45.55 -39.69 45.65 -39.155 ;
      RECT 45.55 -38.365 45.65 -37.83 ;
      RECT 45.55 -36.46 45.65 -35.925 ;
      RECT 45.55 -35.135 45.65 -34.6 ;
      RECT 45.55 -33.23 45.65 -32.695 ;
      RECT 45.55 -31.905 45.65 -31.37 ;
      RECT 45.55 -30 45.65 -29.465 ;
      RECT 45.55 -28.675 45.65 -28.14 ;
      RECT 45.55 -26.77 45.65 -26.235 ;
      RECT 45.55 -25.445 45.65 -24.91 ;
      RECT 45.55 -23.54 45.65 -23.005 ;
      RECT 45.55 -22.215 45.65 -21.68 ;
      RECT 45.55 -20.31 45.65 -19.775 ;
      RECT 45.55 -18.985 45.65 -18.45 ;
      RECT 45.55 -17.08 45.65 -16.545 ;
      RECT 45.55 -15.755 45.65 -15.22 ;
      RECT 45.55 -13.85 45.65 -13.315 ;
      RECT 45.55 -12.525 45.65 -11.99 ;
      RECT 45.55 -10.62 45.65 -10.085 ;
      RECT 45.55 -9.295 45.65 -8.76 ;
      RECT 45.55 -7.39 45.65 -6.855 ;
      RECT 45.55 -6.065 45.65 -5.53 ;
      RECT 45.55 -4.16 45.65 -3.625 ;
      RECT 45.55 -2.835 45.65 -2.3 ;
      RECT 45.55 -0.93 45.65 -0.395 ;
      RECT 45.55 0.395 45.65 0.93 ;
      RECT 45.425 -108.175 45.525 -107.215 ;
      RECT 45.05 -100.19 45.4 -100.07 ;
      RECT 45.05 -96.96 45.4 -96.84 ;
      RECT 45.05 -93.73 45.4 -93.61 ;
      RECT 45.05 -90.5 45.4 -90.38 ;
      RECT 45.05 -87.27 45.4 -87.15 ;
      RECT 45.05 -84.04 45.4 -83.92 ;
      RECT 45.05 -80.81 45.4 -80.69 ;
      RECT 45.05 -77.58 45.4 -77.46 ;
      RECT 45.05 -74.35 45.4 -74.23 ;
      RECT 45.05 -71.12 45.4 -71 ;
      RECT 45.05 -67.89 45.4 -67.77 ;
      RECT 45.05 -64.66 45.4 -64.54 ;
      RECT 45.05 -61.43 45.4 -61.31 ;
      RECT 45.05 -58.2 45.4 -58.08 ;
      RECT 45.05 -54.97 45.4 -54.85 ;
      RECT 45.05 -51.74 45.4 -51.62 ;
      RECT 45.05 -48.51 45.4 -48.39 ;
      RECT 45.05 -45.28 45.4 -45.16 ;
      RECT 45.05 -42.05 45.4 -41.93 ;
      RECT 45.05 -38.82 45.4 -38.7 ;
      RECT 45.05 -35.59 45.4 -35.47 ;
      RECT 45.05 -32.36 45.4 -32.24 ;
      RECT 45.05 -29.13 45.4 -29.01 ;
      RECT 45.05 -25.9 45.4 -25.78 ;
      RECT 45.05 -22.67 45.4 -22.55 ;
      RECT 45.05 -19.44 45.4 -19.32 ;
      RECT 45.05 -16.21 45.4 -16.09 ;
      RECT 45.05 -12.98 45.4 -12.86 ;
      RECT 45.05 -9.75 45.4 -9.63 ;
      RECT 45.05 -6.52 45.4 -6.4 ;
      RECT 45.05 -3.29 45.4 -3.17 ;
      RECT 45.05 -0.06 45.4 0.06 ;
      RECT 45.255 -112.255 45.355 -111.775 ;
      RECT 45.255 -110.765 45.355 -110.295 ;
      RECT 45.165 -108.175 45.265 -107.215 ;
      RECT 45.165 2.175 45.265 3.135 ;
      RECT 44.565 -100.19 44.915 -100.07 ;
      RECT 44.565 -96.96 44.915 -96.84 ;
      RECT 44.565 -93.73 44.915 -93.61 ;
      RECT 44.565 -90.5 44.915 -90.38 ;
      RECT 44.565 -87.27 44.915 -87.15 ;
      RECT 44.565 -84.04 44.915 -83.92 ;
      RECT 44.565 -80.81 44.915 -80.69 ;
      RECT 44.565 -77.58 44.915 -77.46 ;
      RECT 44.565 -74.35 44.915 -74.23 ;
      RECT 44.565 -71.12 44.915 -71 ;
      RECT 44.565 -67.89 44.915 -67.77 ;
      RECT 44.565 -64.66 44.915 -64.54 ;
      RECT 44.565 -61.43 44.915 -61.31 ;
      RECT 44.565 -58.2 44.915 -58.08 ;
      RECT 44.565 -54.97 44.915 -54.85 ;
      RECT 44.565 -51.74 44.915 -51.62 ;
      RECT 44.565 -48.51 44.915 -48.39 ;
      RECT 44.565 -45.28 44.915 -45.16 ;
      RECT 44.565 -42.05 44.915 -41.93 ;
      RECT 44.565 -38.82 44.915 -38.7 ;
      RECT 44.565 -35.59 44.915 -35.47 ;
      RECT 44.565 -32.36 44.915 -32.24 ;
      RECT 44.565 -29.13 44.915 -29.01 ;
      RECT 44.565 -25.9 44.915 -25.78 ;
      RECT 44.565 -22.67 44.915 -22.55 ;
      RECT 44.565 -19.44 44.915 -19.32 ;
      RECT 44.565 -16.21 44.915 -16.09 ;
      RECT 44.565 -12.98 44.915 -12.86 ;
      RECT 44.565 -9.75 44.915 -9.63 ;
      RECT 44.565 -6.52 44.915 -6.4 ;
      RECT 44.565 -3.29 44.915 -3.17 ;
      RECT 44.565 -0.06 44.915 0.06 ;
      RECT 44.735 -108.175 44.835 -107.215 ;
      RECT 44.735 2.175 44.835 3.135 ;
      RECT 44.63 -110.765 44.8 -110.385 ;
      RECT 44.665 -112.245 44.765 -111.775 ;
      RECT 44.475 -108.175 44.575 -107.215 ;
      RECT 44.35 -101.06 44.45 -100.525 ;
      RECT 44.35 -99.735 44.45 -99.2 ;
      RECT 44.35 -97.83 44.45 -97.295 ;
      RECT 44.35 -96.505 44.45 -95.97 ;
      RECT 44.35 -94.6 44.45 -94.065 ;
      RECT 44.35 -93.275 44.45 -92.74 ;
      RECT 44.35 -91.37 44.45 -90.835 ;
      RECT 44.35 -90.045 44.45 -89.51 ;
      RECT 44.35 -88.14 44.45 -87.605 ;
      RECT 44.35 -86.815 44.45 -86.28 ;
      RECT 44.35 -84.91 44.45 -84.375 ;
      RECT 44.35 -83.585 44.45 -83.05 ;
      RECT 44.35 -81.68 44.45 -81.145 ;
      RECT 44.35 -80.355 44.45 -79.82 ;
      RECT 44.35 -78.45 44.45 -77.915 ;
      RECT 44.35 -77.125 44.45 -76.59 ;
      RECT 44.35 -75.22 44.45 -74.685 ;
      RECT 44.35 -73.895 44.45 -73.36 ;
      RECT 44.35 -71.99 44.45 -71.455 ;
      RECT 44.35 -70.665 44.45 -70.13 ;
      RECT 44.35 -68.76 44.45 -68.225 ;
      RECT 44.35 -67.435 44.45 -66.9 ;
      RECT 44.35 -65.53 44.45 -64.995 ;
      RECT 44.35 -64.205 44.45 -63.67 ;
      RECT 44.35 -62.3 44.45 -61.765 ;
      RECT 44.35 -60.975 44.45 -60.44 ;
      RECT 44.35 -59.07 44.45 -58.535 ;
      RECT 44.35 -57.745 44.45 -57.21 ;
      RECT 44.35 -55.84 44.45 -55.305 ;
      RECT 44.35 -54.515 44.45 -53.98 ;
      RECT 44.35 -52.61 44.45 -52.075 ;
      RECT 44.35 -51.285 44.45 -50.75 ;
      RECT 44.35 -49.38 44.45 -48.845 ;
      RECT 44.35 -48.055 44.45 -47.52 ;
      RECT 44.35 -46.15 44.45 -45.615 ;
      RECT 44.35 -44.825 44.45 -44.29 ;
      RECT 44.35 -42.92 44.45 -42.385 ;
      RECT 44.35 -41.595 44.45 -41.06 ;
      RECT 44.35 -39.69 44.45 -39.155 ;
      RECT 44.35 -38.365 44.45 -37.83 ;
      RECT 44.35 -36.46 44.45 -35.925 ;
      RECT 44.35 -35.135 44.45 -34.6 ;
      RECT 44.35 -33.23 44.45 -32.695 ;
      RECT 44.35 -31.905 44.45 -31.37 ;
      RECT 44.35 -30 44.45 -29.465 ;
      RECT 44.35 -28.675 44.45 -28.14 ;
      RECT 44.35 -26.77 44.45 -26.235 ;
      RECT 44.35 -25.445 44.45 -24.91 ;
      RECT 44.35 -23.54 44.45 -23.005 ;
      RECT 44.35 -22.215 44.45 -21.68 ;
      RECT 44.35 -20.31 44.45 -19.775 ;
      RECT 44.35 -18.985 44.45 -18.45 ;
      RECT 44.35 -17.08 44.45 -16.545 ;
      RECT 44.35 -15.755 44.45 -15.22 ;
      RECT 44.35 -13.85 44.45 -13.315 ;
      RECT 44.35 -12.525 44.45 -11.99 ;
      RECT 44.35 -10.62 44.45 -10.085 ;
      RECT 44.35 -9.295 44.45 -8.76 ;
      RECT 44.35 -7.39 44.45 -6.855 ;
      RECT 44.35 -6.065 44.45 -5.53 ;
      RECT 44.35 -4.16 44.45 -3.625 ;
      RECT 44.35 -2.835 44.45 -2.3 ;
      RECT 44.35 -0.93 44.45 -0.395 ;
      RECT 44.35 0.395 44.45 0.93 ;
      RECT 44.225 -108.175 44.325 -107.215 ;
      RECT 43.85 -100.19 44.2 -100.07 ;
      RECT 43.85 -96.96 44.2 -96.84 ;
      RECT 43.85 -93.73 44.2 -93.61 ;
      RECT 43.85 -90.5 44.2 -90.38 ;
      RECT 43.85 -87.27 44.2 -87.15 ;
      RECT 43.85 -84.04 44.2 -83.92 ;
      RECT 43.85 -80.81 44.2 -80.69 ;
      RECT 43.85 -77.58 44.2 -77.46 ;
      RECT 43.85 -74.35 44.2 -74.23 ;
      RECT 43.85 -71.12 44.2 -71 ;
      RECT 43.85 -67.89 44.2 -67.77 ;
      RECT 43.85 -64.66 44.2 -64.54 ;
      RECT 43.85 -61.43 44.2 -61.31 ;
      RECT 43.85 -58.2 44.2 -58.08 ;
      RECT 43.85 -54.97 44.2 -54.85 ;
      RECT 43.85 -51.74 44.2 -51.62 ;
      RECT 43.85 -48.51 44.2 -48.39 ;
      RECT 43.85 -45.28 44.2 -45.16 ;
      RECT 43.85 -42.05 44.2 -41.93 ;
      RECT 43.85 -38.82 44.2 -38.7 ;
      RECT 43.85 -35.59 44.2 -35.47 ;
      RECT 43.85 -32.36 44.2 -32.24 ;
      RECT 43.85 -29.13 44.2 -29.01 ;
      RECT 43.85 -25.9 44.2 -25.78 ;
      RECT 43.85 -22.67 44.2 -22.55 ;
      RECT 43.85 -19.44 44.2 -19.32 ;
      RECT 43.85 -16.21 44.2 -16.09 ;
      RECT 43.85 -12.98 44.2 -12.86 ;
      RECT 43.85 -9.75 44.2 -9.63 ;
      RECT 43.85 -6.52 44.2 -6.4 ;
      RECT 43.85 -3.29 44.2 -3.17 ;
      RECT 43.85 -0.06 44.2 0.06 ;
      RECT 43.965 -108.175 44.065 -107.215 ;
      RECT 43.965 2.175 44.065 3.135 ;
      RECT 43.865 -113.555 43.965 -113.085 ;
      RECT 43.365 -100.19 43.715 -100.07 ;
      RECT 43.365 -96.96 43.715 -96.84 ;
      RECT 43.365 -93.73 43.715 -93.61 ;
      RECT 43.365 -90.5 43.715 -90.38 ;
      RECT 43.365 -87.27 43.715 -87.15 ;
      RECT 43.365 -84.04 43.715 -83.92 ;
      RECT 43.365 -80.81 43.715 -80.69 ;
      RECT 43.365 -77.58 43.715 -77.46 ;
      RECT 43.365 -74.35 43.715 -74.23 ;
      RECT 43.365 -71.12 43.715 -71 ;
      RECT 43.365 -67.89 43.715 -67.77 ;
      RECT 43.365 -64.66 43.715 -64.54 ;
      RECT 43.365 -61.43 43.715 -61.31 ;
      RECT 43.365 -58.2 43.715 -58.08 ;
      RECT 43.365 -54.97 43.715 -54.85 ;
      RECT 43.365 -51.74 43.715 -51.62 ;
      RECT 43.365 -48.51 43.715 -48.39 ;
      RECT 43.365 -45.28 43.715 -45.16 ;
      RECT 43.365 -42.05 43.715 -41.93 ;
      RECT 43.365 -38.82 43.715 -38.7 ;
      RECT 43.365 -35.59 43.715 -35.47 ;
      RECT 43.365 -32.36 43.715 -32.24 ;
      RECT 43.365 -29.13 43.715 -29.01 ;
      RECT 43.365 -25.9 43.715 -25.78 ;
      RECT 43.365 -22.67 43.715 -22.55 ;
      RECT 43.365 -19.44 43.715 -19.32 ;
      RECT 43.365 -16.21 43.715 -16.09 ;
      RECT 43.365 -12.98 43.715 -12.86 ;
      RECT 43.365 -9.75 43.715 -9.63 ;
      RECT 43.365 -6.52 43.715 -6.4 ;
      RECT 43.365 -3.29 43.715 -3.17 ;
      RECT 43.365 -0.06 43.715 0.06 ;
      RECT 43.5 -110.735 43.65 -110.445 ;
      RECT 43.535 -108.175 43.635 -107.215 ;
      RECT 43.535 2.175 43.635 3.135 ;
      RECT 43.515 -112.19 43.615 -111.65 ;
      RECT 43.275 -113.555 43.375 -113.085 ;
      RECT 43.275 -108.175 43.375 -107.215 ;
      RECT 43.15 -101.06 43.25 -100.525 ;
      RECT 43.15 -99.735 43.25 -99.2 ;
      RECT 43.15 -97.83 43.25 -97.295 ;
      RECT 43.15 -96.505 43.25 -95.97 ;
      RECT 43.15 -94.6 43.25 -94.065 ;
      RECT 43.15 -93.275 43.25 -92.74 ;
      RECT 43.15 -91.37 43.25 -90.835 ;
      RECT 43.15 -90.045 43.25 -89.51 ;
      RECT 43.15 -88.14 43.25 -87.605 ;
      RECT 43.15 -86.815 43.25 -86.28 ;
      RECT 43.15 -84.91 43.25 -84.375 ;
      RECT 43.15 -83.585 43.25 -83.05 ;
      RECT 43.15 -81.68 43.25 -81.145 ;
      RECT 43.15 -80.355 43.25 -79.82 ;
      RECT 43.15 -78.45 43.25 -77.915 ;
      RECT 43.15 -77.125 43.25 -76.59 ;
      RECT 43.15 -75.22 43.25 -74.685 ;
      RECT 43.15 -73.895 43.25 -73.36 ;
      RECT 43.15 -71.99 43.25 -71.455 ;
      RECT 43.15 -70.665 43.25 -70.13 ;
      RECT 43.15 -68.76 43.25 -68.225 ;
      RECT 43.15 -67.435 43.25 -66.9 ;
      RECT 43.15 -65.53 43.25 -64.995 ;
      RECT 43.15 -64.205 43.25 -63.67 ;
      RECT 43.15 -62.3 43.25 -61.765 ;
      RECT 43.15 -60.975 43.25 -60.44 ;
      RECT 43.15 -59.07 43.25 -58.535 ;
      RECT 43.15 -57.745 43.25 -57.21 ;
      RECT 43.15 -55.84 43.25 -55.305 ;
      RECT 43.15 -54.515 43.25 -53.98 ;
      RECT 43.15 -52.61 43.25 -52.075 ;
      RECT 43.15 -51.285 43.25 -50.75 ;
      RECT 43.15 -49.38 43.25 -48.845 ;
      RECT 43.15 -48.055 43.25 -47.52 ;
      RECT 43.15 -46.15 43.25 -45.615 ;
      RECT 43.15 -44.825 43.25 -44.29 ;
      RECT 43.15 -42.92 43.25 -42.385 ;
      RECT 43.15 -41.595 43.25 -41.06 ;
      RECT 43.15 -39.69 43.25 -39.155 ;
      RECT 43.15 -38.365 43.25 -37.83 ;
      RECT 43.15 -36.46 43.25 -35.925 ;
      RECT 43.15 -35.135 43.25 -34.6 ;
      RECT 43.15 -33.23 43.25 -32.695 ;
      RECT 43.15 -31.905 43.25 -31.37 ;
      RECT 43.15 -30 43.25 -29.465 ;
      RECT 43.15 -28.675 43.25 -28.14 ;
      RECT 43.15 -26.77 43.25 -26.235 ;
      RECT 43.15 -25.445 43.25 -24.91 ;
      RECT 43.15 -23.54 43.25 -23.005 ;
      RECT 43.15 -22.215 43.25 -21.68 ;
      RECT 43.15 -20.31 43.25 -19.775 ;
      RECT 43.15 -18.985 43.25 -18.45 ;
      RECT 43.15 -17.08 43.25 -16.545 ;
      RECT 43.15 -15.755 43.25 -15.22 ;
      RECT 43.15 -13.85 43.25 -13.315 ;
      RECT 43.15 -12.525 43.25 -11.99 ;
      RECT 43.15 -10.62 43.25 -10.085 ;
      RECT 43.15 -9.295 43.25 -8.76 ;
      RECT 43.15 -7.39 43.25 -6.855 ;
      RECT 43.15 -6.065 43.25 -5.53 ;
      RECT 43.15 -4.16 43.25 -3.625 ;
      RECT 43.15 -2.835 43.25 -2.3 ;
      RECT 43.15 -0.93 43.25 -0.395 ;
      RECT 43.15 0.395 43.25 0.93 ;
      RECT 43.025 -104.945 43.125 -103.985 ;
      RECT 42.65 -100.19 43 -100.07 ;
      RECT 42.65 -96.96 43 -96.84 ;
      RECT 42.65 -93.73 43 -93.61 ;
      RECT 42.65 -90.5 43 -90.38 ;
      RECT 42.65 -87.27 43 -87.15 ;
      RECT 42.65 -84.04 43 -83.92 ;
      RECT 42.65 -80.81 43 -80.69 ;
      RECT 42.65 -77.58 43 -77.46 ;
      RECT 42.65 -74.35 43 -74.23 ;
      RECT 42.65 -71.12 43 -71 ;
      RECT 42.65 -67.89 43 -67.77 ;
      RECT 42.65 -64.66 43 -64.54 ;
      RECT 42.65 -61.43 43 -61.31 ;
      RECT 42.65 -58.2 43 -58.08 ;
      RECT 42.65 -54.97 43 -54.85 ;
      RECT 42.65 -51.74 43 -51.62 ;
      RECT 42.65 -48.51 43 -48.39 ;
      RECT 42.65 -45.28 43 -45.16 ;
      RECT 42.65 -42.05 43 -41.93 ;
      RECT 42.65 -38.82 43 -38.7 ;
      RECT 42.65 -35.59 43 -35.47 ;
      RECT 42.65 -32.36 43 -32.24 ;
      RECT 42.65 -29.13 43 -29.01 ;
      RECT 42.65 -25.9 43 -25.78 ;
      RECT 42.65 -22.67 43 -22.55 ;
      RECT 42.65 -19.44 43 -19.32 ;
      RECT 42.65 -16.21 43 -16.09 ;
      RECT 42.65 -12.98 43 -12.86 ;
      RECT 42.65 -9.75 43 -9.63 ;
      RECT 42.65 -6.52 43 -6.4 ;
      RECT 42.65 -3.29 43 -3.17 ;
      RECT 42.65 -0.06 43 0.06 ;
      RECT 42.765 -104.945 42.865 -103.985 ;
      RECT 42.765 2.175 42.865 3.135 ;
      RECT 42.475 -112.255 42.575 -111.775 ;
      RECT 42.475 -110.765 42.575 -110.295 ;
      RECT 42.165 -100.19 42.515 -100.07 ;
      RECT 42.165 -96.96 42.515 -96.84 ;
      RECT 42.165 -93.73 42.515 -93.61 ;
      RECT 42.165 -90.5 42.515 -90.38 ;
      RECT 42.165 -87.27 42.515 -87.15 ;
      RECT 42.165 -84.04 42.515 -83.92 ;
      RECT 42.165 -80.81 42.515 -80.69 ;
      RECT 42.165 -77.58 42.515 -77.46 ;
      RECT 42.165 -74.35 42.515 -74.23 ;
      RECT 42.165 -71.12 42.515 -71 ;
      RECT 42.165 -67.89 42.515 -67.77 ;
      RECT 42.165 -64.66 42.515 -64.54 ;
      RECT 42.165 -61.43 42.515 -61.31 ;
      RECT 42.165 -58.2 42.515 -58.08 ;
      RECT 42.165 -54.97 42.515 -54.85 ;
      RECT 42.165 -51.74 42.515 -51.62 ;
      RECT 42.165 -48.51 42.515 -48.39 ;
      RECT 42.165 -45.28 42.515 -45.16 ;
      RECT 42.165 -42.05 42.515 -41.93 ;
      RECT 42.165 -38.82 42.515 -38.7 ;
      RECT 42.165 -35.59 42.515 -35.47 ;
      RECT 42.165 -32.36 42.515 -32.24 ;
      RECT 42.165 -29.13 42.515 -29.01 ;
      RECT 42.165 -25.9 42.515 -25.78 ;
      RECT 42.165 -22.67 42.515 -22.55 ;
      RECT 42.165 -19.44 42.515 -19.32 ;
      RECT 42.165 -16.21 42.515 -16.09 ;
      RECT 42.165 -12.98 42.515 -12.86 ;
      RECT 42.165 -9.75 42.515 -9.63 ;
      RECT 42.165 -6.52 42.515 -6.4 ;
      RECT 42.165 -3.29 42.515 -3.17 ;
      RECT 42.165 -0.06 42.515 0.06 ;
      RECT 42.335 -104.945 42.435 -103.985 ;
      RECT 42.335 2.175 42.435 3.135 ;
      RECT 38.435 -108.655 42.215 -108.535 ;
      RECT 42.075 -104.945 42.175 -103.985 ;
      RECT 41.95 -101.06 42.05 -100.525 ;
      RECT 41.95 -99.735 42.05 -99.2 ;
      RECT 41.95 -97.83 42.05 -97.295 ;
      RECT 41.95 -96.505 42.05 -95.97 ;
      RECT 41.95 -94.6 42.05 -94.065 ;
      RECT 41.95 -93.275 42.05 -92.74 ;
      RECT 41.95 -91.37 42.05 -90.835 ;
      RECT 41.95 -90.045 42.05 -89.51 ;
      RECT 41.95 -88.14 42.05 -87.605 ;
      RECT 41.95 -86.815 42.05 -86.28 ;
      RECT 41.95 -84.91 42.05 -84.375 ;
      RECT 41.95 -83.585 42.05 -83.05 ;
      RECT 41.95 -81.68 42.05 -81.145 ;
      RECT 41.95 -80.355 42.05 -79.82 ;
      RECT 41.95 -78.45 42.05 -77.915 ;
      RECT 41.95 -77.125 42.05 -76.59 ;
      RECT 41.95 -75.22 42.05 -74.685 ;
      RECT 41.95 -73.895 42.05 -73.36 ;
      RECT 41.95 -71.99 42.05 -71.455 ;
      RECT 41.95 -70.665 42.05 -70.13 ;
      RECT 41.95 -68.76 42.05 -68.225 ;
      RECT 41.95 -67.435 42.05 -66.9 ;
      RECT 41.95 -65.53 42.05 -64.995 ;
      RECT 41.95 -64.205 42.05 -63.67 ;
      RECT 41.95 -62.3 42.05 -61.765 ;
      RECT 41.95 -60.975 42.05 -60.44 ;
      RECT 41.95 -59.07 42.05 -58.535 ;
      RECT 41.95 -57.745 42.05 -57.21 ;
      RECT 41.95 -55.84 42.05 -55.305 ;
      RECT 41.95 -54.515 42.05 -53.98 ;
      RECT 41.95 -52.61 42.05 -52.075 ;
      RECT 41.95 -51.285 42.05 -50.75 ;
      RECT 41.95 -49.38 42.05 -48.845 ;
      RECT 41.95 -48.055 42.05 -47.52 ;
      RECT 41.95 -46.15 42.05 -45.615 ;
      RECT 41.95 -44.825 42.05 -44.29 ;
      RECT 41.95 -42.92 42.05 -42.385 ;
      RECT 41.95 -41.595 42.05 -41.06 ;
      RECT 41.95 -39.69 42.05 -39.155 ;
      RECT 41.95 -38.365 42.05 -37.83 ;
      RECT 41.95 -36.46 42.05 -35.925 ;
      RECT 41.95 -35.135 42.05 -34.6 ;
      RECT 41.95 -33.23 42.05 -32.695 ;
      RECT 41.95 -31.905 42.05 -31.37 ;
      RECT 41.95 -30 42.05 -29.465 ;
      RECT 41.95 -28.675 42.05 -28.14 ;
      RECT 41.95 -26.77 42.05 -26.235 ;
      RECT 41.95 -25.445 42.05 -24.91 ;
      RECT 41.95 -23.54 42.05 -23.005 ;
      RECT 41.95 -22.215 42.05 -21.68 ;
      RECT 41.95 -20.31 42.05 -19.775 ;
      RECT 41.95 -18.985 42.05 -18.45 ;
      RECT 41.95 -17.08 42.05 -16.545 ;
      RECT 41.95 -15.755 42.05 -15.22 ;
      RECT 41.95 -13.85 42.05 -13.315 ;
      RECT 41.95 -12.525 42.05 -11.99 ;
      RECT 41.95 -10.62 42.05 -10.085 ;
      RECT 41.95 -9.295 42.05 -8.76 ;
      RECT 41.95 -7.39 42.05 -6.855 ;
      RECT 41.95 -6.065 42.05 -5.53 ;
      RECT 41.95 -4.16 42.05 -3.625 ;
      RECT 41.95 -2.835 42.05 -2.3 ;
      RECT 41.95 -0.93 42.05 -0.395 ;
      RECT 41.95 0.395 42.05 0.93 ;
      RECT 41.885 -110.75 42.005 -110.37 ;
      RECT 41.885 -112.245 41.985 -111.775 ;
      RECT 41.825 -104.945 41.925 -103.985 ;
      RECT 41.45 -100.19 41.8 -100.07 ;
      RECT 41.45 -96.96 41.8 -96.84 ;
      RECT 41.45 -93.73 41.8 -93.61 ;
      RECT 41.45 -90.5 41.8 -90.38 ;
      RECT 41.45 -87.27 41.8 -87.15 ;
      RECT 41.45 -84.04 41.8 -83.92 ;
      RECT 41.45 -80.81 41.8 -80.69 ;
      RECT 41.45 -77.58 41.8 -77.46 ;
      RECT 41.45 -74.35 41.8 -74.23 ;
      RECT 41.45 -71.12 41.8 -71 ;
      RECT 41.45 -67.89 41.8 -67.77 ;
      RECT 41.45 -64.66 41.8 -64.54 ;
      RECT 41.45 -61.43 41.8 -61.31 ;
      RECT 41.45 -58.2 41.8 -58.08 ;
      RECT 41.45 -54.97 41.8 -54.85 ;
      RECT 41.45 -51.74 41.8 -51.62 ;
      RECT 41.45 -48.51 41.8 -48.39 ;
      RECT 41.45 -45.28 41.8 -45.16 ;
      RECT 41.45 -42.05 41.8 -41.93 ;
      RECT 41.45 -38.82 41.8 -38.7 ;
      RECT 41.45 -35.59 41.8 -35.47 ;
      RECT 41.45 -32.36 41.8 -32.24 ;
      RECT 41.45 -29.13 41.8 -29.01 ;
      RECT 41.45 -25.9 41.8 -25.78 ;
      RECT 41.45 -22.67 41.8 -22.55 ;
      RECT 41.45 -19.44 41.8 -19.32 ;
      RECT 41.45 -16.21 41.8 -16.09 ;
      RECT 41.45 -12.98 41.8 -12.86 ;
      RECT 41.45 -9.75 41.8 -9.63 ;
      RECT 41.45 -6.52 41.8 -6.4 ;
      RECT 41.45 -3.29 41.8 -3.17 ;
      RECT 41.45 -0.06 41.8 0.06 ;
      RECT 41.565 -104.945 41.665 -103.985 ;
      RECT 41.565 2.175 41.665 3.135 ;
      RECT 41.295 -109.595 41.43 -109.275 ;
      RECT 40.965 -100.19 41.315 -100.07 ;
      RECT 40.965 -96.96 41.315 -96.84 ;
      RECT 40.965 -93.73 41.315 -93.61 ;
      RECT 40.965 -90.5 41.315 -90.38 ;
      RECT 40.965 -87.27 41.315 -87.15 ;
      RECT 40.965 -84.04 41.315 -83.92 ;
      RECT 40.965 -80.81 41.315 -80.69 ;
      RECT 40.965 -77.58 41.315 -77.46 ;
      RECT 40.965 -74.35 41.315 -74.23 ;
      RECT 40.965 -71.12 41.315 -71 ;
      RECT 40.965 -67.89 41.315 -67.77 ;
      RECT 40.965 -64.66 41.315 -64.54 ;
      RECT 40.965 -61.43 41.315 -61.31 ;
      RECT 40.965 -58.2 41.315 -58.08 ;
      RECT 40.965 -54.97 41.315 -54.85 ;
      RECT 40.965 -51.74 41.315 -51.62 ;
      RECT 40.965 -48.51 41.315 -48.39 ;
      RECT 40.965 -45.28 41.315 -45.16 ;
      RECT 40.965 -42.05 41.315 -41.93 ;
      RECT 40.965 -38.82 41.315 -38.7 ;
      RECT 40.965 -35.59 41.315 -35.47 ;
      RECT 40.965 -32.36 41.315 -32.24 ;
      RECT 40.965 -29.13 41.315 -29.01 ;
      RECT 40.965 -25.9 41.315 -25.78 ;
      RECT 40.965 -22.67 41.315 -22.55 ;
      RECT 40.965 -19.44 41.315 -19.32 ;
      RECT 40.965 -16.21 41.315 -16.09 ;
      RECT 40.965 -12.98 41.315 -12.86 ;
      RECT 40.965 -9.75 41.315 -9.63 ;
      RECT 40.965 -6.52 41.315 -6.4 ;
      RECT 40.965 -3.29 41.315 -3.17 ;
      RECT 40.965 -0.06 41.315 0.06 ;
      RECT 41.135 -104.945 41.235 -103.985 ;
      RECT 41.135 2.175 41.235 3.135 ;
      RECT 40.96 -109.595 41.105 -109.275 ;
      RECT 40.875 -104.945 40.975 -103.985 ;
      RECT 40.75 -101.06 40.85 -100.525 ;
      RECT 40.75 -99.735 40.85 -99.2 ;
      RECT 40.75 -97.83 40.85 -97.295 ;
      RECT 40.75 -96.505 40.85 -95.97 ;
      RECT 40.75 -94.6 40.85 -94.065 ;
      RECT 40.75 -93.275 40.85 -92.74 ;
      RECT 40.75 -91.37 40.85 -90.835 ;
      RECT 40.75 -90.045 40.85 -89.51 ;
      RECT 40.75 -88.14 40.85 -87.605 ;
      RECT 40.75 -86.815 40.85 -86.28 ;
      RECT 40.75 -84.91 40.85 -84.375 ;
      RECT 40.75 -83.585 40.85 -83.05 ;
      RECT 40.75 -81.68 40.85 -81.145 ;
      RECT 40.75 -80.355 40.85 -79.82 ;
      RECT 40.75 -78.45 40.85 -77.915 ;
      RECT 40.75 -77.125 40.85 -76.59 ;
      RECT 40.75 -75.22 40.85 -74.685 ;
      RECT 40.75 -73.895 40.85 -73.36 ;
      RECT 40.75 -71.99 40.85 -71.455 ;
      RECT 40.75 -70.665 40.85 -70.13 ;
      RECT 40.75 -68.76 40.85 -68.225 ;
      RECT 40.75 -67.435 40.85 -66.9 ;
      RECT 40.75 -65.53 40.85 -64.995 ;
      RECT 40.75 -64.205 40.85 -63.67 ;
      RECT 40.75 -62.3 40.85 -61.765 ;
      RECT 40.75 -60.975 40.85 -60.44 ;
      RECT 40.75 -59.07 40.85 -58.535 ;
      RECT 40.75 -57.745 40.85 -57.21 ;
      RECT 40.75 -55.84 40.85 -55.305 ;
      RECT 40.75 -54.515 40.85 -53.98 ;
      RECT 40.75 -52.61 40.85 -52.075 ;
      RECT 40.75 -51.285 40.85 -50.75 ;
      RECT 40.75 -49.38 40.85 -48.845 ;
      RECT 40.75 -48.055 40.85 -47.52 ;
      RECT 40.75 -46.15 40.85 -45.615 ;
      RECT 40.75 -44.825 40.85 -44.29 ;
      RECT 40.75 -42.92 40.85 -42.385 ;
      RECT 40.75 -41.595 40.85 -41.06 ;
      RECT 40.75 -39.69 40.85 -39.155 ;
      RECT 40.75 -38.365 40.85 -37.83 ;
      RECT 40.75 -36.46 40.85 -35.925 ;
      RECT 40.75 -35.135 40.85 -34.6 ;
      RECT 40.75 -33.23 40.85 -32.695 ;
      RECT 40.75 -31.905 40.85 -31.37 ;
      RECT 40.75 -30 40.85 -29.465 ;
      RECT 40.75 -28.675 40.85 -28.14 ;
      RECT 40.75 -26.77 40.85 -26.235 ;
      RECT 40.75 -25.445 40.85 -24.91 ;
      RECT 40.75 -23.54 40.85 -23.005 ;
      RECT 40.75 -22.215 40.85 -21.68 ;
      RECT 40.75 -20.31 40.85 -19.775 ;
      RECT 40.75 -18.985 40.85 -18.45 ;
      RECT 40.75 -17.08 40.85 -16.545 ;
      RECT 40.75 -15.755 40.85 -15.22 ;
      RECT 40.75 -13.85 40.85 -13.315 ;
      RECT 40.75 -12.525 40.85 -11.99 ;
      RECT 40.75 -10.62 40.85 -10.085 ;
      RECT 40.75 -9.295 40.85 -8.76 ;
      RECT 40.75 -7.39 40.85 -6.855 ;
      RECT 40.75 -6.065 40.85 -5.53 ;
      RECT 40.75 -4.16 40.85 -3.625 ;
      RECT 40.75 -2.835 40.85 -2.3 ;
      RECT 40.75 -0.93 40.85 -0.395 ;
      RECT 40.75 0.395 40.85 0.93 ;
      RECT 40.625 -108.175 40.725 -107.215 ;
      RECT 40.25 -100.19 40.6 -100.07 ;
      RECT 40.25 -96.96 40.6 -96.84 ;
      RECT 40.25 -93.73 40.6 -93.61 ;
      RECT 40.25 -90.5 40.6 -90.38 ;
      RECT 40.25 -87.27 40.6 -87.15 ;
      RECT 40.25 -84.04 40.6 -83.92 ;
      RECT 40.25 -80.81 40.6 -80.69 ;
      RECT 40.25 -77.58 40.6 -77.46 ;
      RECT 40.25 -74.35 40.6 -74.23 ;
      RECT 40.25 -71.12 40.6 -71 ;
      RECT 40.25 -67.89 40.6 -67.77 ;
      RECT 40.25 -64.66 40.6 -64.54 ;
      RECT 40.25 -61.43 40.6 -61.31 ;
      RECT 40.25 -58.2 40.6 -58.08 ;
      RECT 40.25 -54.97 40.6 -54.85 ;
      RECT 40.25 -51.74 40.6 -51.62 ;
      RECT 40.25 -48.51 40.6 -48.39 ;
      RECT 40.25 -45.28 40.6 -45.16 ;
      RECT 40.25 -42.05 40.6 -41.93 ;
      RECT 40.25 -38.82 40.6 -38.7 ;
      RECT 40.25 -35.59 40.6 -35.47 ;
      RECT 40.25 -32.36 40.6 -32.24 ;
      RECT 40.25 -29.13 40.6 -29.01 ;
      RECT 40.25 -25.9 40.6 -25.78 ;
      RECT 40.25 -22.67 40.6 -22.55 ;
      RECT 40.25 -19.44 40.6 -19.32 ;
      RECT 40.25 -16.21 40.6 -16.09 ;
      RECT 40.25 -12.98 40.6 -12.86 ;
      RECT 40.25 -9.75 40.6 -9.63 ;
      RECT 40.25 -6.52 40.6 -6.4 ;
      RECT 40.25 -3.29 40.6 -3.17 ;
      RECT 40.25 -0.06 40.6 0.06 ;
      RECT 40.455 -112.255 40.555 -111.775 ;
      RECT 40.455 -110.765 40.555 -110.295 ;
      RECT 40.365 -108.175 40.465 -107.215 ;
      RECT 40.365 2.175 40.465 3.135 ;
      RECT 39.765 -100.19 40.115 -100.07 ;
      RECT 39.765 -96.96 40.115 -96.84 ;
      RECT 39.765 -93.73 40.115 -93.61 ;
      RECT 39.765 -90.5 40.115 -90.38 ;
      RECT 39.765 -87.27 40.115 -87.15 ;
      RECT 39.765 -84.04 40.115 -83.92 ;
      RECT 39.765 -80.81 40.115 -80.69 ;
      RECT 39.765 -77.58 40.115 -77.46 ;
      RECT 39.765 -74.35 40.115 -74.23 ;
      RECT 39.765 -71.12 40.115 -71 ;
      RECT 39.765 -67.89 40.115 -67.77 ;
      RECT 39.765 -64.66 40.115 -64.54 ;
      RECT 39.765 -61.43 40.115 -61.31 ;
      RECT 39.765 -58.2 40.115 -58.08 ;
      RECT 39.765 -54.97 40.115 -54.85 ;
      RECT 39.765 -51.74 40.115 -51.62 ;
      RECT 39.765 -48.51 40.115 -48.39 ;
      RECT 39.765 -45.28 40.115 -45.16 ;
      RECT 39.765 -42.05 40.115 -41.93 ;
      RECT 39.765 -38.82 40.115 -38.7 ;
      RECT 39.765 -35.59 40.115 -35.47 ;
      RECT 39.765 -32.36 40.115 -32.24 ;
      RECT 39.765 -29.13 40.115 -29.01 ;
      RECT 39.765 -25.9 40.115 -25.78 ;
      RECT 39.765 -22.67 40.115 -22.55 ;
      RECT 39.765 -19.44 40.115 -19.32 ;
      RECT 39.765 -16.21 40.115 -16.09 ;
      RECT 39.765 -12.98 40.115 -12.86 ;
      RECT 39.765 -9.75 40.115 -9.63 ;
      RECT 39.765 -6.52 40.115 -6.4 ;
      RECT 39.765 -3.29 40.115 -3.17 ;
      RECT 39.765 -0.06 40.115 0.06 ;
      RECT 39.935 -108.175 40.035 -107.215 ;
      RECT 39.935 2.175 40.035 3.135 ;
      RECT 39.83 -110.765 40 -110.385 ;
      RECT 39.865 -112.245 39.965 -111.775 ;
      RECT 39.675 -108.175 39.775 -107.215 ;
      RECT 39.55 -101.06 39.65 -100.525 ;
      RECT 39.55 -99.735 39.65 -99.2 ;
      RECT 39.55 -97.83 39.65 -97.295 ;
      RECT 39.55 -96.505 39.65 -95.97 ;
      RECT 39.55 -94.6 39.65 -94.065 ;
      RECT 39.55 -93.275 39.65 -92.74 ;
      RECT 39.55 -91.37 39.65 -90.835 ;
      RECT 39.55 -90.045 39.65 -89.51 ;
      RECT 39.55 -88.14 39.65 -87.605 ;
      RECT 39.55 -86.815 39.65 -86.28 ;
      RECT 39.55 -84.91 39.65 -84.375 ;
      RECT 39.55 -83.585 39.65 -83.05 ;
      RECT 39.55 -81.68 39.65 -81.145 ;
      RECT 39.55 -80.355 39.65 -79.82 ;
      RECT 39.55 -78.45 39.65 -77.915 ;
      RECT 39.55 -77.125 39.65 -76.59 ;
      RECT 39.55 -75.22 39.65 -74.685 ;
      RECT 39.55 -73.895 39.65 -73.36 ;
      RECT 39.55 -71.99 39.65 -71.455 ;
      RECT 39.55 -70.665 39.65 -70.13 ;
      RECT 39.55 -68.76 39.65 -68.225 ;
      RECT 39.55 -67.435 39.65 -66.9 ;
      RECT 39.55 -65.53 39.65 -64.995 ;
      RECT 39.55 -64.205 39.65 -63.67 ;
      RECT 39.55 -62.3 39.65 -61.765 ;
      RECT 39.55 -60.975 39.65 -60.44 ;
      RECT 39.55 -59.07 39.65 -58.535 ;
      RECT 39.55 -57.745 39.65 -57.21 ;
      RECT 39.55 -55.84 39.65 -55.305 ;
      RECT 39.55 -54.515 39.65 -53.98 ;
      RECT 39.55 -52.61 39.65 -52.075 ;
      RECT 39.55 -51.285 39.65 -50.75 ;
      RECT 39.55 -49.38 39.65 -48.845 ;
      RECT 39.55 -48.055 39.65 -47.52 ;
      RECT 39.55 -46.15 39.65 -45.615 ;
      RECT 39.55 -44.825 39.65 -44.29 ;
      RECT 39.55 -42.92 39.65 -42.385 ;
      RECT 39.55 -41.595 39.65 -41.06 ;
      RECT 39.55 -39.69 39.65 -39.155 ;
      RECT 39.55 -38.365 39.65 -37.83 ;
      RECT 39.55 -36.46 39.65 -35.925 ;
      RECT 39.55 -35.135 39.65 -34.6 ;
      RECT 39.55 -33.23 39.65 -32.695 ;
      RECT 39.55 -31.905 39.65 -31.37 ;
      RECT 39.55 -30 39.65 -29.465 ;
      RECT 39.55 -28.675 39.65 -28.14 ;
      RECT 39.55 -26.77 39.65 -26.235 ;
      RECT 39.55 -25.445 39.65 -24.91 ;
      RECT 39.55 -23.54 39.65 -23.005 ;
      RECT 39.55 -22.215 39.65 -21.68 ;
      RECT 39.55 -20.31 39.65 -19.775 ;
      RECT 39.55 -18.985 39.65 -18.45 ;
      RECT 39.55 -17.08 39.65 -16.545 ;
      RECT 39.55 -15.755 39.65 -15.22 ;
      RECT 39.55 -13.85 39.65 -13.315 ;
      RECT 39.55 -12.525 39.65 -11.99 ;
      RECT 39.55 -10.62 39.65 -10.085 ;
      RECT 39.55 -9.295 39.65 -8.76 ;
      RECT 39.55 -7.39 39.65 -6.855 ;
      RECT 39.55 -6.065 39.65 -5.53 ;
      RECT 39.55 -4.16 39.65 -3.625 ;
      RECT 39.55 -2.835 39.65 -2.3 ;
      RECT 39.55 -0.93 39.65 -0.395 ;
      RECT 39.55 0.395 39.65 0.93 ;
      RECT 39.425 -108.175 39.525 -107.215 ;
      RECT 39.05 -100.19 39.4 -100.07 ;
      RECT 39.05 -96.96 39.4 -96.84 ;
      RECT 39.05 -93.73 39.4 -93.61 ;
      RECT 39.05 -90.5 39.4 -90.38 ;
      RECT 39.05 -87.27 39.4 -87.15 ;
      RECT 39.05 -84.04 39.4 -83.92 ;
      RECT 39.05 -80.81 39.4 -80.69 ;
      RECT 39.05 -77.58 39.4 -77.46 ;
      RECT 39.05 -74.35 39.4 -74.23 ;
      RECT 39.05 -71.12 39.4 -71 ;
      RECT 39.05 -67.89 39.4 -67.77 ;
      RECT 39.05 -64.66 39.4 -64.54 ;
      RECT 39.05 -61.43 39.4 -61.31 ;
      RECT 39.05 -58.2 39.4 -58.08 ;
      RECT 39.05 -54.97 39.4 -54.85 ;
      RECT 39.05 -51.74 39.4 -51.62 ;
      RECT 39.05 -48.51 39.4 -48.39 ;
      RECT 39.05 -45.28 39.4 -45.16 ;
      RECT 39.05 -42.05 39.4 -41.93 ;
      RECT 39.05 -38.82 39.4 -38.7 ;
      RECT 39.05 -35.59 39.4 -35.47 ;
      RECT 39.05 -32.36 39.4 -32.24 ;
      RECT 39.05 -29.13 39.4 -29.01 ;
      RECT 39.05 -25.9 39.4 -25.78 ;
      RECT 39.05 -22.67 39.4 -22.55 ;
      RECT 39.05 -19.44 39.4 -19.32 ;
      RECT 39.05 -16.21 39.4 -16.09 ;
      RECT 39.05 -12.98 39.4 -12.86 ;
      RECT 39.05 -9.75 39.4 -9.63 ;
      RECT 39.05 -6.52 39.4 -6.4 ;
      RECT 39.05 -3.29 39.4 -3.17 ;
      RECT 39.05 -0.06 39.4 0.06 ;
      RECT 39.165 -108.175 39.265 -107.215 ;
      RECT 39.165 2.175 39.265 3.135 ;
      RECT 39.065 -113.555 39.165 -113.085 ;
      RECT 38.565 -100.19 38.915 -100.07 ;
      RECT 38.565 -96.96 38.915 -96.84 ;
      RECT 38.565 -93.73 38.915 -93.61 ;
      RECT 38.565 -90.5 38.915 -90.38 ;
      RECT 38.565 -87.27 38.915 -87.15 ;
      RECT 38.565 -84.04 38.915 -83.92 ;
      RECT 38.565 -80.81 38.915 -80.69 ;
      RECT 38.565 -77.58 38.915 -77.46 ;
      RECT 38.565 -74.35 38.915 -74.23 ;
      RECT 38.565 -71.12 38.915 -71 ;
      RECT 38.565 -67.89 38.915 -67.77 ;
      RECT 38.565 -64.66 38.915 -64.54 ;
      RECT 38.565 -61.43 38.915 -61.31 ;
      RECT 38.565 -58.2 38.915 -58.08 ;
      RECT 38.565 -54.97 38.915 -54.85 ;
      RECT 38.565 -51.74 38.915 -51.62 ;
      RECT 38.565 -48.51 38.915 -48.39 ;
      RECT 38.565 -45.28 38.915 -45.16 ;
      RECT 38.565 -42.05 38.915 -41.93 ;
      RECT 38.565 -38.82 38.915 -38.7 ;
      RECT 38.565 -35.59 38.915 -35.47 ;
      RECT 38.565 -32.36 38.915 -32.24 ;
      RECT 38.565 -29.13 38.915 -29.01 ;
      RECT 38.565 -25.9 38.915 -25.78 ;
      RECT 38.565 -22.67 38.915 -22.55 ;
      RECT 38.565 -19.44 38.915 -19.32 ;
      RECT 38.565 -16.21 38.915 -16.09 ;
      RECT 38.565 -12.98 38.915 -12.86 ;
      RECT 38.565 -9.75 38.915 -9.63 ;
      RECT 38.565 -6.52 38.915 -6.4 ;
      RECT 38.565 -3.29 38.915 -3.17 ;
      RECT 38.565 -0.06 38.915 0.06 ;
      RECT 38.7 -110.735 38.85 -110.445 ;
      RECT 38.735 -108.175 38.835 -107.215 ;
      RECT 38.735 2.175 38.835 3.135 ;
      RECT 38.715 -112.19 38.815 -111.65 ;
      RECT 38.475 -113.555 38.575 -113.085 ;
      RECT 38.475 -108.175 38.575 -107.215 ;
      RECT 38.35 -101.06 38.45 -100.525 ;
      RECT 38.35 -99.735 38.45 -99.2 ;
      RECT 38.35 -97.83 38.45 -97.295 ;
      RECT 38.35 -96.505 38.45 -95.97 ;
      RECT 38.35 -94.6 38.45 -94.065 ;
      RECT 38.35 -93.275 38.45 -92.74 ;
      RECT 38.35 -91.37 38.45 -90.835 ;
      RECT 38.35 -90.045 38.45 -89.51 ;
      RECT 38.35 -88.14 38.45 -87.605 ;
      RECT 38.35 -86.815 38.45 -86.28 ;
      RECT 38.35 -84.91 38.45 -84.375 ;
      RECT 38.35 -83.585 38.45 -83.05 ;
      RECT 38.35 -81.68 38.45 -81.145 ;
      RECT 38.35 -80.355 38.45 -79.82 ;
      RECT 38.35 -78.45 38.45 -77.915 ;
      RECT 38.35 -77.125 38.45 -76.59 ;
      RECT 38.35 -75.22 38.45 -74.685 ;
      RECT 38.35 -73.895 38.45 -73.36 ;
      RECT 38.35 -71.99 38.45 -71.455 ;
      RECT 38.35 -70.665 38.45 -70.13 ;
      RECT 38.35 -68.76 38.45 -68.225 ;
      RECT 38.35 -67.435 38.45 -66.9 ;
      RECT 38.35 -65.53 38.45 -64.995 ;
      RECT 38.35 -64.205 38.45 -63.67 ;
      RECT 38.35 -62.3 38.45 -61.765 ;
      RECT 38.35 -60.975 38.45 -60.44 ;
      RECT 38.35 -59.07 38.45 -58.535 ;
      RECT 38.35 -57.745 38.45 -57.21 ;
      RECT 38.35 -55.84 38.45 -55.305 ;
      RECT 38.35 -54.515 38.45 -53.98 ;
      RECT 38.35 -52.61 38.45 -52.075 ;
      RECT 38.35 -51.285 38.45 -50.75 ;
      RECT 38.35 -49.38 38.45 -48.845 ;
      RECT 38.35 -48.055 38.45 -47.52 ;
      RECT 38.35 -46.15 38.45 -45.615 ;
      RECT 38.35 -44.825 38.45 -44.29 ;
      RECT 38.35 -42.92 38.45 -42.385 ;
      RECT 38.35 -41.595 38.45 -41.06 ;
      RECT 38.35 -39.69 38.45 -39.155 ;
      RECT 38.35 -38.365 38.45 -37.83 ;
      RECT 38.35 -36.46 38.45 -35.925 ;
      RECT 38.35 -35.135 38.45 -34.6 ;
      RECT 38.35 -33.23 38.45 -32.695 ;
      RECT 38.35 -31.905 38.45 -31.37 ;
      RECT 38.35 -30 38.45 -29.465 ;
      RECT 38.35 -28.675 38.45 -28.14 ;
      RECT 38.35 -26.77 38.45 -26.235 ;
      RECT 38.35 -25.445 38.45 -24.91 ;
      RECT 38.35 -23.54 38.45 -23.005 ;
      RECT 38.35 -22.215 38.45 -21.68 ;
      RECT 38.35 -20.31 38.45 -19.775 ;
      RECT 38.35 -18.985 38.45 -18.45 ;
      RECT 38.35 -17.08 38.45 -16.545 ;
      RECT 38.35 -15.755 38.45 -15.22 ;
      RECT 38.35 -13.85 38.45 -13.315 ;
      RECT 38.35 -12.525 38.45 -11.99 ;
      RECT 38.35 -10.62 38.45 -10.085 ;
      RECT 38.35 -9.295 38.45 -8.76 ;
      RECT 38.35 -7.39 38.45 -6.855 ;
      RECT 38.35 -6.065 38.45 -5.53 ;
      RECT 38.35 -4.16 38.45 -3.625 ;
      RECT 38.35 -2.835 38.45 -2.3 ;
      RECT 38.35 -0.93 38.45 -0.395 ;
      RECT 38.35 0.395 38.45 0.93 ;
      RECT 38.225 -104.945 38.325 -103.985 ;
      RECT 37.85 -100.19 38.2 -100.07 ;
      RECT 37.85 -96.96 38.2 -96.84 ;
      RECT 37.85 -93.73 38.2 -93.61 ;
      RECT 37.85 -90.5 38.2 -90.38 ;
      RECT 37.85 -87.27 38.2 -87.15 ;
      RECT 37.85 -84.04 38.2 -83.92 ;
      RECT 37.85 -80.81 38.2 -80.69 ;
      RECT 37.85 -77.58 38.2 -77.46 ;
      RECT 37.85 -74.35 38.2 -74.23 ;
      RECT 37.85 -71.12 38.2 -71 ;
      RECT 37.85 -67.89 38.2 -67.77 ;
      RECT 37.85 -64.66 38.2 -64.54 ;
      RECT 37.85 -61.43 38.2 -61.31 ;
      RECT 37.85 -58.2 38.2 -58.08 ;
      RECT 37.85 -54.97 38.2 -54.85 ;
      RECT 37.85 -51.74 38.2 -51.62 ;
      RECT 37.85 -48.51 38.2 -48.39 ;
      RECT 37.85 -45.28 38.2 -45.16 ;
      RECT 37.85 -42.05 38.2 -41.93 ;
      RECT 37.85 -38.82 38.2 -38.7 ;
      RECT 37.85 -35.59 38.2 -35.47 ;
      RECT 37.85 -32.36 38.2 -32.24 ;
      RECT 37.85 -29.13 38.2 -29.01 ;
      RECT 37.85 -25.9 38.2 -25.78 ;
      RECT 37.85 -22.67 38.2 -22.55 ;
      RECT 37.85 -19.44 38.2 -19.32 ;
      RECT 37.85 -16.21 38.2 -16.09 ;
      RECT 37.85 -12.98 38.2 -12.86 ;
      RECT 37.85 -9.75 38.2 -9.63 ;
      RECT 37.85 -6.52 38.2 -6.4 ;
      RECT 37.85 -3.29 38.2 -3.17 ;
      RECT 37.85 -0.06 38.2 0.06 ;
      RECT 37.965 -104.945 38.065 -103.985 ;
      RECT 37.965 2.175 38.065 3.135 ;
      RECT 37.675 -112.255 37.775 -111.775 ;
      RECT 37.675 -110.765 37.775 -110.295 ;
      RECT 37.365 -100.19 37.715 -100.07 ;
      RECT 37.365 -96.96 37.715 -96.84 ;
      RECT 37.365 -93.73 37.715 -93.61 ;
      RECT 37.365 -90.5 37.715 -90.38 ;
      RECT 37.365 -87.27 37.715 -87.15 ;
      RECT 37.365 -84.04 37.715 -83.92 ;
      RECT 37.365 -80.81 37.715 -80.69 ;
      RECT 37.365 -77.58 37.715 -77.46 ;
      RECT 37.365 -74.35 37.715 -74.23 ;
      RECT 37.365 -71.12 37.715 -71 ;
      RECT 37.365 -67.89 37.715 -67.77 ;
      RECT 37.365 -64.66 37.715 -64.54 ;
      RECT 37.365 -61.43 37.715 -61.31 ;
      RECT 37.365 -58.2 37.715 -58.08 ;
      RECT 37.365 -54.97 37.715 -54.85 ;
      RECT 37.365 -51.74 37.715 -51.62 ;
      RECT 37.365 -48.51 37.715 -48.39 ;
      RECT 37.365 -45.28 37.715 -45.16 ;
      RECT 37.365 -42.05 37.715 -41.93 ;
      RECT 37.365 -38.82 37.715 -38.7 ;
      RECT 37.365 -35.59 37.715 -35.47 ;
      RECT 37.365 -32.36 37.715 -32.24 ;
      RECT 37.365 -29.13 37.715 -29.01 ;
      RECT 37.365 -25.9 37.715 -25.78 ;
      RECT 37.365 -22.67 37.715 -22.55 ;
      RECT 37.365 -19.44 37.715 -19.32 ;
      RECT 37.365 -16.21 37.715 -16.09 ;
      RECT 37.365 -12.98 37.715 -12.86 ;
      RECT 37.365 -9.75 37.715 -9.63 ;
      RECT 37.365 -6.52 37.715 -6.4 ;
      RECT 37.365 -3.29 37.715 -3.17 ;
      RECT 37.365 -0.06 37.715 0.06 ;
      RECT 37.535 -104.945 37.635 -103.985 ;
      RECT 37.535 2.175 37.635 3.135 ;
      RECT 33.635 -108.655 37.415 -108.535 ;
      RECT 37.275 -104.945 37.375 -103.985 ;
      RECT 37.15 -101.06 37.25 -100.525 ;
      RECT 37.15 -99.735 37.25 -99.2 ;
      RECT 37.15 -97.83 37.25 -97.295 ;
      RECT 37.15 -96.505 37.25 -95.97 ;
      RECT 37.15 -94.6 37.25 -94.065 ;
      RECT 37.15 -93.275 37.25 -92.74 ;
      RECT 37.15 -91.37 37.25 -90.835 ;
      RECT 37.15 -90.045 37.25 -89.51 ;
      RECT 37.15 -88.14 37.25 -87.605 ;
      RECT 37.15 -86.815 37.25 -86.28 ;
      RECT 37.15 -84.91 37.25 -84.375 ;
      RECT 37.15 -83.585 37.25 -83.05 ;
      RECT 37.15 -81.68 37.25 -81.145 ;
      RECT 37.15 -80.355 37.25 -79.82 ;
      RECT 37.15 -78.45 37.25 -77.915 ;
      RECT 37.15 -77.125 37.25 -76.59 ;
      RECT 37.15 -75.22 37.25 -74.685 ;
      RECT 37.15 -73.895 37.25 -73.36 ;
      RECT 37.15 -71.99 37.25 -71.455 ;
      RECT 37.15 -70.665 37.25 -70.13 ;
      RECT 37.15 -68.76 37.25 -68.225 ;
      RECT 37.15 -67.435 37.25 -66.9 ;
      RECT 37.15 -65.53 37.25 -64.995 ;
      RECT 37.15 -64.205 37.25 -63.67 ;
      RECT 37.15 -62.3 37.25 -61.765 ;
      RECT 37.15 -60.975 37.25 -60.44 ;
      RECT 37.15 -59.07 37.25 -58.535 ;
      RECT 37.15 -57.745 37.25 -57.21 ;
      RECT 37.15 -55.84 37.25 -55.305 ;
      RECT 37.15 -54.515 37.25 -53.98 ;
      RECT 37.15 -52.61 37.25 -52.075 ;
      RECT 37.15 -51.285 37.25 -50.75 ;
      RECT 37.15 -49.38 37.25 -48.845 ;
      RECT 37.15 -48.055 37.25 -47.52 ;
      RECT 37.15 -46.15 37.25 -45.615 ;
      RECT 37.15 -44.825 37.25 -44.29 ;
      RECT 37.15 -42.92 37.25 -42.385 ;
      RECT 37.15 -41.595 37.25 -41.06 ;
      RECT 37.15 -39.69 37.25 -39.155 ;
      RECT 37.15 -38.365 37.25 -37.83 ;
      RECT 37.15 -36.46 37.25 -35.925 ;
      RECT 37.15 -35.135 37.25 -34.6 ;
      RECT 37.15 -33.23 37.25 -32.695 ;
      RECT 37.15 -31.905 37.25 -31.37 ;
      RECT 37.15 -30 37.25 -29.465 ;
      RECT 37.15 -28.675 37.25 -28.14 ;
      RECT 37.15 -26.77 37.25 -26.235 ;
      RECT 37.15 -25.445 37.25 -24.91 ;
      RECT 37.15 -23.54 37.25 -23.005 ;
      RECT 37.15 -22.215 37.25 -21.68 ;
      RECT 37.15 -20.31 37.25 -19.775 ;
      RECT 37.15 -18.985 37.25 -18.45 ;
      RECT 37.15 -17.08 37.25 -16.545 ;
      RECT 37.15 -15.755 37.25 -15.22 ;
      RECT 37.15 -13.85 37.25 -13.315 ;
      RECT 37.15 -12.525 37.25 -11.99 ;
      RECT 37.15 -10.62 37.25 -10.085 ;
      RECT 37.15 -9.295 37.25 -8.76 ;
      RECT 37.15 -7.39 37.25 -6.855 ;
      RECT 37.15 -6.065 37.25 -5.53 ;
      RECT 37.15 -4.16 37.25 -3.625 ;
      RECT 37.15 -2.835 37.25 -2.3 ;
      RECT 37.15 -0.93 37.25 -0.395 ;
      RECT 37.15 0.395 37.25 0.93 ;
      RECT 37.085 -110.75 37.205 -110.37 ;
      RECT 37.085 -112.245 37.185 -111.775 ;
      RECT 37.025 -104.945 37.125 -103.985 ;
      RECT 36.65 -100.19 37 -100.07 ;
      RECT 36.65 -96.96 37 -96.84 ;
      RECT 36.65 -93.73 37 -93.61 ;
      RECT 36.65 -90.5 37 -90.38 ;
      RECT 36.65 -87.27 37 -87.15 ;
      RECT 36.65 -84.04 37 -83.92 ;
      RECT 36.65 -80.81 37 -80.69 ;
      RECT 36.65 -77.58 37 -77.46 ;
      RECT 36.65 -74.35 37 -74.23 ;
      RECT 36.65 -71.12 37 -71 ;
      RECT 36.65 -67.89 37 -67.77 ;
      RECT 36.65 -64.66 37 -64.54 ;
      RECT 36.65 -61.43 37 -61.31 ;
      RECT 36.65 -58.2 37 -58.08 ;
      RECT 36.65 -54.97 37 -54.85 ;
      RECT 36.65 -51.74 37 -51.62 ;
      RECT 36.65 -48.51 37 -48.39 ;
      RECT 36.65 -45.28 37 -45.16 ;
      RECT 36.65 -42.05 37 -41.93 ;
      RECT 36.65 -38.82 37 -38.7 ;
      RECT 36.65 -35.59 37 -35.47 ;
      RECT 36.65 -32.36 37 -32.24 ;
      RECT 36.65 -29.13 37 -29.01 ;
      RECT 36.65 -25.9 37 -25.78 ;
      RECT 36.65 -22.67 37 -22.55 ;
      RECT 36.65 -19.44 37 -19.32 ;
      RECT 36.65 -16.21 37 -16.09 ;
      RECT 36.65 -12.98 37 -12.86 ;
      RECT 36.65 -9.75 37 -9.63 ;
      RECT 36.65 -6.52 37 -6.4 ;
      RECT 36.65 -3.29 37 -3.17 ;
      RECT 36.65 -0.06 37 0.06 ;
      RECT 36.765 -104.945 36.865 -103.985 ;
      RECT 36.765 2.175 36.865 3.135 ;
      RECT 36.495 -109.595 36.63 -109.275 ;
      RECT 36.165 -100.19 36.515 -100.07 ;
      RECT 36.165 -96.96 36.515 -96.84 ;
      RECT 36.165 -93.73 36.515 -93.61 ;
      RECT 36.165 -90.5 36.515 -90.38 ;
      RECT 36.165 -87.27 36.515 -87.15 ;
      RECT 36.165 -84.04 36.515 -83.92 ;
      RECT 36.165 -80.81 36.515 -80.69 ;
      RECT 36.165 -77.58 36.515 -77.46 ;
      RECT 36.165 -74.35 36.515 -74.23 ;
      RECT 36.165 -71.12 36.515 -71 ;
      RECT 36.165 -67.89 36.515 -67.77 ;
      RECT 36.165 -64.66 36.515 -64.54 ;
      RECT 36.165 -61.43 36.515 -61.31 ;
      RECT 36.165 -58.2 36.515 -58.08 ;
      RECT 36.165 -54.97 36.515 -54.85 ;
      RECT 36.165 -51.74 36.515 -51.62 ;
      RECT 36.165 -48.51 36.515 -48.39 ;
      RECT 36.165 -45.28 36.515 -45.16 ;
      RECT 36.165 -42.05 36.515 -41.93 ;
      RECT 36.165 -38.82 36.515 -38.7 ;
      RECT 36.165 -35.59 36.515 -35.47 ;
      RECT 36.165 -32.36 36.515 -32.24 ;
      RECT 36.165 -29.13 36.515 -29.01 ;
      RECT 36.165 -25.9 36.515 -25.78 ;
      RECT 36.165 -22.67 36.515 -22.55 ;
      RECT 36.165 -19.44 36.515 -19.32 ;
      RECT 36.165 -16.21 36.515 -16.09 ;
      RECT 36.165 -12.98 36.515 -12.86 ;
      RECT 36.165 -9.75 36.515 -9.63 ;
      RECT 36.165 -6.52 36.515 -6.4 ;
      RECT 36.165 -3.29 36.515 -3.17 ;
      RECT 36.165 -0.06 36.515 0.06 ;
      RECT 36.335 -104.945 36.435 -103.985 ;
      RECT 36.335 2.175 36.435 3.135 ;
      RECT 36.16 -109.595 36.305 -109.275 ;
      RECT 36.075 -104.945 36.175 -103.985 ;
      RECT 35.95 -101.06 36.05 -100.525 ;
      RECT 35.95 -99.735 36.05 -99.2 ;
      RECT 35.95 -97.83 36.05 -97.295 ;
      RECT 35.95 -96.505 36.05 -95.97 ;
      RECT 35.95 -94.6 36.05 -94.065 ;
      RECT 35.95 -93.275 36.05 -92.74 ;
      RECT 35.95 -91.37 36.05 -90.835 ;
      RECT 35.95 -90.045 36.05 -89.51 ;
      RECT 35.95 -88.14 36.05 -87.605 ;
      RECT 35.95 -86.815 36.05 -86.28 ;
      RECT 35.95 -84.91 36.05 -84.375 ;
      RECT 35.95 -83.585 36.05 -83.05 ;
      RECT 35.95 -81.68 36.05 -81.145 ;
      RECT 35.95 -80.355 36.05 -79.82 ;
      RECT 35.95 -78.45 36.05 -77.915 ;
      RECT 35.95 -77.125 36.05 -76.59 ;
      RECT 35.95 -75.22 36.05 -74.685 ;
      RECT 35.95 -73.895 36.05 -73.36 ;
      RECT 35.95 -71.99 36.05 -71.455 ;
      RECT 35.95 -70.665 36.05 -70.13 ;
      RECT 35.95 -68.76 36.05 -68.225 ;
      RECT 35.95 -67.435 36.05 -66.9 ;
      RECT 35.95 -65.53 36.05 -64.995 ;
      RECT 35.95 -64.205 36.05 -63.67 ;
      RECT 35.95 -62.3 36.05 -61.765 ;
      RECT 35.95 -60.975 36.05 -60.44 ;
      RECT 35.95 -59.07 36.05 -58.535 ;
      RECT 35.95 -57.745 36.05 -57.21 ;
      RECT 35.95 -55.84 36.05 -55.305 ;
      RECT 35.95 -54.515 36.05 -53.98 ;
      RECT 35.95 -52.61 36.05 -52.075 ;
      RECT 35.95 -51.285 36.05 -50.75 ;
      RECT 35.95 -49.38 36.05 -48.845 ;
      RECT 35.95 -48.055 36.05 -47.52 ;
      RECT 35.95 -46.15 36.05 -45.615 ;
      RECT 35.95 -44.825 36.05 -44.29 ;
      RECT 35.95 -42.92 36.05 -42.385 ;
      RECT 35.95 -41.595 36.05 -41.06 ;
      RECT 35.95 -39.69 36.05 -39.155 ;
      RECT 35.95 -38.365 36.05 -37.83 ;
      RECT 35.95 -36.46 36.05 -35.925 ;
      RECT 35.95 -35.135 36.05 -34.6 ;
      RECT 35.95 -33.23 36.05 -32.695 ;
      RECT 35.95 -31.905 36.05 -31.37 ;
      RECT 35.95 -30 36.05 -29.465 ;
      RECT 35.95 -28.675 36.05 -28.14 ;
      RECT 35.95 -26.77 36.05 -26.235 ;
      RECT 35.95 -25.445 36.05 -24.91 ;
      RECT 35.95 -23.54 36.05 -23.005 ;
      RECT 35.95 -22.215 36.05 -21.68 ;
      RECT 35.95 -20.31 36.05 -19.775 ;
      RECT 35.95 -18.985 36.05 -18.45 ;
      RECT 35.95 -17.08 36.05 -16.545 ;
      RECT 35.95 -15.755 36.05 -15.22 ;
      RECT 35.95 -13.85 36.05 -13.315 ;
      RECT 35.95 -12.525 36.05 -11.99 ;
      RECT 35.95 -10.62 36.05 -10.085 ;
      RECT 35.95 -9.295 36.05 -8.76 ;
      RECT 35.95 -7.39 36.05 -6.855 ;
      RECT 35.95 -6.065 36.05 -5.53 ;
      RECT 35.95 -4.16 36.05 -3.625 ;
      RECT 35.95 -2.835 36.05 -2.3 ;
      RECT 35.95 -0.93 36.05 -0.395 ;
      RECT 35.95 0.395 36.05 0.93 ;
      RECT 35.825 -108.175 35.925 -107.215 ;
      RECT 35.45 -100.19 35.8 -100.07 ;
      RECT 35.45 -96.96 35.8 -96.84 ;
      RECT 35.45 -93.73 35.8 -93.61 ;
      RECT 35.45 -90.5 35.8 -90.38 ;
      RECT 35.45 -87.27 35.8 -87.15 ;
      RECT 35.45 -84.04 35.8 -83.92 ;
      RECT 35.45 -80.81 35.8 -80.69 ;
      RECT 35.45 -77.58 35.8 -77.46 ;
      RECT 35.45 -74.35 35.8 -74.23 ;
      RECT 35.45 -71.12 35.8 -71 ;
      RECT 35.45 -67.89 35.8 -67.77 ;
      RECT 35.45 -64.66 35.8 -64.54 ;
      RECT 35.45 -61.43 35.8 -61.31 ;
      RECT 35.45 -58.2 35.8 -58.08 ;
      RECT 35.45 -54.97 35.8 -54.85 ;
      RECT 35.45 -51.74 35.8 -51.62 ;
      RECT 35.45 -48.51 35.8 -48.39 ;
      RECT 35.45 -45.28 35.8 -45.16 ;
      RECT 35.45 -42.05 35.8 -41.93 ;
      RECT 35.45 -38.82 35.8 -38.7 ;
      RECT 35.45 -35.59 35.8 -35.47 ;
      RECT 35.45 -32.36 35.8 -32.24 ;
      RECT 35.45 -29.13 35.8 -29.01 ;
      RECT 35.45 -25.9 35.8 -25.78 ;
      RECT 35.45 -22.67 35.8 -22.55 ;
      RECT 35.45 -19.44 35.8 -19.32 ;
      RECT 35.45 -16.21 35.8 -16.09 ;
      RECT 35.45 -12.98 35.8 -12.86 ;
      RECT 35.45 -9.75 35.8 -9.63 ;
      RECT 35.45 -6.52 35.8 -6.4 ;
      RECT 35.45 -3.29 35.8 -3.17 ;
      RECT 35.45 -0.06 35.8 0.06 ;
      RECT 35.655 -112.255 35.755 -111.775 ;
      RECT 35.655 -110.765 35.755 -110.295 ;
      RECT 35.565 -108.175 35.665 -107.215 ;
      RECT 35.565 2.175 35.665 3.135 ;
      RECT 34.965 -100.19 35.315 -100.07 ;
      RECT 34.965 -96.96 35.315 -96.84 ;
      RECT 34.965 -93.73 35.315 -93.61 ;
      RECT 34.965 -90.5 35.315 -90.38 ;
      RECT 34.965 -87.27 35.315 -87.15 ;
      RECT 34.965 -84.04 35.315 -83.92 ;
      RECT 34.965 -80.81 35.315 -80.69 ;
      RECT 34.965 -77.58 35.315 -77.46 ;
      RECT 34.965 -74.35 35.315 -74.23 ;
      RECT 34.965 -71.12 35.315 -71 ;
      RECT 34.965 -67.89 35.315 -67.77 ;
      RECT 34.965 -64.66 35.315 -64.54 ;
      RECT 34.965 -61.43 35.315 -61.31 ;
      RECT 34.965 -58.2 35.315 -58.08 ;
      RECT 34.965 -54.97 35.315 -54.85 ;
      RECT 34.965 -51.74 35.315 -51.62 ;
      RECT 34.965 -48.51 35.315 -48.39 ;
      RECT 34.965 -45.28 35.315 -45.16 ;
      RECT 34.965 -42.05 35.315 -41.93 ;
      RECT 34.965 -38.82 35.315 -38.7 ;
      RECT 34.965 -35.59 35.315 -35.47 ;
      RECT 34.965 -32.36 35.315 -32.24 ;
      RECT 34.965 -29.13 35.315 -29.01 ;
      RECT 34.965 -25.9 35.315 -25.78 ;
      RECT 34.965 -22.67 35.315 -22.55 ;
      RECT 34.965 -19.44 35.315 -19.32 ;
      RECT 34.965 -16.21 35.315 -16.09 ;
      RECT 34.965 -12.98 35.315 -12.86 ;
      RECT 34.965 -9.75 35.315 -9.63 ;
      RECT 34.965 -6.52 35.315 -6.4 ;
      RECT 34.965 -3.29 35.315 -3.17 ;
      RECT 34.965 -0.06 35.315 0.06 ;
      RECT 35.135 -108.175 35.235 -107.215 ;
      RECT 35.135 2.175 35.235 3.135 ;
      RECT 35.03 -110.765 35.2 -110.385 ;
      RECT 35.065 -112.245 35.165 -111.775 ;
      RECT 34.875 -108.175 34.975 -107.215 ;
      RECT 34.75 -101.06 34.85 -100.525 ;
      RECT 34.75 -99.735 34.85 -99.2 ;
      RECT 34.75 -97.83 34.85 -97.295 ;
      RECT 34.75 -96.505 34.85 -95.97 ;
      RECT 34.75 -94.6 34.85 -94.065 ;
      RECT 34.75 -93.275 34.85 -92.74 ;
      RECT 34.75 -91.37 34.85 -90.835 ;
      RECT 34.75 -90.045 34.85 -89.51 ;
      RECT 34.75 -88.14 34.85 -87.605 ;
      RECT 34.75 -86.815 34.85 -86.28 ;
      RECT 34.75 -84.91 34.85 -84.375 ;
      RECT 34.75 -83.585 34.85 -83.05 ;
      RECT 34.75 -81.68 34.85 -81.145 ;
      RECT 34.75 -80.355 34.85 -79.82 ;
      RECT 34.75 -78.45 34.85 -77.915 ;
      RECT 34.75 -77.125 34.85 -76.59 ;
      RECT 34.75 -75.22 34.85 -74.685 ;
      RECT 34.75 -73.895 34.85 -73.36 ;
      RECT 34.75 -71.99 34.85 -71.455 ;
      RECT 34.75 -70.665 34.85 -70.13 ;
      RECT 34.75 -68.76 34.85 -68.225 ;
      RECT 34.75 -67.435 34.85 -66.9 ;
      RECT 34.75 -65.53 34.85 -64.995 ;
      RECT 34.75 -64.205 34.85 -63.67 ;
      RECT 34.75 -62.3 34.85 -61.765 ;
      RECT 34.75 -60.975 34.85 -60.44 ;
      RECT 34.75 -59.07 34.85 -58.535 ;
      RECT 34.75 -57.745 34.85 -57.21 ;
      RECT 34.75 -55.84 34.85 -55.305 ;
      RECT 34.75 -54.515 34.85 -53.98 ;
      RECT 34.75 -52.61 34.85 -52.075 ;
      RECT 34.75 -51.285 34.85 -50.75 ;
      RECT 34.75 -49.38 34.85 -48.845 ;
      RECT 34.75 -48.055 34.85 -47.52 ;
      RECT 34.75 -46.15 34.85 -45.615 ;
      RECT 34.75 -44.825 34.85 -44.29 ;
      RECT 34.75 -42.92 34.85 -42.385 ;
      RECT 34.75 -41.595 34.85 -41.06 ;
      RECT 34.75 -39.69 34.85 -39.155 ;
      RECT 34.75 -38.365 34.85 -37.83 ;
      RECT 34.75 -36.46 34.85 -35.925 ;
      RECT 34.75 -35.135 34.85 -34.6 ;
      RECT 34.75 -33.23 34.85 -32.695 ;
      RECT 34.75 -31.905 34.85 -31.37 ;
      RECT 34.75 -30 34.85 -29.465 ;
      RECT 34.75 -28.675 34.85 -28.14 ;
      RECT 34.75 -26.77 34.85 -26.235 ;
      RECT 34.75 -25.445 34.85 -24.91 ;
      RECT 34.75 -23.54 34.85 -23.005 ;
      RECT 34.75 -22.215 34.85 -21.68 ;
      RECT 34.75 -20.31 34.85 -19.775 ;
      RECT 34.75 -18.985 34.85 -18.45 ;
      RECT 34.75 -17.08 34.85 -16.545 ;
      RECT 34.75 -15.755 34.85 -15.22 ;
      RECT 34.75 -13.85 34.85 -13.315 ;
      RECT 34.75 -12.525 34.85 -11.99 ;
      RECT 34.75 -10.62 34.85 -10.085 ;
      RECT 34.75 -9.295 34.85 -8.76 ;
      RECT 34.75 -7.39 34.85 -6.855 ;
      RECT 34.75 -6.065 34.85 -5.53 ;
      RECT 34.75 -4.16 34.85 -3.625 ;
      RECT 34.75 -2.835 34.85 -2.3 ;
      RECT 34.75 -0.93 34.85 -0.395 ;
      RECT 34.75 0.395 34.85 0.93 ;
      RECT 34.625 -108.175 34.725 -107.215 ;
      RECT 34.25 -100.19 34.6 -100.07 ;
      RECT 34.25 -96.96 34.6 -96.84 ;
      RECT 34.25 -93.73 34.6 -93.61 ;
      RECT 34.25 -90.5 34.6 -90.38 ;
      RECT 34.25 -87.27 34.6 -87.15 ;
      RECT 34.25 -84.04 34.6 -83.92 ;
      RECT 34.25 -80.81 34.6 -80.69 ;
      RECT 34.25 -77.58 34.6 -77.46 ;
      RECT 34.25 -74.35 34.6 -74.23 ;
      RECT 34.25 -71.12 34.6 -71 ;
      RECT 34.25 -67.89 34.6 -67.77 ;
      RECT 34.25 -64.66 34.6 -64.54 ;
      RECT 34.25 -61.43 34.6 -61.31 ;
      RECT 34.25 -58.2 34.6 -58.08 ;
      RECT 34.25 -54.97 34.6 -54.85 ;
      RECT 34.25 -51.74 34.6 -51.62 ;
      RECT 34.25 -48.51 34.6 -48.39 ;
      RECT 34.25 -45.28 34.6 -45.16 ;
      RECT 34.25 -42.05 34.6 -41.93 ;
      RECT 34.25 -38.82 34.6 -38.7 ;
      RECT 34.25 -35.59 34.6 -35.47 ;
      RECT 34.25 -32.36 34.6 -32.24 ;
      RECT 34.25 -29.13 34.6 -29.01 ;
      RECT 34.25 -25.9 34.6 -25.78 ;
      RECT 34.25 -22.67 34.6 -22.55 ;
      RECT 34.25 -19.44 34.6 -19.32 ;
      RECT 34.25 -16.21 34.6 -16.09 ;
      RECT 34.25 -12.98 34.6 -12.86 ;
      RECT 34.25 -9.75 34.6 -9.63 ;
      RECT 34.25 -6.52 34.6 -6.4 ;
      RECT 34.25 -3.29 34.6 -3.17 ;
      RECT 34.25 -0.06 34.6 0.06 ;
      RECT 34.365 -108.175 34.465 -107.215 ;
      RECT 34.365 2.175 34.465 3.135 ;
      RECT 34.265 -113.555 34.365 -113.085 ;
      RECT 33.765 -100.19 34.115 -100.07 ;
      RECT 33.765 -96.96 34.115 -96.84 ;
      RECT 33.765 -93.73 34.115 -93.61 ;
      RECT 33.765 -90.5 34.115 -90.38 ;
      RECT 33.765 -87.27 34.115 -87.15 ;
      RECT 33.765 -84.04 34.115 -83.92 ;
      RECT 33.765 -80.81 34.115 -80.69 ;
      RECT 33.765 -77.58 34.115 -77.46 ;
      RECT 33.765 -74.35 34.115 -74.23 ;
      RECT 33.765 -71.12 34.115 -71 ;
      RECT 33.765 -67.89 34.115 -67.77 ;
      RECT 33.765 -64.66 34.115 -64.54 ;
      RECT 33.765 -61.43 34.115 -61.31 ;
      RECT 33.765 -58.2 34.115 -58.08 ;
      RECT 33.765 -54.97 34.115 -54.85 ;
      RECT 33.765 -51.74 34.115 -51.62 ;
      RECT 33.765 -48.51 34.115 -48.39 ;
      RECT 33.765 -45.28 34.115 -45.16 ;
      RECT 33.765 -42.05 34.115 -41.93 ;
      RECT 33.765 -38.82 34.115 -38.7 ;
      RECT 33.765 -35.59 34.115 -35.47 ;
      RECT 33.765 -32.36 34.115 -32.24 ;
      RECT 33.765 -29.13 34.115 -29.01 ;
      RECT 33.765 -25.9 34.115 -25.78 ;
      RECT 33.765 -22.67 34.115 -22.55 ;
      RECT 33.765 -19.44 34.115 -19.32 ;
      RECT 33.765 -16.21 34.115 -16.09 ;
      RECT 33.765 -12.98 34.115 -12.86 ;
      RECT 33.765 -9.75 34.115 -9.63 ;
      RECT 33.765 -6.52 34.115 -6.4 ;
      RECT 33.765 -3.29 34.115 -3.17 ;
      RECT 33.765 -0.06 34.115 0.06 ;
      RECT 33.9 -110.735 34.05 -110.445 ;
      RECT 33.935 -108.175 34.035 -107.215 ;
      RECT 33.935 2.175 34.035 3.135 ;
      RECT 33.915 -112.19 34.015 -111.65 ;
      RECT 33.675 -113.555 33.775 -113.085 ;
      RECT 33.675 -108.175 33.775 -107.215 ;
      RECT 33.55 -101.06 33.65 -100.525 ;
      RECT 33.55 -99.735 33.65 -99.2 ;
      RECT 33.55 -97.83 33.65 -97.295 ;
      RECT 33.55 -96.505 33.65 -95.97 ;
      RECT 33.55 -94.6 33.65 -94.065 ;
      RECT 33.55 -93.275 33.65 -92.74 ;
      RECT 33.55 -91.37 33.65 -90.835 ;
      RECT 33.55 -90.045 33.65 -89.51 ;
      RECT 33.55 -88.14 33.65 -87.605 ;
      RECT 33.55 -86.815 33.65 -86.28 ;
      RECT 33.55 -84.91 33.65 -84.375 ;
      RECT 33.55 -83.585 33.65 -83.05 ;
      RECT 33.55 -81.68 33.65 -81.145 ;
      RECT 33.55 -80.355 33.65 -79.82 ;
      RECT 33.55 -78.45 33.65 -77.915 ;
      RECT 33.55 -77.125 33.65 -76.59 ;
      RECT 33.55 -75.22 33.65 -74.685 ;
      RECT 33.55 -73.895 33.65 -73.36 ;
      RECT 33.55 -71.99 33.65 -71.455 ;
      RECT 33.55 -70.665 33.65 -70.13 ;
      RECT 33.55 -68.76 33.65 -68.225 ;
      RECT 33.55 -67.435 33.65 -66.9 ;
      RECT 33.55 -65.53 33.65 -64.995 ;
      RECT 33.55 -64.205 33.65 -63.67 ;
      RECT 33.55 -62.3 33.65 -61.765 ;
      RECT 33.55 -60.975 33.65 -60.44 ;
      RECT 33.55 -59.07 33.65 -58.535 ;
      RECT 33.55 -57.745 33.65 -57.21 ;
      RECT 33.55 -55.84 33.65 -55.305 ;
      RECT 33.55 -54.515 33.65 -53.98 ;
      RECT 33.55 -52.61 33.65 -52.075 ;
      RECT 33.55 -51.285 33.65 -50.75 ;
      RECT 33.55 -49.38 33.65 -48.845 ;
      RECT 33.55 -48.055 33.65 -47.52 ;
      RECT 33.55 -46.15 33.65 -45.615 ;
      RECT 33.55 -44.825 33.65 -44.29 ;
      RECT 33.55 -42.92 33.65 -42.385 ;
      RECT 33.55 -41.595 33.65 -41.06 ;
      RECT 33.55 -39.69 33.65 -39.155 ;
      RECT 33.55 -38.365 33.65 -37.83 ;
      RECT 33.55 -36.46 33.65 -35.925 ;
      RECT 33.55 -35.135 33.65 -34.6 ;
      RECT 33.55 -33.23 33.65 -32.695 ;
      RECT 33.55 -31.905 33.65 -31.37 ;
      RECT 33.55 -30 33.65 -29.465 ;
      RECT 33.55 -28.675 33.65 -28.14 ;
      RECT 33.55 -26.77 33.65 -26.235 ;
      RECT 33.55 -25.445 33.65 -24.91 ;
      RECT 33.55 -23.54 33.65 -23.005 ;
      RECT 33.55 -22.215 33.65 -21.68 ;
      RECT 33.55 -20.31 33.65 -19.775 ;
      RECT 33.55 -18.985 33.65 -18.45 ;
      RECT 33.55 -17.08 33.65 -16.545 ;
      RECT 33.55 -15.755 33.65 -15.22 ;
      RECT 33.55 -13.85 33.65 -13.315 ;
      RECT 33.55 -12.525 33.65 -11.99 ;
      RECT 33.55 -10.62 33.65 -10.085 ;
      RECT 33.55 -9.295 33.65 -8.76 ;
      RECT 33.55 -7.39 33.65 -6.855 ;
      RECT 33.55 -6.065 33.65 -5.53 ;
      RECT 33.55 -4.16 33.65 -3.625 ;
      RECT 33.55 -2.835 33.65 -2.3 ;
      RECT 33.55 -0.93 33.65 -0.395 ;
      RECT 33.55 0.395 33.65 0.93 ;
      RECT 33.425 -104.945 33.525 -103.985 ;
      RECT 33.05 -100.19 33.4 -100.07 ;
      RECT 33.05 -96.96 33.4 -96.84 ;
      RECT 33.05 -93.73 33.4 -93.61 ;
      RECT 33.05 -90.5 33.4 -90.38 ;
      RECT 33.05 -87.27 33.4 -87.15 ;
      RECT 33.05 -84.04 33.4 -83.92 ;
      RECT 33.05 -80.81 33.4 -80.69 ;
      RECT 33.05 -77.58 33.4 -77.46 ;
      RECT 33.05 -74.35 33.4 -74.23 ;
      RECT 33.05 -71.12 33.4 -71 ;
      RECT 33.05 -67.89 33.4 -67.77 ;
      RECT 33.05 -64.66 33.4 -64.54 ;
      RECT 33.05 -61.43 33.4 -61.31 ;
      RECT 33.05 -58.2 33.4 -58.08 ;
      RECT 33.05 -54.97 33.4 -54.85 ;
      RECT 33.05 -51.74 33.4 -51.62 ;
      RECT 33.05 -48.51 33.4 -48.39 ;
      RECT 33.05 -45.28 33.4 -45.16 ;
      RECT 33.05 -42.05 33.4 -41.93 ;
      RECT 33.05 -38.82 33.4 -38.7 ;
      RECT 33.05 -35.59 33.4 -35.47 ;
      RECT 33.05 -32.36 33.4 -32.24 ;
      RECT 33.05 -29.13 33.4 -29.01 ;
      RECT 33.05 -25.9 33.4 -25.78 ;
      RECT 33.05 -22.67 33.4 -22.55 ;
      RECT 33.05 -19.44 33.4 -19.32 ;
      RECT 33.05 -16.21 33.4 -16.09 ;
      RECT 33.05 -12.98 33.4 -12.86 ;
      RECT 33.05 -9.75 33.4 -9.63 ;
      RECT 33.05 -6.52 33.4 -6.4 ;
      RECT 33.05 -3.29 33.4 -3.17 ;
      RECT 33.05 -0.06 33.4 0.06 ;
      RECT 33.165 -104.945 33.265 -103.985 ;
      RECT 33.165 2.175 33.265 3.135 ;
      RECT 32.875 -112.255 32.975 -111.775 ;
      RECT 32.875 -110.765 32.975 -110.295 ;
      RECT 32.565 -100.19 32.915 -100.07 ;
      RECT 32.565 -96.96 32.915 -96.84 ;
      RECT 32.565 -93.73 32.915 -93.61 ;
      RECT 32.565 -90.5 32.915 -90.38 ;
      RECT 32.565 -87.27 32.915 -87.15 ;
      RECT 32.565 -84.04 32.915 -83.92 ;
      RECT 32.565 -80.81 32.915 -80.69 ;
      RECT 32.565 -77.58 32.915 -77.46 ;
      RECT 32.565 -74.35 32.915 -74.23 ;
      RECT 32.565 -71.12 32.915 -71 ;
      RECT 32.565 -67.89 32.915 -67.77 ;
      RECT 32.565 -64.66 32.915 -64.54 ;
      RECT 32.565 -61.43 32.915 -61.31 ;
      RECT 32.565 -58.2 32.915 -58.08 ;
      RECT 32.565 -54.97 32.915 -54.85 ;
      RECT 32.565 -51.74 32.915 -51.62 ;
      RECT 32.565 -48.51 32.915 -48.39 ;
      RECT 32.565 -45.28 32.915 -45.16 ;
      RECT 32.565 -42.05 32.915 -41.93 ;
      RECT 32.565 -38.82 32.915 -38.7 ;
      RECT 32.565 -35.59 32.915 -35.47 ;
      RECT 32.565 -32.36 32.915 -32.24 ;
      RECT 32.565 -29.13 32.915 -29.01 ;
      RECT 32.565 -25.9 32.915 -25.78 ;
      RECT 32.565 -22.67 32.915 -22.55 ;
      RECT 32.565 -19.44 32.915 -19.32 ;
      RECT 32.565 -16.21 32.915 -16.09 ;
      RECT 32.565 -12.98 32.915 -12.86 ;
      RECT 32.565 -9.75 32.915 -9.63 ;
      RECT 32.565 -6.52 32.915 -6.4 ;
      RECT 32.565 -3.29 32.915 -3.17 ;
      RECT 32.565 -0.06 32.915 0.06 ;
      RECT 32.735 -104.945 32.835 -103.985 ;
      RECT 32.735 2.175 32.835 3.135 ;
      RECT 28.835 -108.655 32.615 -108.535 ;
      RECT 32.475 -104.945 32.575 -103.985 ;
      RECT 32.35 -101.06 32.45 -100.525 ;
      RECT 32.35 -99.735 32.45 -99.2 ;
      RECT 32.35 -97.83 32.45 -97.295 ;
      RECT 32.35 -96.505 32.45 -95.97 ;
      RECT 32.35 -94.6 32.45 -94.065 ;
      RECT 32.35 -93.275 32.45 -92.74 ;
      RECT 32.35 -91.37 32.45 -90.835 ;
      RECT 32.35 -90.045 32.45 -89.51 ;
      RECT 32.35 -88.14 32.45 -87.605 ;
      RECT 32.35 -86.815 32.45 -86.28 ;
      RECT 32.35 -84.91 32.45 -84.375 ;
      RECT 32.35 -83.585 32.45 -83.05 ;
      RECT 32.35 -81.68 32.45 -81.145 ;
      RECT 32.35 -80.355 32.45 -79.82 ;
      RECT 32.35 -78.45 32.45 -77.915 ;
      RECT 32.35 -77.125 32.45 -76.59 ;
      RECT 32.35 -75.22 32.45 -74.685 ;
      RECT 32.35 -73.895 32.45 -73.36 ;
      RECT 32.35 -71.99 32.45 -71.455 ;
      RECT 32.35 -70.665 32.45 -70.13 ;
      RECT 32.35 -68.76 32.45 -68.225 ;
      RECT 32.35 -67.435 32.45 -66.9 ;
      RECT 32.35 -65.53 32.45 -64.995 ;
      RECT 32.35 -64.205 32.45 -63.67 ;
      RECT 32.35 -62.3 32.45 -61.765 ;
      RECT 32.35 -60.975 32.45 -60.44 ;
      RECT 32.35 -59.07 32.45 -58.535 ;
      RECT 32.35 -57.745 32.45 -57.21 ;
      RECT 32.35 -55.84 32.45 -55.305 ;
      RECT 32.35 -54.515 32.45 -53.98 ;
      RECT 32.35 -52.61 32.45 -52.075 ;
      RECT 32.35 -51.285 32.45 -50.75 ;
      RECT 32.35 -49.38 32.45 -48.845 ;
      RECT 32.35 -48.055 32.45 -47.52 ;
      RECT 32.35 -46.15 32.45 -45.615 ;
      RECT 32.35 -44.825 32.45 -44.29 ;
      RECT 32.35 -42.92 32.45 -42.385 ;
      RECT 32.35 -41.595 32.45 -41.06 ;
      RECT 32.35 -39.69 32.45 -39.155 ;
      RECT 32.35 -38.365 32.45 -37.83 ;
      RECT 32.35 -36.46 32.45 -35.925 ;
      RECT 32.35 -35.135 32.45 -34.6 ;
      RECT 32.35 -33.23 32.45 -32.695 ;
      RECT 32.35 -31.905 32.45 -31.37 ;
      RECT 32.35 -30 32.45 -29.465 ;
      RECT 32.35 -28.675 32.45 -28.14 ;
      RECT 32.35 -26.77 32.45 -26.235 ;
      RECT 32.35 -25.445 32.45 -24.91 ;
      RECT 32.35 -23.54 32.45 -23.005 ;
      RECT 32.35 -22.215 32.45 -21.68 ;
      RECT 32.35 -20.31 32.45 -19.775 ;
      RECT 32.35 -18.985 32.45 -18.45 ;
      RECT 32.35 -17.08 32.45 -16.545 ;
      RECT 32.35 -15.755 32.45 -15.22 ;
      RECT 32.35 -13.85 32.45 -13.315 ;
      RECT 32.35 -12.525 32.45 -11.99 ;
      RECT 32.35 -10.62 32.45 -10.085 ;
      RECT 32.35 -9.295 32.45 -8.76 ;
      RECT 32.35 -7.39 32.45 -6.855 ;
      RECT 32.35 -6.065 32.45 -5.53 ;
      RECT 32.35 -4.16 32.45 -3.625 ;
      RECT 32.35 -2.835 32.45 -2.3 ;
      RECT 32.35 -0.93 32.45 -0.395 ;
      RECT 32.35 0.395 32.45 0.93 ;
      RECT 32.285 -110.75 32.405 -110.37 ;
      RECT 32.285 -112.245 32.385 -111.775 ;
      RECT 32.225 -104.945 32.325 -103.985 ;
      RECT 31.85 -100.19 32.2 -100.07 ;
      RECT 31.85 -96.96 32.2 -96.84 ;
      RECT 31.85 -93.73 32.2 -93.61 ;
      RECT 31.85 -90.5 32.2 -90.38 ;
      RECT 31.85 -87.27 32.2 -87.15 ;
      RECT 31.85 -84.04 32.2 -83.92 ;
      RECT 31.85 -80.81 32.2 -80.69 ;
      RECT 31.85 -77.58 32.2 -77.46 ;
      RECT 31.85 -74.35 32.2 -74.23 ;
      RECT 31.85 -71.12 32.2 -71 ;
      RECT 31.85 -67.89 32.2 -67.77 ;
      RECT 31.85 -64.66 32.2 -64.54 ;
      RECT 31.85 -61.43 32.2 -61.31 ;
      RECT 31.85 -58.2 32.2 -58.08 ;
      RECT 31.85 -54.97 32.2 -54.85 ;
      RECT 31.85 -51.74 32.2 -51.62 ;
      RECT 31.85 -48.51 32.2 -48.39 ;
      RECT 31.85 -45.28 32.2 -45.16 ;
      RECT 31.85 -42.05 32.2 -41.93 ;
      RECT 31.85 -38.82 32.2 -38.7 ;
      RECT 31.85 -35.59 32.2 -35.47 ;
      RECT 31.85 -32.36 32.2 -32.24 ;
      RECT 31.85 -29.13 32.2 -29.01 ;
      RECT 31.85 -25.9 32.2 -25.78 ;
      RECT 31.85 -22.67 32.2 -22.55 ;
      RECT 31.85 -19.44 32.2 -19.32 ;
      RECT 31.85 -16.21 32.2 -16.09 ;
      RECT 31.85 -12.98 32.2 -12.86 ;
      RECT 31.85 -9.75 32.2 -9.63 ;
      RECT 31.85 -6.52 32.2 -6.4 ;
      RECT 31.85 -3.29 32.2 -3.17 ;
      RECT 31.85 -0.06 32.2 0.06 ;
      RECT 31.965 -104.945 32.065 -103.985 ;
      RECT 31.965 2.175 32.065 3.135 ;
      RECT 31.695 -109.595 31.83 -109.275 ;
      RECT 31.365 -100.19 31.715 -100.07 ;
      RECT 31.365 -96.96 31.715 -96.84 ;
      RECT 31.365 -93.73 31.715 -93.61 ;
      RECT 31.365 -90.5 31.715 -90.38 ;
      RECT 31.365 -87.27 31.715 -87.15 ;
      RECT 31.365 -84.04 31.715 -83.92 ;
      RECT 31.365 -80.81 31.715 -80.69 ;
      RECT 31.365 -77.58 31.715 -77.46 ;
      RECT 31.365 -74.35 31.715 -74.23 ;
      RECT 31.365 -71.12 31.715 -71 ;
      RECT 31.365 -67.89 31.715 -67.77 ;
      RECT 31.365 -64.66 31.715 -64.54 ;
      RECT 31.365 -61.43 31.715 -61.31 ;
      RECT 31.365 -58.2 31.715 -58.08 ;
      RECT 31.365 -54.97 31.715 -54.85 ;
      RECT 31.365 -51.74 31.715 -51.62 ;
      RECT 31.365 -48.51 31.715 -48.39 ;
      RECT 31.365 -45.28 31.715 -45.16 ;
      RECT 31.365 -42.05 31.715 -41.93 ;
      RECT 31.365 -38.82 31.715 -38.7 ;
      RECT 31.365 -35.59 31.715 -35.47 ;
      RECT 31.365 -32.36 31.715 -32.24 ;
      RECT 31.365 -29.13 31.715 -29.01 ;
      RECT 31.365 -25.9 31.715 -25.78 ;
      RECT 31.365 -22.67 31.715 -22.55 ;
      RECT 31.365 -19.44 31.715 -19.32 ;
      RECT 31.365 -16.21 31.715 -16.09 ;
      RECT 31.365 -12.98 31.715 -12.86 ;
      RECT 31.365 -9.75 31.715 -9.63 ;
      RECT 31.365 -6.52 31.715 -6.4 ;
      RECT 31.365 -3.29 31.715 -3.17 ;
      RECT 31.365 -0.06 31.715 0.06 ;
      RECT 31.535 -104.945 31.635 -103.985 ;
      RECT 31.535 2.175 31.635 3.135 ;
      RECT 31.36 -109.595 31.505 -109.275 ;
      RECT 31.275 -104.945 31.375 -103.985 ;
      RECT 31.15 -101.06 31.25 -100.525 ;
      RECT 31.15 -99.735 31.25 -99.2 ;
      RECT 31.15 -97.83 31.25 -97.295 ;
      RECT 31.15 -96.505 31.25 -95.97 ;
      RECT 31.15 -94.6 31.25 -94.065 ;
      RECT 31.15 -93.275 31.25 -92.74 ;
      RECT 31.15 -91.37 31.25 -90.835 ;
      RECT 31.15 -90.045 31.25 -89.51 ;
      RECT 31.15 -88.14 31.25 -87.605 ;
      RECT 31.15 -86.815 31.25 -86.28 ;
      RECT 31.15 -84.91 31.25 -84.375 ;
      RECT 31.15 -83.585 31.25 -83.05 ;
      RECT 31.15 -81.68 31.25 -81.145 ;
      RECT 31.15 -80.355 31.25 -79.82 ;
      RECT 31.15 -78.45 31.25 -77.915 ;
      RECT 31.15 -77.125 31.25 -76.59 ;
      RECT 31.15 -75.22 31.25 -74.685 ;
      RECT 31.15 -73.895 31.25 -73.36 ;
      RECT 31.15 -71.99 31.25 -71.455 ;
      RECT 31.15 -70.665 31.25 -70.13 ;
      RECT 31.15 -68.76 31.25 -68.225 ;
      RECT 31.15 -67.435 31.25 -66.9 ;
      RECT 31.15 -65.53 31.25 -64.995 ;
      RECT 31.15 -64.205 31.25 -63.67 ;
      RECT 31.15 -62.3 31.25 -61.765 ;
      RECT 31.15 -60.975 31.25 -60.44 ;
      RECT 31.15 -59.07 31.25 -58.535 ;
      RECT 31.15 -57.745 31.25 -57.21 ;
      RECT 31.15 -55.84 31.25 -55.305 ;
      RECT 31.15 -54.515 31.25 -53.98 ;
      RECT 31.15 -52.61 31.25 -52.075 ;
      RECT 31.15 -51.285 31.25 -50.75 ;
      RECT 31.15 -49.38 31.25 -48.845 ;
      RECT 31.15 -48.055 31.25 -47.52 ;
      RECT 31.15 -46.15 31.25 -45.615 ;
      RECT 31.15 -44.825 31.25 -44.29 ;
      RECT 31.15 -42.92 31.25 -42.385 ;
      RECT 31.15 -41.595 31.25 -41.06 ;
      RECT 31.15 -39.69 31.25 -39.155 ;
      RECT 31.15 -38.365 31.25 -37.83 ;
      RECT 31.15 -36.46 31.25 -35.925 ;
      RECT 31.15 -35.135 31.25 -34.6 ;
      RECT 31.15 -33.23 31.25 -32.695 ;
      RECT 31.15 -31.905 31.25 -31.37 ;
      RECT 31.15 -30 31.25 -29.465 ;
      RECT 31.15 -28.675 31.25 -28.14 ;
      RECT 31.15 -26.77 31.25 -26.235 ;
      RECT 31.15 -25.445 31.25 -24.91 ;
      RECT 31.15 -23.54 31.25 -23.005 ;
      RECT 31.15 -22.215 31.25 -21.68 ;
      RECT 31.15 -20.31 31.25 -19.775 ;
      RECT 31.15 -18.985 31.25 -18.45 ;
      RECT 31.15 -17.08 31.25 -16.545 ;
      RECT 31.15 -15.755 31.25 -15.22 ;
      RECT 31.15 -13.85 31.25 -13.315 ;
      RECT 31.15 -12.525 31.25 -11.99 ;
      RECT 31.15 -10.62 31.25 -10.085 ;
      RECT 31.15 -9.295 31.25 -8.76 ;
      RECT 31.15 -7.39 31.25 -6.855 ;
      RECT 31.15 -6.065 31.25 -5.53 ;
      RECT 31.15 -4.16 31.25 -3.625 ;
      RECT 31.15 -2.835 31.25 -2.3 ;
      RECT 31.15 -0.93 31.25 -0.395 ;
      RECT 31.15 0.395 31.25 0.93 ;
      RECT 31.025 -108.175 31.125 -107.215 ;
      RECT 30.65 -100.19 31 -100.07 ;
      RECT 30.65 -96.96 31 -96.84 ;
      RECT 30.65 -93.73 31 -93.61 ;
      RECT 30.65 -90.5 31 -90.38 ;
      RECT 30.65 -87.27 31 -87.15 ;
      RECT 30.65 -84.04 31 -83.92 ;
      RECT 30.65 -80.81 31 -80.69 ;
      RECT 30.65 -77.58 31 -77.46 ;
      RECT 30.65 -74.35 31 -74.23 ;
      RECT 30.65 -71.12 31 -71 ;
      RECT 30.65 -67.89 31 -67.77 ;
      RECT 30.65 -64.66 31 -64.54 ;
      RECT 30.65 -61.43 31 -61.31 ;
      RECT 30.65 -58.2 31 -58.08 ;
      RECT 30.65 -54.97 31 -54.85 ;
      RECT 30.65 -51.74 31 -51.62 ;
      RECT 30.65 -48.51 31 -48.39 ;
      RECT 30.65 -45.28 31 -45.16 ;
      RECT 30.65 -42.05 31 -41.93 ;
      RECT 30.65 -38.82 31 -38.7 ;
      RECT 30.65 -35.59 31 -35.47 ;
      RECT 30.65 -32.36 31 -32.24 ;
      RECT 30.65 -29.13 31 -29.01 ;
      RECT 30.65 -25.9 31 -25.78 ;
      RECT 30.65 -22.67 31 -22.55 ;
      RECT 30.65 -19.44 31 -19.32 ;
      RECT 30.65 -16.21 31 -16.09 ;
      RECT 30.65 -12.98 31 -12.86 ;
      RECT 30.65 -9.75 31 -9.63 ;
      RECT 30.65 -6.52 31 -6.4 ;
      RECT 30.65 -3.29 31 -3.17 ;
      RECT 30.65 -0.06 31 0.06 ;
      RECT 30.855 -112.255 30.955 -111.775 ;
      RECT 30.855 -110.765 30.955 -110.295 ;
      RECT 30.765 -108.175 30.865 -107.215 ;
      RECT 30.765 2.175 30.865 3.135 ;
      RECT 30.165 -100.19 30.515 -100.07 ;
      RECT 30.165 -96.96 30.515 -96.84 ;
      RECT 30.165 -93.73 30.515 -93.61 ;
      RECT 30.165 -90.5 30.515 -90.38 ;
      RECT 30.165 -87.27 30.515 -87.15 ;
      RECT 30.165 -84.04 30.515 -83.92 ;
      RECT 30.165 -80.81 30.515 -80.69 ;
      RECT 30.165 -77.58 30.515 -77.46 ;
      RECT 30.165 -74.35 30.515 -74.23 ;
      RECT 30.165 -71.12 30.515 -71 ;
      RECT 30.165 -67.89 30.515 -67.77 ;
      RECT 30.165 -64.66 30.515 -64.54 ;
      RECT 30.165 -61.43 30.515 -61.31 ;
      RECT 30.165 -58.2 30.515 -58.08 ;
      RECT 30.165 -54.97 30.515 -54.85 ;
      RECT 30.165 -51.74 30.515 -51.62 ;
      RECT 30.165 -48.51 30.515 -48.39 ;
      RECT 30.165 -45.28 30.515 -45.16 ;
      RECT 30.165 -42.05 30.515 -41.93 ;
      RECT 30.165 -38.82 30.515 -38.7 ;
      RECT 30.165 -35.59 30.515 -35.47 ;
      RECT 30.165 -32.36 30.515 -32.24 ;
      RECT 30.165 -29.13 30.515 -29.01 ;
      RECT 30.165 -25.9 30.515 -25.78 ;
      RECT 30.165 -22.67 30.515 -22.55 ;
      RECT 30.165 -19.44 30.515 -19.32 ;
      RECT 30.165 -16.21 30.515 -16.09 ;
      RECT 30.165 -12.98 30.515 -12.86 ;
      RECT 30.165 -9.75 30.515 -9.63 ;
      RECT 30.165 -6.52 30.515 -6.4 ;
      RECT 30.165 -3.29 30.515 -3.17 ;
      RECT 30.165 -0.06 30.515 0.06 ;
      RECT 30.335 -108.175 30.435 -107.215 ;
      RECT 30.335 2.175 30.435 3.135 ;
      RECT 30.23 -110.765 30.4 -110.385 ;
      RECT 30.265 -112.245 30.365 -111.775 ;
      RECT 30.075 -108.175 30.175 -107.215 ;
      RECT 29.95 -101.06 30.05 -100.525 ;
      RECT 29.95 -99.735 30.05 -99.2 ;
      RECT 29.95 -97.83 30.05 -97.295 ;
      RECT 29.95 -96.505 30.05 -95.97 ;
      RECT 29.95 -94.6 30.05 -94.065 ;
      RECT 29.95 -93.275 30.05 -92.74 ;
      RECT 29.95 -91.37 30.05 -90.835 ;
      RECT 29.95 -90.045 30.05 -89.51 ;
      RECT 29.95 -88.14 30.05 -87.605 ;
      RECT 29.95 -86.815 30.05 -86.28 ;
      RECT 29.95 -84.91 30.05 -84.375 ;
      RECT 29.95 -83.585 30.05 -83.05 ;
      RECT 29.95 -81.68 30.05 -81.145 ;
      RECT 29.95 -80.355 30.05 -79.82 ;
      RECT 29.95 -78.45 30.05 -77.915 ;
      RECT 29.95 -77.125 30.05 -76.59 ;
      RECT 29.95 -75.22 30.05 -74.685 ;
      RECT 29.95 -73.895 30.05 -73.36 ;
      RECT 29.95 -71.99 30.05 -71.455 ;
      RECT 29.95 -70.665 30.05 -70.13 ;
      RECT 29.95 -68.76 30.05 -68.225 ;
      RECT 29.95 -67.435 30.05 -66.9 ;
      RECT 29.95 -65.53 30.05 -64.995 ;
      RECT 29.95 -64.205 30.05 -63.67 ;
      RECT 29.95 -62.3 30.05 -61.765 ;
      RECT 29.95 -60.975 30.05 -60.44 ;
      RECT 29.95 -59.07 30.05 -58.535 ;
      RECT 29.95 -57.745 30.05 -57.21 ;
      RECT 29.95 -55.84 30.05 -55.305 ;
      RECT 29.95 -54.515 30.05 -53.98 ;
      RECT 29.95 -52.61 30.05 -52.075 ;
      RECT 29.95 -51.285 30.05 -50.75 ;
      RECT 29.95 -49.38 30.05 -48.845 ;
      RECT 29.95 -48.055 30.05 -47.52 ;
      RECT 29.95 -46.15 30.05 -45.615 ;
      RECT 29.95 -44.825 30.05 -44.29 ;
      RECT 29.95 -42.92 30.05 -42.385 ;
      RECT 29.95 -41.595 30.05 -41.06 ;
      RECT 29.95 -39.69 30.05 -39.155 ;
      RECT 29.95 -38.365 30.05 -37.83 ;
      RECT 29.95 -36.46 30.05 -35.925 ;
      RECT 29.95 -35.135 30.05 -34.6 ;
      RECT 29.95 -33.23 30.05 -32.695 ;
      RECT 29.95 -31.905 30.05 -31.37 ;
      RECT 29.95 -30 30.05 -29.465 ;
      RECT 29.95 -28.675 30.05 -28.14 ;
      RECT 29.95 -26.77 30.05 -26.235 ;
      RECT 29.95 -25.445 30.05 -24.91 ;
      RECT 29.95 -23.54 30.05 -23.005 ;
      RECT 29.95 -22.215 30.05 -21.68 ;
      RECT 29.95 -20.31 30.05 -19.775 ;
      RECT 29.95 -18.985 30.05 -18.45 ;
      RECT 29.95 -17.08 30.05 -16.545 ;
      RECT 29.95 -15.755 30.05 -15.22 ;
      RECT 29.95 -13.85 30.05 -13.315 ;
      RECT 29.95 -12.525 30.05 -11.99 ;
      RECT 29.95 -10.62 30.05 -10.085 ;
      RECT 29.95 -9.295 30.05 -8.76 ;
      RECT 29.95 -7.39 30.05 -6.855 ;
      RECT 29.95 -6.065 30.05 -5.53 ;
      RECT 29.95 -4.16 30.05 -3.625 ;
      RECT 29.95 -2.835 30.05 -2.3 ;
      RECT 29.95 -0.93 30.05 -0.395 ;
      RECT 29.95 0.395 30.05 0.93 ;
      RECT 29.825 -108.175 29.925 -107.215 ;
      RECT 29.45 -100.19 29.8 -100.07 ;
      RECT 29.45 -96.96 29.8 -96.84 ;
      RECT 29.45 -93.73 29.8 -93.61 ;
      RECT 29.45 -90.5 29.8 -90.38 ;
      RECT 29.45 -87.27 29.8 -87.15 ;
      RECT 29.45 -84.04 29.8 -83.92 ;
      RECT 29.45 -80.81 29.8 -80.69 ;
      RECT 29.45 -77.58 29.8 -77.46 ;
      RECT 29.45 -74.35 29.8 -74.23 ;
      RECT 29.45 -71.12 29.8 -71 ;
      RECT 29.45 -67.89 29.8 -67.77 ;
      RECT 29.45 -64.66 29.8 -64.54 ;
      RECT 29.45 -61.43 29.8 -61.31 ;
      RECT 29.45 -58.2 29.8 -58.08 ;
      RECT 29.45 -54.97 29.8 -54.85 ;
      RECT 29.45 -51.74 29.8 -51.62 ;
      RECT 29.45 -48.51 29.8 -48.39 ;
      RECT 29.45 -45.28 29.8 -45.16 ;
      RECT 29.45 -42.05 29.8 -41.93 ;
      RECT 29.45 -38.82 29.8 -38.7 ;
      RECT 29.45 -35.59 29.8 -35.47 ;
      RECT 29.45 -32.36 29.8 -32.24 ;
      RECT 29.45 -29.13 29.8 -29.01 ;
      RECT 29.45 -25.9 29.8 -25.78 ;
      RECT 29.45 -22.67 29.8 -22.55 ;
      RECT 29.45 -19.44 29.8 -19.32 ;
      RECT 29.45 -16.21 29.8 -16.09 ;
      RECT 29.45 -12.98 29.8 -12.86 ;
      RECT 29.45 -9.75 29.8 -9.63 ;
      RECT 29.45 -6.52 29.8 -6.4 ;
      RECT 29.45 -3.29 29.8 -3.17 ;
      RECT 29.45 -0.06 29.8 0.06 ;
      RECT 29.565 -108.175 29.665 -107.215 ;
      RECT 29.565 2.175 29.665 3.135 ;
      RECT 29.465 -113.555 29.565 -113.085 ;
      RECT 28.965 -100.19 29.315 -100.07 ;
      RECT 28.965 -96.96 29.315 -96.84 ;
      RECT 28.965 -93.73 29.315 -93.61 ;
      RECT 28.965 -90.5 29.315 -90.38 ;
      RECT 28.965 -87.27 29.315 -87.15 ;
      RECT 28.965 -84.04 29.315 -83.92 ;
      RECT 28.965 -80.81 29.315 -80.69 ;
      RECT 28.965 -77.58 29.315 -77.46 ;
      RECT 28.965 -74.35 29.315 -74.23 ;
      RECT 28.965 -71.12 29.315 -71 ;
      RECT 28.965 -67.89 29.315 -67.77 ;
      RECT 28.965 -64.66 29.315 -64.54 ;
      RECT 28.965 -61.43 29.315 -61.31 ;
      RECT 28.965 -58.2 29.315 -58.08 ;
      RECT 28.965 -54.97 29.315 -54.85 ;
      RECT 28.965 -51.74 29.315 -51.62 ;
      RECT 28.965 -48.51 29.315 -48.39 ;
      RECT 28.965 -45.28 29.315 -45.16 ;
      RECT 28.965 -42.05 29.315 -41.93 ;
      RECT 28.965 -38.82 29.315 -38.7 ;
      RECT 28.965 -35.59 29.315 -35.47 ;
      RECT 28.965 -32.36 29.315 -32.24 ;
      RECT 28.965 -29.13 29.315 -29.01 ;
      RECT 28.965 -25.9 29.315 -25.78 ;
      RECT 28.965 -22.67 29.315 -22.55 ;
      RECT 28.965 -19.44 29.315 -19.32 ;
      RECT 28.965 -16.21 29.315 -16.09 ;
      RECT 28.965 -12.98 29.315 -12.86 ;
      RECT 28.965 -9.75 29.315 -9.63 ;
      RECT 28.965 -6.52 29.315 -6.4 ;
      RECT 28.965 -3.29 29.315 -3.17 ;
      RECT 28.965 -0.06 29.315 0.06 ;
      RECT 29.1 -110.735 29.25 -110.445 ;
      RECT 29.135 -108.175 29.235 -107.215 ;
      RECT 29.135 2.175 29.235 3.135 ;
      RECT 29.115 -112.19 29.215 -111.65 ;
      RECT 28.875 -113.555 28.975 -113.085 ;
      RECT 28.875 -108.175 28.975 -107.215 ;
      RECT 28.75 -101.06 28.85 -100.525 ;
      RECT 28.75 -99.735 28.85 -99.2 ;
      RECT 28.75 -97.83 28.85 -97.295 ;
      RECT 28.75 -96.505 28.85 -95.97 ;
      RECT 28.75 -94.6 28.85 -94.065 ;
      RECT 28.75 -93.275 28.85 -92.74 ;
      RECT 28.75 -91.37 28.85 -90.835 ;
      RECT 28.75 -90.045 28.85 -89.51 ;
      RECT 28.75 -88.14 28.85 -87.605 ;
      RECT 28.75 -86.815 28.85 -86.28 ;
      RECT 28.75 -84.91 28.85 -84.375 ;
      RECT 28.75 -83.585 28.85 -83.05 ;
      RECT 28.75 -81.68 28.85 -81.145 ;
      RECT 28.75 -80.355 28.85 -79.82 ;
      RECT 28.75 -78.45 28.85 -77.915 ;
      RECT 28.75 -77.125 28.85 -76.59 ;
      RECT 28.75 -75.22 28.85 -74.685 ;
      RECT 28.75 -73.895 28.85 -73.36 ;
      RECT 28.75 -71.99 28.85 -71.455 ;
      RECT 28.75 -70.665 28.85 -70.13 ;
      RECT 28.75 -68.76 28.85 -68.225 ;
      RECT 28.75 -67.435 28.85 -66.9 ;
      RECT 28.75 -65.53 28.85 -64.995 ;
      RECT 28.75 -64.205 28.85 -63.67 ;
      RECT 28.75 -62.3 28.85 -61.765 ;
      RECT 28.75 -60.975 28.85 -60.44 ;
      RECT 28.75 -59.07 28.85 -58.535 ;
      RECT 28.75 -57.745 28.85 -57.21 ;
      RECT 28.75 -55.84 28.85 -55.305 ;
      RECT 28.75 -54.515 28.85 -53.98 ;
      RECT 28.75 -52.61 28.85 -52.075 ;
      RECT 28.75 -51.285 28.85 -50.75 ;
      RECT 28.75 -49.38 28.85 -48.845 ;
      RECT 28.75 -48.055 28.85 -47.52 ;
      RECT 28.75 -46.15 28.85 -45.615 ;
      RECT 28.75 -44.825 28.85 -44.29 ;
      RECT 28.75 -42.92 28.85 -42.385 ;
      RECT 28.75 -41.595 28.85 -41.06 ;
      RECT 28.75 -39.69 28.85 -39.155 ;
      RECT 28.75 -38.365 28.85 -37.83 ;
      RECT 28.75 -36.46 28.85 -35.925 ;
      RECT 28.75 -35.135 28.85 -34.6 ;
      RECT 28.75 -33.23 28.85 -32.695 ;
      RECT 28.75 -31.905 28.85 -31.37 ;
      RECT 28.75 -30 28.85 -29.465 ;
      RECT 28.75 -28.675 28.85 -28.14 ;
      RECT 28.75 -26.77 28.85 -26.235 ;
      RECT 28.75 -25.445 28.85 -24.91 ;
      RECT 28.75 -23.54 28.85 -23.005 ;
      RECT 28.75 -22.215 28.85 -21.68 ;
      RECT 28.75 -20.31 28.85 -19.775 ;
      RECT 28.75 -18.985 28.85 -18.45 ;
      RECT 28.75 -17.08 28.85 -16.545 ;
      RECT 28.75 -15.755 28.85 -15.22 ;
      RECT 28.75 -13.85 28.85 -13.315 ;
      RECT 28.75 -12.525 28.85 -11.99 ;
      RECT 28.75 -10.62 28.85 -10.085 ;
      RECT 28.75 -9.295 28.85 -8.76 ;
      RECT 28.75 -7.39 28.85 -6.855 ;
      RECT 28.75 -6.065 28.85 -5.53 ;
      RECT 28.75 -4.16 28.85 -3.625 ;
      RECT 28.75 -2.835 28.85 -2.3 ;
      RECT 28.75 -0.93 28.85 -0.395 ;
      RECT 28.75 0.395 28.85 0.93 ;
      RECT 28.625 -104.945 28.725 -103.985 ;
      RECT 28.25 -100.19 28.6 -100.07 ;
      RECT 28.25 -96.96 28.6 -96.84 ;
      RECT 28.25 -93.73 28.6 -93.61 ;
      RECT 28.25 -90.5 28.6 -90.38 ;
      RECT 28.25 -87.27 28.6 -87.15 ;
      RECT 28.25 -84.04 28.6 -83.92 ;
      RECT 28.25 -80.81 28.6 -80.69 ;
      RECT 28.25 -77.58 28.6 -77.46 ;
      RECT 28.25 -74.35 28.6 -74.23 ;
      RECT 28.25 -71.12 28.6 -71 ;
      RECT 28.25 -67.89 28.6 -67.77 ;
      RECT 28.25 -64.66 28.6 -64.54 ;
      RECT 28.25 -61.43 28.6 -61.31 ;
      RECT 28.25 -58.2 28.6 -58.08 ;
      RECT 28.25 -54.97 28.6 -54.85 ;
      RECT 28.25 -51.74 28.6 -51.62 ;
      RECT 28.25 -48.51 28.6 -48.39 ;
      RECT 28.25 -45.28 28.6 -45.16 ;
      RECT 28.25 -42.05 28.6 -41.93 ;
      RECT 28.25 -38.82 28.6 -38.7 ;
      RECT 28.25 -35.59 28.6 -35.47 ;
      RECT 28.25 -32.36 28.6 -32.24 ;
      RECT 28.25 -29.13 28.6 -29.01 ;
      RECT 28.25 -25.9 28.6 -25.78 ;
      RECT 28.25 -22.67 28.6 -22.55 ;
      RECT 28.25 -19.44 28.6 -19.32 ;
      RECT 28.25 -16.21 28.6 -16.09 ;
      RECT 28.25 -12.98 28.6 -12.86 ;
      RECT 28.25 -9.75 28.6 -9.63 ;
      RECT 28.25 -6.52 28.6 -6.4 ;
      RECT 28.25 -3.29 28.6 -3.17 ;
      RECT 28.25 -0.06 28.6 0.06 ;
      RECT 28.365 -104.945 28.465 -103.985 ;
      RECT 28.365 2.175 28.465 3.135 ;
      RECT 28.075 -112.255 28.175 -111.775 ;
      RECT 28.075 -110.765 28.175 -110.295 ;
      RECT 27.765 -100.19 28.115 -100.07 ;
      RECT 27.765 -96.96 28.115 -96.84 ;
      RECT 27.765 -93.73 28.115 -93.61 ;
      RECT 27.765 -90.5 28.115 -90.38 ;
      RECT 27.765 -87.27 28.115 -87.15 ;
      RECT 27.765 -84.04 28.115 -83.92 ;
      RECT 27.765 -80.81 28.115 -80.69 ;
      RECT 27.765 -77.58 28.115 -77.46 ;
      RECT 27.765 -74.35 28.115 -74.23 ;
      RECT 27.765 -71.12 28.115 -71 ;
      RECT 27.765 -67.89 28.115 -67.77 ;
      RECT 27.765 -64.66 28.115 -64.54 ;
      RECT 27.765 -61.43 28.115 -61.31 ;
      RECT 27.765 -58.2 28.115 -58.08 ;
      RECT 27.765 -54.97 28.115 -54.85 ;
      RECT 27.765 -51.74 28.115 -51.62 ;
      RECT 27.765 -48.51 28.115 -48.39 ;
      RECT 27.765 -45.28 28.115 -45.16 ;
      RECT 27.765 -42.05 28.115 -41.93 ;
      RECT 27.765 -38.82 28.115 -38.7 ;
      RECT 27.765 -35.59 28.115 -35.47 ;
      RECT 27.765 -32.36 28.115 -32.24 ;
      RECT 27.765 -29.13 28.115 -29.01 ;
      RECT 27.765 -25.9 28.115 -25.78 ;
      RECT 27.765 -22.67 28.115 -22.55 ;
      RECT 27.765 -19.44 28.115 -19.32 ;
      RECT 27.765 -16.21 28.115 -16.09 ;
      RECT 27.765 -12.98 28.115 -12.86 ;
      RECT 27.765 -9.75 28.115 -9.63 ;
      RECT 27.765 -6.52 28.115 -6.4 ;
      RECT 27.765 -3.29 28.115 -3.17 ;
      RECT 27.765 -0.06 28.115 0.06 ;
      RECT 27.935 -104.945 28.035 -103.985 ;
      RECT 27.935 2.175 28.035 3.135 ;
      RECT 24.035 -108.655 27.815 -108.535 ;
      RECT 27.675 -104.945 27.775 -103.985 ;
      RECT 27.55 -101.06 27.65 -100.525 ;
      RECT 27.55 -99.735 27.65 -99.2 ;
      RECT 27.55 -97.83 27.65 -97.295 ;
      RECT 27.55 -96.505 27.65 -95.97 ;
      RECT 27.55 -94.6 27.65 -94.065 ;
      RECT 27.55 -93.275 27.65 -92.74 ;
      RECT 27.55 -91.37 27.65 -90.835 ;
      RECT 27.55 -90.045 27.65 -89.51 ;
      RECT 27.55 -88.14 27.65 -87.605 ;
      RECT 27.55 -86.815 27.65 -86.28 ;
      RECT 27.55 -84.91 27.65 -84.375 ;
      RECT 27.55 -83.585 27.65 -83.05 ;
      RECT 27.55 -81.68 27.65 -81.145 ;
      RECT 27.55 -80.355 27.65 -79.82 ;
      RECT 27.55 -78.45 27.65 -77.915 ;
      RECT 27.55 -77.125 27.65 -76.59 ;
      RECT 27.55 -75.22 27.65 -74.685 ;
      RECT 27.55 -73.895 27.65 -73.36 ;
      RECT 27.55 -71.99 27.65 -71.455 ;
      RECT 27.55 -70.665 27.65 -70.13 ;
      RECT 27.55 -68.76 27.65 -68.225 ;
      RECT 27.55 -67.435 27.65 -66.9 ;
      RECT 27.55 -65.53 27.65 -64.995 ;
      RECT 27.55 -64.205 27.65 -63.67 ;
      RECT 27.55 -62.3 27.65 -61.765 ;
      RECT 27.55 -60.975 27.65 -60.44 ;
      RECT 27.55 -59.07 27.65 -58.535 ;
      RECT 27.55 -57.745 27.65 -57.21 ;
      RECT 27.55 -55.84 27.65 -55.305 ;
      RECT 27.55 -54.515 27.65 -53.98 ;
      RECT 27.55 -52.61 27.65 -52.075 ;
      RECT 27.55 -51.285 27.65 -50.75 ;
      RECT 27.55 -49.38 27.65 -48.845 ;
      RECT 27.55 -48.055 27.65 -47.52 ;
      RECT 27.55 -46.15 27.65 -45.615 ;
      RECT 27.55 -44.825 27.65 -44.29 ;
      RECT 27.55 -42.92 27.65 -42.385 ;
      RECT 27.55 -41.595 27.65 -41.06 ;
      RECT 27.55 -39.69 27.65 -39.155 ;
      RECT 27.55 -38.365 27.65 -37.83 ;
      RECT 27.55 -36.46 27.65 -35.925 ;
      RECT 27.55 -35.135 27.65 -34.6 ;
      RECT 27.55 -33.23 27.65 -32.695 ;
      RECT 27.55 -31.905 27.65 -31.37 ;
      RECT 27.55 -30 27.65 -29.465 ;
      RECT 27.55 -28.675 27.65 -28.14 ;
      RECT 27.55 -26.77 27.65 -26.235 ;
      RECT 27.55 -25.445 27.65 -24.91 ;
      RECT 27.55 -23.54 27.65 -23.005 ;
      RECT 27.55 -22.215 27.65 -21.68 ;
      RECT 27.55 -20.31 27.65 -19.775 ;
      RECT 27.55 -18.985 27.65 -18.45 ;
      RECT 27.55 -17.08 27.65 -16.545 ;
      RECT 27.55 -15.755 27.65 -15.22 ;
      RECT 27.55 -13.85 27.65 -13.315 ;
      RECT 27.55 -12.525 27.65 -11.99 ;
      RECT 27.55 -10.62 27.65 -10.085 ;
      RECT 27.55 -9.295 27.65 -8.76 ;
      RECT 27.55 -7.39 27.65 -6.855 ;
      RECT 27.55 -6.065 27.65 -5.53 ;
      RECT 27.55 -4.16 27.65 -3.625 ;
      RECT 27.55 -2.835 27.65 -2.3 ;
      RECT 27.55 -0.93 27.65 -0.395 ;
      RECT 27.55 0.395 27.65 0.93 ;
      RECT 27.485 -110.75 27.605 -110.37 ;
      RECT 27.485 -112.245 27.585 -111.775 ;
      RECT 27.425 -104.945 27.525 -103.985 ;
      RECT 27.05 -100.19 27.4 -100.07 ;
      RECT 27.05 -96.96 27.4 -96.84 ;
      RECT 27.05 -93.73 27.4 -93.61 ;
      RECT 27.05 -90.5 27.4 -90.38 ;
      RECT 27.05 -87.27 27.4 -87.15 ;
      RECT 27.05 -84.04 27.4 -83.92 ;
      RECT 27.05 -80.81 27.4 -80.69 ;
      RECT 27.05 -77.58 27.4 -77.46 ;
      RECT 27.05 -74.35 27.4 -74.23 ;
      RECT 27.05 -71.12 27.4 -71 ;
      RECT 27.05 -67.89 27.4 -67.77 ;
      RECT 27.05 -64.66 27.4 -64.54 ;
      RECT 27.05 -61.43 27.4 -61.31 ;
      RECT 27.05 -58.2 27.4 -58.08 ;
      RECT 27.05 -54.97 27.4 -54.85 ;
      RECT 27.05 -51.74 27.4 -51.62 ;
      RECT 27.05 -48.51 27.4 -48.39 ;
      RECT 27.05 -45.28 27.4 -45.16 ;
      RECT 27.05 -42.05 27.4 -41.93 ;
      RECT 27.05 -38.82 27.4 -38.7 ;
      RECT 27.05 -35.59 27.4 -35.47 ;
      RECT 27.05 -32.36 27.4 -32.24 ;
      RECT 27.05 -29.13 27.4 -29.01 ;
      RECT 27.05 -25.9 27.4 -25.78 ;
      RECT 27.05 -22.67 27.4 -22.55 ;
      RECT 27.05 -19.44 27.4 -19.32 ;
      RECT 27.05 -16.21 27.4 -16.09 ;
      RECT 27.05 -12.98 27.4 -12.86 ;
      RECT 27.05 -9.75 27.4 -9.63 ;
      RECT 27.05 -6.52 27.4 -6.4 ;
      RECT 27.05 -3.29 27.4 -3.17 ;
      RECT 27.05 -0.06 27.4 0.06 ;
      RECT 27.165 -104.945 27.265 -103.985 ;
      RECT 27.165 2.175 27.265 3.135 ;
      RECT 26.895 -109.595 27.03 -109.275 ;
      RECT 26.565 -100.19 26.915 -100.07 ;
      RECT 26.565 -96.96 26.915 -96.84 ;
      RECT 26.565 -93.73 26.915 -93.61 ;
      RECT 26.565 -90.5 26.915 -90.38 ;
      RECT 26.565 -87.27 26.915 -87.15 ;
      RECT 26.565 -84.04 26.915 -83.92 ;
      RECT 26.565 -80.81 26.915 -80.69 ;
      RECT 26.565 -77.58 26.915 -77.46 ;
      RECT 26.565 -74.35 26.915 -74.23 ;
      RECT 26.565 -71.12 26.915 -71 ;
      RECT 26.565 -67.89 26.915 -67.77 ;
      RECT 26.565 -64.66 26.915 -64.54 ;
      RECT 26.565 -61.43 26.915 -61.31 ;
      RECT 26.565 -58.2 26.915 -58.08 ;
      RECT 26.565 -54.97 26.915 -54.85 ;
      RECT 26.565 -51.74 26.915 -51.62 ;
      RECT 26.565 -48.51 26.915 -48.39 ;
      RECT 26.565 -45.28 26.915 -45.16 ;
      RECT 26.565 -42.05 26.915 -41.93 ;
      RECT 26.565 -38.82 26.915 -38.7 ;
      RECT 26.565 -35.59 26.915 -35.47 ;
      RECT 26.565 -32.36 26.915 -32.24 ;
      RECT 26.565 -29.13 26.915 -29.01 ;
      RECT 26.565 -25.9 26.915 -25.78 ;
      RECT 26.565 -22.67 26.915 -22.55 ;
      RECT 26.565 -19.44 26.915 -19.32 ;
      RECT 26.565 -16.21 26.915 -16.09 ;
      RECT 26.565 -12.98 26.915 -12.86 ;
      RECT 26.565 -9.75 26.915 -9.63 ;
      RECT 26.565 -6.52 26.915 -6.4 ;
      RECT 26.565 -3.29 26.915 -3.17 ;
      RECT 26.565 -0.06 26.915 0.06 ;
      RECT 26.735 -104.945 26.835 -103.985 ;
      RECT 26.735 2.175 26.835 3.135 ;
      RECT 26.56 -109.595 26.705 -109.275 ;
      RECT 26.475 -104.945 26.575 -103.985 ;
      RECT 26.35 -101.06 26.45 -100.525 ;
      RECT 26.35 -99.735 26.45 -99.2 ;
      RECT 26.35 -97.83 26.45 -97.295 ;
      RECT 26.35 -96.505 26.45 -95.97 ;
      RECT 26.35 -94.6 26.45 -94.065 ;
      RECT 26.35 -93.275 26.45 -92.74 ;
      RECT 26.35 -91.37 26.45 -90.835 ;
      RECT 26.35 -90.045 26.45 -89.51 ;
      RECT 26.35 -88.14 26.45 -87.605 ;
      RECT 26.35 -86.815 26.45 -86.28 ;
      RECT 26.35 -84.91 26.45 -84.375 ;
      RECT 26.35 -83.585 26.45 -83.05 ;
      RECT 26.35 -81.68 26.45 -81.145 ;
      RECT 26.35 -80.355 26.45 -79.82 ;
      RECT 26.35 -78.45 26.45 -77.915 ;
      RECT 26.35 -77.125 26.45 -76.59 ;
      RECT 26.35 -75.22 26.45 -74.685 ;
      RECT 26.35 -73.895 26.45 -73.36 ;
      RECT 26.35 -71.99 26.45 -71.455 ;
      RECT 26.35 -70.665 26.45 -70.13 ;
      RECT 26.35 -68.76 26.45 -68.225 ;
      RECT 26.35 -67.435 26.45 -66.9 ;
      RECT 26.35 -65.53 26.45 -64.995 ;
      RECT 26.35 -64.205 26.45 -63.67 ;
      RECT 26.35 -62.3 26.45 -61.765 ;
      RECT 26.35 -60.975 26.45 -60.44 ;
      RECT 26.35 -59.07 26.45 -58.535 ;
      RECT 26.35 -57.745 26.45 -57.21 ;
      RECT 26.35 -55.84 26.45 -55.305 ;
      RECT 26.35 -54.515 26.45 -53.98 ;
      RECT 26.35 -52.61 26.45 -52.075 ;
      RECT 26.35 -51.285 26.45 -50.75 ;
      RECT 26.35 -49.38 26.45 -48.845 ;
      RECT 26.35 -48.055 26.45 -47.52 ;
      RECT 26.35 -46.15 26.45 -45.615 ;
      RECT 26.35 -44.825 26.45 -44.29 ;
      RECT 26.35 -42.92 26.45 -42.385 ;
      RECT 26.35 -41.595 26.45 -41.06 ;
      RECT 26.35 -39.69 26.45 -39.155 ;
      RECT 26.35 -38.365 26.45 -37.83 ;
      RECT 26.35 -36.46 26.45 -35.925 ;
      RECT 26.35 -35.135 26.45 -34.6 ;
      RECT 26.35 -33.23 26.45 -32.695 ;
      RECT 26.35 -31.905 26.45 -31.37 ;
      RECT 26.35 -30 26.45 -29.465 ;
      RECT 26.35 -28.675 26.45 -28.14 ;
      RECT 26.35 -26.77 26.45 -26.235 ;
      RECT 26.35 -25.445 26.45 -24.91 ;
      RECT 26.35 -23.54 26.45 -23.005 ;
      RECT 26.35 -22.215 26.45 -21.68 ;
      RECT 26.35 -20.31 26.45 -19.775 ;
      RECT 26.35 -18.985 26.45 -18.45 ;
      RECT 26.35 -17.08 26.45 -16.545 ;
      RECT 26.35 -15.755 26.45 -15.22 ;
      RECT 26.35 -13.85 26.45 -13.315 ;
      RECT 26.35 -12.525 26.45 -11.99 ;
      RECT 26.35 -10.62 26.45 -10.085 ;
      RECT 26.35 -9.295 26.45 -8.76 ;
      RECT 26.35 -7.39 26.45 -6.855 ;
      RECT 26.35 -6.065 26.45 -5.53 ;
      RECT 26.35 -4.16 26.45 -3.625 ;
      RECT 26.35 -2.835 26.45 -2.3 ;
      RECT 26.35 -0.93 26.45 -0.395 ;
      RECT 26.35 0.395 26.45 0.93 ;
      RECT 26.225 -108.175 26.325 -107.215 ;
      RECT 25.85 -100.19 26.2 -100.07 ;
      RECT 25.85 -96.96 26.2 -96.84 ;
      RECT 25.85 -93.73 26.2 -93.61 ;
      RECT 25.85 -90.5 26.2 -90.38 ;
      RECT 25.85 -87.27 26.2 -87.15 ;
      RECT 25.85 -84.04 26.2 -83.92 ;
      RECT 25.85 -80.81 26.2 -80.69 ;
      RECT 25.85 -77.58 26.2 -77.46 ;
      RECT 25.85 -74.35 26.2 -74.23 ;
      RECT 25.85 -71.12 26.2 -71 ;
      RECT 25.85 -67.89 26.2 -67.77 ;
      RECT 25.85 -64.66 26.2 -64.54 ;
      RECT 25.85 -61.43 26.2 -61.31 ;
      RECT 25.85 -58.2 26.2 -58.08 ;
      RECT 25.85 -54.97 26.2 -54.85 ;
      RECT 25.85 -51.74 26.2 -51.62 ;
      RECT 25.85 -48.51 26.2 -48.39 ;
      RECT 25.85 -45.28 26.2 -45.16 ;
      RECT 25.85 -42.05 26.2 -41.93 ;
      RECT 25.85 -38.82 26.2 -38.7 ;
      RECT 25.85 -35.59 26.2 -35.47 ;
      RECT 25.85 -32.36 26.2 -32.24 ;
      RECT 25.85 -29.13 26.2 -29.01 ;
      RECT 25.85 -25.9 26.2 -25.78 ;
      RECT 25.85 -22.67 26.2 -22.55 ;
      RECT 25.85 -19.44 26.2 -19.32 ;
      RECT 25.85 -16.21 26.2 -16.09 ;
      RECT 25.85 -12.98 26.2 -12.86 ;
      RECT 25.85 -9.75 26.2 -9.63 ;
      RECT 25.85 -6.52 26.2 -6.4 ;
      RECT 25.85 -3.29 26.2 -3.17 ;
      RECT 25.85 -0.06 26.2 0.06 ;
      RECT 26.055 -112.255 26.155 -111.775 ;
      RECT 26.055 -110.765 26.155 -110.295 ;
      RECT 25.965 -108.175 26.065 -107.215 ;
      RECT 25.965 2.175 26.065 3.135 ;
      RECT 25.365 -100.19 25.715 -100.07 ;
      RECT 25.365 -96.96 25.715 -96.84 ;
      RECT 25.365 -93.73 25.715 -93.61 ;
      RECT 25.365 -90.5 25.715 -90.38 ;
      RECT 25.365 -87.27 25.715 -87.15 ;
      RECT 25.365 -84.04 25.715 -83.92 ;
      RECT 25.365 -80.81 25.715 -80.69 ;
      RECT 25.365 -77.58 25.715 -77.46 ;
      RECT 25.365 -74.35 25.715 -74.23 ;
      RECT 25.365 -71.12 25.715 -71 ;
      RECT 25.365 -67.89 25.715 -67.77 ;
      RECT 25.365 -64.66 25.715 -64.54 ;
      RECT 25.365 -61.43 25.715 -61.31 ;
      RECT 25.365 -58.2 25.715 -58.08 ;
      RECT 25.365 -54.97 25.715 -54.85 ;
      RECT 25.365 -51.74 25.715 -51.62 ;
      RECT 25.365 -48.51 25.715 -48.39 ;
      RECT 25.365 -45.28 25.715 -45.16 ;
      RECT 25.365 -42.05 25.715 -41.93 ;
      RECT 25.365 -38.82 25.715 -38.7 ;
      RECT 25.365 -35.59 25.715 -35.47 ;
      RECT 25.365 -32.36 25.715 -32.24 ;
      RECT 25.365 -29.13 25.715 -29.01 ;
      RECT 25.365 -25.9 25.715 -25.78 ;
      RECT 25.365 -22.67 25.715 -22.55 ;
      RECT 25.365 -19.44 25.715 -19.32 ;
      RECT 25.365 -16.21 25.715 -16.09 ;
      RECT 25.365 -12.98 25.715 -12.86 ;
      RECT 25.365 -9.75 25.715 -9.63 ;
      RECT 25.365 -6.52 25.715 -6.4 ;
      RECT 25.365 -3.29 25.715 -3.17 ;
      RECT 25.365 -0.06 25.715 0.06 ;
      RECT 25.535 -108.175 25.635 -107.215 ;
      RECT 25.535 2.175 25.635 3.135 ;
      RECT 25.43 -110.765 25.6 -110.385 ;
      RECT 25.465 -112.245 25.565 -111.775 ;
      RECT 25.275 -108.175 25.375 -107.215 ;
      RECT 25.15 -101.06 25.25 -100.525 ;
      RECT 25.15 -99.735 25.25 -99.2 ;
      RECT 25.15 -97.83 25.25 -97.295 ;
      RECT 25.15 -96.505 25.25 -95.97 ;
      RECT 25.15 -94.6 25.25 -94.065 ;
      RECT 25.15 -93.275 25.25 -92.74 ;
      RECT 25.15 -91.37 25.25 -90.835 ;
      RECT 25.15 -90.045 25.25 -89.51 ;
      RECT 25.15 -88.14 25.25 -87.605 ;
      RECT 25.15 -86.815 25.25 -86.28 ;
      RECT 25.15 -84.91 25.25 -84.375 ;
      RECT 25.15 -83.585 25.25 -83.05 ;
      RECT 25.15 -81.68 25.25 -81.145 ;
      RECT 25.15 -80.355 25.25 -79.82 ;
      RECT 25.15 -78.45 25.25 -77.915 ;
      RECT 25.15 -77.125 25.25 -76.59 ;
      RECT 25.15 -75.22 25.25 -74.685 ;
      RECT 25.15 -73.895 25.25 -73.36 ;
      RECT 25.15 -71.99 25.25 -71.455 ;
      RECT 25.15 -70.665 25.25 -70.13 ;
      RECT 25.15 -68.76 25.25 -68.225 ;
      RECT 25.15 -67.435 25.25 -66.9 ;
      RECT 25.15 -65.53 25.25 -64.995 ;
      RECT 25.15 -64.205 25.25 -63.67 ;
      RECT 25.15 -62.3 25.25 -61.765 ;
      RECT 25.15 -60.975 25.25 -60.44 ;
      RECT 25.15 -59.07 25.25 -58.535 ;
      RECT 25.15 -57.745 25.25 -57.21 ;
      RECT 25.15 -55.84 25.25 -55.305 ;
      RECT 25.15 -54.515 25.25 -53.98 ;
      RECT 25.15 -52.61 25.25 -52.075 ;
      RECT 25.15 -51.285 25.25 -50.75 ;
      RECT 25.15 -49.38 25.25 -48.845 ;
      RECT 25.15 -48.055 25.25 -47.52 ;
      RECT 25.15 -46.15 25.25 -45.615 ;
      RECT 25.15 -44.825 25.25 -44.29 ;
      RECT 25.15 -42.92 25.25 -42.385 ;
      RECT 25.15 -41.595 25.25 -41.06 ;
      RECT 25.15 -39.69 25.25 -39.155 ;
      RECT 25.15 -38.365 25.25 -37.83 ;
      RECT 25.15 -36.46 25.25 -35.925 ;
      RECT 25.15 -35.135 25.25 -34.6 ;
      RECT 25.15 -33.23 25.25 -32.695 ;
      RECT 25.15 -31.905 25.25 -31.37 ;
      RECT 25.15 -30 25.25 -29.465 ;
      RECT 25.15 -28.675 25.25 -28.14 ;
      RECT 25.15 -26.77 25.25 -26.235 ;
      RECT 25.15 -25.445 25.25 -24.91 ;
      RECT 25.15 -23.54 25.25 -23.005 ;
      RECT 25.15 -22.215 25.25 -21.68 ;
      RECT 25.15 -20.31 25.25 -19.775 ;
      RECT 25.15 -18.985 25.25 -18.45 ;
      RECT 25.15 -17.08 25.25 -16.545 ;
      RECT 25.15 -15.755 25.25 -15.22 ;
      RECT 25.15 -13.85 25.25 -13.315 ;
      RECT 25.15 -12.525 25.25 -11.99 ;
      RECT 25.15 -10.62 25.25 -10.085 ;
      RECT 25.15 -9.295 25.25 -8.76 ;
      RECT 25.15 -7.39 25.25 -6.855 ;
      RECT 25.15 -6.065 25.25 -5.53 ;
      RECT 25.15 -4.16 25.25 -3.625 ;
      RECT 25.15 -2.835 25.25 -2.3 ;
      RECT 25.15 -0.93 25.25 -0.395 ;
      RECT 25.15 0.395 25.25 0.93 ;
      RECT 25.025 -108.175 25.125 -107.215 ;
      RECT 24.65 -100.19 25 -100.07 ;
      RECT 24.65 -96.96 25 -96.84 ;
      RECT 24.65 -93.73 25 -93.61 ;
      RECT 24.65 -90.5 25 -90.38 ;
      RECT 24.65 -87.27 25 -87.15 ;
      RECT 24.65 -84.04 25 -83.92 ;
      RECT 24.65 -80.81 25 -80.69 ;
      RECT 24.65 -77.58 25 -77.46 ;
      RECT 24.65 -74.35 25 -74.23 ;
      RECT 24.65 -71.12 25 -71 ;
      RECT 24.65 -67.89 25 -67.77 ;
      RECT 24.65 -64.66 25 -64.54 ;
      RECT 24.65 -61.43 25 -61.31 ;
      RECT 24.65 -58.2 25 -58.08 ;
      RECT 24.65 -54.97 25 -54.85 ;
      RECT 24.65 -51.74 25 -51.62 ;
      RECT 24.65 -48.51 25 -48.39 ;
      RECT 24.65 -45.28 25 -45.16 ;
      RECT 24.65 -42.05 25 -41.93 ;
      RECT 24.65 -38.82 25 -38.7 ;
      RECT 24.65 -35.59 25 -35.47 ;
      RECT 24.65 -32.36 25 -32.24 ;
      RECT 24.65 -29.13 25 -29.01 ;
      RECT 24.65 -25.9 25 -25.78 ;
      RECT 24.65 -22.67 25 -22.55 ;
      RECT 24.65 -19.44 25 -19.32 ;
      RECT 24.65 -16.21 25 -16.09 ;
      RECT 24.65 -12.98 25 -12.86 ;
      RECT 24.65 -9.75 25 -9.63 ;
      RECT 24.65 -6.52 25 -6.4 ;
      RECT 24.65 -3.29 25 -3.17 ;
      RECT 24.65 -0.06 25 0.06 ;
      RECT 24.765 -108.175 24.865 -107.215 ;
      RECT 24.765 2.175 24.865 3.135 ;
      RECT 24.665 -113.555 24.765 -113.085 ;
      RECT 24.165 -100.19 24.515 -100.07 ;
      RECT 24.165 -96.96 24.515 -96.84 ;
      RECT 24.165 -93.73 24.515 -93.61 ;
      RECT 24.165 -90.5 24.515 -90.38 ;
      RECT 24.165 -87.27 24.515 -87.15 ;
      RECT 24.165 -84.04 24.515 -83.92 ;
      RECT 24.165 -80.81 24.515 -80.69 ;
      RECT 24.165 -77.58 24.515 -77.46 ;
      RECT 24.165 -74.35 24.515 -74.23 ;
      RECT 24.165 -71.12 24.515 -71 ;
      RECT 24.165 -67.89 24.515 -67.77 ;
      RECT 24.165 -64.66 24.515 -64.54 ;
      RECT 24.165 -61.43 24.515 -61.31 ;
      RECT 24.165 -58.2 24.515 -58.08 ;
      RECT 24.165 -54.97 24.515 -54.85 ;
      RECT 24.165 -51.74 24.515 -51.62 ;
      RECT 24.165 -48.51 24.515 -48.39 ;
      RECT 24.165 -45.28 24.515 -45.16 ;
      RECT 24.165 -42.05 24.515 -41.93 ;
      RECT 24.165 -38.82 24.515 -38.7 ;
      RECT 24.165 -35.59 24.515 -35.47 ;
      RECT 24.165 -32.36 24.515 -32.24 ;
      RECT 24.165 -29.13 24.515 -29.01 ;
      RECT 24.165 -25.9 24.515 -25.78 ;
      RECT 24.165 -22.67 24.515 -22.55 ;
      RECT 24.165 -19.44 24.515 -19.32 ;
      RECT 24.165 -16.21 24.515 -16.09 ;
      RECT 24.165 -12.98 24.515 -12.86 ;
      RECT 24.165 -9.75 24.515 -9.63 ;
      RECT 24.165 -6.52 24.515 -6.4 ;
      RECT 24.165 -3.29 24.515 -3.17 ;
      RECT 24.165 -0.06 24.515 0.06 ;
      RECT 24.3 -110.735 24.45 -110.445 ;
      RECT 24.335 -108.175 24.435 -107.215 ;
      RECT 24.335 2.175 24.435 3.135 ;
      RECT 24.315 -112.19 24.415 -111.65 ;
      RECT 24.075 -113.555 24.175 -113.085 ;
      RECT 24.075 -108.175 24.175 -107.215 ;
      RECT 23.95 -101.06 24.05 -100.525 ;
      RECT 23.95 -99.735 24.05 -99.2 ;
      RECT 23.95 -97.83 24.05 -97.295 ;
      RECT 23.95 -96.505 24.05 -95.97 ;
      RECT 23.95 -94.6 24.05 -94.065 ;
      RECT 23.95 -93.275 24.05 -92.74 ;
      RECT 23.95 -91.37 24.05 -90.835 ;
      RECT 23.95 -90.045 24.05 -89.51 ;
      RECT 23.95 -88.14 24.05 -87.605 ;
      RECT 23.95 -86.815 24.05 -86.28 ;
      RECT 23.95 -84.91 24.05 -84.375 ;
      RECT 23.95 -83.585 24.05 -83.05 ;
      RECT 23.95 -81.68 24.05 -81.145 ;
      RECT 23.95 -80.355 24.05 -79.82 ;
      RECT 23.95 -78.45 24.05 -77.915 ;
      RECT 23.95 -77.125 24.05 -76.59 ;
      RECT 23.95 -75.22 24.05 -74.685 ;
      RECT 23.95 -73.895 24.05 -73.36 ;
      RECT 23.95 -71.99 24.05 -71.455 ;
      RECT 23.95 -70.665 24.05 -70.13 ;
      RECT 23.95 -68.76 24.05 -68.225 ;
      RECT 23.95 -67.435 24.05 -66.9 ;
      RECT 23.95 -65.53 24.05 -64.995 ;
      RECT 23.95 -64.205 24.05 -63.67 ;
      RECT 23.95 -62.3 24.05 -61.765 ;
      RECT 23.95 -60.975 24.05 -60.44 ;
      RECT 23.95 -59.07 24.05 -58.535 ;
      RECT 23.95 -57.745 24.05 -57.21 ;
      RECT 23.95 -55.84 24.05 -55.305 ;
      RECT 23.95 -54.515 24.05 -53.98 ;
      RECT 23.95 -52.61 24.05 -52.075 ;
      RECT 23.95 -51.285 24.05 -50.75 ;
      RECT 23.95 -49.38 24.05 -48.845 ;
      RECT 23.95 -48.055 24.05 -47.52 ;
      RECT 23.95 -46.15 24.05 -45.615 ;
      RECT 23.95 -44.825 24.05 -44.29 ;
      RECT 23.95 -42.92 24.05 -42.385 ;
      RECT 23.95 -41.595 24.05 -41.06 ;
      RECT 23.95 -39.69 24.05 -39.155 ;
      RECT 23.95 -38.365 24.05 -37.83 ;
      RECT 23.95 -36.46 24.05 -35.925 ;
      RECT 23.95 -35.135 24.05 -34.6 ;
      RECT 23.95 -33.23 24.05 -32.695 ;
      RECT 23.95 -31.905 24.05 -31.37 ;
      RECT 23.95 -30 24.05 -29.465 ;
      RECT 23.95 -28.675 24.05 -28.14 ;
      RECT 23.95 -26.77 24.05 -26.235 ;
      RECT 23.95 -25.445 24.05 -24.91 ;
      RECT 23.95 -23.54 24.05 -23.005 ;
      RECT 23.95 -22.215 24.05 -21.68 ;
      RECT 23.95 -20.31 24.05 -19.775 ;
      RECT 23.95 -18.985 24.05 -18.45 ;
      RECT 23.95 -17.08 24.05 -16.545 ;
      RECT 23.95 -15.755 24.05 -15.22 ;
      RECT 23.95 -13.85 24.05 -13.315 ;
      RECT 23.95 -12.525 24.05 -11.99 ;
      RECT 23.95 -10.62 24.05 -10.085 ;
      RECT 23.95 -9.295 24.05 -8.76 ;
      RECT 23.95 -7.39 24.05 -6.855 ;
      RECT 23.95 -6.065 24.05 -5.53 ;
      RECT 23.95 -4.16 24.05 -3.625 ;
      RECT 23.95 -2.835 24.05 -2.3 ;
      RECT 23.95 -0.93 24.05 -0.395 ;
      RECT 23.95 0.395 24.05 0.93 ;
      RECT 23.825 -104.945 23.925 -103.985 ;
      RECT 23.45 -100.19 23.8 -100.07 ;
      RECT 23.45 -96.96 23.8 -96.84 ;
      RECT 23.45 -93.73 23.8 -93.61 ;
      RECT 23.45 -90.5 23.8 -90.38 ;
      RECT 23.45 -87.27 23.8 -87.15 ;
      RECT 23.45 -84.04 23.8 -83.92 ;
      RECT 23.45 -80.81 23.8 -80.69 ;
      RECT 23.45 -77.58 23.8 -77.46 ;
      RECT 23.45 -74.35 23.8 -74.23 ;
      RECT 23.45 -71.12 23.8 -71 ;
      RECT 23.45 -67.89 23.8 -67.77 ;
      RECT 23.45 -64.66 23.8 -64.54 ;
      RECT 23.45 -61.43 23.8 -61.31 ;
      RECT 23.45 -58.2 23.8 -58.08 ;
      RECT 23.45 -54.97 23.8 -54.85 ;
      RECT 23.45 -51.74 23.8 -51.62 ;
      RECT 23.45 -48.51 23.8 -48.39 ;
      RECT 23.45 -45.28 23.8 -45.16 ;
      RECT 23.45 -42.05 23.8 -41.93 ;
      RECT 23.45 -38.82 23.8 -38.7 ;
      RECT 23.45 -35.59 23.8 -35.47 ;
      RECT 23.45 -32.36 23.8 -32.24 ;
      RECT 23.45 -29.13 23.8 -29.01 ;
      RECT 23.45 -25.9 23.8 -25.78 ;
      RECT 23.45 -22.67 23.8 -22.55 ;
      RECT 23.45 -19.44 23.8 -19.32 ;
      RECT 23.45 -16.21 23.8 -16.09 ;
      RECT 23.45 -12.98 23.8 -12.86 ;
      RECT 23.45 -9.75 23.8 -9.63 ;
      RECT 23.45 -6.52 23.8 -6.4 ;
      RECT 23.45 -3.29 23.8 -3.17 ;
      RECT 23.45 -0.06 23.8 0.06 ;
      RECT 23.565 -104.945 23.665 -103.985 ;
      RECT 23.565 2.175 23.665 3.135 ;
      RECT 23.275 -112.255 23.375 -111.775 ;
      RECT 23.275 -110.765 23.375 -110.295 ;
      RECT 22.965 -100.19 23.315 -100.07 ;
      RECT 22.965 -96.96 23.315 -96.84 ;
      RECT 22.965 -93.73 23.315 -93.61 ;
      RECT 22.965 -90.5 23.315 -90.38 ;
      RECT 22.965 -87.27 23.315 -87.15 ;
      RECT 22.965 -84.04 23.315 -83.92 ;
      RECT 22.965 -80.81 23.315 -80.69 ;
      RECT 22.965 -77.58 23.315 -77.46 ;
      RECT 22.965 -74.35 23.315 -74.23 ;
      RECT 22.965 -71.12 23.315 -71 ;
      RECT 22.965 -67.89 23.315 -67.77 ;
      RECT 22.965 -64.66 23.315 -64.54 ;
      RECT 22.965 -61.43 23.315 -61.31 ;
      RECT 22.965 -58.2 23.315 -58.08 ;
      RECT 22.965 -54.97 23.315 -54.85 ;
      RECT 22.965 -51.74 23.315 -51.62 ;
      RECT 22.965 -48.51 23.315 -48.39 ;
      RECT 22.965 -45.28 23.315 -45.16 ;
      RECT 22.965 -42.05 23.315 -41.93 ;
      RECT 22.965 -38.82 23.315 -38.7 ;
      RECT 22.965 -35.59 23.315 -35.47 ;
      RECT 22.965 -32.36 23.315 -32.24 ;
      RECT 22.965 -29.13 23.315 -29.01 ;
      RECT 22.965 -25.9 23.315 -25.78 ;
      RECT 22.965 -22.67 23.315 -22.55 ;
      RECT 22.965 -19.44 23.315 -19.32 ;
      RECT 22.965 -16.21 23.315 -16.09 ;
      RECT 22.965 -12.98 23.315 -12.86 ;
      RECT 22.965 -9.75 23.315 -9.63 ;
      RECT 22.965 -6.52 23.315 -6.4 ;
      RECT 22.965 -3.29 23.315 -3.17 ;
      RECT 22.965 -0.06 23.315 0.06 ;
      RECT 23.135 -104.945 23.235 -103.985 ;
      RECT 23.135 2.175 23.235 3.135 ;
      RECT 19.235 -108.655 23.015 -108.535 ;
      RECT 22.875 -104.945 22.975 -103.985 ;
      RECT 22.75 -101.06 22.85 -100.525 ;
      RECT 22.75 -99.735 22.85 -99.2 ;
      RECT 22.75 -97.83 22.85 -97.295 ;
      RECT 22.75 -96.505 22.85 -95.97 ;
      RECT 22.75 -94.6 22.85 -94.065 ;
      RECT 22.75 -93.275 22.85 -92.74 ;
      RECT 22.75 -91.37 22.85 -90.835 ;
      RECT 22.75 -90.045 22.85 -89.51 ;
      RECT 22.75 -88.14 22.85 -87.605 ;
      RECT 22.75 -86.815 22.85 -86.28 ;
      RECT 22.75 -84.91 22.85 -84.375 ;
      RECT 22.75 -83.585 22.85 -83.05 ;
      RECT 22.75 -81.68 22.85 -81.145 ;
      RECT 22.75 -80.355 22.85 -79.82 ;
      RECT 22.75 -78.45 22.85 -77.915 ;
      RECT 22.75 -77.125 22.85 -76.59 ;
      RECT 22.75 -75.22 22.85 -74.685 ;
      RECT 22.75 -73.895 22.85 -73.36 ;
      RECT 22.75 -71.99 22.85 -71.455 ;
      RECT 22.75 -70.665 22.85 -70.13 ;
      RECT 22.75 -68.76 22.85 -68.225 ;
      RECT 22.75 -67.435 22.85 -66.9 ;
      RECT 22.75 -65.53 22.85 -64.995 ;
      RECT 22.75 -64.205 22.85 -63.67 ;
      RECT 22.75 -62.3 22.85 -61.765 ;
      RECT 22.75 -60.975 22.85 -60.44 ;
      RECT 22.75 -59.07 22.85 -58.535 ;
      RECT 22.75 -57.745 22.85 -57.21 ;
      RECT 22.75 -55.84 22.85 -55.305 ;
      RECT 22.75 -54.515 22.85 -53.98 ;
      RECT 22.75 -52.61 22.85 -52.075 ;
      RECT 22.75 -51.285 22.85 -50.75 ;
      RECT 22.75 -49.38 22.85 -48.845 ;
      RECT 22.75 -48.055 22.85 -47.52 ;
      RECT 22.75 -46.15 22.85 -45.615 ;
      RECT 22.75 -44.825 22.85 -44.29 ;
      RECT 22.75 -42.92 22.85 -42.385 ;
      RECT 22.75 -41.595 22.85 -41.06 ;
      RECT 22.75 -39.69 22.85 -39.155 ;
      RECT 22.75 -38.365 22.85 -37.83 ;
      RECT 22.75 -36.46 22.85 -35.925 ;
      RECT 22.75 -35.135 22.85 -34.6 ;
      RECT 22.75 -33.23 22.85 -32.695 ;
      RECT 22.75 -31.905 22.85 -31.37 ;
      RECT 22.75 -30 22.85 -29.465 ;
      RECT 22.75 -28.675 22.85 -28.14 ;
      RECT 22.75 -26.77 22.85 -26.235 ;
      RECT 22.75 -25.445 22.85 -24.91 ;
      RECT 22.75 -23.54 22.85 -23.005 ;
      RECT 22.75 -22.215 22.85 -21.68 ;
      RECT 22.75 -20.31 22.85 -19.775 ;
      RECT 22.75 -18.985 22.85 -18.45 ;
      RECT 22.75 -17.08 22.85 -16.545 ;
      RECT 22.75 -15.755 22.85 -15.22 ;
      RECT 22.75 -13.85 22.85 -13.315 ;
      RECT 22.75 -12.525 22.85 -11.99 ;
      RECT 22.75 -10.62 22.85 -10.085 ;
      RECT 22.75 -9.295 22.85 -8.76 ;
      RECT 22.75 -7.39 22.85 -6.855 ;
      RECT 22.75 -6.065 22.85 -5.53 ;
      RECT 22.75 -4.16 22.85 -3.625 ;
      RECT 22.75 -2.835 22.85 -2.3 ;
      RECT 22.75 -0.93 22.85 -0.395 ;
      RECT 22.75 0.395 22.85 0.93 ;
      RECT 22.685 -110.75 22.805 -110.37 ;
      RECT 22.685 -112.245 22.785 -111.775 ;
      RECT 22.625 -104.945 22.725 -103.985 ;
      RECT 22.25 -100.19 22.6 -100.07 ;
      RECT 22.25 -96.96 22.6 -96.84 ;
      RECT 22.25 -93.73 22.6 -93.61 ;
      RECT 22.25 -90.5 22.6 -90.38 ;
      RECT 22.25 -87.27 22.6 -87.15 ;
      RECT 22.25 -84.04 22.6 -83.92 ;
      RECT 22.25 -80.81 22.6 -80.69 ;
      RECT 22.25 -77.58 22.6 -77.46 ;
      RECT 22.25 -74.35 22.6 -74.23 ;
      RECT 22.25 -71.12 22.6 -71 ;
      RECT 22.25 -67.89 22.6 -67.77 ;
      RECT 22.25 -64.66 22.6 -64.54 ;
      RECT 22.25 -61.43 22.6 -61.31 ;
      RECT 22.25 -58.2 22.6 -58.08 ;
      RECT 22.25 -54.97 22.6 -54.85 ;
      RECT 22.25 -51.74 22.6 -51.62 ;
      RECT 22.25 -48.51 22.6 -48.39 ;
      RECT 22.25 -45.28 22.6 -45.16 ;
      RECT 22.25 -42.05 22.6 -41.93 ;
      RECT 22.25 -38.82 22.6 -38.7 ;
      RECT 22.25 -35.59 22.6 -35.47 ;
      RECT 22.25 -32.36 22.6 -32.24 ;
      RECT 22.25 -29.13 22.6 -29.01 ;
      RECT 22.25 -25.9 22.6 -25.78 ;
      RECT 22.25 -22.67 22.6 -22.55 ;
      RECT 22.25 -19.44 22.6 -19.32 ;
      RECT 22.25 -16.21 22.6 -16.09 ;
      RECT 22.25 -12.98 22.6 -12.86 ;
      RECT 22.25 -9.75 22.6 -9.63 ;
      RECT 22.25 -6.52 22.6 -6.4 ;
      RECT 22.25 -3.29 22.6 -3.17 ;
      RECT 22.25 -0.06 22.6 0.06 ;
      RECT 22.365 -104.945 22.465 -103.985 ;
      RECT 22.365 2.175 22.465 3.135 ;
      RECT 22.095 -109.595 22.23 -109.275 ;
      RECT 21.765 -100.19 22.115 -100.07 ;
      RECT 21.765 -96.96 22.115 -96.84 ;
      RECT 21.765 -93.73 22.115 -93.61 ;
      RECT 21.765 -90.5 22.115 -90.38 ;
      RECT 21.765 -87.27 22.115 -87.15 ;
      RECT 21.765 -84.04 22.115 -83.92 ;
      RECT 21.765 -80.81 22.115 -80.69 ;
      RECT 21.765 -77.58 22.115 -77.46 ;
      RECT 21.765 -74.35 22.115 -74.23 ;
      RECT 21.765 -71.12 22.115 -71 ;
      RECT 21.765 -67.89 22.115 -67.77 ;
      RECT 21.765 -64.66 22.115 -64.54 ;
      RECT 21.765 -61.43 22.115 -61.31 ;
      RECT 21.765 -58.2 22.115 -58.08 ;
      RECT 21.765 -54.97 22.115 -54.85 ;
      RECT 21.765 -51.74 22.115 -51.62 ;
      RECT 21.765 -48.51 22.115 -48.39 ;
      RECT 21.765 -45.28 22.115 -45.16 ;
      RECT 21.765 -42.05 22.115 -41.93 ;
      RECT 21.765 -38.82 22.115 -38.7 ;
      RECT 21.765 -35.59 22.115 -35.47 ;
      RECT 21.765 -32.36 22.115 -32.24 ;
      RECT 21.765 -29.13 22.115 -29.01 ;
      RECT 21.765 -25.9 22.115 -25.78 ;
      RECT 21.765 -22.67 22.115 -22.55 ;
      RECT 21.765 -19.44 22.115 -19.32 ;
      RECT 21.765 -16.21 22.115 -16.09 ;
      RECT 21.765 -12.98 22.115 -12.86 ;
      RECT 21.765 -9.75 22.115 -9.63 ;
      RECT 21.765 -6.52 22.115 -6.4 ;
      RECT 21.765 -3.29 22.115 -3.17 ;
      RECT 21.765 -0.06 22.115 0.06 ;
      RECT 21.935 -104.945 22.035 -103.985 ;
      RECT 21.935 2.175 22.035 3.135 ;
      RECT 21.76 -109.595 21.905 -109.275 ;
      RECT 21.675 -104.945 21.775 -103.985 ;
      RECT 21.55 -101.06 21.65 -100.525 ;
      RECT 21.55 -99.735 21.65 -99.2 ;
      RECT 21.55 -97.83 21.65 -97.295 ;
      RECT 21.55 -96.505 21.65 -95.97 ;
      RECT 21.55 -94.6 21.65 -94.065 ;
      RECT 21.55 -93.275 21.65 -92.74 ;
      RECT 21.55 -91.37 21.65 -90.835 ;
      RECT 21.55 -90.045 21.65 -89.51 ;
      RECT 21.55 -88.14 21.65 -87.605 ;
      RECT 21.55 -86.815 21.65 -86.28 ;
      RECT 21.55 -84.91 21.65 -84.375 ;
      RECT 21.55 -83.585 21.65 -83.05 ;
      RECT 21.55 -81.68 21.65 -81.145 ;
      RECT 21.55 -80.355 21.65 -79.82 ;
      RECT 21.55 -78.45 21.65 -77.915 ;
      RECT 21.55 -77.125 21.65 -76.59 ;
      RECT 21.55 -75.22 21.65 -74.685 ;
      RECT 21.55 -73.895 21.65 -73.36 ;
      RECT 21.55 -71.99 21.65 -71.455 ;
      RECT 21.55 -70.665 21.65 -70.13 ;
      RECT 21.55 -68.76 21.65 -68.225 ;
      RECT 21.55 -67.435 21.65 -66.9 ;
      RECT 21.55 -65.53 21.65 -64.995 ;
      RECT 21.55 -64.205 21.65 -63.67 ;
      RECT 21.55 -62.3 21.65 -61.765 ;
      RECT 21.55 -60.975 21.65 -60.44 ;
      RECT 21.55 -59.07 21.65 -58.535 ;
      RECT 21.55 -57.745 21.65 -57.21 ;
      RECT 21.55 -55.84 21.65 -55.305 ;
      RECT 21.55 -54.515 21.65 -53.98 ;
      RECT 21.55 -52.61 21.65 -52.075 ;
      RECT 21.55 -51.285 21.65 -50.75 ;
      RECT 21.55 -49.38 21.65 -48.845 ;
      RECT 21.55 -48.055 21.65 -47.52 ;
      RECT 21.55 -46.15 21.65 -45.615 ;
      RECT 21.55 -44.825 21.65 -44.29 ;
      RECT 21.55 -42.92 21.65 -42.385 ;
      RECT 21.55 -41.595 21.65 -41.06 ;
      RECT 21.55 -39.69 21.65 -39.155 ;
      RECT 21.55 -38.365 21.65 -37.83 ;
      RECT 21.55 -36.46 21.65 -35.925 ;
      RECT 21.55 -35.135 21.65 -34.6 ;
      RECT 21.55 -33.23 21.65 -32.695 ;
      RECT 21.55 -31.905 21.65 -31.37 ;
      RECT 21.55 -30 21.65 -29.465 ;
      RECT 21.55 -28.675 21.65 -28.14 ;
      RECT 21.55 -26.77 21.65 -26.235 ;
      RECT 21.55 -25.445 21.65 -24.91 ;
      RECT 21.55 -23.54 21.65 -23.005 ;
      RECT 21.55 -22.215 21.65 -21.68 ;
      RECT 21.55 -20.31 21.65 -19.775 ;
      RECT 21.55 -18.985 21.65 -18.45 ;
      RECT 21.55 -17.08 21.65 -16.545 ;
      RECT 21.55 -15.755 21.65 -15.22 ;
      RECT 21.55 -13.85 21.65 -13.315 ;
      RECT 21.55 -12.525 21.65 -11.99 ;
      RECT 21.55 -10.62 21.65 -10.085 ;
      RECT 21.55 -9.295 21.65 -8.76 ;
      RECT 21.55 -7.39 21.65 -6.855 ;
      RECT 21.55 -6.065 21.65 -5.53 ;
      RECT 21.55 -4.16 21.65 -3.625 ;
      RECT 21.55 -2.835 21.65 -2.3 ;
      RECT 21.55 -0.93 21.65 -0.395 ;
      RECT 21.55 0.395 21.65 0.93 ;
      RECT 21.425 -108.175 21.525 -107.215 ;
      RECT 21.05 -100.19 21.4 -100.07 ;
      RECT 21.05 -96.96 21.4 -96.84 ;
      RECT 21.05 -93.73 21.4 -93.61 ;
      RECT 21.05 -90.5 21.4 -90.38 ;
      RECT 21.05 -87.27 21.4 -87.15 ;
      RECT 21.05 -84.04 21.4 -83.92 ;
      RECT 21.05 -80.81 21.4 -80.69 ;
      RECT 21.05 -77.58 21.4 -77.46 ;
      RECT 21.05 -74.35 21.4 -74.23 ;
      RECT 21.05 -71.12 21.4 -71 ;
      RECT 21.05 -67.89 21.4 -67.77 ;
      RECT 21.05 -64.66 21.4 -64.54 ;
      RECT 21.05 -61.43 21.4 -61.31 ;
      RECT 21.05 -58.2 21.4 -58.08 ;
      RECT 21.05 -54.97 21.4 -54.85 ;
      RECT 21.05 -51.74 21.4 -51.62 ;
      RECT 21.05 -48.51 21.4 -48.39 ;
      RECT 21.05 -45.28 21.4 -45.16 ;
      RECT 21.05 -42.05 21.4 -41.93 ;
      RECT 21.05 -38.82 21.4 -38.7 ;
      RECT 21.05 -35.59 21.4 -35.47 ;
      RECT 21.05 -32.36 21.4 -32.24 ;
      RECT 21.05 -29.13 21.4 -29.01 ;
      RECT 21.05 -25.9 21.4 -25.78 ;
      RECT 21.05 -22.67 21.4 -22.55 ;
      RECT 21.05 -19.44 21.4 -19.32 ;
      RECT 21.05 -16.21 21.4 -16.09 ;
      RECT 21.05 -12.98 21.4 -12.86 ;
      RECT 21.05 -9.75 21.4 -9.63 ;
      RECT 21.05 -6.52 21.4 -6.4 ;
      RECT 21.05 -3.29 21.4 -3.17 ;
      RECT 21.05 -0.06 21.4 0.06 ;
      RECT 21.255 -112.255 21.355 -111.775 ;
      RECT 21.255 -110.765 21.355 -110.295 ;
      RECT 21.165 -108.175 21.265 -107.215 ;
      RECT 21.165 2.175 21.265 3.135 ;
      RECT 20.565 -100.19 20.915 -100.07 ;
      RECT 20.565 -96.96 20.915 -96.84 ;
      RECT 20.565 -93.73 20.915 -93.61 ;
      RECT 20.565 -90.5 20.915 -90.38 ;
      RECT 20.565 -87.27 20.915 -87.15 ;
      RECT 20.565 -84.04 20.915 -83.92 ;
      RECT 20.565 -80.81 20.915 -80.69 ;
      RECT 20.565 -77.58 20.915 -77.46 ;
      RECT 20.565 -74.35 20.915 -74.23 ;
      RECT 20.565 -71.12 20.915 -71 ;
      RECT 20.565 -67.89 20.915 -67.77 ;
      RECT 20.565 -64.66 20.915 -64.54 ;
      RECT 20.565 -61.43 20.915 -61.31 ;
      RECT 20.565 -58.2 20.915 -58.08 ;
      RECT 20.565 -54.97 20.915 -54.85 ;
      RECT 20.565 -51.74 20.915 -51.62 ;
      RECT 20.565 -48.51 20.915 -48.39 ;
      RECT 20.565 -45.28 20.915 -45.16 ;
      RECT 20.565 -42.05 20.915 -41.93 ;
      RECT 20.565 -38.82 20.915 -38.7 ;
      RECT 20.565 -35.59 20.915 -35.47 ;
      RECT 20.565 -32.36 20.915 -32.24 ;
      RECT 20.565 -29.13 20.915 -29.01 ;
      RECT 20.565 -25.9 20.915 -25.78 ;
      RECT 20.565 -22.67 20.915 -22.55 ;
      RECT 20.565 -19.44 20.915 -19.32 ;
      RECT 20.565 -16.21 20.915 -16.09 ;
      RECT 20.565 -12.98 20.915 -12.86 ;
      RECT 20.565 -9.75 20.915 -9.63 ;
      RECT 20.565 -6.52 20.915 -6.4 ;
      RECT 20.565 -3.29 20.915 -3.17 ;
      RECT 20.565 -0.06 20.915 0.06 ;
      RECT 20.735 -108.175 20.835 -107.215 ;
      RECT 20.735 2.175 20.835 3.135 ;
      RECT 20.63 -110.765 20.8 -110.385 ;
      RECT 20.665 -112.245 20.765 -111.775 ;
      RECT 20.475 -108.175 20.575 -107.215 ;
      RECT 20.35 -101.06 20.45 -100.525 ;
      RECT 20.35 -99.735 20.45 -99.2 ;
      RECT 20.35 -97.83 20.45 -97.295 ;
      RECT 20.35 -96.505 20.45 -95.97 ;
      RECT 20.35 -94.6 20.45 -94.065 ;
      RECT 20.35 -93.275 20.45 -92.74 ;
      RECT 20.35 -91.37 20.45 -90.835 ;
      RECT 20.35 -90.045 20.45 -89.51 ;
      RECT 20.35 -88.14 20.45 -87.605 ;
      RECT 20.35 -86.815 20.45 -86.28 ;
      RECT 20.35 -84.91 20.45 -84.375 ;
      RECT 20.35 -83.585 20.45 -83.05 ;
      RECT 20.35 -81.68 20.45 -81.145 ;
      RECT 20.35 -80.355 20.45 -79.82 ;
      RECT 20.35 -78.45 20.45 -77.915 ;
      RECT 20.35 -77.125 20.45 -76.59 ;
      RECT 20.35 -75.22 20.45 -74.685 ;
      RECT 20.35 -73.895 20.45 -73.36 ;
      RECT 20.35 -71.99 20.45 -71.455 ;
      RECT 20.35 -70.665 20.45 -70.13 ;
      RECT 20.35 -68.76 20.45 -68.225 ;
      RECT 20.35 -67.435 20.45 -66.9 ;
      RECT 20.35 -65.53 20.45 -64.995 ;
      RECT 20.35 -64.205 20.45 -63.67 ;
      RECT 20.35 -62.3 20.45 -61.765 ;
      RECT 20.35 -60.975 20.45 -60.44 ;
      RECT 20.35 -59.07 20.45 -58.535 ;
      RECT 20.35 -57.745 20.45 -57.21 ;
      RECT 20.35 -55.84 20.45 -55.305 ;
      RECT 20.35 -54.515 20.45 -53.98 ;
      RECT 20.35 -52.61 20.45 -52.075 ;
      RECT 20.35 -51.285 20.45 -50.75 ;
      RECT 20.35 -49.38 20.45 -48.845 ;
      RECT 20.35 -48.055 20.45 -47.52 ;
      RECT 20.35 -46.15 20.45 -45.615 ;
      RECT 20.35 -44.825 20.45 -44.29 ;
      RECT 20.35 -42.92 20.45 -42.385 ;
      RECT 20.35 -41.595 20.45 -41.06 ;
      RECT 20.35 -39.69 20.45 -39.155 ;
      RECT 20.35 -38.365 20.45 -37.83 ;
      RECT 20.35 -36.46 20.45 -35.925 ;
      RECT 20.35 -35.135 20.45 -34.6 ;
      RECT 20.35 -33.23 20.45 -32.695 ;
      RECT 20.35 -31.905 20.45 -31.37 ;
      RECT 20.35 -30 20.45 -29.465 ;
      RECT 20.35 -28.675 20.45 -28.14 ;
      RECT 20.35 -26.77 20.45 -26.235 ;
      RECT 20.35 -25.445 20.45 -24.91 ;
      RECT 20.35 -23.54 20.45 -23.005 ;
      RECT 20.35 -22.215 20.45 -21.68 ;
      RECT 20.35 -20.31 20.45 -19.775 ;
      RECT 20.35 -18.985 20.45 -18.45 ;
      RECT 20.35 -17.08 20.45 -16.545 ;
      RECT 20.35 -15.755 20.45 -15.22 ;
      RECT 20.35 -13.85 20.45 -13.315 ;
      RECT 20.35 -12.525 20.45 -11.99 ;
      RECT 20.35 -10.62 20.45 -10.085 ;
      RECT 20.35 -9.295 20.45 -8.76 ;
      RECT 20.35 -7.39 20.45 -6.855 ;
      RECT 20.35 -6.065 20.45 -5.53 ;
      RECT 20.35 -4.16 20.45 -3.625 ;
      RECT 20.35 -2.835 20.45 -2.3 ;
      RECT 20.35 -0.93 20.45 -0.395 ;
      RECT 20.35 0.395 20.45 0.93 ;
      RECT 20.225 -108.175 20.325 -107.215 ;
      RECT 19.85 -100.19 20.2 -100.07 ;
      RECT 19.85 -96.96 20.2 -96.84 ;
      RECT 19.85 -93.73 20.2 -93.61 ;
      RECT 19.85 -90.5 20.2 -90.38 ;
      RECT 19.85 -87.27 20.2 -87.15 ;
      RECT 19.85 -84.04 20.2 -83.92 ;
      RECT 19.85 -80.81 20.2 -80.69 ;
      RECT 19.85 -77.58 20.2 -77.46 ;
      RECT 19.85 -74.35 20.2 -74.23 ;
      RECT 19.85 -71.12 20.2 -71 ;
      RECT 19.85 -67.89 20.2 -67.77 ;
      RECT 19.85 -64.66 20.2 -64.54 ;
      RECT 19.85 -61.43 20.2 -61.31 ;
      RECT 19.85 -58.2 20.2 -58.08 ;
      RECT 19.85 -54.97 20.2 -54.85 ;
      RECT 19.85 -51.74 20.2 -51.62 ;
      RECT 19.85 -48.51 20.2 -48.39 ;
      RECT 19.85 -45.28 20.2 -45.16 ;
      RECT 19.85 -42.05 20.2 -41.93 ;
      RECT 19.85 -38.82 20.2 -38.7 ;
      RECT 19.85 -35.59 20.2 -35.47 ;
      RECT 19.85 -32.36 20.2 -32.24 ;
      RECT 19.85 -29.13 20.2 -29.01 ;
      RECT 19.85 -25.9 20.2 -25.78 ;
      RECT 19.85 -22.67 20.2 -22.55 ;
      RECT 19.85 -19.44 20.2 -19.32 ;
      RECT 19.85 -16.21 20.2 -16.09 ;
      RECT 19.85 -12.98 20.2 -12.86 ;
      RECT 19.85 -9.75 20.2 -9.63 ;
      RECT 19.85 -6.52 20.2 -6.4 ;
      RECT 19.85 -3.29 20.2 -3.17 ;
      RECT 19.85 -0.06 20.2 0.06 ;
      RECT 19.965 -108.175 20.065 -107.215 ;
      RECT 19.965 2.175 20.065 3.135 ;
      RECT 19.865 -113.555 19.965 -113.085 ;
      RECT 19.365 -100.19 19.715 -100.07 ;
      RECT 19.365 -96.96 19.715 -96.84 ;
      RECT 19.365 -93.73 19.715 -93.61 ;
      RECT 19.365 -90.5 19.715 -90.38 ;
      RECT 19.365 -87.27 19.715 -87.15 ;
      RECT 19.365 -84.04 19.715 -83.92 ;
      RECT 19.365 -80.81 19.715 -80.69 ;
      RECT 19.365 -77.58 19.715 -77.46 ;
      RECT 19.365 -74.35 19.715 -74.23 ;
      RECT 19.365 -71.12 19.715 -71 ;
      RECT 19.365 -67.89 19.715 -67.77 ;
      RECT 19.365 -64.66 19.715 -64.54 ;
      RECT 19.365 -61.43 19.715 -61.31 ;
      RECT 19.365 -58.2 19.715 -58.08 ;
      RECT 19.365 -54.97 19.715 -54.85 ;
      RECT 19.365 -51.74 19.715 -51.62 ;
      RECT 19.365 -48.51 19.715 -48.39 ;
      RECT 19.365 -45.28 19.715 -45.16 ;
      RECT 19.365 -42.05 19.715 -41.93 ;
      RECT 19.365 -38.82 19.715 -38.7 ;
      RECT 19.365 -35.59 19.715 -35.47 ;
      RECT 19.365 -32.36 19.715 -32.24 ;
      RECT 19.365 -29.13 19.715 -29.01 ;
      RECT 19.365 -25.9 19.715 -25.78 ;
      RECT 19.365 -22.67 19.715 -22.55 ;
      RECT 19.365 -19.44 19.715 -19.32 ;
      RECT 19.365 -16.21 19.715 -16.09 ;
      RECT 19.365 -12.98 19.715 -12.86 ;
      RECT 19.365 -9.75 19.715 -9.63 ;
      RECT 19.365 -6.52 19.715 -6.4 ;
      RECT 19.365 -3.29 19.715 -3.17 ;
      RECT 19.365 -0.06 19.715 0.06 ;
      RECT 19.5 -110.735 19.65 -110.445 ;
      RECT 19.535 -108.175 19.635 -107.215 ;
      RECT 19.535 2.175 19.635 3.135 ;
      RECT 19.515 -112.19 19.615 -111.65 ;
      RECT 19.275 -113.555 19.375 -113.085 ;
      RECT 19.275 -108.175 19.375 -107.215 ;
      RECT 19.15 -101.06 19.25 -100.525 ;
      RECT 19.15 -99.735 19.25 -99.2 ;
      RECT 19.15 -97.83 19.25 -97.295 ;
      RECT 19.15 -96.505 19.25 -95.97 ;
      RECT 19.15 -94.6 19.25 -94.065 ;
      RECT 19.15 -93.275 19.25 -92.74 ;
      RECT 19.15 -91.37 19.25 -90.835 ;
      RECT 19.15 -90.045 19.25 -89.51 ;
      RECT 19.15 -88.14 19.25 -87.605 ;
      RECT 19.15 -86.815 19.25 -86.28 ;
      RECT 19.15 -84.91 19.25 -84.375 ;
      RECT 19.15 -83.585 19.25 -83.05 ;
      RECT 19.15 -81.68 19.25 -81.145 ;
      RECT 19.15 -80.355 19.25 -79.82 ;
      RECT 19.15 -78.45 19.25 -77.915 ;
      RECT 19.15 -77.125 19.25 -76.59 ;
      RECT 19.15 -75.22 19.25 -74.685 ;
      RECT 19.15 -73.895 19.25 -73.36 ;
      RECT 19.15 -71.99 19.25 -71.455 ;
      RECT 19.15 -70.665 19.25 -70.13 ;
      RECT 19.15 -68.76 19.25 -68.225 ;
      RECT 19.15 -67.435 19.25 -66.9 ;
      RECT 19.15 -65.53 19.25 -64.995 ;
      RECT 19.15 -64.205 19.25 -63.67 ;
      RECT 19.15 -62.3 19.25 -61.765 ;
      RECT 19.15 -60.975 19.25 -60.44 ;
      RECT 19.15 -59.07 19.25 -58.535 ;
      RECT 19.15 -57.745 19.25 -57.21 ;
      RECT 19.15 -55.84 19.25 -55.305 ;
      RECT 19.15 -54.515 19.25 -53.98 ;
      RECT 19.15 -52.61 19.25 -52.075 ;
      RECT 19.15 -51.285 19.25 -50.75 ;
      RECT 19.15 -49.38 19.25 -48.845 ;
      RECT 19.15 -48.055 19.25 -47.52 ;
      RECT 19.15 -46.15 19.25 -45.615 ;
      RECT 19.15 -44.825 19.25 -44.29 ;
      RECT 19.15 -42.92 19.25 -42.385 ;
      RECT 19.15 -41.595 19.25 -41.06 ;
      RECT 19.15 -39.69 19.25 -39.155 ;
      RECT 19.15 -38.365 19.25 -37.83 ;
      RECT 19.15 -36.46 19.25 -35.925 ;
      RECT 19.15 -35.135 19.25 -34.6 ;
      RECT 19.15 -33.23 19.25 -32.695 ;
      RECT 19.15 -31.905 19.25 -31.37 ;
      RECT 19.15 -30 19.25 -29.465 ;
      RECT 19.15 -28.675 19.25 -28.14 ;
      RECT 19.15 -26.77 19.25 -26.235 ;
      RECT 19.15 -25.445 19.25 -24.91 ;
      RECT 19.15 -23.54 19.25 -23.005 ;
      RECT 19.15 -22.215 19.25 -21.68 ;
      RECT 19.15 -20.31 19.25 -19.775 ;
      RECT 19.15 -18.985 19.25 -18.45 ;
      RECT 19.15 -17.08 19.25 -16.545 ;
      RECT 19.15 -15.755 19.25 -15.22 ;
      RECT 19.15 -13.85 19.25 -13.315 ;
      RECT 19.15 -12.525 19.25 -11.99 ;
      RECT 19.15 -10.62 19.25 -10.085 ;
      RECT 19.15 -9.295 19.25 -8.76 ;
      RECT 19.15 -7.39 19.25 -6.855 ;
      RECT 19.15 -6.065 19.25 -5.53 ;
      RECT 19.15 -4.16 19.25 -3.625 ;
      RECT 19.15 -2.835 19.25 -2.3 ;
      RECT 19.15 -0.93 19.25 -0.395 ;
      RECT 19.15 0.395 19.25 0.93 ;
      RECT 19.025 -104.945 19.125 -103.985 ;
      RECT 18.65 -100.19 19 -100.07 ;
      RECT 18.65 -96.96 19 -96.84 ;
      RECT 18.65 -93.73 19 -93.61 ;
      RECT 18.65 -90.5 19 -90.38 ;
      RECT 18.65 -87.27 19 -87.15 ;
      RECT 18.65 -84.04 19 -83.92 ;
      RECT 18.65 -80.81 19 -80.69 ;
      RECT 18.65 -77.58 19 -77.46 ;
      RECT 18.65 -74.35 19 -74.23 ;
      RECT 18.65 -71.12 19 -71 ;
      RECT 18.65 -67.89 19 -67.77 ;
      RECT 18.65 -64.66 19 -64.54 ;
      RECT 18.65 -61.43 19 -61.31 ;
      RECT 18.65 -58.2 19 -58.08 ;
      RECT 18.65 -54.97 19 -54.85 ;
      RECT 18.65 -51.74 19 -51.62 ;
      RECT 18.65 -48.51 19 -48.39 ;
      RECT 18.65 -45.28 19 -45.16 ;
      RECT 18.65 -42.05 19 -41.93 ;
      RECT 18.65 -38.82 19 -38.7 ;
      RECT 18.65 -35.59 19 -35.47 ;
      RECT 18.65 -32.36 19 -32.24 ;
      RECT 18.65 -29.13 19 -29.01 ;
      RECT 18.65 -25.9 19 -25.78 ;
      RECT 18.65 -22.67 19 -22.55 ;
      RECT 18.65 -19.44 19 -19.32 ;
      RECT 18.65 -16.21 19 -16.09 ;
      RECT 18.65 -12.98 19 -12.86 ;
      RECT 18.65 -9.75 19 -9.63 ;
      RECT 18.65 -6.52 19 -6.4 ;
      RECT 18.65 -3.29 19 -3.17 ;
      RECT 18.65 -0.06 19 0.06 ;
      RECT 18.765 -104.945 18.865 -103.985 ;
      RECT 18.765 2.175 18.865 3.135 ;
      RECT 18.475 -112.255 18.575 -111.775 ;
      RECT 18.475 -110.765 18.575 -110.295 ;
      RECT 18.165 -100.19 18.515 -100.07 ;
      RECT 18.165 -96.96 18.515 -96.84 ;
      RECT 18.165 -93.73 18.515 -93.61 ;
      RECT 18.165 -90.5 18.515 -90.38 ;
      RECT 18.165 -87.27 18.515 -87.15 ;
      RECT 18.165 -84.04 18.515 -83.92 ;
      RECT 18.165 -80.81 18.515 -80.69 ;
      RECT 18.165 -77.58 18.515 -77.46 ;
      RECT 18.165 -74.35 18.515 -74.23 ;
      RECT 18.165 -71.12 18.515 -71 ;
      RECT 18.165 -67.89 18.515 -67.77 ;
      RECT 18.165 -64.66 18.515 -64.54 ;
      RECT 18.165 -61.43 18.515 -61.31 ;
      RECT 18.165 -58.2 18.515 -58.08 ;
      RECT 18.165 -54.97 18.515 -54.85 ;
      RECT 18.165 -51.74 18.515 -51.62 ;
      RECT 18.165 -48.51 18.515 -48.39 ;
      RECT 18.165 -45.28 18.515 -45.16 ;
      RECT 18.165 -42.05 18.515 -41.93 ;
      RECT 18.165 -38.82 18.515 -38.7 ;
      RECT 18.165 -35.59 18.515 -35.47 ;
      RECT 18.165 -32.36 18.515 -32.24 ;
      RECT 18.165 -29.13 18.515 -29.01 ;
      RECT 18.165 -25.9 18.515 -25.78 ;
      RECT 18.165 -22.67 18.515 -22.55 ;
      RECT 18.165 -19.44 18.515 -19.32 ;
      RECT 18.165 -16.21 18.515 -16.09 ;
      RECT 18.165 -12.98 18.515 -12.86 ;
      RECT 18.165 -9.75 18.515 -9.63 ;
      RECT 18.165 -6.52 18.515 -6.4 ;
      RECT 18.165 -3.29 18.515 -3.17 ;
      RECT 18.165 -0.06 18.515 0.06 ;
      RECT 18.335 -104.945 18.435 -103.985 ;
      RECT 18.335 2.175 18.435 3.135 ;
      RECT 14.435 -108.655 18.215 -108.535 ;
      RECT 18.075 -104.945 18.175 -103.985 ;
      RECT 17.95 -101.06 18.05 -100.525 ;
      RECT 17.95 -99.735 18.05 -99.2 ;
      RECT 17.95 -97.83 18.05 -97.295 ;
      RECT 17.95 -96.505 18.05 -95.97 ;
      RECT 17.95 -94.6 18.05 -94.065 ;
      RECT 17.95 -93.275 18.05 -92.74 ;
      RECT 17.95 -91.37 18.05 -90.835 ;
      RECT 17.95 -90.045 18.05 -89.51 ;
      RECT 17.95 -88.14 18.05 -87.605 ;
      RECT 17.95 -86.815 18.05 -86.28 ;
      RECT 17.95 -84.91 18.05 -84.375 ;
      RECT 17.95 -83.585 18.05 -83.05 ;
      RECT 17.95 -81.68 18.05 -81.145 ;
      RECT 17.95 -80.355 18.05 -79.82 ;
      RECT 17.95 -78.45 18.05 -77.915 ;
      RECT 17.95 -77.125 18.05 -76.59 ;
      RECT 17.95 -75.22 18.05 -74.685 ;
      RECT 17.95 -73.895 18.05 -73.36 ;
      RECT 17.95 -71.99 18.05 -71.455 ;
      RECT 17.95 -70.665 18.05 -70.13 ;
      RECT 17.95 -68.76 18.05 -68.225 ;
      RECT 17.95 -67.435 18.05 -66.9 ;
      RECT 17.95 -65.53 18.05 -64.995 ;
      RECT 17.95 -64.205 18.05 -63.67 ;
      RECT 17.95 -62.3 18.05 -61.765 ;
      RECT 17.95 -60.975 18.05 -60.44 ;
      RECT 17.95 -59.07 18.05 -58.535 ;
      RECT 17.95 -57.745 18.05 -57.21 ;
      RECT 17.95 -55.84 18.05 -55.305 ;
      RECT 17.95 -54.515 18.05 -53.98 ;
      RECT 17.95 -52.61 18.05 -52.075 ;
      RECT 17.95 -51.285 18.05 -50.75 ;
      RECT 17.95 -49.38 18.05 -48.845 ;
      RECT 17.95 -48.055 18.05 -47.52 ;
      RECT 17.95 -46.15 18.05 -45.615 ;
      RECT 17.95 -44.825 18.05 -44.29 ;
      RECT 17.95 -42.92 18.05 -42.385 ;
      RECT 17.95 -41.595 18.05 -41.06 ;
      RECT 17.95 -39.69 18.05 -39.155 ;
      RECT 17.95 -38.365 18.05 -37.83 ;
      RECT 17.95 -36.46 18.05 -35.925 ;
      RECT 17.95 -35.135 18.05 -34.6 ;
      RECT 17.95 -33.23 18.05 -32.695 ;
      RECT 17.95 -31.905 18.05 -31.37 ;
      RECT 17.95 -30 18.05 -29.465 ;
      RECT 17.95 -28.675 18.05 -28.14 ;
      RECT 17.95 -26.77 18.05 -26.235 ;
      RECT 17.95 -25.445 18.05 -24.91 ;
      RECT 17.95 -23.54 18.05 -23.005 ;
      RECT 17.95 -22.215 18.05 -21.68 ;
      RECT 17.95 -20.31 18.05 -19.775 ;
      RECT 17.95 -18.985 18.05 -18.45 ;
      RECT 17.95 -17.08 18.05 -16.545 ;
      RECT 17.95 -15.755 18.05 -15.22 ;
      RECT 17.95 -13.85 18.05 -13.315 ;
      RECT 17.95 -12.525 18.05 -11.99 ;
      RECT 17.95 -10.62 18.05 -10.085 ;
      RECT 17.95 -9.295 18.05 -8.76 ;
      RECT 17.95 -7.39 18.05 -6.855 ;
      RECT 17.95 -6.065 18.05 -5.53 ;
      RECT 17.95 -4.16 18.05 -3.625 ;
      RECT 17.95 -2.835 18.05 -2.3 ;
      RECT 17.95 -0.93 18.05 -0.395 ;
      RECT 17.95 0.395 18.05 0.93 ;
      RECT 17.885 -110.75 18.005 -110.37 ;
      RECT 17.885 -112.245 17.985 -111.775 ;
      RECT 17.825 -104.945 17.925 -103.985 ;
      RECT 17.45 -100.19 17.8 -100.07 ;
      RECT 17.45 -96.96 17.8 -96.84 ;
      RECT 17.45 -93.73 17.8 -93.61 ;
      RECT 17.45 -90.5 17.8 -90.38 ;
      RECT 17.45 -87.27 17.8 -87.15 ;
      RECT 17.45 -84.04 17.8 -83.92 ;
      RECT 17.45 -80.81 17.8 -80.69 ;
      RECT 17.45 -77.58 17.8 -77.46 ;
      RECT 17.45 -74.35 17.8 -74.23 ;
      RECT 17.45 -71.12 17.8 -71 ;
      RECT 17.45 -67.89 17.8 -67.77 ;
      RECT 17.45 -64.66 17.8 -64.54 ;
      RECT 17.45 -61.43 17.8 -61.31 ;
      RECT 17.45 -58.2 17.8 -58.08 ;
      RECT 17.45 -54.97 17.8 -54.85 ;
      RECT 17.45 -51.74 17.8 -51.62 ;
      RECT 17.45 -48.51 17.8 -48.39 ;
      RECT 17.45 -45.28 17.8 -45.16 ;
      RECT 17.45 -42.05 17.8 -41.93 ;
      RECT 17.45 -38.82 17.8 -38.7 ;
      RECT 17.45 -35.59 17.8 -35.47 ;
      RECT 17.45 -32.36 17.8 -32.24 ;
      RECT 17.45 -29.13 17.8 -29.01 ;
      RECT 17.45 -25.9 17.8 -25.78 ;
      RECT 17.45 -22.67 17.8 -22.55 ;
      RECT 17.45 -19.44 17.8 -19.32 ;
      RECT 17.45 -16.21 17.8 -16.09 ;
      RECT 17.45 -12.98 17.8 -12.86 ;
      RECT 17.45 -9.75 17.8 -9.63 ;
      RECT 17.45 -6.52 17.8 -6.4 ;
      RECT 17.45 -3.29 17.8 -3.17 ;
      RECT 17.45 -0.06 17.8 0.06 ;
      RECT 17.565 -104.945 17.665 -103.985 ;
      RECT 17.565 2.175 17.665 3.135 ;
      RECT 17.295 -109.595 17.43 -109.275 ;
      RECT 16.965 -100.19 17.315 -100.07 ;
      RECT 16.965 -96.96 17.315 -96.84 ;
      RECT 16.965 -93.73 17.315 -93.61 ;
      RECT 16.965 -90.5 17.315 -90.38 ;
      RECT 16.965 -87.27 17.315 -87.15 ;
      RECT 16.965 -84.04 17.315 -83.92 ;
      RECT 16.965 -80.81 17.315 -80.69 ;
      RECT 16.965 -77.58 17.315 -77.46 ;
      RECT 16.965 -74.35 17.315 -74.23 ;
      RECT 16.965 -71.12 17.315 -71 ;
      RECT 16.965 -67.89 17.315 -67.77 ;
      RECT 16.965 -64.66 17.315 -64.54 ;
      RECT 16.965 -61.43 17.315 -61.31 ;
      RECT 16.965 -58.2 17.315 -58.08 ;
      RECT 16.965 -54.97 17.315 -54.85 ;
      RECT 16.965 -51.74 17.315 -51.62 ;
      RECT 16.965 -48.51 17.315 -48.39 ;
      RECT 16.965 -45.28 17.315 -45.16 ;
      RECT 16.965 -42.05 17.315 -41.93 ;
      RECT 16.965 -38.82 17.315 -38.7 ;
      RECT 16.965 -35.59 17.315 -35.47 ;
      RECT 16.965 -32.36 17.315 -32.24 ;
      RECT 16.965 -29.13 17.315 -29.01 ;
      RECT 16.965 -25.9 17.315 -25.78 ;
      RECT 16.965 -22.67 17.315 -22.55 ;
      RECT 16.965 -19.44 17.315 -19.32 ;
      RECT 16.965 -16.21 17.315 -16.09 ;
      RECT 16.965 -12.98 17.315 -12.86 ;
      RECT 16.965 -9.75 17.315 -9.63 ;
      RECT 16.965 -6.52 17.315 -6.4 ;
      RECT 16.965 -3.29 17.315 -3.17 ;
      RECT 16.965 -0.06 17.315 0.06 ;
      RECT 17.135 -104.945 17.235 -103.985 ;
      RECT 17.135 2.175 17.235 3.135 ;
      RECT 16.96 -109.595 17.105 -109.275 ;
      RECT 16.875 -104.945 16.975 -103.985 ;
      RECT 16.75 -101.06 16.85 -100.525 ;
      RECT 16.75 -99.735 16.85 -99.2 ;
      RECT 16.75 -97.83 16.85 -97.295 ;
      RECT 16.75 -96.505 16.85 -95.97 ;
      RECT 16.75 -94.6 16.85 -94.065 ;
      RECT 16.75 -93.275 16.85 -92.74 ;
      RECT 16.75 -91.37 16.85 -90.835 ;
      RECT 16.75 -90.045 16.85 -89.51 ;
      RECT 16.75 -88.14 16.85 -87.605 ;
      RECT 16.75 -86.815 16.85 -86.28 ;
      RECT 16.75 -84.91 16.85 -84.375 ;
      RECT 16.75 -83.585 16.85 -83.05 ;
      RECT 16.75 -81.68 16.85 -81.145 ;
      RECT 16.75 -80.355 16.85 -79.82 ;
      RECT 16.75 -78.45 16.85 -77.915 ;
      RECT 16.75 -77.125 16.85 -76.59 ;
      RECT 16.75 -75.22 16.85 -74.685 ;
      RECT 16.75 -73.895 16.85 -73.36 ;
      RECT 16.75 -71.99 16.85 -71.455 ;
      RECT 16.75 -70.665 16.85 -70.13 ;
      RECT 16.75 -68.76 16.85 -68.225 ;
      RECT 16.75 -67.435 16.85 -66.9 ;
      RECT 16.75 -65.53 16.85 -64.995 ;
      RECT 16.75 -64.205 16.85 -63.67 ;
      RECT 16.75 -62.3 16.85 -61.765 ;
      RECT 16.75 -60.975 16.85 -60.44 ;
      RECT 16.75 -59.07 16.85 -58.535 ;
      RECT 16.75 -57.745 16.85 -57.21 ;
      RECT 16.75 -55.84 16.85 -55.305 ;
      RECT 16.75 -54.515 16.85 -53.98 ;
      RECT 16.75 -52.61 16.85 -52.075 ;
      RECT 16.75 -51.285 16.85 -50.75 ;
      RECT 16.75 -49.38 16.85 -48.845 ;
      RECT 16.75 -48.055 16.85 -47.52 ;
      RECT 16.75 -46.15 16.85 -45.615 ;
      RECT 16.75 -44.825 16.85 -44.29 ;
      RECT 16.75 -42.92 16.85 -42.385 ;
      RECT 16.75 -41.595 16.85 -41.06 ;
      RECT 16.75 -39.69 16.85 -39.155 ;
      RECT 16.75 -38.365 16.85 -37.83 ;
      RECT 16.75 -36.46 16.85 -35.925 ;
      RECT 16.75 -35.135 16.85 -34.6 ;
      RECT 16.75 -33.23 16.85 -32.695 ;
      RECT 16.75 -31.905 16.85 -31.37 ;
      RECT 16.75 -30 16.85 -29.465 ;
      RECT 16.75 -28.675 16.85 -28.14 ;
      RECT 16.75 -26.77 16.85 -26.235 ;
      RECT 16.75 -25.445 16.85 -24.91 ;
      RECT 16.75 -23.54 16.85 -23.005 ;
      RECT 16.75 -22.215 16.85 -21.68 ;
      RECT 16.75 -20.31 16.85 -19.775 ;
      RECT 16.75 -18.985 16.85 -18.45 ;
      RECT 16.75 -17.08 16.85 -16.545 ;
      RECT 16.75 -15.755 16.85 -15.22 ;
      RECT 16.75 -13.85 16.85 -13.315 ;
      RECT 16.75 -12.525 16.85 -11.99 ;
      RECT 16.75 -10.62 16.85 -10.085 ;
      RECT 16.75 -9.295 16.85 -8.76 ;
      RECT 16.75 -7.39 16.85 -6.855 ;
      RECT 16.75 -6.065 16.85 -5.53 ;
      RECT 16.75 -4.16 16.85 -3.625 ;
      RECT 16.75 -2.835 16.85 -2.3 ;
      RECT 16.75 -0.93 16.85 -0.395 ;
      RECT 16.75 0.395 16.85 0.93 ;
      RECT 16.625 -108.175 16.725 -107.215 ;
      RECT 16.25 -100.19 16.6 -100.07 ;
      RECT 16.25 -96.96 16.6 -96.84 ;
      RECT 16.25 -93.73 16.6 -93.61 ;
      RECT 16.25 -90.5 16.6 -90.38 ;
      RECT 16.25 -87.27 16.6 -87.15 ;
      RECT 16.25 -84.04 16.6 -83.92 ;
      RECT 16.25 -80.81 16.6 -80.69 ;
      RECT 16.25 -77.58 16.6 -77.46 ;
      RECT 16.25 -74.35 16.6 -74.23 ;
      RECT 16.25 -71.12 16.6 -71 ;
      RECT 16.25 -67.89 16.6 -67.77 ;
      RECT 16.25 -64.66 16.6 -64.54 ;
      RECT 16.25 -61.43 16.6 -61.31 ;
      RECT 16.25 -58.2 16.6 -58.08 ;
      RECT 16.25 -54.97 16.6 -54.85 ;
      RECT 16.25 -51.74 16.6 -51.62 ;
      RECT 16.25 -48.51 16.6 -48.39 ;
      RECT 16.25 -45.28 16.6 -45.16 ;
      RECT 16.25 -42.05 16.6 -41.93 ;
      RECT 16.25 -38.82 16.6 -38.7 ;
      RECT 16.25 -35.59 16.6 -35.47 ;
      RECT 16.25 -32.36 16.6 -32.24 ;
      RECT 16.25 -29.13 16.6 -29.01 ;
      RECT 16.25 -25.9 16.6 -25.78 ;
      RECT 16.25 -22.67 16.6 -22.55 ;
      RECT 16.25 -19.44 16.6 -19.32 ;
      RECT 16.25 -16.21 16.6 -16.09 ;
      RECT 16.25 -12.98 16.6 -12.86 ;
      RECT 16.25 -9.75 16.6 -9.63 ;
      RECT 16.25 -6.52 16.6 -6.4 ;
      RECT 16.25 -3.29 16.6 -3.17 ;
      RECT 16.25 -0.06 16.6 0.06 ;
      RECT 16.455 -112.255 16.555 -111.775 ;
      RECT 16.455 -110.765 16.555 -110.295 ;
      RECT 16.365 -108.175 16.465 -107.215 ;
      RECT 16.365 2.175 16.465 3.135 ;
      RECT 15.765 -100.19 16.115 -100.07 ;
      RECT 15.765 -96.96 16.115 -96.84 ;
      RECT 15.765 -93.73 16.115 -93.61 ;
      RECT 15.765 -90.5 16.115 -90.38 ;
      RECT 15.765 -87.27 16.115 -87.15 ;
      RECT 15.765 -84.04 16.115 -83.92 ;
      RECT 15.765 -80.81 16.115 -80.69 ;
      RECT 15.765 -77.58 16.115 -77.46 ;
      RECT 15.765 -74.35 16.115 -74.23 ;
      RECT 15.765 -71.12 16.115 -71 ;
      RECT 15.765 -67.89 16.115 -67.77 ;
      RECT 15.765 -64.66 16.115 -64.54 ;
      RECT 15.765 -61.43 16.115 -61.31 ;
      RECT 15.765 -58.2 16.115 -58.08 ;
      RECT 15.765 -54.97 16.115 -54.85 ;
      RECT 15.765 -51.74 16.115 -51.62 ;
      RECT 15.765 -48.51 16.115 -48.39 ;
      RECT 15.765 -45.28 16.115 -45.16 ;
      RECT 15.765 -42.05 16.115 -41.93 ;
      RECT 15.765 -38.82 16.115 -38.7 ;
      RECT 15.765 -35.59 16.115 -35.47 ;
      RECT 15.765 -32.36 16.115 -32.24 ;
      RECT 15.765 -29.13 16.115 -29.01 ;
      RECT 15.765 -25.9 16.115 -25.78 ;
      RECT 15.765 -22.67 16.115 -22.55 ;
      RECT 15.765 -19.44 16.115 -19.32 ;
      RECT 15.765 -16.21 16.115 -16.09 ;
      RECT 15.765 -12.98 16.115 -12.86 ;
      RECT 15.765 -9.75 16.115 -9.63 ;
      RECT 15.765 -6.52 16.115 -6.4 ;
      RECT 15.765 -3.29 16.115 -3.17 ;
      RECT 15.765 -0.06 16.115 0.06 ;
      RECT 15.935 -108.175 16.035 -107.215 ;
      RECT 15.935 2.175 16.035 3.135 ;
      RECT 15.83 -110.765 16 -110.385 ;
      RECT 15.865 -112.245 15.965 -111.775 ;
      RECT 15.675 -108.175 15.775 -107.215 ;
      RECT 15.55 -101.06 15.65 -100.525 ;
      RECT 15.55 -99.735 15.65 -99.2 ;
      RECT 15.55 -97.83 15.65 -97.295 ;
      RECT 15.55 -96.505 15.65 -95.97 ;
      RECT 15.55 -94.6 15.65 -94.065 ;
      RECT 15.55 -93.275 15.65 -92.74 ;
      RECT 15.55 -91.37 15.65 -90.835 ;
      RECT 15.55 -90.045 15.65 -89.51 ;
      RECT 15.55 -88.14 15.65 -87.605 ;
      RECT 15.55 -86.815 15.65 -86.28 ;
      RECT 15.55 -84.91 15.65 -84.375 ;
      RECT 15.55 -83.585 15.65 -83.05 ;
      RECT 15.55 -81.68 15.65 -81.145 ;
      RECT 15.55 -80.355 15.65 -79.82 ;
      RECT 15.55 -78.45 15.65 -77.915 ;
      RECT 15.55 -77.125 15.65 -76.59 ;
      RECT 15.55 -75.22 15.65 -74.685 ;
      RECT 15.55 -73.895 15.65 -73.36 ;
      RECT 15.55 -71.99 15.65 -71.455 ;
      RECT 15.55 -70.665 15.65 -70.13 ;
      RECT 15.55 -68.76 15.65 -68.225 ;
      RECT 15.55 -67.435 15.65 -66.9 ;
      RECT 15.55 -65.53 15.65 -64.995 ;
      RECT 15.55 -64.205 15.65 -63.67 ;
      RECT 15.55 -62.3 15.65 -61.765 ;
      RECT 15.55 -60.975 15.65 -60.44 ;
      RECT 15.55 -59.07 15.65 -58.535 ;
      RECT 15.55 -57.745 15.65 -57.21 ;
      RECT 15.55 -55.84 15.65 -55.305 ;
      RECT 15.55 -54.515 15.65 -53.98 ;
      RECT 15.55 -52.61 15.65 -52.075 ;
      RECT 15.55 -51.285 15.65 -50.75 ;
      RECT 15.55 -49.38 15.65 -48.845 ;
      RECT 15.55 -48.055 15.65 -47.52 ;
      RECT 15.55 -46.15 15.65 -45.615 ;
      RECT 15.55 -44.825 15.65 -44.29 ;
      RECT 15.55 -42.92 15.65 -42.385 ;
      RECT 15.55 -41.595 15.65 -41.06 ;
      RECT 15.55 -39.69 15.65 -39.155 ;
      RECT 15.55 -38.365 15.65 -37.83 ;
      RECT 15.55 -36.46 15.65 -35.925 ;
      RECT 15.55 -35.135 15.65 -34.6 ;
      RECT 15.55 -33.23 15.65 -32.695 ;
      RECT 15.55 -31.905 15.65 -31.37 ;
      RECT 15.55 -30 15.65 -29.465 ;
      RECT 15.55 -28.675 15.65 -28.14 ;
      RECT 15.55 -26.77 15.65 -26.235 ;
      RECT 15.55 -25.445 15.65 -24.91 ;
      RECT 15.55 -23.54 15.65 -23.005 ;
      RECT 15.55 -22.215 15.65 -21.68 ;
      RECT 15.55 -20.31 15.65 -19.775 ;
      RECT 15.55 -18.985 15.65 -18.45 ;
      RECT 15.55 -17.08 15.65 -16.545 ;
      RECT 15.55 -15.755 15.65 -15.22 ;
      RECT 15.55 -13.85 15.65 -13.315 ;
      RECT 15.55 -12.525 15.65 -11.99 ;
      RECT 15.55 -10.62 15.65 -10.085 ;
      RECT 15.55 -9.295 15.65 -8.76 ;
      RECT 15.55 -7.39 15.65 -6.855 ;
      RECT 15.55 -6.065 15.65 -5.53 ;
      RECT 15.55 -4.16 15.65 -3.625 ;
      RECT 15.55 -2.835 15.65 -2.3 ;
      RECT 15.55 -0.93 15.65 -0.395 ;
      RECT 15.55 0.395 15.65 0.93 ;
      RECT 15.425 -108.175 15.525 -107.215 ;
      RECT 15.05 -100.19 15.4 -100.07 ;
      RECT 15.05 -96.96 15.4 -96.84 ;
      RECT 15.05 -93.73 15.4 -93.61 ;
      RECT 15.05 -90.5 15.4 -90.38 ;
      RECT 15.05 -87.27 15.4 -87.15 ;
      RECT 15.05 -84.04 15.4 -83.92 ;
      RECT 15.05 -80.81 15.4 -80.69 ;
      RECT 15.05 -77.58 15.4 -77.46 ;
      RECT 15.05 -74.35 15.4 -74.23 ;
      RECT 15.05 -71.12 15.4 -71 ;
      RECT 15.05 -67.89 15.4 -67.77 ;
      RECT 15.05 -64.66 15.4 -64.54 ;
      RECT 15.05 -61.43 15.4 -61.31 ;
      RECT 15.05 -58.2 15.4 -58.08 ;
      RECT 15.05 -54.97 15.4 -54.85 ;
      RECT 15.05 -51.74 15.4 -51.62 ;
      RECT 15.05 -48.51 15.4 -48.39 ;
      RECT 15.05 -45.28 15.4 -45.16 ;
      RECT 15.05 -42.05 15.4 -41.93 ;
      RECT 15.05 -38.82 15.4 -38.7 ;
      RECT 15.05 -35.59 15.4 -35.47 ;
      RECT 15.05 -32.36 15.4 -32.24 ;
      RECT 15.05 -29.13 15.4 -29.01 ;
      RECT 15.05 -25.9 15.4 -25.78 ;
      RECT 15.05 -22.67 15.4 -22.55 ;
      RECT 15.05 -19.44 15.4 -19.32 ;
      RECT 15.05 -16.21 15.4 -16.09 ;
      RECT 15.05 -12.98 15.4 -12.86 ;
      RECT 15.05 -9.75 15.4 -9.63 ;
      RECT 15.05 -6.52 15.4 -6.4 ;
      RECT 15.05 -3.29 15.4 -3.17 ;
      RECT 15.05 -0.06 15.4 0.06 ;
      RECT 15.165 -108.175 15.265 -107.215 ;
      RECT 15.165 2.175 15.265 3.135 ;
      RECT 15.065 -113.555 15.165 -113.085 ;
      RECT 14.565 -100.19 14.915 -100.07 ;
      RECT 14.565 -96.96 14.915 -96.84 ;
      RECT 14.565 -93.73 14.915 -93.61 ;
      RECT 14.565 -90.5 14.915 -90.38 ;
      RECT 14.565 -87.27 14.915 -87.15 ;
      RECT 14.565 -84.04 14.915 -83.92 ;
      RECT 14.565 -80.81 14.915 -80.69 ;
      RECT 14.565 -77.58 14.915 -77.46 ;
      RECT 14.565 -74.35 14.915 -74.23 ;
      RECT 14.565 -71.12 14.915 -71 ;
      RECT 14.565 -67.89 14.915 -67.77 ;
      RECT 14.565 -64.66 14.915 -64.54 ;
      RECT 14.565 -61.43 14.915 -61.31 ;
      RECT 14.565 -58.2 14.915 -58.08 ;
      RECT 14.565 -54.97 14.915 -54.85 ;
      RECT 14.565 -51.74 14.915 -51.62 ;
      RECT 14.565 -48.51 14.915 -48.39 ;
      RECT 14.565 -45.28 14.915 -45.16 ;
      RECT 14.565 -42.05 14.915 -41.93 ;
      RECT 14.565 -38.82 14.915 -38.7 ;
      RECT 14.565 -35.59 14.915 -35.47 ;
      RECT 14.565 -32.36 14.915 -32.24 ;
      RECT 14.565 -29.13 14.915 -29.01 ;
      RECT 14.565 -25.9 14.915 -25.78 ;
      RECT 14.565 -22.67 14.915 -22.55 ;
      RECT 14.565 -19.44 14.915 -19.32 ;
      RECT 14.565 -16.21 14.915 -16.09 ;
      RECT 14.565 -12.98 14.915 -12.86 ;
      RECT 14.565 -9.75 14.915 -9.63 ;
      RECT 14.565 -6.52 14.915 -6.4 ;
      RECT 14.565 -3.29 14.915 -3.17 ;
      RECT 14.565 -0.06 14.915 0.06 ;
      RECT 14.7 -110.735 14.85 -110.445 ;
      RECT 14.735 -108.175 14.835 -107.215 ;
      RECT 14.735 2.175 14.835 3.135 ;
      RECT 14.715 -112.19 14.815 -111.65 ;
      RECT 14.475 -113.555 14.575 -113.085 ;
      RECT 14.475 -108.175 14.575 -107.215 ;
      RECT 14.35 -101.06 14.45 -100.525 ;
      RECT 14.35 -99.735 14.45 -99.2 ;
      RECT 14.35 -97.83 14.45 -97.295 ;
      RECT 14.35 -96.505 14.45 -95.97 ;
      RECT 14.35 -94.6 14.45 -94.065 ;
      RECT 14.35 -93.275 14.45 -92.74 ;
      RECT 14.35 -91.37 14.45 -90.835 ;
      RECT 14.35 -90.045 14.45 -89.51 ;
      RECT 14.35 -88.14 14.45 -87.605 ;
      RECT 14.35 -86.815 14.45 -86.28 ;
      RECT 14.35 -84.91 14.45 -84.375 ;
      RECT 14.35 -83.585 14.45 -83.05 ;
      RECT 14.35 -81.68 14.45 -81.145 ;
      RECT 14.35 -80.355 14.45 -79.82 ;
      RECT 14.35 -78.45 14.45 -77.915 ;
      RECT 14.35 -77.125 14.45 -76.59 ;
      RECT 14.35 -75.22 14.45 -74.685 ;
      RECT 14.35 -73.895 14.45 -73.36 ;
      RECT 14.35 -71.99 14.45 -71.455 ;
      RECT 14.35 -70.665 14.45 -70.13 ;
      RECT 14.35 -68.76 14.45 -68.225 ;
      RECT 14.35 -67.435 14.45 -66.9 ;
      RECT 14.35 -65.53 14.45 -64.995 ;
      RECT 14.35 -64.205 14.45 -63.67 ;
      RECT 14.35 -62.3 14.45 -61.765 ;
      RECT 14.35 -60.975 14.45 -60.44 ;
      RECT 14.35 -59.07 14.45 -58.535 ;
      RECT 14.35 -57.745 14.45 -57.21 ;
      RECT 14.35 -55.84 14.45 -55.305 ;
      RECT 14.35 -54.515 14.45 -53.98 ;
      RECT 14.35 -52.61 14.45 -52.075 ;
      RECT 14.35 -51.285 14.45 -50.75 ;
      RECT 14.35 -49.38 14.45 -48.845 ;
      RECT 14.35 -48.055 14.45 -47.52 ;
      RECT 14.35 -46.15 14.45 -45.615 ;
      RECT 14.35 -44.825 14.45 -44.29 ;
      RECT 14.35 -42.92 14.45 -42.385 ;
      RECT 14.35 -41.595 14.45 -41.06 ;
      RECT 14.35 -39.69 14.45 -39.155 ;
      RECT 14.35 -38.365 14.45 -37.83 ;
      RECT 14.35 -36.46 14.45 -35.925 ;
      RECT 14.35 -35.135 14.45 -34.6 ;
      RECT 14.35 -33.23 14.45 -32.695 ;
      RECT 14.35 -31.905 14.45 -31.37 ;
      RECT 14.35 -30 14.45 -29.465 ;
      RECT 14.35 -28.675 14.45 -28.14 ;
      RECT 14.35 -26.77 14.45 -26.235 ;
      RECT 14.35 -25.445 14.45 -24.91 ;
      RECT 14.35 -23.54 14.45 -23.005 ;
      RECT 14.35 -22.215 14.45 -21.68 ;
      RECT 14.35 -20.31 14.45 -19.775 ;
      RECT 14.35 -18.985 14.45 -18.45 ;
      RECT 14.35 -17.08 14.45 -16.545 ;
      RECT 14.35 -15.755 14.45 -15.22 ;
      RECT 14.35 -13.85 14.45 -13.315 ;
      RECT 14.35 -12.525 14.45 -11.99 ;
      RECT 14.35 -10.62 14.45 -10.085 ;
      RECT 14.35 -9.295 14.45 -8.76 ;
      RECT 14.35 -7.39 14.45 -6.855 ;
      RECT 14.35 -6.065 14.45 -5.53 ;
      RECT 14.35 -4.16 14.45 -3.625 ;
      RECT 14.35 -2.835 14.45 -2.3 ;
      RECT 14.35 -0.93 14.45 -0.395 ;
      RECT 14.35 0.395 14.45 0.93 ;
      RECT 14.225 -104.945 14.325 -103.985 ;
      RECT 13.85 -100.19 14.2 -100.07 ;
      RECT 13.85 -96.96 14.2 -96.84 ;
      RECT 13.85 -93.73 14.2 -93.61 ;
      RECT 13.85 -90.5 14.2 -90.38 ;
      RECT 13.85 -87.27 14.2 -87.15 ;
      RECT 13.85 -84.04 14.2 -83.92 ;
      RECT 13.85 -80.81 14.2 -80.69 ;
      RECT 13.85 -77.58 14.2 -77.46 ;
      RECT 13.85 -74.35 14.2 -74.23 ;
      RECT 13.85 -71.12 14.2 -71 ;
      RECT 13.85 -67.89 14.2 -67.77 ;
      RECT 13.85 -64.66 14.2 -64.54 ;
      RECT 13.85 -61.43 14.2 -61.31 ;
      RECT 13.85 -58.2 14.2 -58.08 ;
      RECT 13.85 -54.97 14.2 -54.85 ;
      RECT 13.85 -51.74 14.2 -51.62 ;
      RECT 13.85 -48.51 14.2 -48.39 ;
      RECT 13.85 -45.28 14.2 -45.16 ;
      RECT 13.85 -42.05 14.2 -41.93 ;
      RECT 13.85 -38.82 14.2 -38.7 ;
      RECT 13.85 -35.59 14.2 -35.47 ;
      RECT 13.85 -32.36 14.2 -32.24 ;
      RECT 13.85 -29.13 14.2 -29.01 ;
      RECT 13.85 -25.9 14.2 -25.78 ;
      RECT 13.85 -22.67 14.2 -22.55 ;
      RECT 13.85 -19.44 14.2 -19.32 ;
      RECT 13.85 -16.21 14.2 -16.09 ;
      RECT 13.85 -12.98 14.2 -12.86 ;
      RECT 13.85 -9.75 14.2 -9.63 ;
      RECT 13.85 -6.52 14.2 -6.4 ;
      RECT 13.85 -3.29 14.2 -3.17 ;
      RECT 13.85 -0.06 14.2 0.06 ;
      RECT 13.965 -104.945 14.065 -103.985 ;
      RECT 13.965 2.175 14.065 3.135 ;
      RECT 13.675 -112.255 13.775 -111.775 ;
      RECT 13.675 -110.765 13.775 -110.295 ;
      RECT 13.365 -100.19 13.715 -100.07 ;
      RECT 13.365 -96.96 13.715 -96.84 ;
      RECT 13.365 -93.73 13.715 -93.61 ;
      RECT 13.365 -90.5 13.715 -90.38 ;
      RECT 13.365 -87.27 13.715 -87.15 ;
      RECT 13.365 -84.04 13.715 -83.92 ;
      RECT 13.365 -80.81 13.715 -80.69 ;
      RECT 13.365 -77.58 13.715 -77.46 ;
      RECT 13.365 -74.35 13.715 -74.23 ;
      RECT 13.365 -71.12 13.715 -71 ;
      RECT 13.365 -67.89 13.715 -67.77 ;
      RECT 13.365 -64.66 13.715 -64.54 ;
      RECT 13.365 -61.43 13.715 -61.31 ;
      RECT 13.365 -58.2 13.715 -58.08 ;
      RECT 13.365 -54.97 13.715 -54.85 ;
      RECT 13.365 -51.74 13.715 -51.62 ;
      RECT 13.365 -48.51 13.715 -48.39 ;
      RECT 13.365 -45.28 13.715 -45.16 ;
      RECT 13.365 -42.05 13.715 -41.93 ;
      RECT 13.365 -38.82 13.715 -38.7 ;
      RECT 13.365 -35.59 13.715 -35.47 ;
      RECT 13.365 -32.36 13.715 -32.24 ;
      RECT 13.365 -29.13 13.715 -29.01 ;
      RECT 13.365 -25.9 13.715 -25.78 ;
      RECT 13.365 -22.67 13.715 -22.55 ;
      RECT 13.365 -19.44 13.715 -19.32 ;
      RECT 13.365 -16.21 13.715 -16.09 ;
      RECT 13.365 -12.98 13.715 -12.86 ;
      RECT 13.365 -9.75 13.715 -9.63 ;
      RECT 13.365 -6.52 13.715 -6.4 ;
      RECT 13.365 -3.29 13.715 -3.17 ;
      RECT 13.365 -0.06 13.715 0.06 ;
      RECT 13.535 -104.945 13.635 -103.985 ;
      RECT 13.535 2.175 13.635 3.135 ;
      RECT 9.635 -108.655 13.415 -108.535 ;
      RECT 13.275 -104.945 13.375 -103.985 ;
      RECT 13.15 -101.06 13.25 -100.525 ;
      RECT 13.15 -99.735 13.25 -99.2 ;
      RECT 13.15 -97.83 13.25 -97.295 ;
      RECT 13.15 -96.505 13.25 -95.97 ;
      RECT 13.15 -94.6 13.25 -94.065 ;
      RECT 13.15 -93.275 13.25 -92.74 ;
      RECT 13.15 -91.37 13.25 -90.835 ;
      RECT 13.15 -90.045 13.25 -89.51 ;
      RECT 13.15 -88.14 13.25 -87.605 ;
      RECT 13.15 -86.815 13.25 -86.28 ;
      RECT 13.15 -84.91 13.25 -84.375 ;
      RECT 13.15 -83.585 13.25 -83.05 ;
      RECT 13.15 -81.68 13.25 -81.145 ;
      RECT 13.15 -80.355 13.25 -79.82 ;
      RECT 13.15 -78.45 13.25 -77.915 ;
      RECT 13.15 -77.125 13.25 -76.59 ;
      RECT 13.15 -75.22 13.25 -74.685 ;
      RECT 13.15 -73.895 13.25 -73.36 ;
      RECT 13.15 -71.99 13.25 -71.455 ;
      RECT 13.15 -70.665 13.25 -70.13 ;
      RECT 13.15 -68.76 13.25 -68.225 ;
      RECT 13.15 -67.435 13.25 -66.9 ;
      RECT 13.15 -65.53 13.25 -64.995 ;
      RECT 13.15 -64.205 13.25 -63.67 ;
      RECT 13.15 -62.3 13.25 -61.765 ;
      RECT 13.15 -60.975 13.25 -60.44 ;
      RECT 13.15 -59.07 13.25 -58.535 ;
      RECT 13.15 -57.745 13.25 -57.21 ;
      RECT 13.15 -55.84 13.25 -55.305 ;
      RECT 13.15 -54.515 13.25 -53.98 ;
      RECT 13.15 -52.61 13.25 -52.075 ;
      RECT 13.15 -51.285 13.25 -50.75 ;
      RECT 13.15 -49.38 13.25 -48.845 ;
      RECT 13.15 -48.055 13.25 -47.52 ;
      RECT 13.15 -46.15 13.25 -45.615 ;
      RECT 13.15 -44.825 13.25 -44.29 ;
      RECT 13.15 -42.92 13.25 -42.385 ;
      RECT 13.15 -41.595 13.25 -41.06 ;
      RECT 13.15 -39.69 13.25 -39.155 ;
      RECT 13.15 -38.365 13.25 -37.83 ;
      RECT 13.15 -36.46 13.25 -35.925 ;
      RECT 13.15 -35.135 13.25 -34.6 ;
      RECT 13.15 -33.23 13.25 -32.695 ;
      RECT 13.15 -31.905 13.25 -31.37 ;
      RECT 13.15 -30 13.25 -29.465 ;
      RECT 13.15 -28.675 13.25 -28.14 ;
      RECT 13.15 -26.77 13.25 -26.235 ;
      RECT 13.15 -25.445 13.25 -24.91 ;
      RECT 13.15 -23.54 13.25 -23.005 ;
      RECT 13.15 -22.215 13.25 -21.68 ;
      RECT 13.15 -20.31 13.25 -19.775 ;
      RECT 13.15 -18.985 13.25 -18.45 ;
      RECT 13.15 -17.08 13.25 -16.545 ;
      RECT 13.15 -15.755 13.25 -15.22 ;
      RECT 13.15 -13.85 13.25 -13.315 ;
      RECT 13.15 -12.525 13.25 -11.99 ;
      RECT 13.15 -10.62 13.25 -10.085 ;
      RECT 13.15 -9.295 13.25 -8.76 ;
      RECT 13.15 -7.39 13.25 -6.855 ;
      RECT 13.15 -6.065 13.25 -5.53 ;
      RECT 13.15 -4.16 13.25 -3.625 ;
      RECT 13.15 -2.835 13.25 -2.3 ;
      RECT 13.15 -0.93 13.25 -0.395 ;
      RECT 13.15 0.395 13.25 0.93 ;
      RECT 13.085 -110.75 13.205 -110.37 ;
      RECT 13.085 -112.245 13.185 -111.775 ;
      RECT 13.025 -104.945 13.125 -103.985 ;
      RECT 12.65 -100.19 13 -100.07 ;
      RECT 12.65 -96.96 13 -96.84 ;
      RECT 12.65 -93.73 13 -93.61 ;
      RECT 12.65 -90.5 13 -90.38 ;
      RECT 12.65 -87.27 13 -87.15 ;
      RECT 12.65 -84.04 13 -83.92 ;
      RECT 12.65 -80.81 13 -80.69 ;
      RECT 12.65 -77.58 13 -77.46 ;
      RECT 12.65 -74.35 13 -74.23 ;
      RECT 12.65 -71.12 13 -71 ;
      RECT 12.65 -67.89 13 -67.77 ;
      RECT 12.65 -64.66 13 -64.54 ;
      RECT 12.65 -61.43 13 -61.31 ;
      RECT 12.65 -58.2 13 -58.08 ;
      RECT 12.65 -54.97 13 -54.85 ;
      RECT 12.65 -51.74 13 -51.62 ;
      RECT 12.65 -48.51 13 -48.39 ;
      RECT 12.65 -45.28 13 -45.16 ;
      RECT 12.65 -42.05 13 -41.93 ;
      RECT 12.65 -38.82 13 -38.7 ;
      RECT 12.65 -35.59 13 -35.47 ;
      RECT 12.65 -32.36 13 -32.24 ;
      RECT 12.65 -29.13 13 -29.01 ;
      RECT 12.65 -25.9 13 -25.78 ;
      RECT 12.65 -22.67 13 -22.55 ;
      RECT 12.65 -19.44 13 -19.32 ;
      RECT 12.65 -16.21 13 -16.09 ;
      RECT 12.65 -12.98 13 -12.86 ;
      RECT 12.65 -9.75 13 -9.63 ;
      RECT 12.65 -6.52 13 -6.4 ;
      RECT 12.65 -3.29 13 -3.17 ;
      RECT 12.65 -0.06 13 0.06 ;
      RECT 12.765 -104.945 12.865 -103.985 ;
      RECT 12.765 2.175 12.865 3.135 ;
      RECT 12.495 -109.595 12.63 -109.275 ;
      RECT 12.165 -100.19 12.515 -100.07 ;
      RECT 12.165 -96.96 12.515 -96.84 ;
      RECT 12.165 -93.73 12.515 -93.61 ;
      RECT 12.165 -90.5 12.515 -90.38 ;
      RECT 12.165 -87.27 12.515 -87.15 ;
      RECT 12.165 -84.04 12.515 -83.92 ;
      RECT 12.165 -80.81 12.515 -80.69 ;
      RECT 12.165 -77.58 12.515 -77.46 ;
      RECT 12.165 -74.35 12.515 -74.23 ;
      RECT 12.165 -71.12 12.515 -71 ;
      RECT 12.165 -67.89 12.515 -67.77 ;
      RECT 12.165 -64.66 12.515 -64.54 ;
      RECT 12.165 -61.43 12.515 -61.31 ;
      RECT 12.165 -58.2 12.515 -58.08 ;
      RECT 12.165 -54.97 12.515 -54.85 ;
      RECT 12.165 -51.74 12.515 -51.62 ;
      RECT 12.165 -48.51 12.515 -48.39 ;
      RECT 12.165 -45.28 12.515 -45.16 ;
      RECT 12.165 -42.05 12.515 -41.93 ;
      RECT 12.165 -38.82 12.515 -38.7 ;
      RECT 12.165 -35.59 12.515 -35.47 ;
      RECT 12.165 -32.36 12.515 -32.24 ;
      RECT 12.165 -29.13 12.515 -29.01 ;
      RECT 12.165 -25.9 12.515 -25.78 ;
      RECT 12.165 -22.67 12.515 -22.55 ;
      RECT 12.165 -19.44 12.515 -19.32 ;
      RECT 12.165 -16.21 12.515 -16.09 ;
      RECT 12.165 -12.98 12.515 -12.86 ;
      RECT 12.165 -9.75 12.515 -9.63 ;
      RECT 12.165 -6.52 12.515 -6.4 ;
      RECT 12.165 -3.29 12.515 -3.17 ;
      RECT 12.165 -0.06 12.515 0.06 ;
      RECT 12.335 -104.945 12.435 -103.985 ;
      RECT 12.335 2.175 12.435 3.135 ;
      RECT 12.16 -109.595 12.305 -109.275 ;
      RECT 12.075 -104.945 12.175 -103.985 ;
      RECT 11.95 -101.06 12.05 -100.525 ;
      RECT 11.95 -99.735 12.05 -99.2 ;
      RECT 11.95 -97.83 12.05 -97.295 ;
      RECT 11.95 -96.505 12.05 -95.97 ;
      RECT 11.95 -94.6 12.05 -94.065 ;
      RECT 11.95 -93.275 12.05 -92.74 ;
      RECT 11.95 -91.37 12.05 -90.835 ;
      RECT 11.95 -90.045 12.05 -89.51 ;
      RECT 11.95 -88.14 12.05 -87.605 ;
      RECT 11.95 -86.815 12.05 -86.28 ;
      RECT 11.95 -84.91 12.05 -84.375 ;
      RECT 11.95 -83.585 12.05 -83.05 ;
      RECT 11.95 -81.68 12.05 -81.145 ;
      RECT 11.95 -80.355 12.05 -79.82 ;
      RECT 11.95 -78.45 12.05 -77.915 ;
      RECT 11.95 -77.125 12.05 -76.59 ;
      RECT 11.95 -75.22 12.05 -74.685 ;
      RECT 11.95 -73.895 12.05 -73.36 ;
      RECT 11.95 -71.99 12.05 -71.455 ;
      RECT 11.95 -70.665 12.05 -70.13 ;
      RECT 11.95 -68.76 12.05 -68.225 ;
      RECT 11.95 -67.435 12.05 -66.9 ;
      RECT 11.95 -65.53 12.05 -64.995 ;
      RECT 11.95 -64.205 12.05 -63.67 ;
      RECT 11.95 -62.3 12.05 -61.765 ;
      RECT 11.95 -60.975 12.05 -60.44 ;
      RECT 11.95 -59.07 12.05 -58.535 ;
      RECT 11.95 -57.745 12.05 -57.21 ;
      RECT 11.95 -55.84 12.05 -55.305 ;
      RECT 11.95 -54.515 12.05 -53.98 ;
      RECT 11.95 -52.61 12.05 -52.075 ;
      RECT 11.95 -51.285 12.05 -50.75 ;
      RECT 11.95 -49.38 12.05 -48.845 ;
      RECT 11.95 -48.055 12.05 -47.52 ;
      RECT 11.95 -46.15 12.05 -45.615 ;
      RECT 11.95 -44.825 12.05 -44.29 ;
      RECT 11.95 -42.92 12.05 -42.385 ;
      RECT 11.95 -41.595 12.05 -41.06 ;
      RECT 11.95 -39.69 12.05 -39.155 ;
      RECT 11.95 -38.365 12.05 -37.83 ;
      RECT 11.95 -36.46 12.05 -35.925 ;
      RECT 11.95 -35.135 12.05 -34.6 ;
      RECT 11.95 -33.23 12.05 -32.695 ;
      RECT 11.95 -31.905 12.05 -31.37 ;
      RECT 11.95 -30 12.05 -29.465 ;
      RECT 11.95 -28.675 12.05 -28.14 ;
      RECT 11.95 -26.77 12.05 -26.235 ;
      RECT 11.95 -25.445 12.05 -24.91 ;
      RECT 11.95 -23.54 12.05 -23.005 ;
      RECT 11.95 -22.215 12.05 -21.68 ;
      RECT 11.95 -20.31 12.05 -19.775 ;
      RECT 11.95 -18.985 12.05 -18.45 ;
      RECT 11.95 -17.08 12.05 -16.545 ;
      RECT 11.95 -15.755 12.05 -15.22 ;
      RECT 11.95 -13.85 12.05 -13.315 ;
      RECT 11.95 -12.525 12.05 -11.99 ;
      RECT 11.95 -10.62 12.05 -10.085 ;
      RECT 11.95 -9.295 12.05 -8.76 ;
      RECT 11.95 -7.39 12.05 -6.855 ;
      RECT 11.95 -6.065 12.05 -5.53 ;
      RECT 11.95 -4.16 12.05 -3.625 ;
      RECT 11.95 -2.835 12.05 -2.3 ;
      RECT 11.95 -0.93 12.05 -0.395 ;
      RECT 11.95 0.395 12.05 0.93 ;
      RECT 11.825 -108.175 11.925 -107.215 ;
      RECT 11.45 -100.19 11.8 -100.07 ;
      RECT 11.45 -96.96 11.8 -96.84 ;
      RECT 11.45 -93.73 11.8 -93.61 ;
      RECT 11.45 -90.5 11.8 -90.38 ;
      RECT 11.45 -87.27 11.8 -87.15 ;
      RECT 11.45 -84.04 11.8 -83.92 ;
      RECT 11.45 -80.81 11.8 -80.69 ;
      RECT 11.45 -77.58 11.8 -77.46 ;
      RECT 11.45 -74.35 11.8 -74.23 ;
      RECT 11.45 -71.12 11.8 -71 ;
      RECT 11.45 -67.89 11.8 -67.77 ;
      RECT 11.45 -64.66 11.8 -64.54 ;
      RECT 11.45 -61.43 11.8 -61.31 ;
      RECT 11.45 -58.2 11.8 -58.08 ;
      RECT 11.45 -54.97 11.8 -54.85 ;
      RECT 11.45 -51.74 11.8 -51.62 ;
      RECT 11.45 -48.51 11.8 -48.39 ;
      RECT 11.45 -45.28 11.8 -45.16 ;
      RECT 11.45 -42.05 11.8 -41.93 ;
      RECT 11.45 -38.82 11.8 -38.7 ;
      RECT 11.45 -35.59 11.8 -35.47 ;
      RECT 11.45 -32.36 11.8 -32.24 ;
      RECT 11.45 -29.13 11.8 -29.01 ;
      RECT 11.45 -25.9 11.8 -25.78 ;
      RECT 11.45 -22.67 11.8 -22.55 ;
      RECT 11.45 -19.44 11.8 -19.32 ;
      RECT 11.45 -16.21 11.8 -16.09 ;
      RECT 11.45 -12.98 11.8 -12.86 ;
      RECT 11.45 -9.75 11.8 -9.63 ;
      RECT 11.45 -6.52 11.8 -6.4 ;
      RECT 11.45 -3.29 11.8 -3.17 ;
      RECT 11.45 -0.06 11.8 0.06 ;
      RECT 11.655 -112.255 11.755 -111.775 ;
      RECT 11.655 -110.765 11.755 -110.295 ;
      RECT 11.565 -108.175 11.665 -107.215 ;
      RECT 11.565 2.175 11.665 3.135 ;
      RECT 10.965 -100.19 11.315 -100.07 ;
      RECT 10.965 -96.96 11.315 -96.84 ;
      RECT 10.965 -93.73 11.315 -93.61 ;
      RECT 10.965 -90.5 11.315 -90.38 ;
      RECT 10.965 -87.27 11.315 -87.15 ;
      RECT 10.965 -84.04 11.315 -83.92 ;
      RECT 10.965 -80.81 11.315 -80.69 ;
      RECT 10.965 -77.58 11.315 -77.46 ;
      RECT 10.965 -74.35 11.315 -74.23 ;
      RECT 10.965 -71.12 11.315 -71 ;
      RECT 10.965 -67.89 11.315 -67.77 ;
      RECT 10.965 -64.66 11.315 -64.54 ;
      RECT 10.965 -61.43 11.315 -61.31 ;
      RECT 10.965 -58.2 11.315 -58.08 ;
      RECT 10.965 -54.97 11.315 -54.85 ;
      RECT 10.965 -51.74 11.315 -51.62 ;
      RECT 10.965 -48.51 11.315 -48.39 ;
      RECT 10.965 -45.28 11.315 -45.16 ;
      RECT 10.965 -42.05 11.315 -41.93 ;
      RECT 10.965 -38.82 11.315 -38.7 ;
      RECT 10.965 -35.59 11.315 -35.47 ;
      RECT 10.965 -32.36 11.315 -32.24 ;
      RECT 10.965 -29.13 11.315 -29.01 ;
      RECT 10.965 -25.9 11.315 -25.78 ;
      RECT 10.965 -22.67 11.315 -22.55 ;
      RECT 10.965 -19.44 11.315 -19.32 ;
      RECT 10.965 -16.21 11.315 -16.09 ;
      RECT 10.965 -12.98 11.315 -12.86 ;
      RECT 10.965 -9.75 11.315 -9.63 ;
      RECT 10.965 -6.52 11.315 -6.4 ;
      RECT 10.965 -3.29 11.315 -3.17 ;
      RECT 10.965 -0.06 11.315 0.06 ;
      RECT 11.135 -108.175 11.235 -107.215 ;
      RECT 11.135 2.175 11.235 3.135 ;
      RECT 11.03 -110.765 11.2 -110.385 ;
      RECT 11.065 -112.245 11.165 -111.775 ;
      RECT 10.875 -108.175 10.975 -107.215 ;
      RECT 10.75 -101.06 10.85 -100.525 ;
      RECT 10.75 -99.735 10.85 -99.2 ;
      RECT 10.75 -97.83 10.85 -97.295 ;
      RECT 10.75 -96.505 10.85 -95.97 ;
      RECT 10.75 -94.6 10.85 -94.065 ;
      RECT 10.75 -93.275 10.85 -92.74 ;
      RECT 10.75 -91.37 10.85 -90.835 ;
      RECT 10.75 -90.045 10.85 -89.51 ;
      RECT 10.75 -88.14 10.85 -87.605 ;
      RECT 10.75 -86.815 10.85 -86.28 ;
      RECT 10.75 -84.91 10.85 -84.375 ;
      RECT 10.75 -83.585 10.85 -83.05 ;
      RECT 10.75 -81.68 10.85 -81.145 ;
      RECT 10.75 -80.355 10.85 -79.82 ;
      RECT 10.75 -78.45 10.85 -77.915 ;
      RECT 10.75 -77.125 10.85 -76.59 ;
      RECT 10.75 -75.22 10.85 -74.685 ;
      RECT 10.75 -73.895 10.85 -73.36 ;
      RECT 10.75 -71.99 10.85 -71.455 ;
      RECT 10.75 -70.665 10.85 -70.13 ;
      RECT 10.75 -68.76 10.85 -68.225 ;
      RECT 10.75 -67.435 10.85 -66.9 ;
      RECT 10.75 -65.53 10.85 -64.995 ;
      RECT 10.75 -64.205 10.85 -63.67 ;
      RECT 10.75 -62.3 10.85 -61.765 ;
      RECT 10.75 -60.975 10.85 -60.44 ;
      RECT 10.75 -59.07 10.85 -58.535 ;
      RECT 10.75 -57.745 10.85 -57.21 ;
      RECT 10.75 -55.84 10.85 -55.305 ;
      RECT 10.75 -54.515 10.85 -53.98 ;
      RECT 10.75 -52.61 10.85 -52.075 ;
      RECT 10.75 -51.285 10.85 -50.75 ;
      RECT 10.75 -49.38 10.85 -48.845 ;
      RECT 10.75 -48.055 10.85 -47.52 ;
      RECT 10.75 -46.15 10.85 -45.615 ;
      RECT 10.75 -44.825 10.85 -44.29 ;
      RECT 10.75 -42.92 10.85 -42.385 ;
      RECT 10.75 -41.595 10.85 -41.06 ;
      RECT 10.75 -39.69 10.85 -39.155 ;
      RECT 10.75 -38.365 10.85 -37.83 ;
      RECT 10.75 -36.46 10.85 -35.925 ;
      RECT 10.75 -35.135 10.85 -34.6 ;
      RECT 10.75 -33.23 10.85 -32.695 ;
      RECT 10.75 -31.905 10.85 -31.37 ;
      RECT 10.75 -30 10.85 -29.465 ;
      RECT 10.75 -28.675 10.85 -28.14 ;
      RECT 10.75 -26.77 10.85 -26.235 ;
      RECT 10.75 -25.445 10.85 -24.91 ;
      RECT 10.75 -23.54 10.85 -23.005 ;
      RECT 10.75 -22.215 10.85 -21.68 ;
      RECT 10.75 -20.31 10.85 -19.775 ;
      RECT 10.75 -18.985 10.85 -18.45 ;
      RECT 10.75 -17.08 10.85 -16.545 ;
      RECT 10.75 -15.755 10.85 -15.22 ;
      RECT 10.75 -13.85 10.85 -13.315 ;
      RECT 10.75 -12.525 10.85 -11.99 ;
      RECT 10.75 -10.62 10.85 -10.085 ;
      RECT 10.75 -9.295 10.85 -8.76 ;
      RECT 10.75 -7.39 10.85 -6.855 ;
      RECT 10.75 -6.065 10.85 -5.53 ;
      RECT 10.75 -4.16 10.85 -3.625 ;
      RECT 10.75 -2.835 10.85 -2.3 ;
      RECT 10.75 -0.93 10.85 -0.395 ;
      RECT 10.75 0.395 10.85 0.93 ;
      RECT 10.625 -108.175 10.725 -107.215 ;
      RECT 10.25 -100.19 10.6 -100.07 ;
      RECT 10.25 -96.96 10.6 -96.84 ;
      RECT 10.25 -93.73 10.6 -93.61 ;
      RECT 10.25 -90.5 10.6 -90.38 ;
      RECT 10.25 -87.27 10.6 -87.15 ;
      RECT 10.25 -84.04 10.6 -83.92 ;
      RECT 10.25 -80.81 10.6 -80.69 ;
      RECT 10.25 -77.58 10.6 -77.46 ;
      RECT 10.25 -74.35 10.6 -74.23 ;
      RECT 10.25 -71.12 10.6 -71 ;
      RECT 10.25 -67.89 10.6 -67.77 ;
      RECT 10.25 -64.66 10.6 -64.54 ;
      RECT 10.25 -61.43 10.6 -61.31 ;
      RECT 10.25 -58.2 10.6 -58.08 ;
      RECT 10.25 -54.97 10.6 -54.85 ;
      RECT 10.25 -51.74 10.6 -51.62 ;
      RECT 10.25 -48.51 10.6 -48.39 ;
      RECT 10.25 -45.28 10.6 -45.16 ;
      RECT 10.25 -42.05 10.6 -41.93 ;
      RECT 10.25 -38.82 10.6 -38.7 ;
      RECT 10.25 -35.59 10.6 -35.47 ;
      RECT 10.25 -32.36 10.6 -32.24 ;
      RECT 10.25 -29.13 10.6 -29.01 ;
      RECT 10.25 -25.9 10.6 -25.78 ;
      RECT 10.25 -22.67 10.6 -22.55 ;
      RECT 10.25 -19.44 10.6 -19.32 ;
      RECT 10.25 -16.21 10.6 -16.09 ;
      RECT 10.25 -12.98 10.6 -12.86 ;
      RECT 10.25 -9.75 10.6 -9.63 ;
      RECT 10.25 -6.52 10.6 -6.4 ;
      RECT 10.25 -3.29 10.6 -3.17 ;
      RECT 10.25 -0.06 10.6 0.06 ;
      RECT 10.365 -108.175 10.465 -107.215 ;
      RECT 10.365 2.175 10.465 3.135 ;
      RECT 10.265 -113.555 10.365 -113.085 ;
      RECT 9.765 -100.19 10.115 -100.07 ;
      RECT 9.765 -96.96 10.115 -96.84 ;
      RECT 9.765 -93.73 10.115 -93.61 ;
      RECT 9.765 -90.5 10.115 -90.38 ;
      RECT 9.765 -87.27 10.115 -87.15 ;
      RECT 9.765 -84.04 10.115 -83.92 ;
      RECT 9.765 -80.81 10.115 -80.69 ;
      RECT 9.765 -77.58 10.115 -77.46 ;
      RECT 9.765 -74.35 10.115 -74.23 ;
      RECT 9.765 -71.12 10.115 -71 ;
      RECT 9.765 -67.89 10.115 -67.77 ;
      RECT 9.765 -64.66 10.115 -64.54 ;
      RECT 9.765 -61.43 10.115 -61.31 ;
      RECT 9.765 -58.2 10.115 -58.08 ;
      RECT 9.765 -54.97 10.115 -54.85 ;
      RECT 9.765 -51.74 10.115 -51.62 ;
      RECT 9.765 -48.51 10.115 -48.39 ;
      RECT 9.765 -45.28 10.115 -45.16 ;
      RECT 9.765 -42.05 10.115 -41.93 ;
      RECT 9.765 -38.82 10.115 -38.7 ;
      RECT 9.765 -35.59 10.115 -35.47 ;
      RECT 9.765 -32.36 10.115 -32.24 ;
      RECT 9.765 -29.13 10.115 -29.01 ;
      RECT 9.765 -25.9 10.115 -25.78 ;
      RECT 9.765 -22.67 10.115 -22.55 ;
      RECT 9.765 -19.44 10.115 -19.32 ;
      RECT 9.765 -16.21 10.115 -16.09 ;
      RECT 9.765 -12.98 10.115 -12.86 ;
      RECT 9.765 -9.75 10.115 -9.63 ;
      RECT 9.765 -6.52 10.115 -6.4 ;
      RECT 9.765 -3.29 10.115 -3.17 ;
      RECT 9.765 -0.06 10.115 0.06 ;
      RECT 9.9 -110.735 10.05 -110.445 ;
      RECT 9.935 -108.175 10.035 -107.215 ;
      RECT 9.935 2.175 10.035 3.135 ;
      RECT 9.915 -112.19 10.015 -111.65 ;
      RECT 9.675 -113.555 9.775 -113.085 ;
      RECT 9.675 -108.175 9.775 -107.215 ;
      RECT 9.55 -101.06 9.65 -100.525 ;
      RECT 9.55 -99.735 9.65 -99.2 ;
      RECT 9.55 -97.83 9.65 -97.295 ;
      RECT 9.55 -96.505 9.65 -95.97 ;
      RECT 9.55 -94.6 9.65 -94.065 ;
      RECT 9.55 -93.275 9.65 -92.74 ;
      RECT 9.55 -91.37 9.65 -90.835 ;
      RECT 9.55 -90.045 9.65 -89.51 ;
      RECT 9.55 -88.14 9.65 -87.605 ;
      RECT 9.55 -86.815 9.65 -86.28 ;
      RECT 9.55 -84.91 9.65 -84.375 ;
      RECT 9.55 -83.585 9.65 -83.05 ;
      RECT 9.55 -81.68 9.65 -81.145 ;
      RECT 9.55 -80.355 9.65 -79.82 ;
      RECT 9.55 -78.45 9.65 -77.915 ;
      RECT 9.55 -77.125 9.65 -76.59 ;
      RECT 9.55 -75.22 9.65 -74.685 ;
      RECT 9.55 -73.895 9.65 -73.36 ;
      RECT 9.55 -71.99 9.65 -71.455 ;
      RECT 9.55 -70.665 9.65 -70.13 ;
      RECT 9.55 -68.76 9.65 -68.225 ;
      RECT 9.55 -67.435 9.65 -66.9 ;
      RECT 9.55 -65.53 9.65 -64.995 ;
      RECT 9.55 -64.205 9.65 -63.67 ;
      RECT 9.55 -62.3 9.65 -61.765 ;
      RECT 9.55 -60.975 9.65 -60.44 ;
      RECT 9.55 -59.07 9.65 -58.535 ;
      RECT 9.55 -57.745 9.65 -57.21 ;
      RECT 9.55 -55.84 9.65 -55.305 ;
      RECT 9.55 -54.515 9.65 -53.98 ;
      RECT 9.55 -52.61 9.65 -52.075 ;
      RECT 9.55 -51.285 9.65 -50.75 ;
      RECT 9.55 -49.38 9.65 -48.845 ;
      RECT 9.55 -48.055 9.65 -47.52 ;
      RECT 9.55 -46.15 9.65 -45.615 ;
      RECT 9.55 -44.825 9.65 -44.29 ;
      RECT 9.55 -42.92 9.65 -42.385 ;
      RECT 9.55 -41.595 9.65 -41.06 ;
      RECT 9.55 -39.69 9.65 -39.155 ;
      RECT 9.55 -38.365 9.65 -37.83 ;
      RECT 9.55 -36.46 9.65 -35.925 ;
      RECT 9.55 -35.135 9.65 -34.6 ;
      RECT 9.55 -33.23 9.65 -32.695 ;
      RECT 9.55 -31.905 9.65 -31.37 ;
      RECT 9.55 -30 9.65 -29.465 ;
      RECT 9.55 -28.675 9.65 -28.14 ;
      RECT 9.55 -26.77 9.65 -26.235 ;
      RECT 9.55 -25.445 9.65 -24.91 ;
      RECT 9.55 -23.54 9.65 -23.005 ;
      RECT 9.55 -22.215 9.65 -21.68 ;
      RECT 9.55 -20.31 9.65 -19.775 ;
      RECT 9.55 -18.985 9.65 -18.45 ;
      RECT 9.55 -17.08 9.65 -16.545 ;
      RECT 9.55 -15.755 9.65 -15.22 ;
      RECT 9.55 -13.85 9.65 -13.315 ;
      RECT 9.55 -12.525 9.65 -11.99 ;
      RECT 9.55 -10.62 9.65 -10.085 ;
      RECT 9.55 -9.295 9.65 -8.76 ;
      RECT 9.55 -7.39 9.65 -6.855 ;
      RECT 9.55 -6.065 9.65 -5.53 ;
      RECT 9.55 -4.16 9.65 -3.625 ;
      RECT 9.55 -2.835 9.65 -2.3 ;
      RECT 9.55 -0.93 9.65 -0.395 ;
      RECT 9.55 0.395 9.65 0.93 ;
      RECT 9.425 -104.945 9.525 -103.985 ;
      RECT 9.05 -100.19 9.4 -100.07 ;
      RECT 9.05 -96.96 9.4 -96.84 ;
      RECT 9.05 -93.73 9.4 -93.61 ;
      RECT 9.05 -90.5 9.4 -90.38 ;
      RECT 9.05 -87.27 9.4 -87.15 ;
      RECT 9.05 -84.04 9.4 -83.92 ;
      RECT 9.05 -80.81 9.4 -80.69 ;
      RECT 9.05 -77.58 9.4 -77.46 ;
      RECT 9.05 -74.35 9.4 -74.23 ;
      RECT 9.05 -71.12 9.4 -71 ;
      RECT 9.05 -67.89 9.4 -67.77 ;
      RECT 9.05 -64.66 9.4 -64.54 ;
      RECT 9.05 -61.43 9.4 -61.31 ;
      RECT 9.05 -58.2 9.4 -58.08 ;
      RECT 9.05 -54.97 9.4 -54.85 ;
      RECT 9.05 -51.74 9.4 -51.62 ;
      RECT 9.05 -48.51 9.4 -48.39 ;
      RECT 9.05 -45.28 9.4 -45.16 ;
      RECT 9.05 -42.05 9.4 -41.93 ;
      RECT 9.05 -38.82 9.4 -38.7 ;
      RECT 9.05 -35.59 9.4 -35.47 ;
      RECT 9.05 -32.36 9.4 -32.24 ;
      RECT 9.05 -29.13 9.4 -29.01 ;
      RECT 9.05 -25.9 9.4 -25.78 ;
      RECT 9.05 -22.67 9.4 -22.55 ;
      RECT 9.05 -19.44 9.4 -19.32 ;
      RECT 9.05 -16.21 9.4 -16.09 ;
      RECT 9.05 -12.98 9.4 -12.86 ;
      RECT 9.05 -9.75 9.4 -9.63 ;
      RECT 9.05 -6.52 9.4 -6.4 ;
      RECT 9.05 -3.29 9.4 -3.17 ;
      RECT 9.05 -0.06 9.4 0.06 ;
      RECT 9.165 -104.945 9.265 -103.985 ;
      RECT 9.165 2.175 9.265 3.135 ;
      RECT 8.875 -112.255 8.975 -111.775 ;
      RECT 8.875 -110.765 8.975 -110.295 ;
      RECT 8.565 -100.19 8.915 -100.07 ;
      RECT 8.565 -96.96 8.915 -96.84 ;
      RECT 8.565 -93.73 8.915 -93.61 ;
      RECT 8.565 -90.5 8.915 -90.38 ;
      RECT 8.565 -87.27 8.915 -87.15 ;
      RECT 8.565 -84.04 8.915 -83.92 ;
      RECT 8.565 -80.81 8.915 -80.69 ;
      RECT 8.565 -77.58 8.915 -77.46 ;
      RECT 8.565 -74.35 8.915 -74.23 ;
      RECT 8.565 -71.12 8.915 -71 ;
      RECT 8.565 -67.89 8.915 -67.77 ;
      RECT 8.565 -64.66 8.915 -64.54 ;
      RECT 8.565 -61.43 8.915 -61.31 ;
      RECT 8.565 -58.2 8.915 -58.08 ;
      RECT 8.565 -54.97 8.915 -54.85 ;
      RECT 8.565 -51.74 8.915 -51.62 ;
      RECT 8.565 -48.51 8.915 -48.39 ;
      RECT 8.565 -45.28 8.915 -45.16 ;
      RECT 8.565 -42.05 8.915 -41.93 ;
      RECT 8.565 -38.82 8.915 -38.7 ;
      RECT 8.565 -35.59 8.915 -35.47 ;
      RECT 8.565 -32.36 8.915 -32.24 ;
      RECT 8.565 -29.13 8.915 -29.01 ;
      RECT 8.565 -25.9 8.915 -25.78 ;
      RECT 8.565 -22.67 8.915 -22.55 ;
      RECT 8.565 -19.44 8.915 -19.32 ;
      RECT 8.565 -16.21 8.915 -16.09 ;
      RECT 8.565 -12.98 8.915 -12.86 ;
      RECT 8.565 -9.75 8.915 -9.63 ;
      RECT 8.565 -6.52 8.915 -6.4 ;
      RECT 8.565 -3.29 8.915 -3.17 ;
      RECT 8.565 -0.06 8.915 0.06 ;
      RECT 8.735 -104.945 8.835 -103.985 ;
      RECT 8.735 2.175 8.835 3.135 ;
      RECT 4.835 -108.655 8.615 -108.535 ;
      RECT 8.475 -104.945 8.575 -103.985 ;
      RECT 8.35 -101.06 8.45 -100.525 ;
      RECT 8.35 -99.735 8.45 -99.2 ;
      RECT 8.35 -97.83 8.45 -97.295 ;
      RECT 8.35 -96.505 8.45 -95.97 ;
      RECT 8.35 -94.6 8.45 -94.065 ;
      RECT 8.35 -93.275 8.45 -92.74 ;
      RECT 8.35 -91.37 8.45 -90.835 ;
      RECT 8.35 -90.045 8.45 -89.51 ;
      RECT 8.35 -88.14 8.45 -87.605 ;
      RECT 8.35 -86.815 8.45 -86.28 ;
      RECT 8.35 -84.91 8.45 -84.375 ;
      RECT 8.35 -83.585 8.45 -83.05 ;
      RECT 8.35 -81.68 8.45 -81.145 ;
      RECT 8.35 -80.355 8.45 -79.82 ;
      RECT 8.35 -78.45 8.45 -77.915 ;
      RECT 8.35 -77.125 8.45 -76.59 ;
      RECT 8.35 -75.22 8.45 -74.685 ;
      RECT 8.35 -73.895 8.45 -73.36 ;
      RECT 8.35 -71.99 8.45 -71.455 ;
      RECT 8.35 -70.665 8.45 -70.13 ;
      RECT 8.35 -68.76 8.45 -68.225 ;
      RECT 8.35 -67.435 8.45 -66.9 ;
      RECT 8.35 -65.53 8.45 -64.995 ;
      RECT 8.35 -64.205 8.45 -63.67 ;
      RECT 8.35 -62.3 8.45 -61.765 ;
      RECT 8.35 -60.975 8.45 -60.44 ;
      RECT 8.35 -59.07 8.45 -58.535 ;
      RECT 8.35 -57.745 8.45 -57.21 ;
      RECT 8.35 -55.84 8.45 -55.305 ;
      RECT 8.35 -54.515 8.45 -53.98 ;
      RECT 8.35 -52.61 8.45 -52.075 ;
      RECT 8.35 -51.285 8.45 -50.75 ;
      RECT 8.35 -49.38 8.45 -48.845 ;
      RECT 8.35 -48.055 8.45 -47.52 ;
      RECT 8.35 -46.15 8.45 -45.615 ;
      RECT 8.35 -44.825 8.45 -44.29 ;
      RECT 8.35 -42.92 8.45 -42.385 ;
      RECT 8.35 -41.595 8.45 -41.06 ;
      RECT 8.35 -39.69 8.45 -39.155 ;
      RECT 8.35 -38.365 8.45 -37.83 ;
      RECT 8.35 -36.46 8.45 -35.925 ;
      RECT 8.35 -35.135 8.45 -34.6 ;
      RECT 8.35 -33.23 8.45 -32.695 ;
      RECT 8.35 -31.905 8.45 -31.37 ;
      RECT 8.35 -30 8.45 -29.465 ;
      RECT 8.35 -28.675 8.45 -28.14 ;
      RECT 8.35 -26.77 8.45 -26.235 ;
      RECT 8.35 -25.445 8.45 -24.91 ;
      RECT 8.35 -23.54 8.45 -23.005 ;
      RECT 8.35 -22.215 8.45 -21.68 ;
      RECT 8.35 -20.31 8.45 -19.775 ;
      RECT 8.35 -18.985 8.45 -18.45 ;
      RECT 8.35 -17.08 8.45 -16.545 ;
      RECT 8.35 -15.755 8.45 -15.22 ;
      RECT 8.35 -13.85 8.45 -13.315 ;
      RECT 8.35 -12.525 8.45 -11.99 ;
      RECT 8.35 -10.62 8.45 -10.085 ;
      RECT 8.35 -9.295 8.45 -8.76 ;
      RECT 8.35 -7.39 8.45 -6.855 ;
      RECT 8.35 -6.065 8.45 -5.53 ;
      RECT 8.35 -4.16 8.45 -3.625 ;
      RECT 8.35 -2.835 8.45 -2.3 ;
      RECT 8.35 -0.93 8.45 -0.395 ;
      RECT 8.35 0.395 8.45 0.93 ;
      RECT 8.285 -110.75 8.405 -110.37 ;
      RECT 8.285 -112.245 8.385 -111.775 ;
      RECT 8.225 -104.945 8.325 -103.985 ;
      RECT 7.85 -100.19 8.2 -100.07 ;
      RECT 7.85 -96.96 8.2 -96.84 ;
      RECT 7.85 -93.73 8.2 -93.61 ;
      RECT 7.85 -90.5 8.2 -90.38 ;
      RECT 7.85 -87.27 8.2 -87.15 ;
      RECT 7.85 -84.04 8.2 -83.92 ;
      RECT 7.85 -80.81 8.2 -80.69 ;
      RECT 7.85 -77.58 8.2 -77.46 ;
      RECT 7.85 -74.35 8.2 -74.23 ;
      RECT 7.85 -71.12 8.2 -71 ;
      RECT 7.85 -67.89 8.2 -67.77 ;
      RECT 7.85 -64.66 8.2 -64.54 ;
      RECT 7.85 -61.43 8.2 -61.31 ;
      RECT 7.85 -58.2 8.2 -58.08 ;
      RECT 7.85 -54.97 8.2 -54.85 ;
      RECT 7.85 -51.74 8.2 -51.62 ;
      RECT 7.85 -48.51 8.2 -48.39 ;
      RECT 7.85 -45.28 8.2 -45.16 ;
      RECT 7.85 -42.05 8.2 -41.93 ;
      RECT 7.85 -38.82 8.2 -38.7 ;
      RECT 7.85 -35.59 8.2 -35.47 ;
      RECT 7.85 -32.36 8.2 -32.24 ;
      RECT 7.85 -29.13 8.2 -29.01 ;
      RECT 7.85 -25.9 8.2 -25.78 ;
      RECT 7.85 -22.67 8.2 -22.55 ;
      RECT 7.85 -19.44 8.2 -19.32 ;
      RECT 7.85 -16.21 8.2 -16.09 ;
      RECT 7.85 -12.98 8.2 -12.86 ;
      RECT 7.85 -9.75 8.2 -9.63 ;
      RECT 7.85 -6.52 8.2 -6.4 ;
      RECT 7.85 -3.29 8.2 -3.17 ;
      RECT 7.85 -0.06 8.2 0.06 ;
      RECT 7.965 -104.945 8.065 -103.985 ;
      RECT 7.965 2.175 8.065 3.135 ;
      RECT 7.695 -109.595 7.83 -109.275 ;
      RECT 7.365 -100.19 7.715 -100.07 ;
      RECT 7.365 -96.96 7.715 -96.84 ;
      RECT 7.365 -93.73 7.715 -93.61 ;
      RECT 7.365 -90.5 7.715 -90.38 ;
      RECT 7.365 -87.27 7.715 -87.15 ;
      RECT 7.365 -84.04 7.715 -83.92 ;
      RECT 7.365 -80.81 7.715 -80.69 ;
      RECT 7.365 -77.58 7.715 -77.46 ;
      RECT 7.365 -74.35 7.715 -74.23 ;
      RECT 7.365 -71.12 7.715 -71 ;
      RECT 7.365 -67.89 7.715 -67.77 ;
      RECT 7.365 -64.66 7.715 -64.54 ;
      RECT 7.365 -61.43 7.715 -61.31 ;
      RECT 7.365 -58.2 7.715 -58.08 ;
      RECT 7.365 -54.97 7.715 -54.85 ;
      RECT 7.365 -51.74 7.715 -51.62 ;
      RECT 7.365 -48.51 7.715 -48.39 ;
      RECT 7.365 -45.28 7.715 -45.16 ;
      RECT 7.365 -42.05 7.715 -41.93 ;
      RECT 7.365 -38.82 7.715 -38.7 ;
      RECT 7.365 -35.59 7.715 -35.47 ;
      RECT 7.365 -32.36 7.715 -32.24 ;
      RECT 7.365 -29.13 7.715 -29.01 ;
      RECT 7.365 -25.9 7.715 -25.78 ;
      RECT 7.365 -22.67 7.715 -22.55 ;
      RECT 7.365 -19.44 7.715 -19.32 ;
      RECT 7.365 -16.21 7.715 -16.09 ;
      RECT 7.365 -12.98 7.715 -12.86 ;
      RECT 7.365 -9.75 7.715 -9.63 ;
      RECT 7.365 -6.52 7.715 -6.4 ;
      RECT 7.365 -3.29 7.715 -3.17 ;
      RECT 7.365 -0.06 7.715 0.06 ;
      RECT 7.535 -104.945 7.635 -103.985 ;
      RECT 7.535 2.175 7.635 3.135 ;
      RECT 7.36 -109.595 7.505 -109.275 ;
      RECT 7.275 -104.945 7.375 -103.985 ;
      RECT 7.15 -101.06 7.25 -100.525 ;
      RECT 7.15 -99.735 7.25 -99.2 ;
      RECT 7.15 -97.83 7.25 -97.295 ;
      RECT 7.15 -96.505 7.25 -95.97 ;
      RECT 7.15 -94.6 7.25 -94.065 ;
      RECT 7.15 -93.275 7.25 -92.74 ;
      RECT 7.15 -91.37 7.25 -90.835 ;
      RECT 7.15 -90.045 7.25 -89.51 ;
      RECT 7.15 -88.14 7.25 -87.605 ;
      RECT 7.15 -86.815 7.25 -86.28 ;
      RECT 7.15 -84.91 7.25 -84.375 ;
      RECT 7.15 -83.585 7.25 -83.05 ;
      RECT 7.15 -81.68 7.25 -81.145 ;
      RECT 7.15 -80.355 7.25 -79.82 ;
      RECT 7.15 -78.45 7.25 -77.915 ;
      RECT 7.15 -77.125 7.25 -76.59 ;
      RECT 7.15 -75.22 7.25 -74.685 ;
      RECT 7.15 -73.895 7.25 -73.36 ;
      RECT 7.15 -71.99 7.25 -71.455 ;
      RECT 7.15 -70.665 7.25 -70.13 ;
      RECT 7.15 -68.76 7.25 -68.225 ;
      RECT 7.15 -67.435 7.25 -66.9 ;
      RECT 7.15 -65.53 7.25 -64.995 ;
      RECT 7.15 -64.205 7.25 -63.67 ;
      RECT 7.15 -62.3 7.25 -61.765 ;
      RECT 7.15 -60.975 7.25 -60.44 ;
      RECT 7.15 -59.07 7.25 -58.535 ;
      RECT 7.15 -57.745 7.25 -57.21 ;
      RECT 7.15 -55.84 7.25 -55.305 ;
      RECT 7.15 -54.515 7.25 -53.98 ;
      RECT 7.15 -52.61 7.25 -52.075 ;
      RECT 7.15 -51.285 7.25 -50.75 ;
      RECT 7.15 -49.38 7.25 -48.845 ;
      RECT 7.15 -48.055 7.25 -47.52 ;
      RECT 7.15 -46.15 7.25 -45.615 ;
      RECT 7.15 -44.825 7.25 -44.29 ;
      RECT 7.15 -42.92 7.25 -42.385 ;
      RECT 7.15 -41.595 7.25 -41.06 ;
      RECT 7.15 -39.69 7.25 -39.155 ;
      RECT 7.15 -38.365 7.25 -37.83 ;
      RECT 7.15 -36.46 7.25 -35.925 ;
      RECT 7.15 -35.135 7.25 -34.6 ;
      RECT 7.15 -33.23 7.25 -32.695 ;
      RECT 7.15 -31.905 7.25 -31.37 ;
      RECT 7.15 -30 7.25 -29.465 ;
      RECT 7.15 -28.675 7.25 -28.14 ;
      RECT 7.15 -26.77 7.25 -26.235 ;
      RECT 7.15 -25.445 7.25 -24.91 ;
      RECT 7.15 -23.54 7.25 -23.005 ;
      RECT 7.15 -22.215 7.25 -21.68 ;
      RECT 7.15 -20.31 7.25 -19.775 ;
      RECT 7.15 -18.985 7.25 -18.45 ;
      RECT 7.15 -17.08 7.25 -16.545 ;
      RECT 7.15 -15.755 7.25 -15.22 ;
      RECT 7.15 -13.85 7.25 -13.315 ;
      RECT 7.15 -12.525 7.25 -11.99 ;
      RECT 7.15 -10.62 7.25 -10.085 ;
      RECT 7.15 -9.295 7.25 -8.76 ;
      RECT 7.15 -7.39 7.25 -6.855 ;
      RECT 7.15 -6.065 7.25 -5.53 ;
      RECT 7.15 -4.16 7.25 -3.625 ;
      RECT 7.15 -2.835 7.25 -2.3 ;
      RECT 7.15 -0.93 7.25 -0.395 ;
      RECT 7.15 0.395 7.25 0.93 ;
      RECT 7.025 -108.175 7.125 -107.215 ;
      RECT 6.65 -100.19 7 -100.07 ;
      RECT 6.65 -96.96 7 -96.84 ;
      RECT 6.65 -93.73 7 -93.61 ;
      RECT 6.65 -90.5 7 -90.38 ;
      RECT 6.65 -87.27 7 -87.15 ;
      RECT 6.65 -84.04 7 -83.92 ;
      RECT 6.65 -80.81 7 -80.69 ;
      RECT 6.65 -77.58 7 -77.46 ;
      RECT 6.65 -74.35 7 -74.23 ;
      RECT 6.65 -71.12 7 -71 ;
      RECT 6.65 -67.89 7 -67.77 ;
      RECT 6.65 -64.66 7 -64.54 ;
      RECT 6.65 -61.43 7 -61.31 ;
      RECT 6.65 -58.2 7 -58.08 ;
      RECT 6.65 -54.97 7 -54.85 ;
      RECT 6.65 -51.74 7 -51.62 ;
      RECT 6.65 -48.51 7 -48.39 ;
      RECT 6.65 -45.28 7 -45.16 ;
      RECT 6.65 -42.05 7 -41.93 ;
      RECT 6.65 -38.82 7 -38.7 ;
      RECT 6.65 -35.59 7 -35.47 ;
      RECT 6.65 -32.36 7 -32.24 ;
      RECT 6.65 -29.13 7 -29.01 ;
      RECT 6.65 -25.9 7 -25.78 ;
      RECT 6.65 -22.67 7 -22.55 ;
      RECT 6.65 -19.44 7 -19.32 ;
      RECT 6.65 -16.21 7 -16.09 ;
      RECT 6.65 -12.98 7 -12.86 ;
      RECT 6.65 -9.75 7 -9.63 ;
      RECT 6.65 -6.52 7 -6.4 ;
      RECT 6.65 -3.29 7 -3.17 ;
      RECT 6.65 -0.06 7 0.06 ;
      RECT 6.855 -112.255 6.955 -111.775 ;
      RECT 6.855 -110.765 6.955 -110.295 ;
      RECT 6.765 -108.175 6.865 -107.215 ;
      RECT 6.765 2.175 6.865 3.135 ;
      RECT 6.165 -100.19 6.515 -100.07 ;
      RECT 6.165 -96.96 6.515 -96.84 ;
      RECT 6.165 -93.73 6.515 -93.61 ;
      RECT 6.165 -90.5 6.515 -90.38 ;
      RECT 6.165 -87.27 6.515 -87.15 ;
      RECT 6.165 -84.04 6.515 -83.92 ;
      RECT 6.165 -80.81 6.515 -80.69 ;
      RECT 6.165 -77.58 6.515 -77.46 ;
      RECT 6.165 -74.35 6.515 -74.23 ;
      RECT 6.165 -71.12 6.515 -71 ;
      RECT 6.165 -67.89 6.515 -67.77 ;
      RECT 6.165 -64.66 6.515 -64.54 ;
      RECT 6.165 -61.43 6.515 -61.31 ;
      RECT 6.165 -58.2 6.515 -58.08 ;
      RECT 6.165 -54.97 6.515 -54.85 ;
      RECT 6.165 -51.74 6.515 -51.62 ;
      RECT 6.165 -48.51 6.515 -48.39 ;
      RECT 6.165 -45.28 6.515 -45.16 ;
      RECT 6.165 -42.05 6.515 -41.93 ;
      RECT 6.165 -38.82 6.515 -38.7 ;
      RECT 6.165 -35.59 6.515 -35.47 ;
      RECT 6.165 -32.36 6.515 -32.24 ;
      RECT 6.165 -29.13 6.515 -29.01 ;
      RECT 6.165 -25.9 6.515 -25.78 ;
      RECT 6.165 -22.67 6.515 -22.55 ;
      RECT 6.165 -19.44 6.515 -19.32 ;
      RECT 6.165 -16.21 6.515 -16.09 ;
      RECT 6.165 -12.98 6.515 -12.86 ;
      RECT 6.165 -9.75 6.515 -9.63 ;
      RECT 6.165 -6.52 6.515 -6.4 ;
      RECT 6.165 -3.29 6.515 -3.17 ;
      RECT 6.165 -0.06 6.515 0.06 ;
      RECT 6.335 -108.175 6.435 -107.215 ;
      RECT 6.335 2.175 6.435 3.135 ;
      RECT 6.23 -110.765 6.4 -110.385 ;
      RECT 6.265 -112.245 6.365 -111.775 ;
      RECT 6.075 -108.175 6.175 -107.215 ;
      RECT 5.95 -101.06 6.05 -100.525 ;
      RECT 5.95 -99.735 6.05 -99.2 ;
      RECT 5.95 -97.83 6.05 -97.295 ;
      RECT 5.95 -96.505 6.05 -95.97 ;
      RECT 5.95 -94.6 6.05 -94.065 ;
      RECT 5.95 -93.275 6.05 -92.74 ;
      RECT 5.95 -91.37 6.05 -90.835 ;
      RECT 5.95 -90.045 6.05 -89.51 ;
      RECT 5.95 -88.14 6.05 -87.605 ;
      RECT 5.95 -86.815 6.05 -86.28 ;
      RECT 5.95 -84.91 6.05 -84.375 ;
      RECT 5.95 -83.585 6.05 -83.05 ;
      RECT 5.95 -81.68 6.05 -81.145 ;
      RECT 5.95 -80.355 6.05 -79.82 ;
      RECT 5.95 -78.45 6.05 -77.915 ;
      RECT 5.95 -77.125 6.05 -76.59 ;
      RECT 5.95 -75.22 6.05 -74.685 ;
      RECT 5.95 -73.895 6.05 -73.36 ;
      RECT 5.95 -71.99 6.05 -71.455 ;
      RECT 5.95 -70.665 6.05 -70.13 ;
      RECT 5.95 -68.76 6.05 -68.225 ;
      RECT 5.95 -67.435 6.05 -66.9 ;
      RECT 5.95 -65.53 6.05 -64.995 ;
      RECT 5.95 -64.205 6.05 -63.67 ;
      RECT 5.95 -62.3 6.05 -61.765 ;
      RECT 5.95 -60.975 6.05 -60.44 ;
      RECT 5.95 -59.07 6.05 -58.535 ;
      RECT 5.95 -57.745 6.05 -57.21 ;
      RECT 5.95 -55.84 6.05 -55.305 ;
      RECT 5.95 -54.515 6.05 -53.98 ;
      RECT 5.95 -52.61 6.05 -52.075 ;
      RECT 5.95 -51.285 6.05 -50.75 ;
      RECT 5.95 -49.38 6.05 -48.845 ;
      RECT 5.95 -48.055 6.05 -47.52 ;
      RECT 5.95 -46.15 6.05 -45.615 ;
      RECT 5.95 -44.825 6.05 -44.29 ;
      RECT 5.95 -42.92 6.05 -42.385 ;
      RECT 5.95 -41.595 6.05 -41.06 ;
      RECT 5.95 -39.69 6.05 -39.155 ;
      RECT 5.95 -38.365 6.05 -37.83 ;
      RECT 5.95 -36.46 6.05 -35.925 ;
      RECT 5.95 -35.135 6.05 -34.6 ;
      RECT 5.95 -33.23 6.05 -32.695 ;
      RECT 5.95 -31.905 6.05 -31.37 ;
      RECT 5.95 -30 6.05 -29.465 ;
      RECT 5.95 -28.675 6.05 -28.14 ;
      RECT 5.95 -26.77 6.05 -26.235 ;
      RECT 5.95 -25.445 6.05 -24.91 ;
      RECT 5.95 -23.54 6.05 -23.005 ;
      RECT 5.95 -22.215 6.05 -21.68 ;
      RECT 5.95 -20.31 6.05 -19.775 ;
      RECT 5.95 -18.985 6.05 -18.45 ;
      RECT 5.95 -17.08 6.05 -16.545 ;
      RECT 5.95 -15.755 6.05 -15.22 ;
      RECT 5.95 -13.85 6.05 -13.315 ;
      RECT 5.95 -12.525 6.05 -11.99 ;
      RECT 5.95 -10.62 6.05 -10.085 ;
      RECT 5.95 -9.295 6.05 -8.76 ;
      RECT 5.95 -7.39 6.05 -6.855 ;
      RECT 5.95 -6.065 6.05 -5.53 ;
      RECT 5.95 -4.16 6.05 -3.625 ;
      RECT 5.95 -2.835 6.05 -2.3 ;
      RECT 5.95 -0.93 6.05 -0.395 ;
      RECT 5.95 0.395 6.05 0.93 ;
      RECT 5.825 -108.175 5.925 -107.215 ;
      RECT 5.45 -100.19 5.8 -100.07 ;
      RECT 5.45 -96.96 5.8 -96.84 ;
      RECT 5.45 -93.73 5.8 -93.61 ;
      RECT 5.45 -90.5 5.8 -90.38 ;
      RECT 5.45 -87.27 5.8 -87.15 ;
      RECT 5.45 -84.04 5.8 -83.92 ;
      RECT 5.45 -80.81 5.8 -80.69 ;
      RECT 5.45 -77.58 5.8 -77.46 ;
      RECT 5.45 -74.35 5.8 -74.23 ;
      RECT 5.45 -71.12 5.8 -71 ;
      RECT 5.45 -67.89 5.8 -67.77 ;
      RECT 5.45 -64.66 5.8 -64.54 ;
      RECT 5.45 -61.43 5.8 -61.31 ;
      RECT 5.45 -58.2 5.8 -58.08 ;
      RECT 5.45 -54.97 5.8 -54.85 ;
      RECT 5.45 -51.74 5.8 -51.62 ;
      RECT 5.45 -48.51 5.8 -48.39 ;
      RECT 5.45 -45.28 5.8 -45.16 ;
      RECT 5.45 -42.05 5.8 -41.93 ;
      RECT 5.45 -38.82 5.8 -38.7 ;
      RECT 5.45 -35.59 5.8 -35.47 ;
      RECT 5.45 -32.36 5.8 -32.24 ;
      RECT 5.45 -29.13 5.8 -29.01 ;
      RECT 5.45 -25.9 5.8 -25.78 ;
      RECT 5.45 -22.67 5.8 -22.55 ;
      RECT 5.45 -19.44 5.8 -19.32 ;
      RECT 5.45 -16.21 5.8 -16.09 ;
      RECT 5.45 -12.98 5.8 -12.86 ;
      RECT 5.45 -9.75 5.8 -9.63 ;
      RECT 5.45 -6.52 5.8 -6.4 ;
      RECT 5.45 -3.29 5.8 -3.17 ;
      RECT 5.45 -0.06 5.8 0.06 ;
      RECT 5.565 -108.175 5.665 -107.215 ;
      RECT 5.565 2.175 5.665 3.135 ;
      RECT 5.465 -113.555 5.565 -113.085 ;
      RECT 4.965 -100.19 5.315 -100.07 ;
      RECT 4.965 -96.96 5.315 -96.84 ;
      RECT 4.965 -93.73 5.315 -93.61 ;
      RECT 4.965 -90.5 5.315 -90.38 ;
      RECT 4.965 -87.27 5.315 -87.15 ;
      RECT 4.965 -84.04 5.315 -83.92 ;
      RECT 4.965 -80.81 5.315 -80.69 ;
      RECT 4.965 -77.58 5.315 -77.46 ;
      RECT 4.965 -74.35 5.315 -74.23 ;
      RECT 4.965 -71.12 5.315 -71 ;
      RECT 4.965 -67.89 5.315 -67.77 ;
      RECT 4.965 -64.66 5.315 -64.54 ;
      RECT 4.965 -61.43 5.315 -61.31 ;
      RECT 4.965 -58.2 5.315 -58.08 ;
      RECT 4.965 -54.97 5.315 -54.85 ;
      RECT 4.965 -51.74 5.315 -51.62 ;
      RECT 4.965 -48.51 5.315 -48.39 ;
      RECT 4.965 -45.28 5.315 -45.16 ;
      RECT 4.965 -42.05 5.315 -41.93 ;
      RECT 4.965 -38.82 5.315 -38.7 ;
      RECT 4.965 -35.59 5.315 -35.47 ;
      RECT 4.965 -32.36 5.315 -32.24 ;
      RECT 4.965 -29.13 5.315 -29.01 ;
      RECT 4.965 -25.9 5.315 -25.78 ;
      RECT 4.965 -22.67 5.315 -22.55 ;
      RECT 4.965 -19.44 5.315 -19.32 ;
      RECT 4.965 -16.21 5.315 -16.09 ;
      RECT 4.965 -12.98 5.315 -12.86 ;
      RECT 4.965 -9.75 5.315 -9.63 ;
      RECT 4.965 -6.52 5.315 -6.4 ;
      RECT 4.965 -3.29 5.315 -3.17 ;
      RECT 4.965 -0.06 5.315 0.06 ;
      RECT 5.1 -110.735 5.25 -110.445 ;
      RECT 5.135 -108.175 5.235 -107.215 ;
      RECT 5.135 2.175 5.235 3.135 ;
      RECT 5.115 -112.19 5.215 -111.65 ;
      RECT 4.875 -113.555 4.975 -113.085 ;
      RECT 4.875 -108.175 4.975 -107.215 ;
      RECT 4.75 -101.06 4.85 -100.525 ;
      RECT 4.75 -99.735 4.85 -99.2 ;
      RECT 4.75 -97.83 4.85 -97.295 ;
      RECT 4.75 -96.505 4.85 -95.97 ;
      RECT 4.75 -94.6 4.85 -94.065 ;
      RECT 4.75 -93.275 4.85 -92.74 ;
      RECT 4.75 -91.37 4.85 -90.835 ;
      RECT 4.75 -90.045 4.85 -89.51 ;
      RECT 4.75 -88.14 4.85 -87.605 ;
      RECT 4.75 -86.815 4.85 -86.28 ;
      RECT 4.75 -84.91 4.85 -84.375 ;
      RECT 4.75 -83.585 4.85 -83.05 ;
      RECT 4.75 -81.68 4.85 -81.145 ;
      RECT 4.75 -80.355 4.85 -79.82 ;
      RECT 4.75 -78.45 4.85 -77.915 ;
      RECT 4.75 -77.125 4.85 -76.59 ;
      RECT 4.75 -75.22 4.85 -74.685 ;
      RECT 4.75 -73.895 4.85 -73.36 ;
      RECT 4.75 -71.99 4.85 -71.455 ;
      RECT 4.75 -70.665 4.85 -70.13 ;
      RECT 4.75 -68.76 4.85 -68.225 ;
      RECT 4.75 -67.435 4.85 -66.9 ;
      RECT 4.75 -65.53 4.85 -64.995 ;
      RECT 4.75 -64.205 4.85 -63.67 ;
      RECT 4.75 -62.3 4.85 -61.765 ;
      RECT 4.75 -60.975 4.85 -60.44 ;
      RECT 4.75 -59.07 4.85 -58.535 ;
      RECT 4.75 -57.745 4.85 -57.21 ;
      RECT 4.75 -55.84 4.85 -55.305 ;
      RECT 4.75 -54.515 4.85 -53.98 ;
      RECT 4.75 -52.61 4.85 -52.075 ;
      RECT 4.75 -51.285 4.85 -50.75 ;
      RECT 4.75 -49.38 4.85 -48.845 ;
      RECT 4.75 -48.055 4.85 -47.52 ;
      RECT 4.75 -46.15 4.85 -45.615 ;
      RECT 4.75 -44.825 4.85 -44.29 ;
      RECT 4.75 -42.92 4.85 -42.385 ;
      RECT 4.75 -41.595 4.85 -41.06 ;
      RECT 4.75 -39.69 4.85 -39.155 ;
      RECT 4.75 -38.365 4.85 -37.83 ;
      RECT 4.75 -36.46 4.85 -35.925 ;
      RECT 4.75 -35.135 4.85 -34.6 ;
      RECT 4.75 -33.23 4.85 -32.695 ;
      RECT 4.75 -31.905 4.85 -31.37 ;
      RECT 4.75 -30 4.85 -29.465 ;
      RECT 4.75 -28.675 4.85 -28.14 ;
      RECT 4.75 -26.77 4.85 -26.235 ;
      RECT 4.75 -25.445 4.85 -24.91 ;
      RECT 4.75 -23.54 4.85 -23.005 ;
      RECT 4.75 -22.215 4.85 -21.68 ;
      RECT 4.75 -20.31 4.85 -19.775 ;
      RECT 4.75 -18.985 4.85 -18.45 ;
      RECT 4.75 -17.08 4.85 -16.545 ;
      RECT 4.75 -15.755 4.85 -15.22 ;
      RECT 4.75 -13.85 4.85 -13.315 ;
      RECT 4.75 -12.525 4.85 -11.99 ;
      RECT 4.75 -10.62 4.85 -10.085 ;
      RECT 4.75 -9.295 4.85 -8.76 ;
      RECT 4.75 -7.39 4.85 -6.855 ;
      RECT 4.75 -6.065 4.85 -5.53 ;
      RECT 4.75 -4.16 4.85 -3.625 ;
      RECT 4.75 -2.835 4.85 -2.3 ;
      RECT 4.75 -0.93 4.85 -0.395 ;
      RECT 4.75 0.395 4.85 0.93 ;
      RECT 4.625 -104.945 4.725 -103.985 ;
      RECT 4.25 -100.19 4.6 -100.07 ;
      RECT 4.25 -96.96 4.6 -96.84 ;
      RECT 4.25 -93.73 4.6 -93.61 ;
      RECT 4.25 -90.5 4.6 -90.38 ;
      RECT 4.25 -87.27 4.6 -87.15 ;
      RECT 4.25 -84.04 4.6 -83.92 ;
      RECT 4.25 -80.81 4.6 -80.69 ;
      RECT 4.25 -77.58 4.6 -77.46 ;
      RECT 4.25 -74.35 4.6 -74.23 ;
      RECT 4.25 -71.12 4.6 -71 ;
      RECT 4.25 -67.89 4.6 -67.77 ;
      RECT 4.25 -64.66 4.6 -64.54 ;
      RECT 4.25 -61.43 4.6 -61.31 ;
      RECT 4.25 -58.2 4.6 -58.08 ;
      RECT 4.25 -54.97 4.6 -54.85 ;
      RECT 4.25 -51.74 4.6 -51.62 ;
      RECT 4.25 -48.51 4.6 -48.39 ;
      RECT 4.25 -45.28 4.6 -45.16 ;
      RECT 4.25 -42.05 4.6 -41.93 ;
      RECT 4.25 -38.82 4.6 -38.7 ;
      RECT 4.25 -35.59 4.6 -35.47 ;
      RECT 4.25 -32.36 4.6 -32.24 ;
      RECT 4.25 -29.13 4.6 -29.01 ;
      RECT 4.25 -25.9 4.6 -25.78 ;
      RECT 4.25 -22.67 4.6 -22.55 ;
      RECT 4.25 -19.44 4.6 -19.32 ;
      RECT 4.25 -16.21 4.6 -16.09 ;
      RECT 4.25 -12.98 4.6 -12.86 ;
      RECT 4.25 -9.75 4.6 -9.63 ;
      RECT 4.25 -6.52 4.6 -6.4 ;
      RECT 4.25 -3.29 4.6 -3.17 ;
      RECT 4.25 -0.06 4.6 0.06 ;
      RECT 4.365 -104.945 4.465 -103.985 ;
      RECT 4.365 2.175 4.465 3.135 ;
      RECT 4.075 -112.255 4.175 -111.775 ;
      RECT 4.075 -110.765 4.175 -110.295 ;
      RECT 3.765 -100.19 4.115 -100.07 ;
      RECT 3.765 -96.96 4.115 -96.84 ;
      RECT 3.765 -93.73 4.115 -93.61 ;
      RECT 3.765 -90.5 4.115 -90.38 ;
      RECT 3.765 -87.27 4.115 -87.15 ;
      RECT 3.765 -84.04 4.115 -83.92 ;
      RECT 3.765 -80.81 4.115 -80.69 ;
      RECT 3.765 -77.58 4.115 -77.46 ;
      RECT 3.765 -74.35 4.115 -74.23 ;
      RECT 3.765 -71.12 4.115 -71 ;
      RECT 3.765 -67.89 4.115 -67.77 ;
      RECT 3.765 -64.66 4.115 -64.54 ;
      RECT 3.765 -61.43 4.115 -61.31 ;
      RECT 3.765 -58.2 4.115 -58.08 ;
      RECT 3.765 -54.97 4.115 -54.85 ;
      RECT 3.765 -51.74 4.115 -51.62 ;
      RECT 3.765 -48.51 4.115 -48.39 ;
      RECT 3.765 -45.28 4.115 -45.16 ;
      RECT 3.765 -42.05 4.115 -41.93 ;
      RECT 3.765 -38.82 4.115 -38.7 ;
      RECT 3.765 -35.59 4.115 -35.47 ;
      RECT 3.765 -32.36 4.115 -32.24 ;
      RECT 3.765 -29.13 4.115 -29.01 ;
      RECT 3.765 -25.9 4.115 -25.78 ;
      RECT 3.765 -22.67 4.115 -22.55 ;
      RECT 3.765 -19.44 4.115 -19.32 ;
      RECT 3.765 -16.21 4.115 -16.09 ;
      RECT 3.765 -12.98 4.115 -12.86 ;
      RECT 3.765 -9.75 4.115 -9.63 ;
      RECT 3.765 -6.52 4.115 -6.4 ;
      RECT 3.765 -3.29 4.115 -3.17 ;
      RECT 3.765 -0.06 4.115 0.06 ;
      RECT 3.935 -104.945 4.035 -103.985 ;
      RECT 3.935 2.175 4.035 3.135 ;
      RECT 0.035 -108.655 3.815 -108.535 ;
      RECT 3.675 -104.945 3.775 -103.985 ;
      RECT 3.55 -101.06 3.65 -100.525 ;
      RECT 3.55 -99.735 3.65 -99.2 ;
      RECT 3.55 -97.83 3.65 -97.295 ;
      RECT 3.55 -96.505 3.65 -95.97 ;
      RECT 3.55 -94.6 3.65 -94.065 ;
      RECT 3.55 -93.275 3.65 -92.74 ;
      RECT 3.55 -91.37 3.65 -90.835 ;
      RECT 3.55 -90.045 3.65 -89.51 ;
      RECT 3.55 -88.14 3.65 -87.605 ;
      RECT 3.55 -86.815 3.65 -86.28 ;
      RECT 3.55 -84.91 3.65 -84.375 ;
      RECT 3.55 -83.585 3.65 -83.05 ;
      RECT 3.55 -81.68 3.65 -81.145 ;
      RECT 3.55 -80.355 3.65 -79.82 ;
      RECT 3.55 -78.45 3.65 -77.915 ;
      RECT 3.55 -77.125 3.65 -76.59 ;
      RECT 3.55 -75.22 3.65 -74.685 ;
      RECT 3.55 -73.895 3.65 -73.36 ;
      RECT 3.55 -71.99 3.65 -71.455 ;
      RECT 3.55 -70.665 3.65 -70.13 ;
      RECT 3.55 -68.76 3.65 -68.225 ;
      RECT 3.55 -67.435 3.65 -66.9 ;
      RECT 3.55 -65.53 3.65 -64.995 ;
      RECT 3.55 -64.205 3.65 -63.67 ;
      RECT 3.55 -62.3 3.65 -61.765 ;
      RECT 3.55 -60.975 3.65 -60.44 ;
      RECT 3.55 -59.07 3.65 -58.535 ;
      RECT 3.55 -57.745 3.65 -57.21 ;
      RECT 3.55 -55.84 3.65 -55.305 ;
      RECT 3.55 -54.515 3.65 -53.98 ;
      RECT 3.55 -52.61 3.65 -52.075 ;
      RECT 3.55 -51.285 3.65 -50.75 ;
      RECT 3.55 -49.38 3.65 -48.845 ;
      RECT 3.55 -48.055 3.65 -47.52 ;
      RECT 3.55 -46.15 3.65 -45.615 ;
      RECT 3.55 -44.825 3.65 -44.29 ;
      RECT 3.55 -42.92 3.65 -42.385 ;
      RECT 3.55 -41.595 3.65 -41.06 ;
      RECT 3.55 -39.69 3.65 -39.155 ;
      RECT 3.55 -38.365 3.65 -37.83 ;
      RECT 3.55 -36.46 3.65 -35.925 ;
      RECT 3.55 -35.135 3.65 -34.6 ;
      RECT 3.55 -33.23 3.65 -32.695 ;
      RECT 3.55 -31.905 3.65 -31.37 ;
      RECT 3.55 -30 3.65 -29.465 ;
      RECT 3.55 -28.675 3.65 -28.14 ;
      RECT 3.55 -26.77 3.65 -26.235 ;
      RECT 3.55 -25.445 3.65 -24.91 ;
      RECT 3.55 -23.54 3.65 -23.005 ;
      RECT 3.55 -22.215 3.65 -21.68 ;
      RECT 3.55 -20.31 3.65 -19.775 ;
      RECT 3.55 -18.985 3.65 -18.45 ;
      RECT 3.55 -17.08 3.65 -16.545 ;
      RECT 3.55 -15.755 3.65 -15.22 ;
      RECT 3.55 -13.85 3.65 -13.315 ;
      RECT 3.55 -12.525 3.65 -11.99 ;
      RECT 3.55 -10.62 3.65 -10.085 ;
      RECT 3.55 -9.295 3.65 -8.76 ;
      RECT 3.55 -7.39 3.65 -6.855 ;
      RECT 3.55 -6.065 3.65 -5.53 ;
      RECT 3.55 -4.16 3.65 -3.625 ;
      RECT 3.55 -2.835 3.65 -2.3 ;
      RECT 3.55 -0.93 3.65 -0.395 ;
      RECT 3.55 0.395 3.65 0.93 ;
      RECT 3.485 -110.75 3.605 -110.37 ;
      RECT 3.485 -112.245 3.585 -111.775 ;
      RECT 3.425 -104.945 3.525 -103.985 ;
      RECT 3.05 -100.19 3.4 -100.07 ;
      RECT 3.05 -96.96 3.4 -96.84 ;
      RECT 3.05 -93.73 3.4 -93.61 ;
      RECT 3.05 -90.5 3.4 -90.38 ;
      RECT 3.05 -87.27 3.4 -87.15 ;
      RECT 3.05 -84.04 3.4 -83.92 ;
      RECT 3.05 -80.81 3.4 -80.69 ;
      RECT 3.05 -77.58 3.4 -77.46 ;
      RECT 3.05 -74.35 3.4 -74.23 ;
      RECT 3.05 -71.12 3.4 -71 ;
      RECT 3.05 -67.89 3.4 -67.77 ;
      RECT 3.05 -64.66 3.4 -64.54 ;
      RECT 3.05 -61.43 3.4 -61.31 ;
      RECT 3.05 -58.2 3.4 -58.08 ;
      RECT 3.05 -54.97 3.4 -54.85 ;
      RECT 3.05 -51.74 3.4 -51.62 ;
      RECT 3.05 -48.51 3.4 -48.39 ;
      RECT 3.05 -45.28 3.4 -45.16 ;
      RECT 3.05 -42.05 3.4 -41.93 ;
      RECT 3.05 -38.82 3.4 -38.7 ;
      RECT 3.05 -35.59 3.4 -35.47 ;
      RECT 3.05 -32.36 3.4 -32.24 ;
      RECT 3.05 -29.13 3.4 -29.01 ;
      RECT 3.05 -25.9 3.4 -25.78 ;
      RECT 3.05 -22.67 3.4 -22.55 ;
      RECT 3.05 -19.44 3.4 -19.32 ;
      RECT 3.05 -16.21 3.4 -16.09 ;
      RECT 3.05 -12.98 3.4 -12.86 ;
      RECT 3.05 -9.75 3.4 -9.63 ;
      RECT 3.05 -6.52 3.4 -6.4 ;
      RECT 3.05 -3.29 3.4 -3.17 ;
      RECT 3.05 -0.06 3.4 0.06 ;
      RECT 3.165 -104.945 3.265 -103.985 ;
      RECT 3.165 2.175 3.265 3.135 ;
      RECT 2.895 -109.595 3.03 -109.275 ;
      RECT 2.565 -100.19 2.915 -100.07 ;
      RECT 2.565 -96.96 2.915 -96.84 ;
      RECT 2.565 -93.73 2.915 -93.61 ;
      RECT 2.565 -90.5 2.915 -90.38 ;
      RECT 2.565 -87.27 2.915 -87.15 ;
      RECT 2.565 -84.04 2.915 -83.92 ;
      RECT 2.565 -80.81 2.915 -80.69 ;
      RECT 2.565 -77.58 2.915 -77.46 ;
      RECT 2.565 -74.35 2.915 -74.23 ;
      RECT 2.565 -71.12 2.915 -71 ;
      RECT 2.565 -67.89 2.915 -67.77 ;
      RECT 2.565 -64.66 2.915 -64.54 ;
      RECT 2.565 -61.43 2.915 -61.31 ;
      RECT 2.565 -58.2 2.915 -58.08 ;
      RECT 2.565 -54.97 2.915 -54.85 ;
      RECT 2.565 -51.74 2.915 -51.62 ;
      RECT 2.565 -48.51 2.915 -48.39 ;
      RECT 2.565 -45.28 2.915 -45.16 ;
      RECT 2.565 -42.05 2.915 -41.93 ;
      RECT 2.565 -38.82 2.915 -38.7 ;
      RECT 2.565 -35.59 2.915 -35.47 ;
      RECT 2.565 -32.36 2.915 -32.24 ;
      RECT 2.565 -29.13 2.915 -29.01 ;
      RECT 2.565 -25.9 2.915 -25.78 ;
      RECT 2.565 -22.67 2.915 -22.55 ;
      RECT 2.565 -19.44 2.915 -19.32 ;
      RECT 2.565 -16.21 2.915 -16.09 ;
      RECT 2.565 -12.98 2.915 -12.86 ;
      RECT 2.565 -9.75 2.915 -9.63 ;
      RECT 2.565 -6.52 2.915 -6.4 ;
      RECT 2.565 -3.29 2.915 -3.17 ;
      RECT 2.565 -0.06 2.915 0.06 ;
      RECT 2.735 -104.945 2.835 -103.985 ;
      RECT 2.735 2.175 2.835 3.135 ;
      RECT 2.56 -109.595 2.705 -109.275 ;
      RECT 2.475 -104.945 2.575 -103.985 ;
      RECT 2.35 -101.06 2.45 -100.525 ;
      RECT 2.35 -99.735 2.45 -99.2 ;
      RECT 2.35 -97.83 2.45 -97.295 ;
      RECT 2.35 -96.505 2.45 -95.97 ;
      RECT 2.35 -94.6 2.45 -94.065 ;
      RECT 2.35 -93.275 2.45 -92.74 ;
      RECT 2.35 -91.37 2.45 -90.835 ;
      RECT 2.35 -90.045 2.45 -89.51 ;
      RECT 2.35 -88.14 2.45 -87.605 ;
      RECT 2.35 -86.815 2.45 -86.28 ;
      RECT 2.35 -84.91 2.45 -84.375 ;
      RECT 2.35 -83.585 2.45 -83.05 ;
      RECT 2.35 -81.68 2.45 -81.145 ;
      RECT 2.35 -80.355 2.45 -79.82 ;
      RECT 2.35 -78.45 2.45 -77.915 ;
      RECT 2.35 -77.125 2.45 -76.59 ;
      RECT 2.35 -75.22 2.45 -74.685 ;
      RECT 2.35 -73.895 2.45 -73.36 ;
      RECT 2.35 -71.99 2.45 -71.455 ;
      RECT 2.35 -70.665 2.45 -70.13 ;
      RECT 2.35 -68.76 2.45 -68.225 ;
      RECT 2.35 -67.435 2.45 -66.9 ;
      RECT 2.35 -65.53 2.45 -64.995 ;
      RECT 2.35 -64.205 2.45 -63.67 ;
      RECT 2.35 -62.3 2.45 -61.765 ;
      RECT 2.35 -60.975 2.45 -60.44 ;
      RECT 2.35 -59.07 2.45 -58.535 ;
      RECT 2.35 -57.745 2.45 -57.21 ;
      RECT 2.35 -55.84 2.45 -55.305 ;
      RECT 2.35 -54.515 2.45 -53.98 ;
      RECT 2.35 -52.61 2.45 -52.075 ;
      RECT 2.35 -51.285 2.45 -50.75 ;
      RECT 2.35 -49.38 2.45 -48.845 ;
      RECT 2.35 -48.055 2.45 -47.52 ;
      RECT 2.35 -46.15 2.45 -45.615 ;
      RECT 2.35 -44.825 2.45 -44.29 ;
      RECT 2.35 -42.92 2.45 -42.385 ;
      RECT 2.35 -41.595 2.45 -41.06 ;
      RECT 2.35 -39.69 2.45 -39.155 ;
      RECT 2.35 -38.365 2.45 -37.83 ;
      RECT 2.35 -36.46 2.45 -35.925 ;
      RECT 2.35 -35.135 2.45 -34.6 ;
      RECT 2.35 -33.23 2.45 -32.695 ;
      RECT 2.35 -31.905 2.45 -31.37 ;
      RECT 2.35 -30 2.45 -29.465 ;
      RECT 2.35 -28.675 2.45 -28.14 ;
      RECT 2.35 -26.77 2.45 -26.235 ;
      RECT 2.35 -25.445 2.45 -24.91 ;
      RECT 2.35 -23.54 2.45 -23.005 ;
      RECT 2.35 -22.215 2.45 -21.68 ;
      RECT 2.35 -20.31 2.45 -19.775 ;
      RECT 2.35 -18.985 2.45 -18.45 ;
      RECT 2.35 -17.08 2.45 -16.545 ;
      RECT 2.35 -15.755 2.45 -15.22 ;
      RECT 2.35 -13.85 2.45 -13.315 ;
      RECT 2.35 -12.525 2.45 -11.99 ;
      RECT 2.35 -10.62 2.45 -10.085 ;
      RECT 2.35 -9.295 2.45 -8.76 ;
      RECT 2.35 -7.39 2.45 -6.855 ;
      RECT 2.35 -6.065 2.45 -5.53 ;
      RECT 2.35 -4.16 2.45 -3.625 ;
      RECT 2.35 -2.835 2.45 -2.3 ;
      RECT 2.35 -0.93 2.45 -0.395 ;
      RECT 2.35 0.395 2.45 0.93 ;
      RECT 2.225 -108.175 2.325 -107.215 ;
      RECT 1.85 -100.19 2.2 -100.07 ;
      RECT 1.85 -96.96 2.2 -96.84 ;
      RECT 1.85 -93.73 2.2 -93.61 ;
      RECT 1.85 -90.5 2.2 -90.38 ;
      RECT 1.85 -87.27 2.2 -87.15 ;
      RECT 1.85 -84.04 2.2 -83.92 ;
      RECT 1.85 -80.81 2.2 -80.69 ;
      RECT 1.85 -77.58 2.2 -77.46 ;
      RECT 1.85 -74.35 2.2 -74.23 ;
      RECT 1.85 -71.12 2.2 -71 ;
      RECT 1.85 -67.89 2.2 -67.77 ;
      RECT 1.85 -64.66 2.2 -64.54 ;
      RECT 1.85 -61.43 2.2 -61.31 ;
      RECT 1.85 -58.2 2.2 -58.08 ;
      RECT 1.85 -54.97 2.2 -54.85 ;
      RECT 1.85 -51.74 2.2 -51.62 ;
      RECT 1.85 -48.51 2.2 -48.39 ;
      RECT 1.85 -45.28 2.2 -45.16 ;
      RECT 1.85 -42.05 2.2 -41.93 ;
      RECT 1.85 -38.82 2.2 -38.7 ;
      RECT 1.85 -35.59 2.2 -35.47 ;
      RECT 1.85 -32.36 2.2 -32.24 ;
      RECT 1.85 -29.13 2.2 -29.01 ;
      RECT 1.85 -25.9 2.2 -25.78 ;
      RECT 1.85 -22.67 2.2 -22.55 ;
      RECT 1.85 -19.44 2.2 -19.32 ;
      RECT 1.85 -16.21 2.2 -16.09 ;
      RECT 1.85 -12.98 2.2 -12.86 ;
      RECT 1.85 -9.75 2.2 -9.63 ;
      RECT 1.85 -6.52 2.2 -6.4 ;
      RECT 1.85 -3.29 2.2 -3.17 ;
      RECT 1.85 -0.06 2.2 0.06 ;
      RECT 2.055 -112.255 2.155 -111.775 ;
      RECT 2.055 -110.765 2.155 -110.295 ;
      RECT 1.965 -108.175 2.065 -107.215 ;
      RECT 1.965 2.175 2.065 3.135 ;
      RECT 1.365 -100.19 1.715 -100.07 ;
      RECT 1.365 -96.96 1.715 -96.84 ;
      RECT 1.365 -93.73 1.715 -93.61 ;
      RECT 1.365 -90.5 1.715 -90.38 ;
      RECT 1.365 -87.27 1.715 -87.15 ;
      RECT 1.365 -84.04 1.715 -83.92 ;
      RECT 1.365 -80.81 1.715 -80.69 ;
      RECT 1.365 -77.58 1.715 -77.46 ;
      RECT 1.365 -74.35 1.715 -74.23 ;
      RECT 1.365 -71.12 1.715 -71 ;
      RECT 1.365 -67.89 1.715 -67.77 ;
      RECT 1.365 -64.66 1.715 -64.54 ;
      RECT 1.365 -61.43 1.715 -61.31 ;
      RECT 1.365 -58.2 1.715 -58.08 ;
      RECT 1.365 -54.97 1.715 -54.85 ;
      RECT 1.365 -51.74 1.715 -51.62 ;
      RECT 1.365 -48.51 1.715 -48.39 ;
      RECT 1.365 -45.28 1.715 -45.16 ;
      RECT 1.365 -42.05 1.715 -41.93 ;
      RECT 1.365 -38.82 1.715 -38.7 ;
      RECT 1.365 -35.59 1.715 -35.47 ;
      RECT 1.365 -32.36 1.715 -32.24 ;
      RECT 1.365 -29.13 1.715 -29.01 ;
      RECT 1.365 -25.9 1.715 -25.78 ;
      RECT 1.365 -22.67 1.715 -22.55 ;
      RECT 1.365 -19.44 1.715 -19.32 ;
      RECT 1.365 -16.21 1.715 -16.09 ;
      RECT 1.365 -12.98 1.715 -12.86 ;
      RECT 1.365 -9.75 1.715 -9.63 ;
      RECT 1.365 -6.52 1.715 -6.4 ;
      RECT 1.365 -3.29 1.715 -3.17 ;
      RECT 1.365 -0.06 1.715 0.06 ;
      RECT 1.535 -108.175 1.635 -107.215 ;
      RECT 1.535 2.175 1.635 3.135 ;
      RECT 1.43 -110.765 1.6 -110.385 ;
      RECT 1.465 -112.245 1.565 -111.775 ;
      RECT 1.275 -108.175 1.375 -107.215 ;
      RECT 1.15 -101.06 1.25 -100.525 ;
      RECT 1.15 -99.735 1.25 -99.2 ;
      RECT 1.15 -97.83 1.25 -97.295 ;
      RECT 1.15 -96.505 1.25 -95.97 ;
      RECT 1.15 -94.6 1.25 -94.065 ;
      RECT 1.15 -93.275 1.25 -92.74 ;
      RECT 1.15 -91.37 1.25 -90.835 ;
      RECT 1.15 -90.045 1.25 -89.51 ;
      RECT 1.15 -88.14 1.25 -87.605 ;
      RECT 1.15 -86.815 1.25 -86.28 ;
      RECT 1.15 -84.91 1.25 -84.375 ;
      RECT 1.15 -83.585 1.25 -83.05 ;
      RECT 1.15 -81.68 1.25 -81.145 ;
      RECT 1.15 -80.355 1.25 -79.82 ;
      RECT 1.15 -78.45 1.25 -77.915 ;
      RECT 1.15 -77.125 1.25 -76.59 ;
      RECT 1.15 -75.22 1.25 -74.685 ;
      RECT 1.15 -73.895 1.25 -73.36 ;
      RECT 1.15 -71.99 1.25 -71.455 ;
      RECT 1.15 -70.665 1.25 -70.13 ;
      RECT 1.15 -68.76 1.25 -68.225 ;
      RECT 1.15 -67.435 1.25 -66.9 ;
      RECT 1.15 -65.53 1.25 -64.995 ;
      RECT 1.15 -64.205 1.25 -63.67 ;
      RECT 1.15 -62.3 1.25 -61.765 ;
      RECT 1.15 -60.975 1.25 -60.44 ;
      RECT 1.15 -59.07 1.25 -58.535 ;
      RECT 1.15 -57.745 1.25 -57.21 ;
      RECT 1.15 -55.84 1.25 -55.305 ;
      RECT 1.15 -54.515 1.25 -53.98 ;
      RECT 1.15 -52.61 1.25 -52.075 ;
      RECT 1.15 -51.285 1.25 -50.75 ;
      RECT 1.15 -49.38 1.25 -48.845 ;
      RECT 1.15 -48.055 1.25 -47.52 ;
      RECT 1.15 -46.15 1.25 -45.615 ;
      RECT 1.15 -44.825 1.25 -44.29 ;
      RECT 1.15 -42.92 1.25 -42.385 ;
      RECT 1.15 -41.595 1.25 -41.06 ;
      RECT 1.15 -39.69 1.25 -39.155 ;
      RECT 1.15 -38.365 1.25 -37.83 ;
      RECT 1.15 -36.46 1.25 -35.925 ;
      RECT 1.15 -35.135 1.25 -34.6 ;
      RECT 1.15 -33.23 1.25 -32.695 ;
      RECT 1.15 -31.905 1.25 -31.37 ;
      RECT 1.15 -30 1.25 -29.465 ;
      RECT 1.15 -28.675 1.25 -28.14 ;
      RECT 1.15 -26.77 1.25 -26.235 ;
      RECT 1.15 -25.445 1.25 -24.91 ;
      RECT 1.15 -23.54 1.25 -23.005 ;
      RECT 1.15 -22.215 1.25 -21.68 ;
      RECT 1.15 -20.31 1.25 -19.775 ;
      RECT 1.15 -18.985 1.25 -18.45 ;
      RECT 1.15 -17.08 1.25 -16.545 ;
      RECT 1.15 -15.755 1.25 -15.22 ;
      RECT 1.15 -13.85 1.25 -13.315 ;
      RECT 1.15 -12.525 1.25 -11.99 ;
      RECT 1.15 -10.62 1.25 -10.085 ;
      RECT 1.15 -9.295 1.25 -8.76 ;
      RECT 1.15 -7.39 1.25 -6.855 ;
      RECT 1.15 -6.065 1.25 -5.53 ;
      RECT 1.15 -4.16 1.25 -3.625 ;
      RECT 1.15 -2.835 1.25 -2.3 ;
      RECT 1.15 -0.93 1.25 -0.395 ;
      RECT 1.15 0.395 1.25 0.93 ;
      RECT 1.025 -108.175 1.125 -107.215 ;
      RECT 0.65 -100.19 1 -100.07 ;
      RECT 0.65 -96.96 1 -96.84 ;
      RECT 0.65 -93.73 1 -93.61 ;
      RECT 0.65 -90.5 1 -90.38 ;
      RECT 0.65 -87.27 1 -87.15 ;
      RECT 0.65 -84.04 1 -83.92 ;
      RECT 0.65 -80.81 1 -80.69 ;
      RECT 0.65 -77.58 1 -77.46 ;
      RECT 0.65 -74.35 1 -74.23 ;
      RECT 0.65 -71.12 1 -71 ;
      RECT 0.65 -67.89 1 -67.77 ;
      RECT 0.65 -64.66 1 -64.54 ;
      RECT 0.65 -61.43 1 -61.31 ;
      RECT 0.65 -58.2 1 -58.08 ;
      RECT 0.65 -54.97 1 -54.85 ;
      RECT 0.65 -51.74 1 -51.62 ;
      RECT 0.65 -48.51 1 -48.39 ;
      RECT 0.65 -45.28 1 -45.16 ;
      RECT 0.65 -42.05 1 -41.93 ;
      RECT 0.65 -38.82 1 -38.7 ;
      RECT 0.65 -35.59 1 -35.47 ;
      RECT 0.65 -32.36 1 -32.24 ;
      RECT 0.65 -29.13 1 -29.01 ;
      RECT 0.65 -25.9 1 -25.78 ;
      RECT 0.65 -22.67 1 -22.55 ;
      RECT 0.65 -19.44 1 -19.32 ;
      RECT 0.65 -16.21 1 -16.09 ;
      RECT 0.65 -12.98 1 -12.86 ;
      RECT 0.65 -9.75 1 -9.63 ;
      RECT 0.65 -6.52 1 -6.4 ;
      RECT 0.65 -3.29 1 -3.17 ;
      RECT 0.65 -0.06 1 0.06 ;
      RECT 0.765 -108.175 0.865 -107.215 ;
      RECT 0.765 2.175 0.865 3.135 ;
      RECT 0.665 -113.555 0.765 -113.085 ;
      RECT 0.165 -100.19 0.515 -100.07 ;
      RECT 0.165 -96.96 0.515 -96.84 ;
      RECT 0.165 -93.73 0.515 -93.61 ;
      RECT 0.165 -90.5 0.515 -90.38 ;
      RECT 0.165 -87.27 0.515 -87.15 ;
      RECT 0.165 -84.04 0.515 -83.92 ;
      RECT 0.165 -80.81 0.515 -80.69 ;
      RECT 0.165 -77.58 0.515 -77.46 ;
      RECT 0.165 -74.35 0.515 -74.23 ;
      RECT 0.165 -71.12 0.515 -71 ;
      RECT 0.165 -67.89 0.515 -67.77 ;
      RECT 0.165 -64.66 0.515 -64.54 ;
      RECT 0.165 -61.43 0.515 -61.31 ;
      RECT 0.165 -58.2 0.515 -58.08 ;
      RECT 0.165 -54.97 0.515 -54.85 ;
      RECT 0.165 -51.74 0.515 -51.62 ;
      RECT 0.165 -48.51 0.515 -48.39 ;
      RECT 0.165 -45.28 0.515 -45.16 ;
      RECT 0.165 -42.05 0.515 -41.93 ;
      RECT 0.165 -38.82 0.515 -38.7 ;
      RECT 0.165 -35.59 0.515 -35.47 ;
      RECT 0.165 -32.36 0.515 -32.24 ;
      RECT 0.165 -29.13 0.515 -29.01 ;
      RECT 0.165 -25.9 0.515 -25.78 ;
      RECT 0.165 -22.67 0.515 -22.55 ;
      RECT 0.165 -19.44 0.515 -19.32 ;
      RECT 0.165 -16.21 0.515 -16.09 ;
      RECT 0.165 -12.98 0.515 -12.86 ;
      RECT 0.165 -9.75 0.515 -9.63 ;
      RECT 0.165 -6.52 0.515 -6.4 ;
      RECT 0.165 -3.29 0.515 -3.17 ;
      RECT 0.165 -0.06 0.515 0.06 ;
      RECT 0.3 -110.735 0.45 -110.445 ;
      RECT 0.335 -108.175 0.435 -107.215 ;
      RECT 0.335 2.175 0.435 3.135 ;
      RECT 0.315 -112.19 0.415 -111.65 ;
      RECT 0.075 -113.555 0.175 -113.085 ;
      RECT 0.075 -108.175 0.175 -107.215 ;
      RECT -0.05 -101.06 0.05 -100.525 ;
      RECT -0.05 -99.735 0.05 -99.2 ;
      RECT -0.05 -97.83 0.05 -97.295 ;
      RECT -0.05 -96.505 0.05 -95.97 ;
      RECT -0.05 -94.6 0.05 -94.065 ;
      RECT -0.05 -93.275 0.05 -92.74 ;
      RECT -0.05 -91.37 0.05 -90.835 ;
      RECT -0.05 -90.045 0.05 -89.51 ;
      RECT -0.05 -88.14 0.05 -87.605 ;
      RECT -0.05 -86.815 0.05 -86.28 ;
      RECT -0.05 -84.91 0.05 -84.375 ;
      RECT -0.05 -83.585 0.05 -83.05 ;
      RECT -0.05 -81.68 0.05 -81.145 ;
      RECT -0.05 -80.355 0.05 -79.82 ;
      RECT -0.05 -78.45 0.05 -77.915 ;
      RECT -0.05 -77.125 0.05 -76.59 ;
      RECT -0.05 -75.22 0.05 -74.685 ;
      RECT -0.05 -73.895 0.05 -73.36 ;
      RECT -0.05 -71.99 0.05 -71.455 ;
      RECT -0.05 -70.665 0.05 -70.13 ;
      RECT -0.05 -68.76 0.05 -68.225 ;
      RECT -0.05 -67.435 0.05 -66.9 ;
      RECT -0.05 -65.53 0.05 -64.995 ;
      RECT -0.05 -64.205 0.05 -63.67 ;
      RECT -0.05 -62.3 0.05 -61.765 ;
      RECT -0.05 -60.975 0.05 -60.44 ;
      RECT -0.05 -59.07 0.05 -58.535 ;
      RECT -0.05 -57.745 0.05 -57.21 ;
      RECT -0.05 -55.84 0.05 -55.305 ;
      RECT -0.05 -54.515 0.05 -53.98 ;
      RECT -0.05 -52.61 0.05 -52.075 ;
      RECT -0.05 -51.285 0.05 -50.75 ;
      RECT -0.05 -49.38 0.05 -48.845 ;
      RECT -0.05 -48.055 0.05 -47.52 ;
      RECT -0.05 -46.15 0.05 -45.615 ;
      RECT -0.05 -44.825 0.05 -44.29 ;
      RECT -0.05 -42.92 0.05 -42.385 ;
      RECT -0.05 -41.595 0.05 -41.06 ;
      RECT -0.05 -39.69 0.05 -39.155 ;
      RECT -0.05 -38.365 0.05 -37.83 ;
      RECT -0.05 -36.46 0.05 -35.925 ;
      RECT -0.05 -35.135 0.05 -34.6 ;
      RECT -0.05 -33.23 0.05 -32.695 ;
      RECT -0.05 -31.905 0.05 -31.37 ;
      RECT -0.05 -30 0.05 -29.465 ;
      RECT -0.05 -28.675 0.05 -28.14 ;
      RECT -0.05 -26.77 0.05 -26.235 ;
      RECT -0.05 -25.445 0.05 -24.91 ;
      RECT -0.05 -23.54 0.05 -23.005 ;
      RECT -0.05 -22.215 0.05 -21.68 ;
      RECT -0.05 -20.31 0.05 -19.775 ;
      RECT -0.05 -18.985 0.05 -18.45 ;
      RECT -0.05 -17.08 0.05 -16.545 ;
      RECT -0.05 -15.755 0.05 -15.22 ;
      RECT -0.05 -13.85 0.05 -13.315 ;
      RECT -0.05 -12.525 0.05 -11.99 ;
      RECT -0.05 -10.62 0.05 -10.085 ;
      RECT -0.05 -9.295 0.05 -8.76 ;
      RECT -0.05 -7.39 0.05 -6.855 ;
      RECT -0.05 -6.065 0.05 -5.53 ;
      RECT -0.05 -4.16 0.05 -3.625 ;
      RECT -0.05 -2.835 0.05 -2.3 ;
      RECT -0.05 -0.93 0.05 -0.395 ;
      RECT -0.05 0.395 0.05 0.93 ;
      RECT -0.945 -107.655 -0.845 -107.235 ;
      RECT -0.945 -102.895 -0.845 -102.295 ;
      RECT -0.945 -101.195 -0.845 -100.595 ;
      RECT -0.945 -96.255 -0.845 -95.835 ;
      RECT -0.945 -94.735 -0.845 -94.315 ;
      RECT -0.945 -89.975 -0.845 -89.375 ;
      RECT -0.945 -88.275 -0.845 -87.675 ;
      RECT -0.945 -83.335 -0.845 -82.915 ;
      RECT -0.945 -81.815 -0.845 -81.395 ;
      RECT -0.945 -77.055 -0.845 -76.455 ;
      RECT -0.945 -75.355 -0.845 -74.755 ;
      RECT -0.945 -70.415 -0.845 -69.995 ;
      RECT -0.945 -68.895 -0.845 -68.475 ;
      RECT -0.945 -64.135 -0.845 -63.535 ;
      RECT -0.945 -62.435 -0.845 -61.835 ;
      RECT -0.945 -57.495 -0.845 -57.075 ;
      RECT -0.945 -55.975 -0.845 -55.555 ;
      RECT -0.945 -51.215 -0.845 -50.615 ;
      RECT -0.945 -49.515 -0.845 -48.915 ;
      RECT -0.945 -44.575 -0.845 -44.155 ;
      RECT -0.945 -43.055 -0.845 -42.635 ;
      RECT -0.945 -38.295 -0.845 -37.695 ;
      RECT -0.945 -36.595 -0.845 -35.995 ;
      RECT -0.945 -31.655 -0.845 -31.235 ;
      RECT -0.945 -30.135 -0.845 -29.715 ;
      RECT -0.945 -25.375 -0.845 -24.775 ;
      RECT -0.945 -23.675 -0.845 -23.075 ;
      RECT -0.945 -18.735 -0.845 -18.315 ;
      RECT -0.945 -17.215 -0.845 -16.795 ;
      RECT -0.945 -12.455 -0.845 -11.855 ;
      RECT -0.945 -10.755 -0.845 -10.155 ;
      RECT -0.945 -5.815 -0.845 -5.395 ;
      RECT -0.945 -4.295 -0.845 -3.875 ;
      RECT -0.945 0.465 -0.845 1.065 ;
      RECT -2.025 -103.41 -0.94 -103.31 ;
      RECT -2.025 -100.18 -0.94 -100.08 ;
      RECT -2.025 -90.49 -0.94 -90.39 ;
      RECT -2.025 -87.26 -0.94 -87.16 ;
      RECT -2.025 -77.57 -0.94 -77.47 ;
      RECT -2.025 -74.34 -0.94 -74.24 ;
      RECT -2.025 -64.65 -0.94 -64.55 ;
      RECT -2.025 -61.42 -0.94 -61.32 ;
      RECT -2.025 -51.73 -0.94 -51.63 ;
      RECT -2.025 -48.5 -0.94 -48.4 ;
      RECT -2.025 -38.81 -0.94 -38.71 ;
      RECT -2.025 -35.58 -0.94 -35.48 ;
      RECT -2.025 -25.89 -0.94 -25.79 ;
      RECT -2.025 -22.66 -0.94 -22.56 ;
      RECT -2.025 -12.97 -0.94 -12.87 ;
      RECT -2.025 -9.74 -0.94 -9.64 ;
      RECT -2.025 -0.05 -0.94 0.05 ;
      RECT -1.465 -107.655 -1.365 -107.055 ;
      RECT -1.465 -102.895 -1.365 -102.295 ;
      RECT -1.465 -101.195 -1.365 -100.595 ;
      RECT -1.465 -96.435 -1.365 -95.835 ;
      RECT -1.465 -94.735 -1.365 -94.135 ;
      RECT -1.465 -89.975 -1.365 -89.375 ;
      RECT -1.465 -88.275 -1.365 -87.675 ;
      RECT -1.465 -83.515 -1.365 -82.915 ;
      RECT -1.465 -81.815 -1.365 -81.215 ;
      RECT -1.465 -77.055 -1.365 -76.455 ;
      RECT -1.465 -75.355 -1.365 -74.755 ;
      RECT -1.465 -70.595 -1.365 -69.995 ;
      RECT -1.465 -68.895 -1.365 -68.295 ;
      RECT -1.465 -64.135 -1.365 -63.535 ;
      RECT -1.465 -62.435 -1.365 -61.835 ;
      RECT -1.465 -57.675 -1.365 -57.075 ;
      RECT -1.465 -55.975 -1.365 -55.375 ;
      RECT -1.465 -51.215 -1.365 -50.615 ;
      RECT -1.465 -49.515 -1.365 -48.915 ;
      RECT -1.465 -44.755 -1.365 -44.155 ;
      RECT -1.465 -43.055 -1.365 -42.455 ;
      RECT -1.465 -38.295 -1.365 -37.695 ;
      RECT -1.465 -36.595 -1.365 -35.995 ;
      RECT -1.465 -31.835 -1.365 -31.235 ;
      RECT -1.465 -30.135 -1.365 -29.535 ;
      RECT -1.465 -25.375 -1.365 -24.775 ;
      RECT -1.465 -23.675 -1.365 -23.075 ;
      RECT -1.465 -18.915 -1.365 -18.315 ;
      RECT -1.465 -17.215 -1.365 -16.615 ;
      RECT -1.465 -12.455 -1.365 -11.855 ;
      RECT -1.465 -10.755 -1.365 -10.155 ;
      RECT -1.465 -5.995 -1.365 -5.395 ;
      RECT -1.465 -4.295 -1.365 -3.695 ;
      RECT -1.465 0.465 -1.365 1.065 ;
      RECT -8.785 -104.655 -1.46 -104.555 ;
      RECT -19.185 -97.615 -1.46 -97.515 ;
      RECT -19.185 -93.055 -1.46 -92.955 ;
      RECT -19.185 -84.695 -1.46 -84.595 ;
      RECT -19.185 -80.135 -1.46 -80.035 ;
      RECT -19.185 -71.775 -1.46 -71.675 ;
      RECT -19.185 -67.215 -1.46 -67.115 ;
      RECT -19.185 -58.855 -1.46 -58.755 ;
      RECT -19.185 -54.295 -1.46 -54.195 ;
      RECT -19.185 -45.935 -1.46 -45.835 ;
      RECT -19.185 -41.375 -1.46 -41.275 ;
      RECT -19.185 -33.015 -1.46 -32.915 ;
      RECT -19.185 -28.455 -1.46 -28.355 ;
      RECT -19.185 -20.095 -1.46 -19.995 ;
      RECT -19.185 -15.535 -1.46 -15.435 ;
      RECT -19.185 -7.175 -1.46 -7.075 ;
      RECT -19.185 -2.615 -1.46 -2.515 ;
      RECT -1.725 -107.655 -1.625 -107.055 ;
      RECT -1.725 -96.435 -1.625 -95.835 ;
      RECT -1.725 -94.735 -1.625 -94.135 ;
      RECT -1.725 -83.515 -1.625 -82.915 ;
      RECT -1.725 -81.815 -1.625 -81.215 ;
      RECT -1.725 -70.595 -1.625 -69.995 ;
      RECT -1.725 -68.895 -1.625 -68.295 ;
      RECT -1.725 -57.675 -1.625 -57.075 ;
      RECT -1.725 -55.975 -1.625 -55.375 ;
      RECT -1.725 -44.755 -1.625 -44.155 ;
      RECT -1.725 -43.055 -1.625 -42.455 ;
      RECT -1.725 -31.835 -1.625 -31.235 ;
      RECT -1.725 -30.135 -1.625 -29.535 ;
      RECT -1.725 -18.915 -1.625 -18.315 ;
      RECT -1.725 -17.215 -1.625 -16.615 ;
      RECT -1.725 -5.995 -1.625 -5.395 ;
      RECT -1.725 -4.295 -1.625 -3.695 ;
      RECT -6.085 -103.995 -1.72 -103.895 ;
      RECT -6.085 -99.375 -1.72 -99.275 ;
      RECT -6.085 -91.295 -1.72 -91.195 ;
      RECT -6.085 -86.455 -1.72 -86.355 ;
      RECT -6.085 -78.375 -1.72 -78.275 ;
      RECT -6.085 -73.535 -1.72 -73.435 ;
      RECT -6.085 -65.455 -1.72 -65.355 ;
      RECT -6.085 -60.615 -1.72 -60.515 ;
      RECT -6.085 -52.535 -1.72 -52.435 ;
      RECT -6.085 -47.695 -1.72 -47.595 ;
      RECT -6.085 -39.615 -1.72 -39.515 ;
      RECT -6.085 -34.775 -1.72 -34.675 ;
      RECT -6.085 -26.695 -1.72 -26.595 ;
      RECT -6.085 -21.855 -1.72 -21.755 ;
      RECT -6.085 -13.775 -1.72 -13.675 ;
      RECT -6.085 -8.935 -1.72 -8.835 ;
      RECT -6.085 -0.855 -1.72 -0.755 ;
      RECT -1.985 -102.895 -1.885 -102.295 ;
      RECT -1.985 -101.195 -1.885 -100.595 ;
      RECT -1.985 -89.975 -1.885 -89.375 ;
      RECT -1.985 -88.275 -1.885 -87.675 ;
      RECT -1.985 -77.055 -1.885 -76.455 ;
      RECT -1.985 -75.355 -1.885 -74.755 ;
      RECT -1.985 -64.135 -1.885 -63.535 ;
      RECT -1.985 -62.435 -1.885 -61.835 ;
      RECT -1.985 -51.215 -1.885 -50.615 ;
      RECT -1.985 -49.515 -1.885 -48.915 ;
      RECT -1.985 -38.295 -1.885 -37.695 ;
      RECT -1.985 -36.595 -1.885 -35.995 ;
      RECT -1.985 -25.375 -1.885 -24.775 ;
      RECT -1.985 -23.675 -1.885 -23.075 ;
      RECT -1.985 -12.455 -1.885 -11.855 ;
      RECT -1.985 -10.755 -1.885 -10.155 ;
      RECT -1.985 0.465 -1.885 1.065 ;
      RECT -2.245 -107.655 -2.145 -107.235 ;
      RECT -2.245 -102.895 -2.145 -102.295 ;
      RECT -2.245 -101.195 -2.145 -100.595 ;
      RECT -2.245 -96.255 -2.145 -95.835 ;
      RECT -2.245 -94.735 -2.145 -94.315 ;
      RECT -2.245 -89.975 -2.145 -89.375 ;
      RECT -2.245 -88.275 -2.145 -87.675 ;
      RECT -2.245 -83.335 -2.145 -82.915 ;
      RECT -2.245 -81.815 -2.145 -81.395 ;
      RECT -2.245 -77.055 -2.145 -76.455 ;
      RECT -2.245 -75.355 -2.145 -74.755 ;
      RECT -2.245 -70.415 -2.145 -69.995 ;
      RECT -2.245 -68.895 -2.145 -68.475 ;
      RECT -2.245 -64.135 -2.145 -63.535 ;
      RECT -2.245 -62.435 -2.145 -61.835 ;
      RECT -2.245 -57.495 -2.145 -57.075 ;
      RECT -2.245 -55.975 -2.145 -55.555 ;
      RECT -2.245 -51.215 -2.145 -50.615 ;
      RECT -2.245 -49.515 -2.145 -48.915 ;
      RECT -2.245 -44.575 -2.145 -44.155 ;
      RECT -2.245 -43.055 -2.145 -42.635 ;
      RECT -2.245 -38.295 -2.145 -37.695 ;
      RECT -2.245 -36.595 -2.145 -35.995 ;
      RECT -2.245 -31.655 -2.145 -31.235 ;
      RECT -2.245 -30.135 -2.145 -29.715 ;
      RECT -2.245 -25.375 -2.145 -24.775 ;
      RECT -2.245 -23.675 -2.145 -23.075 ;
      RECT -2.245 -18.735 -2.145 -18.315 ;
      RECT -2.245 -17.215 -2.145 -16.795 ;
      RECT -2.245 -12.455 -2.145 -11.855 ;
      RECT -2.245 -10.755 -2.145 -10.155 ;
      RECT -2.245 -5.815 -2.145 -5.395 ;
      RECT -2.245 -4.295 -2.145 -3.875 ;
      RECT -2.245 0.465 -2.145 1.065 ;
      RECT -3.325 -103.41 -2.24 -103.31 ;
      RECT -3.325 -100.18 -2.24 -100.08 ;
      RECT -3.325 -90.49 -2.24 -90.39 ;
      RECT -3.325 -87.26 -2.24 -87.16 ;
      RECT -3.325 -77.57 -2.24 -77.47 ;
      RECT -3.325 -74.34 -2.24 -74.24 ;
      RECT -3.325 -64.65 -2.24 -64.55 ;
      RECT -3.325 -61.42 -2.24 -61.32 ;
      RECT -3.325 -51.73 -2.24 -51.63 ;
      RECT -3.325 -48.5 -2.24 -48.4 ;
      RECT -3.325 -38.81 -2.24 -38.71 ;
      RECT -3.325 -35.58 -2.24 -35.48 ;
      RECT -3.325 -25.89 -2.24 -25.79 ;
      RECT -3.325 -22.66 -2.24 -22.56 ;
      RECT -3.325 -12.97 -2.24 -12.87 ;
      RECT -3.325 -9.74 -2.24 -9.64 ;
      RECT -3.325 -0.05 -2.24 0.05 ;
      RECT -2.765 -107.655 -2.665 -107.055 ;
      RECT -2.765 -102.895 -2.665 -102.295 ;
      RECT -2.765 -101.195 -2.665 -100.595 ;
      RECT -2.765 -96.435 -2.665 -95.835 ;
      RECT -2.765 -94.735 -2.665 -94.135 ;
      RECT -2.765 -89.975 -2.665 -89.375 ;
      RECT -2.765 -88.275 -2.665 -87.675 ;
      RECT -2.765 -83.515 -2.665 -82.915 ;
      RECT -2.765 -81.815 -2.665 -81.215 ;
      RECT -2.765 -77.055 -2.665 -76.455 ;
      RECT -2.765 -75.355 -2.665 -74.755 ;
      RECT -2.765 -70.595 -2.665 -69.995 ;
      RECT -2.765 -68.895 -2.665 -68.295 ;
      RECT -2.765 -64.135 -2.665 -63.535 ;
      RECT -2.765 -62.435 -2.665 -61.835 ;
      RECT -2.765 -57.675 -2.665 -57.075 ;
      RECT -2.765 -55.975 -2.665 -55.375 ;
      RECT -2.765 -51.215 -2.665 -50.615 ;
      RECT -2.765 -49.515 -2.665 -48.915 ;
      RECT -2.765 -44.755 -2.665 -44.155 ;
      RECT -2.765 -43.055 -2.665 -42.455 ;
      RECT -2.765 -38.295 -2.665 -37.695 ;
      RECT -2.765 -36.595 -2.665 -35.995 ;
      RECT -2.765 -31.835 -2.665 -31.235 ;
      RECT -2.765 -30.135 -2.665 -29.535 ;
      RECT -2.765 -25.375 -2.665 -24.775 ;
      RECT -2.765 -23.675 -2.665 -23.075 ;
      RECT -2.765 -18.915 -2.665 -18.315 ;
      RECT -2.765 -17.215 -2.665 -16.615 ;
      RECT -2.765 -12.455 -2.665 -11.855 ;
      RECT -2.765 -10.755 -2.665 -10.155 ;
      RECT -2.765 -5.995 -2.665 -5.395 ;
      RECT -2.765 -4.295 -2.665 -3.695 ;
      RECT -2.765 0.465 -2.665 1.065 ;
      RECT -10.085 -104.435 -2.76 -104.335 ;
      RECT -25.685 -97.835 -2.76 -97.735 ;
      RECT -25.685 -92.835 -2.76 -92.735 ;
      RECT -25.685 -84.915 -2.76 -84.815 ;
      RECT -25.685 -79.915 -2.76 -79.815 ;
      RECT -25.685 -71.995 -2.76 -71.895 ;
      RECT -25.685 -66.995 -2.76 -66.895 ;
      RECT -25.685 -59.075 -2.76 -58.975 ;
      RECT -25.685 -54.075 -2.76 -53.975 ;
      RECT -25.685 -46.155 -2.76 -46.055 ;
      RECT -25.685 -41.155 -2.76 -41.055 ;
      RECT -25.685 -33.235 -2.76 -33.135 ;
      RECT -25.685 -28.235 -2.76 -28.135 ;
      RECT -25.685 -20.315 -2.76 -20.215 ;
      RECT -25.685 -15.315 -2.76 -15.215 ;
      RECT -25.685 -7.395 -2.76 -7.295 ;
      RECT -25.685 -2.395 -2.76 -2.295 ;
      RECT -3.025 -107.655 -2.925 -107.055 ;
      RECT -3.025 -96.435 -2.925 -95.835 ;
      RECT -3.025 -94.735 -2.925 -94.135 ;
      RECT -3.025 -83.515 -2.925 -82.915 ;
      RECT -3.025 -81.815 -2.925 -81.215 ;
      RECT -3.025 -70.595 -2.925 -69.995 ;
      RECT -3.025 -68.895 -2.925 -68.295 ;
      RECT -3.025 -57.675 -2.925 -57.075 ;
      RECT -3.025 -55.975 -2.925 -55.375 ;
      RECT -3.025 -44.755 -2.925 -44.155 ;
      RECT -3.025 -43.055 -2.925 -42.455 ;
      RECT -3.025 -31.835 -2.925 -31.235 ;
      RECT -3.025 -30.135 -2.925 -29.535 ;
      RECT -3.025 -18.915 -2.925 -18.315 ;
      RECT -3.025 -17.215 -2.925 -16.615 ;
      RECT -3.025 -5.995 -2.925 -5.395 ;
      RECT -3.025 -4.295 -2.925 -3.695 ;
      RECT -3.285 -102.895 -3.185 -102.295 ;
      RECT -3.285 -101.195 -3.185 -100.595 ;
      RECT -3.285 -89.975 -3.185 -89.375 ;
      RECT -3.285 -88.275 -3.185 -87.675 ;
      RECT -3.285 -77.055 -3.185 -76.455 ;
      RECT -3.285 -75.355 -3.185 -74.755 ;
      RECT -3.285 -64.135 -3.185 -63.535 ;
      RECT -3.285 -62.435 -3.185 -61.835 ;
      RECT -3.285 -51.215 -3.185 -50.615 ;
      RECT -3.285 -49.515 -3.185 -48.915 ;
      RECT -3.285 -38.295 -3.185 -37.695 ;
      RECT -3.285 -36.595 -3.185 -35.995 ;
      RECT -3.285 -25.375 -3.185 -24.775 ;
      RECT -3.285 -23.675 -3.185 -23.075 ;
      RECT -3.285 -12.455 -3.185 -11.855 ;
      RECT -3.285 -10.755 -3.185 -10.155 ;
      RECT -3.285 0.465 -3.185 1.065 ;
      RECT -3.545 -107.655 -3.445 -107.235 ;
      RECT -3.545 -102.895 -3.445 -102.295 ;
      RECT -3.545 -101.195 -3.445 -100.595 ;
      RECT -3.545 -96.255 -3.445 -95.835 ;
      RECT -3.545 -94.735 -3.445 -94.315 ;
      RECT -3.545 -89.975 -3.445 -89.375 ;
      RECT -3.545 -88.275 -3.445 -87.675 ;
      RECT -3.545 -83.335 -3.445 -82.915 ;
      RECT -3.545 -81.815 -3.445 -81.395 ;
      RECT -3.545 -77.055 -3.445 -76.455 ;
      RECT -3.545 -75.355 -3.445 -74.755 ;
      RECT -3.545 -70.415 -3.445 -69.995 ;
      RECT -3.545 -68.895 -3.445 -68.475 ;
      RECT -3.545 -64.135 -3.445 -63.535 ;
      RECT -3.545 -62.435 -3.445 -61.835 ;
      RECT -3.545 -57.495 -3.445 -57.075 ;
      RECT -3.545 -55.975 -3.445 -55.555 ;
      RECT -3.545 -51.215 -3.445 -50.615 ;
      RECT -3.545 -49.515 -3.445 -48.915 ;
      RECT -3.545 -44.575 -3.445 -44.155 ;
      RECT -3.545 -43.055 -3.445 -42.635 ;
      RECT -3.545 -38.295 -3.445 -37.695 ;
      RECT -3.545 -36.595 -3.445 -35.995 ;
      RECT -3.545 -31.655 -3.445 -31.235 ;
      RECT -3.545 -30.135 -3.445 -29.715 ;
      RECT -3.545 -25.375 -3.445 -24.775 ;
      RECT -3.545 -23.675 -3.445 -23.075 ;
      RECT -3.545 -18.735 -3.445 -18.315 ;
      RECT -3.545 -17.215 -3.445 -16.795 ;
      RECT -3.545 -12.455 -3.445 -11.855 ;
      RECT -3.545 -10.755 -3.445 -10.155 ;
      RECT -3.545 -5.815 -3.445 -5.395 ;
      RECT -3.545 -4.295 -3.445 -3.875 ;
      RECT -3.545 0.465 -3.445 1.065 ;
      RECT -4.625 -103.41 -3.54 -103.31 ;
      RECT -4.625 -100.18 -3.54 -100.08 ;
      RECT -4.625 -90.49 -3.54 -90.39 ;
      RECT -4.625 -87.26 -3.54 -87.16 ;
      RECT -4.625 -77.57 -3.54 -77.47 ;
      RECT -4.625 -74.34 -3.54 -74.24 ;
      RECT -4.625 -64.65 -3.54 -64.55 ;
      RECT -4.625 -61.42 -3.54 -61.32 ;
      RECT -4.625 -51.73 -3.54 -51.63 ;
      RECT -4.625 -48.5 -3.54 -48.4 ;
      RECT -4.625 -38.81 -3.54 -38.71 ;
      RECT -4.625 -35.58 -3.54 -35.48 ;
      RECT -4.625 -25.89 -3.54 -25.79 ;
      RECT -4.625 -22.66 -3.54 -22.56 ;
      RECT -4.625 -12.97 -3.54 -12.87 ;
      RECT -4.625 -9.74 -3.54 -9.64 ;
      RECT -4.625 -0.05 -3.54 0.05 ;
      RECT -4.065 -107.655 -3.965 -107.055 ;
      RECT -4.065 -102.895 -3.965 -102.295 ;
      RECT -4.065 -101.195 -3.965 -100.595 ;
      RECT -4.065 -96.435 -3.965 -95.835 ;
      RECT -4.065 -94.735 -3.965 -94.135 ;
      RECT -4.065 -89.975 -3.965 -89.375 ;
      RECT -4.065 -88.275 -3.965 -87.675 ;
      RECT -4.065 -83.515 -3.965 -82.915 ;
      RECT -4.065 -81.815 -3.965 -81.215 ;
      RECT -4.065 -77.055 -3.965 -76.455 ;
      RECT -4.065 -75.355 -3.965 -74.755 ;
      RECT -4.065 -70.595 -3.965 -69.995 ;
      RECT -4.065 -68.895 -3.965 -68.295 ;
      RECT -4.065 -64.135 -3.965 -63.535 ;
      RECT -4.065 -62.435 -3.965 -61.835 ;
      RECT -4.065 -57.675 -3.965 -57.075 ;
      RECT -4.065 -55.975 -3.965 -55.375 ;
      RECT -4.065 -51.215 -3.965 -50.615 ;
      RECT -4.065 -49.515 -3.965 -48.915 ;
      RECT -4.065 -44.755 -3.965 -44.155 ;
      RECT -4.065 -43.055 -3.965 -42.455 ;
      RECT -4.065 -38.295 -3.965 -37.695 ;
      RECT -4.065 -36.595 -3.965 -35.995 ;
      RECT -4.065 -31.835 -3.965 -31.235 ;
      RECT -4.065 -30.135 -3.965 -29.535 ;
      RECT -4.065 -25.375 -3.965 -24.775 ;
      RECT -4.065 -23.675 -3.965 -23.075 ;
      RECT -4.065 -18.915 -3.965 -18.315 ;
      RECT -4.065 -17.215 -3.965 -16.615 ;
      RECT -4.065 -12.455 -3.965 -11.855 ;
      RECT -4.065 -10.755 -3.965 -10.155 ;
      RECT -4.065 -5.995 -3.965 -5.395 ;
      RECT -4.065 -4.295 -3.965 -3.695 ;
      RECT -4.065 0.465 -3.965 1.065 ;
      RECT -6.185 -104.215 -4.06 -104.115 ;
      RECT -6.185 -98.055 -4.06 -97.955 ;
      RECT -6.185 -92.615 -4.06 -92.515 ;
      RECT -6.185 -85.135 -4.06 -85.035 ;
      RECT -6.185 -79.695 -4.06 -79.595 ;
      RECT -6.185 -72.215 -4.06 -72.115 ;
      RECT -6.185 -66.775 -4.06 -66.675 ;
      RECT -6.185 -59.295 -4.06 -59.195 ;
      RECT -6.185 -53.855 -4.06 -53.755 ;
      RECT -6.185 -46.375 -4.06 -46.275 ;
      RECT -6.185 -40.935 -4.06 -40.835 ;
      RECT -6.185 -33.455 -4.06 -33.355 ;
      RECT -6.185 -28.015 -4.06 -27.915 ;
      RECT -6.185 -20.535 -4.06 -20.435 ;
      RECT -6.185 -15.095 -4.06 -14.995 ;
      RECT -6.185 -7.615 -4.06 -7.515 ;
      RECT -6.185 -2.175 -4.06 -2.075 ;
      RECT -4.325 -107.655 -4.225 -107.055 ;
      RECT -4.325 -96.435 -4.225 -95.835 ;
      RECT -4.325 -94.735 -4.225 -94.135 ;
      RECT -4.325 -83.515 -4.225 -82.915 ;
      RECT -4.325 -81.815 -4.225 -81.215 ;
      RECT -4.325 -70.595 -4.225 -69.995 ;
      RECT -4.325 -68.895 -4.225 -68.295 ;
      RECT -4.325 -57.675 -4.225 -57.075 ;
      RECT -4.325 -55.975 -4.225 -55.375 ;
      RECT -4.325 -44.755 -4.225 -44.155 ;
      RECT -4.325 -43.055 -4.225 -42.455 ;
      RECT -4.325 -31.835 -4.225 -31.235 ;
      RECT -4.325 -30.135 -4.225 -29.535 ;
      RECT -4.325 -18.915 -4.225 -18.315 ;
      RECT -4.325 -17.215 -4.225 -16.615 ;
      RECT -4.325 -5.995 -4.225 -5.395 ;
      RECT -4.325 -4.295 -4.225 -3.695 ;
      RECT -4.585 -102.895 -4.485 -102.295 ;
      RECT -4.585 -101.195 -4.485 -100.595 ;
      RECT -4.585 -89.975 -4.485 -89.375 ;
      RECT -4.585 -88.275 -4.485 -87.675 ;
      RECT -4.585 -77.055 -4.485 -76.455 ;
      RECT -4.585 -75.355 -4.485 -74.755 ;
      RECT -4.585 -64.135 -4.485 -63.535 ;
      RECT -4.585 -62.435 -4.485 -61.835 ;
      RECT -4.585 -51.215 -4.485 -50.615 ;
      RECT -4.585 -49.515 -4.485 -48.915 ;
      RECT -4.585 -38.295 -4.485 -37.695 ;
      RECT -4.585 -36.595 -4.485 -35.995 ;
      RECT -4.585 -25.375 -4.485 -24.775 ;
      RECT -4.585 -23.675 -4.485 -23.075 ;
      RECT -4.585 -12.455 -4.485 -11.855 ;
      RECT -4.585 -10.755 -4.485 -10.155 ;
      RECT -4.585 0.465 -4.485 1.065 ;
      RECT -4.845 -107.655 -4.745 -107.235 ;
      RECT -4.845 -102.895 -4.745 -102.295 ;
      RECT -4.845 -101.195 -4.745 -100.595 ;
      RECT -4.845 -96.255 -4.745 -95.835 ;
      RECT -4.845 -94.735 -4.745 -94.315 ;
      RECT -4.845 -89.975 -4.745 -89.375 ;
      RECT -4.845 -88.275 -4.745 -87.675 ;
      RECT -4.845 -83.335 -4.745 -82.915 ;
      RECT -4.845 -81.815 -4.745 -81.395 ;
      RECT -4.845 -77.055 -4.745 -76.455 ;
      RECT -4.845 -75.355 -4.745 -74.755 ;
      RECT -4.845 -70.415 -4.745 -69.995 ;
      RECT -4.845 -68.895 -4.745 -68.475 ;
      RECT -4.845 -64.135 -4.745 -63.535 ;
      RECT -4.845 -62.435 -4.745 -61.835 ;
      RECT -4.845 -57.495 -4.745 -57.075 ;
      RECT -4.845 -55.975 -4.745 -55.555 ;
      RECT -4.845 -51.215 -4.745 -50.615 ;
      RECT -4.845 -49.515 -4.745 -48.915 ;
      RECT -4.845 -44.575 -4.745 -44.155 ;
      RECT -4.845 -43.055 -4.745 -42.635 ;
      RECT -4.845 -38.295 -4.745 -37.695 ;
      RECT -4.845 -36.595 -4.745 -35.995 ;
      RECT -4.845 -31.655 -4.745 -31.235 ;
      RECT -4.845 -30.135 -4.745 -29.715 ;
      RECT -4.845 -25.375 -4.745 -24.775 ;
      RECT -4.845 -23.675 -4.745 -23.075 ;
      RECT -4.845 -18.735 -4.745 -18.315 ;
      RECT -4.845 -17.215 -4.745 -16.795 ;
      RECT -4.845 -12.455 -4.745 -11.855 ;
      RECT -4.845 -10.755 -4.745 -10.155 ;
      RECT -4.845 -5.815 -4.745 -5.395 ;
      RECT -4.845 -4.295 -4.745 -3.875 ;
      RECT -4.845 0.465 -4.745 1.065 ;
      RECT -5.925 -103.41 -4.84 -103.31 ;
      RECT -5.925 -100.18 -4.84 -100.08 ;
      RECT -5.925 -90.49 -4.84 -90.39 ;
      RECT -5.925 -87.26 -4.84 -87.16 ;
      RECT -5.925 -77.57 -4.84 -77.47 ;
      RECT -5.925 -74.34 -4.84 -74.24 ;
      RECT -5.925 -64.65 -4.84 -64.55 ;
      RECT -5.925 -61.42 -4.84 -61.32 ;
      RECT -5.925 -51.73 -4.84 -51.63 ;
      RECT -5.925 -48.5 -4.84 -48.4 ;
      RECT -5.925 -38.81 -4.84 -38.71 ;
      RECT -5.925 -35.58 -4.84 -35.48 ;
      RECT -5.925 -25.89 -4.84 -25.79 ;
      RECT -5.925 -22.66 -4.84 -22.56 ;
      RECT -5.925 -12.97 -4.84 -12.87 ;
      RECT -5.925 -9.74 -4.84 -9.64 ;
      RECT -5.925 -0.05 -4.84 0.05 ;
      RECT -5.365 -107.655 -5.265 -107.055 ;
      RECT -5.365 -102.895 -5.265 -102.295 ;
      RECT -5.365 -101.195 -5.265 -100.595 ;
      RECT -5.365 -96.435 -5.265 -95.835 ;
      RECT -5.365 -94.735 -5.265 -94.135 ;
      RECT -5.365 -89.975 -5.265 -89.375 ;
      RECT -5.365 -88.275 -5.265 -87.675 ;
      RECT -5.365 -83.515 -5.265 -82.915 ;
      RECT -5.365 -81.815 -5.265 -81.215 ;
      RECT -5.365 -77.055 -5.265 -76.455 ;
      RECT -5.365 -75.355 -5.265 -74.755 ;
      RECT -5.365 -70.595 -5.265 -69.995 ;
      RECT -5.365 -68.895 -5.265 -68.295 ;
      RECT -5.365 -64.135 -5.265 -63.535 ;
      RECT -5.365 -62.435 -5.265 -61.835 ;
      RECT -5.365 -57.675 -5.265 -57.075 ;
      RECT -5.365 -55.975 -5.265 -55.375 ;
      RECT -5.365 -51.215 -5.265 -50.615 ;
      RECT -5.365 -49.515 -5.265 -48.915 ;
      RECT -5.365 -44.755 -5.265 -44.155 ;
      RECT -5.365 -43.055 -5.265 -42.455 ;
      RECT -5.365 -38.295 -5.265 -37.695 ;
      RECT -5.365 -36.595 -5.265 -35.995 ;
      RECT -5.365 -31.835 -5.265 -31.235 ;
      RECT -5.365 -30.135 -5.265 -29.535 ;
      RECT -5.365 -25.375 -5.265 -24.775 ;
      RECT -5.365 -23.675 -5.265 -23.075 ;
      RECT -5.365 -18.915 -5.265 -18.315 ;
      RECT -5.365 -17.215 -5.265 -16.615 ;
      RECT -5.365 -12.455 -5.265 -11.855 ;
      RECT -5.365 -10.755 -5.265 -10.155 ;
      RECT -5.365 -5.995 -5.265 -5.395 ;
      RECT -5.365 -4.295 -5.265 -3.695 ;
      RECT -5.365 0.465 -5.265 1.065 ;
      RECT -7.485 -103.775 -5.36 -103.675 ;
      RECT -12.685 -99.815 -5.36 -99.715 ;
      RECT -12.685 -90.855 -5.36 -90.755 ;
      RECT -12.685 -86.895 -5.36 -86.795 ;
      RECT -12.685 -77.935 -5.36 -77.835 ;
      RECT -12.685 -73.975 -5.36 -73.875 ;
      RECT -12.685 -65.015 -5.36 -64.915 ;
      RECT -12.685 -61.055 -5.36 -60.955 ;
      RECT -12.685 -52.095 -5.36 -51.995 ;
      RECT -12.685 -48.135 -5.36 -48.035 ;
      RECT -12.685 -39.175 -5.36 -39.075 ;
      RECT -12.685 -35.215 -5.36 -35.115 ;
      RECT -12.685 -26.255 -5.36 -26.155 ;
      RECT -12.685 -22.295 -5.36 -22.195 ;
      RECT -12.685 -13.335 -5.36 -13.235 ;
      RECT -12.685 -9.375 -5.36 -9.275 ;
      RECT -12.685 -0.415 -5.36 -0.315 ;
      RECT -5.625 -107.655 -5.525 -107.055 ;
      RECT -5.625 -96.435 -5.525 -95.835 ;
      RECT -5.625 -94.735 -5.525 -94.135 ;
      RECT -5.625 -83.515 -5.525 -82.915 ;
      RECT -5.625 -81.815 -5.525 -81.215 ;
      RECT -5.625 -70.595 -5.525 -69.995 ;
      RECT -5.625 -68.895 -5.525 -68.295 ;
      RECT -5.625 -57.675 -5.525 -57.075 ;
      RECT -5.625 -55.975 -5.525 -55.375 ;
      RECT -5.625 -44.755 -5.525 -44.155 ;
      RECT -5.625 -43.055 -5.525 -42.455 ;
      RECT -5.625 -31.835 -5.525 -31.235 ;
      RECT -5.625 -30.135 -5.525 -29.535 ;
      RECT -5.625 -18.915 -5.525 -18.315 ;
      RECT -5.625 -17.215 -5.525 -16.615 ;
      RECT -5.625 -5.995 -5.525 -5.395 ;
      RECT -5.625 -4.295 -5.525 -3.695 ;
      RECT -5.885 -102.895 -5.785 -102.295 ;
      RECT -5.885 -101.195 -5.785 -100.595 ;
      RECT -5.885 -89.975 -5.785 -89.375 ;
      RECT -5.885 -88.275 -5.785 -87.675 ;
      RECT -5.885 -77.055 -5.785 -76.455 ;
      RECT -5.885 -75.355 -5.785 -74.755 ;
      RECT -5.885 -64.135 -5.785 -63.535 ;
      RECT -5.885 -62.435 -5.785 -61.835 ;
      RECT -5.885 -51.215 -5.785 -50.615 ;
      RECT -5.885 -49.515 -5.785 -48.915 ;
      RECT -5.885 -38.295 -5.785 -37.695 ;
      RECT -5.885 -36.595 -5.785 -35.995 ;
      RECT -5.885 -25.375 -5.785 -24.775 ;
      RECT -5.885 -23.675 -5.785 -23.075 ;
      RECT -5.885 -12.455 -5.785 -11.855 ;
      RECT -5.885 -10.755 -5.785 -10.155 ;
      RECT -5.885 0.465 -5.785 1.065 ;
      RECT -6.145 -107.655 -6.045 -107.235 ;
      RECT -6.145 -102.895 -6.045 -102.295 ;
      RECT -6.145 -101.195 -6.045 -100.595 ;
      RECT -6.145 -96.255 -6.045 -95.835 ;
      RECT -6.145 -94.735 -6.045 -94.315 ;
      RECT -6.145 -89.975 -6.045 -89.375 ;
      RECT -6.145 -88.275 -6.045 -87.675 ;
      RECT -6.145 -83.335 -6.045 -82.915 ;
      RECT -6.145 -81.815 -6.045 -81.395 ;
      RECT -6.145 -77.055 -6.045 -76.455 ;
      RECT -6.145 -75.355 -6.045 -74.755 ;
      RECT -6.145 -70.415 -6.045 -69.995 ;
      RECT -6.145 -68.895 -6.045 -68.475 ;
      RECT -6.145 -64.135 -6.045 -63.535 ;
      RECT -6.145 -62.435 -6.045 -61.835 ;
      RECT -6.145 -57.495 -6.045 -57.075 ;
      RECT -6.145 -55.975 -6.045 -55.555 ;
      RECT -6.145 -51.215 -6.045 -50.615 ;
      RECT -6.145 -49.515 -6.045 -48.915 ;
      RECT -6.145 -44.575 -6.045 -44.155 ;
      RECT -6.145 -43.055 -6.045 -42.635 ;
      RECT -6.145 -38.295 -6.045 -37.695 ;
      RECT -6.145 -36.595 -6.045 -35.995 ;
      RECT -6.145 -31.655 -6.045 -31.235 ;
      RECT -6.145 -30.135 -6.045 -29.715 ;
      RECT -6.145 -25.375 -6.045 -24.775 ;
      RECT -6.145 -23.675 -6.045 -23.075 ;
      RECT -6.145 -18.735 -6.045 -18.315 ;
      RECT -6.145 -17.215 -6.045 -16.795 ;
      RECT -6.145 -12.455 -6.045 -11.855 ;
      RECT -6.145 -10.755 -6.045 -10.155 ;
      RECT -6.145 -5.815 -6.045 -5.395 ;
      RECT -6.145 -4.295 -6.045 -3.875 ;
      RECT -6.145 0.465 -6.045 1.065 ;
      RECT -6.665 -107.655 -6.565 -107.055 ;
      RECT -6.665 -96.435 -6.565 -95.835 ;
      RECT -6.665 -94.735 -6.565 -94.135 ;
      RECT -6.665 -83.515 -6.565 -82.915 ;
      RECT -6.665 -81.815 -6.565 -81.215 ;
      RECT -6.665 -70.595 -6.565 -69.995 ;
      RECT -6.665 -68.895 -6.565 -68.295 ;
      RECT -6.665 -57.675 -6.565 -57.075 ;
      RECT -6.665 -55.975 -6.565 -55.375 ;
      RECT -6.665 -44.755 -6.565 -44.155 ;
      RECT -6.665 -43.055 -6.565 -42.455 ;
      RECT -6.665 -31.835 -6.565 -31.235 ;
      RECT -6.665 -30.135 -6.565 -29.535 ;
      RECT -6.665 -18.915 -6.565 -18.315 ;
      RECT -6.665 -17.215 -6.565 -16.615 ;
      RECT -6.665 -5.995 -6.565 -5.395 ;
      RECT -6.665 -4.295 -6.565 -3.695 ;
      RECT -7.485 -98.495 -6.66 -98.395 ;
      RECT -7.485 -92.175 -6.66 -92.075 ;
      RECT -7.485 -85.575 -6.66 -85.475 ;
      RECT -7.485 -79.255 -6.66 -79.155 ;
      RECT -7.485 -72.655 -6.66 -72.555 ;
      RECT -7.485 -66.335 -6.66 -66.235 ;
      RECT -7.485 -59.735 -6.66 -59.635 ;
      RECT -7.485 -53.415 -6.66 -53.315 ;
      RECT -7.485 -46.815 -6.66 -46.715 ;
      RECT -7.485 -40.495 -6.66 -40.395 ;
      RECT -7.485 -33.895 -6.66 -33.795 ;
      RECT -7.485 -27.575 -6.66 -27.475 ;
      RECT -7.485 -20.975 -6.66 -20.875 ;
      RECT -7.485 -14.655 -6.66 -14.555 ;
      RECT -7.485 -8.055 -6.66 -7.955 ;
      RECT -7.485 -1.735 -6.66 -1.635 ;
      RECT -6.925 -107.655 -6.825 -107.055 ;
      RECT -6.925 -96.435 -6.825 -95.835 ;
      RECT -6.925 -94.735 -6.825 -94.135 ;
      RECT -6.925 -83.515 -6.825 -82.915 ;
      RECT -6.925 -81.815 -6.825 -81.215 ;
      RECT -6.925 -70.595 -6.825 -69.995 ;
      RECT -6.925 -68.895 -6.825 -68.295 ;
      RECT -6.925 -57.675 -6.825 -57.075 ;
      RECT -6.925 -55.975 -6.825 -55.375 ;
      RECT -6.925 -44.755 -6.825 -44.155 ;
      RECT -6.925 -43.055 -6.825 -42.455 ;
      RECT -6.925 -31.835 -6.825 -31.235 ;
      RECT -6.925 -30.135 -6.825 -29.535 ;
      RECT -6.925 -18.915 -6.825 -18.315 ;
      RECT -6.925 -17.215 -6.825 -16.615 ;
      RECT -6.925 -5.995 -6.825 -5.395 ;
      RECT -6.925 -4.295 -6.825 -3.695 ;
      RECT -8.785 -98.055 -6.92 -97.955 ;
      RECT -8.785 -92.615 -6.92 -92.515 ;
      RECT -8.785 -85.135 -6.92 -85.035 ;
      RECT -8.785 -79.695 -6.92 -79.595 ;
      RECT -8.785 -72.215 -6.92 -72.115 ;
      RECT -8.785 -66.775 -6.92 -66.675 ;
      RECT -8.785 -59.295 -6.92 -59.195 ;
      RECT -8.785 -53.855 -6.92 -53.755 ;
      RECT -8.785 -46.375 -6.92 -46.275 ;
      RECT -8.785 -40.935 -6.92 -40.835 ;
      RECT -8.785 -33.455 -6.92 -33.355 ;
      RECT -8.785 -28.015 -6.92 -27.915 ;
      RECT -8.785 -20.535 -6.92 -20.435 ;
      RECT -8.785 -15.095 -6.92 -14.995 ;
      RECT -8.785 -7.615 -6.92 -7.515 ;
      RECT -8.785 -2.175 -6.92 -2.075 ;
      RECT -7.445 -107.655 -7.345 -107.235 ;
      RECT -7.445 -102.895 -7.345 -102.295 ;
      RECT -7.445 -101.195 -7.345 -100.595 ;
      RECT -7.445 -96.255 -7.345 -95.835 ;
      RECT -7.445 -94.735 -7.345 -94.315 ;
      RECT -7.445 -89.975 -7.345 -89.375 ;
      RECT -7.445 -88.275 -7.345 -87.675 ;
      RECT -7.445 -83.335 -7.345 -82.915 ;
      RECT -7.445 -81.815 -7.345 -81.395 ;
      RECT -7.445 -77.055 -7.345 -76.455 ;
      RECT -7.445 -75.355 -7.345 -74.755 ;
      RECT -7.445 -70.415 -7.345 -69.995 ;
      RECT -7.445 -68.895 -7.345 -68.475 ;
      RECT -7.445 -64.135 -7.345 -63.535 ;
      RECT -7.445 -62.435 -7.345 -61.835 ;
      RECT -7.445 -57.495 -7.345 -57.075 ;
      RECT -7.445 -55.975 -7.345 -55.555 ;
      RECT -7.445 -51.215 -7.345 -50.615 ;
      RECT -7.445 -49.515 -7.345 -48.915 ;
      RECT -7.445 -44.575 -7.345 -44.155 ;
      RECT -7.445 -43.055 -7.345 -42.635 ;
      RECT -7.445 -38.295 -7.345 -37.695 ;
      RECT -7.445 -36.595 -7.345 -35.995 ;
      RECT -7.445 -31.655 -7.345 -31.235 ;
      RECT -7.445 -30.135 -7.345 -29.715 ;
      RECT -7.445 -25.375 -7.345 -24.775 ;
      RECT -7.445 -23.675 -7.345 -23.075 ;
      RECT -7.445 -18.735 -7.345 -18.315 ;
      RECT -7.445 -17.215 -7.345 -16.795 ;
      RECT -7.445 -12.455 -7.345 -11.855 ;
      RECT -7.445 -10.755 -7.345 -10.155 ;
      RECT -7.445 -5.815 -7.345 -5.395 ;
      RECT -7.445 -4.295 -7.345 -3.875 ;
      RECT -7.445 0.465 -7.345 1.065 ;
      RECT -7.965 -107.655 -7.865 -107.055 ;
      RECT -7.965 -96.435 -7.865 -95.835 ;
      RECT -7.965 -94.735 -7.865 -94.135 ;
      RECT -7.965 -83.515 -7.865 -82.915 ;
      RECT -7.965 -81.815 -7.865 -81.215 ;
      RECT -7.965 -70.595 -7.865 -69.995 ;
      RECT -7.965 -68.895 -7.865 -68.295 ;
      RECT -7.965 -57.675 -7.865 -57.075 ;
      RECT -7.965 -55.975 -7.865 -55.375 ;
      RECT -7.965 -44.755 -7.865 -44.155 ;
      RECT -7.965 -43.055 -7.865 -42.455 ;
      RECT -7.965 -31.835 -7.865 -31.235 ;
      RECT -7.965 -30.135 -7.865 -29.535 ;
      RECT -7.965 -18.915 -7.865 -18.315 ;
      RECT -7.965 -17.215 -7.865 -16.615 ;
      RECT -7.965 -5.995 -7.865 -5.395 ;
      RECT -7.965 -4.295 -7.865 -3.695 ;
      RECT -10.085 -98.275 -7.96 -98.175 ;
      RECT -10.085 -92.395 -7.96 -92.295 ;
      RECT -10.085 -85.355 -7.96 -85.255 ;
      RECT -10.085 -79.475 -7.96 -79.375 ;
      RECT -10.085 -72.435 -7.96 -72.335 ;
      RECT -10.085 -66.555 -7.96 -66.455 ;
      RECT -10.085 -59.515 -7.96 -59.415 ;
      RECT -10.085 -53.635 -7.96 -53.535 ;
      RECT -10.085 -46.595 -7.96 -46.495 ;
      RECT -10.085 -40.715 -7.96 -40.615 ;
      RECT -10.085 -33.675 -7.96 -33.575 ;
      RECT -10.085 -27.795 -7.96 -27.695 ;
      RECT -10.085 -20.755 -7.96 -20.655 ;
      RECT -10.085 -14.875 -7.96 -14.775 ;
      RECT -10.085 -7.835 -7.96 -7.735 ;
      RECT -10.085 -1.955 -7.96 -1.855 ;
      RECT -8.225 -107.655 -8.125 -107.055 ;
      RECT -8.225 -96.435 -8.125 -95.835 ;
      RECT -8.225 -94.735 -8.125 -94.135 ;
      RECT -8.225 -83.515 -8.125 -82.915 ;
      RECT -8.225 -81.815 -8.125 -81.215 ;
      RECT -8.225 -70.595 -8.125 -69.995 ;
      RECT -8.225 -68.895 -8.125 -68.295 ;
      RECT -8.225 -57.675 -8.125 -57.075 ;
      RECT -8.225 -55.975 -8.125 -55.375 ;
      RECT -8.225 -44.755 -8.125 -44.155 ;
      RECT -8.225 -43.055 -8.125 -42.455 ;
      RECT -8.225 -31.835 -8.125 -31.235 ;
      RECT -8.225 -30.135 -8.125 -29.535 ;
      RECT -8.225 -18.915 -8.125 -18.315 ;
      RECT -8.225 -17.215 -8.125 -16.615 ;
      RECT -8.225 -5.995 -8.125 -5.395 ;
      RECT -8.225 -4.295 -8.125 -3.695 ;
      RECT -12.645 -103.335 -8.22 -103.235 ;
      RECT -11.385 -98.495 -8.22 -98.395 ;
      RECT -11.385 -92.175 -8.22 -92.075 ;
      RECT -11.385 -85.575 -8.22 -85.475 ;
      RECT -11.385 -79.255 -8.22 -79.155 ;
      RECT -11.385 -72.655 -8.22 -72.555 ;
      RECT -11.385 -66.335 -8.22 -66.235 ;
      RECT -11.385 -59.735 -8.22 -59.635 ;
      RECT -11.385 -53.415 -8.22 -53.315 ;
      RECT -11.385 -46.815 -8.22 -46.715 ;
      RECT -11.385 -40.495 -8.22 -40.395 ;
      RECT -11.385 -33.895 -8.22 -33.795 ;
      RECT -11.385 -27.575 -8.22 -27.475 ;
      RECT -11.385 -20.975 -8.22 -20.875 ;
      RECT -11.385 -14.655 -8.22 -14.555 ;
      RECT -11.385 -8.055 -8.22 -7.955 ;
      RECT -11.385 -1.735 -8.22 -1.635 ;
      RECT -8.745 -107.655 -8.645 -107.235 ;
      RECT -8.745 -102.895 -8.645 -102.295 ;
      RECT -8.745 -101.195 -8.645 -100.595 ;
      RECT -8.745 -96.255 -8.645 -95.835 ;
      RECT -8.745 -94.735 -8.645 -94.315 ;
      RECT -8.745 -89.975 -8.645 -89.375 ;
      RECT -8.745 -88.275 -8.645 -87.675 ;
      RECT -8.745 -83.335 -8.645 -82.915 ;
      RECT -8.745 -81.815 -8.645 -81.395 ;
      RECT -8.745 -77.055 -8.645 -76.455 ;
      RECT -8.745 -75.355 -8.645 -74.755 ;
      RECT -8.745 -70.415 -8.645 -69.995 ;
      RECT -8.745 -68.895 -8.645 -68.475 ;
      RECT -8.745 -64.135 -8.645 -63.535 ;
      RECT -8.745 -62.435 -8.645 -61.835 ;
      RECT -8.745 -57.495 -8.645 -57.075 ;
      RECT -8.745 -55.975 -8.645 -55.555 ;
      RECT -8.745 -51.215 -8.645 -50.615 ;
      RECT -8.745 -49.515 -8.645 -48.915 ;
      RECT -8.745 -44.575 -8.645 -44.155 ;
      RECT -8.745 -43.055 -8.645 -42.635 ;
      RECT -8.745 -38.295 -8.645 -37.695 ;
      RECT -8.745 -36.595 -8.645 -35.995 ;
      RECT -8.745 -31.655 -8.645 -31.235 ;
      RECT -8.745 -30.135 -8.645 -29.715 ;
      RECT -8.745 -25.375 -8.645 -24.775 ;
      RECT -8.745 -23.675 -8.645 -23.075 ;
      RECT -8.745 -18.735 -8.645 -18.315 ;
      RECT -8.745 -17.215 -8.645 -16.795 ;
      RECT -8.745 -12.455 -8.645 -11.855 ;
      RECT -8.745 -10.755 -8.645 -10.155 ;
      RECT -8.745 -5.815 -8.645 -5.395 ;
      RECT -8.745 -4.295 -8.645 -3.875 ;
      RECT -8.745 0.465 -8.645 1.065 ;
      RECT -9.265 -107.655 -9.165 -107.055 ;
      RECT -9.265 -96.435 -9.165 -95.835 ;
      RECT -9.265 -94.735 -9.165 -94.135 ;
      RECT -9.265 -83.515 -9.165 -82.915 ;
      RECT -9.265 -81.815 -9.165 -81.215 ;
      RECT -9.265 -70.595 -9.165 -69.995 ;
      RECT -9.265 -68.895 -9.165 -68.295 ;
      RECT -9.265 -57.675 -9.165 -57.075 ;
      RECT -9.265 -55.975 -9.165 -55.375 ;
      RECT -9.265 -44.755 -9.165 -44.155 ;
      RECT -9.265 -43.055 -9.165 -42.455 ;
      RECT -9.265 -31.835 -9.165 -31.235 ;
      RECT -9.265 -30.135 -9.165 -29.535 ;
      RECT -9.265 -18.915 -9.165 -18.315 ;
      RECT -9.265 -17.215 -9.165 -16.615 ;
      RECT -9.265 -5.995 -9.165 -5.395 ;
      RECT -9.265 -4.295 -9.165 -3.695 ;
      RECT -12.645 -103.775 -9.26 -103.675 ;
      RECT -35.845 -47.035 -9.26 -46.935 ;
      RECT -35.845 -40.275 -9.26 -40.175 ;
      RECT -35.845 -34.115 -9.26 -34.015 ;
      RECT -35.845 -27.355 -9.26 -27.255 ;
      RECT -35.845 -21.195 -9.26 -21.095 ;
      RECT -35.845 -14.435 -9.26 -14.335 ;
      RECT -35.845 -8.275 -9.26 -8.175 ;
      RECT -35.845 -1.515 -9.26 -1.415 ;
      RECT -9.525 -107.655 -9.425 -107.055 ;
      RECT -9.525 -96.435 -9.425 -95.835 ;
      RECT -9.525 -94.735 -9.425 -94.135 ;
      RECT -9.525 -83.515 -9.425 -82.915 ;
      RECT -9.525 -81.815 -9.425 -81.215 ;
      RECT -9.525 -70.595 -9.425 -69.995 ;
      RECT -9.525 -68.895 -9.425 -68.295 ;
      RECT -9.525 -57.675 -9.425 -57.075 ;
      RECT -9.525 -55.975 -9.425 -55.375 ;
      RECT -9.525 -44.755 -9.425 -44.155 ;
      RECT -9.525 -43.055 -9.425 -42.455 ;
      RECT -9.525 -31.835 -9.425 -31.235 ;
      RECT -9.525 -30.135 -9.425 -29.535 ;
      RECT -9.525 -18.915 -9.425 -18.315 ;
      RECT -9.525 -17.215 -9.425 -16.615 ;
      RECT -9.525 -5.995 -9.425 -5.395 ;
      RECT -9.525 -4.295 -9.425 -3.695 ;
      RECT -35.845 -73.095 -9.52 -72.995 ;
      RECT -35.845 -65.895 -9.52 -65.795 ;
      RECT -35.845 -60.175 -9.52 -60.075 ;
      RECT -35.845 -52.975 -9.52 -52.875 ;
      RECT -35.845 -21.415 -9.52 -21.315 ;
      RECT -35.845 -14.215 -9.52 -14.115 ;
      RECT -35.845 -8.495 -9.52 -8.395 ;
      RECT -35.845 -1.295 -9.52 -1.195 ;
      RECT -10.045 -107.655 -9.945 -107.235 ;
      RECT -10.045 -102.895 -9.945 -102.295 ;
      RECT -10.045 -101.195 -9.945 -100.595 ;
      RECT -10.045 -96.255 -9.945 -95.835 ;
      RECT -10.045 -94.735 -9.945 -94.315 ;
      RECT -10.045 -89.975 -9.945 -89.375 ;
      RECT -10.045 -88.275 -9.945 -87.675 ;
      RECT -10.045 -83.335 -9.945 -82.915 ;
      RECT -10.045 -81.815 -9.945 -81.395 ;
      RECT -10.045 -77.055 -9.945 -76.455 ;
      RECT -10.045 -75.355 -9.945 -74.755 ;
      RECT -10.045 -70.415 -9.945 -69.995 ;
      RECT -10.045 -68.895 -9.945 -68.475 ;
      RECT -10.045 -64.135 -9.945 -63.535 ;
      RECT -10.045 -62.435 -9.945 -61.835 ;
      RECT -10.045 -57.495 -9.945 -57.075 ;
      RECT -10.045 -55.975 -9.945 -55.555 ;
      RECT -10.045 -51.215 -9.945 -50.615 ;
      RECT -10.045 -49.515 -9.945 -48.915 ;
      RECT -10.045 -44.575 -9.945 -44.155 ;
      RECT -10.045 -43.055 -9.945 -42.635 ;
      RECT -10.045 -38.295 -9.945 -37.695 ;
      RECT -10.045 -36.595 -9.945 -35.995 ;
      RECT -10.045 -31.655 -9.945 -31.235 ;
      RECT -10.045 -30.135 -9.945 -29.715 ;
      RECT -10.045 -25.375 -9.945 -24.775 ;
      RECT -10.045 -23.675 -9.945 -23.075 ;
      RECT -10.045 -18.735 -9.945 -18.315 ;
      RECT -10.045 -17.215 -9.945 -16.795 ;
      RECT -10.045 -12.455 -9.945 -11.855 ;
      RECT -10.045 -10.755 -9.945 -10.155 ;
      RECT -10.045 -5.815 -9.945 -5.395 ;
      RECT -10.045 -4.295 -9.945 -3.875 ;
      RECT -10.045 0.465 -9.945 1.065 ;
      RECT -10.565 -107.655 -10.465 -107.055 ;
      RECT -10.565 -96.435 -10.465 -95.835 ;
      RECT -10.565 -94.735 -10.465 -94.135 ;
      RECT -10.565 -83.515 -10.465 -82.915 ;
      RECT -10.565 -81.815 -10.465 -81.215 ;
      RECT -10.565 -70.595 -10.465 -69.995 ;
      RECT -10.565 -68.895 -10.465 -68.295 ;
      RECT -10.565 -57.675 -10.465 -57.075 ;
      RECT -10.565 -55.975 -10.465 -55.375 ;
      RECT -10.565 -44.755 -10.465 -44.155 ;
      RECT -10.565 -43.055 -10.465 -42.455 ;
      RECT -10.565 -31.835 -10.465 -31.235 ;
      RECT -10.565 -30.135 -10.465 -29.535 ;
      RECT -10.565 -18.915 -10.465 -18.315 ;
      RECT -10.565 -17.215 -10.465 -16.615 ;
      RECT -10.565 -5.995 -10.465 -5.395 ;
      RECT -10.565 -4.295 -10.465 -3.695 ;
      RECT -35.845 -86.235 -10.56 -86.135 ;
      RECT -35.845 -78.595 -10.56 -78.495 ;
      RECT -35.845 -60.395 -10.56 -60.295 ;
      RECT -35.845 -52.755 -10.56 -52.655 ;
      RECT -35.845 -34.555 -10.56 -34.455 ;
      RECT -35.845 -26.915 -10.56 -26.815 ;
      RECT -35.845 -8.715 -10.56 -8.615 ;
      RECT -35.845 -1.075 -10.56 -0.975 ;
      RECT -10.825 -107.655 -10.725 -107.055 ;
      RECT -10.825 -96.435 -10.725 -95.835 ;
      RECT -10.825 -94.735 -10.725 -94.135 ;
      RECT -10.825 -83.515 -10.725 -82.915 ;
      RECT -10.825 -81.815 -10.725 -81.215 ;
      RECT -10.825 -70.595 -10.725 -69.995 ;
      RECT -10.825 -68.895 -10.725 -68.295 ;
      RECT -10.825 -57.675 -10.725 -57.075 ;
      RECT -10.825 -55.975 -10.725 -55.375 ;
      RECT -10.825 -44.755 -10.725 -44.155 ;
      RECT -10.825 -43.055 -10.725 -42.455 ;
      RECT -10.825 -31.835 -10.725 -31.235 ;
      RECT -10.825 -30.135 -10.725 -29.535 ;
      RECT -10.825 -18.915 -10.725 -18.315 ;
      RECT -10.825 -17.215 -10.725 -16.615 ;
      RECT -10.825 -5.995 -10.725 -5.395 ;
      RECT -10.825 -4.295 -10.725 -3.695 ;
      RECT -35.845 -91.295 -10.82 -91.195 ;
      RECT -35.845 -78.375 -10.82 -78.275 ;
      RECT -35.845 -65.455 -10.82 -65.355 ;
      RECT -35.845 -52.535 -10.82 -52.435 ;
      RECT -35.845 -39.615 -10.82 -39.515 ;
      RECT -35.845 -26.695 -10.82 -26.595 ;
      RECT -35.845 -13.775 -10.82 -13.675 ;
      RECT -35.845 -0.855 -10.82 -0.755 ;
      RECT -11.345 -101.195 -11.245 -100.595 ;
      RECT -11.345 -96.255 -11.245 -95.835 ;
      RECT -11.345 -94.735 -11.245 -94.315 ;
      RECT -11.345 -89.975 -11.245 -89.375 ;
      RECT -11.345 -88.275 -11.245 -87.675 ;
      RECT -11.345 -83.335 -11.245 -82.915 ;
      RECT -11.345 -81.815 -11.245 -81.395 ;
      RECT -11.345 -77.055 -11.245 -76.455 ;
      RECT -11.345 -75.355 -11.245 -74.755 ;
      RECT -11.345 -70.415 -11.245 -69.995 ;
      RECT -11.345 -68.895 -11.245 -68.475 ;
      RECT -11.345 -64.135 -11.245 -63.535 ;
      RECT -11.345 -62.435 -11.245 -61.835 ;
      RECT -11.345 -57.495 -11.245 -57.075 ;
      RECT -11.345 -55.975 -11.245 -55.555 ;
      RECT -11.345 -51.215 -11.245 -50.615 ;
      RECT -11.345 -49.515 -11.245 -48.915 ;
      RECT -11.345 -44.575 -11.245 -44.155 ;
      RECT -11.345 -43.055 -11.245 -42.635 ;
      RECT -11.345 -38.295 -11.245 -37.695 ;
      RECT -11.345 -36.595 -11.245 -35.995 ;
      RECT -11.345 -31.655 -11.245 -31.235 ;
      RECT -11.345 -30.135 -11.245 -29.715 ;
      RECT -11.345 -25.375 -11.245 -24.775 ;
      RECT -11.345 -23.675 -11.245 -23.075 ;
      RECT -11.345 -18.735 -11.245 -18.315 ;
      RECT -11.345 -17.215 -11.245 -16.795 ;
      RECT -11.345 -12.455 -11.245 -11.855 ;
      RECT -11.345 -10.755 -11.245 -10.155 ;
      RECT -11.345 -5.815 -11.245 -5.395 ;
      RECT -11.345 -4.295 -11.245 -3.875 ;
      RECT -11.345 0.465 -11.245 1.065 ;
      RECT -11.445 -110.635 -11.345 -110.155 ;
      RECT -11.445 -109.175 -11.345 -108.755 ;
      RECT -11.865 -96.435 -11.765 -95.835 ;
      RECT -11.865 -94.735 -11.765 -94.135 ;
      RECT -11.865 -83.515 -11.765 -82.915 ;
      RECT -11.865 -81.815 -11.765 -81.215 ;
      RECT -11.865 -70.595 -11.765 -69.995 ;
      RECT -11.865 -68.895 -11.765 -68.295 ;
      RECT -11.865 -57.675 -11.765 -57.075 ;
      RECT -11.865 -55.975 -11.765 -55.375 ;
      RECT -11.865 -44.755 -11.765 -44.155 ;
      RECT -11.865 -43.055 -11.765 -42.455 ;
      RECT -11.865 -31.835 -11.765 -31.235 ;
      RECT -11.865 -30.135 -11.765 -29.535 ;
      RECT -11.865 -18.915 -11.765 -18.315 ;
      RECT -11.865 -17.215 -11.765 -16.615 ;
      RECT -11.865 -5.995 -11.765 -5.395 ;
      RECT -11.865 -4.295 -11.765 -3.695 ;
      RECT -12.045 -110.635 -11.945 -110.155 ;
      RECT -12.045 -109.175 -11.945 -108.755 ;
      RECT -12.125 -96.435 -12.025 -95.835 ;
      RECT -12.125 -94.735 -12.025 -94.135 ;
      RECT -12.125 -83.515 -12.025 -82.915 ;
      RECT -12.125 -81.815 -12.025 -81.215 ;
      RECT -12.125 -70.595 -12.025 -69.995 ;
      RECT -12.125 -68.895 -12.025 -68.295 ;
      RECT -12.125 -57.675 -12.025 -57.075 ;
      RECT -12.125 -55.975 -12.025 -55.375 ;
      RECT -12.125 -44.755 -12.025 -44.155 ;
      RECT -12.125 -43.055 -12.025 -42.455 ;
      RECT -12.125 -31.835 -12.025 -31.235 ;
      RECT -12.125 -30.135 -12.025 -29.535 ;
      RECT -12.125 -18.915 -12.025 -18.315 ;
      RECT -12.125 -17.215 -12.025 -16.615 ;
      RECT -12.125 -5.995 -12.025 -5.395 ;
      RECT -12.125 -4.295 -12.025 -3.695 ;
      RECT -12.645 -101.195 -12.545 -100.595 ;
      RECT -12.645 -96.255 -12.545 -95.835 ;
      RECT -12.645 -94.735 -12.545 -94.315 ;
      RECT -12.645 -89.975 -12.545 -89.375 ;
      RECT -12.645 -88.275 -12.545 -87.675 ;
      RECT -12.645 -83.335 -12.545 -82.915 ;
      RECT -12.645 -81.815 -12.545 -81.395 ;
      RECT -12.645 -77.055 -12.545 -76.455 ;
      RECT -12.645 -75.355 -12.545 -74.755 ;
      RECT -12.645 -70.415 -12.545 -69.995 ;
      RECT -12.645 -68.895 -12.545 -68.475 ;
      RECT -12.645 -64.135 -12.545 -63.535 ;
      RECT -12.645 -62.435 -12.545 -61.835 ;
      RECT -12.645 -57.495 -12.545 -57.075 ;
      RECT -12.645 -55.975 -12.545 -55.555 ;
      RECT -12.645 -51.215 -12.545 -50.615 ;
      RECT -12.645 -49.515 -12.545 -48.915 ;
      RECT -12.645 -44.575 -12.545 -44.155 ;
      RECT -12.645 -43.055 -12.545 -42.635 ;
      RECT -12.645 -38.295 -12.545 -37.695 ;
      RECT -12.645 -36.595 -12.545 -35.995 ;
      RECT -12.645 -31.655 -12.545 -31.235 ;
      RECT -12.645 -30.135 -12.545 -29.715 ;
      RECT -12.645 -25.375 -12.545 -24.775 ;
      RECT -12.645 -23.675 -12.545 -23.075 ;
      RECT -12.645 -18.735 -12.545 -18.315 ;
      RECT -12.645 -17.215 -12.545 -16.795 ;
      RECT -12.645 -12.455 -12.545 -11.855 ;
      RECT -12.645 -10.755 -12.545 -10.155 ;
      RECT -12.645 -5.815 -12.545 -5.395 ;
      RECT -12.645 -4.295 -12.545 -3.875 ;
      RECT -12.645 0.465 -12.545 1.065 ;
      RECT -13.165 -96.435 -13.065 -95.835 ;
      RECT -13.165 -94.735 -13.065 -94.135 ;
      RECT -13.165 -83.515 -13.065 -82.915 ;
      RECT -13.165 -81.815 -13.065 -81.215 ;
      RECT -13.165 -70.595 -13.065 -69.995 ;
      RECT -13.165 -68.895 -13.065 -68.295 ;
      RECT -13.165 -57.675 -13.065 -57.075 ;
      RECT -13.165 -55.975 -13.065 -55.375 ;
      RECT -13.165 -44.755 -13.065 -44.155 ;
      RECT -13.165 -43.055 -13.065 -42.455 ;
      RECT -13.165 -31.835 -13.065 -31.235 ;
      RECT -13.165 -30.135 -13.065 -29.535 ;
      RECT -13.165 -18.915 -13.065 -18.315 ;
      RECT -13.165 -17.215 -13.065 -16.615 ;
      RECT -13.165 -5.995 -13.065 -5.395 ;
      RECT -13.165 -4.295 -13.065 -3.695 ;
      RECT -13.985 -98.495 -13.16 -98.395 ;
      RECT -13.985 -92.175 -13.16 -92.075 ;
      RECT -13.985 -85.575 -13.16 -85.475 ;
      RECT -13.985 -79.255 -13.16 -79.155 ;
      RECT -13.985 -72.655 -13.16 -72.555 ;
      RECT -13.985 -66.335 -13.16 -66.235 ;
      RECT -13.985 -59.735 -13.16 -59.635 ;
      RECT -13.985 -53.415 -13.16 -53.315 ;
      RECT -13.985 -46.815 -13.16 -46.715 ;
      RECT -13.985 -40.495 -13.16 -40.395 ;
      RECT -13.985 -33.895 -13.16 -33.795 ;
      RECT -13.985 -27.575 -13.16 -27.475 ;
      RECT -13.985 -20.975 -13.16 -20.875 ;
      RECT -13.985 -14.655 -13.16 -14.555 ;
      RECT -13.985 -8.055 -13.16 -7.955 ;
      RECT -13.985 -1.735 -13.16 -1.635 ;
      RECT -13.425 -96.435 -13.325 -95.835 ;
      RECT -13.425 -94.735 -13.325 -94.135 ;
      RECT -13.425 -83.515 -13.325 -82.915 ;
      RECT -13.425 -81.815 -13.325 -81.215 ;
      RECT -13.425 -70.595 -13.325 -69.995 ;
      RECT -13.425 -68.895 -13.325 -68.295 ;
      RECT -13.425 -57.675 -13.325 -57.075 ;
      RECT -13.425 -55.975 -13.325 -55.375 ;
      RECT -13.425 -44.755 -13.325 -44.155 ;
      RECT -13.425 -43.055 -13.325 -42.455 ;
      RECT -13.425 -31.835 -13.325 -31.235 ;
      RECT -13.425 -30.135 -13.325 -29.535 ;
      RECT -13.425 -18.915 -13.325 -18.315 ;
      RECT -13.425 -17.215 -13.325 -16.615 ;
      RECT -13.425 -5.995 -13.325 -5.395 ;
      RECT -13.425 -4.295 -13.325 -3.695 ;
      RECT -15.285 -98.055 -13.42 -97.955 ;
      RECT -15.285 -92.615 -13.42 -92.515 ;
      RECT -15.285 -85.135 -13.42 -85.035 ;
      RECT -15.285 -79.695 -13.42 -79.595 ;
      RECT -15.285 -72.215 -13.42 -72.115 ;
      RECT -15.285 -66.775 -13.42 -66.675 ;
      RECT -15.285 -59.295 -13.42 -59.195 ;
      RECT -15.285 -53.855 -13.42 -53.755 ;
      RECT -15.285 -46.375 -13.42 -46.275 ;
      RECT -15.285 -40.935 -13.42 -40.835 ;
      RECT -15.285 -33.455 -13.42 -33.355 ;
      RECT -15.285 -28.015 -13.42 -27.915 ;
      RECT -15.285 -20.535 -13.42 -20.435 ;
      RECT -15.285 -15.095 -13.42 -14.995 ;
      RECT -15.285 -7.615 -13.42 -7.515 ;
      RECT -15.285 -2.175 -13.42 -2.075 ;
      RECT -13.945 -101.195 -13.845 -100.595 ;
      RECT -13.945 -96.255 -13.845 -95.835 ;
      RECT -13.945 -94.735 -13.845 -94.315 ;
      RECT -13.945 -89.975 -13.845 -89.375 ;
      RECT -13.945 -88.275 -13.845 -87.675 ;
      RECT -13.945 -83.335 -13.845 -82.915 ;
      RECT -13.945 -81.815 -13.845 -81.395 ;
      RECT -13.945 -77.055 -13.845 -76.455 ;
      RECT -13.945 -75.355 -13.845 -74.755 ;
      RECT -13.945 -70.415 -13.845 -69.995 ;
      RECT -13.945 -68.895 -13.845 -68.475 ;
      RECT -13.945 -64.135 -13.845 -63.535 ;
      RECT -13.945 -62.435 -13.845 -61.835 ;
      RECT -13.945 -57.495 -13.845 -57.075 ;
      RECT -13.945 -55.975 -13.845 -55.555 ;
      RECT -13.945 -51.215 -13.845 -50.615 ;
      RECT -13.945 -49.515 -13.845 -48.915 ;
      RECT -13.945 -44.575 -13.845 -44.155 ;
      RECT -13.945 -43.055 -13.845 -42.635 ;
      RECT -13.945 -38.295 -13.845 -37.695 ;
      RECT -13.945 -36.595 -13.845 -35.995 ;
      RECT -13.945 -31.655 -13.845 -31.235 ;
      RECT -13.945 -30.135 -13.845 -29.715 ;
      RECT -13.945 -25.375 -13.845 -24.775 ;
      RECT -13.945 -23.675 -13.845 -23.075 ;
      RECT -13.945 -18.735 -13.845 -18.315 ;
      RECT -13.945 -17.215 -13.845 -16.795 ;
      RECT -13.945 -12.455 -13.845 -11.855 ;
      RECT -13.945 -10.755 -13.845 -10.155 ;
      RECT -13.945 -5.815 -13.845 -5.395 ;
      RECT -13.945 -4.295 -13.845 -3.875 ;
      RECT -13.945 0.465 -13.845 1.065 ;
      RECT -14.465 -96.435 -14.365 -95.835 ;
      RECT -14.465 -94.735 -14.365 -94.135 ;
      RECT -14.465 -83.515 -14.365 -82.915 ;
      RECT -14.465 -81.815 -14.365 -81.215 ;
      RECT -14.465 -70.595 -14.365 -69.995 ;
      RECT -14.465 -68.895 -14.365 -68.295 ;
      RECT -14.465 -57.675 -14.365 -57.075 ;
      RECT -14.465 -55.975 -14.365 -55.375 ;
      RECT -14.465 -44.755 -14.365 -44.155 ;
      RECT -14.465 -43.055 -14.365 -42.455 ;
      RECT -14.465 -31.835 -14.365 -31.235 ;
      RECT -14.465 -30.135 -14.365 -29.535 ;
      RECT -14.465 -18.915 -14.365 -18.315 ;
      RECT -14.465 -17.215 -14.365 -16.615 ;
      RECT -14.465 -5.995 -14.365 -5.395 ;
      RECT -14.465 -4.295 -14.365 -3.695 ;
      RECT -16.585 -98.275 -14.46 -98.175 ;
      RECT -16.585 -92.395 -14.46 -92.295 ;
      RECT -16.585 -85.355 -14.46 -85.255 ;
      RECT -16.585 -79.475 -14.46 -79.375 ;
      RECT -16.585 -72.435 -14.46 -72.335 ;
      RECT -16.585 -66.555 -14.46 -66.455 ;
      RECT -16.585 -59.515 -14.46 -59.415 ;
      RECT -16.585 -53.635 -14.46 -53.535 ;
      RECT -16.585 -46.595 -14.46 -46.495 ;
      RECT -16.585 -40.715 -14.46 -40.615 ;
      RECT -16.585 -33.675 -14.46 -33.575 ;
      RECT -16.585 -27.795 -14.46 -27.695 ;
      RECT -16.585 -20.755 -14.46 -20.655 ;
      RECT -16.585 -14.875 -14.46 -14.775 ;
      RECT -16.585 -7.835 -14.46 -7.735 ;
      RECT -16.585 -1.955 -14.46 -1.855 ;
      RECT -14.725 -96.435 -14.625 -95.835 ;
      RECT -14.725 -94.735 -14.625 -94.135 ;
      RECT -14.725 -83.515 -14.625 -82.915 ;
      RECT -14.725 -81.815 -14.625 -81.215 ;
      RECT -14.725 -70.595 -14.625 -69.995 ;
      RECT -14.725 -68.895 -14.625 -68.295 ;
      RECT -14.725 -57.675 -14.625 -57.075 ;
      RECT -14.725 -55.975 -14.625 -55.375 ;
      RECT -14.725 -44.755 -14.625 -44.155 ;
      RECT -14.725 -43.055 -14.625 -42.455 ;
      RECT -14.725 -31.835 -14.625 -31.235 ;
      RECT -14.725 -30.135 -14.625 -29.535 ;
      RECT -14.725 -18.915 -14.625 -18.315 ;
      RECT -14.725 -17.215 -14.625 -16.615 ;
      RECT -14.725 -5.995 -14.625 -5.395 ;
      RECT -14.725 -4.295 -14.625 -3.695 ;
      RECT -17.885 -98.495 -14.72 -98.395 ;
      RECT -17.885 -92.175 -14.72 -92.075 ;
      RECT -17.885 -85.575 -14.72 -85.475 ;
      RECT -17.885 -79.255 -14.72 -79.155 ;
      RECT -17.885 -72.655 -14.72 -72.555 ;
      RECT -17.885 -66.335 -14.72 -66.235 ;
      RECT -17.885 -59.735 -14.72 -59.635 ;
      RECT -17.885 -53.415 -14.72 -53.315 ;
      RECT -17.885 -46.815 -14.72 -46.715 ;
      RECT -17.885 -40.495 -14.72 -40.395 ;
      RECT -17.885 -33.895 -14.72 -33.795 ;
      RECT -17.885 -27.575 -14.72 -27.475 ;
      RECT -17.885 -20.975 -14.72 -20.875 ;
      RECT -17.885 -14.655 -14.72 -14.555 ;
      RECT -17.885 -8.055 -14.72 -7.955 ;
      RECT -17.885 -1.735 -14.72 -1.635 ;
      RECT -15.245 -101.195 -15.145 -100.595 ;
      RECT -15.245 -96.255 -15.145 -95.835 ;
      RECT -15.245 -94.735 -15.145 -94.315 ;
      RECT -15.245 -89.975 -15.145 -89.375 ;
      RECT -15.245 -88.275 -15.145 -87.675 ;
      RECT -15.245 -83.335 -15.145 -82.915 ;
      RECT -15.245 -81.815 -15.145 -81.395 ;
      RECT -15.245 -77.055 -15.145 -76.455 ;
      RECT -15.245 -75.355 -15.145 -74.755 ;
      RECT -15.245 -70.415 -15.145 -69.995 ;
      RECT -15.245 -68.895 -15.145 -68.475 ;
      RECT -15.245 -64.135 -15.145 -63.535 ;
      RECT -15.245 -62.435 -15.145 -61.835 ;
      RECT -15.245 -57.495 -15.145 -57.075 ;
      RECT -15.245 -55.975 -15.145 -55.555 ;
      RECT -15.245 -51.215 -15.145 -50.615 ;
      RECT -15.245 -49.515 -15.145 -48.915 ;
      RECT -15.245 -44.575 -15.145 -44.155 ;
      RECT -15.245 -43.055 -15.145 -42.635 ;
      RECT -15.245 -38.295 -15.145 -37.695 ;
      RECT -15.245 -36.595 -15.145 -35.995 ;
      RECT -15.245 -31.655 -15.145 -31.235 ;
      RECT -15.245 -30.135 -15.145 -29.715 ;
      RECT -15.245 -25.375 -15.145 -24.775 ;
      RECT -15.245 -23.675 -15.145 -23.075 ;
      RECT -15.245 -18.735 -15.145 -18.315 ;
      RECT -15.245 -17.215 -15.145 -16.795 ;
      RECT -15.245 -12.455 -15.145 -11.855 ;
      RECT -15.245 -10.755 -15.145 -10.155 ;
      RECT -15.245 -5.815 -15.145 -5.395 ;
      RECT -15.245 -4.295 -15.145 -3.875 ;
      RECT -15.245 0.465 -15.145 1.065 ;
      RECT -15.765 -96.435 -15.665 -95.835 ;
      RECT -15.765 -94.735 -15.665 -94.135 ;
      RECT -15.765 -83.515 -15.665 -82.915 ;
      RECT -15.765 -81.815 -15.665 -81.215 ;
      RECT -15.765 -70.595 -15.665 -69.995 ;
      RECT -15.765 -68.895 -15.665 -68.295 ;
      RECT -15.765 -57.675 -15.665 -57.075 ;
      RECT -15.765 -55.975 -15.665 -55.375 ;
      RECT -15.765 -44.755 -15.665 -44.155 ;
      RECT -15.765 -43.055 -15.665 -42.455 ;
      RECT -15.765 -31.835 -15.665 -31.235 ;
      RECT -15.765 -30.135 -15.665 -29.535 ;
      RECT -15.765 -18.915 -15.665 -18.315 ;
      RECT -15.765 -17.215 -15.665 -16.615 ;
      RECT -15.765 -5.995 -15.665 -5.395 ;
      RECT -15.765 -4.295 -15.665 -3.695 ;
      RECT -16.025 -96.435 -15.925 -95.835 ;
      RECT -16.025 -94.735 -15.925 -94.135 ;
      RECT -16.025 -83.515 -15.925 -82.915 ;
      RECT -16.025 -81.815 -15.925 -81.215 ;
      RECT -16.025 -70.595 -15.925 -69.995 ;
      RECT -16.025 -68.895 -15.925 -68.295 ;
      RECT -16.025 -57.675 -15.925 -57.075 ;
      RECT -16.025 -55.975 -15.925 -55.375 ;
      RECT -16.025 -44.755 -15.925 -44.155 ;
      RECT -16.025 -43.055 -15.925 -42.455 ;
      RECT -16.025 -31.835 -15.925 -31.235 ;
      RECT -16.025 -30.135 -15.925 -29.535 ;
      RECT -16.025 -18.915 -15.925 -18.315 ;
      RECT -16.025 -17.215 -15.925 -16.615 ;
      RECT -16.025 -5.995 -15.925 -5.395 ;
      RECT -16.025 -4.295 -15.925 -3.695 ;
      RECT -16.545 -101.195 -16.445 -100.595 ;
      RECT -16.545 -96.255 -16.445 -95.835 ;
      RECT -16.545 -94.735 -16.445 -94.315 ;
      RECT -16.545 -89.975 -16.445 -89.375 ;
      RECT -16.545 -88.275 -16.445 -87.675 ;
      RECT -16.545 -83.335 -16.445 -82.915 ;
      RECT -16.545 -81.815 -16.445 -81.395 ;
      RECT -16.545 -77.055 -16.445 -76.455 ;
      RECT -16.545 -75.355 -16.445 -74.755 ;
      RECT -16.545 -70.415 -16.445 -69.995 ;
      RECT -16.545 -68.895 -16.445 -68.475 ;
      RECT -16.545 -64.135 -16.445 -63.535 ;
      RECT -16.545 -62.435 -16.445 -61.835 ;
      RECT -16.545 -57.495 -16.445 -57.075 ;
      RECT -16.545 -55.975 -16.445 -55.555 ;
      RECT -16.545 -51.215 -16.445 -50.615 ;
      RECT -16.545 -49.515 -16.445 -48.915 ;
      RECT -16.545 -44.575 -16.445 -44.155 ;
      RECT -16.545 -43.055 -16.445 -42.635 ;
      RECT -16.545 -38.295 -16.445 -37.695 ;
      RECT -16.545 -36.595 -16.445 -35.995 ;
      RECT -16.545 -31.655 -16.445 -31.235 ;
      RECT -16.545 -30.135 -16.445 -29.715 ;
      RECT -16.545 -25.375 -16.445 -24.775 ;
      RECT -16.545 -23.675 -16.445 -23.075 ;
      RECT -16.545 -18.735 -16.445 -18.315 ;
      RECT -16.545 -17.215 -16.445 -16.795 ;
      RECT -16.545 -12.455 -16.445 -11.855 ;
      RECT -16.545 -10.755 -16.445 -10.155 ;
      RECT -16.545 -5.815 -16.445 -5.395 ;
      RECT -16.545 -4.295 -16.445 -3.875 ;
      RECT -16.545 0.465 -16.445 1.065 ;
      RECT -17.065 -96.435 -16.965 -95.835 ;
      RECT -17.065 -94.735 -16.965 -94.135 ;
      RECT -17.065 -83.515 -16.965 -82.915 ;
      RECT -17.065 -81.815 -16.965 -81.215 ;
      RECT -17.065 -70.595 -16.965 -69.995 ;
      RECT -17.065 -68.895 -16.965 -68.295 ;
      RECT -17.065 -57.675 -16.965 -57.075 ;
      RECT -17.065 -55.975 -16.965 -55.375 ;
      RECT -17.065 -44.755 -16.965 -44.155 ;
      RECT -17.065 -43.055 -16.965 -42.455 ;
      RECT -17.065 -31.835 -16.965 -31.235 ;
      RECT -17.065 -30.135 -16.965 -29.535 ;
      RECT -17.065 -18.915 -16.965 -18.315 ;
      RECT -17.065 -17.215 -16.965 -16.615 ;
      RECT -17.065 -5.995 -16.965 -5.395 ;
      RECT -17.065 -4.295 -16.965 -3.695 ;
      RECT -17.325 -96.435 -17.225 -95.835 ;
      RECT -17.325 -94.735 -17.225 -94.135 ;
      RECT -17.325 -83.515 -17.225 -82.915 ;
      RECT -17.325 -81.815 -17.225 -81.215 ;
      RECT -17.325 -70.595 -17.225 -69.995 ;
      RECT -17.325 -68.895 -17.225 -68.295 ;
      RECT -17.325 -57.675 -17.225 -57.075 ;
      RECT -17.325 -55.975 -17.225 -55.375 ;
      RECT -17.325 -44.755 -17.225 -44.155 ;
      RECT -17.325 -43.055 -17.225 -42.455 ;
      RECT -17.325 -31.835 -17.225 -31.235 ;
      RECT -17.325 -30.135 -17.225 -29.535 ;
      RECT -17.325 -18.915 -17.225 -18.315 ;
      RECT -17.325 -17.215 -17.225 -16.615 ;
      RECT -17.325 -5.995 -17.225 -5.395 ;
      RECT -17.325 -4.295 -17.225 -3.695 ;
      RECT -17.845 -101.195 -17.745 -100.595 ;
      RECT -17.845 -96.255 -17.745 -95.835 ;
      RECT -17.845 -94.735 -17.745 -94.315 ;
      RECT -17.845 -89.975 -17.745 -89.375 ;
      RECT -17.845 -88.275 -17.745 -87.675 ;
      RECT -17.845 -83.335 -17.745 -82.915 ;
      RECT -17.845 -81.815 -17.745 -81.395 ;
      RECT -17.845 -77.055 -17.745 -76.455 ;
      RECT -17.845 -75.355 -17.745 -74.755 ;
      RECT -17.845 -70.415 -17.745 -69.995 ;
      RECT -17.845 -68.895 -17.745 -68.475 ;
      RECT -17.845 -64.135 -17.745 -63.535 ;
      RECT -17.845 -62.435 -17.745 -61.835 ;
      RECT -17.845 -57.495 -17.745 -57.075 ;
      RECT -17.845 -55.975 -17.745 -55.555 ;
      RECT -17.845 -51.215 -17.745 -50.615 ;
      RECT -17.845 -49.515 -17.745 -48.915 ;
      RECT -17.845 -44.575 -17.745 -44.155 ;
      RECT -17.845 -43.055 -17.745 -42.635 ;
      RECT -17.845 -38.295 -17.745 -37.695 ;
      RECT -17.845 -36.595 -17.745 -35.995 ;
      RECT -17.845 -31.655 -17.745 -31.235 ;
      RECT -17.845 -30.135 -17.745 -29.715 ;
      RECT -17.845 -25.375 -17.745 -24.775 ;
      RECT -17.845 -23.675 -17.745 -23.075 ;
      RECT -17.845 -18.735 -17.745 -18.315 ;
      RECT -17.845 -17.215 -17.745 -16.795 ;
      RECT -17.845 -12.455 -17.745 -11.855 ;
      RECT -17.845 -10.755 -17.745 -10.155 ;
      RECT -17.845 -5.815 -17.745 -5.395 ;
      RECT -17.845 -4.295 -17.745 -3.875 ;
      RECT -17.845 0.465 -17.745 1.065 ;
      RECT -18.365 -96.435 -18.265 -95.835 ;
      RECT -18.365 -94.735 -18.265 -94.135 ;
      RECT -18.365 -83.515 -18.265 -82.915 ;
      RECT -18.365 -81.815 -18.265 -81.215 ;
      RECT -18.365 -70.595 -18.265 -69.995 ;
      RECT -18.365 -68.895 -18.265 -68.295 ;
      RECT -18.365 -57.675 -18.265 -57.075 ;
      RECT -18.365 -55.975 -18.265 -55.375 ;
      RECT -18.365 -44.755 -18.265 -44.155 ;
      RECT -18.365 -43.055 -18.265 -42.455 ;
      RECT -18.365 -31.835 -18.265 -31.235 ;
      RECT -18.365 -30.135 -18.265 -29.535 ;
      RECT -18.365 -18.915 -18.265 -18.315 ;
      RECT -18.365 -17.215 -18.265 -16.615 ;
      RECT -18.365 -5.995 -18.265 -5.395 ;
      RECT -18.365 -4.295 -18.265 -3.695 ;
      RECT -18.625 -96.435 -18.525 -95.835 ;
      RECT -18.625 -94.735 -18.525 -94.135 ;
      RECT -18.625 -83.515 -18.525 -82.915 ;
      RECT -18.625 -81.815 -18.525 -81.215 ;
      RECT -18.625 -70.595 -18.525 -69.995 ;
      RECT -18.625 -68.895 -18.525 -68.295 ;
      RECT -18.625 -57.675 -18.525 -57.075 ;
      RECT -18.625 -55.975 -18.525 -55.375 ;
      RECT -18.625 -44.755 -18.525 -44.155 ;
      RECT -18.625 -43.055 -18.525 -42.455 ;
      RECT -18.625 -31.835 -18.525 -31.235 ;
      RECT -18.625 -30.135 -18.525 -29.535 ;
      RECT -18.625 -18.915 -18.525 -18.315 ;
      RECT -18.625 -17.215 -18.525 -16.615 ;
      RECT -18.625 -5.995 -18.525 -5.395 ;
      RECT -18.625 -4.295 -18.525 -3.695 ;
      RECT -35.845 -100.255 -18.62 -100.155 ;
      RECT -35.845 -90.415 -18.62 -90.315 ;
      RECT -35.845 -87.335 -18.62 -87.235 ;
      RECT -35.845 -77.495 -18.62 -77.395 ;
      RECT -35.845 -74.415 -18.62 -74.315 ;
      RECT -35.845 -64.575 -18.62 -64.475 ;
      RECT -35.845 -61.495 -18.62 -61.395 ;
      RECT -35.845 -51.655 -18.62 -51.555 ;
      RECT -35.845 -48.575 -18.62 -48.475 ;
      RECT -35.845 -38.735 -18.62 -38.635 ;
      RECT -35.845 -35.655 -18.62 -35.555 ;
      RECT -35.845 -25.815 -18.62 -25.715 ;
      RECT -35.845 -22.735 -18.62 -22.635 ;
      RECT -35.845 -12.895 -18.62 -12.795 ;
      RECT -35.845 -9.815 -18.62 -9.715 ;
      RECT -35.845 0.025 -18.62 0.125 ;
      RECT -19.145 -101.195 -19.045 -100.595 ;
      RECT -19.145 -96.255 -19.045 -95.835 ;
      RECT -19.145 -94.735 -19.045 -94.315 ;
      RECT -19.145 -89.975 -19.045 -89.375 ;
      RECT -19.145 -88.275 -19.045 -87.675 ;
      RECT -19.145 -83.335 -19.045 -82.915 ;
      RECT -19.145 -81.815 -19.045 -81.395 ;
      RECT -19.145 -77.055 -19.045 -76.455 ;
      RECT -19.145 -75.355 -19.045 -74.755 ;
      RECT -19.145 -70.415 -19.045 -69.995 ;
      RECT -19.145 -68.895 -19.045 -68.475 ;
      RECT -19.145 -64.135 -19.045 -63.535 ;
      RECT -19.145 -62.435 -19.045 -61.835 ;
      RECT -19.145 -57.495 -19.045 -57.075 ;
      RECT -19.145 -55.975 -19.045 -55.555 ;
      RECT -19.145 -51.215 -19.045 -50.615 ;
      RECT -19.145 -49.515 -19.045 -48.915 ;
      RECT -19.145 -44.575 -19.045 -44.155 ;
      RECT -19.145 -43.055 -19.045 -42.635 ;
      RECT -19.145 -38.295 -19.045 -37.695 ;
      RECT -19.145 -36.595 -19.045 -35.995 ;
      RECT -19.145 -31.655 -19.045 -31.235 ;
      RECT -19.145 -30.135 -19.045 -29.715 ;
      RECT -19.145 -25.375 -19.045 -24.775 ;
      RECT -19.145 -23.675 -19.045 -23.075 ;
      RECT -19.145 -18.735 -19.045 -18.315 ;
      RECT -19.145 -17.215 -19.045 -16.795 ;
      RECT -19.145 -12.455 -19.045 -11.855 ;
      RECT -19.145 -10.755 -19.045 -10.155 ;
      RECT -19.145 -5.815 -19.045 -5.395 ;
      RECT -19.145 -4.295 -19.045 -3.875 ;
      RECT -19.145 0.465 -19.045 1.065 ;
      RECT -19.665 -96.435 -19.565 -95.835 ;
      RECT -19.665 -94.735 -19.565 -94.135 ;
      RECT -19.665 -83.515 -19.565 -82.915 ;
      RECT -19.665 -81.815 -19.565 -81.215 ;
      RECT -19.665 -70.595 -19.565 -69.995 ;
      RECT -19.665 -68.895 -19.565 -68.295 ;
      RECT -19.665 -57.675 -19.565 -57.075 ;
      RECT -19.665 -55.975 -19.565 -55.375 ;
      RECT -19.665 -44.755 -19.565 -44.155 ;
      RECT -19.665 -43.055 -19.565 -42.455 ;
      RECT -19.665 -31.835 -19.565 -31.235 ;
      RECT -19.665 -30.135 -19.565 -29.535 ;
      RECT -19.665 -18.915 -19.565 -18.315 ;
      RECT -19.665 -17.215 -19.565 -16.615 ;
      RECT -19.665 -5.995 -19.565 -5.395 ;
      RECT -19.665 -4.295 -19.565 -3.695 ;
      RECT -20.485 -98.495 -19.66 -98.395 ;
      RECT -20.485 -92.175 -19.66 -92.075 ;
      RECT -20.485 -85.575 -19.66 -85.475 ;
      RECT -20.485 -79.255 -19.66 -79.155 ;
      RECT -20.485 -72.655 -19.66 -72.555 ;
      RECT -20.485 -66.335 -19.66 -66.235 ;
      RECT -20.485 -59.735 -19.66 -59.635 ;
      RECT -20.485 -53.415 -19.66 -53.315 ;
      RECT -20.485 -46.815 -19.66 -46.715 ;
      RECT -20.485 -40.495 -19.66 -40.395 ;
      RECT -20.485 -33.895 -19.66 -33.795 ;
      RECT -20.485 -27.575 -19.66 -27.475 ;
      RECT -20.485 -20.975 -19.66 -20.875 ;
      RECT -20.485 -14.655 -19.66 -14.555 ;
      RECT -20.485 -8.055 -19.66 -7.955 ;
      RECT -20.485 -1.735 -19.66 -1.635 ;
      RECT -19.925 -96.435 -19.825 -95.835 ;
      RECT -19.925 -94.735 -19.825 -94.135 ;
      RECT -19.925 -83.515 -19.825 -82.915 ;
      RECT -19.925 -81.815 -19.825 -81.215 ;
      RECT -19.925 -70.595 -19.825 -69.995 ;
      RECT -19.925 -68.895 -19.825 -68.295 ;
      RECT -19.925 -57.675 -19.825 -57.075 ;
      RECT -19.925 -55.975 -19.825 -55.375 ;
      RECT -19.925 -44.755 -19.825 -44.155 ;
      RECT -19.925 -43.055 -19.825 -42.455 ;
      RECT -19.925 -31.835 -19.825 -31.235 ;
      RECT -19.925 -30.135 -19.825 -29.535 ;
      RECT -19.925 -18.915 -19.825 -18.315 ;
      RECT -19.925 -17.215 -19.825 -16.615 ;
      RECT -19.925 -5.995 -19.825 -5.395 ;
      RECT -19.925 -4.295 -19.825 -3.695 ;
      RECT -21.785 -98.055 -19.92 -97.955 ;
      RECT -21.785 -92.615 -19.92 -92.515 ;
      RECT -21.785 -85.135 -19.92 -85.035 ;
      RECT -21.785 -79.695 -19.92 -79.595 ;
      RECT -21.785 -72.215 -19.92 -72.115 ;
      RECT -21.785 -66.775 -19.92 -66.675 ;
      RECT -21.785 -59.295 -19.92 -59.195 ;
      RECT -21.785 -53.855 -19.92 -53.755 ;
      RECT -21.785 -46.375 -19.92 -46.275 ;
      RECT -21.785 -40.935 -19.92 -40.835 ;
      RECT -21.785 -33.455 -19.92 -33.355 ;
      RECT -21.785 -28.015 -19.92 -27.915 ;
      RECT -21.785 -20.535 -19.92 -20.435 ;
      RECT -21.785 -15.095 -19.92 -14.995 ;
      RECT -21.785 -7.615 -19.92 -7.515 ;
      RECT -21.785 -2.175 -19.92 -2.075 ;
      RECT -20.445 -101.195 -20.345 -100.595 ;
      RECT -20.445 -96.255 -20.345 -95.835 ;
      RECT -20.445 -94.735 -20.345 -94.315 ;
      RECT -20.445 -89.975 -20.345 -89.375 ;
      RECT -20.445 -88.275 -20.345 -87.675 ;
      RECT -20.445 -83.335 -20.345 -82.915 ;
      RECT -20.445 -81.815 -20.345 -81.395 ;
      RECT -20.445 -77.055 -20.345 -76.455 ;
      RECT -20.445 -75.355 -20.345 -74.755 ;
      RECT -20.445 -70.415 -20.345 -69.995 ;
      RECT -20.445 -68.895 -20.345 -68.475 ;
      RECT -20.445 -64.135 -20.345 -63.535 ;
      RECT -20.445 -62.435 -20.345 -61.835 ;
      RECT -20.445 -57.495 -20.345 -57.075 ;
      RECT -20.445 -55.975 -20.345 -55.555 ;
      RECT -20.445 -51.215 -20.345 -50.615 ;
      RECT -20.445 -49.515 -20.345 -48.915 ;
      RECT -20.445 -44.575 -20.345 -44.155 ;
      RECT -20.445 -43.055 -20.345 -42.635 ;
      RECT -20.445 -38.295 -20.345 -37.695 ;
      RECT -20.445 -36.595 -20.345 -35.995 ;
      RECT -20.445 -31.655 -20.345 -31.235 ;
      RECT -20.445 -30.135 -20.345 -29.715 ;
      RECT -20.445 -25.375 -20.345 -24.775 ;
      RECT -20.445 -23.675 -20.345 -23.075 ;
      RECT -20.445 -18.735 -20.345 -18.315 ;
      RECT -20.445 -17.215 -20.345 -16.795 ;
      RECT -20.445 -12.455 -20.345 -11.855 ;
      RECT -20.445 -10.755 -20.345 -10.155 ;
      RECT -20.445 -5.815 -20.345 -5.395 ;
      RECT -20.445 -4.295 -20.345 -3.875 ;
      RECT -20.445 0.465 -20.345 1.065 ;
      RECT -20.965 -96.435 -20.865 -95.835 ;
      RECT -20.965 -94.735 -20.865 -94.135 ;
      RECT -20.965 -83.515 -20.865 -82.915 ;
      RECT -20.965 -81.815 -20.865 -81.215 ;
      RECT -20.965 -70.595 -20.865 -69.995 ;
      RECT -20.965 -68.895 -20.865 -68.295 ;
      RECT -20.965 -57.675 -20.865 -57.075 ;
      RECT -20.965 -55.975 -20.865 -55.375 ;
      RECT -20.965 -44.755 -20.865 -44.155 ;
      RECT -20.965 -43.055 -20.865 -42.455 ;
      RECT -20.965 -31.835 -20.865 -31.235 ;
      RECT -20.965 -30.135 -20.865 -29.535 ;
      RECT -20.965 -18.915 -20.865 -18.315 ;
      RECT -20.965 -17.215 -20.865 -16.615 ;
      RECT -20.965 -5.995 -20.865 -5.395 ;
      RECT -20.965 -4.295 -20.865 -3.695 ;
      RECT -23.085 -98.275 -20.96 -98.175 ;
      RECT -23.085 -92.395 -20.96 -92.295 ;
      RECT -23.085 -85.355 -20.96 -85.255 ;
      RECT -23.085 -79.475 -20.96 -79.375 ;
      RECT -23.085 -72.435 -20.96 -72.335 ;
      RECT -23.085 -66.555 -20.96 -66.455 ;
      RECT -23.085 -59.515 -20.96 -59.415 ;
      RECT -23.085 -53.635 -20.96 -53.535 ;
      RECT -23.085 -46.595 -20.96 -46.495 ;
      RECT -23.085 -40.715 -20.96 -40.615 ;
      RECT -23.085 -33.675 -20.96 -33.575 ;
      RECT -23.085 -27.795 -20.96 -27.695 ;
      RECT -23.085 -20.755 -20.96 -20.655 ;
      RECT -23.085 -14.875 -20.96 -14.775 ;
      RECT -23.085 -7.835 -20.96 -7.735 ;
      RECT -23.085 -1.955 -20.96 -1.855 ;
      RECT -21.225 -96.435 -21.125 -95.835 ;
      RECT -21.225 -94.735 -21.125 -94.135 ;
      RECT -21.225 -83.515 -21.125 -82.915 ;
      RECT -21.225 -81.815 -21.125 -81.215 ;
      RECT -21.225 -70.595 -21.125 -69.995 ;
      RECT -21.225 -68.895 -21.125 -68.295 ;
      RECT -21.225 -57.675 -21.125 -57.075 ;
      RECT -21.225 -55.975 -21.125 -55.375 ;
      RECT -21.225 -44.755 -21.125 -44.155 ;
      RECT -21.225 -43.055 -21.125 -42.455 ;
      RECT -21.225 -31.835 -21.125 -31.235 ;
      RECT -21.225 -30.135 -21.125 -29.535 ;
      RECT -21.225 -18.915 -21.125 -18.315 ;
      RECT -21.225 -17.215 -21.125 -16.615 ;
      RECT -21.225 -5.995 -21.125 -5.395 ;
      RECT -21.225 -4.295 -21.125 -3.695 ;
      RECT -24.385 -98.495 -21.22 -98.395 ;
      RECT -24.385 -92.175 -21.22 -92.075 ;
      RECT -24.385 -85.575 -21.22 -85.475 ;
      RECT -24.385 -79.255 -21.22 -79.155 ;
      RECT -24.385 -72.655 -21.22 -72.555 ;
      RECT -24.385 -66.335 -21.22 -66.235 ;
      RECT -24.385 -59.735 -21.22 -59.635 ;
      RECT -24.385 -53.415 -21.22 -53.315 ;
      RECT -24.385 -46.815 -21.22 -46.715 ;
      RECT -24.385 -40.495 -21.22 -40.395 ;
      RECT -24.385 -33.895 -21.22 -33.795 ;
      RECT -24.385 -27.575 -21.22 -27.475 ;
      RECT -24.385 -20.975 -21.22 -20.875 ;
      RECT -24.385 -14.655 -21.22 -14.555 ;
      RECT -24.385 -8.055 -21.22 -7.955 ;
      RECT -24.385 -1.735 -21.22 -1.635 ;
      RECT -21.745 -101.195 -21.645 -100.595 ;
      RECT -21.745 -96.255 -21.645 -95.835 ;
      RECT -21.745 -94.735 -21.645 -94.315 ;
      RECT -21.745 -89.975 -21.645 -89.375 ;
      RECT -21.745 -88.275 -21.645 -87.675 ;
      RECT -21.745 -83.335 -21.645 -82.915 ;
      RECT -21.745 -81.815 -21.645 -81.395 ;
      RECT -21.745 -77.055 -21.645 -76.455 ;
      RECT -21.745 -75.355 -21.645 -74.755 ;
      RECT -21.745 -70.415 -21.645 -69.995 ;
      RECT -21.745 -68.895 -21.645 -68.475 ;
      RECT -21.745 -64.135 -21.645 -63.535 ;
      RECT -21.745 -62.435 -21.645 -61.835 ;
      RECT -21.745 -57.495 -21.645 -57.075 ;
      RECT -21.745 -55.975 -21.645 -55.555 ;
      RECT -21.745 -51.215 -21.645 -50.615 ;
      RECT -21.745 -49.515 -21.645 -48.915 ;
      RECT -21.745 -44.575 -21.645 -44.155 ;
      RECT -21.745 -43.055 -21.645 -42.635 ;
      RECT -21.745 -38.295 -21.645 -37.695 ;
      RECT -21.745 -36.595 -21.645 -35.995 ;
      RECT -21.745 -31.655 -21.645 -31.235 ;
      RECT -21.745 -30.135 -21.645 -29.715 ;
      RECT -21.745 -25.375 -21.645 -24.775 ;
      RECT -21.745 -23.675 -21.645 -23.075 ;
      RECT -21.745 -18.735 -21.645 -18.315 ;
      RECT -21.745 -17.215 -21.645 -16.795 ;
      RECT -21.745 -12.455 -21.645 -11.855 ;
      RECT -21.745 -10.755 -21.645 -10.155 ;
      RECT -21.745 -5.815 -21.645 -5.395 ;
      RECT -21.745 -4.295 -21.645 -3.875 ;
      RECT -21.745 0.465 -21.645 1.065 ;
      RECT -22.265 -96.435 -22.165 -95.835 ;
      RECT -22.265 -94.735 -22.165 -94.135 ;
      RECT -22.265 -83.515 -22.165 -82.915 ;
      RECT -22.265 -81.815 -22.165 -81.215 ;
      RECT -22.265 -70.595 -22.165 -69.995 ;
      RECT -22.265 -68.895 -22.165 -68.295 ;
      RECT -22.265 -57.675 -22.165 -57.075 ;
      RECT -22.265 -55.975 -22.165 -55.375 ;
      RECT -22.265 -44.755 -22.165 -44.155 ;
      RECT -22.265 -43.055 -22.165 -42.455 ;
      RECT -22.265 -31.835 -22.165 -31.235 ;
      RECT -22.265 -30.135 -22.165 -29.535 ;
      RECT -22.265 -18.915 -22.165 -18.315 ;
      RECT -22.265 -17.215 -22.165 -16.615 ;
      RECT -22.265 -5.995 -22.165 -5.395 ;
      RECT -22.265 -4.295 -22.165 -3.695 ;
      RECT -22.525 -96.435 -22.425 -95.835 ;
      RECT -22.525 -94.735 -22.425 -94.135 ;
      RECT -22.525 -83.515 -22.425 -82.915 ;
      RECT -22.525 -81.815 -22.425 -81.215 ;
      RECT -22.525 -70.595 -22.425 -69.995 ;
      RECT -22.525 -68.895 -22.425 -68.295 ;
      RECT -22.525 -57.675 -22.425 -57.075 ;
      RECT -22.525 -55.975 -22.425 -55.375 ;
      RECT -22.525 -44.755 -22.425 -44.155 ;
      RECT -22.525 -43.055 -22.425 -42.455 ;
      RECT -22.525 -31.835 -22.425 -31.235 ;
      RECT -22.525 -30.135 -22.425 -29.535 ;
      RECT -22.525 -18.915 -22.425 -18.315 ;
      RECT -22.525 -17.215 -22.425 -16.615 ;
      RECT -22.525 -5.995 -22.425 -5.395 ;
      RECT -22.525 -4.295 -22.425 -3.695 ;
      RECT -23.045 -101.195 -22.945 -100.595 ;
      RECT -23.045 -96.255 -22.945 -95.835 ;
      RECT -23.045 -94.735 -22.945 -94.315 ;
      RECT -23.045 -89.975 -22.945 -89.375 ;
      RECT -23.045 -88.275 -22.945 -87.675 ;
      RECT -23.045 -83.335 -22.945 -82.915 ;
      RECT -23.045 -81.815 -22.945 -81.395 ;
      RECT -23.045 -77.055 -22.945 -76.455 ;
      RECT -23.045 -75.355 -22.945 -74.755 ;
      RECT -23.045 -70.415 -22.945 -69.995 ;
      RECT -23.045 -68.895 -22.945 -68.475 ;
      RECT -23.045 -64.135 -22.945 -63.535 ;
      RECT -23.045 -62.435 -22.945 -61.835 ;
      RECT -23.045 -57.495 -22.945 -57.075 ;
      RECT -23.045 -55.975 -22.945 -55.555 ;
      RECT -23.045 -51.215 -22.945 -50.615 ;
      RECT -23.045 -49.515 -22.945 -48.915 ;
      RECT -23.045 -44.575 -22.945 -44.155 ;
      RECT -23.045 -43.055 -22.945 -42.635 ;
      RECT -23.045 -38.295 -22.945 -37.695 ;
      RECT -23.045 -36.595 -22.945 -35.995 ;
      RECT -23.045 -31.655 -22.945 -31.235 ;
      RECT -23.045 -30.135 -22.945 -29.715 ;
      RECT -23.045 -25.375 -22.945 -24.775 ;
      RECT -23.045 -23.675 -22.945 -23.075 ;
      RECT -23.045 -18.735 -22.945 -18.315 ;
      RECT -23.045 -17.215 -22.945 -16.795 ;
      RECT -23.045 -12.455 -22.945 -11.855 ;
      RECT -23.045 -10.755 -22.945 -10.155 ;
      RECT -23.045 -5.815 -22.945 -5.395 ;
      RECT -23.045 -4.295 -22.945 -3.875 ;
      RECT -23.045 0.465 -22.945 1.065 ;
      RECT -23.565 -96.435 -23.465 -95.835 ;
      RECT -23.565 -94.735 -23.465 -94.135 ;
      RECT -23.565 -83.515 -23.465 -82.915 ;
      RECT -23.565 -81.815 -23.465 -81.215 ;
      RECT -23.565 -70.595 -23.465 -69.995 ;
      RECT -23.565 -68.895 -23.465 -68.295 ;
      RECT -23.565 -57.675 -23.465 -57.075 ;
      RECT -23.565 -55.975 -23.465 -55.375 ;
      RECT -23.565 -44.755 -23.465 -44.155 ;
      RECT -23.565 -43.055 -23.465 -42.455 ;
      RECT -23.565 -31.835 -23.465 -31.235 ;
      RECT -23.565 -30.135 -23.465 -29.535 ;
      RECT -23.565 -18.915 -23.465 -18.315 ;
      RECT -23.565 -17.215 -23.465 -16.615 ;
      RECT -23.565 -5.995 -23.465 -5.395 ;
      RECT -23.565 -4.295 -23.465 -3.695 ;
      RECT -23.825 -96.435 -23.725 -95.835 ;
      RECT -23.825 -94.735 -23.725 -94.135 ;
      RECT -23.825 -83.515 -23.725 -82.915 ;
      RECT -23.825 -81.815 -23.725 -81.215 ;
      RECT -23.825 -70.595 -23.725 -69.995 ;
      RECT -23.825 -68.895 -23.725 -68.295 ;
      RECT -23.825 -57.675 -23.725 -57.075 ;
      RECT -23.825 -55.975 -23.725 -55.375 ;
      RECT -23.825 -44.755 -23.725 -44.155 ;
      RECT -23.825 -43.055 -23.725 -42.455 ;
      RECT -23.825 -31.835 -23.725 -31.235 ;
      RECT -23.825 -30.135 -23.725 -29.535 ;
      RECT -23.825 -18.915 -23.725 -18.315 ;
      RECT -23.825 -17.215 -23.725 -16.615 ;
      RECT -23.825 -5.995 -23.725 -5.395 ;
      RECT -23.825 -4.295 -23.725 -3.695 ;
      RECT -24.345 -101.195 -24.245 -100.595 ;
      RECT -24.345 -96.255 -24.245 -95.835 ;
      RECT -24.345 -94.735 -24.245 -94.315 ;
      RECT -24.345 -89.975 -24.245 -89.375 ;
      RECT -24.345 -88.275 -24.245 -87.675 ;
      RECT -24.345 -83.335 -24.245 -82.915 ;
      RECT -24.345 -81.815 -24.245 -81.395 ;
      RECT -24.345 -77.055 -24.245 -76.455 ;
      RECT -24.345 -75.355 -24.245 -74.755 ;
      RECT -24.345 -70.415 -24.245 -69.995 ;
      RECT -24.345 -68.895 -24.245 -68.475 ;
      RECT -24.345 -64.135 -24.245 -63.535 ;
      RECT -24.345 -62.435 -24.245 -61.835 ;
      RECT -24.345 -57.495 -24.245 -57.075 ;
      RECT -24.345 -55.975 -24.245 -55.555 ;
      RECT -24.345 -51.215 -24.245 -50.615 ;
      RECT -24.345 -49.515 -24.245 -48.915 ;
      RECT -24.345 -44.575 -24.245 -44.155 ;
      RECT -24.345 -43.055 -24.245 -42.635 ;
      RECT -24.345 -38.295 -24.245 -37.695 ;
      RECT -24.345 -36.595 -24.245 -35.995 ;
      RECT -24.345 -31.655 -24.245 -31.235 ;
      RECT -24.345 -30.135 -24.245 -29.715 ;
      RECT -24.345 -25.375 -24.245 -24.775 ;
      RECT -24.345 -23.675 -24.245 -23.075 ;
      RECT -24.345 -18.735 -24.245 -18.315 ;
      RECT -24.345 -17.215 -24.245 -16.795 ;
      RECT -24.345 -12.455 -24.245 -11.855 ;
      RECT -24.345 -10.755 -24.245 -10.155 ;
      RECT -24.345 -5.815 -24.245 -5.395 ;
      RECT -24.345 -4.295 -24.245 -3.875 ;
      RECT -24.345 0.465 -24.245 1.065 ;
      RECT -24.865 -96.435 -24.765 -95.835 ;
      RECT -24.865 -94.735 -24.765 -94.135 ;
      RECT -24.865 -83.515 -24.765 -82.915 ;
      RECT -24.865 -81.815 -24.765 -81.215 ;
      RECT -24.865 -70.595 -24.765 -69.995 ;
      RECT -24.865 -68.895 -24.765 -68.295 ;
      RECT -24.865 -57.675 -24.765 -57.075 ;
      RECT -24.865 -55.975 -24.765 -55.375 ;
      RECT -24.865 -44.755 -24.765 -44.155 ;
      RECT -24.865 -43.055 -24.765 -42.455 ;
      RECT -24.865 -31.835 -24.765 -31.235 ;
      RECT -24.865 -30.135 -24.765 -29.535 ;
      RECT -24.865 -18.915 -24.765 -18.315 ;
      RECT -24.865 -17.215 -24.765 -16.615 ;
      RECT -24.865 -5.995 -24.765 -5.395 ;
      RECT -24.865 -4.295 -24.765 -3.695 ;
      RECT -35.845 -99.815 -24.86 -99.715 ;
      RECT -35.845 -90.855 -24.86 -90.755 ;
      RECT -35.845 -86.895 -24.86 -86.795 ;
      RECT -35.845 -77.935 -24.86 -77.835 ;
      RECT -35.845 -73.975 -24.86 -73.875 ;
      RECT -35.845 -65.015 -24.86 -64.915 ;
      RECT -35.845 -61.055 -24.86 -60.955 ;
      RECT -35.845 -52.095 -24.86 -51.995 ;
      RECT -35.845 -48.135 -24.86 -48.035 ;
      RECT -35.845 -39.175 -24.86 -39.075 ;
      RECT -35.845 -35.215 -24.86 -35.115 ;
      RECT -35.845 -26.255 -24.86 -26.155 ;
      RECT -35.845 -22.295 -24.86 -22.195 ;
      RECT -35.845 -13.335 -24.86 -13.235 ;
      RECT -35.845 -9.375 -24.86 -9.275 ;
      RECT -35.845 -0.415 -24.86 -0.315 ;
      RECT -25.125 -96.435 -25.025 -95.835 ;
      RECT -25.125 -94.735 -25.025 -94.135 ;
      RECT -25.125 -83.515 -25.025 -82.915 ;
      RECT -25.125 -81.815 -25.025 -81.215 ;
      RECT -25.125 -70.595 -25.025 -69.995 ;
      RECT -25.125 -68.895 -25.025 -68.295 ;
      RECT -25.125 -57.675 -25.025 -57.075 ;
      RECT -25.125 -55.975 -25.025 -55.375 ;
      RECT -25.125 -44.755 -25.025 -44.155 ;
      RECT -25.125 -43.055 -25.025 -42.455 ;
      RECT -25.125 -31.835 -25.025 -31.235 ;
      RECT -25.125 -30.135 -25.025 -29.535 ;
      RECT -25.125 -18.915 -25.025 -18.315 ;
      RECT -25.125 -17.215 -25.025 -16.615 ;
      RECT -25.125 -5.995 -25.025 -5.395 ;
      RECT -25.125 -4.295 -25.025 -3.695 ;
      RECT -25.645 -101.195 -25.545 -100.595 ;
      RECT -25.645 -96.255 -25.545 -95.835 ;
      RECT -25.645 -94.735 -25.545 -94.315 ;
      RECT -25.645 -89.975 -25.545 -89.375 ;
      RECT -25.645 -88.275 -25.545 -87.675 ;
      RECT -25.645 -83.335 -25.545 -82.915 ;
      RECT -25.645 -81.815 -25.545 -81.395 ;
      RECT -25.645 -77.055 -25.545 -76.455 ;
      RECT -25.645 -75.355 -25.545 -74.755 ;
      RECT -25.645 -70.415 -25.545 -69.995 ;
      RECT -25.645 -68.895 -25.545 -68.475 ;
      RECT -25.645 -64.135 -25.545 -63.535 ;
      RECT -25.645 -62.435 -25.545 -61.835 ;
      RECT -25.645 -57.495 -25.545 -57.075 ;
      RECT -25.645 -55.975 -25.545 -55.555 ;
      RECT -25.645 -51.215 -25.545 -50.615 ;
      RECT -25.645 -49.515 -25.545 -48.915 ;
      RECT -25.645 -44.575 -25.545 -44.155 ;
      RECT -25.645 -43.055 -25.545 -42.635 ;
      RECT -25.645 -38.295 -25.545 -37.695 ;
      RECT -25.645 -36.595 -25.545 -35.995 ;
      RECT -25.645 -31.655 -25.545 -31.235 ;
      RECT -25.645 -30.135 -25.545 -29.715 ;
      RECT -25.645 -25.375 -25.545 -24.775 ;
      RECT -25.645 -23.675 -25.545 -23.075 ;
      RECT -25.645 -18.735 -25.545 -18.315 ;
      RECT -25.645 -17.215 -25.545 -16.795 ;
      RECT -25.645 -12.455 -25.545 -11.855 ;
      RECT -25.645 -10.755 -25.545 -10.155 ;
      RECT -25.645 -5.815 -25.545 -5.395 ;
      RECT -25.645 -4.295 -25.545 -3.875 ;
      RECT -25.645 0.465 -25.545 1.065 ;
      RECT -26.165 -96.435 -26.065 -95.835 ;
      RECT -26.165 -94.735 -26.065 -94.135 ;
      RECT -26.165 -83.515 -26.065 -82.915 ;
      RECT -26.165 -81.815 -26.065 -81.215 ;
      RECT -26.165 -70.595 -26.065 -69.995 ;
      RECT -26.165 -68.895 -26.065 -68.295 ;
      RECT -26.165 -57.675 -26.065 -57.075 ;
      RECT -26.165 -55.975 -26.065 -55.375 ;
      RECT -26.165 -44.755 -26.065 -44.155 ;
      RECT -26.165 -43.055 -26.065 -42.455 ;
      RECT -26.165 -31.835 -26.065 -31.235 ;
      RECT -26.165 -30.135 -26.065 -29.535 ;
      RECT -26.165 -18.915 -26.065 -18.315 ;
      RECT -26.165 -17.215 -26.065 -16.615 ;
      RECT -26.165 -5.995 -26.065 -5.395 ;
      RECT -26.165 -4.295 -26.065 -3.695 ;
      RECT -26.985 -98.495 -26.16 -98.395 ;
      RECT -26.985 -92.175 -26.16 -92.075 ;
      RECT -26.985 -85.575 -26.16 -85.475 ;
      RECT -26.985 -79.255 -26.16 -79.155 ;
      RECT -26.985 -72.655 -26.16 -72.555 ;
      RECT -26.985 -66.335 -26.16 -66.235 ;
      RECT -26.985 -59.735 -26.16 -59.635 ;
      RECT -26.985 -53.415 -26.16 -53.315 ;
      RECT -26.985 -46.815 -26.16 -46.715 ;
      RECT -26.985 -40.495 -26.16 -40.395 ;
      RECT -26.985 -33.895 -26.16 -33.795 ;
      RECT -26.985 -27.575 -26.16 -27.475 ;
      RECT -26.985 -20.975 -26.16 -20.875 ;
      RECT -26.985 -14.655 -26.16 -14.555 ;
      RECT -26.985 -8.055 -26.16 -7.955 ;
      RECT -26.985 -1.735 -26.16 -1.635 ;
      RECT -26.425 -96.435 -26.325 -95.835 ;
      RECT -26.425 -94.735 -26.325 -94.135 ;
      RECT -26.425 -83.515 -26.325 -82.915 ;
      RECT -26.425 -81.815 -26.325 -81.215 ;
      RECT -26.425 -70.595 -26.325 -69.995 ;
      RECT -26.425 -68.895 -26.325 -68.295 ;
      RECT -26.425 -57.675 -26.325 -57.075 ;
      RECT -26.425 -55.975 -26.325 -55.375 ;
      RECT -26.425 -44.755 -26.325 -44.155 ;
      RECT -26.425 -43.055 -26.325 -42.455 ;
      RECT -26.425 -31.835 -26.325 -31.235 ;
      RECT -26.425 -30.135 -26.325 -29.535 ;
      RECT -26.425 -18.915 -26.325 -18.315 ;
      RECT -26.425 -17.215 -26.325 -16.615 ;
      RECT -26.425 -5.995 -26.325 -5.395 ;
      RECT -26.425 -4.295 -26.325 -3.695 ;
      RECT -28.285 -98.055 -26.42 -97.955 ;
      RECT -28.285 -92.615 -26.42 -92.515 ;
      RECT -28.285 -85.135 -26.42 -85.035 ;
      RECT -28.285 -79.695 -26.42 -79.595 ;
      RECT -28.285 -72.215 -26.42 -72.115 ;
      RECT -28.285 -66.775 -26.42 -66.675 ;
      RECT -28.285 -59.295 -26.42 -59.195 ;
      RECT -28.285 -53.855 -26.42 -53.755 ;
      RECT -28.285 -46.375 -26.42 -46.275 ;
      RECT -28.285 -40.935 -26.42 -40.835 ;
      RECT -28.285 -33.455 -26.42 -33.355 ;
      RECT -28.285 -28.015 -26.42 -27.915 ;
      RECT -28.285 -20.535 -26.42 -20.435 ;
      RECT -28.285 -15.095 -26.42 -14.995 ;
      RECT -28.285 -7.615 -26.42 -7.515 ;
      RECT -28.285 -2.175 -26.42 -2.075 ;
      RECT -26.945 -101.195 -26.845 -100.595 ;
      RECT -26.945 -96.255 -26.845 -95.835 ;
      RECT -26.945 -94.735 -26.845 -94.315 ;
      RECT -26.945 -89.975 -26.845 -89.375 ;
      RECT -26.945 -88.275 -26.845 -87.675 ;
      RECT -26.945 -83.335 -26.845 -82.915 ;
      RECT -26.945 -81.815 -26.845 -81.395 ;
      RECT -26.945 -77.055 -26.845 -76.455 ;
      RECT -26.945 -75.355 -26.845 -74.755 ;
      RECT -26.945 -70.415 -26.845 -69.995 ;
      RECT -26.945 -68.895 -26.845 -68.475 ;
      RECT -26.945 -64.135 -26.845 -63.535 ;
      RECT -26.945 -62.435 -26.845 -61.835 ;
      RECT -26.945 -57.495 -26.845 -57.075 ;
      RECT -26.945 -55.975 -26.845 -55.555 ;
      RECT -26.945 -51.215 -26.845 -50.615 ;
      RECT -26.945 -49.515 -26.845 -48.915 ;
      RECT -26.945 -44.575 -26.845 -44.155 ;
      RECT -26.945 -43.055 -26.845 -42.635 ;
      RECT -26.945 -38.295 -26.845 -37.695 ;
      RECT -26.945 -36.595 -26.845 -35.995 ;
      RECT -26.945 -31.655 -26.845 -31.235 ;
      RECT -26.945 -30.135 -26.845 -29.715 ;
      RECT -26.945 -25.375 -26.845 -24.775 ;
      RECT -26.945 -23.675 -26.845 -23.075 ;
      RECT -26.945 -18.735 -26.845 -18.315 ;
      RECT -26.945 -17.215 -26.845 -16.795 ;
      RECT -26.945 -12.455 -26.845 -11.855 ;
      RECT -26.945 -10.755 -26.845 -10.155 ;
      RECT -26.945 -5.815 -26.845 -5.395 ;
      RECT -26.945 -4.295 -26.845 -3.875 ;
      RECT -26.945 0.465 -26.845 1.065 ;
      RECT -27.465 -96.435 -27.365 -95.835 ;
      RECT -27.465 -94.735 -27.365 -94.135 ;
      RECT -27.465 -83.515 -27.365 -82.915 ;
      RECT -27.465 -81.815 -27.365 -81.215 ;
      RECT -27.465 -70.595 -27.365 -69.995 ;
      RECT -27.465 -68.895 -27.365 -68.295 ;
      RECT -27.465 -57.675 -27.365 -57.075 ;
      RECT -27.465 -55.975 -27.365 -55.375 ;
      RECT -27.465 -44.755 -27.365 -44.155 ;
      RECT -27.465 -43.055 -27.365 -42.455 ;
      RECT -27.465 -31.835 -27.365 -31.235 ;
      RECT -27.465 -30.135 -27.365 -29.535 ;
      RECT -27.465 -18.915 -27.365 -18.315 ;
      RECT -27.465 -17.215 -27.365 -16.615 ;
      RECT -27.465 -5.995 -27.365 -5.395 ;
      RECT -27.465 -4.295 -27.365 -3.695 ;
      RECT -29.585 -98.275 -27.46 -98.175 ;
      RECT -29.585 -92.395 -27.46 -92.295 ;
      RECT -29.585 -85.355 -27.46 -85.255 ;
      RECT -29.585 -79.475 -27.46 -79.375 ;
      RECT -29.585 -72.435 -27.46 -72.335 ;
      RECT -29.585 -66.555 -27.46 -66.455 ;
      RECT -29.585 -59.515 -27.46 -59.415 ;
      RECT -29.585 -53.635 -27.46 -53.535 ;
      RECT -29.585 -46.595 -27.46 -46.495 ;
      RECT -29.585 -40.715 -27.46 -40.615 ;
      RECT -29.585 -33.675 -27.46 -33.575 ;
      RECT -29.585 -27.795 -27.46 -27.695 ;
      RECT -29.585 -20.755 -27.46 -20.655 ;
      RECT -29.585 -14.875 -27.46 -14.775 ;
      RECT -29.585 -7.835 -27.46 -7.735 ;
      RECT -29.585 -1.955 -27.46 -1.855 ;
      RECT -27.725 -96.435 -27.625 -95.835 ;
      RECT -27.725 -94.735 -27.625 -94.135 ;
      RECT -27.725 -83.515 -27.625 -82.915 ;
      RECT -27.725 -81.815 -27.625 -81.215 ;
      RECT -27.725 -70.595 -27.625 -69.995 ;
      RECT -27.725 -68.895 -27.625 -68.295 ;
      RECT -27.725 -57.675 -27.625 -57.075 ;
      RECT -27.725 -55.975 -27.625 -55.375 ;
      RECT -27.725 -44.755 -27.625 -44.155 ;
      RECT -27.725 -43.055 -27.625 -42.455 ;
      RECT -27.725 -31.835 -27.625 -31.235 ;
      RECT -27.725 -30.135 -27.625 -29.535 ;
      RECT -27.725 -18.915 -27.625 -18.315 ;
      RECT -27.725 -17.215 -27.625 -16.615 ;
      RECT -27.725 -5.995 -27.625 -5.395 ;
      RECT -27.725 -4.295 -27.625 -3.695 ;
      RECT -30.885 -98.495 -27.72 -98.395 ;
      RECT -30.885 -92.175 -27.72 -92.075 ;
      RECT -30.885 -85.575 -27.72 -85.475 ;
      RECT -30.885 -79.255 -27.72 -79.155 ;
      RECT -30.885 -72.655 -27.72 -72.555 ;
      RECT -30.885 -66.335 -27.72 -66.235 ;
      RECT -30.885 -59.735 -27.72 -59.635 ;
      RECT -30.885 -53.415 -27.72 -53.315 ;
      RECT -30.885 -46.815 -27.72 -46.715 ;
      RECT -30.885 -40.495 -27.72 -40.395 ;
      RECT -30.885 -33.895 -27.72 -33.795 ;
      RECT -30.885 -27.575 -27.72 -27.475 ;
      RECT -30.885 -20.975 -27.72 -20.875 ;
      RECT -30.885 -14.655 -27.72 -14.555 ;
      RECT -30.885 -8.055 -27.72 -7.955 ;
      RECT -30.885 -1.735 -27.72 -1.635 ;
      RECT -28.245 -101.195 -28.145 -100.595 ;
      RECT -28.245 -96.255 -28.145 -95.835 ;
      RECT -28.245 -94.735 -28.145 -94.315 ;
      RECT -28.245 -89.975 -28.145 -89.375 ;
      RECT -28.245 -88.275 -28.145 -87.675 ;
      RECT -28.245 -83.335 -28.145 -82.915 ;
      RECT -28.245 -81.815 -28.145 -81.395 ;
      RECT -28.245 -77.055 -28.145 -76.455 ;
      RECT -28.245 -75.355 -28.145 -74.755 ;
      RECT -28.245 -70.415 -28.145 -69.995 ;
      RECT -28.245 -68.895 -28.145 -68.475 ;
      RECT -28.245 -64.135 -28.145 -63.535 ;
      RECT -28.245 -62.435 -28.145 -61.835 ;
      RECT -28.245 -57.495 -28.145 -57.075 ;
      RECT -28.245 -55.975 -28.145 -55.555 ;
      RECT -28.245 -51.215 -28.145 -50.615 ;
      RECT -28.245 -49.515 -28.145 -48.915 ;
      RECT -28.245 -44.575 -28.145 -44.155 ;
      RECT -28.245 -43.055 -28.145 -42.635 ;
      RECT -28.245 -38.295 -28.145 -37.695 ;
      RECT -28.245 -36.595 -28.145 -35.995 ;
      RECT -28.245 -31.655 -28.145 -31.235 ;
      RECT -28.245 -30.135 -28.145 -29.715 ;
      RECT -28.245 -25.375 -28.145 -24.775 ;
      RECT -28.245 -23.675 -28.145 -23.075 ;
      RECT -28.245 -18.735 -28.145 -18.315 ;
      RECT -28.245 -17.215 -28.145 -16.795 ;
      RECT -28.245 -12.455 -28.145 -11.855 ;
      RECT -28.245 -10.755 -28.145 -10.155 ;
      RECT -28.245 -5.815 -28.145 -5.395 ;
      RECT -28.245 -4.295 -28.145 -3.875 ;
      RECT -28.245 0.465 -28.145 1.065 ;
      RECT -28.765 -96.435 -28.665 -95.835 ;
      RECT -28.765 -94.735 -28.665 -94.135 ;
      RECT -28.765 -83.515 -28.665 -82.915 ;
      RECT -28.765 -81.815 -28.665 -81.215 ;
      RECT -28.765 -70.595 -28.665 -69.995 ;
      RECT -28.765 -68.895 -28.665 -68.295 ;
      RECT -28.765 -57.675 -28.665 -57.075 ;
      RECT -28.765 -55.975 -28.665 -55.375 ;
      RECT -28.765 -44.755 -28.665 -44.155 ;
      RECT -28.765 -43.055 -28.665 -42.455 ;
      RECT -28.765 -31.835 -28.665 -31.235 ;
      RECT -28.765 -30.135 -28.665 -29.535 ;
      RECT -28.765 -18.915 -28.665 -18.315 ;
      RECT -28.765 -17.215 -28.665 -16.615 ;
      RECT -28.765 -5.995 -28.665 -5.395 ;
      RECT -28.765 -4.295 -28.665 -3.695 ;
      RECT -29.025 -96.435 -28.925 -95.835 ;
      RECT -29.025 -94.735 -28.925 -94.135 ;
      RECT -29.025 -83.515 -28.925 -82.915 ;
      RECT -29.025 -81.815 -28.925 -81.215 ;
      RECT -29.025 -70.595 -28.925 -69.995 ;
      RECT -29.025 -68.895 -28.925 -68.295 ;
      RECT -29.025 -57.675 -28.925 -57.075 ;
      RECT -29.025 -55.975 -28.925 -55.375 ;
      RECT -29.025 -44.755 -28.925 -44.155 ;
      RECT -29.025 -43.055 -28.925 -42.455 ;
      RECT -29.025 -31.835 -28.925 -31.235 ;
      RECT -29.025 -30.135 -28.925 -29.535 ;
      RECT -29.025 -18.915 -28.925 -18.315 ;
      RECT -29.025 -17.215 -28.925 -16.615 ;
      RECT -29.025 -5.995 -28.925 -5.395 ;
      RECT -29.025 -4.295 -28.925 -3.695 ;
      RECT -29.545 -101.195 -29.445 -100.595 ;
      RECT -29.545 -96.255 -29.445 -95.835 ;
      RECT -29.545 -94.735 -29.445 -94.315 ;
      RECT -29.545 -89.975 -29.445 -89.375 ;
      RECT -29.545 -88.275 -29.445 -87.675 ;
      RECT -29.545 -83.335 -29.445 -82.915 ;
      RECT -29.545 -81.815 -29.445 -81.395 ;
      RECT -29.545 -77.055 -29.445 -76.455 ;
      RECT -29.545 -75.355 -29.445 -74.755 ;
      RECT -29.545 -70.415 -29.445 -69.995 ;
      RECT -29.545 -68.895 -29.445 -68.475 ;
      RECT -29.545 -64.135 -29.445 -63.535 ;
      RECT -29.545 -62.435 -29.445 -61.835 ;
      RECT -29.545 -57.495 -29.445 -57.075 ;
      RECT -29.545 -55.975 -29.445 -55.555 ;
      RECT -29.545 -51.215 -29.445 -50.615 ;
      RECT -29.545 -49.515 -29.445 -48.915 ;
      RECT -29.545 -44.575 -29.445 -44.155 ;
      RECT -29.545 -43.055 -29.445 -42.635 ;
      RECT -29.545 -38.295 -29.445 -37.695 ;
      RECT -29.545 -36.595 -29.445 -35.995 ;
      RECT -29.545 -31.655 -29.445 -31.235 ;
      RECT -29.545 -30.135 -29.445 -29.715 ;
      RECT -29.545 -25.375 -29.445 -24.775 ;
      RECT -29.545 -23.675 -29.445 -23.075 ;
      RECT -29.545 -18.735 -29.445 -18.315 ;
      RECT -29.545 -17.215 -29.445 -16.795 ;
      RECT -29.545 -12.455 -29.445 -11.855 ;
      RECT -29.545 -10.755 -29.445 -10.155 ;
      RECT -29.545 -5.815 -29.445 -5.395 ;
      RECT -29.545 -4.295 -29.445 -3.875 ;
      RECT -29.545 0.465 -29.445 1.065 ;
      RECT -30.065 -96.435 -29.965 -95.835 ;
      RECT -30.065 -94.735 -29.965 -94.135 ;
      RECT -30.065 -83.515 -29.965 -82.915 ;
      RECT -30.065 -81.815 -29.965 -81.215 ;
      RECT -30.065 -70.595 -29.965 -69.995 ;
      RECT -30.065 -68.895 -29.965 -68.295 ;
      RECT -30.065 -57.675 -29.965 -57.075 ;
      RECT -30.065 -55.975 -29.965 -55.375 ;
      RECT -30.065 -44.755 -29.965 -44.155 ;
      RECT -30.065 -43.055 -29.965 -42.455 ;
      RECT -30.065 -31.835 -29.965 -31.235 ;
      RECT -30.065 -30.135 -29.965 -29.535 ;
      RECT -30.065 -18.915 -29.965 -18.315 ;
      RECT -30.065 -17.215 -29.965 -16.615 ;
      RECT -30.065 -5.995 -29.965 -5.395 ;
      RECT -30.065 -4.295 -29.965 -3.695 ;
      RECT -30.325 -96.435 -30.225 -95.835 ;
      RECT -30.325 -94.735 -30.225 -94.135 ;
      RECT -30.325 -83.515 -30.225 -82.915 ;
      RECT -30.325 -81.815 -30.225 -81.215 ;
      RECT -30.325 -70.595 -30.225 -69.995 ;
      RECT -30.325 -68.895 -30.225 -68.295 ;
      RECT -30.325 -57.675 -30.225 -57.075 ;
      RECT -30.325 -55.975 -30.225 -55.375 ;
      RECT -30.325 -44.755 -30.225 -44.155 ;
      RECT -30.325 -43.055 -30.225 -42.455 ;
      RECT -30.325 -31.835 -30.225 -31.235 ;
      RECT -30.325 -30.135 -30.225 -29.535 ;
      RECT -30.325 -18.915 -30.225 -18.315 ;
      RECT -30.325 -17.215 -30.225 -16.615 ;
      RECT -30.325 -5.995 -30.225 -5.395 ;
      RECT -30.325 -4.295 -30.225 -3.695 ;
      RECT -30.845 -101.195 -30.745 -100.595 ;
      RECT -30.845 -96.255 -30.745 -95.835 ;
      RECT -30.845 -94.735 -30.745 -94.315 ;
      RECT -30.845 -89.975 -30.745 -89.375 ;
      RECT -30.845 -88.275 -30.745 -87.675 ;
      RECT -30.845 -83.335 -30.745 -82.915 ;
      RECT -30.845 -81.815 -30.745 -81.395 ;
      RECT -30.845 -77.055 -30.745 -76.455 ;
      RECT -30.845 -75.355 -30.745 -74.755 ;
      RECT -30.845 -70.415 -30.745 -69.995 ;
      RECT -30.845 -68.895 -30.745 -68.475 ;
      RECT -30.845 -64.135 -30.745 -63.535 ;
      RECT -30.845 -62.435 -30.745 -61.835 ;
      RECT -30.845 -57.495 -30.745 -57.075 ;
      RECT -30.845 -55.975 -30.745 -55.555 ;
      RECT -30.845 -51.215 -30.745 -50.615 ;
      RECT -30.845 -49.515 -30.745 -48.915 ;
      RECT -30.845 -44.575 -30.745 -44.155 ;
      RECT -30.845 -43.055 -30.745 -42.635 ;
      RECT -30.845 -38.295 -30.745 -37.695 ;
      RECT -30.845 -36.595 -30.745 -35.995 ;
      RECT -30.845 -31.655 -30.745 -31.235 ;
      RECT -30.845 -30.135 -30.745 -29.715 ;
      RECT -30.845 -25.375 -30.745 -24.775 ;
      RECT -30.845 -23.675 -30.745 -23.075 ;
      RECT -30.845 -18.735 -30.745 -18.315 ;
      RECT -30.845 -17.215 -30.745 -16.795 ;
      RECT -30.845 -12.455 -30.745 -11.855 ;
      RECT -30.845 -10.755 -30.745 -10.155 ;
      RECT -30.845 -5.815 -30.745 -5.395 ;
      RECT -30.845 -4.295 -30.745 -3.875 ;
      RECT -30.845 0.465 -30.745 1.065 ;
      RECT -31.365 -96.435 -31.265 -95.835 ;
      RECT -31.365 -94.735 -31.265 -94.135 ;
      RECT -31.365 -83.515 -31.265 -82.915 ;
      RECT -31.365 -81.815 -31.265 -81.215 ;
      RECT -31.365 -70.595 -31.265 -69.995 ;
      RECT -31.365 -68.895 -31.265 -68.295 ;
      RECT -31.365 -57.675 -31.265 -57.075 ;
      RECT -31.365 -55.975 -31.265 -55.375 ;
      RECT -31.365 -44.755 -31.265 -44.155 ;
      RECT -31.365 -43.055 -31.265 -42.455 ;
      RECT -31.365 -31.835 -31.265 -31.235 ;
      RECT -31.365 -30.135 -31.265 -29.535 ;
      RECT -31.365 -18.915 -31.265 -18.315 ;
      RECT -31.365 -17.215 -31.265 -16.615 ;
      RECT -31.365 -5.995 -31.265 -5.395 ;
      RECT -31.365 -4.295 -31.265 -3.695 ;
      RECT -31.625 -96.435 -31.525 -95.835 ;
      RECT -31.625 -94.735 -31.525 -94.135 ;
      RECT -31.625 -83.515 -31.525 -82.915 ;
      RECT -31.625 -81.815 -31.525 -81.215 ;
      RECT -31.625 -70.595 -31.525 -69.995 ;
      RECT -31.625 -68.895 -31.525 -68.295 ;
      RECT -31.625 -57.675 -31.525 -57.075 ;
      RECT -31.625 -55.975 -31.525 -55.375 ;
      RECT -31.625 -44.755 -31.525 -44.155 ;
      RECT -31.625 -43.055 -31.525 -42.455 ;
      RECT -31.625 -31.835 -31.525 -31.235 ;
      RECT -31.625 -30.135 -31.525 -29.535 ;
      RECT -31.625 -18.915 -31.525 -18.315 ;
      RECT -31.625 -17.215 -31.525 -16.615 ;
      RECT -31.625 -5.995 -31.525 -5.395 ;
      RECT -31.625 -4.295 -31.525 -3.695 ;
      RECT -32.245 2.165 -32.145 2.645 ;
      RECT -32.245 4.985 -32.145 5.405 ;
      RECT -32.845 2.165 -32.745 2.645 ;
      RECT -32.845 4.985 -32.745 5.405 ;
      RECT -33.445 2.165 -33.345 2.645 ;
      RECT -33.445 4.985 -33.345 5.405 ;
      RECT -34.045 2.165 -33.945 2.645 ;
      RECT -34.045 4.985 -33.945 5.405 ;
      RECT -34.645 2.165 -34.545 2.645 ;
      RECT -34.645 4.985 -34.545 5.405 ;
      RECT -35.245 2.165 -35.145 2.645 ;
      RECT -35.245 4.985 -35.145 5.405 ;
    LAYER M2 SPACING 0.16 ;
      RECT 151.695 -109.775 151.83 -109.275 ;
      RECT 151.695 -109.775 152.975 -109.67 ;
      RECT 152.875 -112.205 152.975 -109.67 ;
      RECT 151.36 -109.775 151.505 -109.275 ;
      RECT 150.855 -109.775 151.505 -109.67 ;
      RECT 150.855 -112.205 150.955 -109.67 ;
      RECT 149.825 -113 149.925 -107.215 ;
      RECT 149.465 -113 149.925 -112.9 ;
      RECT 149.465 -113.47 149.565 -112.9 ;
      RECT 149.115 -112.015 149.215 -110.555 ;
      RECT 149.075 -111.495 149.255 -111.395 ;
      RECT 146.895 -109.775 147.03 -109.275 ;
      RECT 146.895 -109.775 148.175 -109.67 ;
      RECT 148.075 -112.205 148.175 -109.67 ;
      RECT 146.56 -109.775 146.705 -109.275 ;
      RECT 146.055 -109.775 146.705 -109.67 ;
      RECT 146.055 -112.205 146.155 -109.67 ;
      RECT 145.025 -113 145.125 -107.215 ;
      RECT 144.665 -113 145.125 -112.9 ;
      RECT 144.665 -113.47 144.765 -112.9 ;
      RECT 144.315 -112.015 144.415 -110.555 ;
      RECT 144.275 -111.495 144.455 -111.395 ;
      RECT 142.095 -109.775 142.23 -109.275 ;
      RECT 142.095 -109.775 143.375 -109.67 ;
      RECT 143.275 -112.205 143.375 -109.67 ;
      RECT 141.76 -109.775 141.905 -109.275 ;
      RECT 141.255 -109.775 141.905 -109.67 ;
      RECT 141.255 -112.205 141.355 -109.67 ;
      RECT 140.225 -113 140.325 -107.215 ;
      RECT 139.865 -113 140.325 -112.9 ;
      RECT 139.865 -113.47 139.965 -112.9 ;
      RECT 139.515 -112.015 139.615 -110.555 ;
      RECT 139.475 -111.495 139.655 -111.395 ;
      RECT 137.295 -109.775 137.43 -109.275 ;
      RECT 137.295 -109.775 138.575 -109.67 ;
      RECT 138.475 -112.205 138.575 -109.67 ;
      RECT 136.96 -109.775 137.105 -109.275 ;
      RECT 136.455 -109.775 137.105 -109.67 ;
      RECT 136.455 -112.205 136.555 -109.67 ;
      RECT 135.425 -113 135.525 -107.215 ;
      RECT 135.065 -113 135.525 -112.9 ;
      RECT 135.065 -113.47 135.165 -112.9 ;
      RECT 134.715 -112.015 134.815 -110.555 ;
      RECT 134.675 -111.495 134.855 -111.395 ;
      RECT 132.495 -109.775 132.63 -109.275 ;
      RECT 132.495 -109.775 133.775 -109.67 ;
      RECT 133.675 -112.205 133.775 -109.67 ;
      RECT 132.16 -109.775 132.305 -109.275 ;
      RECT 131.655 -109.775 132.305 -109.67 ;
      RECT 131.655 -112.205 131.755 -109.67 ;
      RECT 130.625 -113 130.725 -107.215 ;
      RECT 130.265 -113 130.725 -112.9 ;
      RECT 130.265 -113.47 130.365 -112.9 ;
      RECT 129.915 -112.015 130.015 -110.555 ;
      RECT 129.875 -111.495 130.055 -111.395 ;
      RECT 127.695 -109.775 127.83 -109.275 ;
      RECT 127.695 -109.775 128.975 -109.67 ;
      RECT 128.875 -112.205 128.975 -109.67 ;
      RECT 127.36 -109.775 127.505 -109.275 ;
      RECT 126.855 -109.775 127.505 -109.67 ;
      RECT 126.855 -112.205 126.955 -109.67 ;
      RECT 125.825 -113 125.925 -107.215 ;
      RECT 125.465 -113 125.925 -112.9 ;
      RECT 125.465 -113.47 125.565 -112.9 ;
      RECT 125.115 -112.015 125.215 -110.555 ;
      RECT 125.075 -111.495 125.255 -111.395 ;
      RECT 122.895 -109.775 123.03 -109.275 ;
      RECT 122.895 -109.775 124.175 -109.67 ;
      RECT 124.075 -112.205 124.175 -109.67 ;
      RECT 122.56 -109.775 122.705 -109.275 ;
      RECT 122.055 -109.775 122.705 -109.67 ;
      RECT 122.055 -112.205 122.155 -109.67 ;
      RECT 121.025 -113 121.125 -107.215 ;
      RECT 120.665 -113 121.125 -112.9 ;
      RECT 120.665 -113.47 120.765 -112.9 ;
      RECT 120.315 -112.015 120.415 -110.555 ;
      RECT 120.275 -111.495 120.455 -111.395 ;
      RECT 118.095 -109.775 118.23 -109.275 ;
      RECT 118.095 -109.775 119.375 -109.67 ;
      RECT 119.275 -112.205 119.375 -109.67 ;
      RECT 117.76 -109.775 117.905 -109.275 ;
      RECT 117.255 -109.775 117.905 -109.67 ;
      RECT 117.255 -112.205 117.355 -109.67 ;
      RECT 116.225 -113 116.325 -107.215 ;
      RECT 115.865 -113 116.325 -112.9 ;
      RECT 115.865 -113.47 115.965 -112.9 ;
      RECT 115.515 -112.015 115.615 -110.555 ;
      RECT 115.475 -111.495 115.655 -111.395 ;
      RECT 113.295 -109.775 113.43 -109.275 ;
      RECT 113.295 -109.775 114.575 -109.67 ;
      RECT 114.475 -112.205 114.575 -109.67 ;
      RECT 112.96 -109.775 113.105 -109.275 ;
      RECT 112.455 -109.775 113.105 -109.67 ;
      RECT 112.455 -112.205 112.555 -109.67 ;
      RECT 111.425 -113 111.525 -107.215 ;
      RECT 111.065 -113 111.525 -112.9 ;
      RECT 111.065 -113.47 111.165 -112.9 ;
      RECT 110.715 -112.015 110.815 -110.555 ;
      RECT 110.675 -111.495 110.855 -111.395 ;
      RECT 108.495 -109.775 108.63 -109.275 ;
      RECT 108.495 -109.775 109.775 -109.67 ;
      RECT 109.675 -112.205 109.775 -109.67 ;
      RECT 108.16 -109.775 108.305 -109.275 ;
      RECT 107.655 -109.775 108.305 -109.67 ;
      RECT 107.655 -112.205 107.755 -109.67 ;
      RECT 106.625 -113 106.725 -107.215 ;
      RECT 106.265 -113 106.725 -112.9 ;
      RECT 106.265 -113.47 106.365 -112.9 ;
      RECT 105.915 -112.015 106.015 -110.555 ;
      RECT 105.875 -111.495 106.055 -111.395 ;
      RECT 103.695 -109.775 103.83 -109.275 ;
      RECT 103.695 -109.775 104.975 -109.67 ;
      RECT 104.875 -112.205 104.975 -109.67 ;
      RECT 103.36 -109.775 103.505 -109.275 ;
      RECT 102.855 -109.775 103.505 -109.67 ;
      RECT 102.855 -112.205 102.955 -109.67 ;
      RECT 101.825 -113 101.925 -107.215 ;
      RECT 101.465 -113 101.925 -112.9 ;
      RECT 101.465 -113.47 101.565 -112.9 ;
      RECT 101.115 -112.015 101.215 -110.555 ;
      RECT 101.075 -111.495 101.255 -111.395 ;
      RECT 98.895 -109.775 99.03 -109.275 ;
      RECT 98.895 -109.775 100.175 -109.67 ;
      RECT 100.075 -112.205 100.175 -109.67 ;
      RECT 98.56 -109.775 98.705 -109.275 ;
      RECT 98.055 -109.775 98.705 -109.67 ;
      RECT 98.055 -112.205 98.155 -109.67 ;
      RECT 97.025 -113 97.125 -107.215 ;
      RECT 96.665 -113 97.125 -112.9 ;
      RECT 96.665 -113.47 96.765 -112.9 ;
      RECT 96.315 -112.015 96.415 -110.555 ;
      RECT 96.275 -111.495 96.455 -111.395 ;
      RECT 94.095 -109.775 94.23 -109.275 ;
      RECT 94.095 -109.775 95.375 -109.67 ;
      RECT 95.275 -112.205 95.375 -109.67 ;
      RECT 93.76 -109.775 93.905 -109.275 ;
      RECT 93.255 -109.775 93.905 -109.67 ;
      RECT 93.255 -112.205 93.355 -109.67 ;
      RECT 92.225 -113 92.325 -107.215 ;
      RECT 91.865 -113 92.325 -112.9 ;
      RECT 91.865 -113.47 91.965 -112.9 ;
      RECT 91.515 -112.015 91.615 -110.555 ;
      RECT 91.475 -111.495 91.655 -111.395 ;
      RECT 89.295 -109.775 89.43 -109.275 ;
      RECT 89.295 -109.775 90.575 -109.67 ;
      RECT 90.475 -112.205 90.575 -109.67 ;
      RECT 88.96 -109.775 89.105 -109.275 ;
      RECT 88.455 -109.775 89.105 -109.67 ;
      RECT 88.455 -112.205 88.555 -109.67 ;
      RECT 87.425 -113 87.525 -107.215 ;
      RECT 87.065 -113 87.525 -112.9 ;
      RECT 87.065 -113.47 87.165 -112.9 ;
      RECT 86.715 -112.015 86.815 -110.555 ;
      RECT 86.675 -111.495 86.855 -111.395 ;
      RECT 84.495 -109.775 84.63 -109.275 ;
      RECT 84.495 -109.775 85.775 -109.67 ;
      RECT 85.675 -112.205 85.775 -109.67 ;
      RECT 84.16 -109.775 84.305 -109.275 ;
      RECT 83.655 -109.775 84.305 -109.67 ;
      RECT 83.655 -112.205 83.755 -109.67 ;
      RECT 82.625 -113 82.725 -107.215 ;
      RECT 82.265 -113 82.725 -112.9 ;
      RECT 82.265 -113.47 82.365 -112.9 ;
      RECT 81.915 -112.015 82.015 -110.555 ;
      RECT 81.875 -111.495 82.055 -111.395 ;
      RECT 79.695 -109.775 79.83 -109.275 ;
      RECT 79.695 -109.775 80.975 -109.67 ;
      RECT 80.875 -112.205 80.975 -109.67 ;
      RECT 79.36 -109.775 79.505 -109.275 ;
      RECT 78.855 -109.775 79.505 -109.67 ;
      RECT 78.855 -112.205 78.955 -109.67 ;
      RECT 77.825 -113 77.925 -107.215 ;
      RECT 77.465 -113 77.925 -112.9 ;
      RECT 77.465 -113.47 77.565 -112.9 ;
      RECT 77.115 -112.015 77.215 -110.555 ;
      RECT 77.075 -111.495 77.255 -111.395 ;
      RECT 74.895 -109.775 75.03 -109.275 ;
      RECT 74.895 -109.775 76.175 -109.67 ;
      RECT 76.075 -112.205 76.175 -109.67 ;
      RECT 74.56 -109.775 74.705 -109.275 ;
      RECT 74.055 -109.775 74.705 -109.67 ;
      RECT 74.055 -112.205 74.155 -109.67 ;
      RECT 73.025 -113 73.125 -107.215 ;
      RECT 72.665 -113 73.125 -112.9 ;
      RECT 72.665 -113.47 72.765 -112.9 ;
      RECT 72.315 -112.015 72.415 -110.555 ;
      RECT 72.275 -111.495 72.455 -111.395 ;
      RECT 70.095 -109.775 70.23 -109.275 ;
      RECT 70.095 -109.775 71.375 -109.67 ;
      RECT 71.275 -112.205 71.375 -109.67 ;
      RECT 69.76 -109.775 69.905 -109.275 ;
      RECT 69.255 -109.775 69.905 -109.67 ;
      RECT 69.255 -112.205 69.355 -109.67 ;
      RECT 68.225 -113 68.325 -107.215 ;
      RECT 67.865 -113 68.325 -112.9 ;
      RECT 67.865 -113.47 67.965 -112.9 ;
      RECT 67.515 -112.015 67.615 -110.555 ;
      RECT 67.475 -111.495 67.655 -111.395 ;
      RECT 65.295 -109.775 65.43 -109.275 ;
      RECT 65.295 -109.775 66.575 -109.67 ;
      RECT 66.475 -112.205 66.575 -109.67 ;
      RECT 64.96 -109.775 65.105 -109.275 ;
      RECT 64.455 -109.775 65.105 -109.67 ;
      RECT 64.455 -112.205 64.555 -109.67 ;
      RECT 63.425 -113 63.525 -107.215 ;
      RECT 63.065 -113 63.525 -112.9 ;
      RECT 63.065 -113.47 63.165 -112.9 ;
      RECT 62.715 -112.015 62.815 -110.555 ;
      RECT 62.675 -111.495 62.855 -111.395 ;
      RECT 60.495 -109.775 60.63 -109.275 ;
      RECT 60.495 -109.775 61.775 -109.67 ;
      RECT 61.675 -112.205 61.775 -109.67 ;
      RECT 60.16 -109.775 60.305 -109.275 ;
      RECT 59.655 -109.775 60.305 -109.67 ;
      RECT 59.655 -112.205 59.755 -109.67 ;
      RECT 58.625 -113 58.725 -107.215 ;
      RECT 58.265 -113 58.725 -112.9 ;
      RECT 58.265 -113.47 58.365 -112.9 ;
      RECT 57.915 -112.015 58.015 -110.555 ;
      RECT 57.875 -111.495 58.055 -111.395 ;
      RECT 55.695 -109.775 55.83 -109.275 ;
      RECT 55.695 -109.775 56.975 -109.67 ;
      RECT 56.875 -112.205 56.975 -109.67 ;
      RECT 55.36 -109.775 55.505 -109.275 ;
      RECT 54.855 -109.775 55.505 -109.67 ;
      RECT 54.855 -112.205 54.955 -109.67 ;
      RECT 53.825 -113 53.925 -107.215 ;
      RECT 53.465 -113 53.925 -112.9 ;
      RECT 53.465 -113.47 53.565 -112.9 ;
      RECT 53.115 -112.015 53.215 -110.555 ;
      RECT 53.075 -111.495 53.255 -111.395 ;
      RECT 50.895 -109.775 51.03 -109.275 ;
      RECT 50.895 -109.775 52.175 -109.67 ;
      RECT 52.075 -112.205 52.175 -109.67 ;
      RECT 50.56 -109.775 50.705 -109.275 ;
      RECT 50.055 -109.775 50.705 -109.67 ;
      RECT 50.055 -112.205 50.155 -109.67 ;
      RECT 49.025 -113 49.125 -107.215 ;
      RECT 48.665 -113 49.125 -112.9 ;
      RECT 48.665 -113.47 48.765 -112.9 ;
      RECT 48.315 -112.015 48.415 -110.555 ;
      RECT 48.275 -111.495 48.455 -111.395 ;
      RECT 46.095 -109.775 46.23 -109.275 ;
      RECT 46.095 -109.775 47.375 -109.67 ;
      RECT 47.275 -112.205 47.375 -109.67 ;
      RECT 45.76 -109.775 45.905 -109.275 ;
      RECT 45.255 -109.775 45.905 -109.67 ;
      RECT 45.255 -112.205 45.355 -109.67 ;
      RECT 44.225 -113 44.325 -107.215 ;
      RECT 43.865 -113 44.325 -112.9 ;
      RECT 43.865 -113.47 43.965 -112.9 ;
      RECT 43.515 -112.015 43.615 -110.555 ;
      RECT 43.475 -111.495 43.655 -111.395 ;
      RECT 41.295 -109.775 41.43 -109.275 ;
      RECT 41.295 -109.775 42.575 -109.67 ;
      RECT 42.475 -112.205 42.575 -109.67 ;
      RECT 40.96 -109.775 41.105 -109.275 ;
      RECT 40.455 -109.775 41.105 -109.67 ;
      RECT 40.455 -112.205 40.555 -109.67 ;
      RECT 39.425 -113 39.525 -107.215 ;
      RECT 39.065 -113 39.525 -112.9 ;
      RECT 39.065 -113.47 39.165 -112.9 ;
      RECT 38.715 -112.015 38.815 -110.555 ;
      RECT 38.675 -111.495 38.855 -111.395 ;
      RECT 36.495 -109.775 36.63 -109.275 ;
      RECT 36.495 -109.775 37.775 -109.67 ;
      RECT 37.675 -112.205 37.775 -109.67 ;
      RECT 36.16 -109.775 36.305 -109.275 ;
      RECT 35.655 -109.775 36.305 -109.67 ;
      RECT 35.655 -112.205 35.755 -109.67 ;
      RECT 34.625 -113 34.725 -107.215 ;
      RECT 34.265 -113 34.725 -112.9 ;
      RECT 34.265 -113.47 34.365 -112.9 ;
      RECT 33.915 -112.015 34.015 -110.555 ;
      RECT 33.875 -111.495 34.055 -111.395 ;
      RECT 31.695 -109.775 31.83 -109.275 ;
      RECT 31.695 -109.775 32.975 -109.67 ;
      RECT 32.875 -112.205 32.975 -109.67 ;
      RECT 31.36 -109.775 31.505 -109.275 ;
      RECT 30.855 -109.775 31.505 -109.67 ;
      RECT 30.855 -112.205 30.955 -109.67 ;
      RECT 29.825 -113 29.925 -107.215 ;
      RECT 29.465 -113 29.925 -112.9 ;
      RECT 29.465 -113.47 29.565 -112.9 ;
      RECT 29.115 -112.015 29.215 -110.555 ;
      RECT 29.075 -111.495 29.255 -111.395 ;
      RECT 26.895 -109.775 27.03 -109.275 ;
      RECT 26.895 -109.775 28.175 -109.67 ;
      RECT 28.075 -112.205 28.175 -109.67 ;
      RECT 26.56 -109.775 26.705 -109.275 ;
      RECT 26.055 -109.775 26.705 -109.67 ;
      RECT 26.055 -112.205 26.155 -109.67 ;
      RECT 25.025 -113 25.125 -107.215 ;
      RECT 24.665 -113 25.125 -112.9 ;
      RECT 24.665 -113.47 24.765 -112.9 ;
      RECT 24.315 -112.015 24.415 -110.555 ;
      RECT 24.275 -111.495 24.455 -111.395 ;
      RECT 22.095 -109.775 22.23 -109.275 ;
      RECT 22.095 -109.775 23.375 -109.67 ;
      RECT 23.275 -112.205 23.375 -109.67 ;
      RECT 21.76 -109.775 21.905 -109.275 ;
      RECT 21.255 -109.775 21.905 -109.67 ;
      RECT 21.255 -112.205 21.355 -109.67 ;
      RECT 20.225 -113 20.325 -107.215 ;
      RECT 19.865 -113 20.325 -112.9 ;
      RECT 19.865 -113.47 19.965 -112.9 ;
      RECT 19.515 -112.015 19.615 -110.555 ;
      RECT 19.475 -111.495 19.655 -111.395 ;
      RECT 17.295 -109.775 17.43 -109.275 ;
      RECT 17.295 -109.775 18.575 -109.67 ;
      RECT 18.475 -112.205 18.575 -109.67 ;
      RECT 16.96 -109.775 17.105 -109.275 ;
      RECT 16.455 -109.775 17.105 -109.67 ;
      RECT 16.455 -112.205 16.555 -109.67 ;
      RECT 15.425 -113 15.525 -107.215 ;
      RECT 15.065 -113 15.525 -112.9 ;
      RECT 15.065 -113.47 15.165 -112.9 ;
      RECT 14.715 -112.015 14.815 -110.555 ;
      RECT 14.675 -111.495 14.855 -111.395 ;
      RECT 12.495 -109.775 12.63 -109.275 ;
      RECT 12.495 -109.775 13.775 -109.67 ;
      RECT 13.675 -112.205 13.775 -109.67 ;
      RECT 12.16 -109.775 12.305 -109.275 ;
      RECT 11.655 -109.775 12.305 -109.67 ;
      RECT 11.655 -112.205 11.755 -109.67 ;
      RECT 10.625 -113 10.725 -107.215 ;
      RECT 10.265 -113 10.725 -112.9 ;
      RECT 10.265 -113.47 10.365 -112.9 ;
      RECT 9.915 -112.015 10.015 -110.555 ;
      RECT 9.875 -111.495 10.055 -111.395 ;
      RECT 7.695 -109.775 7.83 -109.275 ;
      RECT 7.695 -109.775 8.975 -109.67 ;
      RECT 8.875 -112.205 8.975 -109.67 ;
      RECT 7.36 -109.775 7.505 -109.275 ;
      RECT 6.855 -109.775 7.505 -109.67 ;
      RECT 6.855 -112.205 6.955 -109.67 ;
      RECT 5.825 -113 5.925 -107.215 ;
      RECT 5.465 -113 5.925 -112.9 ;
      RECT 5.465 -113.47 5.565 -112.9 ;
      RECT 5.115 -112.015 5.215 -110.555 ;
      RECT 5.075 -111.495 5.255 -111.395 ;
      RECT 2.895 -109.775 3.03 -109.275 ;
      RECT 2.895 -109.775 4.175 -109.67 ;
      RECT 4.075 -112.205 4.175 -109.67 ;
      RECT 2.56 -109.775 2.705 -109.275 ;
      RECT 2.055 -109.775 2.705 -109.67 ;
      RECT 2.055 -112.205 2.155 -109.67 ;
      RECT 1.025 -113 1.125 -107.215 ;
      RECT 0.665 -113 1.125 -112.9 ;
      RECT 0.665 -113.47 0.765 -112.9 ;
      RECT 0.315 -112.015 0.415 -110.555 ;
      RECT 0.275 -111.495 0.455 -111.395 ;
      RECT -11.445 -107.175 -11.265 -102.715 ;
      RECT -11.445 -110.635 -11.345 -102.715 ;
      RECT -12.045 -107.175 -11.865 -102.715 ;
      RECT -12.045 -110.635 -11.945 -102.715 ;
      RECT -32.245 -100.715 -32.145 5.405 ;
      RECT -32.245 -100.715 -32.065 0.645 ;
      RECT -32.845 -100.715 -32.745 5.405 ;
      RECT -32.845 -100.715 -32.665 0.645 ;
      RECT -33.445 -100.715 -33.345 5.405 ;
      RECT -33.445 -100.715 -33.265 0.645 ;
      RECT -34.045 -100.715 -33.945 5.405 ;
      RECT -34.045 -100.715 -33.865 0.645 ;
      RECT -34.645 -100.715 -34.545 5.405 ;
      RECT -34.645 -100.715 -34.465 0.645 ;
      RECT -35.245 -100.715 -35.145 5.405 ;
      RECT -35.245 -100.715 -35.065 0.645 ;
      RECT 157.465 -116.645 158.465 9.895 ;
      RECT 155.465 -120.365 156.465 5.175 ;
      RECT 153.55 -101.845 153.65 9.895 ;
      RECT 153.425 -108.965 153.525 -103.985 ;
      RECT 153.165 -104.945 153.265 3.135 ;
      RECT 152.735 -104.945 152.835 3.135 ;
      RECT 152.475 -108.685 152.575 -103.985 ;
      RECT 152.35 -101.845 152.45 9.895 ;
      RECT 152.285 -111.985 152.385 -110.37 ;
      RECT 152.225 -108.965 152.325 -103.985 ;
      RECT 151.985 -109.19 152.085 -108.505 ;
      RECT 151.965 -104.945 152.065 3.135 ;
      RECT 151.535 -104.945 151.635 3.135 ;
      RECT 151.275 -108.685 151.375 -103.985 ;
      RECT 151.15 -101.845 151.25 9.895 ;
      RECT 151.025 -108.965 151.125 -107.215 ;
      RECT 150.765 -108.175 150.865 3.135 ;
      RECT 150.335 -108.175 150.435 3.135 ;
      RECT 150.265 -111.985 150.365 -110.385 ;
      RECT 150.075 -108.685 150.175 -107.215 ;
      RECT 149.95 -101.845 150.05 9.895 ;
      RECT 149.565 -108.175 149.665 3.135 ;
      RECT 149.135 -108.175 149.235 3.135 ;
      RECT 148.875 -113.47 148.975 -107.215 ;
      RECT 148.75 -101.845 148.85 9.895 ;
      RECT 148.625 -108.965 148.725 -103.985 ;
      RECT 148.365 -104.945 148.465 3.135 ;
      RECT 147.935 -104.945 148.035 3.135 ;
      RECT 147.675 -108.685 147.775 -103.985 ;
      RECT 147.55 -101.845 147.65 9.895 ;
      RECT 147.485 -111.985 147.585 -110.37 ;
      RECT 147.425 -108.965 147.525 -103.985 ;
      RECT 147.185 -109.19 147.285 -108.505 ;
      RECT 147.165 -104.945 147.265 3.135 ;
      RECT 146.735 -104.945 146.835 3.135 ;
      RECT 146.475 -108.685 146.575 -103.985 ;
      RECT 146.35 -101.845 146.45 9.895 ;
      RECT 146.225 -108.965 146.325 -107.215 ;
      RECT 145.965 -108.175 146.065 3.135 ;
      RECT 145.535 -108.175 145.635 3.135 ;
      RECT 145.465 -111.985 145.565 -110.385 ;
      RECT 145.275 -108.685 145.375 -107.215 ;
      RECT 145.15 -101.845 145.25 9.895 ;
      RECT 144.765 -108.175 144.865 3.135 ;
      RECT 144.335 -108.175 144.435 3.135 ;
      RECT 144.075 -113.47 144.175 -107.215 ;
      RECT 143.95 -101.845 144.05 9.895 ;
      RECT 143.825 -108.965 143.925 -103.985 ;
      RECT 143.565 -104.945 143.665 3.135 ;
      RECT 143.135 -104.945 143.235 3.135 ;
      RECT 142.875 -108.685 142.975 -103.985 ;
      RECT 142.75 -101.845 142.85 9.895 ;
      RECT 142.685 -111.985 142.785 -110.37 ;
      RECT 142.625 -108.965 142.725 -103.985 ;
      RECT 142.385 -109.19 142.485 -108.505 ;
      RECT 142.365 -104.945 142.465 3.135 ;
      RECT 141.935 -104.945 142.035 3.135 ;
      RECT 141.675 -108.685 141.775 -103.985 ;
      RECT 141.55 -101.845 141.65 9.895 ;
      RECT 141.425 -108.965 141.525 -107.215 ;
      RECT 141.165 -108.175 141.265 3.135 ;
      RECT 140.735 -108.175 140.835 3.135 ;
      RECT 140.665 -111.985 140.765 -110.385 ;
      RECT 140.475 -108.685 140.575 -107.215 ;
      RECT 140.35 -101.845 140.45 9.895 ;
      RECT 139.965 -108.175 140.065 3.135 ;
      RECT 139.535 -108.175 139.635 3.135 ;
      RECT 139.275 -113.47 139.375 -107.215 ;
      RECT 139.15 -101.845 139.25 9.895 ;
      RECT 139.025 -108.965 139.125 -103.985 ;
      RECT 138.765 -104.945 138.865 3.135 ;
      RECT 138.335 -104.945 138.435 3.135 ;
      RECT 138.075 -108.685 138.175 -103.985 ;
      RECT 137.95 -101.845 138.05 9.895 ;
      RECT 137.885 -111.985 137.985 -110.37 ;
      RECT 137.825 -108.965 137.925 -103.985 ;
      RECT 137.585 -109.19 137.685 -108.505 ;
      RECT 137.565 -104.945 137.665 3.135 ;
      RECT 137.135 -104.945 137.235 3.135 ;
      RECT 136.875 -108.685 136.975 -103.985 ;
      RECT 136.75 -101.845 136.85 9.895 ;
      RECT 136.625 -108.965 136.725 -107.215 ;
      RECT 136.365 -108.175 136.465 3.135 ;
      RECT 135.935 -108.175 136.035 3.135 ;
      RECT 135.865 -111.985 135.965 -110.385 ;
      RECT 135.675 -108.685 135.775 -107.215 ;
      RECT 135.55 -101.845 135.65 9.895 ;
      RECT 135.165 -108.175 135.265 3.135 ;
      RECT 134.735 -108.175 134.835 3.135 ;
      RECT 134.475 -113.47 134.575 -107.215 ;
      RECT 134.35 -101.845 134.45 9.895 ;
      RECT 134.225 -108.965 134.325 -103.985 ;
      RECT 133.965 -104.945 134.065 3.135 ;
      RECT 133.535 -104.945 133.635 3.135 ;
      RECT 133.275 -108.685 133.375 -103.985 ;
      RECT 133.15 -101.845 133.25 9.895 ;
      RECT 133.085 -111.985 133.185 -110.37 ;
      RECT 133.025 -108.965 133.125 -103.985 ;
      RECT 132.785 -109.19 132.885 -108.505 ;
      RECT 132.765 -104.945 132.865 3.135 ;
      RECT 132.335 -104.945 132.435 3.135 ;
      RECT 132.075 -108.685 132.175 -103.985 ;
      RECT 131.95 -101.845 132.05 9.895 ;
      RECT 131.825 -108.965 131.925 -107.215 ;
      RECT 131.565 -108.175 131.665 3.135 ;
      RECT 131.135 -108.175 131.235 3.135 ;
      RECT 131.065 -111.985 131.165 -110.385 ;
      RECT 130.875 -108.685 130.975 -107.215 ;
      RECT 130.75 -101.845 130.85 9.895 ;
      RECT 130.365 -108.175 130.465 3.135 ;
      RECT 129.935 -108.175 130.035 3.135 ;
      RECT 129.675 -113.47 129.775 -107.215 ;
      RECT 129.55 -101.845 129.65 9.895 ;
      RECT 129.425 -108.965 129.525 -103.985 ;
      RECT 129.165 -104.945 129.265 3.135 ;
      RECT 128.735 -104.945 128.835 3.135 ;
      RECT 128.475 -108.685 128.575 -103.985 ;
      RECT 128.35 -101.845 128.45 9.895 ;
      RECT 128.285 -111.985 128.385 -110.37 ;
      RECT 128.225 -108.965 128.325 -103.985 ;
      RECT 127.985 -109.19 128.085 -108.505 ;
      RECT 127.965 -104.945 128.065 3.135 ;
      RECT 127.535 -104.945 127.635 3.135 ;
      RECT 127.275 -108.685 127.375 -103.985 ;
      RECT 127.15 -101.845 127.25 9.895 ;
      RECT 127.025 -108.965 127.125 -107.215 ;
      RECT 126.765 -108.175 126.865 3.135 ;
      RECT 126.335 -108.175 126.435 3.135 ;
      RECT 126.265 -111.985 126.365 -110.385 ;
      RECT 126.075 -108.685 126.175 -107.215 ;
      RECT 125.95 -101.845 126.05 9.895 ;
      RECT 125.565 -108.175 125.665 3.135 ;
      RECT 125.135 -108.175 125.235 3.135 ;
      RECT 124.875 -113.47 124.975 -107.215 ;
      RECT 124.75 -101.845 124.85 9.895 ;
      RECT 124.625 -108.965 124.725 -103.985 ;
      RECT 124.365 -104.945 124.465 3.135 ;
      RECT 123.935 -104.945 124.035 3.135 ;
      RECT 123.675 -108.685 123.775 -103.985 ;
      RECT 123.55 -101.845 123.65 9.895 ;
      RECT 123.485 -111.985 123.585 -110.37 ;
      RECT 123.425 -108.965 123.525 -103.985 ;
      RECT 123.185 -109.19 123.285 -108.505 ;
      RECT 123.165 -104.945 123.265 3.135 ;
      RECT 122.735 -104.945 122.835 3.135 ;
      RECT 122.475 -108.685 122.575 -103.985 ;
      RECT 122.35 -101.845 122.45 9.895 ;
      RECT 122.225 -108.965 122.325 -107.215 ;
      RECT 121.965 -108.175 122.065 3.135 ;
      RECT 121.535 -108.175 121.635 3.135 ;
      RECT 121.465 -111.985 121.565 -110.385 ;
      RECT 121.275 -108.685 121.375 -107.215 ;
      RECT 121.15 -101.845 121.25 9.895 ;
      RECT 120.765 -108.175 120.865 3.135 ;
      RECT 120.335 -108.175 120.435 3.135 ;
      RECT 120.075 -113.47 120.175 -107.215 ;
      RECT 119.95 -101.845 120.05 9.895 ;
      RECT 119.825 -108.965 119.925 -103.985 ;
      RECT 119.565 -104.945 119.665 3.135 ;
      RECT 119.135 -104.945 119.235 3.135 ;
      RECT 118.875 -108.685 118.975 -103.985 ;
      RECT 118.75 -101.845 118.85 9.895 ;
      RECT 118.685 -111.985 118.785 -110.37 ;
      RECT 118.625 -108.965 118.725 -103.985 ;
      RECT 118.385 -109.19 118.485 -108.505 ;
      RECT 118.365 -104.945 118.465 3.135 ;
      RECT 117.935 -104.945 118.035 3.135 ;
      RECT 117.675 -108.685 117.775 -103.985 ;
      RECT 117.55 -101.845 117.65 9.895 ;
      RECT 117.425 -108.965 117.525 -107.215 ;
      RECT 117.165 -108.175 117.265 3.135 ;
      RECT 116.735 -108.175 116.835 3.135 ;
      RECT 116.665 -111.985 116.765 -110.385 ;
      RECT 116.475 -108.685 116.575 -107.215 ;
      RECT 116.35 -101.845 116.45 9.895 ;
      RECT 115.965 -108.175 116.065 3.135 ;
      RECT 115.535 -108.175 115.635 3.135 ;
      RECT 115.275 -113.47 115.375 -107.215 ;
      RECT 115.15 -101.845 115.25 9.895 ;
      RECT 115.025 -108.965 115.125 -103.985 ;
      RECT 114.765 -104.945 114.865 3.135 ;
      RECT 114.335 -104.945 114.435 3.135 ;
      RECT 114.075 -108.685 114.175 -103.985 ;
      RECT 113.95 -101.845 114.05 9.895 ;
      RECT 113.885 -111.985 113.985 -110.37 ;
      RECT 113.825 -108.965 113.925 -103.985 ;
      RECT 113.585 -109.19 113.685 -108.505 ;
      RECT 113.565 -104.945 113.665 3.135 ;
      RECT 113.135 -104.945 113.235 3.135 ;
      RECT 112.875 -108.685 112.975 -103.985 ;
      RECT 112.75 -101.845 112.85 9.895 ;
      RECT 112.625 -108.965 112.725 -107.215 ;
      RECT 112.365 -108.175 112.465 3.135 ;
      RECT 111.935 -108.175 112.035 3.135 ;
      RECT 111.865 -111.985 111.965 -110.385 ;
      RECT 111.675 -108.685 111.775 -107.215 ;
      RECT 111.55 -101.845 111.65 9.895 ;
      RECT 111.165 -108.175 111.265 3.135 ;
      RECT 110.735 -108.175 110.835 3.135 ;
      RECT 110.475 -113.47 110.575 -107.215 ;
      RECT 110.35 -101.845 110.45 9.895 ;
      RECT 110.225 -108.965 110.325 -103.985 ;
      RECT 109.965 -104.945 110.065 3.135 ;
      RECT 109.535 -104.945 109.635 3.135 ;
      RECT 109.275 -108.685 109.375 -103.985 ;
      RECT 109.15 -101.845 109.25 9.895 ;
      RECT 109.085 -111.985 109.185 -110.37 ;
      RECT 109.025 -108.965 109.125 -103.985 ;
      RECT 108.785 -109.19 108.885 -108.505 ;
      RECT 108.765 -104.945 108.865 3.135 ;
      RECT 108.335 -104.945 108.435 3.135 ;
      RECT 108.075 -108.685 108.175 -103.985 ;
      RECT 107.95 -101.845 108.05 9.895 ;
      RECT 107.825 -108.965 107.925 -107.215 ;
      RECT 107.565 -108.175 107.665 3.135 ;
      RECT 107.135 -108.175 107.235 3.135 ;
      RECT 107.065 -111.985 107.165 -110.385 ;
      RECT 106.875 -108.685 106.975 -107.215 ;
      RECT 106.75 -101.845 106.85 9.895 ;
      RECT 106.365 -108.175 106.465 3.135 ;
      RECT 105.935 -108.175 106.035 3.135 ;
      RECT 105.675 -113.47 105.775 -107.215 ;
      RECT 105.55 -101.845 105.65 9.895 ;
      RECT 105.425 -108.965 105.525 -103.985 ;
      RECT 105.165 -104.945 105.265 3.135 ;
      RECT 104.735 -104.945 104.835 3.135 ;
      RECT 104.475 -108.685 104.575 -103.985 ;
      RECT 104.35 -101.845 104.45 9.895 ;
      RECT 104.285 -111.985 104.385 -110.37 ;
      RECT 104.225 -108.965 104.325 -103.985 ;
      RECT 103.985 -109.19 104.085 -108.505 ;
      RECT 103.965 -104.945 104.065 3.135 ;
      RECT 103.535 -104.945 103.635 3.135 ;
      RECT 103.275 -108.685 103.375 -103.985 ;
      RECT 103.15 -101.845 103.25 9.895 ;
      RECT 103.025 -108.965 103.125 -107.215 ;
      RECT 102.765 -108.175 102.865 3.135 ;
      RECT 102.335 -108.175 102.435 3.135 ;
      RECT 102.265 -111.985 102.365 -110.385 ;
      RECT 102.075 -108.685 102.175 -107.215 ;
      RECT 101.95 -101.845 102.05 9.895 ;
      RECT 101.565 -108.175 101.665 3.135 ;
      RECT 101.135 -108.175 101.235 3.135 ;
      RECT 100.875 -113.47 100.975 -107.215 ;
      RECT 100.75 -101.845 100.85 9.895 ;
      RECT 100.625 -108.965 100.725 -103.985 ;
      RECT 100.365 -104.945 100.465 3.135 ;
      RECT 99.935 -104.945 100.035 3.135 ;
      RECT 99.675 -108.685 99.775 -103.985 ;
      RECT 99.55 -101.845 99.65 9.895 ;
      RECT 99.485 -111.985 99.585 -110.37 ;
      RECT 99.425 -108.965 99.525 -103.985 ;
      RECT 99.185 -109.19 99.285 -108.505 ;
      RECT 99.165 -104.945 99.265 3.135 ;
      RECT 98.735 -104.945 98.835 3.135 ;
      RECT 98.475 -108.685 98.575 -103.985 ;
      RECT 98.35 -101.845 98.45 9.895 ;
      RECT 98.225 -108.965 98.325 -107.215 ;
      RECT 97.965 -108.175 98.065 3.135 ;
      RECT 97.535 -108.175 97.635 3.135 ;
      RECT 97.465 -111.985 97.565 -110.385 ;
      RECT 97.275 -108.685 97.375 -107.215 ;
      RECT 97.15 -101.845 97.25 9.895 ;
      RECT 96.765 -108.175 96.865 3.135 ;
      RECT 96.335 -108.175 96.435 3.135 ;
      RECT 96.075 -113.47 96.175 -107.215 ;
      RECT 95.95 -101.845 96.05 9.895 ;
      RECT 95.825 -108.965 95.925 -103.985 ;
      RECT 95.565 -104.945 95.665 3.135 ;
      RECT 95.135 -104.945 95.235 3.135 ;
      RECT 94.875 -108.685 94.975 -103.985 ;
      RECT 94.75 -101.845 94.85 9.895 ;
      RECT 94.685 -111.985 94.785 -110.37 ;
      RECT 94.625 -108.965 94.725 -103.985 ;
      RECT 94.385 -109.19 94.485 -108.505 ;
      RECT 94.365 -104.945 94.465 3.135 ;
      RECT 93.935 -104.945 94.035 3.135 ;
      RECT 93.675 -108.685 93.775 -103.985 ;
      RECT 93.55 -101.845 93.65 9.895 ;
      RECT 93.425 -108.965 93.525 -107.215 ;
      RECT 93.165 -108.175 93.265 3.135 ;
      RECT 92.735 -108.175 92.835 3.135 ;
      RECT 92.665 -111.985 92.765 -110.385 ;
      RECT 92.475 -108.685 92.575 -107.215 ;
      RECT 92.35 -101.845 92.45 9.895 ;
      RECT 91.965 -108.175 92.065 3.135 ;
      RECT 91.535 -108.175 91.635 3.135 ;
      RECT 91.275 -113.47 91.375 -107.215 ;
      RECT 91.15 -101.845 91.25 9.895 ;
      RECT 91.025 -108.965 91.125 -103.985 ;
      RECT 90.765 -104.945 90.865 3.135 ;
      RECT 90.335 -104.945 90.435 3.135 ;
      RECT 90.075 -108.685 90.175 -103.985 ;
      RECT 89.95 -101.845 90.05 9.895 ;
      RECT 89.885 -111.985 89.985 -110.37 ;
      RECT 89.825 -108.965 89.925 -103.985 ;
      RECT 89.585 -109.19 89.685 -108.505 ;
      RECT 89.565 -104.945 89.665 3.135 ;
      RECT 89.135 -104.945 89.235 3.135 ;
      RECT 88.875 -108.685 88.975 -103.985 ;
      RECT 88.75 -101.845 88.85 9.895 ;
      RECT 88.625 -108.965 88.725 -107.215 ;
      RECT 88.365 -108.175 88.465 3.135 ;
      RECT 87.935 -108.175 88.035 3.135 ;
      RECT 87.865 -111.985 87.965 -110.385 ;
      RECT 87.675 -108.685 87.775 -107.215 ;
      RECT 87.55 -101.845 87.65 9.895 ;
      RECT 87.165 -108.175 87.265 3.135 ;
      RECT 86.735 -108.175 86.835 3.135 ;
      RECT 86.475 -113.47 86.575 -107.215 ;
      RECT 86.35 -101.845 86.45 9.895 ;
      RECT 86.225 -108.965 86.325 -103.985 ;
      RECT 85.965 -104.945 86.065 3.135 ;
      RECT 85.535 -104.945 85.635 3.135 ;
      RECT 85.275 -108.685 85.375 -103.985 ;
      RECT 85.15 -101.845 85.25 9.895 ;
      RECT 85.085 -111.985 85.185 -110.37 ;
      RECT 85.025 -108.965 85.125 -103.985 ;
      RECT 84.785 -109.19 84.885 -108.505 ;
      RECT 84.765 -104.945 84.865 3.135 ;
      RECT 84.335 -104.945 84.435 3.135 ;
      RECT 84.075 -108.685 84.175 -103.985 ;
      RECT 83.95 -101.845 84.05 9.895 ;
      RECT 83.825 -108.965 83.925 -107.215 ;
      RECT 83.565 -108.175 83.665 3.135 ;
      RECT 83.135 -108.175 83.235 3.135 ;
      RECT 83.065 -111.985 83.165 -110.385 ;
      RECT 82.875 -108.685 82.975 -107.215 ;
      RECT 82.75 -101.845 82.85 9.895 ;
      RECT 82.365 -108.175 82.465 3.135 ;
      RECT 81.935 -108.175 82.035 3.135 ;
      RECT 81.675 -113.47 81.775 -107.215 ;
      RECT 81.55 -101.845 81.65 9.895 ;
      RECT 81.425 -108.965 81.525 -103.985 ;
      RECT 81.165 -104.945 81.265 3.135 ;
      RECT 80.735 -104.945 80.835 3.135 ;
      RECT 80.475 -108.685 80.575 -103.985 ;
      RECT 80.35 -101.845 80.45 9.895 ;
      RECT 80.285 -111.985 80.385 -110.37 ;
      RECT 80.225 -108.965 80.325 -103.985 ;
      RECT 79.985 -109.19 80.085 -108.505 ;
      RECT 79.965 -104.945 80.065 3.135 ;
      RECT 79.535 -104.945 79.635 3.135 ;
      RECT 79.275 -108.685 79.375 -103.985 ;
      RECT 79.15 -101.845 79.25 9.895 ;
      RECT 79.025 -108.965 79.125 -107.215 ;
      RECT 78.765 -108.175 78.865 3.135 ;
      RECT 78.335 -108.175 78.435 3.135 ;
      RECT 78.265 -111.985 78.365 -110.385 ;
      RECT 78.075 -108.685 78.175 -107.215 ;
      RECT 77.95 -101.845 78.05 9.895 ;
      RECT 77.565 -108.175 77.665 3.135 ;
      RECT 77.135 -108.175 77.235 3.135 ;
      RECT 76.875 -113.47 76.975 -107.215 ;
      RECT 76.75 -101.845 76.85 9.895 ;
      RECT 76.625 -108.965 76.725 -103.985 ;
      RECT 76.365 -104.945 76.465 3.135 ;
      RECT 75.935 -104.945 76.035 3.135 ;
      RECT 75.675 -108.685 75.775 -103.985 ;
      RECT 75.55 -101.845 75.65 9.895 ;
      RECT 75.485 -111.985 75.585 -110.37 ;
      RECT 75.425 -108.965 75.525 -103.985 ;
      RECT 75.185 -109.19 75.285 -108.505 ;
      RECT 75.165 -104.945 75.265 3.135 ;
      RECT 74.735 -104.945 74.835 3.135 ;
      RECT 74.475 -108.685 74.575 -103.985 ;
      RECT 74.35 -101.845 74.45 9.895 ;
      RECT 74.225 -108.965 74.325 -107.215 ;
      RECT 73.965 -108.175 74.065 3.135 ;
      RECT 73.535 -108.175 73.635 3.135 ;
      RECT 73.465 -111.985 73.565 -110.385 ;
      RECT 73.275 -108.685 73.375 -107.215 ;
      RECT 73.15 -101.845 73.25 9.895 ;
      RECT 72.765 -108.175 72.865 3.135 ;
      RECT 72.335 -108.175 72.435 3.135 ;
      RECT 72.075 -113.47 72.175 -107.215 ;
      RECT 71.95 -101.845 72.05 9.895 ;
      RECT 71.825 -108.965 71.925 -103.985 ;
      RECT 71.565 -104.945 71.665 3.135 ;
      RECT 71.135 -104.945 71.235 3.135 ;
      RECT 70.875 -108.685 70.975 -103.985 ;
      RECT 70.75 -101.845 70.85 9.895 ;
      RECT 70.685 -111.985 70.785 -110.37 ;
      RECT 70.625 -108.965 70.725 -103.985 ;
      RECT 70.385 -109.19 70.485 -108.505 ;
      RECT 70.365 -104.945 70.465 3.135 ;
      RECT 69.935 -104.945 70.035 3.135 ;
      RECT 69.675 -108.685 69.775 -103.985 ;
      RECT 69.55 -101.845 69.65 9.895 ;
      RECT 69.425 -108.965 69.525 -107.215 ;
      RECT 69.165 -108.175 69.265 3.135 ;
      RECT 68.735 -108.175 68.835 3.135 ;
      RECT 68.665 -111.985 68.765 -110.385 ;
      RECT 68.475 -108.685 68.575 -107.215 ;
      RECT 68.35 -101.845 68.45 9.895 ;
      RECT 67.965 -108.175 68.065 3.135 ;
      RECT 67.535 -108.175 67.635 3.135 ;
      RECT 67.275 -113.47 67.375 -107.215 ;
      RECT 67.15 -101.845 67.25 9.895 ;
      RECT 67.025 -108.965 67.125 -103.985 ;
      RECT 66.765 -104.945 66.865 3.135 ;
      RECT 66.335 -104.945 66.435 3.135 ;
      RECT 66.075 -108.685 66.175 -103.985 ;
      RECT 65.95 -101.845 66.05 9.895 ;
      RECT 65.885 -111.985 65.985 -110.37 ;
      RECT 65.825 -108.965 65.925 -103.985 ;
      RECT 65.585 -109.19 65.685 -108.505 ;
      RECT 65.565 -104.945 65.665 3.135 ;
      RECT 65.135 -104.945 65.235 3.135 ;
      RECT 64.875 -108.685 64.975 -103.985 ;
      RECT 64.75 -101.845 64.85 9.895 ;
      RECT 64.625 -108.965 64.725 -107.215 ;
      RECT 64.365 -108.175 64.465 3.135 ;
      RECT 63.935 -108.175 64.035 3.135 ;
      RECT 63.865 -111.985 63.965 -110.385 ;
      RECT 63.675 -108.685 63.775 -107.215 ;
      RECT 63.55 -101.845 63.65 9.895 ;
      RECT 63.165 -108.175 63.265 3.135 ;
      RECT 62.735 -108.175 62.835 3.135 ;
      RECT 62.475 -113.47 62.575 -107.215 ;
      RECT 62.35 -101.845 62.45 9.895 ;
      RECT 62.225 -108.965 62.325 -103.985 ;
      RECT 61.965 -104.945 62.065 3.135 ;
      RECT 61.535 -104.945 61.635 3.135 ;
      RECT 61.275 -108.685 61.375 -103.985 ;
      RECT 61.15 -101.845 61.25 9.895 ;
      RECT 61.085 -111.985 61.185 -110.37 ;
      RECT 61.025 -108.965 61.125 -103.985 ;
      RECT 60.785 -109.19 60.885 -108.505 ;
      RECT 60.765 -104.945 60.865 3.135 ;
      RECT 60.335 -104.945 60.435 3.135 ;
      RECT 60.075 -108.685 60.175 -103.985 ;
      RECT 59.95 -101.845 60.05 9.895 ;
      RECT 59.825 -108.965 59.925 -107.215 ;
      RECT 59.565 -108.175 59.665 3.135 ;
      RECT 59.135 -108.175 59.235 3.135 ;
      RECT 59.065 -111.985 59.165 -110.385 ;
      RECT 58.875 -108.685 58.975 -107.215 ;
      RECT 58.75 -101.845 58.85 9.895 ;
      RECT 58.365 -108.175 58.465 3.135 ;
      RECT 57.935 -108.175 58.035 3.135 ;
      RECT 57.675 -113.47 57.775 -107.215 ;
      RECT 57.55 -101.845 57.65 9.895 ;
      RECT 57.425 -108.965 57.525 -103.985 ;
      RECT 57.165 -104.945 57.265 3.135 ;
      RECT 56.735 -104.945 56.835 3.135 ;
      RECT 56.475 -108.685 56.575 -103.985 ;
      RECT 56.35 -101.845 56.45 9.895 ;
      RECT 56.285 -111.985 56.385 -110.37 ;
      RECT 56.225 -108.965 56.325 -103.985 ;
      RECT 55.985 -109.19 56.085 -108.505 ;
      RECT 55.965 -104.945 56.065 3.135 ;
      RECT 55.535 -104.945 55.635 3.135 ;
      RECT 55.275 -108.685 55.375 -103.985 ;
      RECT 55.15 -101.845 55.25 9.895 ;
      RECT 55.025 -108.965 55.125 -107.215 ;
      RECT 54.765 -108.175 54.865 3.135 ;
      RECT 54.335 -108.175 54.435 3.135 ;
      RECT 54.265 -111.985 54.365 -110.385 ;
      RECT 54.075 -108.685 54.175 -107.215 ;
      RECT 53.95 -101.845 54.05 9.895 ;
      RECT 53.565 -108.175 53.665 3.135 ;
      RECT 53.135 -108.175 53.235 3.135 ;
      RECT 52.875 -113.47 52.975 -107.215 ;
      RECT 52.75 -101.845 52.85 9.895 ;
      RECT 52.625 -108.965 52.725 -103.985 ;
      RECT 52.365 -104.945 52.465 3.135 ;
      RECT 51.935 -104.945 52.035 3.135 ;
      RECT 51.675 -108.685 51.775 -103.985 ;
      RECT 51.55 -101.845 51.65 9.895 ;
      RECT 51.485 -111.985 51.585 -110.37 ;
      RECT 51.425 -108.965 51.525 -103.985 ;
      RECT 51.185 -109.19 51.285 -108.505 ;
      RECT 51.165 -104.945 51.265 3.135 ;
      RECT 50.735 -104.945 50.835 3.135 ;
      RECT 50.475 -108.685 50.575 -103.985 ;
      RECT 50.35 -101.845 50.45 9.895 ;
      RECT 50.225 -108.965 50.325 -107.215 ;
      RECT 49.965 -108.175 50.065 3.135 ;
      RECT 49.535 -108.175 49.635 3.135 ;
      RECT 49.465 -111.985 49.565 -110.385 ;
      RECT 49.275 -108.685 49.375 -107.215 ;
      RECT 49.15 -101.845 49.25 9.895 ;
      RECT 48.765 -108.175 48.865 3.135 ;
      RECT 48.335 -108.175 48.435 3.135 ;
      RECT 48.075 -113.47 48.175 -107.215 ;
      RECT 47.95 -101.845 48.05 9.895 ;
      RECT 47.825 -108.965 47.925 -103.985 ;
      RECT 47.565 -104.945 47.665 3.135 ;
      RECT 47.135 -104.945 47.235 3.135 ;
      RECT 46.875 -108.685 46.975 -103.985 ;
      RECT 46.75 -101.845 46.85 9.895 ;
      RECT 46.685 -111.985 46.785 -110.37 ;
      RECT 46.625 -108.965 46.725 -103.985 ;
      RECT 46.385 -109.19 46.485 -108.505 ;
      RECT 46.365 -104.945 46.465 3.135 ;
      RECT 45.935 -104.945 46.035 3.135 ;
      RECT 45.675 -108.685 45.775 -103.985 ;
      RECT 45.55 -101.845 45.65 9.895 ;
      RECT 45.425 -108.965 45.525 -107.215 ;
      RECT 45.165 -108.175 45.265 3.135 ;
      RECT 44.735 -108.175 44.835 3.135 ;
      RECT 44.665 -111.985 44.765 -110.385 ;
      RECT 44.475 -108.685 44.575 -107.215 ;
      RECT 44.35 -101.845 44.45 9.895 ;
      RECT 43.965 -108.175 44.065 3.135 ;
      RECT 43.535 -108.175 43.635 3.135 ;
      RECT 43.275 -113.47 43.375 -107.215 ;
      RECT 43.15 -101.845 43.25 9.895 ;
      RECT 43.025 -108.965 43.125 -103.985 ;
      RECT 42.765 -104.945 42.865 3.135 ;
      RECT 42.335 -104.945 42.435 3.135 ;
      RECT 42.075 -108.685 42.175 -103.985 ;
      RECT 41.95 -101.845 42.05 9.895 ;
      RECT 41.885 -111.985 41.985 -110.37 ;
      RECT 41.825 -108.965 41.925 -103.985 ;
      RECT 41.585 -109.19 41.685 -108.505 ;
      RECT 41.565 -104.945 41.665 3.135 ;
      RECT 41.135 -104.945 41.235 3.135 ;
      RECT 40.875 -108.685 40.975 -103.985 ;
      RECT 40.75 -101.845 40.85 9.895 ;
      RECT 40.625 -108.965 40.725 -107.215 ;
      RECT 40.365 -108.175 40.465 3.135 ;
      RECT 39.935 -108.175 40.035 3.135 ;
      RECT 39.865 -111.985 39.965 -110.385 ;
      RECT 39.675 -108.685 39.775 -107.215 ;
      RECT 39.55 -101.845 39.65 9.895 ;
      RECT 39.165 -108.175 39.265 3.135 ;
      RECT 38.735 -108.175 38.835 3.135 ;
      RECT 38.475 -113.47 38.575 -107.215 ;
      RECT 38.35 -101.845 38.45 9.895 ;
      RECT 38.225 -108.965 38.325 -103.985 ;
      RECT 37.965 -104.945 38.065 3.135 ;
      RECT 37.535 -104.945 37.635 3.135 ;
      RECT 37.275 -108.685 37.375 -103.985 ;
      RECT 37.15 -101.845 37.25 9.895 ;
      RECT 37.085 -111.985 37.185 -110.37 ;
      RECT 37.025 -108.965 37.125 -103.985 ;
      RECT 36.785 -109.19 36.885 -108.505 ;
      RECT 36.765 -104.945 36.865 3.135 ;
      RECT 36.335 -104.945 36.435 3.135 ;
      RECT 36.075 -108.685 36.175 -103.985 ;
      RECT 35.95 -101.845 36.05 9.895 ;
      RECT 35.825 -108.965 35.925 -107.215 ;
      RECT 35.565 -108.175 35.665 3.135 ;
      RECT 35.135 -108.175 35.235 3.135 ;
      RECT 35.065 -111.985 35.165 -110.385 ;
      RECT 34.875 -108.685 34.975 -107.215 ;
      RECT 34.75 -101.845 34.85 9.895 ;
      RECT 34.365 -108.175 34.465 3.135 ;
      RECT 33.935 -108.175 34.035 3.135 ;
      RECT 33.675 -113.47 33.775 -107.215 ;
      RECT 33.55 -101.845 33.65 9.895 ;
      RECT 33.425 -108.965 33.525 -103.985 ;
      RECT 33.165 -104.945 33.265 3.135 ;
      RECT 32.735 -104.945 32.835 3.135 ;
      RECT 32.475 -108.685 32.575 -103.985 ;
      RECT 32.35 -101.845 32.45 9.895 ;
      RECT 32.285 -111.985 32.385 -110.37 ;
      RECT 32.225 -108.965 32.325 -103.985 ;
      RECT 31.985 -109.19 32.085 -108.505 ;
      RECT 31.965 -104.945 32.065 3.135 ;
      RECT 31.535 -104.945 31.635 3.135 ;
      RECT 31.275 -108.685 31.375 -103.985 ;
      RECT 31.15 -101.845 31.25 9.895 ;
      RECT 31.025 -108.965 31.125 -107.215 ;
      RECT 30.765 -108.175 30.865 3.135 ;
      RECT 30.335 -108.175 30.435 3.135 ;
      RECT 30.265 -111.985 30.365 -110.385 ;
      RECT 30.075 -108.685 30.175 -107.215 ;
      RECT 29.95 -101.845 30.05 9.895 ;
      RECT 29.565 -108.175 29.665 3.135 ;
      RECT 29.135 -108.175 29.235 3.135 ;
      RECT 28.875 -113.47 28.975 -107.215 ;
      RECT 28.75 -101.845 28.85 9.895 ;
      RECT 28.625 -108.965 28.725 -103.985 ;
      RECT 28.365 -104.945 28.465 3.135 ;
      RECT 27.935 -104.945 28.035 3.135 ;
      RECT 27.675 -108.685 27.775 -103.985 ;
      RECT 27.55 -101.845 27.65 9.895 ;
      RECT 27.485 -111.985 27.585 -110.37 ;
      RECT 27.425 -108.965 27.525 -103.985 ;
      RECT 27.185 -109.19 27.285 -108.505 ;
      RECT 27.165 -104.945 27.265 3.135 ;
      RECT 26.735 -104.945 26.835 3.135 ;
      RECT 26.475 -108.685 26.575 -103.985 ;
      RECT 26.35 -101.845 26.45 9.895 ;
      RECT 26.225 -108.965 26.325 -107.215 ;
      RECT 25.965 -108.175 26.065 3.135 ;
      RECT 25.535 -108.175 25.635 3.135 ;
      RECT 25.465 -111.985 25.565 -110.385 ;
      RECT 25.275 -108.685 25.375 -107.215 ;
      RECT 25.15 -101.845 25.25 9.895 ;
      RECT 24.765 -108.175 24.865 3.135 ;
      RECT 24.335 -108.175 24.435 3.135 ;
      RECT 24.075 -113.47 24.175 -107.215 ;
      RECT 23.95 -101.845 24.05 9.895 ;
      RECT 23.825 -108.965 23.925 -103.985 ;
      RECT 23.565 -104.945 23.665 3.135 ;
      RECT 23.135 -104.945 23.235 3.135 ;
      RECT 22.875 -108.685 22.975 -103.985 ;
      RECT 22.75 -101.845 22.85 9.895 ;
      RECT 22.685 -111.985 22.785 -110.37 ;
      RECT 22.625 -108.965 22.725 -103.985 ;
      RECT 22.385 -109.19 22.485 -108.505 ;
      RECT 22.365 -104.945 22.465 3.135 ;
      RECT 21.935 -104.945 22.035 3.135 ;
      RECT 21.675 -108.685 21.775 -103.985 ;
      RECT 21.55 -101.845 21.65 9.895 ;
      RECT 21.425 -108.965 21.525 -107.215 ;
      RECT 21.165 -108.175 21.265 3.135 ;
      RECT 20.735 -108.175 20.835 3.135 ;
      RECT 20.665 -111.985 20.765 -110.385 ;
      RECT 20.475 -108.685 20.575 -107.215 ;
      RECT 20.35 -101.845 20.45 9.895 ;
      RECT 19.965 -108.175 20.065 3.135 ;
      RECT 19.535 -108.175 19.635 3.135 ;
      RECT 19.275 -113.47 19.375 -107.215 ;
      RECT 19.15 -101.845 19.25 9.895 ;
      RECT 19.025 -108.965 19.125 -103.985 ;
      RECT 18.765 -104.945 18.865 3.135 ;
      RECT 18.335 -104.945 18.435 3.135 ;
      RECT 18.075 -108.685 18.175 -103.985 ;
      RECT 17.95 -101.845 18.05 9.895 ;
      RECT 17.885 -111.985 17.985 -110.37 ;
      RECT 17.825 -108.965 17.925 -103.985 ;
      RECT 17.585 -109.19 17.685 -108.505 ;
      RECT 17.565 -104.945 17.665 3.135 ;
      RECT 17.135 -104.945 17.235 3.135 ;
      RECT 16.875 -108.685 16.975 -103.985 ;
      RECT 16.75 -101.845 16.85 9.895 ;
      RECT 16.625 -108.965 16.725 -107.215 ;
      RECT 16.365 -108.175 16.465 3.135 ;
      RECT 15.935 -108.175 16.035 3.135 ;
      RECT 15.865 -111.985 15.965 -110.385 ;
      RECT 15.675 -108.685 15.775 -107.215 ;
      RECT 15.55 -101.845 15.65 9.895 ;
      RECT 15.165 -108.175 15.265 3.135 ;
      RECT 14.735 -108.175 14.835 3.135 ;
      RECT 14.475 -113.47 14.575 -107.215 ;
      RECT 14.35 -101.845 14.45 9.895 ;
      RECT 14.225 -108.965 14.325 -103.985 ;
      RECT 13.965 -104.945 14.065 3.135 ;
      RECT 13.535 -104.945 13.635 3.135 ;
      RECT 13.275 -108.685 13.375 -103.985 ;
      RECT 13.15 -101.845 13.25 9.895 ;
      RECT 13.085 -111.985 13.185 -110.37 ;
      RECT 13.025 -108.965 13.125 -103.985 ;
      RECT 12.785 -109.19 12.885 -108.505 ;
      RECT 12.765 -104.945 12.865 3.135 ;
      RECT 12.335 -104.945 12.435 3.135 ;
      RECT 12.075 -108.685 12.175 -103.985 ;
      RECT 11.95 -101.845 12.05 9.895 ;
      RECT 11.825 -108.965 11.925 -107.215 ;
      RECT 11.565 -108.175 11.665 3.135 ;
      RECT 11.135 -108.175 11.235 3.135 ;
      RECT 11.065 -111.985 11.165 -110.385 ;
      RECT 10.875 -108.685 10.975 -107.215 ;
      RECT 10.75 -101.845 10.85 9.895 ;
      RECT 10.365 -108.175 10.465 3.135 ;
      RECT 9.935 -108.175 10.035 3.135 ;
      RECT 9.675 -113.47 9.775 -107.215 ;
      RECT 9.55 -101.845 9.65 9.895 ;
      RECT 9.425 -108.965 9.525 -103.985 ;
      RECT 9.165 -104.945 9.265 3.135 ;
      RECT 8.735 -104.945 8.835 3.135 ;
      RECT 8.475 -108.685 8.575 -103.985 ;
      RECT 8.35 -101.845 8.45 9.895 ;
      RECT 8.285 -111.985 8.385 -110.37 ;
      RECT 8.225 -108.965 8.325 -103.985 ;
      RECT 7.985 -109.19 8.085 -108.505 ;
      RECT 7.965 -104.945 8.065 3.135 ;
      RECT 7.535 -104.945 7.635 3.135 ;
      RECT 7.275 -108.685 7.375 -103.985 ;
      RECT 7.15 -101.845 7.25 9.895 ;
      RECT 7.025 -108.965 7.125 -107.215 ;
      RECT 6.765 -108.175 6.865 3.135 ;
      RECT 6.335 -108.175 6.435 3.135 ;
      RECT 6.265 -111.985 6.365 -110.385 ;
      RECT 6.075 -108.685 6.175 -107.215 ;
      RECT 5.95 -101.845 6.05 9.895 ;
      RECT 5.565 -108.175 5.665 3.135 ;
      RECT 5.135 -108.175 5.235 3.135 ;
      RECT 4.875 -113.47 4.975 -107.215 ;
      RECT 4.75 -101.845 4.85 9.895 ;
      RECT 4.625 -108.965 4.725 -103.985 ;
      RECT 4.365 -104.945 4.465 3.135 ;
      RECT 3.935 -104.945 4.035 3.135 ;
      RECT 3.675 -108.685 3.775 -103.985 ;
      RECT 3.55 -101.845 3.65 9.895 ;
      RECT 3.485 -111.985 3.585 -110.37 ;
      RECT 3.425 -108.965 3.525 -103.985 ;
      RECT 3.185 -109.19 3.285 -108.505 ;
      RECT 3.165 -104.945 3.265 3.135 ;
      RECT 2.735 -104.945 2.835 3.135 ;
      RECT 2.475 -108.685 2.575 -103.985 ;
      RECT 2.35 -101.845 2.45 9.895 ;
      RECT 2.225 -108.965 2.325 -107.215 ;
      RECT 1.965 -108.175 2.065 3.135 ;
      RECT 1.535 -108.175 1.635 3.135 ;
      RECT 1.465 -111.985 1.565 -110.385 ;
      RECT 1.275 -108.685 1.375 -107.215 ;
      RECT 1.15 -101.845 1.25 9.895 ;
      RECT 0.765 -108.175 0.865 3.135 ;
      RECT 0.335 -108.175 0.435 3.135 ;
      RECT 0.075 -113.47 0.175 -107.215 ;
      RECT -0.05 -101.845 0.05 9.895 ;
      RECT -0.565 1.895 -0.465 4.275 ;
      RECT -0.945 -107.655 -0.845 -102.295 ;
      RECT -0.945 -101.195 -0.845 -95.835 ;
      RECT -0.945 -94.735 -0.845 -89.375 ;
      RECT -0.945 -88.275 -0.845 -82.915 ;
      RECT -0.945 -81.815 -0.845 -76.455 ;
      RECT -0.945 -75.355 -0.845 -69.995 ;
      RECT -0.945 -68.895 -0.845 -63.535 ;
      RECT -0.945 -62.435 -0.845 -57.075 ;
      RECT -0.945 -55.975 -0.845 -50.615 ;
      RECT -0.945 -49.515 -0.845 -44.155 ;
      RECT -0.945 -43.055 -0.845 -37.695 ;
      RECT -0.945 -36.595 -0.845 -31.235 ;
      RECT -0.945 -30.135 -0.845 -24.775 ;
      RECT -0.945 -23.675 -0.845 -18.315 ;
      RECT -0.945 -17.215 -0.845 -11.855 ;
      RECT -0.945 -10.755 -0.845 -5.395 ;
      RECT -0.945 -4.295 -0.845 1.065 ;
      RECT -1.465 -107.655 -1.365 -102.295 ;
      RECT -1.465 -101.195 -1.365 -95.835 ;
      RECT -1.465 -94.735 -1.365 -89.375 ;
      RECT -1.465 -88.275 -1.365 -82.915 ;
      RECT -1.465 -81.815 -1.365 -76.455 ;
      RECT -1.465 -75.355 -1.365 -69.995 ;
      RECT -1.465 -68.895 -1.365 -63.535 ;
      RECT -1.465 -62.435 -1.365 -57.075 ;
      RECT -1.465 -55.975 -1.365 -50.615 ;
      RECT -1.465 -49.515 -1.365 -44.155 ;
      RECT -1.465 -43.055 -1.365 -37.695 ;
      RECT -1.465 -36.595 -1.365 -31.235 ;
      RECT -1.465 -30.135 -1.365 -24.775 ;
      RECT -1.465 -23.675 -1.365 -18.315 ;
      RECT -1.465 -17.215 -1.365 -11.855 ;
      RECT -1.465 -10.755 -1.365 -5.395 ;
      RECT -1.465 -4.295 -1.365 1.065 ;
      RECT -1.985 -107.655 -1.885 -107.055 ;
      RECT -1.985 -103.45 -1.885 -102.295 ;
      RECT -1.985 -101.195 -1.885 -100.04 ;
      RECT -1.985 -96.435 -1.885 -95.835 ;
      RECT -1.985 -94.735 -1.885 -94.135 ;
      RECT -1.985 -90.53 -1.885 -89.375 ;
      RECT -1.985 -88.275 -1.885 -87.12 ;
      RECT -1.985 -83.515 -1.885 -82.915 ;
      RECT -1.985 -81.815 -1.885 -81.215 ;
      RECT -1.985 -77.61 -1.885 -76.455 ;
      RECT -1.985 -75.355 -1.885 -74.2 ;
      RECT -1.985 -70.595 -1.885 -69.995 ;
      RECT -1.985 -68.895 -1.885 -68.295 ;
      RECT -1.985 -64.69 -1.885 -63.535 ;
      RECT -1.985 -62.435 -1.885 -61.28 ;
      RECT -1.985 -57.675 -1.885 -57.075 ;
      RECT -1.985 -55.975 -1.885 -55.375 ;
      RECT -1.985 -51.77 -1.885 -50.615 ;
      RECT -1.985 -49.515 -1.885 -48.36 ;
      RECT -1.985 -44.755 -1.885 -44.155 ;
      RECT -1.985 -43.055 -1.885 -42.455 ;
      RECT -1.985 -38.85 -1.885 -37.695 ;
      RECT -1.985 -36.595 -1.885 -35.44 ;
      RECT -1.985 -31.835 -1.885 -31.235 ;
      RECT -1.985 -30.135 -1.885 -29.535 ;
      RECT -1.985 -25.93 -1.885 -24.775 ;
      RECT -1.985 -23.675 -1.885 -22.52 ;
      RECT -1.985 -18.915 -1.885 -18.315 ;
      RECT -1.985 -17.215 -1.885 -16.615 ;
      RECT -1.985 -13.01 -1.885 -11.855 ;
      RECT -1.985 -10.755 -1.885 -9.6 ;
      RECT -1.985 -5.995 -1.885 -5.395 ;
      RECT -1.985 -4.295 -1.885 -3.695 ;
      RECT -1.985 -0.09 -1.885 1.065 ;
      RECT -2.245 -107.655 -2.145 -102.295 ;
      RECT -2.245 -101.195 -2.145 -95.835 ;
      RECT -2.245 -94.735 -2.145 -89.375 ;
      RECT -2.245 -88.275 -2.145 -82.915 ;
      RECT -2.245 -81.815 -2.145 -76.455 ;
      RECT -2.245 -75.355 -2.145 -69.995 ;
      RECT -2.245 -68.895 -2.145 -63.535 ;
      RECT -2.245 -62.435 -2.145 -57.075 ;
      RECT -2.245 -55.975 -2.145 -50.615 ;
      RECT -2.245 -49.515 -2.145 -44.155 ;
      RECT -2.245 -43.055 -2.145 -37.695 ;
      RECT -2.245 -36.595 -2.145 -31.235 ;
      RECT -2.245 -30.135 -2.145 -24.775 ;
      RECT -2.245 -23.675 -2.145 -18.315 ;
      RECT -2.245 -17.215 -2.145 -11.855 ;
      RECT -2.245 -10.755 -2.145 -5.395 ;
      RECT -2.245 -4.295 -2.145 1.065 ;
      RECT -2.765 -107.655 -2.665 -102.295 ;
      RECT -2.765 -101.195 -2.665 -95.835 ;
      RECT -2.765 -94.735 -2.665 -89.375 ;
      RECT -2.765 -88.275 -2.665 -82.915 ;
      RECT -2.765 -81.815 -2.665 -76.455 ;
      RECT -2.765 -75.355 -2.665 -69.995 ;
      RECT -2.765 -68.895 -2.665 -63.535 ;
      RECT -2.765 -62.435 -2.665 -57.075 ;
      RECT -2.765 -55.975 -2.665 -50.615 ;
      RECT -2.765 -49.515 -2.665 -44.155 ;
      RECT -2.765 -43.055 -2.665 -37.695 ;
      RECT -2.765 -36.595 -2.665 -31.235 ;
      RECT -2.765 -30.135 -2.665 -24.775 ;
      RECT -2.765 -23.675 -2.665 -18.315 ;
      RECT -2.765 -17.215 -2.665 -11.855 ;
      RECT -2.765 -10.755 -2.665 -5.395 ;
      RECT -2.765 -4.295 -2.665 1.065 ;
      RECT -3.285 -107.655 -3.185 -107.055 ;
      RECT -3.285 -103.45 -3.185 -102.295 ;
      RECT -3.285 -101.195 -3.185 -100.04 ;
      RECT -3.285 -96.435 -3.185 -95.835 ;
      RECT -3.285 -94.735 -3.185 -94.135 ;
      RECT -3.285 -90.53 -3.185 -89.375 ;
      RECT -3.285 -88.275 -3.185 -87.12 ;
      RECT -3.285 -83.515 -3.185 -82.915 ;
      RECT -3.285 -81.815 -3.185 -81.215 ;
      RECT -3.285 -77.61 -3.185 -76.455 ;
      RECT -3.285 -75.355 -3.185 -74.2 ;
      RECT -3.285 -70.595 -3.185 -69.995 ;
      RECT -3.285 -68.895 -3.185 -68.295 ;
      RECT -3.285 -64.69 -3.185 -63.535 ;
      RECT -3.285 -62.435 -3.185 -61.28 ;
      RECT -3.285 -57.675 -3.185 -57.075 ;
      RECT -3.285 -55.975 -3.185 -55.375 ;
      RECT -3.285 -51.77 -3.185 -50.615 ;
      RECT -3.285 -49.515 -3.185 -48.36 ;
      RECT -3.285 -44.755 -3.185 -44.155 ;
      RECT -3.285 -43.055 -3.185 -42.455 ;
      RECT -3.285 -38.85 -3.185 -37.695 ;
      RECT -3.285 -36.595 -3.185 -35.44 ;
      RECT -3.285 -31.835 -3.185 -31.235 ;
      RECT -3.285 -30.135 -3.185 -29.535 ;
      RECT -3.285 -25.93 -3.185 -24.775 ;
      RECT -3.285 -23.675 -3.185 -22.52 ;
      RECT -3.285 -18.915 -3.185 -18.315 ;
      RECT -3.285 -17.215 -3.185 -16.615 ;
      RECT -3.285 -13.01 -3.185 -11.855 ;
      RECT -3.285 -10.755 -3.185 -9.6 ;
      RECT -3.285 -5.995 -3.185 -5.395 ;
      RECT -3.285 -4.295 -3.185 -3.695 ;
      RECT -3.285 -0.09 -3.185 1.065 ;
      RECT -3.545 -107.655 -3.445 -102.295 ;
      RECT -3.545 -101.195 -3.445 -95.835 ;
      RECT -3.545 -94.735 -3.445 -89.375 ;
      RECT -3.545 -88.275 -3.445 -82.915 ;
      RECT -3.545 -81.815 -3.445 -76.455 ;
      RECT -3.545 -75.355 -3.445 -69.995 ;
      RECT -3.545 -68.895 -3.445 -63.535 ;
      RECT -3.545 -62.435 -3.445 -57.075 ;
      RECT -3.545 -55.975 -3.445 -50.615 ;
      RECT -3.545 -49.515 -3.445 -44.155 ;
      RECT -3.545 -43.055 -3.445 -37.695 ;
      RECT -3.545 -36.595 -3.445 -31.235 ;
      RECT -3.545 -30.135 -3.445 -24.775 ;
      RECT -3.545 -23.675 -3.445 -18.315 ;
      RECT -3.545 -17.215 -3.445 -11.855 ;
      RECT -3.545 -10.755 -3.445 -5.395 ;
      RECT -3.545 -4.295 -3.445 1.065 ;
      RECT -4.065 -107.655 -3.965 -102.295 ;
      RECT -4.065 -101.195 -3.965 -95.835 ;
      RECT -4.065 -94.735 -3.965 -89.375 ;
      RECT -4.065 -88.275 -3.965 -82.915 ;
      RECT -4.065 -81.815 -3.965 -76.455 ;
      RECT -4.065 -75.355 -3.965 -69.995 ;
      RECT -4.065 -68.895 -3.965 -63.535 ;
      RECT -4.065 -62.435 -3.965 -57.075 ;
      RECT -4.065 -55.975 -3.965 -50.615 ;
      RECT -4.065 -49.515 -3.965 -44.155 ;
      RECT -4.065 -43.055 -3.965 -37.695 ;
      RECT -4.065 -36.595 -3.965 -31.235 ;
      RECT -4.065 -30.135 -3.965 -24.775 ;
      RECT -4.065 -23.675 -3.965 -18.315 ;
      RECT -4.065 -17.215 -3.965 -11.855 ;
      RECT -4.065 -10.755 -3.965 -5.395 ;
      RECT -4.065 -4.295 -3.965 1.065 ;
      RECT -4.585 -107.655 -4.485 -107.055 ;
      RECT -4.585 -103.45 -4.485 -102.295 ;
      RECT -4.585 -101.195 -4.485 -100.04 ;
      RECT -4.585 -96.435 -4.485 -95.835 ;
      RECT -4.585 -94.735 -4.485 -94.135 ;
      RECT -4.585 -90.53 -4.485 -89.375 ;
      RECT -4.585 -88.275 -4.485 -87.12 ;
      RECT -4.585 -83.515 -4.485 -82.915 ;
      RECT -4.585 -81.815 -4.485 -81.215 ;
      RECT -4.585 -77.61 -4.485 -76.455 ;
      RECT -4.585 -75.355 -4.485 -74.2 ;
      RECT -4.585 -70.595 -4.485 -69.995 ;
      RECT -4.585 -68.895 -4.485 -68.295 ;
      RECT -4.585 -64.69 -4.485 -63.535 ;
      RECT -4.585 -62.435 -4.485 -61.28 ;
      RECT -4.585 -57.675 -4.485 -57.075 ;
      RECT -4.585 -55.975 -4.485 -55.375 ;
      RECT -4.585 -51.77 -4.485 -50.615 ;
      RECT -4.585 -49.515 -4.485 -48.36 ;
      RECT -4.585 -44.755 -4.485 -44.155 ;
      RECT -4.585 -43.055 -4.485 -42.455 ;
      RECT -4.585 -38.85 -4.485 -37.695 ;
      RECT -4.585 -36.595 -4.485 -35.44 ;
      RECT -4.585 -31.835 -4.485 -31.235 ;
      RECT -4.585 -30.135 -4.485 -29.535 ;
      RECT -4.585 -25.93 -4.485 -24.775 ;
      RECT -4.585 -23.675 -4.485 -22.52 ;
      RECT -4.585 -18.915 -4.485 -18.315 ;
      RECT -4.585 -17.215 -4.485 -16.615 ;
      RECT -4.585 -13.01 -4.485 -11.855 ;
      RECT -4.585 -10.755 -4.485 -9.6 ;
      RECT -4.585 -5.995 -4.485 -5.395 ;
      RECT -4.585 -4.295 -4.485 -3.695 ;
      RECT -4.585 -0.09 -4.485 1.065 ;
      RECT -4.845 -107.655 -4.745 -102.295 ;
      RECT -4.845 -101.195 -4.745 -95.835 ;
      RECT -4.845 -94.735 -4.745 -89.375 ;
      RECT -4.845 -88.275 -4.745 -82.915 ;
      RECT -4.845 -81.815 -4.745 -76.455 ;
      RECT -4.845 -75.355 -4.745 -69.995 ;
      RECT -4.845 -68.895 -4.745 -63.535 ;
      RECT -4.845 -62.435 -4.745 -57.075 ;
      RECT -4.845 -55.975 -4.745 -50.615 ;
      RECT -4.845 -49.515 -4.745 -44.155 ;
      RECT -4.845 -43.055 -4.745 -37.695 ;
      RECT -4.845 -36.595 -4.745 -31.235 ;
      RECT -4.845 -30.135 -4.745 -24.775 ;
      RECT -4.845 -23.675 -4.745 -18.315 ;
      RECT -4.845 -17.215 -4.745 -11.855 ;
      RECT -4.845 -10.755 -4.745 -5.395 ;
      RECT -4.845 -4.295 -4.745 1.065 ;
      RECT -5.105 -111.215 -5.005 4.275 ;
      RECT -5.365 -107.655 -5.265 -102.295 ;
      RECT -5.365 -101.195 -5.265 -95.835 ;
      RECT -5.365 -94.735 -5.265 -89.375 ;
      RECT -5.365 -88.275 -5.265 -82.915 ;
      RECT -5.365 -81.815 -5.265 -76.455 ;
      RECT -5.365 -75.355 -5.265 -69.995 ;
      RECT -5.365 -68.895 -5.265 -63.535 ;
      RECT -5.365 -62.435 -5.265 -57.075 ;
      RECT -5.365 -55.975 -5.265 -50.615 ;
      RECT -5.365 -49.515 -5.265 -44.155 ;
      RECT -5.365 -43.055 -5.265 -37.695 ;
      RECT -5.365 -36.595 -5.265 -31.235 ;
      RECT -5.365 -30.135 -5.265 -24.775 ;
      RECT -5.365 -23.675 -5.265 -18.315 ;
      RECT -5.365 -17.215 -5.265 -11.855 ;
      RECT -5.365 -10.755 -5.265 -5.395 ;
      RECT -5.365 -4.295 -5.265 1.065 ;
      RECT -5.885 -107.655 -5.785 -107.055 ;
      RECT -5.885 -103.45 -5.785 -102.295 ;
      RECT -5.885 -101.195 -5.785 -100.04 ;
      RECT -5.885 -96.435 -5.785 -95.835 ;
      RECT -5.885 -94.735 -5.785 -94.135 ;
      RECT -5.885 -90.53 -5.785 -89.375 ;
      RECT -5.885 -88.275 -5.785 -87.12 ;
      RECT -5.885 -83.515 -5.785 -82.915 ;
      RECT -5.885 -81.815 -5.785 -81.215 ;
      RECT -5.885 -77.61 -5.785 -76.455 ;
      RECT -5.885 -75.355 -5.785 -74.2 ;
      RECT -5.885 -70.595 -5.785 -69.995 ;
      RECT -5.885 -68.895 -5.785 -68.295 ;
      RECT -5.885 -64.69 -5.785 -63.535 ;
      RECT -5.885 -62.435 -5.785 -61.28 ;
      RECT -5.885 -57.675 -5.785 -57.075 ;
      RECT -5.885 -55.975 -5.785 -55.375 ;
      RECT -5.885 -51.77 -5.785 -50.615 ;
      RECT -5.885 -49.515 -5.785 -48.36 ;
      RECT -5.885 -44.755 -5.785 -44.155 ;
      RECT -5.885 -43.055 -5.785 -42.455 ;
      RECT -5.885 -38.85 -5.785 -37.695 ;
      RECT -5.885 -36.595 -5.785 -35.44 ;
      RECT -5.885 -31.835 -5.785 -31.235 ;
      RECT -5.885 -30.135 -5.785 -29.535 ;
      RECT -5.885 -25.93 -5.785 -24.775 ;
      RECT -5.885 -23.675 -5.785 -22.52 ;
      RECT -5.885 -18.915 -5.785 -18.315 ;
      RECT -5.885 -17.215 -5.785 -16.615 ;
      RECT -5.885 -13.01 -5.785 -11.855 ;
      RECT -5.885 -10.755 -5.785 -9.6 ;
      RECT -5.885 -5.995 -5.785 -5.395 ;
      RECT -5.885 -4.295 -5.785 -3.695 ;
      RECT -5.885 -0.09 -5.785 1.065 ;
      RECT -6.145 -107.655 -6.045 -102.295 ;
      RECT -6.145 -101.195 -6.045 -95.835 ;
      RECT -6.145 -94.735 -6.045 -89.375 ;
      RECT -6.145 -88.275 -6.045 -82.915 ;
      RECT -6.145 -81.815 -6.045 -76.455 ;
      RECT -6.145 -75.355 -6.045 -69.995 ;
      RECT -6.145 -68.895 -6.045 -63.535 ;
      RECT -6.145 -62.435 -6.045 -57.075 ;
      RECT -6.145 -55.975 -6.045 -50.615 ;
      RECT -6.145 -49.515 -6.045 -44.155 ;
      RECT -6.145 -43.055 -6.045 -37.695 ;
      RECT -6.145 -36.595 -6.045 -31.235 ;
      RECT -6.145 -30.135 -6.045 -24.775 ;
      RECT -6.145 -23.675 -6.045 -18.315 ;
      RECT -6.145 -17.215 -6.045 -11.855 ;
      RECT -6.145 -10.755 -6.045 -5.395 ;
      RECT -6.145 -4.295 -6.045 1.065 ;
      RECT -6.665 -107.655 -6.565 -102.295 ;
      RECT -6.665 -101.195 -6.565 -95.835 ;
      RECT -6.665 -94.735 -6.565 -89.375 ;
      RECT -6.665 -88.275 -6.565 -82.915 ;
      RECT -6.665 -81.815 -6.565 -76.455 ;
      RECT -6.665 -75.355 -6.565 -69.995 ;
      RECT -6.665 -68.895 -6.565 -63.535 ;
      RECT -6.665 -62.435 -6.565 -57.075 ;
      RECT -6.665 -55.975 -6.565 -50.615 ;
      RECT -6.665 -49.515 -6.565 -44.155 ;
      RECT -6.665 -43.055 -6.565 -37.695 ;
      RECT -6.665 -36.595 -6.565 -31.235 ;
      RECT -6.665 -30.135 -6.565 -24.775 ;
      RECT -6.665 -23.675 -6.565 -18.315 ;
      RECT -6.665 -17.215 -6.565 -11.855 ;
      RECT -6.665 -10.755 -6.565 -5.395 ;
      RECT -6.665 -4.295 -6.565 1.065 ;
      RECT -7.445 -107.655 -7.345 -102.295 ;
      RECT -7.445 -101.195 -7.345 -95.835 ;
      RECT -7.445 -94.735 -7.345 -89.375 ;
      RECT -7.445 -88.275 -7.345 -82.915 ;
      RECT -7.445 -81.815 -7.345 -76.455 ;
      RECT -7.445 -75.355 -7.345 -69.995 ;
      RECT -7.445 -68.895 -7.345 -63.535 ;
      RECT -7.445 -62.435 -7.345 -57.075 ;
      RECT -7.445 -55.975 -7.345 -50.615 ;
      RECT -7.445 -49.515 -7.345 -44.155 ;
      RECT -7.445 -43.055 -7.345 -37.695 ;
      RECT -7.445 -36.595 -7.345 -31.235 ;
      RECT -7.445 -30.135 -7.345 -24.775 ;
      RECT -7.445 -23.675 -7.345 -18.315 ;
      RECT -7.445 -17.215 -7.345 -11.855 ;
      RECT -7.445 -10.755 -7.345 -5.395 ;
      RECT -7.445 -4.295 -7.345 1.065 ;
      RECT -7.965 -107.655 -7.865 -102.295 ;
      RECT -7.965 -101.195 -7.865 -95.835 ;
      RECT -7.965 -94.735 -7.865 -89.375 ;
      RECT -7.965 -88.275 -7.865 -82.915 ;
      RECT -7.965 -81.815 -7.865 -76.455 ;
      RECT -7.965 -75.355 -7.865 -69.995 ;
      RECT -7.965 -68.895 -7.865 -63.535 ;
      RECT -7.965 -62.435 -7.865 -57.075 ;
      RECT -7.965 -55.975 -7.865 -50.615 ;
      RECT -7.965 -49.515 -7.865 -44.155 ;
      RECT -7.965 -43.055 -7.865 -37.695 ;
      RECT -7.965 -36.595 -7.865 -31.235 ;
      RECT -7.965 -30.135 -7.865 -24.775 ;
      RECT -7.965 -23.675 -7.865 -18.315 ;
      RECT -7.965 -17.215 -7.865 -11.855 ;
      RECT -7.965 -10.755 -7.865 -5.395 ;
      RECT -7.965 -4.295 -7.865 1.065 ;
      RECT -8.745 -107.655 -8.645 -102.295 ;
      RECT -8.745 -101.195 -8.645 -95.835 ;
      RECT -8.745 -94.735 -8.645 -89.375 ;
      RECT -8.745 -88.275 -8.645 -82.915 ;
      RECT -8.745 -81.815 -8.645 -76.455 ;
      RECT -8.745 -75.355 -8.645 -69.995 ;
      RECT -8.745 -68.895 -8.645 -63.535 ;
      RECT -8.745 -62.435 -8.645 -57.075 ;
      RECT -8.745 -55.975 -8.645 -50.615 ;
      RECT -8.745 -49.515 -8.645 -44.155 ;
      RECT -8.745 -43.055 -8.645 -37.695 ;
      RECT -8.745 -36.595 -8.645 -31.235 ;
      RECT -8.745 -30.135 -8.645 -24.775 ;
      RECT -8.745 -23.675 -8.645 -18.315 ;
      RECT -8.745 -17.215 -8.645 -11.855 ;
      RECT -8.745 -10.755 -8.645 -5.395 ;
      RECT -8.745 -4.295 -8.645 1.065 ;
      RECT -9.265 -107.655 -9.165 -102.295 ;
      RECT -9.265 -101.195 -9.165 -95.835 ;
      RECT -9.265 -94.735 -9.165 -89.375 ;
      RECT -9.265 -88.275 -9.165 -82.915 ;
      RECT -9.265 -81.815 -9.165 -76.455 ;
      RECT -9.265 -75.355 -9.165 -69.995 ;
      RECT -9.265 -68.895 -9.165 -63.535 ;
      RECT -9.265 -62.435 -9.165 -57.075 ;
      RECT -9.265 -55.975 -9.165 -50.615 ;
      RECT -9.265 -49.515 -9.165 -44.155 ;
      RECT -9.265 -43.055 -9.165 -37.695 ;
      RECT -9.265 -36.595 -9.165 -31.235 ;
      RECT -9.265 -30.135 -9.165 -24.775 ;
      RECT -9.265 -23.675 -9.165 -18.315 ;
      RECT -9.265 -17.215 -9.165 -11.855 ;
      RECT -9.265 -10.755 -9.165 -5.395 ;
      RECT -9.265 -4.295 -9.165 1.065 ;
      RECT -10.045 -107.655 -9.945 -102.295 ;
      RECT -10.045 -101.195 -9.945 -95.835 ;
      RECT -10.045 -94.735 -9.945 -89.375 ;
      RECT -10.045 -88.275 -9.945 -82.915 ;
      RECT -10.045 -81.815 -9.945 -76.455 ;
      RECT -10.045 -75.355 -9.945 -69.995 ;
      RECT -10.045 -68.895 -9.945 -63.535 ;
      RECT -10.045 -62.435 -9.945 -57.075 ;
      RECT -10.045 -55.975 -9.945 -50.615 ;
      RECT -10.045 -49.515 -9.945 -44.155 ;
      RECT -10.045 -43.055 -9.945 -37.695 ;
      RECT -10.045 -36.595 -9.945 -31.235 ;
      RECT -10.045 -30.135 -9.945 -24.775 ;
      RECT -10.045 -23.675 -9.945 -18.315 ;
      RECT -10.045 -17.215 -9.945 -11.855 ;
      RECT -10.045 -10.755 -9.945 -5.395 ;
      RECT -10.045 -4.295 -9.945 1.065 ;
      RECT -10.565 -107.655 -10.465 -102.295 ;
      RECT -10.565 -101.195 -10.465 -95.835 ;
      RECT -10.565 -94.735 -10.465 -89.375 ;
      RECT -10.565 -88.275 -10.465 -82.915 ;
      RECT -10.565 -81.815 -10.465 -76.455 ;
      RECT -10.565 -75.355 -10.465 -69.995 ;
      RECT -10.565 -68.895 -10.465 -63.535 ;
      RECT -10.565 -62.435 -10.465 -57.075 ;
      RECT -10.565 -55.975 -10.465 -50.615 ;
      RECT -10.565 -49.515 -10.465 -44.155 ;
      RECT -10.565 -43.055 -10.465 -37.695 ;
      RECT -10.565 -36.595 -10.465 -31.235 ;
      RECT -10.565 -30.135 -10.465 -24.775 ;
      RECT -10.565 -23.675 -10.465 -18.315 ;
      RECT -10.565 -17.215 -10.465 -11.855 ;
      RECT -10.565 -10.755 -10.465 -5.395 ;
      RECT -10.565 -4.295 -10.465 1.065 ;
      RECT -11.345 -101.195 -11.245 -95.835 ;
      RECT -11.345 -94.735 -11.245 -89.375 ;
      RECT -11.345 -88.275 -11.245 -82.915 ;
      RECT -11.345 -81.815 -11.245 -76.455 ;
      RECT -11.345 -75.355 -11.245 -69.995 ;
      RECT -11.345 -68.895 -11.245 -63.535 ;
      RECT -11.345 -62.435 -11.245 -57.075 ;
      RECT -11.345 -55.975 -11.245 -50.615 ;
      RECT -11.345 -49.515 -11.245 -44.155 ;
      RECT -11.345 -43.055 -11.245 -37.695 ;
      RECT -11.345 -36.595 -11.245 -31.235 ;
      RECT -11.345 -30.135 -11.245 -24.775 ;
      RECT -11.345 -23.675 -11.245 -18.315 ;
      RECT -11.345 -17.215 -11.245 -11.855 ;
      RECT -11.345 -10.755 -11.245 -5.395 ;
      RECT -11.345 -4.295 -11.245 1.065 ;
      RECT -11.865 -101.195 -11.765 -95.835 ;
      RECT -11.865 -94.735 -11.765 -89.375 ;
      RECT -11.865 -88.275 -11.765 -82.915 ;
      RECT -11.865 -81.815 -11.765 -76.455 ;
      RECT -11.865 -75.355 -11.765 -69.995 ;
      RECT -11.865 -68.895 -11.765 -63.535 ;
      RECT -11.865 -62.435 -11.765 -57.075 ;
      RECT -11.865 -55.975 -11.765 -50.615 ;
      RECT -11.865 -49.515 -11.765 -44.155 ;
      RECT -11.865 -43.055 -11.765 -37.695 ;
      RECT -11.865 -36.595 -11.765 -31.235 ;
      RECT -11.865 -30.135 -11.765 -24.775 ;
      RECT -11.865 -23.675 -11.765 -18.315 ;
      RECT -11.865 -17.215 -11.765 -11.855 ;
      RECT -11.865 -10.755 -11.765 -5.395 ;
      RECT -11.865 -4.295 -11.765 1.065 ;
      RECT -12.645 -101.195 -12.545 -95.835 ;
      RECT -12.645 -94.735 -12.545 -89.375 ;
      RECT -12.645 -88.275 -12.545 -82.915 ;
      RECT -12.645 -81.815 -12.545 -76.455 ;
      RECT -12.645 -75.355 -12.545 -69.995 ;
      RECT -12.645 -68.895 -12.545 -63.535 ;
      RECT -12.645 -62.435 -12.545 -57.075 ;
      RECT -12.645 -55.975 -12.545 -50.615 ;
      RECT -12.645 -49.515 -12.545 -44.155 ;
      RECT -12.645 -43.055 -12.545 -37.695 ;
      RECT -12.645 -36.595 -12.545 -31.235 ;
      RECT -12.645 -30.135 -12.545 -24.775 ;
      RECT -12.645 -23.675 -12.545 -18.315 ;
      RECT -12.645 -17.215 -12.545 -11.855 ;
      RECT -12.645 -10.755 -12.545 -5.395 ;
      RECT -12.645 -4.295 -12.545 1.065 ;
      RECT -13.165 -101.195 -13.065 -95.835 ;
      RECT -13.165 -94.735 -13.065 -89.375 ;
      RECT -13.165 -88.275 -13.065 -82.915 ;
      RECT -13.165 -81.815 -13.065 -76.455 ;
      RECT -13.165 -75.355 -13.065 -69.995 ;
      RECT -13.165 -68.895 -13.065 -63.535 ;
      RECT -13.165 -62.435 -13.065 -57.075 ;
      RECT -13.165 -55.975 -13.065 -50.615 ;
      RECT -13.165 -49.515 -13.065 -44.155 ;
      RECT -13.165 -43.055 -13.065 -37.695 ;
      RECT -13.165 -36.595 -13.065 -31.235 ;
      RECT -13.165 -30.135 -13.065 -24.775 ;
      RECT -13.165 -23.675 -13.065 -18.315 ;
      RECT -13.165 -17.215 -13.065 -11.855 ;
      RECT -13.165 -10.755 -13.065 -5.395 ;
      RECT -13.165 -4.295 -13.065 1.065 ;
      RECT -13.945 -101.195 -13.845 -95.835 ;
      RECT -13.945 -94.735 -13.845 -89.375 ;
      RECT -13.945 -88.275 -13.845 -82.915 ;
      RECT -13.945 -81.815 -13.845 -76.455 ;
      RECT -13.945 -75.355 -13.845 -69.995 ;
      RECT -13.945 -68.895 -13.845 -63.535 ;
      RECT -13.945 -62.435 -13.845 -57.075 ;
      RECT -13.945 -55.975 -13.845 -50.615 ;
      RECT -13.945 -49.515 -13.845 -44.155 ;
      RECT -13.945 -43.055 -13.845 -37.695 ;
      RECT -13.945 -36.595 -13.845 -31.235 ;
      RECT -13.945 -30.135 -13.845 -24.775 ;
      RECT -13.945 -23.675 -13.845 -18.315 ;
      RECT -13.945 -17.215 -13.845 -11.855 ;
      RECT -13.945 -10.755 -13.845 -5.395 ;
      RECT -13.945 -4.295 -13.845 1.065 ;
      RECT -14.465 -101.195 -14.365 -95.835 ;
      RECT -14.465 -94.735 -14.365 -89.375 ;
      RECT -14.465 -88.275 -14.365 -82.915 ;
      RECT -14.465 -81.815 -14.365 -76.455 ;
      RECT -14.465 -75.355 -14.365 -69.995 ;
      RECT -14.465 -68.895 -14.365 -63.535 ;
      RECT -14.465 -62.435 -14.365 -57.075 ;
      RECT -14.465 -55.975 -14.365 -50.615 ;
      RECT -14.465 -49.515 -14.365 -44.155 ;
      RECT -14.465 -43.055 -14.365 -37.695 ;
      RECT -14.465 -36.595 -14.365 -31.235 ;
      RECT -14.465 -30.135 -14.365 -24.775 ;
      RECT -14.465 -23.675 -14.365 -18.315 ;
      RECT -14.465 -17.215 -14.365 -11.855 ;
      RECT -14.465 -10.755 -14.365 -5.395 ;
      RECT -14.465 -4.295 -14.365 1.065 ;
      RECT -15.245 -101.195 -15.145 -95.835 ;
      RECT -15.245 -94.735 -15.145 -89.375 ;
      RECT -15.245 -88.275 -15.145 -82.915 ;
      RECT -15.245 -81.815 -15.145 -76.455 ;
      RECT -15.245 -75.355 -15.145 -69.995 ;
      RECT -15.245 -68.895 -15.145 -63.535 ;
      RECT -15.245 -62.435 -15.145 -57.075 ;
      RECT -15.245 -55.975 -15.145 -50.615 ;
      RECT -15.245 -49.515 -15.145 -44.155 ;
      RECT -15.245 -43.055 -15.145 -37.695 ;
      RECT -15.245 -36.595 -15.145 -31.235 ;
      RECT -15.245 -30.135 -15.145 -24.775 ;
      RECT -15.245 -23.675 -15.145 -18.315 ;
      RECT -15.245 -17.215 -15.145 -11.855 ;
      RECT -15.245 -10.755 -15.145 -5.395 ;
      RECT -15.245 -4.295 -15.145 1.065 ;
      RECT -15.765 -101.195 -15.665 -95.835 ;
      RECT -15.765 -94.735 -15.665 -89.375 ;
      RECT -15.765 -88.275 -15.665 -82.915 ;
      RECT -15.765 -81.815 -15.665 -76.455 ;
      RECT -15.765 -75.355 -15.665 -69.995 ;
      RECT -15.765 -68.895 -15.665 -63.535 ;
      RECT -15.765 -62.435 -15.665 -57.075 ;
      RECT -15.765 -55.975 -15.665 -50.615 ;
      RECT -15.765 -49.515 -15.665 -44.155 ;
      RECT -15.765 -43.055 -15.665 -37.695 ;
      RECT -15.765 -36.595 -15.665 -31.235 ;
      RECT -15.765 -30.135 -15.665 -24.775 ;
      RECT -15.765 -23.675 -15.665 -18.315 ;
      RECT -15.765 -17.215 -15.665 -11.855 ;
      RECT -15.765 -10.755 -15.665 -5.395 ;
      RECT -15.765 -4.295 -15.665 1.065 ;
      RECT -16.545 -101.195 -16.445 -95.835 ;
      RECT -16.545 -94.735 -16.445 -89.375 ;
      RECT -16.545 -88.275 -16.445 -82.915 ;
      RECT -16.545 -81.815 -16.445 -76.455 ;
      RECT -16.545 -75.355 -16.445 -69.995 ;
      RECT -16.545 -68.895 -16.445 -63.535 ;
      RECT -16.545 -62.435 -16.445 -57.075 ;
      RECT -16.545 -55.975 -16.445 -50.615 ;
      RECT -16.545 -49.515 -16.445 -44.155 ;
      RECT -16.545 -43.055 -16.445 -37.695 ;
      RECT -16.545 -36.595 -16.445 -31.235 ;
      RECT -16.545 -30.135 -16.445 -24.775 ;
      RECT -16.545 -23.675 -16.445 -18.315 ;
      RECT -16.545 -17.215 -16.445 -11.855 ;
      RECT -16.545 -10.755 -16.445 -5.395 ;
      RECT -16.545 -4.295 -16.445 1.065 ;
      RECT -17.065 -101.195 -16.965 -95.835 ;
      RECT -17.065 -94.735 -16.965 -89.375 ;
      RECT -17.065 -88.275 -16.965 -82.915 ;
      RECT -17.065 -81.815 -16.965 -76.455 ;
      RECT -17.065 -75.355 -16.965 -69.995 ;
      RECT -17.065 -68.895 -16.965 -63.535 ;
      RECT -17.065 -62.435 -16.965 -57.075 ;
      RECT -17.065 -55.975 -16.965 -50.615 ;
      RECT -17.065 -49.515 -16.965 -44.155 ;
      RECT -17.065 -43.055 -16.965 -37.695 ;
      RECT -17.065 -36.595 -16.965 -31.235 ;
      RECT -17.065 -30.135 -16.965 -24.775 ;
      RECT -17.065 -23.675 -16.965 -18.315 ;
      RECT -17.065 -17.215 -16.965 -11.855 ;
      RECT -17.065 -10.755 -16.965 -5.395 ;
      RECT -17.065 -4.295 -16.965 1.065 ;
      RECT -17.845 -101.195 -17.745 -95.835 ;
      RECT -17.845 -94.735 -17.745 -89.375 ;
      RECT -17.845 -88.275 -17.745 -82.915 ;
      RECT -17.845 -81.815 -17.745 -76.455 ;
      RECT -17.845 -75.355 -17.745 -69.995 ;
      RECT -17.845 -68.895 -17.745 -63.535 ;
      RECT -17.845 -62.435 -17.745 -57.075 ;
      RECT -17.845 -55.975 -17.745 -50.615 ;
      RECT -17.845 -49.515 -17.745 -44.155 ;
      RECT -17.845 -43.055 -17.745 -37.695 ;
      RECT -17.845 -36.595 -17.745 -31.235 ;
      RECT -17.845 -30.135 -17.745 -24.775 ;
      RECT -17.845 -23.675 -17.745 -18.315 ;
      RECT -17.845 -17.215 -17.745 -11.855 ;
      RECT -17.845 -10.755 -17.745 -5.395 ;
      RECT -17.845 -4.295 -17.745 1.065 ;
      RECT -18.365 -101.195 -18.265 -95.835 ;
      RECT -18.365 -94.735 -18.265 -89.375 ;
      RECT -18.365 -88.275 -18.265 -82.915 ;
      RECT -18.365 -81.815 -18.265 -76.455 ;
      RECT -18.365 -75.355 -18.265 -69.995 ;
      RECT -18.365 -68.895 -18.265 -63.535 ;
      RECT -18.365 -62.435 -18.265 -57.075 ;
      RECT -18.365 -55.975 -18.265 -50.615 ;
      RECT -18.365 -49.515 -18.265 -44.155 ;
      RECT -18.365 -43.055 -18.265 -37.695 ;
      RECT -18.365 -36.595 -18.265 -31.235 ;
      RECT -18.365 -30.135 -18.265 -24.775 ;
      RECT -18.365 -23.675 -18.265 -18.315 ;
      RECT -18.365 -17.215 -18.265 -11.855 ;
      RECT -18.365 -10.755 -18.265 -5.395 ;
      RECT -18.365 -4.295 -18.265 1.065 ;
      RECT -19.145 -101.195 -19.045 -95.835 ;
      RECT -19.145 -94.735 -19.045 -89.375 ;
      RECT -19.145 -88.275 -19.045 -82.915 ;
      RECT -19.145 -81.815 -19.045 -76.455 ;
      RECT -19.145 -75.355 -19.045 -69.995 ;
      RECT -19.145 -68.895 -19.045 -63.535 ;
      RECT -19.145 -62.435 -19.045 -57.075 ;
      RECT -19.145 -55.975 -19.045 -50.615 ;
      RECT -19.145 -49.515 -19.045 -44.155 ;
      RECT -19.145 -43.055 -19.045 -37.695 ;
      RECT -19.145 -36.595 -19.045 -31.235 ;
      RECT -19.145 -30.135 -19.045 -24.775 ;
      RECT -19.145 -23.675 -19.045 -18.315 ;
      RECT -19.145 -17.215 -19.045 -11.855 ;
      RECT -19.145 -10.755 -19.045 -5.395 ;
      RECT -19.145 -4.295 -19.045 1.065 ;
      RECT -19.665 -101.195 -19.565 -95.835 ;
      RECT -19.665 -94.735 -19.565 -89.375 ;
      RECT -19.665 -88.275 -19.565 -82.915 ;
      RECT -19.665 -81.815 -19.565 -76.455 ;
      RECT -19.665 -75.355 -19.565 -69.995 ;
      RECT -19.665 -68.895 -19.565 -63.535 ;
      RECT -19.665 -62.435 -19.565 -57.075 ;
      RECT -19.665 -55.975 -19.565 -50.615 ;
      RECT -19.665 -49.515 -19.565 -44.155 ;
      RECT -19.665 -43.055 -19.565 -37.695 ;
      RECT -19.665 -36.595 -19.565 -31.235 ;
      RECT -19.665 -30.135 -19.565 -24.775 ;
      RECT -19.665 -23.675 -19.565 -18.315 ;
      RECT -19.665 -17.215 -19.565 -11.855 ;
      RECT -19.665 -10.755 -19.565 -5.395 ;
      RECT -19.665 -4.295 -19.565 1.065 ;
      RECT -20.445 -101.195 -20.345 -95.835 ;
      RECT -20.445 -94.735 -20.345 -89.375 ;
      RECT -20.445 -88.275 -20.345 -82.915 ;
      RECT -20.445 -81.815 -20.345 -76.455 ;
      RECT -20.445 -75.355 -20.345 -69.995 ;
      RECT -20.445 -68.895 -20.345 -63.535 ;
      RECT -20.445 -62.435 -20.345 -57.075 ;
      RECT -20.445 -55.975 -20.345 -50.615 ;
      RECT -20.445 -49.515 -20.345 -44.155 ;
      RECT -20.445 -43.055 -20.345 -37.695 ;
      RECT -20.445 -36.595 -20.345 -31.235 ;
      RECT -20.445 -30.135 -20.345 -24.775 ;
      RECT -20.445 -23.675 -20.345 -18.315 ;
      RECT -20.445 -17.215 -20.345 -11.855 ;
      RECT -20.445 -10.755 -20.345 -5.395 ;
      RECT -20.445 -4.295 -20.345 1.065 ;
      RECT -20.965 -101.195 -20.865 -95.835 ;
      RECT -20.965 -94.735 -20.865 -89.375 ;
      RECT -20.965 -88.275 -20.865 -82.915 ;
      RECT -20.965 -81.815 -20.865 -76.455 ;
      RECT -20.965 -75.355 -20.865 -69.995 ;
      RECT -20.965 -68.895 -20.865 -63.535 ;
      RECT -20.965 -62.435 -20.865 -57.075 ;
      RECT -20.965 -55.975 -20.865 -50.615 ;
      RECT -20.965 -49.515 -20.865 -44.155 ;
      RECT -20.965 -43.055 -20.865 -37.695 ;
      RECT -20.965 -36.595 -20.865 -31.235 ;
      RECT -20.965 -30.135 -20.865 -24.775 ;
      RECT -20.965 -23.675 -20.865 -18.315 ;
      RECT -20.965 -17.215 -20.865 -11.855 ;
      RECT -20.965 -10.755 -20.865 -5.395 ;
      RECT -20.965 -4.295 -20.865 1.065 ;
      RECT -21.745 -101.195 -21.645 -95.835 ;
      RECT -21.745 -94.735 -21.645 -89.375 ;
      RECT -21.745 -88.275 -21.645 -82.915 ;
      RECT -21.745 -81.815 -21.645 -76.455 ;
      RECT -21.745 -75.355 -21.645 -69.995 ;
      RECT -21.745 -68.895 -21.645 -63.535 ;
      RECT -21.745 -62.435 -21.645 -57.075 ;
      RECT -21.745 -55.975 -21.645 -50.615 ;
      RECT -21.745 -49.515 -21.645 -44.155 ;
      RECT -21.745 -43.055 -21.645 -37.695 ;
      RECT -21.745 -36.595 -21.645 -31.235 ;
      RECT -21.745 -30.135 -21.645 -24.775 ;
      RECT -21.745 -23.675 -21.645 -18.315 ;
      RECT -21.745 -17.215 -21.645 -11.855 ;
      RECT -21.745 -10.755 -21.645 -5.395 ;
      RECT -21.745 -4.295 -21.645 1.065 ;
      RECT -22.265 -101.195 -22.165 -95.835 ;
      RECT -22.265 -94.735 -22.165 -89.375 ;
      RECT -22.265 -88.275 -22.165 -82.915 ;
      RECT -22.265 -81.815 -22.165 -76.455 ;
      RECT -22.265 -75.355 -22.165 -69.995 ;
      RECT -22.265 -68.895 -22.165 -63.535 ;
      RECT -22.265 -62.435 -22.165 -57.075 ;
      RECT -22.265 -55.975 -22.165 -50.615 ;
      RECT -22.265 -49.515 -22.165 -44.155 ;
      RECT -22.265 -43.055 -22.165 -37.695 ;
      RECT -22.265 -36.595 -22.165 -31.235 ;
      RECT -22.265 -30.135 -22.165 -24.775 ;
      RECT -22.265 -23.675 -22.165 -18.315 ;
      RECT -22.265 -17.215 -22.165 -11.855 ;
      RECT -22.265 -10.755 -22.165 -5.395 ;
      RECT -22.265 -4.295 -22.165 1.065 ;
      RECT -23.045 -101.195 -22.945 -95.835 ;
      RECT -23.045 -94.735 -22.945 -89.375 ;
      RECT -23.045 -88.275 -22.945 -82.915 ;
      RECT -23.045 -81.815 -22.945 -76.455 ;
      RECT -23.045 -75.355 -22.945 -69.995 ;
      RECT -23.045 -68.895 -22.945 -63.535 ;
      RECT -23.045 -62.435 -22.945 -57.075 ;
      RECT -23.045 -55.975 -22.945 -50.615 ;
      RECT -23.045 -49.515 -22.945 -44.155 ;
      RECT -23.045 -43.055 -22.945 -37.695 ;
      RECT -23.045 -36.595 -22.945 -31.235 ;
      RECT -23.045 -30.135 -22.945 -24.775 ;
      RECT -23.045 -23.675 -22.945 -18.315 ;
      RECT -23.045 -17.215 -22.945 -11.855 ;
      RECT -23.045 -10.755 -22.945 -5.395 ;
      RECT -23.045 -4.295 -22.945 1.065 ;
      RECT -23.565 -101.195 -23.465 -95.835 ;
      RECT -23.565 -94.735 -23.465 -89.375 ;
      RECT -23.565 -88.275 -23.465 -82.915 ;
      RECT -23.565 -81.815 -23.465 -76.455 ;
      RECT -23.565 -75.355 -23.465 -69.995 ;
      RECT -23.565 -68.895 -23.465 -63.535 ;
      RECT -23.565 -62.435 -23.465 -57.075 ;
      RECT -23.565 -55.975 -23.465 -50.615 ;
      RECT -23.565 -49.515 -23.465 -44.155 ;
      RECT -23.565 -43.055 -23.465 -37.695 ;
      RECT -23.565 -36.595 -23.465 -31.235 ;
      RECT -23.565 -30.135 -23.465 -24.775 ;
      RECT -23.565 -23.675 -23.465 -18.315 ;
      RECT -23.565 -17.215 -23.465 -11.855 ;
      RECT -23.565 -10.755 -23.465 -5.395 ;
      RECT -23.565 -4.295 -23.465 1.065 ;
      RECT -24.345 -101.195 -24.245 -95.835 ;
      RECT -24.345 -94.735 -24.245 -89.375 ;
      RECT -24.345 -88.275 -24.245 -82.915 ;
      RECT -24.345 -81.815 -24.245 -76.455 ;
      RECT -24.345 -75.355 -24.245 -69.995 ;
      RECT -24.345 -68.895 -24.245 -63.535 ;
      RECT -24.345 -62.435 -24.245 -57.075 ;
      RECT -24.345 -55.975 -24.245 -50.615 ;
      RECT -24.345 -49.515 -24.245 -44.155 ;
      RECT -24.345 -43.055 -24.245 -37.695 ;
      RECT -24.345 -36.595 -24.245 -31.235 ;
      RECT -24.345 -30.135 -24.245 -24.775 ;
      RECT -24.345 -23.675 -24.245 -18.315 ;
      RECT -24.345 -17.215 -24.245 -11.855 ;
      RECT -24.345 -10.755 -24.245 -5.395 ;
      RECT -24.345 -4.295 -24.245 1.065 ;
      RECT -24.865 -101.195 -24.765 -95.835 ;
      RECT -24.865 -94.735 -24.765 -89.375 ;
      RECT -24.865 -88.275 -24.765 -82.915 ;
      RECT -24.865 -81.815 -24.765 -76.455 ;
      RECT -24.865 -75.355 -24.765 -69.995 ;
      RECT -24.865 -68.895 -24.765 -63.535 ;
      RECT -24.865 -62.435 -24.765 -57.075 ;
      RECT -24.865 -55.975 -24.765 -50.615 ;
      RECT -24.865 -49.515 -24.765 -44.155 ;
      RECT -24.865 -43.055 -24.765 -37.695 ;
      RECT -24.865 -36.595 -24.765 -31.235 ;
      RECT -24.865 -30.135 -24.765 -24.775 ;
      RECT -24.865 -23.675 -24.765 -18.315 ;
      RECT -24.865 -17.215 -24.765 -11.855 ;
      RECT -24.865 -10.755 -24.765 -5.395 ;
      RECT -24.865 -4.295 -24.765 1.065 ;
      RECT -25.645 -101.195 -25.545 -95.835 ;
      RECT -25.645 -94.735 -25.545 -89.375 ;
      RECT -25.645 -88.275 -25.545 -82.915 ;
      RECT -25.645 -81.815 -25.545 -76.455 ;
      RECT -25.645 -75.355 -25.545 -69.995 ;
      RECT -25.645 -68.895 -25.545 -63.535 ;
      RECT -25.645 -62.435 -25.545 -57.075 ;
      RECT -25.645 -55.975 -25.545 -50.615 ;
      RECT -25.645 -49.515 -25.545 -44.155 ;
      RECT -25.645 -43.055 -25.545 -37.695 ;
      RECT -25.645 -36.595 -25.545 -31.235 ;
      RECT -25.645 -30.135 -25.545 -24.775 ;
      RECT -25.645 -23.675 -25.545 -18.315 ;
      RECT -25.645 -17.215 -25.545 -11.855 ;
      RECT -25.645 -10.755 -25.545 -5.395 ;
      RECT -25.645 -4.295 -25.545 1.065 ;
      RECT -26.165 -101.195 -26.065 -95.835 ;
      RECT -26.165 -94.735 -26.065 -89.375 ;
      RECT -26.165 -88.275 -26.065 -82.915 ;
      RECT -26.165 -81.815 -26.065 -76.455 ;
      RECT -26.165 -75.355 -26.065 -69.995 ;
      RECT -26.165 -68.895 -26.065 -63.535 ;
      RECT -26.165 -62.435 -26.065 -57.075 ;
      RECT -26.165 -55.975 -26.065 -50.615 ;
      RECT -26.165 -49.515 -26.065 -44.155 ;
      RECT -26.165 -43.055 -26.065 -37.695 ;
      RECT -26.165 -36.595 -26.065 -31.235 ;
      RECT -26.165 -30.135 -26.065 -24.775 ;
      RECT -26.165 -23.675 -26.065 -18.315 ;
      RECT -26.165 -17.215 -26.065 -11.855 ;
      RECT -26.165 -10.755 -26.065 -5.395 ;
      RECT -26.165 -4.295 -26.065 1.065 ;
      RECT -26.945 -101.195 -26.845 -95.835 ;
      RECT -26.945 -94.735 -26.845 -89.375 ;
      RECT -26.945 -88.275 -26.845 -82.915 ;
      RECT -26.945 -81.815 -26.845 -76.455 ;
      RECT -26.945 -75.355 -26.845 -69.995 ;
      RECT -26.945 -68.895 -26.845 -63.535 ;
      RECT -26.945 -62.435 -26.845 -57.075 ;
      RECT -26.945 -55.975 -26.845 -50.615 ;
      RECT -26.945 -49.515 -26.845 -44.155 ;
      RECT -26.945 -43.055 -26.845 -37.695 ;
      RECT -26.945 -36.595 -26.845 -31.235 ;
      RECT -26.945 -30.135 -26.845 -24.775 ;
      RECT -26.945 -23.675 -26.845 -18.315 ;
      RECT -26.945 -17.215 -26.845 -11.855 ;
      RECT -26.945 -10.755 -26.845 -5.395 ;
      RECT -26.945 -4.295 -26.845 1.065 ;
      RECT -27.465 -101.195 -27.365 -95.835 ;
      RECT -27.465 -94.735 -27.365 -89.375 ;
      RECT -27.465 -88.275 -27.365 -82.915 ;
      RECT -27.465 -81.815 -27.365 -76.455 ;
      RECT -27.465 -75.355 -27.365 -69.995 ;
      RECT -27.465 -68.895 -27.365 -63.535 ;
      RECT -27.465 -62.435 -27.365 -57.075 ;
      RECT -27.465 -55.975 -27.365 -50.615 ;
      RECT -27.465 -49.515 -27.365 -44.155 ;
      RECT -27.465 -43.055 -27.365 -37.695 ;
      RECT -27.465 -36.595 -27.365 -31.235 ;
      RECT -27.465 -30.135 -27.365 -24.775 ;
      RECT -27.465 -23.675 -27.365 -18.315 ;
      RECT -27.465 -17.215 -27.365 -11.855 ;
      RECT -27.465 -10.755 -27.365 -5.395 ;
      RECT -27.465 -4.295 -27.365 1.065 ;
      RECT -28.245 -101.195 -28.145 -95.835 ;
      RECT -28.245 -94.735 -28.145 -89.375 ;
      RECT -28.245 -88.275 -28.145 -82.915 ;
      RECT -28.245 -81.815 -28.145 -76.455 ;
      RECT -28.245 -75.355 -28.145 -69.995 ;
      RECT -28.245 -68.895 -28.145 -63.535 ;
      RECT -28.245 -62.435 -28.145 -57.075 ;
      RECT -28.245 -55.975 -28.145 -50.615 ;
      RECT -28.245 -49.515 -28.145 -44.155 ;
      RECT -28.245 -43.055 -28.145 -37.695 ;
      RECT -28.245 -36.595 -28.145 -31.235 ;
      RECT -28.245 -30.135 -28.145 -24.775 ;
      RECT -28.245 -23.675 -28.145 -18.315 ;
      RECT -28.245 -17.215 -28.145 -11.855 ;
      RECT -28.245 -10.755 -28.145 -5.395 ;
      RECT -28.245 -4.295 -28.145 1.065 ;
      RECT -28.765 -101.195 -28.665 -95.835 ;
      RECT -28.765 -94.735 -28.665 -89.375 ;
      RECT -28.765 -88.275 -28.665 -82.915 ;
      RECT -28.765 -81.815 -28.665 -76.455 ;
      RECT -28.765 -75.355 -28.665 -69.995 ;
      RECT -28.765 -68.895 -28.665 -63.535 ;
      RECT -28.765 -62.435 -28.665 -57.075 ;
      RECT -28.765 -55.975 -28.665 -50.615 ;
      RECT -28.765 -49.515 -28.665 -44.155 ;
      RECT -28.765 -43.055 -28.665 -37.695 ;
      RECT -28.765 -36.595 -28.665 -31.235 ;
      RECT -28.765 -30.135 -28.665 -24.775 ;
      RECT -28.765 -23.675 -28.665 -18.315 ;
      RECT -28.765 -17.215 -28.665 -11.855 ;
      RECT -28.765 -10.755 -28.665 -5.395 ;
      RECT -28.765 -4.295 -28.665 1.065 ;
      RECT -29.545 -101.195 -29.445 -95.835 ;
      RECT -29.545 -94.735 -29.445 -89.375 ;
      RECT -29.545 -88.275 -29.445 -82.915 ;
      RECT -29.545 -81.815 -29.445 -76.455 ;
      RECT -29.545 -75.355 -29.445 -69.995 ;
      RECT -29.545 -68.895 -29.445 -63.535 ;
      RECT -29.545 -62.435 -29.445 -57.075 ;
      RECT -29.545 -55.975 -29.445 -50.615 ;
      RECT -29.545 -49.515 -29.445 -44.155 ;
      RECT -29.545 -43.055 -29.445 -37.695 ;
      RECT -29.545 -36.595 -29.445 -31.235 ;
      RECT -29.545 -30.135 -29.445 -24.775 ;
      RECT -29.545 -23.675 -29.445 -18.315 ;
      RECT -29.545 -17.215 -29.445 -11.855 ;
      RECT -29.545 -10.755 -29.445 -5.395 ;
      RECT -29.545 -4.295 -29.445 1.065 ;
      RECT -30.065 -101.195 -29.965 -95.835 ;
      RECT -30.065 -94.735 -29.965 -89.375 ;
      RECT -30.065 -88.275 -29.965 -82.915 ;
      RECT -30.065 -81.815 -29.965 -76.455 ;
      RECT -30.065 -75.355 -29.965 -69.995 ;
      RECT -30.065 -68.895 -29.965 -63.535 ;
      RECT -30.065 -62.435 -29.965 -57.075 ;
      RECT -30.065 -55.975 -29.965 -50.615 ;
      RECT -30.065 -49.515 -29.965 -44.155 ;
      RECT -30.065 -43.055 -29.965 -37.695 ;
      RECT -30.065 -36.595 -29.965 -31.235 ;
      RECT -30.065 -30.135 -29.965 -24.775 ;
      RECT -30.065 -23.675 -29.965 -18.315 ;
      RECT -30.065 -17.215 -29.965 -11.855 ;
      RECT -30.065 -10.755 -29.965 -5.395 ;
      RECT -30.065 -4.295 -29.965 1.065 ;
      RECT -30.845 -101.195 -30.745 -95.835 ;
      RECT -30.845 -94.735 -30.745 -89.375 ;
      RECT -30.845 -88.275 -30.745 -82.915 ;
      RECT -30.845 -81.815 -30.745 -76.455 ;
      RECT -30.845 -75.355 -30.745 -69.995 ;
      RECT -30.845 -68.895 -30.745 -63.535 ;
      RECT -30.845 -62.435 -30.745 -57.075 ;
      RECT -30.845 -55.975 -30.745 -50.615 ;
      RECT -30.845 -49.515 -30.745 -44.155 ;
      RECT -30.845 -43.055 -30.745 -37.695 ;
      RECT -30.845 -36.595 -30.745 -31.235 ;
      RECT -30.845 -30.135 -30.745 -24.775 ;
      RECT -30.845 -23.675 -30.745 -18.315 ;
      RECT -30.845 -17.215 -30.745 -11.855 ;
      RECT -30.845 -10.755 -30.745 -5.395 ;
      RECT -30.845 -4.295 -30.745 1.065 ;
      RECT -31.365 -101.195 -31.265 -95.835 ;
      RECT -31.365 -94.735 -31.265 -89.375 ;
      RECT -31.365 -88.275 -31.265 -82.915 ;
      RECT -31.365 -81.815 -31.265 -76.455 ;
      RECT -31.365 -75.355 -31.265 -69.995 ;
      RECT -31.365 -68.895 -31.265 -63.535 ;
      RECT -31.365 -62.435 -31.265 -57.075 ;
      RECT -31.365 -55.975 -31.265 -50.615 ;
      RECT -31.365 -49.515 -31.265 -44.155 ;
      RECT -31.365 -43.055 -31.265 -37.695 ;
      RECT -31.365 -36.595 -31.265 -31.235 ;
      RECT -31.365 -30.135 -31.265 -24.775 ;
      RECT -31.365 -23.675 -31.265 -18.315 ;
      RECT -31.365 -17.215 -31.265 -11.855 ;
      RECT -31.365 -10.755 -31.265 -5.395 ;
      RECT -31.365 -4.295 -31.265 1.065 ;
      RECT -37.505 -120.605 -36.505 5.645 ;
      RECT -39.505 -115.155 -38.505 9.895 ;
  END
END sram_1kb_64x128x32

END LIBRARY
